// Benchmark "amba5c5y_cert" written by ABC on Sat Jul 29 16:29:14 2017

module amba5c5y_cert ( 
    n55, reg_controllable_hgrant2_out, reg_controllable_hmaster1_out,
    reg_controllable_hgrant3_out, next_env_fair_out,
    reg_controllable_hmaster2_out, reg_controllable_hgrant4_out,
    reg_stateG3_0_out, reg_stateG3_1_out, reg_controllable_locked_out,
    reg_controllable_ndecide_out, reg_stateG3_2_out,
    reg_controllable_busreq_out, reg_i_hlock4_out,
    reg_controllable_nstart_out, reg_i_hbusreq0_out, reg_i_hlock3_out,
    reg_stateG2_out, reg_stateG10_1_out, reg_i_hbusreq1_out,
    reg_i_hlock2_out, reg_controllable_hmastlock_out, reg_stateG10_2_out,
    reg_controllable_nhgrant0_out, reg_i_hbusreq2_out, reg_stateA1_out,
    reg_i_hlock1_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , next_sys_fair<0>_out , next_sys_fair<1>_out ,
    next_sys_fair<2>_out , next_sys_fair<3>_out , reg_stateG10_3_out,
    reg_i_hbusreq3_out, reg_i_hlock0_out, reg_i_hready_out,
    env_safe_err_happened_out, reg_stateG10_4_out, reg_i_hbusreq4_out,
    reg_controllable_hgrant1_out, reg_controllable_hmaster0_out, i_hlock0,
    i_hlock1, i_hlock2, i_hlock3, i_hlock4, i_hready, i_hburst1, i_hburst0,
    i_hbusreq0, i_hbusreq1, i_hbusreq2, i_hbusreq3, i_hbusreq4,
    controllable_nhgrant0, controllable_hgrant1, controllable_locked,
    controllable_nstart, controllable_hgrant2, controllable_hgrant3,
    controllable_hgrant4, controllable_busreq, controllable_ndecide,
    controllable_hmaster2, controllable_hmaster1, controllable_hmaster0,
    controllable_hmastlock,
    inductivity_check   );
  input  n55, reg_controllable_hgrant2_out,
    reg_controllable_hmaster1_out, reg_controllable_hgrant3_out,
    next_env_fair_out, reg_controllable_hmaster2_out,
    reg_controllable_hgrant4_out, reg_stateG3_0_out, reg_stateG3_1_out,
    reg_controllable_locked_out, reg_controllable_ndecide_out,
    reg_stateG3_2_out, reg_controllable_busreq_out, reg_i_hlock4_out,
    reg_controllable_nstart_out, reg_i_hbusreq0_out, reg_i_hlock3_out,
    reg_stateG2_out, reg_stateG10_1_out, reg_i_hbusreq1_out,
    reg_i_hlock2_out, reg_controllable_hmastlock_out, reg_stateG10_2_out,
    reg_controllable_nhgrant0_out, reg_i_hbusreq2_out, reg_stateA1_out,
    reg_i_hlock1_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , next_sys_fair<0>_out , next_sys_fair<1>_out ,
    next_sys_fair<2>_out , next_sys_fair<3>_out , reg_stateG10_3_out,
    reg_i_hbusreq3_out, reg_i_hlock0_out, reg_i_hready_out,
    env_safe_err_happened_out, reg_stateG10_4_out, reg_i_hbusreq4_out,
    reg_controllable_hgrant1_out, reg_controllable_hmaster0_out, i_hlock0,
    i_hlock1, i_hlock2, i_hlock3, i_hlock4, i_hready, i_hburst1, i_hburst0,
    i_hbusreq0, i_hbusreq1, i_hbusreq2, i_hbusreq3, i_hbusreq4,
    controllable_nhgrant0, controllable_hgrant1, controllable_locked,
    controllable_nstart, controllable_hgrant2, controllable_hgrant3,
    controllable_hgrant4, controllable_busreq, controllable_ndecide,
    controllable_hmaster2, controllable_hmaster1, controllable_hmaster0,
    controllable_hmastlock;
  output inductivity_check ;
  wire n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
    n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
    n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
    n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
    n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
    n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
    n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
    n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
    n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
    n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
    n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
    n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
    n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
    n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
    n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
    n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
    n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
    n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
    n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
    n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
    n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
    n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
    n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
    n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
    n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
    n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
    n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
    n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
    n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
    n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
    n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
    n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
    n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
    n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
    n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
    n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
    n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
    n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
    n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
    n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
    n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
    n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
    n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
    n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
    n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
    n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
    n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
    n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
    n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
    n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
    n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
    n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
    n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
    n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
    n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
    n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
    n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
    n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
    n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
    n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
    n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
    n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
    n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
    n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
    n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
    n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
    n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
    n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
    n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
    n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
    n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
    n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
    n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
    n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
    n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
    n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
    n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
    n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
    n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
    n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
    n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
    n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
    n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
    n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
    n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
    n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
    n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
    n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
    n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
    n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
    n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
    n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
    n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
    n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
    n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
    n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
    n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
    n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
    n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
    n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
    n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
    n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
    n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
    n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
    n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
    n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
    n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
    n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
    n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
    n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
    n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
    n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
    n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
    n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
    n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
    n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
    n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
    n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
    n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
    n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
    n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
    n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
    n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
    n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
    n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
    n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
    n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
    n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
    n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
    n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
    n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
    n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
    n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
    n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
    n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
    n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
    n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
    n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
    n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
    n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
    n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
    n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
    n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
    n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
    n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
    n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
    n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
    n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
    n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
    n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
    n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
    n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
    n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
    n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
    n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
    n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
    n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
    n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
    n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
    n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
    n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
    n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
    n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
    n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
    n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
    n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
    n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
    n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
    n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
    n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
    n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
    n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
    n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
    n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
    n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
    n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
    n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
    n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
    n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
    n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
    n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
    n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
    n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
    n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
    n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
    n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
    n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
    n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
    n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
    n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
    n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
    n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
    n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
    n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
    n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
    n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
    n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
    n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
    n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
    n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
    n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
    n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
    n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
    n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
    n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
    n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
    n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
    n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
    n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
    n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
    n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
    n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
    n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
    n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
    n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
    n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
    n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
    n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
    n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
    n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
    n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
    n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
    n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
    n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
    n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
    n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
    n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
    n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
    n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
    n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
    n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
    n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
    n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
    n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
    n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
    n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
    n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
    n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
    n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
    n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
    n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
    n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
    n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
    n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
    n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
    n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
    n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
    n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
    n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
    n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
    n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
    n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
    n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
    n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
    n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
    n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
    n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
    n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
    n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
    n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
    n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
    n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
    n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
    n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
    n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
    n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
    n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
    n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
    n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
    n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
    n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
    n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
    n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
    n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
    n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
    n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
    n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
    n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
    n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
    n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
    n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
    n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
    n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
    n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
    n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
    n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
    n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
    n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
    n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
    n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
    n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
    n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
    n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
    n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
    n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
    n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
    n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
    n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
    n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
    n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
    n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
    n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
    n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
    n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
    n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
    n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
    n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
    n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
    n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
    n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
    n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
    n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
    n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
    n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
    n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
    n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
    n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
    n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
    n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
    n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
    n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
    n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
    n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
    n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
    n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
    n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
    n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
    n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
    n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
    n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
    n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
    n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
    n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
    n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
    n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
    n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
    n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
    n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
    n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
    n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
    n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
    n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
    n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
    n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
    n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
    n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
    n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
    n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
    n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
    n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
    n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
    n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
    n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
    n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
    n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
    n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
    n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
    n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
    n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
    n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
    n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
    n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
    n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
    n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
    n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
    n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
    n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
    n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
    n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
    n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
    n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
    n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
    n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
    n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
    n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
    n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
    n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
    n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
    n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
    n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
    n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
    n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
    n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
    n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
    n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
    n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
    n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
    n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
    n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
    n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
    n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
    n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
    n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
    n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
    n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
    n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
    n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
    n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
    n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
    n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
    n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
    n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
    n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
    n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
    n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
    n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
    n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
    n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
    n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
    n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
    n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
    n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
    n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
    n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
    n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
    n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
    n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
    n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
    n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
    n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
    n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
    n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
    n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
    n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
    n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
    n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
    n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
    n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
    n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
    n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
    n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
    n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
    n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
    n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
    n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
    n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
    n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
    n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
    n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
    n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
    n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
    n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
    n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
    n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
    n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
    n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
    n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
    n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
    n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
    n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
    n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
    n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
    n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
    n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
    n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
    n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
    n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
    n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
    n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
    n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
    n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
    n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
    n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
    n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
    n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
    n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
    n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
    n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
    n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
    n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
    n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
    n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
    n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
    n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
    n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
    n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
    n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
    n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
    n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
    n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
    n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
    n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
    n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
    n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
    n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
    n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
    n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
    n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
    n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
    n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
    n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
    n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
    n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
    n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
    n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
    n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
    n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
    n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
    n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
    n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
    n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
    n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
    n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
    n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
    n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
    n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
    n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
    n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
    n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
    n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
    n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
    n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
    n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
    n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
    n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
    n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
    n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
    n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
    n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
    n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
    n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
    n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
    n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
    n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
    n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
    n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
    n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
    n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
    n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
    n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
    n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
    n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
    n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
    n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
    n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
    n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
    n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
    n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
    n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
    n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
    n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
    n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
    n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
    n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
    n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
    n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
    n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
    n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
    n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
    n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
    n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
    n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
    n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
    n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
    n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
    n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
    n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
    n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
    n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
    n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
    n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
    n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
    n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
    n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
    n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
    n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
    n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
    n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
    n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
    n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
    n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
    n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
    n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
    n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
    n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
    n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
    n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
    n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
    n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
    n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
    n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
    n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
    n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
    n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
    n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
    n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
    n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
    n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
    n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
    n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
    n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
    n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
    n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
    n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
    n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
    n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
    n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
    n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
    n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
    n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
    n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
    n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
    n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
    n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
    n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
    n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
    n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
    n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
    n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
    n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
    n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
    n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
    n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
    n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
    n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
    n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
    n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
    n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
    n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
    n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
    n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
    n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
    n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
    n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
    n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
    n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
    n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
    n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016,
    n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
    n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
    n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
    n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
    n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
    n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
    n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
    n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088,
    n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
    n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
    n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
    n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
    n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
    n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
    n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
    n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160,
    n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
    n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
    n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
    n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
    n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
    n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
    n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
    n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
    n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
    n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
    n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
    n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
    n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
    n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
    n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
    n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
    n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
    n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
    n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
    n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
    n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
    n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
    n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
    n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
    n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
    n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
    n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
    n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
    n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
    n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
    n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
    n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
    n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
    n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
    n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
    n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
    n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
    n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
    n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
    n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
    n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
    n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
    n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
    n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
    n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
    n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
    n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
    n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
    n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
    n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
    n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
    n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997,
    n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
    n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
    n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
    n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
    n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
    n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
    n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
    n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069,
    n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
    n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
    n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
    n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
    n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
    n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
    n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
    n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
    n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
    n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
    n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
    n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
    n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204,
    n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213,
    n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
    n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
    n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
    n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
    n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
    n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
    n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
    n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
    n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357,
    n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
    n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
    n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
    n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
    n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
    n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
    n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
    n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501,
    n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
    n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
    n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
    n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573,
    n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
    n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
    n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
    n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645,
    n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
    n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
    n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
    n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
    n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
    n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708,
    n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
    n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
    n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
    n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
    n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
    n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
    n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
    n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
    n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
    n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
    n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852,
    n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861,
    n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
    n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
    n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
    n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
    n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
    n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
    n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924,
    n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933,
    n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
    n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
    n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
    n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996,
    n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005,
    n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
    n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
    n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
    n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
    n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
    n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
    n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
    n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077,
    n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
    n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
    n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
    n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
    n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
    n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
    n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
    n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
    n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
    n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
    n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
    n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212,
    n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221,
    n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
    n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
    n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
    n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
    n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
    n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
    n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284,
    n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
    n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
    n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
    n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
    n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
    n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
    n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
    n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356,
    n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365,
    n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
    n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
    n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
    n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428,
    n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
    n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
    n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
    n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
    n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
    n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
    n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
    n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509,
    n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
    n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
    n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
    n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
    n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572,
    n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581,
    n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
    n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
    n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
    n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
    n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
    n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
    n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644,
    n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653,
    n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
    n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
    n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
    n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
    n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
    n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
    n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716,
    n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
    n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
    n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
    n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
    n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
    n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
    n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
    n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860,
    n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869,
    n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
    n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
    n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
    n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
    n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
    n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
    n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
    n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
    n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
    n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
    n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
    n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
    n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013,
    n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
    n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
    n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
    n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
    n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
    n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
    n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
    n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085,
    n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
    n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
    n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
    n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
    n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
    n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
    n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
    n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157,
    n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
    n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
    n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
    n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
    n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
    n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
    n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
    n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229,
    n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
    n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
    n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
    n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
    n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
    n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
    n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301,
    n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
    n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
    n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
    n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
    n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
    n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
    n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
    n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373,
    n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
    n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
    n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
    n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
    n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
    n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
    n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445,
    n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
    n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
    n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
    n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
    n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517,
    n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
    n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
    n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
    n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
    n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589,
    n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
    n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
    n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
    n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661,
    n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
    n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
    n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
    n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
    n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
    n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
    n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733,
    n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
    n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
    n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
    n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
    n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805,
    n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
    n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
    n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
    n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
    n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
    n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
    n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
    n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877,
    n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
    n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
    n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
    n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
    n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
    n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
    n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949,
    n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
    n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
    n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
    n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
    n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
    n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
    n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
    n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021,
    n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
    n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039,
    n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
    n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
    n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
    n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
    n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
    n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
    n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
    n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
    n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
    n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
    n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
    n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165,
    n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
    n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
    n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
    n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237,
    n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
    n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264,
    n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
    n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
    n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
    n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
    n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309,
    n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
    n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
    n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336,
    n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
    n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
    n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
    n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
    n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381,
    n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
    n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
    n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
    n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453,
    n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471,
    n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
    n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
    n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
    n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
    n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
    n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525,
    n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
    n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
    n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
    n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
    n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
    n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
    n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
    n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597,
    n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
    n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615,
    n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
    n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
    n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
    n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
    n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
    n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669,
    n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
    n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
    n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
    n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
    n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
    n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
    n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
    n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
    n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
    n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
    n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
    n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
    n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
    n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813,
    n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
    n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
    n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
    n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
    n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
    n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
    n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885,
    n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
    n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
    n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
    n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
    n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
    n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
    n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957,
    n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
    n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
    n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
    n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
    n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
    n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
    n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
    n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029,
    n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
    n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
    n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
    n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
    n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
    n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
    n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101,
    n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
    n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
    n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
    n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
    n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
    n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
    n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173,
    n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
    n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
    n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
    n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245,
    n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
    n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263,
    n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
    n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
    n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
    n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
    n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
    n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317,
    n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
    n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
    n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
    n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
    n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
    n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
    n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
    n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389,
    n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
    n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407,
    n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
    n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
    n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
    n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
    n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
    n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
    n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
    n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
    n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
    n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
    n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
    n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
    n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
    n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
    n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
    n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
    n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
    n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
    n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
    n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
    n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605,
    n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
    n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623,
    n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
    n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
    n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
    n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
    n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
    n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677,
    n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
    n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695,
    n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
    n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
    n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
    n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
    n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
    n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749,
    n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
    n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767,
    n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
    n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
    n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
    n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
    n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
    n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821,
    n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
    n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839,
    n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
    n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
    n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
    n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
    n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
    n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893,
    n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
    n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
    n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
    n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
    n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965,
    n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
    n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
    n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
    n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
    n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037,
    n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
    n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
    n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
    n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
    n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
    n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
    n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109,
    n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
    n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
    n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
    n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
    n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
    n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
    n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
    n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181,
    n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
    n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
    n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
    n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
    n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
    n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
    n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
    n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253,
    n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
    n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
    n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
    n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
    n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
    n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
    n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
    n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325,
    n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
    n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
    n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
    n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
    n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
    n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
    n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
    n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397,
    n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
    n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
    n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
    n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
    n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
    n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
    n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
    n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469,
    n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
    n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
    n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
    n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
    n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
    n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
    n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
    n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541,
    n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
    n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
    n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
    n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
    n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
    n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
    n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
    n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613,
    n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
    n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
    n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
    n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
    n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
    n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
    n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685,
    n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
    n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
    n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
    n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
    n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
    n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
    n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757,
    n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
    n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
    n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
    n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
    n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
    n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
    n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
    n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829,
    n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
    n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
    n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856,
    n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
    n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
    n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
    n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892,
    n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901,
    n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
    n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
    n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928,
    n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
    n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
    n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
    n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964,
    n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973,
    n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
    n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
    n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000,
    n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
    n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
    n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
    n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036,
    n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045,
    n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
    n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
    n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
    n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
    n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
    n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
    n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
    n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117,
    n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
    n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
    n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
    n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
    n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
    n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
    n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180,
    n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189,
    n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
    n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
    n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
    n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
    n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
    n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
    n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
    n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261,
    n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
    n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
    n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
    n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
    n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
    n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324,
    n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
    n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
    n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
    n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
    n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
    n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
    n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
    n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405,
    n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
    n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
    n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
    n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
    n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
    n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
    n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468,
    n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477,
    n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
    n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
    n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
    n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
    n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
    n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
    n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
    n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549,
    n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
    n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
    n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
    n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
    n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
    n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
    n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621,
    n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
    n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
    n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
    n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
    n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
    n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693,
    n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
    n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
    n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720,
    n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
    n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
    n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
    n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756,
    n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765,
    n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
    n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
    n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
    n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
    n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837,
    n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
    n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
    n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
    n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900,
    n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909,
    n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
    n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
    n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
    n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
    n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
    n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
    n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972,
    n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981,
    n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
    n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
    n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008,
    n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
    n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
    n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
    n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044,
    n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053,
    n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
    n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080,
    n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
    n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
    n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
    n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116,
    n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125,
    n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143,
    n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
    n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
    n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
    n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188,
    n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197,
    n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
    n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
    n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
    n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260,
    n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269,
    n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
    n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296,
    n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
    n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
    n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
    n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332,
    n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341,
    n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
    n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359,
    n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368,
    n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
    n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
    n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
    n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404,
    n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413,
    n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
    n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431,
    n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
    n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
    n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
    n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
    n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476,
    n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485,
    n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
    n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
    n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512,
    n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
    n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
    n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
    n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548,
    n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557,
    n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
    n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
    n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584,
    n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
    n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
    n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629,
    n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
    n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
    n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
    n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
    n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692,
    n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701,
    n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
    n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719,
    n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728,
    n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
    n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
    n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
    n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764,
    n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773,
    n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
    n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791,
    n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800,
    n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
    n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
    n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
    n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836,
    n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845,
    n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
    n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863,
    n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
    n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
    n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
    n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
    n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908,
    n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917,
    n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
    n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935,
    n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
    n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980,
    n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989,
    n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
    n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007,
    n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
    n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
    n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
    n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
    n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052,
    n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061,
    n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
    n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079,
    n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
    n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
    n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
    n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133,
    n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151,
    n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
    n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
    n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196,
    n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205,
    n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
    n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223,
    n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
    n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
    n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
    n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
    n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268,
    n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277,
    n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
    n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
    n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
    n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
    n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
    n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
    n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340,
    n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349,
    n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
    n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367,
    n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
    n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
    n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
    n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
    n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412,
    n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421,
    n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
    n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439,
    n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
    n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
    n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
    n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
    n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484,
    n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493,
    n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
    n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511,
    n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
    n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
    n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
    n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556,
    n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565,
    n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
    n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583,
    n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
    n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
    n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
    n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
    n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628,
    n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637,
    n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
    n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
    n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
    n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
    n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
    n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
    n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709,
    n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
    n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
    n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
    n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
    n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
    n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
    n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772,
    n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781,
    n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
    n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799,
    n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
    n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
    n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
    n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
    n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844,
    n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853,
    n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
    n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871,
    n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
    n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
    n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
    n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
    n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916,
    n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925,
    n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
    n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
    n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
    n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
    n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
    n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
    n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997,
    n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
    n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
    n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
    n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
    n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
    n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
    n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
    n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
    n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
    n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
    n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
    n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
    n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
    n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
    n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204,
    n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
    n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
    n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276,
    n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285,
    n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
    n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
    n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
    n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
    n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348,
    n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
    n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
    n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
    n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420,
    n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
    n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
    n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
    n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483,
    n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492,
    n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501,
    n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
    n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519,
    n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
    n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
    n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
    n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
    n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564,
    n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573,
    n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
    n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591,
    n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
    n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
    n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
    n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
    n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636,
    n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645,
    n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
    n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663,
    n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
    n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
    n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
    n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699,
    n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708,
    n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717,
    n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
    n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735,
    n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
    n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
    n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
    n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771,
    n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780,
    n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789,
    n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
    n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
    n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
    n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
    n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
    n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
    n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852,
    n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861,
    n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
    n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879,
    n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
    n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
    n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
    n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
    n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924,
    n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933,
    n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
    n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951,
    n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
    n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
    n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
    n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
    n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996,
    n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005,
    n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
    n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
    n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
    n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
    n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
    n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
    n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068,
    n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077,
    n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
    n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
    n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
    n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
    n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
    n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
    n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140,
    n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149,
    n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
    n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167,
    n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
    n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
    n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
    n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
    n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212,
    n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221,
    n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
    n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239,
    n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
    n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
    n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
    n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
    n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284,
    n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293,
    n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
    n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
    n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
    n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
    n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
    n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
    n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356,
    n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365,
    n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
    n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383,
    n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
    n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
    n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
    n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
    n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428,
    n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437,
    n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
    n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
    n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
    n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
    n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
    n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
    n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500,
    n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509,
    n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
    n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527,
    n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
    n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
    n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
    n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
    n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572,
    n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581,
    n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
    n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
    n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
    n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
    n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
    n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
    n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644,
    n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653,
    n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
    n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671,
    n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
    n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
    n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
    n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
    n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
    n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725,
    n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
    n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743,
    n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
    n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
    n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
    n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788,
    n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797,
    n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
    n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815,
    n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
    n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
    n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
    n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
    n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860,
    n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869,
    n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
    n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887,
    n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
    n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
    n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
    n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
    n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932,
    n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941,
    n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
    n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
    n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
    n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
    n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
    n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
    n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004,
    n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013,
    n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
    n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
    n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
    n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
    n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
    n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
    n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085,
    n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
    n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
    n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
    n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
    n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
    n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148,
    n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157,
    n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
    n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
    n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
    n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
    n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
    n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
    n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220,
    n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229,
    n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
    n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
    n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
    n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
    n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
    n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
    n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301,
    n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
    n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
    n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
    n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
    n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373,
    n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
    n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
    n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
    n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
    n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
    n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445,
    n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
    n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
    n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
    n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
    n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
    n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508,
    n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517,
    n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
    n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
    n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
    n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
    n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
    n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
    n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580,
    n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589,
    n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
    n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607,
    n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
    n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
    n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
    n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652,
    n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661,
    n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
    n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679,
    n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
    n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
    n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
    n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
    n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
    n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733,
    n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
    n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751,
    n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
    n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
    n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
    n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
    n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796,
    n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805,
    n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
    n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823,
    n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
    n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
    n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
    n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
    n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868,
    n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877,
    n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
    n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895,
    n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
    n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
    n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949,
    n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
    n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967,
    n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
    n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
    n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
    n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
    n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021,
    n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
    n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
    n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
    n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
    n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
    n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
    n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093,
    n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102,
    n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
    n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
    n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
    n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
    n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
    n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156,
    n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165,
    n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174,
    n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183,
    n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
    n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
    n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
    n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
    n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228,
    n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237,
    n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246,
    n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255,
    n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
    n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
    n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
    n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
    n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300,
    n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309,
    n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318,
    n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327,
    n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
    n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
    n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
    n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
    n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
    n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381,
    n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390,
    n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
    n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
    n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
    n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
    n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
    n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444,
    n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453,
    n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462,
    n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
    n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
    n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
    n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
    n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525,
    n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
    n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
    n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
    n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
    n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
    n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588,
    n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597,
    n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606,
    n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615,
    n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
    n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
    n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
    n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
    n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660,
    n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669,
    n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
    n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687,
    n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
    n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
    n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
    n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
    n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732,
    n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741,
    n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
    n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759,
    n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
    n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
    n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
    n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
    n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804,
    n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813,
    n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
    n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831,
    n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
    n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
    n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
    n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
    n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876,
    n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885,
    n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903,
    n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
    n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
    n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
    n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
    n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948,
    n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957,
    n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
    n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975,
    n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
    n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
    n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
    n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
    n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020,
    n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029,
    n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047,
    n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
    n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
    n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
    n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
    n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092,
    n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101,
    n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
    n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119,
    n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
    n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
    n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
    n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173,
    n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
    n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191,
    n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
    n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
    n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
    n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
    n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
    n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245,
    n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
    n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263,
    n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
    n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
    n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
    n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
    n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
    n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317,
    n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
    n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335,
    n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
    n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
    n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
    n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
    n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380,
    n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389,
    n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
    n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407,
    n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
    n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
    n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
    n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
    n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452,
    n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461,
    n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
    n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479,
    n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488,
    n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
    n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
    n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
    n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524,
    n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533,
    n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
    n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551,
    n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560,
    n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
    n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
    n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596,
    n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605,
    n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623,
    n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
    n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
    n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
    n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668,
    n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677,
    n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
    n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695,
    n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704,
    n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
    n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
    n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
    n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740,
    n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749,
    n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
    n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767,
    n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
    n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
    n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
    n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
    n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812,
    n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821,
    n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
    n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839,
    n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848,
    n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
    n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
    n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
    n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884,
    n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893,
    n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
    n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911,
    n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920,
    n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
    n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
    n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
    n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956,
    n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965,
    n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
    n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983,
    n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992,
    n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
    n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
    n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
    n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028,
    n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037,
    n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
    n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055,
    n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
    n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
    n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
    n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
    n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100,
    n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109,
    n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
    n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127,
    n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
    n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
    n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
    n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
    n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172,
    n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181,
    n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
    n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199,
    n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
    n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
    n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
    n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
    n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244,
    n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253,
    n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
    n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271,
    n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
    n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
    n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
    n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
    n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316,
    n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325,
    n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
    n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343,
    n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
    n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
    n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397,
    n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415,
    n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
    n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
    n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469,
    n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487,
    n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
    n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
    n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541,
    n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
    n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559,
    n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568,
    n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
    n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
    n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
    n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604,
    n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613,
    n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
    n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631,
    n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640,
    n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
    n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
    n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
    n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676,
    n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685,
    n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
    n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703,
    n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712,
    n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
    n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
    n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
    n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748,
    n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757,
    n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
    n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775,
    n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
    n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
    n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
    n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
    n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820,
    n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829,
    n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847,
    n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856,
    n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
    n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
    n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
    n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892,
    n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901,
    n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
    n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919,
    n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928,
    n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
    n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
    n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
    n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964,
    n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973,
    n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
    n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991,
    n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000,
    n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
    n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
    n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
    n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036,
    n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045,
    n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
    n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063,
    n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072,
    n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
    n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
    n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
    n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108,
    n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117,
    n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
    n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135,
    n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144,
    n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
    n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
    n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
    n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180,
    n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189,
    n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
    n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207,
    n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216,
    n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
    n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
    n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
    n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252,
    n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261,
    n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
    n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279,
    n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288,
    n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
    n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
    n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
    n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324,
    n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333,
    n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
    n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351,
    n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
    n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
    n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
    n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
    n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396,
    n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405,
    n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
    n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423,
    n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
    n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
    n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
    n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468,
    n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477,
    n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
    n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495,
    n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504,
    n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
    n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
    n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
    n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540,
    n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549,
    n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
    n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567,
    n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
    n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
    n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
    n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
    n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612,
    n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621,
    n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
    n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639,
    n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648,
    n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
    n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
    n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
    n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684,
    n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693,
    n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
    n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711,
    n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720,
    n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729,
    n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
    n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
    n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756,
    n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765,
    n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
    n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783,
    n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792,
    n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801,
    n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
    n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
    n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828,
    n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837,
    n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
    n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855,
    n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
    n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873,
    n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
    n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
    n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900,
    n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909,
    n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
    n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927,
    n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936,
    n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945,
    n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
    n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
    n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972,
    n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
    n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999,
    n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008,
    n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
    n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
    n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
    n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044,
    n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053,
    n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
    n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071,
    n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080,
    n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089,
    n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
    n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
    n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116,
    n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125,
    n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
    n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143,
    n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
    n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161,
    n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
    n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
    n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188,
    n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197,
    n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
    n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215,
    n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224,
    n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233,
    n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
    n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
    n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260,
    n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269,
    n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
    n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287,
    n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296,
    n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
    n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
    n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
    n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332,
    n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341,
    n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
    n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359,
    n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
    n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
    n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
    n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
    n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404,
    n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413,
    n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
    n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431,
    n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440,
    n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
    n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
    n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
    n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476,
    n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485,
    n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503,
    n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521,
    n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
    n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539,
    n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548,
    n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557,
    n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
    n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575,
    n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584,
    n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593,
    n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
    n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611,
    n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620,
    n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629,
    n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
    n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647,
    n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656,
    n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665,
    n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
    n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683,
    n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692,
    n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701,
    n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
    n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719,
    n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
    n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737,
    n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
    n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755,
    n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764,
    n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773,
    n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
    n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791,
    n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
    n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
    n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
    n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
    n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836,
    n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845,
    n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
    n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863,
    n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
    n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
    n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
    n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
    n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908,
    n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917,
    n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
    n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935,
    n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
    n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
    n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
    n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989,
    n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
    n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007,
    n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
    n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
    n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
    n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
    n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052,
    n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061,
    n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
    n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079,
    n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
    n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
    n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
    n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
    n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124,
    n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133,
    n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
    n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151,
    n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
    n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
    n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
    n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
    n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196,
    n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205,
    n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
    n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223,
    n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
    n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
    n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
    n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
    n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268,
    n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277,
    n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
    n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295,
    n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
    n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
    n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
    n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
    n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340,
    n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349,
    n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
    n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367,
    n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
    n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
    n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
    n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
    n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412,
    n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
    n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
    n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439,
    n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
    n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
    n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
    n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
    n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484,
    n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493,
    n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
    n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511,
    n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
    n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
    n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
    n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
    n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556,
    n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565,
    n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
    n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583,
    n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
    n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
    n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
    n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
    n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628,
    n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637,
    n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
    n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655,
    n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
    n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
    n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
    n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
    n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700,
    n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709,
    n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
    n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727,
    n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736,
    n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
    n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
    n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
    n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772,
    n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781,
    n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790,
    n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799,
    n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808,
    n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
    n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
    n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835,
    n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844,
    n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853,
    n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862,
    n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871,
    n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
    n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
    n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
    n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
    n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916,
    n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925,
    n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934,
    n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943,
    n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952,
    n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
    n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
    n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
    n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988,
    n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997,
    n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
    n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015,
    n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
    n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
    n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
    n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051,
    n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060,
    n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069,
    n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078,
    n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087,
    n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096,
    n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
    n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
    n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123,
    n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132,
    n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141,
    n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150,
    n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159,
    n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168,
    n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
    n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
    n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195,
    n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204,
    n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213,
    n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222,
    n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231,
    n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240,
    n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
    n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
    n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267,
    n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276,
    n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285,
    n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
    n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303,
    n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
    n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
    n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
    n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
    n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348,
    n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357,
    n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366,
    n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375,
    n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384,
    n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
    n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
    n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
    n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420,
    n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429,
    n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438,
    n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447,
    n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456,
    n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
    n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
    n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
    n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492,
    n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501,
    n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510,
    n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519,
    n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528,
    n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537,
    n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
    n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
    n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564,
    n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573,
    n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
    n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591,
    n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600,
    n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609,
    n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
    n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
    n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636,
    n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645,
    n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
    n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663,
    n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
    n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
    n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
    n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
    n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708,
    n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
    n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735,
    n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744,
    n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753,
    n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
    n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
    n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780,
    n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789,
    n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798,
    n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807,
    n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816,
    n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825,
    n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
    n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
    n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852,
    n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861,
    n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
    n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879,
    n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888,
    n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897,
    n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
    n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915,
    n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924,
    n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933,
    n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942,
    n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951,
    n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960,
    n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969,
    n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
    n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
    n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996,
    n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005,
    n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014,
    n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023,
    n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032,
    n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041,
    n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
    n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059,
    n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068,
    n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077,
    n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
    n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095,
    n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104,
    n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113,
    n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
    n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131,
    n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140,
    n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149,
    n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
    n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167,
    n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176,
    n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185,
    n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
    n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203,
    n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212,
    n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221,
    n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
    n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239,
    n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
    n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
    n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
    n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
    n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284,
    n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293,
    n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
    n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311,
    n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
    n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329,
    n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
    n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347,
    n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356,
    n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365,
    n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374,
    n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383,
    n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392,
    n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401,
    n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
    n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419,
    n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428,
    n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437,
    n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446,
    n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455,
    n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
    n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473,
    n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
    n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491,
    n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500,
    n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509,
    n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
    n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527,
    n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536,
    n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545,
    n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
    n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563,
    n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572,
    n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581,
    n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
    n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599,
    n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608,
    n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617,
    n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
    n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635,
    n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644,
    n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653,
    n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
    n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671,
    n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680,
    n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689,
    n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
    n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707,
    n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716,
    n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725,
    n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734,
    n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743,
    n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752,
    n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761,
    n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
    n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
    n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788,
    n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797,
    n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806,
    n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815,
    n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824,
    n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833,
    n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
    n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851,
    n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860,
    n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869,
    n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
    n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887,
    n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896,
    n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905,
    n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
    n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923,
    n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932,
    n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941,
    n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
    n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959,
    n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
    n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977,
    n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
    n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
    n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004,
    n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013,
    n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
    n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031,
    n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
    n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049,
    n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
    n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067,
    n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076,
    n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085,
    n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094,
    n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103,
    n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112,
    n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121,
    n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
    n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139,
    n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148,
    n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157,
    n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166,
    n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175,
    n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
    n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193,
    n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
    n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211,
    n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220,
    n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229,
    n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238,
    n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247,
    n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256,
    n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265,
    n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
    n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283,
    n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292,
    n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301,
    n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310,
    n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319,
    n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
    n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337,
    n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
    n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355,
    n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364,
    n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373,
    n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382,
    n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391,
    n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400,
    n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409,
    n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
    n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
    n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436,
    n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445,
    n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
    n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463,
    n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472,
    n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481,
    n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
    n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499,
    n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508,
    n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517,
    n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
    n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535,
    n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544,
    n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553,
    n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
    n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571,
    n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580,
    n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589,
    n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
    n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607,
    n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616,
    n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625,
    n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
    n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
    n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652,
    n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661,
    n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
    n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679,
    n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688,
    n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697,
    n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
    n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715,
    n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724,
    n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733,
    n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
    n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751,
    n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
    n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769,
    n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
    n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787,
    n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796,
    n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805,
    n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
    n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823,
    n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
    n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841,
    n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
    n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859,
    n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868,
    n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877,
    n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
    n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895,
    n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904,
    n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913,
    n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
    n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
    n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940,
    n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949,
    n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
    n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967,
    n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976,
    n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985,
    n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
    n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003,
    n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012,
    n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021,
    n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
    n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039,
    n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
    n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057,
    n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
    n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
    n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084,
    n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093,
    n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
    n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111,
    n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
    n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129,
    n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
    n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147,
    n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156,
    n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165,
    n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174,
    n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183,
    n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
    n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201,
    n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
    n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219,
    n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228,
    n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237,
    n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
    n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255,
    n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
    n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273,
    n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
    n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
    n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300,
    n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309,
    n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
    n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327,
    n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
    n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345,
    n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
    n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363,
    n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372,
    n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381,
    n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390,
    n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399,
    n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
    n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417,
    n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
    n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435,
    n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444,
    n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453,
    n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462,
    n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471,
    n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
    n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489,
    n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
    n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
    n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
    n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525,
    n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534,
    n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543,
    n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
    n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561,
    n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
    n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
    n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588,
    n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597,
    n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606,
    n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615,
    n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
    n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633,
    n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
    n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
    n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660,
    n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669,
    n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678,
    n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687,
    n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696,
    n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705,
    n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
    n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723,
    n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732,
    n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741,
    n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
    n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759,
    n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768,
    n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777,
    n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
    n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795,
    n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804,
    n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813,
    n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822,
    n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831,
    n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840,
    n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
    n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
    n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867,
    n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876,
    n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885,
    n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894,
    n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903,
    n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
    n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921,
    n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
    n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939,
    n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948,
    n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957,
    n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966,
    n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975,
    n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984,
    n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993,
    n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
    n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011,
    n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020,
    n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029,
    n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
    n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047,
    n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
    n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065,
    n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
    n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083,
    n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092,
    n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101,
    n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
    n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119,
    n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
    n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137,
    n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
    n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155,
    n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164,
    n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173,
    n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182,
    n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191,
    n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200,
    n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209,
    n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
    n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227,
    n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236,
    n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245,
    n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254,
    n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263,
    n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272,
    n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281,
    n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
    n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299,
    n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308,
    n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317,
    n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326,
    n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335,
    n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
    n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353,
    n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
    n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371,
    n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380,
    n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389,
    n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398,
    n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407,
    n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
    n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425,
    n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
    n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443,
    n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452,
    n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461,
    n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470,
    n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479,
    n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488,
    n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497,
    n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
    n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515,
    n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524,
    n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533,
    n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542,
    n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551,
    n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560,
    n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569,
    n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
    n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587,
    n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
    n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605,
    n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614,
    n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623,
    n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
    n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641,
    n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
    n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659,
    n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
    n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677,
    n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686,
    n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695,
    n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704,
    n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713,
    n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
    n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731,
    n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740,
    n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748, n51749,
    n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758,
    n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767,
    n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776,
    n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785,
    n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
    n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803,
    n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812,
    n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820, n51821,
    n51822, n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830,
    n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838, n51839,
    n51840, n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848,
    n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857,
    n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
    n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875,
    n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884,
    n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893,
    n51894, n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902,
    n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911,
    n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920,
    n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929,
    n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
    n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947,
    n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956,
    n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965,
    n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974,
    n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983,
    n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
    n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001,
    n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
    n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019,
    n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028,
    n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037,
    n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
    n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055,
    n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
    n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073,
    n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
    n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091,
    n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100,
    n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109,
    n52110, n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118,
    n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127,
    n52128, n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136,
    n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145,
    n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
    n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163,
    n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172,
    n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180, n52181,
    n52182, n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190,
    n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198, n52199,
    n52200, n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208,
    n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217,
    n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
    n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235,
    n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244,
    n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252, n52253,
    n52254, n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262,
    n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270, n52271,
    n52272, n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280,
    n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289,
    n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
    n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307,
    n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316,
    n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325,
    n52326, n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334,
    n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342, n52343,
    n52344, n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352,
    n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361,
    n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
    n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379,
    n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388,
    n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397,
    n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406,
    n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415,
    n52416, n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424,
    n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433,
    n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
    n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451,
    n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460,
    n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469,
    n52470, n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478,
    n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487,
    n52488, n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496,
    n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505,
    n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
    n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523,
    n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532,
    n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540, n52541,
    n52542, n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550,
    n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558, n52559,
    n52560, n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568,
    n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577,
    n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
    n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595,
    n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604,
    n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612, n52613,
    n52614, n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622,
    n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631,
    n52632, n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640,
    n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649,
    n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
    n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667,
    n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676,
    n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684, n52685,
    n52686, n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694,
    n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702, n52703,
    n52704, n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712,
    n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721,
    n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
    n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739,
    n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748,
    n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756, n52757,
    n52758, n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766,
    n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774, n52775,
    n52776, n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784,
    n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793,
    n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
    n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811,
    n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820,
    n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828, n52829,
    n52830, n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838,
    n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846, n52847,
    n52848, n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856,
    n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865,
    n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
    n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883,
    n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892,
    n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900, n52901,
    n52902, n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910,
    n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918, n52919,
    n52920, n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928,
    n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937,
    n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
    n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955,
    n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964,
    n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972, n52973,
    n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982,
    n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990, n52991,
    n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000,
    n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009,
    n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
    n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027,
    n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
    n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045,
    n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054,
    n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063,
    n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072,
    n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081,
    n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
    n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099,
    n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
    n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117,
    n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126,
    n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135,
    n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144,
    n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153,
    n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
    n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171,
    n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180,
    n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189,
    n53190, n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198,
    n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206, n53207,
    n53208, n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216,
    n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225,
    n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
    n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243,
    n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252,
    n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260, n53261,
    n53262, n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270,
    n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279,
    n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288,
    n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297,
    n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
    n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315,
    n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324,
    n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332, n53333,
    n53334, n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342,
    n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350, n53351,
    n53352, n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360,
    n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369,
    n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
    n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387,
    n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396,
    n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405,
    n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414,
    n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422, n53423,
    n53424, n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432,
    n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441,
    n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
    n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459,
    n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468,
    n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477,
    n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486,
    n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494, n53495,
    n53496, n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504,
    n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513,
    n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
    n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531,
    n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540,
    n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549,
    n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558,
    n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, n53567,
    n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576,
    n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585,
    n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
    n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603,
    n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612,
    n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621,
    n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630,
    n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639,
    n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648,
    n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657,
    n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
    n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675,
    n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684,
    n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693,
    n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702,
    n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710, n53711,
    n53712, n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720,
    n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729,
    n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
    n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747,
    n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756,
    n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765,
    n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774,
    n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783,
    n53784, n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792,
    n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801,
    n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
    n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819,
    n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828,
    n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837,
    n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846,
    n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855,
    n53856, n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864,
    n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873,
    n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
    n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891,
    n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900,
    n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909,
    n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918,
    n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927,
    n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936,
    n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945,
    n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
    n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963,
    n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972,
    n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981,
    n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990,
    n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999,
    n54000, n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008,
    n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017,
    n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
    n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035,
    n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044,
    n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053,
    n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062,
    n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070, n54071,
    n54072, n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080,
    n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089,
    n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
    n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107,
    n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116,
    n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124, n54125,
    n54126, n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134,
    n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143,
    n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152,
    n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161,
    n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
    n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179,
    n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188,
    n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197,
    n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206,
    n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215,
    n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224,
    n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233,
    n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
    n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251,
    n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260,
    n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269,
    n54270, n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278,
    n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287,
    n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296,
    n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305,
    n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
    n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323,
    n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332,
    n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340, n54341,
    n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349, n54350,
    n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359,
    n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368,
    n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377,
    n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
    n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395,
    n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404,
    n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413,
    n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422,
    n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431,
    n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440,
    n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449,
    n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
    n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467,
    n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476,
    n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485,
    n54486, n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494,
    n54495, n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503,
    n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512,
    n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521,
    n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
    n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539,
    n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548,
    n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54557,
    n54558, n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566,
    n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575,
    n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584,
    n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593,
    n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
    n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611,
    n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620,
    n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629,
    n54630, n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638,
    n54639, n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647,
    n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656,
    n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665,
    n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
    n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683,
    n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692,
    n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700, n54701,
    n54702, n54703, n54704, n54705, n54706, n54707, n54708, n54709, n54710,
    n54711, n54712, n54713, n54714, n54715, n54716, n54717, n54718, n54719,
    n54720, n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728,
    n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737,
    n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
    n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755,
    n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764,
    n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772, n54773,
    n54774, n54775, n54776, n54777, n54778, n54779, n54780, n54781, n54782,
    n54783, n54784, n54785, n54786, n54787, n54788, n54789, n54790, n54791,
    n54792, n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800,
    n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809,
    n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
    n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827,
    n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836,
    n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844, n54845,
    n54846, n54847, n54848, n54849, n54850, n54851, n54852, n54853, n54854,
    n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862, n54863,
    n54864, n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872,
    n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
    n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
    n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899,
    n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908,
    n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916, n54917,
    n54918, n54919, n54920, n54921, n54922, n54923, n54924, n54925, n54926,
    n54927, n54928, n54929, n54930, n54931, n54932, n54933, n54934, n54935,
    n54936, n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944,
    n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953,
    n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962,
    n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971,
    n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980,
    n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988, n54989,
    n54990, n54991, n54992, n54993, n54994, n54995, n54996, n54997, n54998,
    n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007,
    n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016,
    n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025,
    n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034,
    n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043,
    n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052,
    n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061,
    n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070,
    n55071, n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079,
    n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088,
    n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097,
    n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106,
    n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115,
    n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124,
    n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132, n55133,
    n55134, n55135, n55136, n55137, n55138, n55139, n55140, n55141, n55142,
    n55143, n55144, n55145, n55146, n55147, n55148, n55149, n55150, n55151,
    n55152, n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160,
    n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169,
    n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178,
    n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187,
    n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196,
    n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205,
    n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55213, n55214,
    n55215, n55216, n55217, n55218, n55219, n55220, n55221, n55222, n55223,
    n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232,
    n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241,
    n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250,
    n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259,
    n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268,
    n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277,
    n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285, n55286,
    n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295,
    n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304,
    n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313,
    n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322,
    n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331,
    n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340,
    n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349,
    n55350, n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358,
    n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366, n55367,
    n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376,
    n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385,
    n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394,
    n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403,
    n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412,
    n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420, n55421,
    n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430,
    n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439,
    n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448,
    n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457,
    n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
    n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475,
    n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484,
    n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492, n55493,
    n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502,
    n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511,
    n55512, n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520,
    n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529,
    n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538,
    n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547,
    n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556,
    n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565,
    n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574,
    n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582, n55583,
    n55584, n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592,
    n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601,
    n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610,
    n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619,
    n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628,
    n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636, n55637,
    n55638, n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646,
    n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655,
    n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664,
    n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673,
    n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682,
    n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691,
    n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700,
    n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708, n55709,
    n55710, n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718,
    n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726, n55727,
    n55728, n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736,
    n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745,
    n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754,
    n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763,
    n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772,
    n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780, n55781,
    n55782, n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790,
    n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799,
    n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808,
    n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817,
    n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826,
    n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835,
    n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844,
    n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852, n55853,
    n55854, n55855, n55856, n55857, n55858, n55859, n55860, n55861, n55862,
    n55863, n55864, n55865, n55866, n55867, n55868, n55869, n55870, n55871,
    n55872, n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880,
    n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889,
    n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898,
    n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907,
    n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916,
    n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924, n55925,
    n55926, n55927, n55928, n55929, n55930, n55931, n55932, n55933, n55934,
    n55935, n55936, n55937, n55938, n55939, n55940, n55941, n55942, n55943,
    n55944, n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952,
    n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961,
    n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970,
    n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979,
    n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988,
    n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996, n55997,
    n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006,
    n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015,
    n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024,
    n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033,
    n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
    n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051,
    n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060,
    n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069,
    n56070, n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078,
    n56079, n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087,
    n56088, n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096,
    n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105,
    n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114,
    n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123,
    n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132,
    n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140, n56141,
    n56142, n56143, n56144, n56145, n56146, n56147, n56148, n56149, n56150,
    n56151, n56152, n56153, n56154, n56155, n56156, n56157, n56158, n56159,
    n56160, n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168,
    n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177,
    n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186,
    n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195,
    n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204,
    n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212, n56213,
    n56214, n56215, n56216, n56217, n56218, n56219, n56220, n56221, n56222,
    n56223, n56224, n56225, n56226, n56227, n56228, n56229, n56230, n56231,
    n56232, n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240,
    n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249,
    n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258,
    n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267,
    n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276,
    n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285,
    n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293, n56294,
    n56295, n56296, n56297, n56298, n56299, n56300, n56301, n56302, n56303,
    n56304, n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312,
    n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321,
    n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330,
    n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339,
    n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348,
    n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356, n56357,
    n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365, n56366,
    n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374, n56375,
    n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384,
    n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393,
    n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402,
    n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410, n56411,
    n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420,
    n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428, n56429,
    n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437, n56438,
    n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446, n56447,
    n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456,
    n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465,
    n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474,
    n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483,
    n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492,
    n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500, n56501,
    n56502, n56503, n56504, n56505, n56506, n56507, n56508, n56509, n56510,
    n56511, n56512, n56513, n56514, n56515, n56516, n56517, n56518, n56519,
    n56520, n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528,
    n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537,
    n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
    n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555,
    n56556, n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564,
    n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572, n56573,
    n56574, n56575, n56576, n56577, n56578, n56579, n56580, n56581, n56582,
    n56583, n56584, n56585, n56586, n56587, n56588, n56589, n56590, n56591,
    n56592, n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600,
    n56601, n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609,
    n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618,
    n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626, n56627,
    n56628, n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636,
    n56637, n56638, n56639, n56640, n56641, n56642, n56643, n56644, n56645,
    n56646, n56647, n56648, n56649, n56650, n56651, n56652, n56653, n56654,
    n56655, n56656, n56657, n56658, n56659, n56660, n56661, n56662, n56663,
    n56664, n56665, n56666, n56667, n56668, n56669, n56670, n56671, n56672,
    n56673, n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681,
    n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690,
    n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698, n56699,
    n56700, n56701, n56702, n56703, n56704, n56705, n56706, n56707, n56708,
    n56709, n56710, n56711, n56712, n56713, n56714, n56715, n56716, n56717,
    n56718, n56719, n56720, n56721, n56722, n56723, n56724, n56725, n56726,
    n56727, n56728, n56729, n56730, n56731, n56732, n56733, n56734, n56735,
    n56736, n56737, n56738, n56739, n56740, n56741, n56742, n56743, n56744,
    n56745, n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753,
    n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762,
    n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770, n56771,
    n56772, n56773, n56774, n56775, n56776, n56777, n56778, n56779, n56780,
    n56781, n56782, n56783, n56784, n56785, n56786, n56787, n56788, n56789,
    n56790, n56791, n56792, n56793, n56794, n56795, n56796, n56797, n56798,
    n56799, n56800, n56801, n56802, n56803, n56804, n56805, n56806, n56807,
    n56808, n56809, n56810, n56811, n56812, n56813, n56814, n56815, n56816,
    n56817, n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825,
    n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834,
    n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842, n56843,
    n56844, n56845, n56846, n56847, n56848, n56849, n56850, n56851, n56852,
    n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860, n56861,
    n56862, n56863, n56864, n56865, n56866, n56867, n56868, n56869, n56870,
    n56871, n56872, n56873, n56874, n56875, n56876, n56877, n56878, n56879,
    n56880, n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888,
    n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897,
    n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
    n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914, n56915,
    n56916, n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924,
    n56925, n56926, n56927, n56928, n56929, n56930, n56931, n56932, n56933,
    n56934, n56935, n56936, n56937, n56938, n56939, n56940, n56941, n56942,
    n56943, n56944, n56945, n56946, n56947, n56948, n56949, n56950, n56951,
    n56952, n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960,
    n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969,
    n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978,
    n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986, n56987,
    n56988, n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996,
    n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004, n57005,
    n57006, n57007, n57008, n57009, n57010, n57011, n57012, n57013, n57014,
    n57015, n57016, n57017, n57018, n57019, n57020, n57021, n57022, n57023,
    n57024, n57025, n57026, n57027, n57028, n57029, n57030, n57031, n57032,
    n57033, n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041,
    n57042, n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050,
    n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058, n57059,
    n57060, n57061, n57062, n57063, n57064, n57065, n57066, n57067, n57068,
    n57069, n57070, n57071, n57072, n57073, n57074, n57075, n57076, n57077,
    n57078, n57079, n57080, n57081, n57082, n57083, n57084, n57085, n57086,
    n57087, n57088, n57089, n57090, n57091, n57092, n57093, n57094, n57095,
    n57096, n57097, n57098, n57099, n57100, n57101, n57102, n57103, n57104,
    n57105, n57106, n57107, n57108, n57109, n57110, n57111, n57112, n57113,
    n57114, n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122,
    n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130, n57131,
    n57132, n57133, n57134, n57135, n57136, n57137, n57138, n57139, n57140,
    n57141, n57142, n57143, n57144, n57145, n57146, n57147, n57148, n57149,
    n57150, n57151, n57152, n57153, n57154, n57155, n57156, n57157, n57158,
    n57159, n57160, n57161, n57162, n57163, n57164, n57165, n57166, n57167,
    n57168, n57169, n57170, n57171, n57172, n57173, n57174, n57175, n57176,
    n57177, n57178, n57179, n57180, n57181, n57182, n57183, n57184, n57185,
    n57186, n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194,
    n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202, n57203,
    n57204, n57205, n57206, n57207, n57208, n57209, n57210, n57211, n57212,
    n57213, n57214, n57215, n57216, n57217, n57218, n57219, n57220, n57221,
    n57222, n57223, n57224, n57225, n57226, n57227, n57228, n57229, n57230,
    n57231, n57232, n57233, n57234, n57235, n57236, n57237, n57238, n57239,
    n57240, n57241, n57242, n57243, n57244, n57245, n57246, n57247, n57248,
    n57249, n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257,
    n57258, n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266,
    n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274, n57275,
    n57276, n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57284,
    n57285, n57286, n57287, n57288, n57289, n57290, n57291, n57292, n57293,
    n57294, n57295, n57296, n57297, n57298, n57299, n57300, n57301, n57302,
    n57303, n57304, n57305, n57306, n57307, n57308, n57309, n57310, n57311,
    n57312, n57313, n57314, n57315, n57316, n57317, n57318, n57319, n57320,
    n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328, n57329,
    n57330, n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338,
    n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346, n57347,
    n57348, n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356,
    n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364, n57365,
    n57366, n57367, n57368, n57369, n57370, n57371, n57372, n57373, n57374,
    n57375, n57376, n57377, n57378, n57379, n57380, n57381, n57382, n57383,
    n57384, n57385, n57386, n57387, n57388, n57389, n57390, n57391, n57392,
    n57393, n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401,
    n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410,
    n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418, n57419,
    n57420, n57421, n57422, n57423, n57424, n57425, n57426, n57427, n57428,
    n57429, n57430, n57431, n57432, n57433, n57434, n57435, n57436, n57437,
    n57438, n57439, n57440, n57441, n57442, n57443, n57444, n57445, n57446,
    n57447, n57448, n57449, n57450, n57451, n57452, n57453, n57454, n57455,
    n57456, n57457, n57458, n57459, n57460, n57461, n57462, n57463, n57464,
    n57465, n57466, n57467, n57468, n57469, n57470, n57471, n57472, n57473,
    n57474, n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482,
    n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490, n57491,
    n57492, n57493, n57494, n57495, n57496, n57497, n57498, n57499, n57500,
    n57501, n57502, n57503, n57504, n57505, n57506, n57507, n57508, n57509,
    n57510, n57511, n57512, n57513, n57514, n57515, n57516, n57517, n57518,
    n57519, n57520, n57521, n57522, n57523, n57524, n57525, n57526, n57527,
    n57528, n57529, n57530, n57531, n57532, n57533, n57534, n57535, n57536,
    n57537, n57538, n57539, n57540, n57541, n57542, n57543, n57544, n57545,
    n57546, n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554,
    n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562, n57563,
    n57564, n57565, n57566, n57567, n57568, n57569, n57570, n57571, n57572,
    n57573, n57574, n57575, n57576, n57577, n57578, n57579, n57580, n57581,
    n57582, n57583, n57584, n57585, n57586, n57587, n57588, n57589, n57590,
    n57591, n57592, n57593, n57594, n57595, n57596, n57597, n57598, n57599,
    n57600, n57601, n57602, n57603, n57604, n57605, n57606, n57607, n57608,
    n57609, n57610, n57611, n57612, n57613, n57614, n57615, n57616, n57617,
    n57618, n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626,
    n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634, n57635,
    n57636, n57637, n57638, n57639, n57640, n57641, n57642, n57643, n57644,
    n57645, n57646, n57647, n57648, n57649, n57650, n57651, n57652, n57653,
    n57654, n57655, n57656, n57657, n57658, n57659, n57660, n57661, n57662,
    n57663, n57664, n57665, n57666, n57667, n57668, n57669, n57670, n57671,
    n57672, n57673, n57674, n57675, n57676, n57677, n57678, n57679, n57680,
    n57681, n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689,
    n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698,
    n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706, n57707,
    n57708, n57709, n57710, n57711, n57712, n57713, n57714, n57715, n57716,
    n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724, n57725,
    n57726, n57727, n57728, n57729, n57730, n57731, n57732, n57733, n57734,
    n57735, n57736, n57737, n57738, n57739, n57740, n57741, n57742, n57743,
    n57744, n57745, n57746, n57747, n57748, n57749, n57750, n57751, n57752,
    n57753, n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761,
    n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
    n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778, n57779,
    n57780, n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788,
    n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796, n57797,
    n57798, n57799, n57800, n57801, n57802, n57803, n57804, n57805, n57806,
    n57807, n57808, n57809, n57810, n57811, n57812, n57813, n57814, n57815,
    n57816, n57817, n57818, n57819, n57820, n57821, n57822, n57823, n57824,
    n57825, n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833,
    n57834, n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842,
    n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850, n57851,
    n57852, n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860,
    n57861, n57862, n57863, n57864, n57865, n57866, n57867, n57868, n57869,
    n57870, n57871, n57872, n57873, n57874, n57875, n57876, n57877, n57878,
    n57879, n57880, n57881, n57882, n57883, n57884, n57885, n57886, n57887,
    n57888, n57889, n57890, n57891, n57892, n57893, n57894, n57895, n57896,
    n57897, n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905,
    n57906, n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
    n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922, n57923,
    n57924, n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932,
    n57933, n57934, n57935, n57936, n57937, n57938, n57939, n57940, n57941,
    n57942, n57943, n57944, n57945, n57946, n57947, n57948, n57949, n57950,
    n57951, n57952, n57953, n57954, n57955, n57956, n57957, n57958, n57959,
    n57960, n57961, n57962, n57963, n57964, n57965, n57966, n57967, n57968,
    n57969, n57970, n57971, n57972, n57973, n57974, n57975, n57976, n57977,
    n57978, n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
    n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994, n57995,
    n57996, n57997, n57998, n57999, n58000, n58001, n58002, n58003, n58004,
    n58005, n58006, n58007, n58008, n58009, n58010, n58011, n58012, n58013,
    n58014, n58015, n58016, n58017, n58018, n58019, n58020, n58021, n58022,
    n58023, n58024, n58025, n58026, n58027, n58028, n58029, n58030, n58031,
    n58032, n58033, n58034, n58035, n58036, n58037, n58038, n58039, n58040,
    n58041, n58042, n58043, n58044, n58045, n58046, n58047, n58048, n58049,
    n58050, n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058,
    n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066, n58067,
    n58068, n58069, n58070, n58071, n58072, n58073, n58074, n58075, n58076,
    n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084, n58085,
    n58086, n58087, n58088, n58089, n58090, n58091, n58092, n58093, n58094,
    n58095, n58096, n58097, n58098, n58099, n58100, n58101, n58102, n58103,
    n58104, n58105, n58106, n58107, n58108, n58109, n58110, n58111, n58112,
    n58113, n58114, n58115, n58116, n58117, n58118, n58119, n58120, n58121,
    n58122, n58123, n58124, n58125;
  assign n71 = ~reg_stateA1_out & ~fair_cnt<0>_out ;
  assign n72 = ~fair_cnt<0>_out  & ~n71;
  assign n73 = ~fair_cnt<1>_out  & ~n72;
  assign n74 = ~fair_cnt<1>_out  & ~n73;
  assign n75 = ~next_env_fair_out & ~n74;
  assign n76 = ~next_env_fair_out & ~n75;
  assign n77 = fair_cnt<2>_out  & ~n76;
  assign n78 = ~reg_stateA1_out & ~fair_cnt<2>_out ;
  assign n79 = ~n77 & ~n78;
  assign n80 = reg_controllable_hmastlock_out & ~n79;
  assign n81 = reg_stateG3_0_out & ~reg_stateG3_1_out;
  assign n82 = ~reg_stateG3_1_out & ~n81;
  assign n83 = ~reg_stateG3_2_out & ~n82;
  assign n84 = ~reg_stateG3_2_out & ~n83;
  assign n85 = ~reg_stateG2_out & ~n84;
  assign n86 = ~reg_stateG2_out & ~n85;
  assign n87 = reg_stateA1_out & ~n86;
  assign n88 = reg_stateA1_out & ~n87;
  assign n89 = ~fair_cnt<0>_out  & ~n88;
  assign n90 = ~fair_cnt<0>_out  & ~n89;
  assign n91 = ~fair_cnt<1>_out  & ~n90;
  assign n92 = ~fair_cnt<1>_out  & ~n91;
  assign n93 = ~next_env_fair_out & ~n92;
  assign n94 = ~next_env_fair_out & ~n93;
  assign n95 = fair_cnt<2>_out  & ~n94;
  assign n96 = ~fair_cnt<2>_out  & ~n88;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~reg_controllable_hmastlock_out & ~n97;
  assign n99 = ~n80 & ~n98;
  assign n100 = reg_controllable_locked_out & ~n99;
  assign n101 = reg_controllable_hmastlock_out & ~n97;
  assign n102 = ~reg_controllable_hmastlock_out & ~n79;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~reg_controllable_locked_out & ~n103;
  assign n105 = ~n100 & ~n104;
  assign n106 = ~reg_controllable_hgrant1_out & ~n105;
  assign n107 = ~reg_controllable_hgrant1_out & ~n106;
  assign n108 = reg_controllable_hmaster2_out & ~n107;
  assign n109 = ~reg_controllable_hgrant1_out & ~n97;
  assign n110 = ~reg_controllable_hgrant1_out & ~n109;
  assign n111 = ~reg_controllable_hmaster2_out & ~n110;
  assign n112 = ~n108 & ~n111;
  assign n113 = reg_controllable_hmaster0_out & ~n112;
  assign n114 = reg_controllable_hmaster1_out & ~n112;
  assign n115 = ~reg_controllable_hmaster1_out & ~n110;
  assign n116 = ~n114 & ~n115;
  assign n117 = ~reg_controllable_hmaster0_out & ~n116;
  assign n118 = ~n113 & ~n117;
  assign n119 = ~reg_controllable_hgrant2_out & ~n118;
  assign n120 = ~reg_controllable_hgrant2_out & ~n119;
  assign n121 = ~reg_controllable_hgrant3_out & ~n120;
  assign n122 = ~reg_controllable_hgrant3_out & ~n121;
  assign n123 = ~reg_controllable_hgrant4_out & ~n122;
  assign n124 = ~reg_controllable_hgrant4_out & ~n123;
  assign n125 = reg_controllable_nhgrant0_out & ~n124;
  assign n126 = reg_controllable_nhgrant0_out & ~n125;
  assign n127 = reg_i_hready_out & ~n126;
  assign n128 = ~reg_stateG2_out & ~n82;
  assign n129 = ~reg_stateG2_out & ~n128;
  assign n130 = reg_stateA1_out & ~n129;
  assign n131 = reg_stateA1_out & ~n130;
  assign n132 = ~fair_cnt<0>_out  & ~n131;
  assign n133 = ~fair_cnt<0>_out  & ~n132;
  assign n134 = ~fair_cnt<1>_out  & ~n133;
  assign n135 = ~fair_cnt<1>_out  & ~n134;
  assign n136 = ~next_env_fair_out & ~n135;
  assign n137 = ~next_env_fair_out & ~n136;
  assign n138 = fair_cnt<2>_out  & ~n137;
  assign n139 = ~fair_cnt<2>_out  & ~n131;
  assign n140 = ~n138 & ~n139;
  assign n141 = ~reg_controllable_hmastlock_out & ~n140;
  assign n142 = ~n80 & ~n141;
  assign n143 = reg_controllable_locked_out & ~n142;
  assign n144 = reg_controllable_hmastlock_out & ~n140;
  assign n145 = ~n102 & ~n144;
  assign n146 = ~reg_controllable_locked_out & ~n145;
  assign n147 = ~n143 & ~n146;
  assign n148 = ~reg_controllable_hgrant1_out & ~n147;
  assign n149 = ~reg_controllable_hgrant1_out & ~n148;
  assign n150 = reg_controllable_hmaster2_out & ~n149;
  assign n151 = reg_controllable_hmaster2_out & ~n150;
  assign n152 = reg_controllable_hmaster0_out & ~n151;
  assign n153 = reg_controllable_hmaster1_out & ~n151;
  assign n154 = reg_controllable_hmaster1_out & ~n153;
  assign n155 = ~reg_controllable_hmaster0_out & ~n154;
  assign n156 = ~n152 & ~n155;
  assign n157 = ~reg_controllable_hgrant2_out & ~n156;
  assign n158 = ~reg_controllable_hgrant2_out & ~n157;
  assign n159 = ~reg_controllable_hgrant3_out & ~n158;
  assign n160 = ~reg_controllable_hgrant3_out & ~n159;
  assign n161 = ~reg_controllable_hgrant4_out & ~n160;
  assign n162 = ~reg_controllable_hgrant4_out & ~n161;
  assign n163 = reg_controllable_nhgrant0_out & ~n162;
  assign n164 = reg_controllable_nhgrant0_out & ~n163;
  assign n165 = ~reg_i_hready_out & ~n164;
  assign n166 = ~n127 & ~n165;
  assign n167 = next_sys_fair<3>_out  & ~n166;
  assign n168 = ~reg_stateA1_out & ~n86;
  assign n169 = ~reg_stateA1_out & ~n168;
  assign n170 = ~fair_cnt<0>_out  & ~n169;
  assign n171 = ~fair_cnt<0>_out  & ~n170;
  assign n172 = ~fair_cnt<1>_out  & ~n171;
  assign n173 = ~fair_cnt<1>_out  & ~n172;
  assign n174 = fair_cnt<2>_out  & ~n173;
  assign n175 = ~fair_cnt<2>_out  & ~n169;
  assign n176 = ~n174 & ~n175;
  assign n177 = reg_controllable_locked_out & ~n176;
  assign n178 = ~fair_cnt<0>_out  & ~n86;
  assign n179 = ~fair_cnt<0>_out  & ~n178;
  assign n180 = ~fair_cnt<1>_out  & ~n179;
  assign n181 = ~fair_cnt<1>_out  & ~n180;
  assign n182 = fair_cnt<2>_out  & ~n181;
  assign n183 = ~fair_cnt<2>_out  & ~n86;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~reg_controllable_locked_out & ~n184;
  assign n186 = ~n177 & ~n185;
  assign n187 = ~reg_controllable_hgrant1_out & ~n186;
  assign n188 = ~reg_controllable_hgrant1_out & ~n187;
  assign n189 = ~reg_stateG10_4_out & ~n188;
  assign n190 = ~reg_stateG10_4_out & ~n189;
  assign n191 = ~next_sys_fair<0>_out  & ~n190;
  assign n192 = ~next_sys_fair<0>_out  & ~n191;
  assign n193 = next_sys_fair<1>_out  & ~n192;
  assign n194 = ~fair_cnt<2>_out  & ~n173;
  assign n195 = ~fair_cnt<2>_out  & ~n194;
  assign n196 = reg_controllable_locked_out & ~n195;
  assign n197 = fair_cnt<1>_out  & ~n179;
  assign n198 = ~fair_cnt<1>_out  & ~n86;
  assign n199 = ~n197 & ~n198;
  assign n200 = next_env_fair_out & ~n199;
  assign n201 = ~next_env_fair_out & ~n86;
  assign n202 = ~n200 & ~n201;
  assign n203 = ~fair_cnt<2>_out  & ~n202;
  assign n204 = ~fair_cnt<2>_out  & ~n203;
  assign n205 = ~reg_controllable_locked_out & ~n204;
  assign n206 = ~n196 & ~n205;
  assign n207 = ~reg_controllable_hgrant1_out & ~n206;
  assign n208 = ~reg_controllable_hgrant1_out & ~n207;
  assign n209 = ~reg_stateG10_4_out & ~n208;
  assign n210 = ~reg_stateG10_4_out & ~n209;
  assign n211 = ~next_sys_fair<1>_out  & ~n210;
  assign n212 = ~n193 & ~n211;
  assign n213 = reg_controllable_hmaster0_out & ~n212;
  assign n214 = reg_controllable_hmaster1_out & ~n212;
  assign n215 = reg_stateG3_2_out & ~n82;
  assign n216 = reg_stateA1_out & n215;
  assign n217 = ~reg_stateG2_out & n215;
  assign n218 = ~reg_stateG2_out & ~n217;
  assign n219 = ~reg_stateA1_out & ~n218;
  assign n220 = ~n216 & ~n219;
  assign n221 = ~fair_cnt<0>_out  & ~n220;
  assign n222 = ~fair_cnt<0>_out  & ~n221;
  assign n223 = ~fair_cnt<1>_out  & ~n222;
  assign n224 = ~fair_cnt<1>_out  & ~n223;
  assign n225 = fair_cnt<2>_out  & ~n224;
  assign n226 = ~fair_cnt<2>_out  & ~n220;
  assign n227 = ~n225 & ~n226;
  assign n228 = reg_controllable_hmastlock_out & ~n227;
  assign n229 = ~reg_controllable_hmastlock_out & ~n176;
  assign n230 = ~n228 & ~n229;
  assign n231 = reg_controllable_locked_out & ~n230;
  assign n232 = reg_controllable_hmastlock_out & ~n184;
  assign n233 = ~reg_controllable_hmastlock_out & ~n227;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~reg_controllable_locked_out & ~n234;
  assign n236 = ~n231 & ~n235;
  assign n237 = ~reg_controllable_hgrant1_out & ~n236;
  assign n238 = ~reg_controllable_hgrant1_out & ~n237;
  assign n239 = ~reg_stateG10_4_out & ~n238;
  assign n240 = ~reg_stateG10_4_out & ~n239;
  assign n241 = ~next_sys_fair<0>_out  & ~n240;
  assign n242 = ~next_sys_fair<0>_out  & ~n241;
  assign n243 = next_sys_fair<1>_out  & ~n242;
  assign n244 = reg_stateG3_0_out & reg_stateG3_1_out;
  assign n245 = ~reg_stateG3_0_out & ~reg_stateG3_1_out;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~reg_stateG3_2_out & n246;
  assign n248 = ~n215 & ~n247;
  assign n249 = reg_stateA1_out & ~n248;
  assign n250 = ~reg_stateG2_out & ~n248;
  assign n251 = ~reg_stateG2_out & ~n250;
  assign n252 = ~reg_stateA1_out & ~n251;
  assign n253 = ~n249 & ~n252;
  assign n254 = ~fair_cnt<0>_out  & ~n253;
  assign n255 = ~fair_cnt<0>_out  & ~n254;
  assign n256 = fair_cnt<1>_out  & ~n255;
  assign n257 = ~reg_stateG3_1_out & ~n245;
  assign n258 = ~reg_stateG3_2_out & n257;
  assign n259 = ~n215 & ~n258;
  assign n260 = reg_stateA1_out & ~n259;
  assign n261 = ~reg_stateG2_out & ~n259;
  assign n262 = ~reg_stateG2_out & ~n261;
  assign n263 = ~reg_stateA1_out & ~n262;
  assign n264 = ~n260 & ~n263;
  assign n265 = fair_cnt<0>_out  & ~n264;
  assign n266 = ~n221 & ~n265;
  assign n267 = ~fair_cnt<1>_out  & ~n266;
  assign n268 = ~n256 & ~n267;
  assign n269 = next_env_fair_out & ~n268;
  assign n270 = reg_stateA1_out & ~n82;
  assign n271 = ~reg_stateA1_out & ~n129;
  assign n272 = ~n270 & ~n271;
  assign n273 = fair_cnt<0>_out  & ~n272;
  assign n274 = ~n254 & ~n273;
  assign n275 = fair_cnt<1>_out  & ~n274;
  assign n276 = ~n267 & ~n275;
  assign n277 = ~next_env_fair_out & ~n276;
  assign n278 = ~n269 & ~n277;
  assign n279 = ~fair_cnt<2>_out  & ~n278;
  assign n280 = ~fair_cnt<2>_out  & ~n279;
  assign n281 = reg_controllable_hmastlock_out & ~n280;
  assign n282 = ~reg_controllable_hmastlock_out & ~n195;
  assign n283 = ~n281 & ~n282;
  assign n284 = reg_controllable_locked_out & ~n283;
  assign n285 = reg_controllable_hmastlock_out & ~n204;
  assign n286 = ~reg_controllable_hmastlock_out & ~n280;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~reg_controllable_locked_out & ~n287;
  assign n289 = ~n284 & ~n288;
  assign n290 = ~reg_controllable_hgrant1_out & ~n289;
  assign n291 = ~reg_controllable_hgrant1_out & ~n290;
  assign n292 = ~reg_stateG10_4_out & ~n291;
  assign n293 = ~reg_stateG10_4_out & ~n292;
  assign n294 = ~next_sys_fair<1>_out  & ~n293;
  assign n295 = ~n243 & ~n294;
  assign n296 = reg_controllable_hmaster2_out & ~n295;
  assign n297 = ~reg_controllable_hmaster2_out & ~n212;
  assign n298 = ~n296 & ~n297;
  assign n299 = ~reg_controllable_hmaster1_out & ~n298;
  assign n300 = ~n214 & ~n299;
  assign n301 = ~reg_controllable_hmaster0_out & ~n300;
  assign n302 = ~n213 & ~n301;
  assign n303 = next_sys_fair<2>_out  & ~n302;
  assign n304 = next_sys_fair<1>_out  & ~n210;
  assign n305 = ~next_sys_fair<1>_out  & ~n190;
  assign n306 = ~n304 & ~n305;
  assign n307 = reg_controllable_hmaster0_out & ~n306;
  assign n308 = reg_controllable_hmaster1_out & ~n306;
  assign n309 = next_sys_fair<1>_out  & ~n293;
  assign n310 = reg_stateA1_out & ~n84;
  assign n311 = ~n168 & ~n310;
  assign n312 = ~fair_cnt<0>_out  & ~n311;
  assign n313 = ~fair_cnt<0>_out  & ~n312;
  assign n314 = ~fair_cnt<1>_out  & ~n313;
  assign n315 = ~fair_cnt<1>_out  & ~n314;
  assign n316 = fair_cnt<2>_out  & ~n315;
  assign n317 = ~fair_cnt<2>_out  & ~n276;
  assign n318 = ~n316 & ~n317;
  assign n319 = reg_controllable_hmastlock_out & ~n318;
  assign n320 = ~n229 & ~n319;
  assign n321 = reg_controllable_locked_out & ~n320;
  assign n322 = ~reg_controllable_hmastlock_out & ~n318;
  assign n323 = ~n232 & ~n322;
  assign n324 = ~reg_controllable_locked_out & ~n323;
  assign n325 = ~n321 & ~n324;
  assign n326 = ~reg_controllable_hgrant1_out & ~n325;
  assign n327 = ~reg_controllable_hgrant1_out & ~n326;
  assign n328 = ~reg_stateG10_4_out & ~n327;
  assign n329 = ~reg_stateG10_4_out & ~n328;
  assign n330 = next_sys_fair<0>_out  & ~n329;
  assign n331 = ~fair_cnt<0>_out  & ~n218;
  assign n332 = ~fair_cnt<0>_out  & ~n331;
  assign n333 = ~fair_cnt<1>_out  & ~n332;
  assign n334 = ~fair_cnt<1>_out  & ~n333;
  assign n335 = next_env_fair_out & ~n334;
  assign n336 = ~next_env_fair_out & ~n224;
  assign n337 = ~n335 & ~n336;
  assign n338 = fair_cnt<2>_out  & ~n337;
  assign n339 = ~n226 & ~n338;
  assign n340 = reg_controllable_hmastlock_out & ~n339;
  assign n341 = ~n229 & ~n340;
  assign n342 = reg_controllable_locked_out & ~n341;
  assign n343 = ~reg_controllable_hmastlock_out & ~n339;
  assign n344 = ~n232 & ~n343;
  assign n345 = ~reg_controllable_locked_out & ~n344;
  assign n346 = ~n342 & ~n345;
  assign n347 = ~reg_controllable_hgrant1_out & ~n346;
  assign n348 = ~reg_controllable_hgrant1_out & ~n347;
  assign n349 = ~reg_stateG10_4_out & ~n348;
  assign n350 = ~reg_stateG10_4_out & ~n349;
  assign n351 = ~next_sys_fair<0>_out  & ~n350;
  assign n352 = ~n330 & ~n351;
  assign n353 = ~next_sys_fair<1>_out  & ~n352;
  assign n354 = ~n309 & ~n353;
  assign n355 = reg_controllable_hmaster2_out & ~n354;
  assign n356 = ~reg_controllable_hmaster2_out & ~n306;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~reg_controllable_hmaster1_out & ~n357;
  assign n359 = ~n308 & ~n358;
  assign n360 = ~reg_controllable_hmaster0_out & ~n359;
  assign n361 = ~n307 & ~n360;
  assign n362 = ~next_sys_fair<2>_out  & ~n361;
  assign n363 = ~n303 & ~n362;
  assign n364 = ~reg_controllable_hgrant2_out & ~n363;
  assign n365 = ~reg_controllable_hgrant2_out & ~n364;
  assign n366 = ~reg_controllable_hgrant3_out & ~n365;
  assign n367 = ~reg_controllable_hgrant3_out & ~n366;
  assign n368 = reg_controllable_hgrant4_out & ~n367;
  assign n369 = ~next_sys_fair<0>_out  & ~n208;
  assign n370 = ~next_sys_fair<0>_out  & ~n369;
  assign n371 = next_sys_fair<1>_out  & ~n370;
  assign n372 = next_sys_fair<0>_out  & ~n188;
  assign n373 = ~n369 & ~n372;
  assign n374 = ~next_sys_fair<1>_out  & ~n373;
  assign n375 = ~n371 & ~n374;
  assign n376 = reg_controllable_hmaster2_out & ~n375;
  assign n377 = ~next_sys_fair<0>_out  & ~n291;
  assign n378 = ~next_sys_fair<0>_out  & ~n377;
  assign n379 = next_sys_fair<1>_out  & ~n378;
  assign n380 = next_sys_fair<0>_out  & ~n238;
  assign n381 = ~n377 & ~n380;
  assign n382 = ~next_sys_fair<1>_out  & ~n381;
  assign n383 = ~n379 & ~n382;
  assign n384 = ~reg_controllable_hmaster2_out & ~n383;
  assign n385 = ~n376 & ~n384;
  assign n386 = reg_controllable_hmaster1_out & ~n385;
  assign n387 = ~reg_controllable_hmaster1_out & ~n375;
  assign n388 = ~n386 & ~n387;
  assign n389 = reg_controllable_hmaster0_out & ~n388;
  assign n390 = ~reg_controllable_hmaster0_out & ~n375;
  assign n391 = ~n389 & ~n390;
  assign n392 = next_sys_fair<2>_out  & ~n391;
  assign n393 = next_sys_fair<1>_out  & ~n208;
  assign n394 = ~next_sys_fair<1>_out  & ~n188;
  assign n395 = ~n393 & ~n394;
  assign n396 = reg_controllable_hmaster2_out & ~n395;
  assign n397 = next_sys_fair<1>_out  & ~n291;
  assign n398 = next_sys_fair<0>_out  & ~n327;
  assign n399 = ~next_sys_fair<0>_out  & ~n348;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~next_sys_fair<1>_out  & ~n400;
  assign n402 = ~n397 & ~n401;
  assign n403 = ~reg_controllable_hmaster2_out & ~n402;
  assign n404 = ~n396 & ~n403;
  assign n405 = reg_controllable_hmaster1_out & ~n404;
  assign n406 = ~reg_controllable_hmaster1_out & ~n395;
  assign n407 = ~n405 & ~n406;
  assign n408 = reg_controllable_hmaster0_out & ~n407;
  assign n409 = ~reg_controllable_hmaster0_out & ~n395;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~next_sys_fair<2>_out  & ~n410;
  assign n412 = ~n392 & ~n411;
  assign n413 = ~reg_stateG10_3_out & ~n412;
  assign n414 = ~reg_stateG10_3_out & ~n413;
  assign n415 = ~reg_controllable_hgrant2_out & ~n414;
  assign n416 = ~reg_controllable_hgrant2_out & ~n415;
  assign n417 = reg_controllable_hgrant3_out & ~n416;
  assign n418 = next_sys_fair<0>_out  & ~n208;
  assign n419 = ~next_sys_fair<0>_out  & ~n188;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~next_sys_fair<1>_out  & ~n420;
  assign n422 = ~n371 & ~n421;
  assign n423 = reg_controllable_hmaster0_out & ~n422;
  assign n424 = reg_controllable_hmaster2_out & ~n422;
  assign n425 = next_sys_fair<0>_out  & ~n291;
  assign n426 = ~next_sys_fair<0>_out  & ~n238;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~next_sys_fair<1>_out  & ~n427;
  assign n429 = ~n379 & ~n428;
  assign n430 = ~reg_controllable_hmaster2_out & ~n429;
  assign n431 = ~n424 & ~n430;
  assign n432 = reg_controllable_hmaster1_out & ~n431;
  assign n433 = ~reg_controllable_hmaster1_out & ~n422;
  assign n434 = ~n432 & ~n433;
  assign n435 = ~reg_controllable_hmaster0_out & ~n434;
  assign n436 = ~n423 & ~n435;
  assign n437 = ~reg_stateG10_2_out & ~n436;
  assign n438 = ~reg_stateG10_2_out & ~n437;
  assign n439 = next_sys_fair<2>_out  & ~n438;
  assign n440 = reg_controllable_hmaster0_out & ~n395;
  assign n441 = ~reg_controllable_hmaster0_out & ~n407;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~reg_stateG10_2_out & ~n442;
  assign n444 = ~reg_stateG10_2_out & ~n443;
  assign n445 = ~next_sys_fair<2>_out  & ~n444;
  assign n446 = ~n439 & ~n445;
  assign n447 = reg_controllable_hgrant2_out & ~n446;
  assign n448 = next_sys_fair<0>_out  & ~n107;
  assign n449 = ~reg_stateG10_1_out & ~n206;
  assign n450 = ~reg_stateG10_1_out & ~n449;
  assign n451 = reg_controllable_hgrant1_out & ~n450;
  assign n452 = reg_stateA1_out & fair_cnt<0>_out ;
  assign n453 = ~reg_stateA1_out & n248;
  assign n454 = ~reg_stateA1_out & ~n453;
  assign n455 = ~fair_cnt<0>_out  & ~n454;
  assign n456 = ~n452 & ~n455;
  assign n457 = fair_cnt<1>_out  & ~n456;
  assign n458 = ~reg_stateA1_out & n259;
  assign n459 = ~reg_stateA1_out & ~n458;
  assign n460 = fair_cnt<0>_out  & ~n459;
  assign n461 = ~reg_stateA1_out & ~n215;
  assign n462 = ~reg_stateA1_out & ~n461;
  assign n463 = ~fair_cnt<0>_out  & ~n462;
  assign n464 = ~n460 & ~n463;
  assign n465 = ~fair_cnt<1>_out  & ~n464;
  assign n466 = ~n457 & ~n465;
  assign n467 = next_env_fair_out & ~n466;
  assign n468 = ~reg_stateA1_out & n82;
  assign n469 = ~reg_stateA1_out & ~n468;
  assign n470 = fair_cnt<0>_out  & ~n469;
  assign n471 = ~n455 & ~n470;
  assign n472 = fair_cnt<1>_out  & ~n471;
  assign n473 = ~n465 & ~n472;
  assign n474 = ~next_env_fair_out & ~n473;
  assign n475 = ~n467 & ~n474;
  assign n476 = ~fair_cnt<2>_out  & n475;
  assign n477 = ~n77 & ~n476;
  assign n478 = reg_controllable_hmastlock_out & ~n477;
  assign n479 = fair_cnt<1>_out  & ~n88;
  assign n480 = fair_cnt<0>_out  & ~n88;
  assign n481 = ~n178 & ~n480;
  assign n482 = ~fair_cnt<1>_out  & ~n481;
  assign n483 = ~n479 & ~n482;
  assign n484 = ~fair_cnt<2>_out  & ~n483;
  assign n485 = ~n95 & ~n484;
  assign n486 = ~reg_controllable_hmastlock_out & ~n485;
  assign n487 = ~n478 & ~n486;
  assign n488 = reg_controllable_locked_out & ~n487;
  assign n489 = fair_cnt<1>_out  & ~n481;
  assign n490 = ~n198 & ~n489;
  assign n491 = next_env_fair_out & ~n490;
  assign n492 = ~n201 & ~n491;
  assign n493 = ~fair_cnt<2>_out  & ~n492;
  assign n494 = ~n95 & ~n493;
  assign n495 = reg_controllable_hmastlock_out & ~n494;
  assign n496 = ~reg_controllable_hmastlock_out & ~n477;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~reg_controllable_locked_out & ~n497;
  assign n499 = ~n488 & ~n498;
  assign n500 = ~reg_controllable_hgrant1_out & ~n499;
  assign n501 = ~n451 & ~n500;
  assign n502 = ~next_sys_fair<0>_out  & ~n501;
  assign n503 = ~n448 & ~n502;
  assign n504 = next_sys_fair<1>_out  & ~n503;
  assign n505 = ~next_sys_fair<1>_out  & ~n501;
  assign n506 = ~n504 & ~n505;
  assign n507 = reg_controllable_hmaster2_out & ~n506;
  assign n508 = next_sys_fair<0>_out  & ~n110;
  assign n509 = reg_controllable_locked_out & ~n485;
  assign n510 = ~reg_controllable_locked_out & ~n494;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~reg_controllable_hgrant1_out & ~n511;
  assign n513 = ~n451 & ~n512;
  assign n514 = ~next_sys_fair<0>_out  & ~n513;
  assign n515 = ~n508 & ~n514;
  assign n516 = next_sys_fair<1>_out  & ~n515;
  assign n517 = ~next_sys_fair<1>_out  & ~n513;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~reg_controllable_hmaster2_out & ~n518;
  assign n520 = ~n507 & ~n519;
  assign n521 = reg_controllable_hmaster1_out & ~n520;
  assign n522 = ~reg_stateG10_1_out & ~n289;
  assign n523 = ~reg_stateG10_1_out & ~n522;
  assign n524 = reg_controllable_hgrant1_out & ~n523;
  assign n525 = ~n512 & ~n524;
  assign n526 = ~next_sys_fair<0>_out  & ~n525;
  assign n527 = ~n508 & ~n526;
  assign n528 = next_sys_fair<1>_out  & ~n527;
  assign n529 = ~next_sys_fair<1>_out  & ~n525;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~reg_controllable_hmaster2_out & ~n530;
  assign n532 = ~n507 & ~n531;
  assign n533 = ~reg_controllable_hmaster1_out & ~n532;
  assign n534 = ~n521 & ~n533;
  assign n535 = reg_controllable_hmaster0_out & ~n534;
  assign n536 = ~reg_controllable_hmaster1_out & ~n518;
  assign n537 = ~n521 & ~n536;
  assign n538 = ~reg_controllable_hmaster0_out & ~n537;
  assign n539 = ~n535 & ~n538;
  assign n540 = next_sys_fair<2>_out  & ~n539;
  assign n541 = ~reg_stateG10_1_out & ~n186;
  assign n542 = ~reg_stateG10_1_out & ~n541;
  assign n543 = reg_controllable_hgrant1_out & ~n542;
  assign n544 = ~n500 & ~n543;
  assign n545 = next_sys_fair<0>_out  & ~n544;
  assign n546 = ~n502 & ~n545;
  assign n547 = next_sys_fair<1>_out  & ~n546;
  assign n548 = ~fair_cnt<0>_out  & ~n84;
  assign n549 = ~fair_cnt<0>_out  & ~n548;
  assign n550 = ~fair_cnt<1>_out  & ~n549;
  assign n551 = ~fair_cnt<1>_out  & ~n550;
  assign n552 = next_env_fair_out & ~n551;
  assign n553 = ~reg_stateA1_out & n84;
  assign n554 = ~reg_stateA1_out & ~n553;
  assign n555 = ~fair_cnt<0>_out  & n554;
  assign n556 = ~fair_cnt<0>_out  & ~n555;
  assign n557 = ~fair_cnt<1>_out  & ~n556;
  assign n558 = ~fair_cnt<1>_out  & ~n557;
  assign n559 = ~next_env_fair_out & ~n558;
  assign n560 = ~n552 & ~n559;
  assign n561 = fair_cnt<2>_out  & ~n560;
  assign n562 = ~fair_cnt<2>_out  & n473;
  assign n563 = ~n561 & ~n562;
  assign n564 = reg_controllable_hmastlock_out & ~n563;
  assign n565 = ~reg_controllable_hmastlock_out & ~n184;
  assign n566 = ~n564 & ~n565;
  assign n567 = reg_controllable_locked_out & ~n566;
  assign n568 = ~reg_controllable_hmastlock_out & ~n563;
  assign n569 = ~n232 & ~n568;
  assign n570 = ~reg_controllable_locked_out & ~n569;
  assign n571 = ~n567 & ~n570;
  assign n572 = ~reg_controllable_hgrant1_out & ~n571;
  assign n573 = ~n543 & ~n572;
  assign n574 = next_sys_fair<0>_out  & ~n573;
  assign n575 = reg_stateG2_out & reg_stateA1_out;
  assign n576 = ~n219 & ~n575;
  assign n577 = ~fair_cnt<0>_out  & ~n576;
  assign n578 = ~fair_cnt<0>_out  & ~n577;
  assign n579 = ~fair_cnt<1>_out  & ~n578;
  assign n580 = ~fair_cnt<1>_out  & ~n579;
  assign n581 = next_env_fair_out & ~n580;
  assign n582 = ~fair_cnt<0>_out  & n462;
  assign n583 = ~fair_cnt<0>_out  & ~n582;
  assign n584 = ~fair_cnt<1>_out  & ~n583;
  assign n585 = ~fair_cnt<1>_out  & ~n584;
  assign n586 = ~next_env_fair_out & ~n585;
  assign n587 = ~n581 & ~n586;
  assign n588 = fair_cnt<2>_out  & ~n587;
  assign n589 = ~fair_cnt<2>_out  & n462;
  assign n590 = ~n588 & ~n589;
  assign n591 = reg_controllable_hmastlock_out & ~n590;
  assign n592 = ~n565 & ~n591;
  assign n593 = reg_controllable_locked_out & ~n592;
  assign n594 = ~reg_controllable_hmastlock_out & ~n590;
  assign n595 = ~n232 & ~n594;
  assign n596 = ~reg_controllable_locked_out & ~n595;
  assign n597 = ~n593 & ~n596;
  assign n598 = ~reg_controllable_hgrant1_out & ~n597;
  assign n599 = ~n543 & ~n598;
  assign n600 = ~next_sys_fair<0>_out  & ~n599;
  assign n601 = ~n574 & ~n600;
  assign n602 = ~next_sys_fair<1>_out  & ~n601;
  assign n603 = ~n547 & ~n602;
  assign n604 = reg_controllable_hmaster2_out & ~n603;
  assign n605 = ~n512 & ~n543;
  assign n606 = next_sys_fair<0>_out  & ~n605;
  assign n607 = ~n514 & ~n606;
  assign n608 = next_sys_fair<1>_out  & ~n607;
  assign n609 = ~reg_controllable_hgrant1_out & ~n184;
  assign n610 = ~n543 & ~n609;
  assign n611 = ~next_sys_fair<1>_out  & ~n610;
  assign n612 = ~n608 & ~n611;
  assign n613 = ~reg_controllable_hmaster2_out & ~n612;
  assign n614 = ~n604 & ~n613;
  assign n615 = reg_controllable_hmaster1_out & ~n614;
  assign n616 = ~reg_stateG10_1_out & ~n236;
  assign n617 = ~reg_stateG10_1_out & ~n616;
  assign n618 = reg_controllable_hgrant1_out & ~n617;
  assign n619 = ~n512 & ~n618;
  assign n620 = next_sys_fair<0>_out  & ~n619;
  assign n621 = ~n526 & ~n620;
  assign n622 = next_sys_fair<1>_out  & ~n621;
  assign n623 = ~reg_stateG10_1_out & ~n325;
  assign n624 = ~reg_stateG10_1_out & ~n623;
  assign n625 = reg_controllable_hgrant1_out & ~n624;
  assign n626 = ~n609 & ~n625;
  assign n627 = next_sys_fair<0>_out  & ~n626;
  assign n628 = ~reg_stateG10_1_out & ~n346;
  assign n629 = ~reg_stateG10_1_out & ~n628;
  assign n630 = reg_controllable_hgrant1_out & ~n629;
  assign n631 = ~n609 & ~n630;
  assign n632 = ~next_sys_fair<0>_out  & ~n631;
  assign n633 = ~n627 & ~n632;
  assign n634 = ~next_sys_fair<1>_out  & ~n633;
  assign n635 = ~n622 & ~n634;
  assign n636 = ~reg_controllable_hmaster2_out & ~n635;
  assign n637 = ~n604 & ~n636;
  assign n638 = ~reg_controllable_hmaster1_out & ~n637;
  assign n639 = ~n615 & ~n638;
  assign n640 = reg_controllable_hmaster0_out & ~n639;
  assign n641 = ~reg_controllable_hmaster1_out & ~n612;
  assign n642 = ~n615 & ~n641;
  assign n643 = ~reg_controllable_hmaster0_out & ~n642;
  assign n644 = ~n640 & ~n643;
  assign n645 = ~next_sys_fair<2>_out  & ~n644;
  assign n646 = ~n540 & ~n645;
  assign n647 = ~reg_controllable_hgrant2_out & ~n646;
  assign n648 = ~n447 & ~n647;
  assign n649 = ~reg_controllable_hgrant3_out & ~n648;
  assign n650 = ~n417 & ~n649;
  assign n651 = ~reg_controllable_hgrant4_out & ~n650;
  assign n652 = ~n368 & ~n651;
  assign n653 = reg_controllable_nhgrant0_out & ~n652;
  assign n654 = ~next_sys_fair<1>_out  & ~n208;
  assign n655 = ~n371 & ~n654;
  assign n656 = reg_controllable_hmaster0_out & ~n655;
  assign n657 = reg_controllable_hmaster1_out & ~n655;
  assign n658 = reg_controllable_hmaster2_out & ~n655;
  assign n659 = ~next_sys_fair<1>_out  & ~n291;
  assign n660 = ~n379 & ~n659;
  assign n661 = ~reg_controllable_hmaster2_out & ~n660;
  assign n662 = ~n658 & ~n661;
  assign n663 = ~reg_controllable_hmaster1_out & ~n662;
  assign n664 = ~n657 & ~n663;
  assign n665 = ~reg_controllable_hmaster0_out & ~n664;
  assign n666 = ~n656 & ~n665;
  assign n667 = next_sys_fair<2>_out  & ~n666;
  assign n668 = next_sys_fair<1>_out  & ~n420;
  assign n669 = ~n394 & ~n668;
  assign n670 = reg_controllable_hmaster0_out & ~n669;
  assign n671 = reg_controllable_hmaster1_out & ~n669;
  assign n672 = reg_controllable_hmaster2_out & ~n669;
  assign n673 = next_sys_fair<1>_out  & ~n427;
  assign n674 = ~n401 & ~n673;
  assign n675 = ~reg_controllable_hmaster2_out & ~n674;
  assign n676 = ~n672 & ~n675;
  assign n677 = ~reg_controllable_hmaster1_out & ~n676;
  assign n678 = ~n671 & ~n677;
  assign n679 = ~reg_controllable_hmaster0_out & ~n678;
  assign n680 = ~n670 & ~n679;
  assign n681 = ~next_sys_fair<2>_out  & ~n680;
  assign n682 = ~n667 & ~n681;
  assign n683 = ~reg_controllable_hgrant2_out & ~n682;
  assign n684 = ~reg_controllable_hgrant2_out & ~n683;
  assign n685 = ~reg_controllable_hgrant3_out & ~n684;
  assign n686 = ~reg_controllable_hgrant3_out & ~n685;
  assign n687 = ~reg_controllable_hgrant4_out & ~n686;
  assign n688 = ~reg_controllable_hgrant4_out & ~n687;
  assign n689 = ~reg_controllable_nhgrant0_out & ~n688;
  assign n690 = ~n653 & ~n689;
  assign n691 = reg_i_hready_out & ~n690;
  assign n692 = reg_stateA1_out & ~n270;
  assign n693 = ~fair_cnt<0>_out  & ~n692;
  assign n694 = ~fair_cnt<0>_out  & ~n693;
  assign n695 = ~fair_cnt<1>_out  & ~n694;
  assign n696 = ~fair_cnt<1>_out  & ~n695;
  assign n697 = ~next_env_fair_out & ~n696;
  assign n698 = ~next_env_fair_out & ~n697;
  assign n699 = fair_cnt<2>_out  & ~n698;
  assign n700 = ~fair_cnt<2>_out  & ~n692;
  assign n701 = ~n699 & ~n700;
  assign n702 = reg_controllable_hmastlock_out & ~n701;
  assign n703 = ~fair_cnt<2>_out  & ~n82;
  assign n704 = ~n699 & ~n703;
  assign n705 = ~reg_controllable_hmastlock_out & ~n704;
  assign n706 = ~n702 & ~n705;
  assign n707 = reg_controllable_locked_out & ~n706;
  assign n708 = ~reg_controllable_locked_out & ~n704;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~reg_controllable_hgrant1_out & ~n709;
  assign n711 = ~reg_controllable_hgrant1_out & ~n710;
  assign n712 = ~reg_stateG10_4_out & ~n711;
  assign n713 = ~reg_stateG10_4_out & ~n712;
  assign n714 = ~next_sys_fair<0>_out  & ~n713;
  assign n715 = ~next_sys_fair<0>_out  & ~n714;
  assign n716 = next_sys_fair<1>_out  & ~n715;
  assign n717 = ~fair_cnt<2>_out  & ~n698;
  assign n718 = ~fair_cnt<2>_out  & ~n717;
  assign n719 = reg_controllable_hmastlock_out & ~n718;
  assign n720 = ~fair_cnt<0>_out  & ~n82;
  assign n721 = ~fair_cnt<0>_out  & ~n720;
  assign n722 = ~fair_cnt<1>_out  & ~n721;
  assign n723 = ~fair_cnt<1>_out  & ~n722;
  assign n724 = ~next_env_fair_out & ~n723;
  assign n725 = ~next_env_fair_out & ~n724;
  assign n726 = ~fair_cnt<2>_out  & ~n725;
  assign n727 = ~fair_cnt<2>_out  & ~n726;
  assign n728 = ~reg_controllable_hmastlock_out & ~n727;
  assign n729 = ~n719 & ~n728;
  assign n730 = reg_controllable_locked_out & ~n729;
  assign n731 = fair_cnt<1>_out  & ~n721;
  assign n732 = ~fair_cnt<1>_out  & ~n82;
  assign n733 = ~n731 & ~n732;
  assign n734 = next_env_fair_out & ~n733;
  assign n735 = ~next_env_fair_out & ~n82;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~fair_cnt<2>_out  & ~n736;
  assign n738 = ~fair_cnt<2>_out  & ~n737;
  assign n739 = ~reg_controllable_locked_out & ~n738;
  assign n740 = ~n730 & ~n739;
  assign n741 = ~reg_controllable_hgrant1_out & ~n740;
  assign n742 = ~reg_controllable_hgrant1_out & ~n741;
  assign n743 = ~reg_stateG10_4_out & ~n742;
  assign n744 = ~reg_stateG10_4_out & ~n743;
  assign n745 = ~next_sys_fair<1>_out  & ~n744;
  assign n746 = ~n716 & ~n745;
  assign n747 = reg_controllable_hmaster2_out & ~n746;
  assign n748 = ~reg_stateA1_out & ~n271;
  assign n749 = ~fair_cnt<2>_out  & ~n748;
  assign n750 = ~fair_cnt<2>_out  & ~n749;
  assign n751 = ~reg_controllable_hmastlock_out & ~n750;
  assign n752 = ~reg_controllable_hmastlock_out & ~n751;
  assign n753 = reg_controllable_locked_out & ~n752;
  assign n754 = ~fair_cnt<2>_out  & ~n129;
  assign n755 = ~fair_cnt<2>_out  & ~n754;
  assign n756 = ~reg_controllable_locked_out & ~n755;
  assign n757 = ~n753 & ~n756;
  assign n758 = ~reg_controllable_hgrant1_out & ~n757;
  assign n759 = ~reg_controllable_hgrant1_out & ~n758;
  assign n760 = ~reg_stateG10_4_out & ~n759;
  assign n761 = ~reg_stateG10_4_out & ~n760;
  assign n762 = ~next_sys_fair<0>_out  & ~n761;
  assign n763 = ~next_sys_fair<0>_out  & ~n762;
  assign n764 = next_sys_fair<1>_out  & ~n763;
  assign n765 = ~fair_cnt<0>_out  & ~n748;
  assign n766 = ~fair_cnt<0>_out  & ~n765;
  assign n767 = ~fair_cnt<1>_out  & ~n766;
  assign n768 = ~fair_cnt<1>_out  & ~n767;
  assign n769 = fair_cnt<2>_out  & ~n768;
  assign n770 = ~n749 & ~n769;
  assign n771 = ~reg_controllable_hmastlock_out & ~n770;
  assign n772 = ~reg_controllable_hmastlock_out & ~n771;
  assign n773 = reg_controllable_locked_out & ~n772;
  assign n774 = ~fair_cnt<0>_out  & ~n129;
  assign n775 = ~fair_cnt<0>_out  & ~n774;
  assign n776 = ~fair_cnt<1>_out  & ~n775;
  assign n777 = ~fair_cnt<1>_out  & ~n776;
  assign n778 = fair_cnt<2>_out  & ~n777;
  assign n779 = ~n754 & ~n778;
  assign n780 = ~reg_controllable_locked_out & ~n779;
  assign n781 = ~n773 & ~n780;
  assign n782 = ~reg_controllable_hgrant1_out & ~n781;
  assign n783 = ~reg_controllable_hgrant1_out & ~n782;
  assign n784 = ~reg_stateG10_4_out & ~n783;
  assign n785 = ~reg_stateG10_4_out & ~n784;
  assign n786 = next_sys_fair<0>_out  & ~n785;
  assign n787 = ~next_env_fair_out & ~n768;
  assign n788 = ~next_env_fair_out & ~n787;
  assign n789 = ~fair_cnt<2>_out  & ~n788;
  assign n790 = ~fair_cnt<2>_out  & ~n789;
  assign n791 = ~reg_controllable_hmastlock_out & ~n790;
  assign n792 = ~reg_controllable_hmastlock_out & ~n791;
  assign n793 = reg_controllable_locked_out & ~n792;
  assign n794 = fair_cnt<1>_out  & ~n775;
  assign n795 = ~fair_cnt<1>_out  & ~n129;
  assign n796 = ~n794 & ~n795;
  assign n797 = next_env_fair_out & ~n796;
  assign n798 = ~next_env_fair_out & ~n129;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~fair_cnt<2>_out  & ~n799;
  assign n801 = ~fair_cnt<2>_out  & ~n800;
  assign n802 = ~reg_controllable_locked_out & ~n801;
  assign n803 = ~n793 & ~n802;
  assign n804 = ~reg_controllable_hgrant1_out & ~n803;
  assign n805 = ~reg_controllable_hgrant1_out & ~n804;
  assign n806 = ~reg_stateG10_4_out & ~n805;
  assign n807 = ~reg_stateG10_4_out & ~n806;
  assign n808 = ~next_sys_fair<0>_out  & ~n807;
  assign n809 = ~n786 & ~n808;
  assign n810 = ~next_sys_fair<1>_out  & ~n809;
  assign n811 = ~n764 & ~n810;
  assign n812 = ~reg_controllable_hmaster2_out & ~n811;
  assign n813 = ~n747 & ~n812;
  assign n814 = reg_controllable_hmaster1_out & ~n813;
  assign n815 = ~next_sys_fair<1>_out  & ~n807;
  assign n816 = ~n764 & ~n815;
  assign n817 = ~reg_controllable_hmaster2_out & ~n816;
  assign n818 = ~n747 & ~n817;
  assign n819 = ~reg_controllable_hmaster1_out & ~n818;
  assign n820 = ~n814 & ~n819;
  assign n821 = reg_controllable_hmaster0_out & ~n820;
  assign n822 = next_sys_fair<0>_out  & ~n807;
  assign n823 = ~next_sys_fair<0>_out  & ~n785;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~next_sys_fair<1>_out  & ~n824;
  assign n826 = ~n764 & ~n825;
  assign n827 = ~reg_controllable_hmaster2_out & ~n826;
  assign n828 = ~n747 & ~n827;
  assign n829 = reg_controllable_hmaster1_out & ~n828;
  assign n830 = ~n228 & ~n771;
  assign n831 = reg_controllable_locked_out & ~n830;
  assign n832 = reg_controllable_hmastlock_out & ~n779;
  assign n833 = ~n233 & ~n832;
  assign n834 = ~reg_controllable_locked_out & ~n833;
  assign n835 = ~n831 & ~n834;
  assign n836 = ~reg_controllable_hgrant1_out & ~n835;
  assign n837 = ~reg_controllable_hgrant1_out & ~n836;
  assign n838 = ~reg_stateG10_4_out & ~n837;
  assign n839 = ~reg_stateG10_4_out & ~n838;
  assign n840 = ~next_sys_fair<0>_out  & ~n839;
  assign n841 = ~next_sys_fair<0>_out  & ~n840;
  assign n842 = next_sys_fair<1>_out  & ~n841;
  assign n843 = ~n281 & ~n791;
  assign n844 = reg_controllable_locked_out & ~n843;
  assign n845 = reg_controllable_hmastlock_out & ~n801;
  assign n846 = ~n286 & ~n845;
  assign n847 = ~reg_controllable_locked_out & ~n846;
  assign n848 = ~n844 & ~n847;
  assign n849 = ~reg_controllable_hgrant1_out & ~n848;
  assign n850 = ~reg_controllable_hgrant1_out & ~n849;
  assign n851 = ~reg_stateG10_4_out & ~n850;
  assign n852 = ~reg_stateG10_4_out & ~n851;
  assign n853 = ~next_sys_fair<1>_out  & ~n852;
  assign n854 = ~n842 & ~n853;
  assign n855 = reg_controllable_hmaster2_out & ~n854;
  assign n856 = ~n817 & ~n855;
  assign n857 = ~reg_controllable_hmaster1_out & ~n856;
  assign n858 = ~n829 & ~n857;
  assign n859 = ~reg_controllable_hmaster0_out & ~n858;
  assign n860 = ~n821 & ~n859;
  assign n861 = next_sys_fair<2>_out  & ~n860;
  assign n862 = next_sys_fair<1>_out  & ~n744;
  assign n863 = reg_stateA1_out & ~n310;
  assign n864 = ~fair_cnt<0>_out  & ~n863;
  assign n865 = ~fair_cnt<0>_out  & ~n864;
  assign n866 = ~fair_cnt<1>_out  & ~n865;
  assign n867 = ~fair_cnt<1>_out  & ~n866;
  assign n868 = next_env_fair_out & ~n867;
  assign n869 = ~n697 & ~n868;
  assign n870 = fair_cnt<2>_out  & ~n869;
  assign n871 = ~n700 & ~n870;
  assign n872 = reg_controllable_hmastlock_out & ~n871;
  assign n873 = ~reg_stateA1_out & ~n84;
  assign n874 = ~n270 & ~n873;
  assign n875 = ~fair_cnt<0>_out  & ~n874;
  assign n876 = ~fair_cnt<0>_out  & ~n875;
  assign n877 = ~fair_cnt<1>_out  & ~n876;
  assign n878 = ~fair_cnt<1>_out  & ~n877;
  assign n879 = ~next_env_fair_out & ~n878;
  assign n880 = ~n552 & ~n879;
  assign n881 = fair_cnt<2>_out  & ~n880;
  assign n882 = ~n703 & ~n881;
  assign n883 = ~reg_controllable_hmastlock_out & ~n882;
  assign n884 = ~n872 & ~n883;
  assign n885 = reg_controllable_locked_out & ~n884;
  assign n886 = ~reg_controllable_locked_out & ~n882;
  assign n887 = ~n885 & ~n886;
  assign n888 = ~reg_controllable_hgrant1_out & ~n887;
  assign n889 = ~reg_controllable_hgrant1_out & ~n888;
  assign n890 = ~reg_stateG10_4_out & ~n889;
  assign n891 = ~reg_stateG10_4_out & ~n890;
  assign n892 = next_sys_fair<0>_out  & ~n891;
  assign n893 = next_env_fair_out & ~n135;
  assign n894 = ~n697 & ~n893;
  assign n895 = fair_cnt<2>_out  & ~n894;
  assign n896 = ~n700 & ~n895;
  assign n897 = reg_controllable_hmastlock_out & ~n896;
  assign n898 = next_env_fair_out & ~n777;
  assign n899 = ~n724 & ~n898;
  assign n900 = fair_cnt<2>_out  & ~n899;
  assign n901 = ~n703 & ~n900;
  assign n902 = ~reg_controllable_hmastlock_out & ~n901;
  assign n903 = ~n897 & ~n902;
  assign n904 = reg_controllable_locked_out & ~n903;
  assign n905 = ~reg_controllable_locked_out & ~n901;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~reg_controllable_hgrant1_out & ~n906;
  assign n908 = ~reg_controllable_hgrant1_out & ~n907;
  assign n909 = ~reg_stateG10_4_out & ~n908;
  assign n910 = ~reg_stateG10_4_out & ~n909;
  assign n911 = ~next_sys_fair<0>_out  & ~n910;
  assign n912 = ~n892 & ~n911;
  assign n913 = ~next_sys_fair<1>_out  & ~n912;
  assign n914 = ~n862 & ~n913;
  assign n915 = reg_controllable_hmaster2_out & ~n914;
  assign n916 = next_sys_fair<1>_out  & ~n807;
  assign n917 = ~n174 & ~n749;
  assign n918 = ~reg_controllable_hmastlock_out & ~n917;
  assign n919 = ~reg_controllable_hmastlock_out & ~n918;
  assign n920 = reg_controllable_locked_out & ~n919;
  assign n921 = ~n182 & ~n754;
  assign n922 = ~reg_controllable_locked_out & ~n921;
  assign n923 = ~n920 & ~n922;
  assign n924 = ~reg_controllable_hgrant1_out & ~n923;
  assign n925 = ~reg_controllable_hgrant1_out & ~n924;
  assign n926 = ~reg_stateG10_4_out & ~n925;
  assign n927 = ~reg_stateG10_4_out & ~n926;
  assign n928 = next_sys_fair<0>_out  & ~n927;
  assign n929 = ~n823 & ~n928;
  assign n930 = ~next_sys_fair<1>_out  & ~n929;
  assign n931 = ~n916 & ~n930;
  assign n932 = ~reg_controllable_hmaster2_out & ~n931;
  assign n933 = ~n915 & ~n932;
  assign n934 = reg_controllable_hmaster1_out & ~n933;
  assign n935 = next_sys_fair<1>_out  & ~n809;
  assign n936 = ~n930 & ~n935;
  assign n937 = ~reg_controllable_hmaster2_out & ~n936;
  assign n938 = ~n915 & ~n937;
  assign n939 = ~reg_controllable_hmaster1_out & ~n938;
  assign n940 = ~n934 & ~n939;
  assign n941 = reg_controllable_hmaster0_out & ~n940;
  assign n942 = next_sys_fair<1>_out  & ~n852;
  assign n943 = ~n319 & ~n918;
  assign n944 = reg_controllable_locked_out & ~n943;
  assign n945 = reg_controllable_hmastlock_out & ~n921;
  assign n946 = ~n322 & ~n945;
  assign n947 = ~reg_controllable_locked_out & ~n946;
  assign n948 = ~n944 & ~n947;
  assign n949 = ~reg_controllable_hgrant1_out & ~n948;
  assign n950 = ~reg_controllable_hgrant1_out & ~n949;
  assign n951 = ~reg_stateG10_4_out & ~n950;
  assign n952 = ~reg_stateG10_4_out & ~n951;
  assign n953 = next_sys_fair<0>_out  & ~n952;
  assign n954 = ~n340 & ~n771;
  assign n955 = reg_controllable_locked_out & ~n954;
  assign n956 = ~n343 & ~n832;
  assign n957 = ~reg_controllable_locked_out & ~n956;
  assign n958 = ~n955 & ~n957;
  assign n959 = ~reg_controllable_hgrant1_out & ~n958;
  assign n960 = ~reg_controllable_hgrant1_out & ~n959;
  assign n961 = ~reg_stateG10_4_out & ~n960;
  assign n962 = ~reg_stateG10_4_out & ~n961;
  assign n963 = ~next_sys_fair<0>_out  & ~n962;
  assign n964 = ~n953 & ~n963;
  assign n965 = ~next_sys_fair<1>_out  & ~n964;
  assign n966 = ~n942 & ~n965;
  assign n967 = reg_controllable_hmaster2_out & ~n966;
  assign n968 = next_sys_fair<1>_out  & ~n824;
  assign n969 = ~n930 & ~n968;
  assign n970 = ~reg_controllable_hmaster2_out & ~n969;
  assign n971 = ~n967 & ~n970;
  assign n972 = ~reg_controllable_hmaster1_out & ~n971;
  assign n973 = ~n934 & ~n972;
  assign n974 = ~reg_controllable_hmaster0_out & ~n973;
  assign n975 = ~n941 & ~n974;
  assign n976 = ~next_sys_fair<2>_out  & ~n975;
  assign n977 = ~n861 & ~n976;
  assign n978 = ~reg_controllable_hgrant2_out & ~n977;
  assign n979 = ~reg_controllable_hgrant2_out & ~n978;
  assign n980 = ~reg_controllable_hgrant3_out & ~n979;
  assign n981 = ~reg_controllable_hgrant3_out & ~n980;
  assign n982 = reg_controllable_hgrant4_out & ~n981;
  assign n983 = ~next_sys_fair<0>_out  & ~n742;
  assign n984 = ~next_sys_fair<0>_out  & ~n983;
  assign n985 = next_sys_fair<1>_out  & ~n984;
  assign n986 = next_sys_fair<0>_out  & ~n711;
  assign n987 = ~n983 & ~n986;
  assign n988 = ~next_sys_fair<1>_out  & ~n987;
  assign n989 = ~n985 & ~n988;
  assign n990 = reg_controllable_hmaster2_out & ~n989;
  assign n991 = ~next_sys_fair<0>_out  & ~n850;
  assign n992 = ~next_sys_fair<0>_out  & ~n991;
  assign n993 = next_sys_fair<1>_out  & ~n992;
  assign n994 = next_sys_fair<0>_out  & ~n837;
  assign n995 = ~n991 & ~n994;
  assign n996 = ~next_sys_fair<1>_out  & ~n995;
  assign n997 = ~n993 & ~n996;
  assign n998 = ~reg_controllable_hmaster2_out & ~n997;
  assign n999 = ~n990 & ~n998;
  assign n1000 = reg_controllable_hmaster1_out & ~n999;
  assign n1001 = ~next_sys_fair<0>_out  & ~n805;
  assign n1002 = ~next_sys_fair<0>_out  & ~n1001;
  assign n1003 = next_sys_fair<1>_out  & ~n1002;
  assign n1004 = next_sys_fair<0>_out  & ~n759;
  assign n1005 = ~n1001 & ~n1004;
  assign n1006 = ~next_sys_fair<1>_out  & ~n1005;
  assign n1007 = ~n1003 & ~n1006;
  assign n1008 = ~reg_controllable_hmaster2_out & ~n1007;
  assign n1009 = ~n990 & ~n1008;
  assign n1010 = ~reg_controllable_hmaster1_out & ~n1009;
  assign n1011 = ~n1000 & ~n1010;
  assign n1012 = reg_controllable_hmaster0_out & ~n1011;
  assign n1013 = ~next_sys_fair<0>_out  & ~n783;
  assign n1014 = ~n1004 & ~n1013;
  assign n1015 = ~next_sys_fair<1>_out  & ~n1014;
  assign n1016 = ~n1003 & ~n1015;
  assign n1017 = ~reg_controllable_hmaster2_out & ~n1016;
  assign n1018 = ~n990 & ~n1017;
  assign n1019 = reg_controllable_hmaster1_out & ~n1018;
  assign n1020 = ~next_sys_fair<0>_out  & ~n1013;
  assign n1021 = next_sys_fair<1>_out  & ~n1020;
  assign n1022 = ~n1006 & ~n1021;
  assign n1023 = reg_controllable_hmaster2_out & ~n1022;
  assign n1024 = ~n1008 & ~n1023;
  assign n1025 = ~reg_controllable_hmaster1_out & ~n1024;
  assign n1026 = ~n1019 & ~n1025;
  assign n1027 = ~reg_controllable_hmaster0_out & ~n1026;
  assign n1028 = ~n1012 & ~n1027;
  assign n1029 = next_sys_fair<2>_out  & ~n1028;
  assign n1030 = next_sys_fair<1>_out  & ~n742;
  assign n1031 = next_sys_fair<0>_out  & ~n889;
  assign n1032 = ~next_sys_fair<0>_out  & ~n908;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = ~next_sys_fair<1>_out  & ~n1033;
  assign n1035 = ~n1030 & ~n1034;
  assign n1036 = reg_controllable_hmaster2_out & ~n1035;
  assign n1037 = next_sys_fair<1>_out  & ~n850;
  assign n1038 = next_sys_fair<0>_out  & ~n950;
  assign n1039 = ~next_sys_fair<0>_out  & ~n960;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = ~next_sys_fair<1>_out  & ~n1040;
  assign n1042 = ~n1037 & ~n1041;
  assign n1043 = ~reg_controllable_hmaster2_out & ~n1042;
  assign n1044 = ~n1036 & ~n1043;
  assign n1045 = reg_controllable_hmaster1_out & ~n1044;
  assign n1046 = next_sys_fair<0>_out  & ~n783;
  assign n1047 = ~n1001 & ~n1046;
  assign n1048 = next_sys_fair<1>_out  & ~n1047;
  assign n1049 = next_sys_fair<0>_out  & ~n925;
  assign n1050 = ~n1013 & ~n1049;
  assign n1051 = ~next_sys_fair<1>_out  & ~n1050;
  assign n1052 = ~n1048 & ~n1051;
  assign n1053 = ~reg_controllable_hmaster2_out & ~n1052;
  assign n1054 = ~n1036 & ~n1053;
  assign n1055 = ~reg_controllable_hmaster1_out & ~n1054;
  assign n1056 = ~n1045 & ~n1055;
  assign n1057 = reg_controllable_hmaster0_out & ~n1056;
  assign n1058 = next_sys_fair<1>_out  & ~n805;
  assign n1059 = ~n1051 & ~n1058;
  assign n1060 = ~reg_controllable_hmaster2_out & ~n1059;
  assign n1061 = ~n1036 & ~n1060;
  assign n1062 = reg_controllable_hmaster1_out & ~n1061;
  assign n1063 = reg_controllable_hmaster2_out & ~n1059;
  assign n1064 = next_sys_fair<0>_out  & ~n805;
  assign n1065 = ~n1013 & ~n1064;
  assign n1066 = next_sys_fair<1>_out  & ~n1065;
  assign n1067 = ~n1051 & ~n1066;
  assign n1068 = ~reg_controllable_hmaster2_out & ~n1067;
  assign n1069 = ~n1063 & ~n1068;
  assign n1070 = ~reg_controllable_hmaster1_out & ~n1069;
  assign n1071 = ~n1062 & ~n1070;
  assign n1072 = ~reg_controllable_hmaster0_out & ~n1071;
  assign n1073 = ~n1057 & ~n1072;
  assign n1074 = ~next_sys_fair<2>_out  & ~n1073;
  assign n1075 = ~n1029 & ~n1074;
  assign n1076 = ~reg_stateG10_3_out & ~n1075;
  assign n1077 = ~reg_stateG10_3_out & ~n1076;
  assign n1078 = ~reg_controllable_hgrant2_out & ~n1077;
  assign n1079 = ~reg_controllable_hgrant2_out & ~n1078;
  assign n1080 = reg_controllable_hgrant3_out & ~n1079;
  assign n1081 = next_sys_fair<0>_out  & ~n742;
  assign n1082 = ~next_sys_fair<0>_out  & ~n711;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~next_sys_fair<1>_out  & ~n1083;
  assign n1085 = ~n985 & ~n1084;
  assign n1086 = reg_controllable_hmaster2_out & ~n1085;
  assign n1087 = ~next_sys_fair<0>_out  & ~n759;
  assign n1088 = ~n1046 & ~n1087;
  assign n1089 = ~next_sys_fair<1>_out  & ~n1088;
  assign n1090 = ~n1003 & ~n1089;
  assign n1091 = ~reg_controllable_hmaster2_out & ~n1090;
  assign n1092 = ~n1086 & ~n1091;
  assign n1093 = reg_controllable_hmaster1_out & ~n1092;
  assign n1094 = ~n1064 & ~n1087;
  assign n1095 = ~next_sys_fair<1>_out  & ~n1094;
  assign n1096 = ~n1003 & ~n1095;
  assign n1097 = ~reg_controllable_hmaster2_out & ~n1096;
  assign n1098 = ~n1086 & ~n1097;
  assign n1099 = ~reg_controllable_hmaster1_out & ~n1098;
  assign n1100 = ~n1093 & ~n1099;
  assign n1101 = reg_controllable_hmaster0_out & ~n1100;
  assign n1102 = next_sys_fair<0>_out  & ~n850;
  assign n1103 = ~next_sys_fair<0>_out  & ~n837;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~next_sys_fair<1>_out  & ~n1104;
  assign n1106 = ~n993 & ~n1105;
  assign n1107 = ~reg_controllable_hmaster2_out & ~n1106;
  assign n1108 = ~n1086 & ~n1107;
  assign n1109 = reg_controllable_hmaster1_out & ~n1108;
  assign n1110 = ~n1021 & ~n1095;
  assign n1111 = reg_controllable_hmaster2_out & ~n1110;
  assign n1112 = ~n1097 & ~n1111;
  assign n1113 = ~reg_controllable_hmaster1_out & ~n1112;
  assign n1114 = ~n1109 & ~n1113;
  assign n1115 = ~reg_controllable_hmaster0_out & ~n1114;
  assign n1116 = ~n1101 & ~n1115;
  assign n1117 = ~reg_stateG10_2_out & ~n1116;
  assign n1118 = ~reg_stateG10_2_out & ~n1117;
  assign n1119 = next_sys_fair<2>_out  & ~n1118;
  assign n1120 = ~n1055 & ~n1062;
  assign n1121 = reg_controllable_hmaster0_out & ~n1120;
  assign n1122 = ~n1045 & ~n1070;
  assign n1123 = ~reg_controllable_hmaster0_out & ~n1122;
  assign n1124 = ~n1121 & ~n1123;
  assign n1125 = ~reg_stateG10_2_out & ~n1124;
  assign n1126 = ~reg_stateG10_2_out & ~n1125;
  assign n1127 = ~next_sys_fair<2>_out  & ~n1126;
  assign n1128 = ~n1119 & ~n1127;
  assign n1129 = reg_controllable_hgrant2_out & ~n1128;
  assign n1130 = next_sys_fair<0>_out  & ~n149;
  assign n1131 = ~reg_stateG10_1_out & ~n740;
  assign n1132 = ~reg_stateG10_1_out & ~n1131;
  assign n1133 = reg_controllable_hgrant1_out & ~n1132;
  assign n1134 = next_env_fair_out & ~n131;
  assign n1135 = fair_cnt<1>_out  & ~n131;
  assign n1136 = fair_cnt<0>_out  & ~n131;
  assign n1137 = ~n720 & ~n1136;
  assign n1138 = ~fair_cnt<1>_out  & ~n1137;
  assign n1139 = ~n1135 & ~n1138;
  assign n1140 = ~next_env_fair_out & ~n1139;
  assign n1141 = ~n1134 & ~n1140;
  assign n1142 = ~fair_cnt<2>_out  & ~n1141;
  assign n1143 = ~n138 & ~n1142;
  assign n1144 = ~reg_controllable_hmastlock_out & ~n1143;
  assign n1145 = ~n478 & ~n1144;
  assign n1146 = reg_controllable_locked_out & ~n1145;
  assign n1147 = fair_cnt<1>_out  & ~n1137;
  assign n1148 = ~n732 & ~n1147;
  assign n1149 = next_env_fair_out & ~n1148;
  assign n1150 = ~n735 & ~n1149;
  assign n1151 = ~fair_cnt<2>_out  & ~n1150;
  assign n1152 = ~n138 & ~n1151;
  assign n1153 = reg_controllable_hmastlock_out & ~n1152;
  assign n1154 = ~n496 & ~n1153;
  assign n1155 = ~reg_controllable_locked_out & ~n1154;
  assign n1156 = ~n1146 & ~n1155;
  assign n1157 = ~reg_controllable_hgrant1_out & ~n1156;
  assign n1158 = ~n1133 & ~n1157;
  assign n1159 = ~next_sys_fair<0>_out  & ~n1158;
  assign n1160 = ~n1130 & ~n1159;
  assign n1161 = next_sys_fair<1>_out  & ~n1160;
  assign n1162 = ~next_sys_fair<1>_out  & ~n1158;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = reg_controllable_hmaster2_out & ~n1163;
  assign n1165 = ~reg_stateG10_1_out & ~n803;
  assign n1166 = ~reg_stateG10_1_out & ~n1165;
  assign n1167 = reg_controllable_hgrant1_out & ~n1166;
  assign n1168 = ~next_env_fair_out & ~n777;
  assign n1169 = ~next_env_fair_out & ~n1168;
  assign n1170 = ~fair_cnt<2>_out  & ~n1169;
  assign n1171 = ~fair_cnt<2>_out  & ~n1170;
  assign n1172 = reg_controllable_locked_out & ~n1171;
  assign n1173 = ~n802 & ~n1172;
  assign n1174 = ~reg_controllable_hgrant1_out & ~n1173;
  assign n1175 = ~n1167 & ~n1174;
  assign n1176 = ~next_sys_fair<0>_out  & ~n1175;
  assign n1177 = ~next_sys_fair<0>_out  & ~n1176;
  assign n1178 = next_sys_fair<1>_out  & ~n1177;
  assign n1179 = ~reg_stateG10_1_out & ~n781;
  assign n1180 = ~reg_stateG10_1_out & ~n1179;
  assign n1181 = reg_controllable_hgrant1_out & ~n1180;
  assign n1182 = ~reg_controllable_hgrant1_out & ~n779;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = next_sys_fair<0>_out  & ~n1183;
  assign n1185 = ~n1176 & ~n1184;
  assign n1186 = ~next_sys_fair<1>_out  & ~n1185;
  assign n1187 = ~n1178 & ~n1186;
  assign n1188 = ~reg_controllable_hmaster2_out & ~n1187;
  assign n1189 = ~n1164 & ~n1188;
  assign n1190 = reg_controllable_hmaster1_out & ~n1189;
  assign n1191 = ~reg_stateG10_1_out & ~n848;
  assign n1192 = ~reg_stateG10_1_out & ~n1191;
  assign n1193 = reg_controllable_hgrant1_out & ~n1192;
  assign n1194 = ~n1174 & ~n1193;
  assign n1195 = ~next_sys_fair<0>_out  & ~n1194;
  assign n1196 = ~next_sys_fair<0>_out  & ~n1195;
  assign n1197 = next_sys_fair<1>_out  & ~n1196;
  assign n1198 = ~next_sys_fair<1>_out  & ~n1194;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~reg_controllable_hmaster2_out & ~n1199;
  assign n1201 = ~n1164 & ~n1200;
  assign n1202 = ~reg_controllable_hmaster1_out & ~n1201;
  assign n1203 = ~n1190 & ~n1202;
  assign n1204 = reg_controllable_hmaster0_out & ~n1203;
  assign n1205 = next_sys_fair<0>_out  & ~n1175;
  assign n1206 = ~next_sys_fair<0>_out  & ~n1183;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~next_sys_fair<1>_out  & ~n1207;
  assign n1209 = ~n1178 & ~n1208;
  assign n1210 = ~reg_controllable_hmaster2_out & ~n1209;
  assign n1211 = ~n1164 & ~n1210;
  assign n1212 = reg_controllable_hmaster1_out & ~n1211;
  assign n1213 = ~next_sys_fair<0>_out  & ~n1206;
  assign n1214 = next_sys_fair<1>_out  & ~n1213;
  assign n1215 = ~next_sys_fair<1>_out  & ~n1175;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = reg_controllable_hmaster2_out & ~n1216;
  assign n1218 = ~n1178 & ~n1215;
  assign n1219 = ~reg_controllable_hmaster2_out & ~n1218;
  assign n1220 = ~n1217 & ~n1219;
  assign n1221 = ~reg_controllable_hmaster1_out & ~n1220;
  assign n1222 = ~n1212 & ~n1221;
  assign n1223 = ~reg_controllable_hmaster0_out & ~n1222;
  assign n1224 = ~n1204 & ~n1223;
  assign n1225 = next_sys_fair<2>_out  & ~n1224;
  assign n1226 = ~reg_stateG10_1_out & ~n709;
  assign n1227 = ~reg_stateG10_1_out & ~n1226;
  assign n1228 = reg_controllable_hgrant1_out & ~n1227;
  assign n1229 = ~n1157 & ~n1228;
  assign n1230 = next_sys_fair<0>_out  & ~n1229;
  assign n1231 = ~n1159 & ~n1230;
  assign n1232 = next_sys_fair<1>_out  & ~n1231;
  assign n1233 = ~reg_stateG10_1_out & ~n887;
  assign n1234 = ~reg_stateG10_1_out & ~n1233;
  assign n1235 = reg_controllable_hgrant1_out & ~n1234;
  assign n1236 = ~n564 & ~n883;
  assign n1237 = reg_controllable_locked_out & ~n1236;
  assign n1238 = reg_controllable_hmastlock_out & ~n882;
  assign n1239 = ~n568 & ~n1238;
  assign n1240 = ~reg_controllable_locked_out & ~n1239;
  assign n1241 = ~n1237 & ~n1240;
  assign n1242 = ~reg_controllable_hgrant1_out & ~n1241;
  assign n1243 = ~n1235 & ~n1242;
  assign n1244 = next_sys_fair<0>_out  & ~n1243;
  assign n1245 = ~reg_stateG10_1_out & ~n906;
  assign n1246 = ~reg_stateG10_1_out & ~n1245;
  assign n1247 = reg_controllable_hgrant1_out & ~n1246;
  assign n1248 = ~n591 & ~n902;
  assign n1249 = reg_controllable_locked_out & ~n1248;
  assign n1250 = reg_controllable_hmastlock_out & ~n901;
  assign n1251 = ~n594 & ~n1250;
  assign n1252 = ~reg_controllable_locked_out & ~n1251;
  assign n1253 = ~n1249 & ~n1252;
  assign n1254 = ~reg_controllable_hgrant1_out & ~n1253;
  assign n1255 = ~n1247 & ~n1254;
  assign n1256 = ~next_sys_fair<0>_out  & ~n1255;
  assign n1257 = ~n1244 & ~n1256;
  assign n1258 = ~next_sys_fair<1>_out  & ~n1257;
  assign n1259 = ~n1232 & ~n1258;
  assign n1260 = reg_controllable_hmaster2_out & ~n1259;
  assign n1261 = ~reg_stateG10_1_out & ~n757;
  assign n1262 = ~reg_stateG10_1_out & ~n1261;
  assign n1263 = reg_controllable_hgrant1_out & ~n1262;
  assign n1264 = ~n1174 & ~n1263;
  assign n1265 = next_sys_fair<0>_out  & ~n1264;
  assign n1266 = ~n1176 & ~n1265;
  assign n1267 = next_sys_fair<1>_out  & ~n1266;
  assign n1268 = ~reg_stateG10_1_out & ~n923;
  assign n1269 = ~reg_stateG10_1_out & ~n1268;
  assign n1270 = reg_controllable_hgrant1_out & ~n1269;
  assign n1271 = ~reg_controllable_hgrant1_out & ~n921;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = next_sys_fair<0>_out  & ~n1272;
  assign n1274 = ~n1206 & ~n1273;
  assign n1275 = ~next_sys_fair<1>_out  & ~n1274;
  assign n1276 = ~n1267 & ~n1275;
  assign n1277 = ~reg_controllable_hmaster2_out & ~n1276;
  assign n1278 = ~n1260 & ~n1277;
  assign n1279 = reg_controllable_hmaster1_out & ~n1278;
  assign n1280 = ~reg_stateG10_1_out & ~n835;
  assign n1281 = ~reg_stateG10_1_out & ~n1280;
  assign n1282 = reg_controllable_hgrant1_out & ~n1281;
  assign n1283 = ~n1182 & ~n1282;
  assign n1284 = next_sys_fair<0>_out  & ~n1283;
  assign n1285 = ~n1195 & ~n1284;
  assign n1286 = next_sys_fair<1>_out  & ~n1285;
  assign n1287 = ~reg_stateG10_1_out & ~n948;
  assign n1288 = ~reg_stateG10_1_out & ~n1287;
  assign n1289 = reg_controllable_hgrant1_out & ~n1288;
  assign n1290 = ~n1271 & ~n1289;
  assign n1291 = next_sys_fair<0>_out  & ~n1290;
  assign n1292 = ~reg_stateG10_1_out & ~n958;
  assign n1293 = ~reg_stateG10_1_out & ~n1292;
  assign n1294 = reg_controllable_hgrant1_out & ~n1293;
  assign n1295 = ~n1182 & ~n1294;
  assign n1296 = ~next_sys_fair<0>_out  & ~n1295;
  assign n1297 = ~n1291 & ~n1296;
  assign n1298 = ~next_sys_fair<1>_out  & ~n1297;
  assign n1299 = ~n1286 & ~n1298;
  assign n1300 = ~reg_controllable_hmaster2_out & ~n1299;
  assign n1301 = ~n1260 & ~n1300;
  assign n1302 = ~reg_controllable_hmaster1_out & ~n1301;
  assign n1303 = ~n1279 & ~n1302;
  assign n1304 = reg_controllable_hmaster0_out & ~n1303;
  assign n1305 = reg_controllable_hmaster2_out & ~n1276;
  assign n1306 = ~n1206 & ~n1265;
  assign n1307 = next_sys_fair<1>_out  & ~n1306;
  assign n1308 = ~n1275 & ~n1307;
  assign n1309 = ~reg_controllable_hmaster2_out & ~n1308;
  assign n1310 = ~n1305 & ~n1309;
  assign n1311 = ~reg_controllable_hmaster1_out & ~n1310;
  assign n1312 = ~n1279 & ~n1311;
  assign n1313 = ~reg_controllable_hmaster0_out & ~n1312;
  assign n1314 = ~n1304 & ~n1313;
  assign n1315 = ~next_sys_fair<2>_out  & ~n1314;
  assign n1316 = ~n1225 & ~n1315;
  assign n1317 = ~reg_controllable_hgrant2_out & ~n1316;
  assign n1318 = ~n1129 & ~n1317;
  assign n1319 = ~reg_controllable_hgrant3_out & ~n1318;
  assign n1320 = ~n1080 & ~n1319;
  assign n1321 = ~reg_controllable_hgrant4_out & ~n1320;
  assign n1322 = ~n982 & ~n1321;
  assign n1323 = reg_controllable_nhgrant0_out & ~n1322;
  assign n1324 = ~next_sys_fair<1>_out  & ~n742;
  assign n1325 = ~n985 & ~n1324;
  assign n1326 = reg_controllable_hmaster2_out & ~n1325;
  assign n1327 = ~next_sys_fair<1>_out  & ~n1047;
  assign n1328 = ~n1003 & ~n1327;
  assign n1329 = ~reg_controllable_hmaster2_out & ~n1328;
  assign n1330 = ~n1326 & ~n1329;
  assign n1331 = reg_controllable_hmaster1_out & ~n1330;
  assign n1332 = ~next_sys_fair<1>_out  & ~n805;
  assign n1333 = ~n1003 & ~n1332;
  assign n1334 = ~reg_controllable_hmaster2_out & ~n1333;
  assign n1335 = ~n1326 & ~n1334;
  assign n1336 = ~reg_controllable_hmaster1_out & ~n1335;
  assign n1337 = ~n1331 & ~n1336;
  assign n1338 = reg_controllable_hmaster0_out & ~n1337;
  assign n1339 = ~next_sys_fair<1>_out  & ~n1065;
  assign n1340 = ~n1003 & ~n1339;
  assign n1341 = ~reg_controllable_hmaster2_out & ~n1340;
  assign n1342 = ~n1326 & ~n1341;
  assign n1343 = reg_controllable_hmaster1_out & ~n1342;
  assign n1344 = ~n1021 & ~n1332;
  assign n1345 = reg_controllable_hmaster2_out & ~n1344;
  assign n1346 = ~next_sys_fair<1>_out  & ~n850;
  assign n1347 = ~n993 & ~n1346;
  assign n1348 = ~reg_controllable_hmaster2_out & ~n1347;
  assign n1349 = ~n1345 & ~n1348;
  assign n1350 = ~reg_controllable_hmaster1_out & ~n1349;
  assign n1351 = ~n1343 & ~n1350;
  assign n1352 = ~reg_controllable_hmaster0_out & ~n1351;
  assign n1353 = ~n1338 & ~n1352;
  assign n1354 = next_sys_fair<2>_out  & ~n1353;
  assign n1355 = next_sys_fair<1>_out  & ~n1083;
  assign n1356 = ~n1034 & ~n1355;
  assign n1357 = reg_controllable_hmaster2_out & ~n1356;
  assign n1358 = next_sys_fair<1>_out  & ~n1094;
  assign n1359 = ~n1051 & ~n1358;
  assign n1360 = ~reg_controllable_hmaster2_out & ~n1359;
  assign n1361 = ~n1357 & ~n1360;
  assign n1362 = reg_controllable_hmaster1_out & ~n1361;
  assign n1363 = next_sys_fair<1>_out  & ~n1088;
  assign n1364 = ~n1051 & ~n1363;
  assign n1365 = ~reg_controllable_hmaster2_out & ~n1364;
  assign n1366 = ~n1357 & ~n1365;
  assign n1367 = ~reg_controllable_hmaster1_out & ~n1366;
  assign n1368 = ~n1362 & ~n1367;
  assign n1369 = reg_controllable_hmaster0_out & ~n1368;
  assign n1370 = reg_controllable_hmaster2_out & ~n1359;
  assign n1371 = next_sys_fair<1>_out  & ~n1104;
  assign n1372 = ~n1041 & ~n1371;
  assign n1373 = ~reg_controllable_hmaster2_out & ~n1372;
  assign n1374 = ~n1370 & ~n1373;
  assign n1375 = ~reg_controllable_hmaster1_out & ~n1374;
  assign n1376 = ~n1362 & ~n1375;
  assign n1377 = ~reg_controllable_hmaster0_out & ~n1376;
  assign n1378 = ~n1369 & ~n1377;
  assign n1379 = ~next_sys_fair<2>_out  & ~n1378;
  assign n1380 = ~n1354 & ~n1379;
  assign n1381 = ~reg_controllable_hgrant2_out & ~n1380;
  assign n1382 = ~reg_controllable_hgrant2_out & ~n1381;
  assign n1383 = ~reg_controllable_hgrant3_out & ~n1382;
  assign n1384 = ~reg_controllable_hgrant3_out & ~n1383;
  assign n1385 = ~reg_controllable_hgrant4_out & ~n1384;
  assign n1386 = ~reg_controllable_hgrant4_out & ~n1385;
  assign n1387 = ~reg_controllable_nhgrant0_out & ~n1386;
  assign n1388 = ~n1323 & ~n1387;
  assign n1389 = ~reg_i_hready_out & ~n1388;
  assign n1390 = ~n691 & ~n1389;
  assign n1391 = ~next_sys_fair<3>_out  & ~n1390;
  assign n1392 = ~n167 & ~n1391;
  assign n1393 = reg_controllable_ndecide_out & ~n1392;
  assign n1394 = reg_controllable_hmaster2_out & ~n79;
  assign n1395 = reg_controllable_hmaster2_out & ~n1394;
  assign n1396 = reg_controllable_hmaster0_out & ~n1395;
  assign n1397 = reg_controllable_hmaster1_out & ~n1395;
  assign n1398 = reg_controllable_hmaster1_out & ~n1397;
  assign n1399 = ~reg_controllable_hmaster0_out & ~n1398;
  assign n1400 = ~n1396 & ~n1399;
  assign n1401 = ~reg_i_hready_out & ~n1400;
  assign n1402 = ~n127 & ~n1401;
  assign n1403 = next_sys_fair<3>_out  & ~n1402;
  assign n1404 = ~reg_controllable_locked_out & ~n185;
  assign n1405 = ~reg_controllable_hgrant1_out & ~n1404;
  assign n1406 = ~reg_controllable_hgrant1_out & ~n1405;
  assign n1407 = reg_stateG10_4_out & ~n1406;
  assign n1408 = ~n189 & ~n1407;
  assign n1409 = reg_i_hlock4_out & ~n1408;
  assign n1410 = ~reg_i_hlock4_out & ~n1406;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~next_sys_fair<0>_out  & ~n1411;
  assign n1413 = ~next_sys_fair<0>_out  & ~n1412;
  assign n1414 = next_sys_fair<1>_out  & ~n1413;
  assign n1415 = ~fair_cnt<2>_out  & ~n183;
  assign n1416 = ~reg_controllable_locked_out & ~n1415;
  assign n1417 = ~reg_controllable_locked_out & ~n1416;
  assign n1418 = ~reg_controllable_hgrant1_out & ~n1417;
  assign n1419 = ~reg_controllable_hgrant1_out & ~n1418;
  assign n1420 = reg_stateG10_4_out & ~n1419;
  assign n1421 = ~n196 & ~n1416;
  assign n1422 = ~reg_controllable_hgrant1_out & ~n1421;
  assign n1423 = ~reg_controllable_hgrant1_out & ~n1422;
  assign n1424 = ~reg_stateG10_4_out & ~n1423;
  assign n1425 = ~n1420 & ~n1424;
  assign n1426 = reg_i_hlock4_out & ~n1425;
  assign n1427 = ~reg_i_hlock4_out & ~n1419;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = ~next_sys_fair<1>_out  & ~n1428;
  assign n1430 = ~n1414 & ~n1429;
  assign n1431 = reg_controllable_hmaster0_out & ~n1430;
  assign n1432 = reg_controllable_hmaster1_out & ~n1430;
  assign n1433 = ~fair_cnt<0>_out  & ~n272;
  assign n1434 = ~fair_cnt<0>_out  & ~n1433;
  assign n1435 = ~fair_cnt<1>_out  & ~n1434;
  assign n1436 = ~fair_cnt<1>_out  & ~n1435;
  assign n1437 = fair_cnt<2>_out  & ~n1436;
  assign n1438 = ~fair_cnt<2>_out  & ~n272;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = reg_controllable_hmastlock_out & ~n1439;
  assign n1441 = reg_controllable_hmastlock_out & ~n1440;
  assign n1442 = reg_controllable_locked_out & ~n1441;
  assign n1443 = ~reg_controllable_hmastlock_out & ~n779;
  assign n1444 = ~n232 & ~n1443;
  assign n1445 = ~reg_controllable_locked_out & ~n1444;
  assign n1446 = ~n1442 & ~n1445;
  assign n1447 = ~reg_controllable_hgrant1_out & ~n1446;
  assign n1448 = ~reg_controllable_hgrant1_out & ~n1447;
  assign n1449 = reg_stateG10_4_out & ~n1448;
  assign n1450 = ~n231 & ~n1445;
  assign n1451 = ~reg_controllable_hgrant1_out & ~n1450;
  assign n1452 = ~reg_controllable_hgrant1_out & ~n1451;
  assign n1453 = ~reg_stateG10_4_out & ~n1452;
  assign n1454 = ~n1449 & ~n1453;
  assign n1455 = reg_i_hlock4_out & ~n1454;
  assign n1456 = reg_controllable_hmastlock_out & ~n832;
  assign n1457 = reg_controllable_locked_out & ~n1456;
  assign n1458 = ~reg_controllable_hmastlock_out & ~n1439;
  assign n1459 = ~n232 & ~n1458;
  assign n1460 = ~reg_controllable_locked_out & ~n1459;
  assign n1461 = ~n1457 & ~n1460;
  assign n1462 = ~reg_controllable_hgrant1_out & ~n1461;
  assign n1463 = ~reg_controllable_hgrant1_out & ~n1462;
  assign n1464 = reg_stateG10_4_out & ~n1463;
  assign n1465 = ~n235 & ~n1457;
  assign n1466 = ~reg_controllable_hgrant1_out & ~n1465;
  assign n1467 = ~reg_controllable_hgrant1_out & ~n1466;
  assign n1468 = ~reg_stateG10_4_out & ~n1467;
  assign n1469 = ~n1464 & ~n1468;
  assign n1470 = ~reg_i_hlock4_out & ~n1469;
  assign n1471 = ~n1455 & ~n1470;
  assign n1472 = ~next_sys_fair<0>_out  & ~n1471;
  assign n1473 = ~next_sys_fair<0>_out  & ~n1472;
  assign n1474 = next_sys_fair<1>_out  & ~n1473;
  assign n1475 = fair_cnt<0>_out  & ~n129;
  assign n1476 = ~n1433 & ~n1475;
  assign n1477 = fair_cnt<1>_out  & ~n1476;
  assign n1478 = ~fair_cnt<1>_out  & ~n272;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = next_env_fair_out & ~n1479;
  assign n1481 = ~next_env_fair_out & ~n272;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~fair_cnt<2>_out  & ~n1482;
  assign n1484 = ~fair_cnt<2>_out  & ~n1483;
  assign n1485 = reg_controllable_hmastlock_out & ~n1484;
  assign n1486 = reg_controllable_hmastlock_out & ~n1485;
  assign n1487 = reg_controllable_locked_out & ~n1486;
  assign n1488 = reg_controllable_hmastlock_out & ~n1415;
  assign n1489 = ~reg_controllable_hmastlock_out & ~n755;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~reg_controllable_locked_out & ~n1490;
  assign n1492 = ~n1487 & ~n1491;
  assign n1493 = ~reg_controllable_hgrant1_out & ~n1492;
  assign n1494 = ~reg_controllable_hgrant1_out & ~n1493;
  assign n1495 = reg_stateG10_4_out & ~n1494;
  assign n1496 = ~n254 & ~n1475;
  assign n1497 = fair_cnt<1>_out  & ~n1496;
  assign n1498 = ~n267 & ~n1497;
  assign n1499 = next_env_fair_out & ~n1498;
  assign n1500 = ~n277 & ~n1499;
  assign n1501 = ~fair_cnt<2>_out  & ~n1500;
  assign n1502 = ~fair_cnt<2>_out  & ~n1501;
  assign n1503 = reg_controllable_hmastlock_out & ~n1502;
  assign n1504 = ~n282 & ~n1503;
  assign n1505 = reg_controllable_locked_out & ~n1504;
  assign n1506 = ~n1491 & ~n1505;
  assign n1507 = ~reg_controllable_hgrant1_out & ~n1506;
  assign n1508 = ~reg_controllable_hgrant1_out & ~n1507;
  assign n1509 = ~reg_stateG10_4_out & ~n1508;
  assign n1510 = ~n1495 & ~n1509;
  assign n1511 = reg_i_hlock4_out & ~n1510;
  assign n1512 = reg_controllable_hmastlock_out & ~n755;
  assign n1513 = reg_controllable_hmastlock_out & ~n1512;
  assign n1514 = reg_controllable_locked_out & ~n1513;
  assign n1515 = ~reg_controllable_hmastlock_out & ~n1484;
  assign n1516 = ~n1488 & ~n1515;
  assign n1517 = ~reg_controllable_locked_out & ~n1516;
  assign n1518 = ~n1514 & ~n1517;
  assign n1519 = ~reg_controllable_hgrant1_out & ~n1518;
  assign n1520 = ~reg_controllable_hgrant1_out & ~n1519;
  assign n1521 = reg_stateG10_4_out & ~n1520;
  assign n1522 = ~reg_controllable_hmastlock_out & ~n1502;
  assign n1523 = ~n1488 & ~n1522;
  assign n1524 = ~reg_controllable_locked_out & ~n1523;
  assign n1525 = ~n1514 & ~n1524;
  assign n1526 = ~reg_controllable_hgrant1_out & ~n1525;
  assign n1527 = ~reg_controllable_hgrant1_out & ~n1526;
  assign n1528 = ~reg_stateG10_4_out & ~n1527;
  assign n1529 = ~n1521 & ~n1528;
  assign n1530 = ~reg_i_hlock4_out & ~n1529;
  assign n1531 = ~n1511 & ~n1530;
  assign n1532 = ~next_sys_fair<1>_out  & ~n1531;
  assign n1533 = ~n1474 & ~n1532;
  assign n1534 = reg_controllable_hmaster2_out & ~n1533;
  assign n1535 = ~reg_controllable_hmaster2_out & ~n1430;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~reg_controllable_hmaster1_out & ~n1536;
  assign n1538 = ~n1432 & ~n1537;
  assign n1539 = ~reg_controllable_hmaster0_out & ~n1538;
  assign n1540 = ~n1431 & ~n1539;
  assign n1541 = next_sys_fair<2>_out  & ~n1540;
  assign n1542 = next_sys_fair<1>_out  & ~n1428;
  assign n1543 = ~next_sys_fair<1>_out  & ~n1411;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = reg_controllable_hmaster0_out & ~n1544;
  assign n1546 = reg_controllable_hmaster1_out & ~n1544;
  assign n1547 = next_sys_fair<1>_out  & ~n1531;
  assign n1548 = ~n316 & ~n1438;
  assign n1549 = reg_controllable_hmastlock_out & ~n1548;
  assign n1550 = reg_controllable_hmastlock_out & ~n1549;
  assign n1551 = reg_controllable_locked_out & ~n1550;
  assign n1552 = ~reg_controllable_hmastlock_out & ~n921;
  assign n1553 = ~n232 & ~n1552;
  assign n1554 = ~reg_controllable_locked_out & ~n1553;
  assign n1555 = ~n1551 & ~n1554;
  assign n1556 = ~reg_controllable_hgrant1_out & ~n1555;
  assign n1557 = ~reg_controllable_hgrant1_out & ~n1556;
  assign n1558 = reg_stateG10_4_out & ~n1557;
  assign n1559 = ~n321 & ~n1554;
  assign n1560 = ~reg_controllable_hgrant1_out & ~n1559;
  assign n1561 = ~reg_controllable_hgrant1_out & ~n1560;
  assign n1562 = ~reg_stateG10_4_out & ~n1561;
  assign n1563 = ~n1558 & ~n1562;
  assign n1564 = reg_i_hlock4_out & ~n1563;
  assign n1565 = reg_controllable_hmastlock_out & ~n945;
  assign n1566 = reg_controllable_locked_out & ~n1565;
  assign n1567 = ~reg_controllable_hmastlock_out & ~n1548;
  assign n1568 = ~n232 & ~n1567;
  assign n1569 = ~reg_controllable_locked_out & ~n1568;
  assign n1570 = ~n1566 & ~n1569;
  assign n1571 = ~reg_controllable_hgrant1_out & ~n1570;
  assign n1572 = ~reg_controllable_hgrant1_out & ~n1571;
  assign n1573 = reg_stateG10_4_out & ~n1572;
  assign n1574 = ~n324 & ~n1566;
  assign n1575 = ~reg_controllable_hgrant1_out & ~n1574;
  assign n1576 = ~reg_controllable_hgrant1_out & ~n1575;
  assign n1577 = ~reg_stateG10_4_out & ~n1576;
  assign n1578 = ~n1573 & ~n1577;
  assign n1579 = ~reg_i_hlock4_out & ~n1578;
  assign n1580 = ~n1564 & ~n1579;
  assign n1581 = next_sys_fair<0>_out  & ~n1580;
  assign n1582 = ~next_env_fair_out & ~n1436;
  assign n1583 = ~n898 & ~n1582;
  assign n1584 = fair_cnt<2>_out  & ~n1583;
  assign n1585 = ~n1438 & ~n1584;
  assign n1586 = reg_controllable_hmastlock_out & ~n1585;
  assign n1587 = reg_controllable_hmastlock_out & ~n1586;
  assign n1588 = reg_controllable_locked_out & ~n1587;
  assign n1589 = ~n1445 & ~n1588;
  assign n1590 = ~reg_controllable_hgrant1_out & ~n1589;
  assign n1591 = ~reg_controllable_hgrant1_out & ~n1590;
  assign n1592 = reg_stateG10_4_out & ~n1591;
  assign n1593 = ~n342 & ~n1445;
  assign n1594 = ~reg_controllable_hgrant1_out & ~n1593;
  assign n1595 = ~reg_controllable_hgrant1_out & ~n1594;
  assign n1596 = ~reg_stateG10_4_out & ~n1595;
  assign n1597 = ~n1592 & ~n1596;
  assign n1598 = reg_i_hlock4_out & ~n1597;
  assign n1599 = ~reg_controllable_hmastlock_out & ~n1585;
  assign n1600 = ~n232 & ~n1599;
  assign n1601 = ~reg_controllable_locked_out & ~n1600;
  assign n1602 = ~n1457 & ~n1601;
  assign n1603 = ~reg_controllable_hgrant1_out & ~n1602;
  assign n1604 = ~reg_controllable_hgrant1_out & ~n1603;
  assign n1605 = reg_stateG10_4_out & ~n1604;
  assign n1606 = ~n345 & ~n1457;
  assign n1607 = ~reg_controllable_hgrant1_out & ~n1606;
  assign n1608 = ~reg_controllable_hgrant1_out & ~n1607;
  assign n1609 = ~reg_stateG10_4_out & ~n1608;
  assign n1610 = ~n1605 & ~n1609;
  assign n1611 = ~reg_i_hlock4_out & ~n1610;
  assign n1612 = ~n1598 & ~n1611;
  assign n1613 = ~next_sys_fair<0>_out  & ~n1612;
  assign n1614 = ~n1581 & ~n1613;
  assign n1615 = ~next_sys_fair<1>_out  & ~n1614;
  assign n1616 = ~n1547 & ~n1615;
  assign n1617 = reg_controllable_hmaster2_out & ~n1616;
  assign n1618 = ~reg_controllable_hmaster2_out & ~n1544;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~reg_controllable_hmaster1_out & ~n1619;
  assign n1621 = ~n1546 & ~n1620;
  assign n1622 = ~reg_controllable_hmaster0_out & ~n1621;
  assign n1623 = ~n1545 & ~n1622;
  assign n1624 = ~next_sys_fair<2>_out  & ~n1623;
  assign n1625 = ~n1541 & ~n1624;
  assign n1626 = ~reg_controllable_hgrant2_out & ~n1625;
  assign n1627 = ~reg_controllable_hgrant2_out & ~n1626;
  assign n1628 = ~reg_controllable_hgrant3_out & ~n1627;
  assign n1629 = ~reg_controllable_hgrant3_out & ~n1628;
  assign n1630 = reg_controllable_hgrant4_out & ~n1629;
  assign n1631 = ~next_sys_fair<0>_out  & ~n1419;
  assign n1632 = ~next_sys_fair<0>_out  & ~n1631;
  assign n1633 = next_sys_fair<1>_out  & ~n1632;
  assign n1634 = next_sys_fair<0>_out  & ~n1406;
  assign n1635 = ~n1631 & ~n1634;
  assign n1636 = ~next_sys_fair<1>_out  & ~n1635;
  assign n1637 = ~n1633 & ~n1636;
  assign n1638 = reg_controllable_hmaster2_out & ~n1637;
  assign n1639 = ~next_sys_fair<0>_out  & ~n1494;
  assign n1640 = ~next_sys_fair<0>_out  & ~n1639;
  assign n1641 = next_sys_fair<1>_out  & ~n1640;
  assign n1642 = next_sys_fair<0>_out  & ~n1448;
  assign n1643 = ~n1639 & ~n1642;
  assign n1644 = ~next_sys_fair<1>_out  & ~n1643;
  assign n1645 = ~n1641 & ~n1644;
  assign n1646 = ~reg_controllable_hmaster2_out & ~n1645;
  assign n1647 = ~n1638 & ~n1646;
  assign n1648 = reg_controllable_hmaster1_out & ~n1647;
  assign n1649 = ~reg_controllable_hmaster1_out & ~n1637;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = reg_controllable_hmaster0_out & ~n1650;
  assign n1652 = ~reg_controllable_hmaster0_out & ~n1637;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = next_sys_fair<2>_out  & ~n1653;
  assign n1655 = next_sys_fair<1>_out  & ~n1419;
  assign n1656 = ~next_sys_fair<1>_out  & ~n1406;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = reg_controllable_hmaster2_out & ~n1657;
  assign n1659 = next_sys_fair<1>_out  & ~n1494;
  assign n1660 = next_sys_fair<0>_out  & ~n1557;
  assign n1661 = ~next_sys_fair<0>_out  & ~n1591;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = ~next_sys_fair<1>_out  & ~n1662;
  assign n1664 = ~n1659 & ~n1663;
  assign n1665 = ~reg_controllable_hmaster2_out & ~n1664;
  assign n1666 = ~n1658 & ~n1665;
  assign n1667 = reg_controllable_hmaster1_out & ~n1666;
  assign n1668 = ~reg_controllable_hmaster1_out & ~n1657;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = reg_controllable_hmaster0_out & ~n1669;
  assign n1671 = ~reg_controllable_hmaster0_out & ~n1657;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~next_sys_fair<2>_out  & ~n1672;
  assign n1674 = ~n1654 & ~n1673;
  assign n1675 = reg_stateG10_3_out & ~n1674;
  assign n1676 = ~next_sys_fair<0>_out  & ~n1423;
  assign n1677 = ~next_sys_fair<0>_out  & ~n1676;
  assign n1678 = next_sys_fair<1>_out  & ~n1677;
  assign n1679 = ~n372 & ~n1676;
  assign n1680 = ~next_sys_fair<1>_out  & ~n1679;
  assign n1681 = ~n1678 & ~n1680;
  assign n1682 = reg_controllable_hmaster2_out & ~n1681;
  assign n1683 = ~next_sys_fair<0>_out  & ~n1508;
  assign n1684 = ~next_sys_fair<0>_out  & ~n1683;
  assign n1685 = next_sys_fair<1>_out  & ~n1684;
  assign n1686 = next_sys_fair<0>_out  & ~n1452;
  assign n1687 = ~n1683 & ~n1686;
  assign n1688 = ~next_sys_fair<1>_out  & ~n1687;
  assign n1689 = ~n1685 & ~n1688;
  assign n1690 = ~reg_controllable_hmaster2_out & ~n1689;
  assign n1691 = ~n1682 & ~n1690;
  assign n1692 = reg_controllable_hmaster1_out & ~n1691;
  assign n1693 = ~reg_controllable_hmaster1_out & ~n1681;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = reg_controllable_hmaster0_out & ~n1694;
  assign n1696 = ~reg_controllable_hmaster0_out & ~n1681;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = next_sys_fair<2>_out  & ~n1697;
  assign n1699 = next_sys_fair<1>_out  & ~n1423;
  assign n1700 = ~n394 & ~n1699;
  assign n1701 = reg_controllable_hmaster2_out & ~n1700;
  assign n1702 = next_sys_fair<1>_out  & ~n1508;
  assign n1703 = next_sys_fair<0>_out  & ~n1561;
  assign n1704 = ~next_sys_fair<0>_out  & ~n1595;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~next_sys_fair<1>_out  & ~n1705;
  assign n1707 = ~n1702 & ~n1706;
  assign n1708 = ~reg_controllable_hmaster2_out & ~n1707;
  assign n1709 = ~n1701 & ~n1708;
  assign n1710 = reg_controllable_hmaster1_out & ~n1709;
  assign n1711 = ~reg_controllable_hmaster1_out & ~n1700;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = reg_controllable_hmaster0_out & ~n1712;
  assign n1714 = ~reg_controllable_hmaster0_out & ~n1700;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~next_sys_fair<2>_out  & ~n1715;
  assign n1717 = ~n1698 & ~n1716;
  assign n1718 = ~reg_stateG10_3_out & ~n1717;
  assign n1719 = ~n1675 & ~n1718;
  assign n1720 = ~reg_controllable_hgrant2_out & ~n1719;
  assign n1721 = ~reg_controllable_hgrant2_out & ~n1720;
  assign n1722 = reg_i_hlock3_out & ~n1721;
  assign n1723 = ~next_sys_fair<0>_out  & ~n1520;
  assign n1724 = ~next_sys_fair<0>_out  & ~n1723;
  assign n1725 = next_sys_fair<1>_out  & ~n1724;
  assign n1726 = next_sys_fair<0>_out  & ~n1463;
  assign n1727 = ~n1723 & ~n1726;
  assign n1728 = ~next_sys_fair<1>_out  & ~n1727;
  assign n1729 = ~n1725 & ~n1728;
  assign n1730 = ~reg_controllable_hmaster2_out & ~n1729;
  assign n1731 = ~n1638 & ~n1730;
  assign n1732 = reg_controllable_hmaster1_out & ~n1731;
  assign n1733 = ~n1649 & ~n1732;
  assign n1734 = reg_controllable_hmaster0_out & ~n1733;
  assign n1735 = ~n1652 & ~n1734;
  assign n1736 = next_sys_fair<2>_out  & ~n1735;
  assign n1737 = next_sys_fair<1>_out  & ~n1520;
  assign n1738 = next_sys_fair<0>_out  & ~n1572;
  assign n1739 = ~next_sys_fair<0>_out  & ~n1604;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = ~next_sys_fair<1>_out  & ~n1740;
  assign n1742 = ~n1737 & ~n1741;
  assign n1743 = ~reg_controllable_hmaster2_out & ~n1742;
  assign n1744 = ~n1658 & ~n1743;
  assign n1745 = reg_controllable_hmaster1_out & ~n1744;
  assign n1746 = ~n1668 & ~n1745;
  assign n1747 = reg_controllable_hmaster0_out & ~n1746;
  assign n1748 = ~n1671 & ~n1747;
  assign n1749 = ~next_sys_fair<2>_out  & ~n1748;
  assign n1750 = ~n1736 & ~n1749;
  assign n1751 = reg_stateG10_3_out & ~n1750;
  assign n1752 = ~next_sys_fair<0>_out  & ~n1527;
  assign n1753 = ~next_sys_fair<0>_out  & ~n1752;
  assign n1754 = next_sys_fair<1>_out  & ~n1753;
  assign n1755 = next_sys_fair<0>_out  & ~n1467;
  assign n1756 = ~n1752 & ~n1755;
  assign n1757 = ~next_sys_fair<1>_out  & ~n1756;
  assign n1758 = ~n1754 & ~n1757;
  assign n1759 = ~reg_controllable_hmaster2_out & ~n1758;
  assign n1760 = ~n1638 & ~n1759;
  assign n1761 = reg_controllable_hmaster1_out & ~n1760;
  assign n1762 = ~n1649 & ~n1761;
  assign n1763 = reg_controllable_hmaster0_out & ~n1762;
  assign n1764 = ~n1652 & ~n1763;
  assign n1765 = next_sys_fair<2>_out  & ~n1764;
  assign n1766 = next_sys_fair<1>_out  & ~n1527;
  assign n1767 = next_sys_fair<0>_out  & ~n1576;
  assign n1768 = ~next_sys_fair<0>_out  & ~n1608;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = ~next_sys_fair<1>_out  & ~n1769;
  assign n1771 = ~n1766 & ~n1770;
  assign n1772 = ~reg_controllable_hmaster2_out & ~n1771;
  assign n1773 = ~n1658 & ~n1772;
  assign n1774 = reg_controllable_hmaster1_out & ~n1773;
  assign n1775 = ~n1668 & ~n1774;
  assign n1776 = reg_controllable_hmaster0_out & ~n1775;
  assign n1777 = ~n1671 & ~n1776;
  assign n1778 = ~next_sys_fair<2>_out  & ~n1777;
  assign n1779 = ~n1765 & ~n1778;
  assign n1780 = ~reg_stateG10_3_out & ~n1779;
  assign n1781 = ~n1751 & ~n1780;
  assign n1782 = ~reg_controllable_hgrant2_out & ~n1781;
  assign n1783 = ~reg_controllable_hgrant2_out & ~n1782;
  assign n1784 = ~reg_i_hlock3_out & ~n1783;
  assign n1785 = ~n1722 & ~n1784;
  assign n1786 = reg_controllable_hgrant3_out & ~n1785;
  assign n1787 = next_sys_fair<0>_out  & ~n1419;
  assign n1788 = ~next_sys_fair<0>_out  & ~n1406;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~next_sys_fair<1>_out  & ~n1789;
  assign n1791 = ~n1633 & ~n1790;
  assign n1792 = reg_controllable_hmaster0_out & ~n1791;
  assign n1793 = reg_controllable_hmaster2_out & ~n1791;
  assign n1794 = next_sys_fair<0>_out  & ~n1494;
  assign n1795 = ~next_sys_fair<0>_out  & ~n1448;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~next_sys_fair<1>_out  & ~n1796;
  assign n1798 = ~n1641 & ~n1797;
  assign n1799 = ~reg_controllable_hmaster2_out & ~n1798;
  assign n1800 = ~n1793 & ~n1799;
  assign n1801 = reg_controllable_hmaster1_out & ~n1800;
  assign n1802 = ~reg_controllable_hmaster1_out & ~n1791;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = ~reg_controllable_hmaster0_out & ~n1803;
  assign n1805 = ~n1792 & ~n1804;
  assign n1806 = reg_stateG10_2_out & ~n1805;
  assign n1807 = next_sys_fair<0>_out  & ~n1423;
  assign n1808 = ~n419 & ~n1807;
  assign n1809 = ~next_sys_fair<1>_out  & ~n1808;
  assign n1810 = ~n1678 & ~n1809;
  assign n1811 = reg_controllable_hmaster0_out & ~n1810;
  assign n1812 = reg_controllable_hmaster2_out & ~n1810;
  assign n1813 = next_sys_fair<0>_out  & ~n1508;
  assign n1814 = ~next_sys_fair<0>_out  & ~n1452;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~next_sys_fair<1>_out  & ~n1815;
  assign n1817 = ~n1685 & ~n1816;
  assign n1818 = ~reg_controllable_hmaster2_out & ~n1817;
  assign n1819 = ~n1812 & ~n1818;
  assign n1820 = reg_controllable_hmaster1_out & ~n1819;
  assign n1821 = ~reg_controllable_hmaster1_out & ~n1810;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~reg_controllable_hmaster0_out & ~n1822;
  assign n1824 = ~n1811 & ~n1823;
  assign n1825 = ~reg_stateG10_2_out & ~n1824;
  assign n1826 = ~n1806 & ~n1825;
  assign n1827 = reg_i_hlock2_out & ~n1826;
  assign n1828 = next_sys_fair<0>_out  & ~n1520;
  assign n1829 = ~next_sys_fair<0>_out  & ~n1463;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~next_sys_fair<1>_out  & ~n1830;
  assign n1832 = ~n1725 & ~n1831;
  assign n1833 = ~reg_controllable_hmaster2_out & ~n1832;
  assign n1834 = ~n1793 & ~n1833;
  assign n1835 = reg_controllable_hmaster1_out & ~n1834;
  assign n1836 = ~n1802 & ~n1835;
  assign n1837 = ~reg_controllable_hmaster0_out & ~n1836;
  assign n1838 = ~n1792 & ~n1837;
  assign n1839 = reg_stateG10_2_out & ~n1838;
  assign n1840 = next_sys_fair<0>_out  & ~n1527;
  assign n1841 = ~next_sys_fair<0>_out  & ~n1467;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~next_sys_fair<1>_out  & ~n1842;
  assign n1844 = ~n1754 & ~n1843;
  assign n1845 = ~reg_controllable_hmaster2_out & ~n1844;
  assign n1846 = ~n1793 & ~n1845;
  assign n1847 = reg_controllable_hmaster1_out & ~n1846;
  assign n1848 = ~n1802 & ~n1847;
  assign n1849 = ~reg_controllable_hmaster0_out & ~n1848;
  assign n1850 = ~n1792 & ~n1849;
  assign n1851 = ~reg_stateG10_2_out & ~n1850;
  assign n1852 = ~n1839 & ~n1851;
  assign n1853 = ~reg_i_hlock2_out & ~n1852;
  assign n1854 = ~n1827 & ~n1853;
  assign n1855 = next_sys_fair<2>_out  & ~n1854;
  assign n1856 = reg_controllable_hmaster0_out & ~n1657;
  assign n1857 = ~reg_controllable_hmaster0_out & ~n1669;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = reg_stateG10_2_out & ~n1858;
  assign n1860 = reg_controllable_hmaster0_out & ~n1700;
  assign n1861 = ~reg_controllable_hmaster0_out & ~n1712;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = ~reg_stateG10_2_out & ~n1862;
  assign n1864 = ~n1859 & ~n1863;
  assign n1865 = reg_i_hlock2_out & ~n1864;
  assign n1866 = ~reg_controllable_hmaster0_out & ~n1746;
  assign n1867 = ~n1856 & ~n1866;
  assign n1868 = reg_stateG10_2_out & ~n1867;
  assign n1869 = ~reg_controllable_hmaster0_out & ~n1775;
  assign n1870 = ~n1856 & ~n1869;
  assign n1871 = ~reg_stateG10_2_out & ~n1870;
  assign n1872 = ~n1868 & ~n1871;
  assign n1873 = ~reg_i_hlock2_out & ~n1872;
  assign n1874 = ~n1865 & ~n1873;
  assign n1875 = ~next_sys_fair<2>_out  & ~n1874;
  assign n1876 = ~n1855 & ~n1875;
  assign n1877 = reg_controllable_hgrant2_out & ~n1876;
  assign n1878 = reg_stateG10_1_out & ~n1417;
  assign n1879 = reg_i_hlock1_out & ~n1421;
  assign n1880 = ~reg_i_hlock1_out & ~n1417;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~reg_stateG10_1_out & ~n1881;
  assign n1883 = ~n1878 & ~n1882;
  assign n1884 = reg_controllable_hgrant1_out & ~n1883;
  assign n1885 = ~n77 & ~n562;
  assign n1886 = reg_controllable_hmastlock_out & ~n1885;
  assign n1887 = ~n486 & ~n1886;
  assign n1888 = reg_controllable_locked_out & ~n1887;
  assign n1889 = ~n95 & ~n183;
  assign n1890 = reg_controllable_hmastlock_out & ~n1889;
  assign n1891 = ~reg_controllable_hmastlock_out & ~n1885;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = ~reg_controllable_locked_out & ~n1892;
  assign n1894 = ~n1888 & ~n1893;
  assign n1895 = ~reg_controllable_hgrant1_out & ~n1894;
  assign n1896 = ~n1884 & ~n1895;
  assign n1897 = ~next_sys_fair<0>_out  & ~n1896;
  assign n1898 = ~n448 & ~n1897;
  assign n1899 = next_sys_fair<1>_out  & ~n1898;
  assign n1900 = ~next_sys_fair<1>_out  & ~n1896;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = reg_controllable_hmaster2_out & ~n1901;
  assign n1903 = ~reg_controllable_locked_out & ~n1889;
  assign n1904 = ~n509 & ~n1903;
  assign n1905 = ~reg_controllable_hgrant1_out & ~n1904;
  assign n1906 = ~n1884 & ~n1905;
  assign n1907 = ~next_sys_fair<0>_out  & ~n1906;
  assign n1908 = ~n508 & ~n1907;
  assign n1909 = next_sys_fair<1>_out  & ~n1908;
  assign n1910 = ~next_sys_fair<1>_out  & ~n1906;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~reg_controllable_hmaster2_out & ~n1911;
  assign n1913 = ~n1902 & ~n1912;
  assign n1914 = reg_controllable_hmaster1_out & ~n1913;
  assign n1915 = reg_i_hlock1_out & ~n1492;
  assign n1916 = ~reg_i_hlock1_out & ~n1518;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = reg_stateG10_1_out & ~n1917;
  assign n1919 = reg_i_hlock1_out & ~n1506;
  assign n1920 = ~reg_i_hlock1_out & ~n1525;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = ~reg_stateG10_1_out & ~n1921;
  assign n1923 = ~n1918 & ~n1922;
  assign n1924 = reg_controllable_hgrant1_out & ~n1923;
  assign n1925 = ~n1905 & ~n1924;
  assign n1926 = ~next_sys_fair<0>_out  & ~n1925;
  assign n1927 = ~n508 & ~n1926;
  assign n1928 = next_sys_fair<1>_out  & ~n1927;
  assign n1929 = ~next_sys_fair<1>_out  & ~n1925;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = ~reg_controllable_hmaster2_out & ~n1930;
  assign n1932 = ~n1902 & ~n1931;
  assign n1933 = ~reg_controllable_hmaster1_out & ~n1932;
  assign n1934 = ~n1914 & ~n1933;
  assign n1935 = reg_controllable_hmaster0_out & ~n1934;
  assign n1936 = ~reg_controllable_hmaster1_out & ~n1911;
  assign n1937 = ~n1914 & ~n1936;
  assign n1938 = ~reg_controllable_hmaster0_out & ~n1937;
  assign n1939 = ~n1935 & ~n1938;
  assign n1940 = next_sys_fair<2>_out  & ~n1939;
  assign n1941 = reg_stateG10_1_out & ~n1404;
  assign n1942 = reg_i_hlock1_out & ~n186;
  assign n1943 = ~reg_i_hlock1_out & ~n1404;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~reg_stateG10_1_out & ~n1944;
  assign n1946 = ~n1941 & ~n1945;
  assign n1947 = reg_controllable_hgrant1_out & ~n1946;
  assign n1948 = ~n1895 & ~n1947;
  assign n1949 = next_sys_fair<0>_out  & ~n1948;
  assign n1950 = ~n1897 & ~n1949;
  assign n1951 = next_sys_fair<1>_out  & ~n1950;
  assign n1952 = ~n572 & ~n1947;
  assign n1953 = next_sys_fair<0>_out  & ~n1952;
  assign n1954 = ~n598 & ~n1947;
  assign n1955 = ~next_sys_fair<0>_out  & ~n1954;
  assign n1956 = ~n1953 & ~n1955;
  assign n1957 = ~next_sys_fair<1>_out  & ~n1956;
  assign n1958 = ~n1951 & ~n1957;
  assign n1959 = reg_controllable_hmaster2_out & ~n1958;
  assign n1960 = ~n1905 & ~n1947;
  assign n1961 = next_sys_fair<0>_out  & ~n1960;
  assign n1962 = ~n1907 & ~n1961;
  assign n1963 = next_sys_fair<1>_out  & ~n1962;
  assign n1964 = ~n609 & ~n1947;
  assign n1965 = ~next_sys_fair<1>_out  & ~n1964;
  assign n1966 = ~n1963 & ~n1965;
  assign n1967 = ~reg_controllable_hmaster2_out & ~n1966;
  assign n1968 = ~n1959 & ~n1967;
  assign n1969 = reg_controllable_hmaster1_out & ~n1968;
  assign n1970 = reg_i_hlock1_out & ~n1446;
  assign n1971 = ~reg_i_hlock1_out & ~n1461;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = reg_stateG10_1_out & ~n1972;
  assign n1974 = reg_i_hlock1_out & ~n1450;
  assign n1975 = ~reg_i_hlock1_out & ~n1465;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~reg_stateG10_1_out & ~n1976;
  assign n1978 = ~n1973 & ~n1977;
  assign n1979 = reg_controllable_hgrant1_out & ~n1978;
  assign n1980 = ~n1905 & ~n1979;
  assign n1981 = next_sys_fair<0>_out  & ~n1980;
  assign n1982 = ~n1926 & ~n1981;
  assign n1983 = next_sys_fair<1>_out  & ~n1982;
  assign n1984 = reg_i_hlock1_out & ~n1555;
  assign n1985 = ~reg_i_hlock1_out & ~n1570;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = reg_stateG10_1_out & ~n1986;
  assign n1988 = reg_i_hlock1_out & ~n1559;
  assign n1989 = ~reg_i_hlock1_out & ~n1574;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = ~reg_stateG10_1_out & ~n1990;
  assign n1992 = ~n1987 & ~n1991;
  assign n1993 = reg_controllable_hgrant1_out & ~n1992;
  assign n1994 = ~n609 & ~n1993;
  assign n1995 = next_sys_fair<0>_out  & ~n1994;
  assign n1996 = reg_i_hlock1_out & ~n1589;
  assign n1997 = ~reg_i_hlock1_out & ~n1602;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = reg_stateG10_1_out & ~n1998;
  assign n2000 = reg_i_hlock1_out & ~n1593;
  assign n2001 = ~reg_i_hlock1_out & ~n1606;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~reg_stateG10_1_out & ~n2002;
  assign n2004 = ~n1999 & ~n2003;
  assign n2005 = reg_controllable_hgrant1_out & ~n2004;
  assign n2006 = ~n609 & ~n2005;
  assign n2007 = ~next_sys_fair<0>_out  & ~n2006;
  assign n2008 = ~n1995 & ~n2007;
  assign n2009 = ~next_sys_fair<1>_out  & ~n2008;
  assign n2010 = ~n1983 & ~n2009;
  assign n2011 = ~reg_controllable_hmaster2_out & ~n2010;
  assign n2012 = ~n1959 & ~n2011;
  assign n2013 = ~reg_controllable_hmaster1_out & ~n2012;
  assign n2014 = ~n1969 & ~n2013;
  assign n2015 = reg_controllable_hmaster0_out & ~n2014;
  assign n2016 = ~reg_controllable_hmaster1_out & ~n1966;
  assign n2017 = ~n1969 & ~n2016;
  assign n2018 = ~reg_controllable_hmaster0_out & ~n2017;
  assign n2019 = ~n2015 & ~n2018;
  assign n2020 = ~next_sys_fair<2>_out  & ~n2019;
  assign n2021 = ~n1940 & ~n2020;
  assign n2022 = ~reg_controllable_hgrant2_out & ~n2021;
  assign n2023 = ~n1877 & ~n2022;
  assign n2024 = ~reg_controllable_hgrant3_out & ~n2023;
  assign n2025 = ~n1786 & ~n2024;
  assign n2026 = ~reg_controllable_hgrant4_out & ~n2025;
  assign n2027 = ~n1630 & ~n2026;
  assign n2028 = reg_controllable_nhgrant0_out & ~n2027;
  assign n2029 = ~next_sys_fair<1>_out  & ~n1423;
  assign n2030 = ~n1678 & ~n2029;
  assign n2031 = reg_i_hlock0_out & ~n2030;
  assign n2032 = ~next_sys_fair<1>_out  & ~n1419;
  assign n2033 = ~n1633 & ~n2032;
  assign n2034 = ~reg_i_hlock0_out & ~n2033;
  assign n2035 = ~n2031 & ~n2034;
  assign n2036 = reg_controllable_hmaster0_out & ~n2035;
  assign n2037 = reg_controllable_hmaster1_out & ~n2035;
  assign n2038 = reg_controllable_hmaster2_out & ~n2035;
  assign n2039 = ~next_sys_fair<1>_out  & ~n1508;
  assign n2040 = ~n1685 & ~n2039;
  assign n2041 = reg_i_hlock0_out & ~n2040;
  assign n2042 = ~next_sys_fair<1>_out  & ~n1527;
  assign n2043 = ~n1754 & ~n2042;
  assign n2044 = ~reg_i_hlock0_out & ~n2043;
  assign n2045 = ~n2041 & ~n2044;
  assign n2046 = ~reg_controllable_hmaster2_out & ~n2045;
  assign n2047 = ~n2038 & ~n2046;
  assign n2048 = ~reg_controllable_hmaster1_out & ~n2047;
  assign n2049 = ~n2037 & ~n2048;
  assign n2050 = ~reg_controllable_hmaster0_out & ~n2049;
  assign n2051 = ~n2036 & ~n2050;
  assign n2052 = next_sys_fair<2>_out  & ~n2051;
  assign n2053 = next_sys_fair<1>_out  & ~n1808;
  assign n2054 = ~n394 & ~n2053;
  assign n2055 = reg_i_hlock0_out & ~n2054;
  assign n2056 = next_sys_fair<1>_out  & ~n1789;
  assign n2057 = ~n1656 & ~n2056;
  assign n2058 = ~reg_i_hlock0_out & ~n2057;
  assign n2059 = ~n2055 & ~n2058;
  assign n2060 = reg_controllable_hmaster0_out & ~n2059;
  assign n2061 = reg_controllable_hmaster1_out & ~n2059;
  assign n2062 = reg_controllable_hmaster2_out & ~n2059;
  assign n2063 = next_sys_fair<1>_out  & ~n1815;
  assign n2064 = ~n1706 & ~n2063;
  assign n2065 = reg_i_hlock0_out & ~n2064;
  assign n2066 = next_sys_fair<1>_out  & ~n1842;
  assign n2067 = ~n1770 & ~n2066;
  assign n2068 = ~reg_i_hlock0_out & ~n2067;
  assign n2069 = ~n2065 & ~n2068;
  assign n2070 = ~reg_controllable_hmaster2_out & ~n2069;
  assign n2071 = ~n2062 & ~n2070;
  assign n2072 = ~reg_controllable_hmaster1_out & ~n2071;
  assign n2073 = ~n2061 & ~n2072;
  assign n2074 = ~reg_controllable_hmaster0_out & ~n2073;
  assign n2075 = ~n2060 & ~n2074;
  assign n2076 = ~next_sys_fair<2>_out  & ~n2075;
  assign n2077 = ~n2052 & ~n2076;
  assign n2078 = ~reg_controllable_hgrant2_out & ~n2077;
  assign n2079 = ~reg_controllable_hgrant2_out & ~n2078;
  assign n2080 = ~reg_controllable_hgrant3_out & ~n2079;
  assign n2081 = ~reg_controllable_hgrant3_out & ~n2080;
  assign n2082 = ~reg_controllable_hgrant4_out & ~n2081;
  assign n2083 = ~reg_controllable_hgrant4_out & ~n2082;
  assign n2084 = ~reg_controllable_nhgrant0_out & ~n2083;
  assign n2085 = ~n2028 & ~n2084;
  assign n2086 = reg_i_hready_out & ~n2085;
  assign n2087 = next_sys_fair<0>_out  & ~n79;
  assign n2088 = ~next_sys_fair<0>_out  & ~n1885;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = next_sys_fair<1>_out  & ~n2089;
  assign n2091 = ~next_sys_fair<1>_out  & ~n1885;
  assign n2092 = ~n2090 & ~n2091;
  assign n2093 = reg_controllable_hmaster2_out & ~n2092;
  assign n2094 = ~n1485 & ~n1489;
  assign n2095 = ~next_sys_fair<0>_out  & ~n2094;
  assign n2096 = ~next_sys_fair<0>_out  & ~n2095;
  assign n2097 = next_sys_fair<1>_out  & ~n2096;
  assign n2098 = ~n1440 & ~n1443;
  assign n2099 = next_sys_fair<0>_out  & ~n2098;
  assign n2100 = ~n2095 & ~n2099;
  assign n2101 = ~next_sys_fair<1>_out  & ~n2100;
  assign n2102 = ~n2097 & ~n2101;
  assign n2103 = ~reg_controllable_hmaster2_out & ~n2102;
  assign n2104 = ~n2093 & ~n2103;
  assign n2105 = reg_controllable_hmaster1_out & ~n2104;
  assign n2106 = reg_i_hlock1_out & ~n2094;
  assign n2107 = ~n1512 & ~n1515;
  assign n2108 = ~reg_i_hlock1_out & ~n2107;
  assign n2109 = ~n2106 & ~n2108;
  assign n2110 = reg_stateG10_1_out & ~n2109;
  assign n2111 = ~n1489 & ~n1503;
  assign n2112 = reg_i_hlock1_out & ~n2111;
  assign n2113 = ~n1512 & ~n1522;
  assign n2114 = ~reg_i_hlock1_out & ~n2113;
  assign n2115 = ~n2112 & ~n2114;
  assign n2116 = ~reg_stateG10_1_out & ~n2115;
  assign n2117 = ~n2110 & ~n2116;
  assign n2118 = ~next_sys_fair<0>_out  & ~n2117;
  assign n2119 = ~next_sys_fair<0>_out  & ~n2118;
  assign n2120 = next_sys_fair<1>_out  & ~n2119;
  assign n2121 = ~next_sys_fair<1>_out  & ~n2117;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~reg_controllable_hmaster2_out & ~n2122;
  assign n2124 = ~n2093 & ~n2123;
  assign n2125 = ~reg_controllable_hmaster1_out & ~n2124;
  assign n2126 = ~n2105 & ~n2125;
  assign n2127 = reg_controllable_hmaster0_out & ~n2126;
  assign n2128 = next_sys_fair<0>_out  & ~n2094;
  assign n2129 = ~next_sys_fair<0>_out  & ~n2098;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~next_sys_fair<1>_out  & ~n2130;
  assign n2132 = ~n2097 & ~n2131;
  assign n2133 = ~reg_controllable_hmaster2_out & ~n2132;
  assign n2134 = ~n2093 & ~n2133;
  assign n2135 = reg_controllable_hmaster1_out & ~n2134;
  assign n2136 = reg_stateG10_4_out & ~n2098;
  assign n2137 = ~n228 & ~n1443;
  assign n2138 = ~reg_stateG10_4_out & ~n2137;
  assign n2139 = ~n2136 & ~n2138;
  assign n2140 = reg_i_hlock4_out & ~n2139;
  assign n2141 = ~n832 & ~n1458;
  assign n2142 = reg_stateG10_4_out & ~n2141;
  assign n2143 = ~reg_stateG10_4_out & ~n833;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~reg_i_hlock4_out & ~n2144;
  assign n2146 = ~n2140 & ~n2145;
  assign n2147 = ~next_sys_fair<0>_out  & ~n2146;
  assign n2148 = ~next_sys_fair<0>_out  & ~n2147;
  assign n2149 = next_sys_fair<1>_out  & ~n2148;
  assign n2150 = reg_stateG10_4_out & ~n2094;
  assign n2151 = ~reg_stateG10_4_out & ~n2111;
  assign n2152 = ~n2150 & ~n2151;
  assign n2153 = reg_i_hlock4_out & ~n2152;
  assign n2154 = reg_stateG10_4_out & ~n2107;
  assign n2155 = ~reg_stateG10_4_out & ~n2113;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~reg_i_hlock4_out & ~n2156;
  assign n2158 = ~n2153 & ~n2157;
  assign n2159 = ~next_sys_fair<1>_out  & ~n2158;
  assign n2160 = ~n2149 & ~n2159;
  assign n2161 = reg_controllable_hmaster2_out & ~n2160;
  assign n2162 = ~next_sys_fair<0>_out  & ~n2111;
  assign n2163 = ~next_sys_fair<0>_out  & ~n2162;
  assign n2164 = next_sys_fair<1>_out  & ~n2163;
  assign n2165 = ~next_sys_fair<1>_out  & ~n2111;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = reg_i_hlock0_out & ~n2166;
  assign n2168 = ~next_sys_fair<0>_out  & ~n2113;
  assign n2169 = ~next_sys_fair<0>_out  & ~n2168;
  assign n2170 = next_sys_fair<1>_out  & ~n2169;
  assign n2171 = ~next_sys_fair<1>_out  & ~n2113;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~reg_i_hlock0_out & ~n2172;
  assign n2174 = ~n2167 & ~n2173;
  assign n2175 = ~reg_controllable_hmaster2_out & ~n2174;
  assign n2176 = ~n2161 & ~n2175;
  assign n2177 = ~reg_controllable_hmaster1_out & ~n2176;
  assign n2178 = ~n2135 & ~n2177;
  assign n2179 = ~reg_controllable_hmaster0_out & ~n2178;
  assign n2180 = ~n2127 & ~n2179;
  assign n2181 = reg_stateG10_2_out & ~n2180;
  assign n2182 = next_sys_fair<0>_out  & ~n2111;
  assign n2183 = ~next_sys_fair<0>_out  & ~n2137;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~next_sys_fair<1>_out  & ~n2184;
  assign n2186 = ~n2164 & ~n2185;
  assign n2187 = ~reg_controllable_hmaster2_out & ~n2186;
  assign n2188 = ~n2093 & ~n2187;
  assign n2189 = reg_controllable_hmaster1_out & ~n2188;
  assign n2190 = ~n2177 & ~n2189;
  assign n2191 = ~reg_controllable_hmaster0_out & ~n2190;
  assign n2192 = ~n2127 & ~n2191;
  assign n2193 = ~reg_stateG10_2_out & ~n2192;
  assign n2194 = ~n2181 & ~n2193;
  assign n2195 = reg_i_hlock2_out & ~n2194;
  assign n2196 = ~next_sys_fair<0>_out  & ~n2107;
  assign n2197 = ~next_sys_fair<0>_out  & ~n2196;
  assign n2198 = next_sys_fair<1>_out  & ~n2197;
  assign n2199 = next_sys_fair<0>_out  & ~n2107;
  assign n2200 = ~next_sys_fair<0>_out  & ~n2141;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~next_sys_fair<1>_out  & ~n2201;
  assign n2203 = ~n2198 & ~n2202;
  assign n2204 = ~reg_controllable_hmaster2_out & ~n2203;
  assign n2205 = ~n2093 & ~n2204;
  assign n2206 = reg_controllable_hmaster1_out & ~n2205;
  assign n2207 = ~n2177 & ~n2206;
  assign n2208 = ~reg_controllable_hmaster0_out & ~n2207;
  assign n2209 = ~n2127 & ~n2208;
  assign n2210 = reg_stateG10_2_out & ~n2209;
  assign n2211 = next_sys_fair<0>_out  & ~n2113;
  assign n2212 = ~next_sys_fair<0>_out  & ~n833;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = ~next_sys_fair<1>_out  & ~n2213;
  assign n2215 = ~n2170 & ~n2214;
  assign n2216 = ~reg_controllable_hmaster2_out & ~n2215;
  assign n2217 = ~n2093 & ~n2216;
  assign n2218 = reg_controllable_hmaster1_out & ~n2217;
  assign n2219 = ~n2177 & ~n2218;
  assign n2220 = ~reg_controllable_hmaster0_out & ~n2219;
  assign n2221 = ~n2127 & ~n2220;
  assign n2222 = ~reg_stateG10_2_out & ~n2221;
  assign n2223 = ~n2210 & ~n2222;
  assign n2224 = ~reg_i_hlock2_out & ~n2223;
  assign n2225 = ~n2195 & ~n2224;
  assign n2226 = next_sys_fair<2>_out  & ~n2225;
  assign n2227 = next_sys_fair<1>_out  & ~n1885;
  assign n2228 = next_sys_fair<0>_out  & ~n563;
  assign n2229 = ~next_sys_fair<0>_out  & ~n590;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = ~next_sys_fair<1>_out  & ~n2230;
  assign n2232 = ~n2227 & ~n2231;
  assign n2233 = reg_controllable_hmaster2_out & ~n2232;
  assign n2234 = next_sys_fair<1>_out  & ~n2094;
  assign n2235 = ~n1549 & ~n1552;
  assign n2236 = next_sys_fair<0>_out  & ~n2235;
  assign n2237 = ~n1443 & ~n1586;
  assign n2238 = ~next_sys_fair<0>_out  & ~n2237;
  assign n2239 = ~n2236 & ~n2238;
  assign n2240 = ~next_sys_fair<1>_out  & ~n2239;
  assign n2241 = ~n2234 & ~n2240;
  assign n2242 = ~reg_controllable_hmaster2_out & ~n2241;
  assign n2243 = ~n2233 & ~n2242;
  assign n2244 = reg_controllable_hmaster1_out & ~n2243;
  assign n2245 = reg_i_hlock1_out & ~n2098;
  assign n2246 = ~reg_i_hlock1_out & ~n2141;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = reg_stateG10_1_out & ~n2247;
  assign n2249 = reg_i_hlock1_out & ~n2137;
  assign n2250 = ~reg_i_hlock1_out & ~n833;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = ~reg_stateG10_1_out & ~n2251;
  assign n2253 = ~n2248 & ~n2252;
  assign n2254 = next_sys_fair<0>_out  & ~n2253;
  assign n2255 = ~n2118 & ~n2254;
  assign n2256 = next_sys_fair<1>_out  & ~n2255;
  assign n2257 = reg_i_hlock1_out & ~n2235;
  assign n2258 = ~n945 & ~n1567;
  assign n2259 = ~reg_i_hlock1_out & ~n2258;
  assign n2260 = ~n2257 & ~n2259;
  assign n2261 = reg_stateG10_1_out & ~n2260;
  assign n2262 = ~n319 & ~n1552;
  assign n2263 = reg_i_hlock1_out & ~n2262;
  assign n2264 = ~reg_i_hlock1_out & ~n946;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = ~reg_stateG10_1_out & ~n2265;
  assign n2267 = ~n2261 & ~n2266;
  assign n2268 = next_sys_fair<0>_out  & ~n2267;
  assign n2269 = reg_i_hlock1_out & ~n2237;
  assign n2270 = ~n832 & ~n1599;
  assign n2271 = ~reg_i_hlock1_out & ~n2270;
  assign n2272 = ~n2269 & ~n2271;
  assign n2273 = reg_stateG10_1_out & ~n2272;
  assign n2274 = ~n340 & ~n1443;
  assign n2275 = reg_i_hlock1_out & ~n2274;
  assign n2276 = ~reg_i_hlock1_out & ~n956;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~reg_stateG10_1_out & ~n2277;
  assign n2279 = ~n2273 & ~n2278;
  assign n2280 = ~next_sys_fair<0>_out  & ~n2279;
  assign n2281 = ~n2268 & ~n2280;
  assign n2282 = ~next_sys_fair<1>_out  & ~n2281;
  assign n2283 = ~n2256 & ~n2282;
  assign n2284 = ~reg_controllable_hmaster2_out & ~n2283;
  assign n2285 = ~n2233 & ~n2284;
  assign n2286 = ~reg_controllable_hmaster1_out & ~n2285;
  assign n2287 = ~n2244 & ~n2286;
  assign n2288 = reg_controllable_hmaster0_out & ~n2287;
  assign n2289 = next_sys_fair<1>_out  & ~n2158;
  assign n2290 = reg_stateG10_4_out & ~n2235;
  assign n2291 = ~reg_stateG10_4_out & ~n2262;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = reg_i_hlock4_out & ~n2292;
  assign n2294 = reg_stateG10_4_out & ~n2258;
  assign n2295 = ~reg_stateG10_4_out & ~n946;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = ~reg_i_hlock4_out & ~n2296;
  assign n2298 = ~n2293 & ~n2297;
  assign n2299 = next_sys_fair<0>_out  & ~n2298;
  assign n2300 = reg_stateG10_4_out & ~n2237;
  assign n2301 = ~reg_stateG10_4_out & ~n2274;
  assign n2302 = ~n2300 & ~n2301;
  assign n2303 = reg_i_hlock4_out & ~n2302;
  assign n2304 = reg_stateG10_4_out & ~n2270;
  assign n2305 = ~reg_stateG10_4_out & ~n956;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = ~reg_i_hlock4_out & ~n2306;
  assign n2308 = ~n2303 & ~n2307;
  assign n2309 = ~next_sys_fair<0>_out  & ~n2308;
  assign n2310 = ~n2299 & ~n2309;
  assign n2311 = ~next_sys_fair<1>_out  & ~n2310;
  assign n2312 = ~n2289 & ~n2311;
  assign n2313 = reg_controllable_hmaster2_out & ~n2312;
  assign n2314 = next_sys_fair<1>_out  & ~n2184;
  assign n2315 = next_sys_fair<0>_out  & ~n2262;
  assign n2316 = ~next_sys_fair<0>_out  & ~n2274;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~next_sys_fair<1>_out  & ~n2317;
  assign n2319 = ~n2314 & ~n2318;
  assign n2320 = reg_i_hlock0_out & ~n2319;
  assign n2321 = next_sys_fair<1>_out  & ~n2213;
  assign n2322 = next_sys_fair<0>_out  & ~n946;
  assign n2323 = ~next_sys_fair<0>_out  & ~n956;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~next_sys_fair<1>_out  & ~n2324;
  assign n2326 = ~n2321 & ~n2325;
  assign n2327 = ~reg_i_hlock0_out & ~n2326;
  assign n2328 = ~n2320 & ~n2327;
  assign n2329 = ~reg_controllable_hmaster2_out & ~n2328;
  assign n2330 = ~n2313 & ~n2329;
  assign n2331 = ~reg_controllable_hmaster1_out & ~n2330;
  assign n2332 = ~n2244 & ~n2331;
  assign n2333 = ~reg_controllable_hmaster0_out & ~n2332;
  assign n2334 = ~n2288 & ~n2333;
  assign n2335 = reg_stateG10_2_out & ~n2334;
  assign n2336 = next_sys_fair<1>_out  & ~n2111;
  assign n2337 = ~n2318 & ~n2336;
  assign n2338 = ~reg_controllable_hmaster2_out & ~n2337;
  assign n2339 = ~n2233 & ~n2338;
  assign n2340 = reg_controllable_hmaster1_out & ~n2339;
  assign n2341 = ~n2331 & ~n2340;
  assign n2342 = ~reg_controllable_hmaster0_out & ~n2341;
  assign n2343 = ~n2288 & ~n2342;
  assign n2344 = ~reg_stateG10_2_out & ~n2343;
  assign n2345 = ~n2335 & ~n2344;
  assign n2346 = reg_i_hlock2_out & ~n2345;
  assign n2347 = next_sys_fair<1>_out  & ~n2107;
  assign n2348 = next_sys_fair<0>_out  & ~n2258;
  assign n2349 = ~next_sys_fair<0>_out  & ~n2270;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~next_sys_fair<1>_out  & ~n2350;
  assign n2352 = ~n2347 & ~n2351;
  assign n2353 = ~reg_controllable_hmaster2_out & ~n2352;
  assign n2354 = ~n2233 & ~n2353;
  assign n2355 = reg_controllable_hmaster1_out & ~n2354;
  assign n2356 = ~n2331 & ~n2355;
  assign n2357 = ~reg_controllable_hmaster0_out & ~n2356;
  assign n2358 = ~n2288 & ~n2357;
  assign n2359 = reg_stateG10_2_out & ~n2358;
  assign n2360 = next_sys_fair<1>_out  & ~n2113;
  assign n2361 = ~n2325 & ~n2360;
  assign n2362 = ~reg_controllable_hmaster2_out & ~n2361;
  assign n2363 = ~n2233 & ~n2362;
  assign n2364 = reg_controllable_hmaster1_out & ~n2363;
  assign n2365 = ~n2331 & ~n2364;
  assign n2366 = ~reg_controllable_hmaster0_out & ~n2365;
  assign n2367 = ~n2288 & ~n2366;
  assign n2368 = ~reg_stateG10_2_out & ~n2367;
  assign n2369 = ~n2359 & ~n2368;
  assign n2370 = ~reg_i_hlock2_out & ~n2369;
  assign n2371 = ~n2346 & ~n2370;
  assign n2372 = ~next_sys_fair<2>_out  & ~n2371;
  assign n2373 = ~n2226 & ~n2372;
  assign n2374 = reg_stateG10_3_out & ~n2373;
  assign n2375 = next_sys_fair<0>_out  & ~n2137;
  assign n2376 = ~n2162 & ~n2375;
  assign n2377 = ~next_sys_fair<1>_out  & ~n2376;
  assign n2378 = ~n2164 & ~n2377;
  assign n2379 = ~reg_controllable_hmaster2_out & ~n2378;
  assign n2380 = ~n2093 & ~n2379;
  assign n2381 = reg_controllable_hmaster1_out & ~n2380;
  assign n2382 = ~n2125 & ~n2381;
  assign n2383 = reg_controllable_hmaster0_out & ~n2382;
  assign n2384 = ~n2179 & ~n2383;
  assign n2385 = reg_stateG10_2_out & ~n2384;
  assign n2386 = ~n2191 & ~n2383;
  assign n2387 = ~reg_stateG10_2_out & ~n2386;
  assign n2388 = ~n2385 & ~n2387;
  assign n2389 = reg_i_hlock2_out & ~n2388;
  assign n2390 = ~n2208 & ~n2383;
  assign n2391 = reg_stateG10_2_out & ~n2390;
  assign n2392 = ~n2220 & ~n2383;
  assign n2393 = ~reg_stateG10_2_out & ~n2392;
  assign n2394 = ~n2391 & ~n2393;
  assign n2395 = ~reg_i_hlock2_out & ~n2394;
  assign n2396 = ~n2389 & ~n2395;
  assign n2397 = next_sys_fair<2>_out  & ~n2396;
  assign n2398 = ~n2286 & ~n2340;
  assign n2399 = reg_controllable_hmaster0_out & ~n2398;
  assign n2400 = ~n2333 & ~n2399;
  assign n2401 = reg_stateG10_2_out & ~n2400;
  assign n2402 = ~n2342 & ~n2399;
  assign n2403 = ~reg_stateG10_2_out & ~n2402;
  assign n2404 = ~n2401 & ~n2403;
  assign n2405 = reg_i_hlock2_out & ~n2404;
  assign n2406 = ~n2357 & ~n2399;
  assign n2407 = reg_stateG10_2_out & ~n2406;
  assign n2408 = ~n2366 & ~n2399;
  assign n2409 = ~reg_stateG10_2_out & ~n2408;
  assign n2410 = ~n2407 & ~n2409;
  assign n2411 = ~reg_i_hlock2_out & ~n2410;
  assign n2412 = ~n2405 & ~n2411;
  assign n2413 = ~next_sys_fair<2>_out  & ~n2412;
  assign n2414 = ~n2397 & ~n2413;
  assign n2415 = ~reg_stateG10_3_out & ~n2414;
  assign n2416 = ~n2374 & ~n2415;
  assign n2417 = reg_i_hlock3_out & ~n2416;
  assign n2418 = next_sys_fair<0>_out  & ~n2141;
  assign n2419 = ~n2196 & ~n2418;
  assign n2420 = ~next_sys_fair<1>_out  & ~n2419;
  assign n2421 = ~n2198 & ~n2420;
  assign n2422 = ~reg_controllable_hmaster2_out & ~n2421;
  assign n2423 = ~n2093 & ~n2422;
  assign n2424 = reg_controllable_hmaster1_out & ~n2423;
  assign n2425 = ~n2125 & ~n2424;
  assign n2426 = reg_controllable_hmaster0_out & ~n2425;
  assign n2427 = ~n2179 & ~n2426;
  assign n2428 = reg_stateG10_2_out & ~n2427;
  assign n2429 = ~n2191 & ~n2426;
  assign n2430 = ~reg_stateG10_2_out & ~n2429;
  assign n2431 = ~n2428 & ~n2430;
  assign n2432 = reg_i_hlock2_out & ~n2431;
  assign n2433 = ~n2208 & ~n2426;
  assign n2434 = reg_stateG10_2_out & ~n2433;
  assign n2435 = ~n2220 & ~n2426;
  assign n2436 = ~reg_stateG10_2_out & ~n2435;
  assign n2437 = ~n2434 & ~n2436;
  assign n2438 = ~reg_i_hlock2_out & ~n2437;
  assign n2439 = ~n2432 & ~n2438;
  assign n2440 = next_sys_fair<2>_out  & ~n2439;
  assign n2441 = ~n2286 & ~n2355;
  assign n2442 = reg_controllable_hmaster0_out & ~n2441;
  assign n2443 = ~n2333 & ~n2442;
  assign n2444 = reg_stateG10_2_out & ~n2443;
  assign n2445 = ~n2342 & ~n2442;
  assign n2446 = ~reg_stateG10_2_out & ~n2445;
  assign n2447 = ~n2444 & ~n2446;
  assign n2448 = reg_i_hlock2_out & ~n2447;
  assign n2449 = ~n2357 & ~n2442;
  assign n2450 = reg_stateG10_2_out & ~n2449;
  assign n2451 = ~n2366 & ~n2442;
  assign n2452 = ~reg_stateG10_2_out & ~n2451;
  assign n2453 = ~n2450 & ~n2452;
  assign n2454 = ~reg_i_hlock2_out & ~n2453;
  assign n2455 = ~n2448 & ~n2454;
  assign n2456 = ~next_sys_fair<2>_out  & ~n2455;
  assign n2457 = ~n2440 & ~n2456;
  assign n2458 = reg_stateG10_3_out & ~n2457;
  assign n2459 = next_sys_fair<0>_out  & ~n833;
  assign n2460 = ~n2168 & ~n2459;
  assign n2461 = ~next_sys_fair<1>_out  & ~n2460;
  assign n2462 = ~n2170 & ~n2461;
  assign n2463 = ~reg_controllable_hmaster2_out & ~n2462;
  assign n2464 = ~n2093 & ~n2463;
  assign n2465 = reg_controllable_hmaster1_out & ~n2464;
  assign n2466 = ~n2125 & ~n2465;
  assign n2467 = reg_controllable_hmaster0_out & ~n2466;
  assign n2468 = ~n2179 & ~n2467;
  assign n2469 = reg_stateG10_2_out & ~n2468;
  assign n2470 = ~n2191 & ~n2467;
  assign n2471 = ~reg_stateG10_2_out & ~n2470;
  assign n2472 = ~n2469 & ~n2471;
  assign n2473 = reg_i_hlock2_out & ~n2472;
  assign n2474 = ~n2208 & ~n2467;
  assign n2475 = reg_stateG10_2_out & ~n2474;
  assign n2476 = ~n2220 & ~n2467;
  assign n2477 = ~reg_stateG10_2_out & ~n2476;
  assign n2478 = ~n2475 & ~n2477;
  assign n2479 = ~reg_i_hlock2_out & ~n2478;
  assign n2480 = ~n2473 & ~n2479;
  assign n2481 = next_sys_fair<2>_out  & ~n2480;
  assign n2482 = ~n2286 & ~n2364;
  assign n2483 = reg_controllable_hmaster0_out & ~n2482;
  assign n2484 = ~n2333 & ~n2483;
  assign n2485 = reg_stateG10_2_out & ~n2484;
  assign n2486 = ~n2342 & ~n2483;
  assign n2487 = ~reg_stateG10_2_out & ~n2486;
  assign n2488 = ~n2485 & ~n2487;
  assign n2489 = reg_i_hlock2_out & ~n2488;
  assign n2490 = ~n2357 & ~n2483;
  assign n2491 = reg_stateG10_2_out & ~n2490;
  assign n2492 = ~n2366 & ~n2483;
  assign n2493 = ~reg_stateG10_2_out & ~n2492;
  assign n2494 = ~n2491 & ~n2493;
  assign n2495 = ~reg_i_hlock2_out & ~n2494;
  assign n2496 = ~n2489 & ~n2495;
  assign n2497 = ~next_sys_fair<2>_out  & ~n2496;
  assign n2498 = ~n2481 & ~n2497;
  assign n2499 = ~reg_stateG10_3_out & ~n2498;
  assign n2500 = ~n2458 & ~n2499;
  assign n2501 = ~reg_i_hlock3_out & ~n2500;
  assign n2502 = ~n2417 & ~n2501;
  assign n2503 = ~reg_i_hready_out & ~n2502;
  assign n2504 = ~n2086 & ~n2503;
  assign n2505 = ~next_sys_fair<3>_out  & ~n2504;
  assign n2506 = ~n1403 & ~n2505;
  assign n2507 = reg_i_hbusreq0_out & ~n2506;
  assign n2508 = reg_i_hbusreq4_out & ~n2506;
  assign n2509 = reg_i_hbusreq1_out & ~n2506;
  assign n2510 = reg_i_hbusreq2_out & ~n2506;
  assign n2511 = reg_i_hbusreq3_out & ~n2506;
  assign n2512 = ~reg_controllable_locked_out & ~n176;
  assign n2513 = ~reg_controllable_locked_out & ~n2512;
  assign n2514 = ~reg_controllable_hgrant1_out & ~n2513;
  assign n2515 = ~reg_controllable_hgrant1_out & ~n2514;
  assign n2516 = ~next_sys_fair<0>_out  & ~n2515;
  assign n2517 = ~next_sys_fair<0>_out  & ~n2516;
  assign n2518 = next_sys_fair<1>_out  & ~n2517;
  assign n2519 = ~next_env_fair_out & ~n173;
  assign n2520 = ~next_env_fair_out & ~n2519;
  assign n2521 = ~fair_cnt<2>_out  & ~n2520;
  assign n2522 = ~fair_cnt<2>_out  & ~n2521;
  assign n2523 = ~reg_controllable_locked_out & ~n2522;
  assign n2524 = ~reg_controllable_locked_out & ~n2523;
  assign n2525 = ~reg_controllable_hgrant1_out & ~n2524;
  assign n2526 = ~reg_controllable_hgrant1_out & ~n2525;
  assign n2527 = ~next_sys_fair<1>_out  & ~n2526;
  assign n2528 = ~n2518 & ~n2527;
  assign n2529 = reg_i_hlock0_out & ~n2528;
  assign n2530 = ~next_sys_fair<0>_out  & ~n1788;
  assign n2531 = next_sys_fair<1>_out  & ~n2530;
  assign n2532 = ~reg_controllable_locked_out & ~n205;
  assign n2533 = ~reg_controllable_hgrant1_out & ~n2532;
  assign n2534 = ~reg_controllable_hgrant1_out & ~n2533;
  assign n2535 = ~next_sys_fair<1>_out  & ~n2534;
  assign n2536 = ~n2531 & ~n2535;
  assign n2537 = ~reg_i_hlock0_out & ~n2536;
  assign n2538 = ~n2529 & ~n2537;
  assign n2539 = reg_controllable_hmaster0_out & ~n2538;
  assign n2540 = reg_controllable_hmaster1_out & ~n2538;
  assign n2541 = reg_controllable_hmastlock_out & ~n176;
  assign n2542 = ~n771 & ~n2541;
  assign n2543 = ~reg_controllable_locked_out & ~n2542;
  assign n2544 = ~reg_controllable_locked_out & ~n2543;
  assign n2545 = ~reg_controllable_hgrant1_out & ~n2544;
  assign n2546 = ~reg_controllable_hgrant1_out & ~n2545;
  assign n2547 = ~next_sys_fair<0>_out  & ~n2546;
  assign n2548 = ~next_sys_fair<0>_out  & ~n2547;
  assign n2549 = next_sys_fair<1>_out  & ~n2548;
  assign n2550 = reg_controllable_hmastlock_out & ~n2522;
  assign n2551 = ~n791 & ~n2550;
  assign n2552 = ~reg_controllable_locked_out & ~n2551;
  assign n2553 = ~reg_controllable_locked_out & ~n2552;
  assign n2554 = ~reg_controllable_hgrant1_out & ~n2553;
  assign n2555 = ~reg_controllable_hgrant1_out & ~n2554;
  assign n2556 = ~next_sys_fair<1>_out  & ~n2555;
  assign n2557 = ~n2549 & ~n2556;
  assign n2558 = reg_i_hlock0_out & ~n2557;
  assign n2559 = ~n1445 & ~n1457;
  assign n2560 = ~reg_controllable_hgrant1_out & ~n2559;
  assign n2561 = ~reg_controllable_hgrant1_out & ~n2560;
  assign n2562 = ~next_sys_fair<0>_out  & ~n2561;
  assign n2563 = ~next_sys_fair<0>_out  & ~n2562;
  assign n2564 = next_sys_fair<1>_out  & ~n2563;
  assign n2565 = reg_controllable_hmastlock_out & ~n845;
  assign n2566 = reg_controllable_locked_out & ~n2565;
  assign n2567 = ~reg_controllable_hmastlock_out & ~n801;
  assign n2568 = ~n285 & ~n2567;
  assign n2569 = ~reg_controllable_locked_out & ~n2568;
  assign n2570 = ~n2566 & ~n2569;
  assign n2571 = ~reg_controllable_hgrant1_out & ~n2570;
  assign n2572 = ~reg_controllable_hgrant1_out & ~n2571;
  assign n2573 = ~next_sys_fair<1>_out  & ~n2572;
  assign n2574 = ~n2564 & ~n2573;
  assign n2575 = ~reg_i_hlock0_out & ~n2574;
  assign n2576 = ~n2558 & ~n2575;
  assign n2577 = reg_controllable_hmaster2_out & ~n2576;
  assign n2578 = ~reg_controllable_hmaster2_out & ~n2538;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = ~reg_controllable_hmaster1_out & ~n2579;
  assign n2581 = ~n2540 & ~n2580;
  assign n2582 = ~reg_controllable_hmaster0_out & ~n2581;
  assign n2583 = ~n2539 & ~n2582;
  assign n2584 = next_sys_fair<2>_out  & ~n2583;
  assign n2585 = next_sys_fair<0>_out  & ~n2526;
  assign n2586 = ~fair_cnt<2>_out  & ~n175;
  assign n2587 = ~reg_controllable_locked_out & ~n2586;
  assign n2588 = ~reg_controllable_locked_out & ~n2587;
  assign n2589 = ~reg_controllable_hgrant1_out & ~n2588;
  assign n2590 = ~reg_controllable_hgrant1_out & ~n2589;
  assign n2591 = ~next_sys_fair<0>_out  & ~n2590;
  assign n2592 = ~n2585 & ~n2591;
  assign n2593 = next_sys_fair<1>_out  & ~n2592;
  assign n2594 = ~next_sys_fair<1>_out  & ~n2515;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = reg_i_hlock0_out & ~n2595;
  assign n2597 = next_sys_fair<0>_out  & ~n2534;
  assign n2598 = ~n1631 & ~n2597;
  assign n2599 = next_sys_fair<1>_out  & ~n2598;
  assign n2600 = ~n1656 & ~n2599;
  assign n2601 = ~reg_i_hlock0_out & ~n2600;
  assign n2602 = ~n2596 & ~n2601;
  assign n2603 = reg_controllable_hmaster0_out & ~n2602;
  assign n2604 = reg_controllable_hmaster1_out & ~n2602;
  assign n2605 = next_sys_fair<0>_out  & ~n2555;
  assign n2606 = reg_controllable_hmastlock_out & ~n2586;
  assign n2607 = ~n751 & ~n2606;
  assign n2608 = ~reg_controllable_locked_out & ~n2607;
  assign n2609 = ~reg_controllable_locked_out & ~n2608;
  assign n2610 = ~reg_controllable_hgrant1_out & ~n2609;
  assign n2611 = ~reg_controllable_hgrant1_out & ~n2610;
  assign n2612 = ~next_sys_fair<0>_out  & ~n2611;
  assign n2613 = ~n2605 & ~n2612;
  assign n2614 = next_sys_fair<1>_out  & ~n2613;
  assign n2615 = ~n918 & ~n2541;
  assign n2616 = ~reg_controllable_locked_out & ~n2615;
  assign n2617 = ~reg_controllable_locked_out & ~n2616;
  assign n2618 = ~reg_controllable_hgrant1_out & ~n2617;
  assign n2619 = ~reg_controllable_hgrant1_out & ~n2618;
  assign n2620 = next_sys_fair<0>_out  & ~n2619;
  assign n2621 = ~n2547 & ~n2620;
  assign n2622 = ~next_sys_fair<1>_out  & ~n2621;
  assign n2623 = ~n2614 & ~n2622;
  assign n2624 = reg_i_hlock0_out & ~n2623;
  assign n2625 = next_sys_fair<0>_out  & ~n2572;
  assign n2626 = ~n1491 & ~n1514;
  assign n2627 = ~reg_controllable_hgrant1_out & ~n2626;
  assign n2628 = ~reg_controllable_hgrant1_out & ~n2627;
  assign n2629 = ~next_sys_fair<0>_out  & ~n2628;
  assign n2630 = ~n2625 & ~n2629;
  assign n2631 = next_sys_fair<1>_out  & ~n2630;
  assign n2632 = ~n1554 & ~n1566;
  assign n2633 = ~reg_controllable_hgrant1_out & ~n2632;
  assign n2634 = ~reg_controllable_hgrant1_out & ~n2633;
  assign n2635 = next_sys_fair<0>_out  & ~n2634;
  assign n2636 = ~n2562 & ~n2635;
  assign n2637 = ~next_sys_fair<1>_out  & ~n2636;
  assign n2638 = ~n2631 & ~n2637;
  assign n2639 = ~reg_i_hlock0_out & ~n2638;
  assign n2640 = ~n2624 & ~n2639;
  assign n2641 = reg_controllable_hmaster2_out & ~n2640;
  assign n2642 = ~reg_controllable_hmaster2_out & ~n2602;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = ~reg_controllable_hmaster1_out & ~n2643;
  assign n2645 = ~n2604 & ~n2644;
  assign n2646 = ~reg_controllable_hmaster0_out & ~n2645;
  assign n2647 = ~n2603 & ~n2646;
  assign n2648 = ~next_sys_fair<2>_out  & ~n2647;
  assign n2649 = ~n2584 & ~n2648;
  assign n2650 = ~reg_controllable_hgrant2_out & ~n2649;
  assign n2651 = ~reg_controllable_hgrant2_out & ~n2650;
  assign n2652 = ~reg_controllable_hgrant3_out & ~n2651;
  assign n2653 = ~reg_controllable_hgrant3_out & ~n2652;
  assign n2654 = reg_controllable_hgrant4_out & ~n2653;
  assign n2655 = ~next_sys_fair<0>_out  & ~n2526;
  assign n2656 = ~next_sys_fair<0>_out  & ~n2655;
  assign n2657 = next_sys_fair<1>_out  & ~n2656;
  assign n2658 = next_sys_fair<0>_out  & ~n2515;
  assign n2659 = ~n2655 & ~n2658;
  assign n2660 = ~next_sys_fair<1>_out  & ~n2659;
  assign n2661 = ~n2657 & ~n2660;
  assign n2662 = reg_i_hlock0_out & ~n2661;
  assign n2663 = ~next_sys_fair<0>_out  & ~n2534;
  assign n2664 = ~next_sys_fair<0>_out  & ~n2663;
  assign n2665 = next_sys_fair<1>_out  & ~n2664;
  assign n2666 = ~n1634 & ~n2663;
  assign n2667 = ~next_sys_fair<1>_out  & ~n2666;
  assign n2668 = ~n2665 & ~n2667;
  assign n2669 = ~reg_i_hlock0_out & ~n2668;
  assign n2670 = ~n2662 & ~n2669;
  assign n2671 = reg_controllable_hmaster2_out & ~n2670;
  assign n2672 = ~next_sys_fair<0>_out  & ~n2555;
  assign n2673 = ~next_sys_fair<0>_out  & ~n2672;
  assign n2674 = next_sys_fair<1>_out  & ~n2673;
  assign n2675 = next_sys_fair<0>_out  & ~n2546;
  assign n2676 = ~n2672 & ~n2675;
  assign n2677 = ~next_sys_fair<1>_out  & ~n2676;
  assign n2678 = ~n2674 & ~n2677;
  assign n2679 = reg_i_hlock0_out & ~n2678;
  assign n2680 = ~next_sys_fair<0>_out  & ~n2572;
  assign n2681 = ~next_sys_fair<0>_out  & ~n2680;
  assign n2682 = next_sys_fair<1>_out  & ~n2681;
  assign n2683 = next_sys_fair<0>_out  & ~n2561;
  assign n2684 = ~n2680 & ~n2683;
  assign n2685 = ~next_sys_fair<1>_out  & ~n2684;
  assign n2686 = ~n2682 & ~n2685;
  assign n2687 = ~reg_i_hlock0_out & ~n2686;
  assign n2688 = ~n2679 & ~n2687;
  assign n2689 = ~reg_controllable_hmaster2_out & ~n2688;
  assign n2690 = ~n2671 & ~n2689;
  assign n2691 = reg_controllable_hmaster1_out & ~n2690;
  assign n2692 = ~reg_controllable_hmaster1_out & ~n2670;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = reg_controllable_hmaster0_out & ~n2693;
  assign n2695 = ~reg_controllable_hmaster0_out & ~n2670;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = next_sys_fair<2>_out  & ~n2696;
  assign n2698 = reg_controllable_hmaster2_out & ~n2602;
  assign n2699 = ~reg_controllable_hmaster2_out & ~n2640;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = reg_controllable_hmaster1_out & ~n2700;
  assign n2702 = ~reg_controllable_hmaster1_out & ~n2602;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = reg_controllable_hmaster0_out & ~n2703;
  assign n2705 = ~reg_controllable_hmaster0_out & ~n2602;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~next_sys_fair<2>_out  & ~n2706;
  assign n2708 = ~n2697 & ~n2707;
  assign n2709 = ~reg_controllable_hgrant2_out & ~n2708;
  assign n2710 = ~reg_controllable_hgrant2_out & ~n2709;
  assign n2711 = reg_controllable_hgrant3_out & ~n2710;
  assign n2712 = ~n2516 & ~n2585;
  assign n2713 = ~next_sys_fair<1>_out  & ~n2712;
  assign n2714 = ~n2657 & ~n2713;
  assign n2715 = reg_i_hlock0_out & ~n2714;
  assign n2716 = ~n1788 & ~n2597;
  assign n2717 = ~next_sys_fair<1>_out  & ~n2716;
  assign n2718 = ~n2665 & ~n2717;
  assign n2719 = ~reg_i_hlock0_out & ~n2718;
  assign n2720 = ~n2715 & ~n2719;
  assign n2721 = reg_controllable_hmaster0_out & ~n2720;
  assign n2722 = reg_controllable_hmaster2_out & ~n2720;
  assign n2723 = ~n2547 & ~n2605;
  assign n2724 = ~next_sys_fair<1>_out  & ~n2723;
  assign n2725 = ~n2674 & ~n2724;
  assign n2726 = reg_i_hlock0_out & ~n2725;
  assign n2727 = ~n2562 & ~n2625;
  assign n2728 = ~next_sys_fair<1>_out  & ~n2727;
  assign n2729 = ~n2682 & ~n2728;
  assign n2730 = ~reg_i_hlock0_out & ~n2729;
  assign n2731 = ~n2726 & ~n2730;
  assign n2732 = ~reg_controllable_hmaster2_out & ~n2731;
  assign n2733 = ~n2722 & ~n2732;
  assign n2734 = reg_controllable_hmaster1_out & ~n2733;
  assign n2735 = ~reg_controllable_hmaster1_out & ~n2720;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = ~reg_controllable_hmaster0_out & ~n2736;
  assign n2738 = ~n2721 & ~n2737;
  assign n2739 = next_sys_fair<2>_out  & ~n2738;
  assign n2740 = ~reg_controllable_hmaster0_out & ~n2703;
  assign n2741 = ~n2603 & ~n2740;
  assign n2742 = ~next_sys_fair<2>_out  & ~n2741;
  assign n2743 = ~n2739 & ~n2742;
  assign n2744 = reg_controllable_hgrant2_out & ~n2743;
  assign n2745 = reg_controllable_hgrant1_out & ~n2524;
  assign n2746 = reg_controllable_hmastlock_out & ~n719;
  assign n2747 = reg_controllable_locked_out & ~n2746;
  assign n2748 = ~next_env_fair_out & ~n181;
  assign n2749 = ~next_env_fair_out & ~n2748;
  assign n2750 = ~fair_cnt<2>_out  & ~n2749;
  assign n2751 = ~fair_cnt<2>_out  & ~n2750;
  assign n2752 = reg_controllable_hmastlock_out & ~n2751;
  assign n2753 = ~n728 & ~n2752;
  assign n2754 = ~reg_controllable_locked_out & ~n2753;
  assign n2755 = ~n2747 & ~n2754;
  assign n2756 = ~reg_controllable_hgrant1_out & ~n2755;
  assign n2757 = ~n2745 & ~n2756;
  assign n2758 = ~next_sys_fair<0>_out  & ~n2757;
  assign n2759 = ~next_sys_fair<0>_out  & ~n2758;
  assign n2760 = next_sys_fair<1>_out  & ~n2759;
  assign n2761 = ~next_sys_fair<1>_out  & ~n2757;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = reg_i_hlock0_out & ~n2762;
  assign n2764 = reg_controllable_hgrant1_out & ~n2532;
  assign n2765 = reg_controllable_hmastlock_out & ~n738;
  assign n2766 = reg_controllable_hmastlock_out & ~n2765;
  assign n2767 = reg_controllable_locked_out & ~n2766;
  assign n2768 = ~reg_controllable_hmastlock_out & ~n738;
  assign n2769 = ~n285 & ~n2768;
  assign n2770 = ~reg_controllable_locked_out & ~n2769;
  assign n2771 = ~n2767 & ~n2770;
  assign n2772 = ~reg_controllable_hgrant1_out & ~n2771;
  assign n2773 = ~n2764 & ~n2772;
  assign n2774 = ~next_sys_fair<0>_out  & ~n2773;
  assign n2775 = ~next_sys_fair<0>_out  & ~n2774;
  assign n2776 = next_sys_fair<1>_out  & ~n2775;
  assign n2777 = ~next_sys_fair<1>_out  & ~n2773;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = ~reg_i_hlock0_out & ~n2778;
  assign n2780 = ~n2763 & ~n2779;
  assign n2781 = reg_controllable_hmaster2_out & ~n2780;
  assign n2782 = ~reg_controllable_locked_out & ~n2751;
  assign n2783 = ~reg_controllable_locked_out & ~n2782;
  assign n2784 = ~reg_controllable_hgrant1_out & ~n2783;
  assign n2785 = ~n2745 & ~n2784;
  assign n2786 = ~next_sys_fair<0>_out  & ~n2785;
  assign n2787 = ~next_sys_fair<0>_out  & ~n2786;
  assign n2788 = next_sys_fair<1>_out  & ~n2787;
  assign n2789 = ~next_sys_fair<1>_out  & ~n2785;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = reg_i_hlock0_out & ~n2790;
  assign n2792 = ~next_sys_fair<0>_out  & ~n2532;
  assign n2793 = ~next_sys_fair<0>_out  & ~n2792;
  assign n2794 = next_sys_fair<1>_out  & ~n2793;
  assign n2795 = ~next_sys_fair<1>_out  & ~n2532;
  assign n2796 = ~n2794 & ~n2795;
  assign n2797 = ~reg_i_hlock0_out & ~n2796;
  assign n2798 = ~n2791 & ~n2797;
  assign n2799 = ~reg_controllable_hmaster2_out & ~n2798;
  assign n2800 = ~n2781 & ~n2799;
  assign n2801 = reg_controllable_hmaster1_out & ~n2800;
  assign n2802 = reg_controllable_hgrant1_out & ~n2553;
  assign n2803 = ~n2784 & ~n2802;
  assign n2804 = ~next_sys_fair<0>_out  & ~n2803;
  assign n2805 = ~next_sys_fair<0>_out  & ~n2804;
  assign n2806 = next_sys_fair<1>_out  & ~n2805;
  assign n2807 = ~next_sys_fair<1>_out  & ~n2803;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = reg_i_hlock0_out & ~n2808;
  assign n2810 = reg_controllable_hgrant1_out & ~n2570;
  assign n2811 = ~n2533 & ~n2810;
  assign n2812 = ~next_sys_fair<0>_out  & ~n2811;
  assign n2813 = ~next_sys_fair<0>_out  & ~n2812;
  assign n2814 = next_sys_fair<1>_out  & ~n2813;
  assign n2815 = ~next_sys_fair<1>_out  & ~n2811;
  assign n2816 = ~n2814 & ~n2815;
  assign n2817 = ~reg_i_hlock0_out & ~n2816;
  assign n2818 = ~n2809 & ~n2817;
  assign n2819 = ~reg_controllable_hmaster2_out & ~n2818;
  assign n2820 = ~n2781 & ~n2819;
  assign n2821 = ~reg_controllable_hmaster1_out & ~n2820;
  assign n2822 = ~n2801 & ~n2821;
  assign n2823 = reg_controllable_hmaster0_out & ~n2822;
  assign n2824 = ~reg_controllable_hmaster1_out & ~n2798;
  assign n2825 = ~n2801 & ~n2824;
  assign n2826 = ~reg_controllable_hmaster0_out & ~n2825;
  assign n2827 = ~n2823 & ~n2826;
  assign n2828 = next_sys_fair<2>_out  & ~n2827;
  assign n2829 = reg_controllable_hgrant1_out & ~n2513;
  assign n2830 = ~n2756 & ~n2829;
  assign n2831 = next_sys_fair<0>_out  & ~n2830;
  assign n2832 = reg_controllable_hgrant1_out & ~n2588;
  assign n2833 = reg_controllable_hmastlock_out & ~n702;
  assign n2834 = reg_controllable_locked_out & ~n2833;
  assign n2835 = ~n705 & ~n1890;
  assign n2836 = ~reg_controllable_locked_out & ~n2835;
  assign n2837 = ~n2834 & ~n2836;
  assign n2838 = ~reg_controllable_hgrant1_out & ~n2837;
  assign n2839 = ~n2832 & ~n2838;
  assign n2840 = ~next_sys_fair<0>_out  & ~n2839;
  assign n2841 = ~n2831 & ~n2840;
  assign n2842 = next_sys_fair<1>_out  & ~n2841;
  assign n2843 = reg_controllable_hmastlock_out & ~n872;
  assign n2844 = reg_controllable_locked_out & ~n2843;
  assign n2845 = ~n232 & ~n883;
  assign n2846 = ~reg_controllable_locked_out & ~n2845;
  assign n2847 = ~n2844 & ~n2846;
  assign n2848 = ~reg_controllable_hgrant1_out & ~n2847;
  assign n2849 = ~n2829 & ~n2848;
  assign n2850 = next_sys_fair<0>_out  & ~n2849;
  assign n2851 = reg_controllable_hmastlock_out & ~n897;
  assign n2852 = reg_controllable_locked_out & ~n2851;
  assign n2853 = ~n232 & ~n902;
  assign n2854 = ~reg_controllable_locked_out & ~n2853;
  assign n2855 = ~n2852 & ~n2854;
  assign n2856 = ~reg_controllable_hgrant1_out & ~n2855;
  assign n2857 = ~n2829 & ~n2856;
  assign n2858 = ~next_sys_fair<0>_out  & ~n2857;
  assign n2859 = ~n2850 & ~n2858;
  assign n2860 = ~next_sys_fair<1>_out  & ~n2859;
  assign n2861 = ~n2842 & ~n2860;
  assign n2862 = reg_i_hlock0_out & ~n2861;
  assign n2863 = reg_controllable_hgrant1_out & ~n1404;
  assign n2864 = ~n2772 & ~n2863;
  assign n2865 = next_sys_fair<0>_out  & ~n2864;
  assign n2866 = reg_controllable_hgrant1_out & ~n1417;
  assign n2867 = reg_controllable_hmastlock_out & ~n704;
  assign n2868 = reg_controllable_hmastlock_out & ~n2867;
  assign n2869 = reg_controllable_locked_out & ~n2868;
  assign n2870 = ~n2836 & ~n2869;
  assign n2871 = ~reg_controllable_hgrant1_out & ~n2870;
  assign n2872 = ~n2866 & ~n2871;
  assign n2873 = ~next_sys_fair<0>_out  & ~n2872;
  assign n2874 = ~n2865 & ~n2873;
  assign n2875 = next_sys_fair<1>_out  & ~n2874;
  assign n2876 = reg_controllable_hmastlock_out & ~n1238;
  assign n2877 = reg_controllable_locked_out & ~n2876;
  assign n2878 = ~n2846 & ~n2877;
  assign n2879 = ~reg_controllable_hgrant1_out & ~n2878;
  assign n2880 = ~n2863 & ~n2879;
  assign n2881 = next_sys_fair<0>_out  & ~n2880;
  assign n2882 = reg_controllable_hmastlock_out & ~n1250;
  assign n2883 = reg_controllable_locked_out & ~n2882;
  assign n2884 = ~n2854 & ~n2883;
  assign n2885 = ~reg_controllable_hgrant1_out & ~n2884;
  assign n2886 = ~n2863 & ~n2885;
  assign n2887 = ~next_sys_fair<0>_out  & ~n2886;
  assign n2888 = ~n2881 & ~n2887;
  assign n2889 = ~next_sys_fair<1>_out  & ~n2888;
  assign n2890 = ~n2875 & ~n2889;
  assign n2891 = ~reg_i_hlock0_out & ~n2890;
  assign n2892 = ~n2862 & ~n2891;
  assign n2893 = reg_controllable_hmaster2_out & ~n2892;
  assign n2894 = ~n2784 & ~n2829;
  assign n2895 = next_sys_fair<0>_out  & ~n2894;
  assign n2896 = ~reg_controllable_locked_out & ~n1903;
  assign n2897 = ~reg_controllable_hgrant1_out & ~n2896;
  assign n2898 = ~n2832 & ~n2897;
  assign n2899 = ~next_sys_fair<0>_out  & ~n2898;
  assign n2900 = ~n2895 & ~n2899;
  assign n2901 = next_sys_fair<1>_out  & ~n2900;
  assign n2902 = ~n1405 & ~n2829;
  assign n2903 = ~next_sys_fair<1>_out  & ~n2902;
  assign n2904 = ~n2901 & ~n2903;
  assign n2905 = reg_i_hlock0_out & ~n2904;
  assign n2906 = ~n2533 & ~n2863;
  assign n2907 = next_sys_fair<0>_out  & ~n2906;
  assign n2908 = ~n2866 & ~n2897;
  assign n2909 = ~next_sys_fair<0>_out  & ~n2908;
  assign n2910 = ~n2907 & ~n2909;
  assign n2911 = next_sys_fair<1>_out  & ~n2910;
  assign n2912 = ~next_sys_fair<1>_out  & ~n1404;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = ~reg_i_hlock0_out & ~n2913;
  assign n2915 = ~n2905 & ~n2914;
  assign n2916 = ~reg_controllable_hmaster2_out & ~n2915;
  assign n2917 = ~n2893 & ~n2916;
  assign n2918 = reg_controllable_hmaster1_out & ~n2917;
  assign n2919 = reg_controllable_hgrant1_out & ~n2544;
  assign n2920 = ~n2784 & ~n2919;
  assign n2921 = next_sys_fair<0>_out  & ~n2920;
  assign n2922 = reg_controllable_hgrant1_out & ~n2609;
  assign n2923 = ~n2897 & ~n2922;
  assign n2924 = ~next_sys_fair<0>_out  & ~n2923;
  assign n2925 = ~n2921 & ~n2924;
  assign n2926 = next_sys_fair<1>_out  & ~n2925;
  assign n2927 = reg_controllable_hgrant1_out & ~n2617;
  assign n2928 = ~n1405 & ~n2927;
  assign n2929 = next_sys_fair<0>_out  & ~n2928;
  assign n2930 = ~n1405 & ~n2919;
  assign n2931 = ~next_sys_fair<0>_out  & ~n2930;
  assign n2932 = ~n2929 & ~n2931;
  assign n2933 = ~next_sys_fair<1>_out  & ~n2932;
  assign n2934 = ~n2926 & ~n2933;
  assign n2935 = reg_i_hlock0_out & ~n2934;
  assign n2936 = reg_controllable_hgrant1_out & ~n2559;
  assign n2937 = ~n2533 & ~n2936;
  assign n2938 = next_sys_fair<0>_out  & ~n2937;
  assign n2939 = reg_controllable_hgrant1_out & ~n2626;
  assign n2940 = ~n2897 & ~n2939;
  assign n2941 = ~next_sys_fair<0>_out  & ~n2940;
  assign n2942 = ~n2938 & ~n2941;
  assign n2943 = next_sys_fair<1>_out  & ~n2942;
  assign n2944 = reg_controllable_hgrant1_out & ~n2632;
  assign n2945 = ~n1405 & ~n2944;
  assign n2946 = next_sys_fair<0>_out  & ~n2945;
  assign n2947 = ~n1405 & ~n2936;
  assign n2948 = ~next_sys_fair<0>_out  & ~n2947;
  assign n2949 = ~n2946 & ~n2948;
  assign n2950 = ~next_sys_fair<1>_out  & ~n2949;
  assign n2951 = ~n2943 & ~n2950;
  assign n2952 = ~reg_i_hlock0_out & ~n2951;
  assign n2953 = ~n2935 & ~n2952;
  assign n2954 = ~reg_controllable_hmaster2_out & ~n2953;
  assign n2955 = ~n2893 & ~n2954;
  assign n2956 = ~reg_controllable_hmaster1_out & ~n2955;
  assign n2957 = ~n2918 & ~n2956;
  assign n2958 = reg_controllable_hmaster0_out & ~n2957;
  assign n2959 = ~reg_controllable_hmaster1_out & ~n2915;
  assign n2960 = ~n2918 & ~n2959;
  assign n2961 = ~reg_controllable_hmaster0_out & ~n2960;
  assign n2962 = ~n2958 & ~n2961;
  assign n2963 = ~next_sys_fair<2>_out  & ~n2962;
  assign n2964 = ~n2828 & ~n2963;
  assign n2965 = ~reg_controllable_hgrant2_out & ~n2964;
  assign n2966 = ~n2744 & ~n2965;
  assign n2967 = ~reg_controllable_hgrant3_out & ~n2966;
  assign n2968 = ~n2711 & ~n2967;
  assign n2969 = ~reg_controllable_hgrant4_out & ~n2968;
  assign n2970 = ~n2654 & ~n2969;
  assign n2971 = reg_controllable_nhgrant0_out & ~n2970;
  assign n2972 = ~n196 & ~n2523;
  assign n2973 = ~reg_controllable_hgrant1_out & ~n2972;
  assign n2974 = ~reg_controllable_hgrant1_out & ~n2973;
  assign n2975 = ~next_sys_fair<0>_out  & ~n2974;
  assign n2976 = ~next_sys_fair<0>_out  & ~n2975;
  assign n2977 = next_sys_fair<1>_out  & ~n2976;
  assign n2978 = ~next_sys_fair<1>_out  & ~n2974;
  assign n2979 = ~n2977 & ~n2978;
  assign n2980 = reg_i_hlock0_out & ~n2979;
  assign n2981 = ~n2535 & ~n2665;
  assign n2982 = ~reg_i_hlock0_out & ~n2981;
  assign n2983 = ~n2980 & ~n2982;
  assign n2984 = reg_controllable_hmaster0_out & ~n2983;
  assign n2985 = reg_controllable_hmaster1_out & ~n2983;
  assign n2986 = reg_controllable_hmaster2_out & ~n2983;
  assign n2987 = ~n284 & ~n2552;
  assign n2988 = ~reg_controllable_hgrant1_out & ~n2987;
  assign n2989 = ~reg_controllable_hgrant1_out & ~n2988;
  assign n2990 = ~next_sys_fair<0>_out  & ~n2989;
  assign n2991 = ~next_sys_fair<0>_out  & ~n2990;
  assign n2992 = next_sys_fair<1>_out  & ~n2991;
  assign n2993 = ~next_sys_fair<1>_out  & ~n2989;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = reg_i_hlock0_out & ~n2994;
  assign n2996 = ~n288 & ~n2566;
  assign n2997 = ~reg_controllable_hgrant1_out & ~n2996;
  assign n2998 = ~reg_controllable_hgrant1_out & ~n2997;
  assign n2999 = ~next_sys_fair<0>_out  & ~n2998;
  assign n3000 = ~next_sys_fair<0>_out  & ~n2999;
  assign n3001 = next_sys_fair<1>_out  & ~n3000;
  assign n3002 = ~next_sys_fair<1>_out  & ~n2998;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = ~reg_i_hlock0_out & ~n3003;
  assign n3005 = ~n2995 & ~n3004;
  assign n3006 = ~reg_controllable_hmaster2_out & ~n3005;
  assign n3007 = ~n2986 & ~n3006;
  assign n3008 = ~reg_controllable_hmaster1_out & ~n3007;
  assign n3009 = ~n2985 & ~n3008;
  assign n3010 = ~reg_controllable_hmaster0_out & ~n3009;
  assign n3011 = ~n2984 & ~n3010;
  assign n3012 = next_sys_fair<2>_out  & ~n3011;
  assign n3013 = next_sys_fair<0>_out  & ~n2974;
  assign n3014 = ~reg_controllable_hgrant1_out & ~n176;
  assign n3015 = ~reg_controllable_hgrant1_out & ~n3014;
  assign n3016 = ~next_sys_fair<0>_out  & ~n3015;
  assign n3017 = ~n3013 & ~n3016;
  assign n3018 = next_sys_fair<1>_out  & ~n3017;
  assign n3019 = ~next_sys_fair<1>_out  & ~n3015;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = reg_i_hlock0_out & ~n3020;
  assign n3022 = next_sys_fair<1>_out  & ~n2716;
  assign n3023 = ~n1656 & ~n3022;
  assign n3024 = ~reg_i_hlock0_out & ~n3023;
  assign n3025 = ~n3021 & ~n3024;
  assign n3026 = reg_controllable_hmaster0_out & ~n3025;
  assign n3027 = reg_controllable_hmaster1_out & ~n3025;
  assign n3028 = reg_controllable_hmaster2_out & ~n3025;
  assign n3029 = next_sys_fair<0>_out  & ~n2989;
  assign n3030 = ~n231 & ~n2543;
  assign n3031 = ~reg_controllable_hgrant1_out & ~n3030;
  assign n3032 = ~reg_controllable_hgrant1_out & ~n3031;
  assign n3033 = ~next_sys_fair<0>_out  & ~n3032;
  assign n3034 = ~n3029 & ~n3033;
  assign n3035 = next_sys_fair<1>_out  & ~n3034;
  assign n3036 = ~n321 & ~n2616;
  assign n3037 = ~reg_controllable_hgrant1_out & ~n3036;
  assign n3038 = ~reg_controllable_hgrant1_out & ~n3037;
  assign n3039 = next_sys_fair<0>_out  & ~n3038;
  assign n3040 = ~n342 & ~n2543;
  assign n3041 = ~reg_controllable_hgrant1_out & ~n3040;
  assign n3042 = ~reg_controllable_hgrant1_out & ~n3041;
  assign n3043 = ~next_sys_fair<0>_out  & ~n3042;
  assign n3044 = ~n3039 & ~n3043;
  assign n3045 = ~next_sys_fair<1>_out  & ~n3044;
  assign n3046 = ~n3035 & ~n3045;
  assign n3047 = reg_i_hlock0_out & ~n3046;
  assign n3048 = next_sys_fair<0>_out  & ~n2998;
  assign n3049 = ~n1841 & ~n3048;
  assign n3050 = next_sys_fair<1>_out  & ~n3049;
  assign n3051 = ~n1770 & ~n3050;
  assign n3052 = ~reg_i_hlock0_out & ~n3051;
  assign n3053 = ~n3047 & ~n3052;
  assign n3054 = ~reg_controllable_hmaster2_out & ~n3053;
  assign n3055 = ~n3028 & ~n3054;
  assign n3056 = ~reg_controllable_hmaster1_out & ~n3055;
  assign n3057 = ~n3027 & ~n3056;
  assign n3058 = ~reg_controllable_hmaster0_out & ~n3057;
  assign n3059 = ~n3026 & ~n3058;
  assign n3060 = ~next_sys_fair<2>_out  & ~n3059;
  assign n3061 = ~n3012 & ~n3060;
  assign n3062 = ~reg_controllable_hgrant2_out & ~n3061;
  assign n3063 = ~reg_controllable_hgrant2_out & ~n3062;
  assign n3064 = ~reg_controllable_hgrant3_out & ~n3063;
  assign n3065 = ~reg_controllable_hgrant3_out & ~n3064;
  assign n3066 = ~reg_controllable_hgrant4_out & ~n3065;
  assign n3067 = ~reg_controllable_hgrant4_out & ~n3066;
  assign n3068 = ~reg_controllable_nhgrant0_out & ~n3067;
  assign n3069 = ~n2971 & ~n3068;
  assign n3070 = reg_i_hready_out & ~n3069;
  assign n3071 = ~next_sys_fair<0>_out  & ~n729;
  assign n3072 = ~next_sys_fair<0>_out  & ~n3071;
  assign n3073 = next_sys_fair<1>_out  & ~n3072;
  assign n3074 = ~next_sys_fair<1>_out  & ~n729;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = reg_i_hlock0_out & ~n3075;
  assign n3077 = ~next_sys_fair<0>_out  & ~n738;
  assign n3078 = ~next_sys_fair<0>_out  & ~n3077;
  assign n3079 = next_sys_fair<1>_out  & ~n3078;
  assign n3080 = ~next_sys_fair<1>_out  & ~n738;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = ~reg_i_hlock0_out & ~n3081;
  assign n3083 = ~n3076 & ~n3082;
  assign n3084 = reg_controllable_hmaster2_out & ~n3083;
  assign n3085 = ~next_sys_fair<0>_out  & ~n792;
  assign n3086 = ~next_sys_fair<0>_out  & ~n3085;
  assign n3087 = next_sys_fair<1>_out  & ~n3086;
  assign n3088 = next_sys_fair<0>_out  & ~n772;
  assign n3089 = ~n3085 & ~n3088;
  assign n3090 = ~next_sys_fair<1>_out  & ~n3089;
  assign n3091 = ~n3087 & ~n3090;
  assign n3092 = reg_i_hlock0_out & ~n3091;
  assign n3093 = ~next_sys_fair<0>_out  & ~n801;
  assign n3094 = ~next_sys_fair<0>_out  & ~n3093;
  assign n3095 = next_sys_fair<1>_out  & ~n3094;
  assign n3096 = next_sys_fair<0>_out  & ~n779;
  assign n3097 = ~n3093 & ~n3096;
  assign n3098 = ~next_sys_fair<1>_out  & ~n3097;
  assign n3099 = ~n3095 & ~n3098;
  assign n3100 = ~reg_i_hlock0_out & ~n3099;
  assign n3101 = ~n3092 & ~n3100;
  assign n3102 = ~reg_controllable_hmaster2_out & ~n3101;
  assign n3103 = ~n3084 & ~n3102;
  assign n3104 = reg_controllable_hmaster1_out & ~n3103;
  assign n3105 = ~next_sys_fair<1>_out  & ~n792;
  assign n3106 = ~n3087 & ~n3105;
  assign n3107 = reg_i_hlock0_out & ~n3106;
  assign n3108 = ~next_sys_fair<1>_out  & ~n801;
  assign n3109 = ~n3095 & ~n3108;
  assign n3110 = ~reg_i_hlock0_out & ~n3109;
  assign n3111 = ~n3107 & ~n3110;
  assign n3112 = ~reg_controllable_hmaster2_out & ~n3111;
  assign n3113 = ~n3084 & ~n3112;
  assign n3114 = ~reg_controllable_hmaster1_out & ~n3113;
  assign n3115 = ~n3104 & ~n3114;
  assign n3116 = reg_controllable_hmaster0_out & ~n3115;
  assign n3117 = next_sys_fair<0>_out  & ~n792;
  assign n3118 = ~next_sys_fair<0>_out  & ~n772;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = ~next_sys_fair<1>_out  & ~n3119;
  assign n3121 = ~n3087 & ~n3120;
  assign n3122 = reg_i_hlock0_out & ~n3121;
  assign n3123 = next_sys_fair<0>_out  & ~n801;
  assign n3124 = ~next_sys_fair<0>_out  & ~n779;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~next_sys_fair<1>_out  & ~n3125;
  assign n3127 = ~n3095 & ~n3126;
  assign n3128 = ~reg_i_hlock0_out & ~n3127;
  assign n3129 = ~n3122 & ~n3128;
  assign n3130 = ~reg_controllable_hmaster2_out & ~n3129;
  assign n3131 = ~n3084 & ~n3130;
  assign n3132 = reg_controllable_hmaster1_out & ~n3131;
  assign n3133 = ~next_sys_fair<0>_out  & ~n3118;
  assign n3134 = next_sys_fair<1>_out  & ~n3133;
  assign n3135 = ~n3105 & ~n3134;
  assign n3136 = reg_i_hlock0_out & ~n3135;
  assign n3137 = ~next_sys_fair<0>_out  & ~n3124;
  assign n3138 = next_sys_fair<1>_out  & ~n3137;
  assign n3139 = ~n3108 & ~n3138;
  assign n3140 = ~reg_i_hlock0_out & ~n3139;
  assign n3141 = ~n3136 & ~n3140;
  assign n3142 = reg_controllable_hmaster2_out & ~n3141;
  assign n3143 = ~next_sys_fair<0>_out  & ~n843;
  assign n3144 = ~next_sys_fair<0>_out  & ~n3143;
  assign n3145 = next_sys_fair<1>_out  & ~n3144;
  assign n3146 = ~next_sys_fair<1>_out  & ~n843;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = reg_i_hlock0_out & ~n3147;
  assign n3149 = ~next_sys_fair<0>_out  & ~n846;
  assign n3150 = ~next_sys_fair<0>_out  & ~n3149;
  assign n3151 = next_sys_fair<1>_out  & ~n3150;
  assign n3152 = ~next_sys_fair<1>_out  & ~n846;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = ~reg_i_hlock0_out & ~n3153;
  assign n3155 = ~n3148 & ~n3154;
  assign n3156 = ~reg_controllable_hmaster2_out & ~n3155;
  assign n3157 = ~n3142 & ~n3156;
  assign n3158 = ~reg_controllable_hmaster1_out & ~n3157;
  assign n3159 = ~n3132 & ~n3158;
  assign n3160 = ~reg_controllable_hmaster0_out & ~n3159;
  assign n3161 = ~n3116 & ~n3160;
  assign n3162 = next_sys_fair<2>_out  & ~n3161;
  assign n3163 = next_sys_fair<0>_out  & ~n729;
  assign n3164 = ~next_sys_fair<0>_out  & ~n706;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = next_sys_fair<1>_out  & ~n3165;
  assign n3167 = next_sys_fair<0>_out  & ~n884;
  assign n3168 = ~next_sys_fair<0>_out  & ~n903;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~next_sys_fair<1>_out  & ~n3169;
  assign n3171 = ~n3166 & ~n3170;
  assign n3172 = reg_i_hlock0_out & ~n3171;
  assign n3173 = next_sys_fair<0>_out  & ~n738;
  assign n3174 = ~next_sys_fair<0>_out  & ~n704;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = next_sys_fair<1>_out  & ~n3175;
  assign n3177 = next_sys_fair<0>_out  & ~n882;
  assign n3178 = ~next_sys_fair<0>_out  & ~n901;
  assign n3179 = ~n3177 & ~n3178;
  assign n3180 = ~next_sys_fair<1>_out  & ~n3179;
  assign n3181 = ~n3176 & ~n3180;
  assign n3182 = ~reg_i_hlock0_out & ~n3181;
  assign n3183 = ~n3172 & ~n3182;
  assign n3184 = reg_controllable_hmaster2_out & ~n3183;
  assign n3185 = ~next_sys_fair<0>_out  & ~n752;
  assign n3186 = ~n3117 & ~n3185;
  assign n3187 = next_sys_fair<1>_out  & ~n3186;
  assign n3188 = next_sys_fair<0>_out  & ~n919;
  assign n3189 = ~n3118 & ~n3188;
  assign n3190 = ~next_sys_fair<1>_out  & ~n3189;
  assign n3191 = ~n3187 & ~n3190;
  assign n3192 = reg_i_hlock0_out & ~n3191;
  assign n3193 = ~next_sys_fair<0>_out  & ~n755;
  assign n3194 = ~n3123 & ~n3193;
  assign n3195 = next_sys_fair<1>_out  & ~n3194;
  assign n3196 = next_sys_fair<0>_out  & ~n921;
  assign n3197 = ~n3124 & ~n3196;
  assign n3198 = ~next_sys_fair<1>_out  & ~n3197;
  assign n3199 = ~n3195 & ~n3198;
  assign n3200 = ~reg_i_hlock0_out & ~n3199;
  assign n3201 = ~n3192 & ~n3200;
  assign n3202 = ~reg_controllable_hmaster2_out & ~n3201;
  assign n3203 = ~n3184 & ~n3202;
  assign n3204 = reg_controllable_hmaster1_out & ~n3203;
  assign n3205 = ~n3088 & ~n3185;
  assign n3206 = next_sys_fair<1>_out  & ~n3205;
  assign n3207 = ~n3190 & ~n3206;
  assign n3208 = reg_i_hlock0_out & ~n3207;
  assign n3209 = ~n3096 & ~n3193;
  assign n3210 = next_sys_fair<1>_out  & ~n3209;
  assign n3211 = ~n3198 & ~n3210;
  assign n3212 = ~reg_i_hlock0_out & ~n3211;
  assign n3213 = ~n3208 & ~n3212;
  assign n3214 = ~reg_controllable_hmaster2_out & ~n3213;
  assign n3215 = ~n3184 & ~n3214;
  assign n3216 = ~reg_controllable_hmaster1_out & ~n3215;
  assign n3217 = ~n3204 & ~n3216;
  assign n3218 = reg_controllable_hmaster0_out & ~n3217;
  assign n3219 = reg_controllable_hmaster2_out & ~n3201;
  assign n3220 = next_sys_fair<0>_out  & ~n843;
  assign n3221 = ~next_sys_fair<0>_out  & ~n830;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = next_sys_fair<1>_out  & ~n3222;
  assign n3224 = next_sys_fair<0>_out  & ~n943;
  assign n3225 = ~next_sys_fair<0>_out  & ~n954;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = ~next_sys_fair<1>_out  & ~n3226;
  assign n3228 = ~n3223 & ~n3227;
  assign n3229 = reg_i_hlock0_out & ~n3228;
  assign n3230 = next_sys_fair<0>_out  & ~n846;
  assign n3231 = ~n2212 & ~n3230;
  assign n3232 = next_sys_fair<1>_out  & ~n3231;
  assign n3233 = ~n2325 & ~n3232;
  assign n3234 = ~reg_i_hlock0_out & ~n3233;
  assign n3235 = ~n3229 & ~n3234;
  assign n3236 = ~reg_controllable_hmaster2_out & ~n3235;
  assign n3237 = ~n3219 & ~n3236;
  assign n3238 = ~reg_controllable_hmaster1_out & ~n3237;
  assign n3239 = ~n3204 & ~n3238;
  assign n3240 = ~reg_controllable_hmaster0_out & ~n3239;
  assign n3241 = ~n3218 & ~n3240;
  assign n3242 = ~next_sys_fair<2>_out  & ~n3241;
  assign n3243 = ~n3162 & ~n3242;
  assign n3244 = ~reg_i_hready_out & ~n3243;
  assign n3245 = ~n3070 & ~n3244;
  assign n3246 = ~next_sys_fair<3>_out  & ~n3245;
  assign n3247 = ~next_sys_fair<3>_out  & ~n3246;
  assign n3248 = ~reg_i_hbusreq3_out & ~n3247;
  assign n3249 = ~n2511 & ~n3248;
  assign n3250 = ~reg_i_hbusreq2_out & ~n3249;
  assign n3251 = ~n2510 & ~n3250;
  assign n3252 = ~reg_i_hbusreq1_out & ~n3251;
  assign n3253 = ~n2509 & ~n3252;
  assign n3254 = ~reg_i_hbusreq4_out & ~n3253;
  assign n3255 = ~n2508 & ~n3254;
  assign n3256 = ~reg_i_hbusreq0_out & ~n3255;
  assign n3257 = ~n2507 & ~n3256;
  assign n3258 = ~reg_controllable_ndecide_out & ~n3257;
  assign n3259 = ~n1393 & ~n3258;
  assign n3260 = ~env_safe_err_happened_out & n3259;
  assign n3261 = ~env_safe_err_happened_out & ~n3260;
  assign n3262 = n55 & ~n3261;
  assign n3263 = n55 & ~n3262;
  assign n3264 = n55 & reg_stateG10_4_out;
  assign n3265 = controllable_hgrant4 & ~n3264;
  assign n3266 = ~i_hbusreq4 & ~n3265;
  assign n3267 = i_hlock0 & ~i_hbusreq0;
  assign n3268 = i_hlock1 & ~i_hbusreq1;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = i_hlock2 & ~i_hbusreq2;
  assign n3271 = n3269 & ~n3270;
  assign n3272 = i_hlock3 & ~i_hbusreq3;
  assign n3273 = n3271 & ~n3272;
  assign n3274 = i_hlock4 & ~i_hbusreq4;
  assign n3275 = n3273 & ~n3274;
  assign n3276 = n55 & env_safe_err_happened_out;
  assign n3277 = n3275 & ~n3276;
  assign n3278 = n55 & reg_stateG10_3_out;
  assign n3279 = controllable_hgrant3 & ~n3278;
  assign n3280 = ~i_hbusreq3 & ~n3279;
  assign n3281 = n55 & next_sys_fair<3>_out ;
  assign n3282 = n55 & next_sys_fair<2>_out ;
  assign n3283 = n55 & next_sys_fair<0>_out ;
  assign n3284 = n55 & next_sys_fair<1>_out ;
  assign n3285 = n3283 & ~n3284;
  assign n3286 = n3282 & n3285;
  assign n3287 = ~n3281 & n3286;
  assign n3288 = controllable_hmaster1 & controllable_hmaster0;
  assign n3289 = ~controllable_hmaster2 & n3288;
  assign n3290 = i_hbusreq3 & ~n3289;
  assign n3291 = n3287 & ~n3290;
  assign n3292 = ~n3283 & ~n3284;
  assign n3293 = n3282 & n3292;
  assign n3294 = ~n3281 & n3293;
  assign n3295 = controllable_hmaster1 & ~controllable_hmaster0;
  assign n3296 = ~controllable_hmaster2 & n3295;
  assign n3297 = i_hbusreq2 & ~n3296;
  assign n3298 = n3294 & ~n3297;
  assign n3299 = n3283 & n3284;
  assign n3300 = ~n3282 & n3299;
  assign n3301 = ~n3281 & n3300;
  assign n3302 = ~controllable_hmaster1 & controllable_hmaster0;
  assign n3303 = ~controllable_hmaster2 & n3302;
  assign n3304 = i_hbusreq1 & ~n3303;
  assign n3305 = n3301 & ~n3304;
  assign n3306 = ~n3298 & ~n3305;
  assign n3307 = ~n3291 & n3306;
  assign n3308 = ~n3283 & n3284;
  assign n3309 = n3282 & n3308;
  assign n3310 = ~n3281 & n3309;
  assign n3311 = ~controllable_hmaster1 & ~controllable_hmaster0;
  assign n3312 = controllable_hmaster2 & n3311;
  assign n3313 = i_hbusreq4 & ~n3312;
  assign n3314 = n3310 & ~n3313;
  assign n3315 = ~n3282 & n3308;
  assign n3316 = ~n3281 & n3315;
  assign n3317 = ~controllable_hmaster2 & n3311;
  assign n3318 = i_hbusreq0 & ~n3317;
  assign n3319 = n3316 & ~n3318;
  assign n3320 = n55 & reg_stateG2_out;
  assign n3321 = ~n3282 & n3292;
  assign n3322 = ~n3281 & n3321;
  assign n3323 = ~n3320 & n3322;
  assign n3324 = n55 & reg_stateG3_0_out;
  assign n3325 = n55 & reg_stateG3_1_out;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = n55 & reg_stateG3_2_out;
  assign n3328 = n3326 & ~n3327;
  assign n3329 = ~n3282 & n3285;
  assign n3330 = ~n3281 & n3329;
  assign n3331 = n3328 & n3330;
  assign n3332 = ~n3323 & ~n3331;
  assign n3333 = ~n3319 & n3332;
  assign n3334 = n3307 & n3333;
  assign n3335 = ~n3314 & n3334;
  assign n3336 = n3282 & n3335;
  assign n3337 = n3307 & ~n3336;
  assign n3338 = n3284 & n3335;
  assign n3339 = ~n3291 & ~n3319;
  assign n3340 = ~n3331 & n3339;
  assign n3341 = ~n3338 & n3340;
  assign n3342 = n3283 & n3335;
  assign n3343 = ~n3298 & ~n3319;
  assign n3344 = ~n3323 & n3343;
  assign n3345 = ~n3342 & n3344;
  assign n3346 = n55 & fair_cnt<0>_out ;
  assign n3347 = n55 & next_env_fair_out;
  assign n3348 = i_hready & n3347;
  assign n3349 = n3346 & n3348;
  assign n3350 = n55 & fair_cnt<1>_out ;
  assign n3351 = n3349 & n3350;
  assign n3352 = n55 & fair_cnt<2>_out ;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = n3351 & n3352;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = n3335 & n3355;
  assign n3357 = ~n3349 & ~n3350;
  assign n3358 = ~n3351 & ~n3357;
  assign n3359 = n3335 & n3358;
  assign n3360 = ~n3346 & ~n3348;
  assign n3361 = ~n3349 & ~n3360;
  assign n3362 = n3335 & n3361;
  assign n3363 = n55 & reg_stateA1_out;
  assign n3364 = controllable_hmastlock & ~n3363;
  assign n3365 = ~i_hburst1 & ~i_hburst0;
  assign n3366 = n3364 & n3365;
  assign n3367 = controllable_busreq & n3363;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = controllable_busreq & n3320;
  assign n3370 = ~controllable_nstart & controllable_hmastlock;
  assign n3371 = ~i_hburst0 & n3370;
  assign n3372 = ~i_hburst1 & ~n3320;
  assign n3373 = n3371 & n3372;
  assign n3374 = ~n3369 & ~n3373;
  assign n3375 = ~n3347 & ~n3363;
  assign n3376 = ~i_hready & n3347;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = n3335 & ~n3377;
  assign n3379 = ~i_hready & controllable_ndecide;
  assign n3380 = ~i_hready & ~n3379;
  assign n3381 = controllable_hmaster1 & ~n3380;
  assign n3382 = controllable_hmaster0 & ~n3380;
  assign n3383 = controllable_hmaster0 & ~n3382;
  assign n3384 = ~controllable_hmaster1 & ~n3383;
  assign n3385 = ~n3381 & ~n3384;
  assign n3386 = i_hbusreq3 & ~n3385;
  assign n3387 = i_hbusreq2 & ~n3380;
  assign n3388 = i_hbusreq4 & ~n3380;
  assign n3389 = i_hbusreq0 & ~n3380;
  assign n3390 = ~i_hbusreq1 & ~controllable_ndecide;
  assign n3391 = ~controllable_ndecide & ~n3390;
  assign n3392 = ~i_hready & ~n3391;
  assign n3393 = ~i_hready & ~n3392;
  assign n3394 = ~i_hbusreq0 & ~n3393;
  assign n3395 = ~n3389 & ~n3394;
  assign n3396 = ~i_hbusreq4 & ~n3395;
  assign n3397 = ~n3388 & ~n3396;
  assign n3398 = ~i_hbusreq2 & ~n3397;
  assign n3399 = ~n3387 & ~n3398;
  assign n3400 = controllable_hmaster1 & ~n3399;
  assign n3401 = controllable_hmaster0 & ~n3399;
  assign n3402 = controllable_hmaster0 & ~n3401;
  assign n3403 = ~controllable_hmaster1 & ~n3402;
  assign n3404 = ~n3400 & ~n3403;
  assign n3405 = ~i_hbusreq3 & ~n3404;
  assign n3406 = ~n3386 & ~n3405;
  assign n3407 = controllable_hmaster2 & ~n3406;
  assign n3408 = controllable_hmaster2 & ~n3407;
  assign n3409 = controllable_hgrant3 & ~n3408;
  assign n3410 = controllable_hgrant2 & ~n3380;
  assign n3411 = controllable_hgrant4 & ~n3380;
  assign n3412 = controllable_locked & controllable_hmastlock;
  assign n3413 = ~controllable_locked & ~controllable_hmastlock;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~controllable_hgrant1 & n3414;
  assign n3416 = ~controllable_hgrant1 & ~n3415;
  assign n3417 = i_hready & ~n3416;
  assign n3418 = controllable_ndecide & ~n3416;
  assign n3419 = ~i_hready & n3418;
  assign n3420 = ~n3417 & ~n3419;
  assign n3421 = ~controllable_hgrant4 & ~n3420;
  assign n3422 = ~n3411 & ~n3421;
  assign n3423 = ~controllable_hgrant2 & ~n3422;
  assign n3424 = ~n3410 & ~n3423;
  assign n3425 = controllable_hmaster1 & ~n3424;
  assign n3426 = controllable_hmaster0 & ~n3424;
  assign n3427 = controllable_hmaster0 & ~n3426;
  assign n3428 = ~controllable_hmaster1 & ~n3427;
  assign n3429 = ~n3425 & ~n3428;
  assign n3430 = i_hbusreq3 & ~n3429;
  assign n3431 = controllable_hgrant2 & ~n3399;
  assign n3432 = i_hbusreq2 & ~n3422;
  assign n3433 = controllable_hgrant4 & ~n3397;
  assign n3434 = i_hbusreq4 & ~n3420;
  assign n3435 = i_hbusreq0 & ~n3420;
  assign n3436 = i_hbusreq1 & ~n3416;
  assign n3437 = i_hbusreq1 & ~n3436;
  assign n3438 = ~controllable_ndecide & ~n3437;
  assign n3439 = ~n3418 & ~n3438;
  assign n3440 = i_hready & ~n3439;
  assign n3441 = ~n3390 & ~n3418;
  assign n3442 = ~i_hready & ~n3441;
  assign n3443 = ~n3440 & ~n3442;
  assign n3444 = ~i_hbusreq0 & ~n3443;
  assign n3445 = ~n3435 & ~n3444;
  assign n3446 = ~i_hbusreq4 & ~n3445;
  assign n3447 = ~n3434 & ~n3446;
  assign n3448 = ~controllable_hgrant4 & ~n3447;
  assign n3449 = ~n3433 & ~n3448;
  assign n3450 = ~i_hbusreq2 & ~n3449;
  assign n3451 = ~n3432 & ~n3450;
  assign n3452 = ~controllable_hgrant2 & ~n3451;
  assign n3453 = ~n3431 & ~n3452;
  assign n3454 = controllable_hmaster1 & ~n3453;
  assign n3455 = controllable_hmaster0 & ~n3453;
  assign n3456 = controllable_hmaster0 & ~n3455;
  assign n3457 = ~controllable_hmaster1 & ~n3456;
  assign n3458 = ~n3454 & ~n3457;
  assign n3459 = ~i_hbusreq3 & ~n3458;
  assign n3460 = ~n3430 & ~n3459;
  assign n3461 = controllable_hmaster2 & ~n3460;
  assign n3462 = controllable_hmaster2 & ~n3461;
  assign n3463 = ~controllable_hgrant3 & ~n3462;
  assign n3464 = ~n3409 & ~n3463;
  assign n3465 = controllable_nhgrant0 & ~n3464;
  assign n3466 = ~controllable_nhgrant0 & ~n3408;
  assign n3467 = ~n3465 & ~n3466;
  assign n3468 = ~n3378 & ~n3467;
  assign n3469 = ~n3378 & ~n3468;
  assign n3470 = ~n3374 & ~n3469;
  assign n3471 = n3324 & n3325;
  assign n3472 = ~n3327 & n3471;
  assign n3473 = i_hready & n3472;
  assign n3474 = i_hready & n3326;
  assign n3475 = n3327 & ~n3474;
  assign n3476 = ~n3473 & ~n3475;
  assign n3477 = n3328 & n3371;
  assign n3478 = i_hburst1 & n3477;
  assign n3479 = i_hready & n3478;
  assign n3480 = n3325 & ~n3473;
  assign n3481 = i_hready & ~n3327;
  assign n3482 = n3324 & ~n3325;
  assign n3483 = n3481 & n3482;
  assign n3484 = ~n3480 & ~n3483;
  assign n3485 = ~n3479 & n3484;
  assign n3486 = ~n3469 & ~n3485;
  assign n3487 = ~i_hready & n3478;
  assign n3488 = ~n3324 & ~n3481;
  assign n3489 = n3324 & n3481;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = ~n3326 & n3490;
  assign n3492 = ~n3487 & ~n3491;
  assign n3493 = ~n3469 & ~n3492;
  assign n3494 = controllable_hgrant1 & controllable_ndecide;
  assign n3495 = ~i_hready & n3494;
  assign n3496 = ~n3417 & ~n3495;
  assign n3497 = ~controllable_hgrant4 & ~n3496;
  assign n3498 = ~n3411 & ~n3497;
  assign n3499 = ~controllable_hgrant2 & ~n3498;
  assign n3500 = ~n3410 & ~n3499;
  assign n3501 = controllable_hmaster1 & ~n3500;
  assign n3502 = controllable_hmaster0 & ~n3500;
  assign n3503 = controllable_hmaster0 & ~n3502;
  assign n3504 = ~controllable_hmaster1 & ~n3503;
  assign n3505 = ~n3501 & ~n3504;
  assign n3506 = i_hbusreq3 & ~n3505;
  assign n3507 = i_hbusreq2 & ~n3498;
  assign n3508 = i_hbusreq4 & ~n3496;
  assign n3509 = i_hbusreq0 & ~n3496;
  assign n3510 = ~n3390 & ~n3494;
  assign n3511 = ~i_hready & ~n3510;
  assign n3512 = ~n3440 & ~n3511;
  assign n3513 = ~i_hbusreq0 & ~n3512;
  assign n3514 = ~n3509 & ~n3513;
  assign n3515 = ~i_hbusreq4 & ~n3514;
  assign n3516 = ~n3508 & ~n3515;
  assign n3517 = ~controllable_hgrant4 & ~n3516;
  assign n3518 = ~n3433 & ~n3517;
  assign n3519 = ~i_hbusreq2 & ~n3518;
  assign n3520 = ~n3507 & ~n3519;
  assign n3521 = ~controllable_hgrant2 & ~n3520;
  assign n3522 = ~n3431 & ~n3521;
  assign n3523 = controllable_hmaster1 & ~n3522;
  assign n3524 = controllable_hmaster0 & ~n3522;
  assign n3525 = controllable_hmaster0 & ~n3524;
  assign n3526 = ~controllable_hmaster1 & ~n3525;
  assign n3527 = ~n3523 & ~n3526;
  assign n3528 = ~i_hbusreq3 & ~n3527;
  assign n3529 = ~n3506 & ~n3528;
  assign n3530 = controllable_hmaster2 & ~n3529;
  assign n3531 = controllable_hmaster2 & ~n3530;
  assign n3532 = ~controllable_hgrant3 & ~n3531;
  assign n3533 = ~n3409 & ~n3532;
  assign n3534 = controllable_nhgrant0 & ~n3533;
  assign n3535 = ~n3466 & ~n3534;
  assign n3536 = ~n3378 & ~n3535;
  assign n3537 = ~n3378 & ~n3536;
  assign n3538 = n3492 & ~n3537;
  assign n3539 = ~n3493 & ~n3538;
  assign n3540 = n3485 & ~n3539;
  assign n3541 = ~n3486 & ~n3540;
  assign n3542 = ~n3476 & ~n3541;
  assign n3543 = i_hready & controllable_hgrant1;
  assign n3544 = ~n3495 & ~n3543;
  assign n3545 = ~controllable_hgrant4 & ~n3544;
  assign n3546 = ~n3411 & ~n3545;
  assign n3547 = ~controllable_hgrant2 & ~n3546;
  assign n3548 = ~n3410 & ~n3547;
  assign n3549 = controllable_hmaster1 & ~n3548;
  assign n3550 = controllable_hmaster0 & ~n3548;
  assign n3551 = i_hready & ~n3543;
  assign n3552 = ~controllable_hgrant4 & ~n3551;
  assign n3553 = ~controllable_hgrant4 & ~n3552;
  assign n3554 = ~controllable_hgrant2 & ~n3553;
  assign n3555 = ~controllable_hgrant2 & ~n3554;
  assign n3556 = ~controllable_hmaster0 & ~n3555;
  assign n3557 = ~n3550 & ~n3556;
  assign n3558 = ~controllable_hmaster1 & ~n3557;
  assign n3559 = ~n3549 & ~n3558;
  assign n3560 = i_hbusreq3 & ~n3559;
  assign n3561 = i_hbusreq2 & ~n3546;
  assign n3562 = i_hbusreq4 & ~n3544;
  assign n3563 = i_hbusreq0 & ~n3544;
  assign n3564 = i_hbusreq1 & controllable_hgrant1;
  assign n3565 = i_hbusreq1 & ~n3564;
  assign n3566 = ~controllable_ndecide & ~n3565;
  assign n3567 = ~n3494 & ~n3566;
  assign n3568 = i_hready & ~n3567;
  assign n3569 = ~n3511 & ~n3568;
  assign n3570 = ~i_hbusreq0 & ~n3569;
  assign n3571 = ~n3563 & ~n3570;
  assign n3572 = ~i_hbusreq4 & ~n3571;
  assign n3573 = ~n3562 & ~n3572;
  assign n3574 = ~controllable_hgrant4 & ~n3573;
  assign n3575 = ~n3433 & ~n3574;
  assign n3576 = ~i_hbusreq2 & ~n3575;
  assign n3577 = ~n3561 & ~n3576;
  assign n3578 = ~controllable_hgrant2 & ~n3577;
  assign n3579 = ~n3431 & ~n3578;
  assign n3580 = controllable_hmaster1 & ~n3579;
  assign n3581 = controllable_hmaster0 & ~n3579;
  assign n3582 = i_hbusreq2 & ~n3553;
  assign n3583 = i_hbusreq4 & ~n3551;
  assign n3584 = i_hbusreq0 & ~n3551;
  assign n3585 = i_hready & ~n3568;
  assign n3586 = ~i_hbusreq0 & ~n3585;
  assign n3587 = ~n3584 & ~n3586;
  assign n3588 = ~i_hbusreq4 & ~n3587;
  assign n3589 = ~n3583 & ~n3588;
  assign n3590 = ~controllable_hgrant4 & ~n3589;
  assign n3591 = ~controllable_hgrant4 & ~n3590;
  assign n3592 = ~i_hbusreq2 & ~n3591;
  assign n3593 = ~n3582 & ~n3592;
  assign n3594 = ~controllable_hgrant2 & ~n3593;
  assign n3595 = ~controllable_hgrant2 & ~n3594;
  assign n3596 = ~controllable_hmaster0 & ~n3595;
  assign n3597 = ~n3581 & ~n3596;
  assign n3598 = ~controllable_hmaster1 & ~n3597;
  assign n3599 = ~n3580 & ~n3598;
  assign n3600 = ~i_hbusreq3 & ~n3599;
  assign n3601 = ~n3560 & ~n3600;
  assign n3602 = controllable_hmaster2 & ~n3601;
  assign n3603 = i_hbusreq3 & ~n3555;
  assign n3604 = ~i_hbusreq3 & ~n3595;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~controllable_hmaster2 & ~n3605;
  assign n3607 = ~n3602 & ~n3606;
  assign n3608 = ~controllable_hgrant3 & ~n3607;
  assign n3609 = ~n3409 & ~n3608;
  assign n3610 = controllable_nhgrant0 & ~n3609;
  assign n3611 = ~n3466 & ~n3610;
  assign n3612 = ~n3378 & ~n3611;
  assign n3613 = ~n3378 & ~n3612;
  assign n3614 = n3492 & ~n3613;
  assign n3615 = ~n3493 & ~n3614;
  assign n3616 = n3485 & ~n3615;
  assign n3617 = ~n3486 & ~n3616;
  assign n3618 = n3476 & ~n3617;
  assign n3619 = ~n3542 & ~n3618;
  assign n3620 = n3374 & ~n3619;
  assign n3621 = ~n3470 & ~n3620;
  assign n3622 = ~n3368 & ~n3621;
  assign n3623 = ~n3368 & ~n3622;
  assign n3624 = ~n3362 & ~n3623;
  assign n3625 = ~n3362 & ~n3624;
  assign n3626 = ~n3359 & ~n3625;
  assign n3627 = ~n3359 & ~n3626;
  assign n3628 = n3356 & ~n3627;
  assign n3629 = ~n3374 & ~n3467;
  assign n3630 = ~n3467 & ~n3485;
  assign n3631 = ~n3467 & ~n3492;
  assign n3632 = n3492 & ~n3535;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = n3485 & ~n3633;
  assign n3635 = ~n3630 & ~n3634;
  assign n3636 = ~n3476 & ~n3635;
  assign n3637 = n3492 & ~n3611;
  assign n3638 = ~n3631 & ~n3637;
  assign n3639 = n3485 & ~n3638;
  assign n3640 = ~n3630 & ~n3639;
  assign n3641 = n3476 & ~n3640;
  assign n3642 = ~n3636 & ~n3641;
  assign n3643 = n3374 & ~n3642;
  assign n3644 = ~n3629 & ~n3643;
  assign n3645 = ~n3368 & ~n3644;
  assign n3646 = ~n3368 & ~n3645;
  assign n3647 = ~n3356 & ~n3646;
  assign n3648 = ~n3628 & ~n3647;
  assign n3649 = ~n3345 & ~n3648;
  assign n3650 = n55 & reg_stateG10_2_out;
  assign n3651 = controllable_hgrant2 & ~n3650;
  assign n3652 = ~i_hbusreq2 & ~n3651;
  assign n3653 = n55 & reg_stateG10_1_out;
  assign n3654 = controllable_hgrant1 & ~n3653;
  assign n3655 = ~i_hbusreq1 & ~n3654;
  assign n3656 = ~controllable_ndecide & ~controllable_hmastlock;
  assign n3657 = ~controllable_ndecide & ~n3656;
  assign n3658 = ~i_hready & ~n3657;
  assign n3659 = ~i_hready & ~n3658;
  assign n3660 = i_hlock4 & ~n3659;
  assign n3661 = ~controllable_ndecide & controllable_hmastlock;
  assign n3662 = ~controllable_ndecide & ~n3661;
  assign n3663 = ~i_hready & ~n3662;
  assign n3664 = ~i_hready & ~n3663;
  assign n3665 = ~i_hlock4 & ~n3664;
  assign n3666 = ~n3660 & ~n3665;
  assign n3667 = ~controllable_hmaster0 & ~n3666;
  assign n3668 = ~controllable_hmaster0 & ~n3667;
  assign n3669 = ~controllable_hmaster1 & ~n3668;
  assign n3670 = ~controllable_hmaster1 & ~n3669;
  assign n3671 = i_hbusreq3 & ~n3670;
  assign n3672 = i_hbusreq2 & ~n3666;
  assign n3673 = i_hbusreq4 & ~n3666;
  assign n3674 = i_hbusreq0 & ~n3659;
  assign n3675 = i_hbusreq1 & controllable_hmastlock;
  assign n3676 = ~controllable_ndecide & ~n3675;
  assign n3677 = ~controllable_ndecide & ~n3676;
  assign n3678 = ~i_hready & ~n3677;
  assign n3679 = ~i_hready & ~n3678;
  assign n3680 = ~i_hbusreq0 & ~n3679;
  assign n3681 = ~n3674 & ~n3680;
  assign n3682 = i_hlock4 & ~n3681;
  assign n3683 = i_hbusreq0 & ~n3664;
  assign n3684 = i_hbusreq1 & ~n3675;
  assign n3685 = ~controllable_ndecide & ~n3684;
  assign n3686 = ~controllable_ndecide & ~n3685;
  assign n3687 = ~i_hready & ~n3686;
  assign n3688 = ~i_hready & ~n3687;
  assign n3689 = ~i_hbusreq0 & ~n3688;
  assign n3690 = ~n3683 & ~n3689;
  assign n3691 = ~i_hlock4 & ~n3690;
  assign n3692 = ~n3682 & ~n3691;
  assign n3693 = ~i_hbusreq4 & ~n3692;
  assign n3694 = ~n3673 & ~n3693;
  assign n3695 = ~i_hbusreq2 & ~n3694;
  assign n3696 = ~n3672 & ~n3695;
  assign n3697 = ~controllable_hmaster0 & ~n3696;
  assign n3698 = ~controllable_hmaster0 & ~n3697;
  assign n3699 = ~controllable_hmaster1 & ~n3698;
  assign n3700 = ~controllable_hmaster1 & ~n3699;
  assign n3701 = ~i_hbusreq3 & ~n3700;
  assign n3702 = ~n3671 & ~n3701;
  assign n3703 = controllable_hmaster2 & ~n3702;
  assign n3704 = controllable_hmaster2 & ~n3703;
  assign n3705 = controllable_hgrant3 & ~n3704;
  assign n3706 = controllable_hgrant2 & ~n3666;
  assign n3707 = ~controllable_hgrant1 & ~n3412;
  assign n3708 = ~controllable_hgrant1 & ~n3707;
  assign n3709 = ~controllable_ndecide & ~n3708;
  assign n3710 = ~controllable_ndecide & ~n3709;
  assign n3711 = i_hready & ~n3710;
  assign n3712 = ~n3658 & ~n3711;
  assign n3713 = i_hlock4 & ~n3712;
  assign n3714 = ~controllable_locked & controllable_hmastlock;
  assign n3715 = ~controllable_locked & ~n3714;
  assign n3716 = ~controllable_hgrant1 & ~n3715;
  assign n3717 = ~controllable_hgrant1 & ~n3716;
  assign n3718 = ~controllable_ndecide & ~n3717;
  assign n3719 = ~controllable_ndecide & ~n3718;
  assign n3720 = i_hready & ~n3719;
  assign n3721 = ~n3663 & ~n3720;
  assign n3722 = ~i_hlock4 & ~n3721;
  assign n3723 = ~n3713 & ~n3722;
  assign n3724 = controllable_hgrant4 & ~n3723;
  assign n3725 = ~controllable_hgrant4 & ~n3666;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = ~controllable_hgrant2 & ~n3726;
  assign n3728 = ~n3706 & ~n3727;
  assign n3729 = ~controllable_hmaster0 & ~n3728;
  assign n3730 = ~controllable_hmaster0 & ~n3729;
  assign n3731 = ~controllable_hmaster1 & ~n3730;
  assign n3732 = ~controllable_hmaster1 & ~n3731;
  assign n3733 = i_hbusreq3 & ~n3732;
  assign n3734 = controllable_hgrant2 & ~n3696;
  assign n3735 = i_hbusreq2 & ~n3726;
  assign n3736 = i_hbusreq4 & ~n3723;
  assign n3737 = i_hbusreq0 & ~n3712;
  assign n3738 = i_hbusreq1 & ~n3708;
  assign n3739 = i_hbusreq1 & ~n3738;
  assign n3740 = ~controllable_ndecide & ~n3739;
  assign n3741 = ~controllable_ndecide & ~n3740;
  assign n3742 = i_hready & ~n3741;
  assign n3743 = ~n3678 & ~n3742;
  assign n3744 = ~i_hbusreq0 & ~n3743;
  assign n3745 = ~n3737 & ~n3744;
  assign n3746 = i_hlock4 & ~n3745;
  assign n3747 = i_hbusreq0 & ~n3721;
  assign n3748 = i_hbusreq1 & ~n3717;
  assign n3749 = i_hbusreq1 & ~n3748;
  assign n3750 = ~controllable_ndecide & ~n3749;
  assign n3751 = ~controllable_ndecide & ~n3750;
  assign n3752 = i_hready & ~n3751;
  assign n3753 = ~n3687 & ~n3752;
  assign n3754 = ~i_hbusreq0 & ~n3753;
  assign n3755 = ~n3747 & ~n3754;
  assign n3756 = ~i_hlock4 & ~n3755;
  assign n3757 = ~n3746 & ~n3756;
  assign n3758 = ~i_hbusreq4 & ~n3757;
  assign n3759 = ~n3736 & ~n3758;
  assign n3760 = controllable_hgrant4 & ~n3759;
  assign n3761 = ~controllable_hgrant4 & ~n3694;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = ~i_hbusreq2 & ~n3762;
  assign n3764 = ~n3735 & ~n3763;
  assign n3765 = ~controllable_hgrant2 & ~n3764;
  assign n3766 = ~n3734 & ~n3765;
  assign n3767 = ~controllable_hmaster0 & ~n3766;
  assign n3768 = ~controllable_hmaster0 & ~n3767;
  assign n3769 = ~controllable_hmaster1 & ~n3768;
  assign n3770 = ~controllable_hmaster1 & ~n3769;
  assign n3771 = ~i_hbusreq3 & ~n3770;
  assign n3772 = ~n3733 & ~n3771;
  assign n3773 = controllable_hmaster2 & ~n3772;
  assign n3774 = controllable_hmaster2 & ~n3773;
  assign n3775 = ~controllable_hgrant3 & ~n3774;
  assign n3776 = ~n3705 & ~n3775;
  assign n3777 = controllable_nhgrant0 & ~n3776;
  assign n3778 = ~controllable_nhgrant0 & ~n3704;
  assign n3779 = ~n3777 & ~n3778;
  assign n3780 = ~n3281 & ~n3779;
  assign n3781 = ~n3281 & ~n3780;
  assign n3782 = n3378 & ~n3781;
  assign n3783 = n3281 & ~n3467;
  assign n3784 = ~n3382 & ~n3667;
  assign n3785 = ~controllable_hmaster1 & ~n3784;
  assign n3786 = ~n3381 & ~n3785;
  assign n3787 = i_hbusreq3 & ~n3786;
  assign n3788 = ~n3401 & ~n3697;
  assign n3789 = ~controllable_hmaster1 & ~n3788;
  assign n3790 = ~n3400 & ~n3789;
  assign n3791 = ~i_hbusreq3 & ~n3790;
  assign n3792 = ~n3787 & ~n3791;
  assign n3793 = controllable_hmaster2 & ~n3792;
  assign n3794 = controllable_hmaster2 & ~n3793;
  assign n3795 = controllable_hgrant3 & ~n3794;
  assign n3796 = ~n3426 & ~n3729;
  assign n3797 = ~controllable_hmaster1 & ~n3796;
  assign n3798 = ~n3425 & ~n3797;
  assign n3799 = i_hbusreq3 & ~n3798;
  assign n3800 = ~n3455 & ~n3767;
  assign n3801 = ~controllable_hmaster1 & ~n3800;
  assign n3802 = ~n3454 & ~n3801;
  assign n3803 = ~i_hbusreq3 & ~n3802;
  assign n3804 = ~n3799 & ~n3803;
  assign n3805 = controllable_hmaster2 & ~n3804;
  assign n3806 = controllable_hmaster2 & ~n3805;
  assign n3807 = ~controllable_hgrant3 & ~n3806;
  assign n3808 = ~n3795 & ~n3807;
  assign n3809 = controllable_nhgrant0 & ~n3808;
  assign n3810 = ~controllable_nhgrant0 & ~n3794;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = ~n3281 & ~n3811;
  assign n3813 = ~n3783 & ~n3812;
  assign n3814 = ~n3378 & ~n3813;
  assign n3815 = ~n3782 & ~n3814;
  assign n3816 = n3492 & ~n3815;
  assign n3817 = ~n3493 & ~n3816;
  assign n3818 = n3485 & ~n3817;
  assign n3819 = ~n3486 & ~n3818;
  assign n3820 = ~n3374 & ~n3819;
  assign n3821 = ~controllable_hmaster0 & ~n3380;
  assign n3822 = ~controllable_hmaster0 & ~n3821;
  assign n3823 = ~controllable_hmaster1 & ~n3822;
  assign n3824 = ~controllable_hmaster1 & ~n3823;
  assign n3825 = i_hbusreq3 & ~n3824;
  assign n3826 = i_hlock0 & ~n3393;
  assign n3827 = ~i_hlock0 & ~n3380;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~i_hbusreq0 & ~n3828;
  assign n3830 = ~n3389 & ~n3829;
  assign n3831 = ~i_hbusreq4 & ~n3830;
  assign n3832 = ~n3388 & ~n3831;
  assign n3833 = ~i_hbusreq2 & ~n3832;
  assign n3834 = ~n3387 & ~n3833;
  assign n3835 = ~controllable_hmaster0 & ~n3834;
  assign n3836 = ~controllable_hmaster0 & ~n3835;
  assign n3837 = ~controllable_hmaster1 & ~n3836;
  assign n3838 = ~controllable_hmaster1 & ~n3837;
  assign n3839 = ~i_hbusreq3 & ~n3838;
  assign n3840 = ~n3825 & ~n3839;
  assign n3841 = controllable_hmaster2 & ~n3840;
  assign n3842 = controllable_hmaster2 & ~n3841;
  assign n3843 = controllable_hgrant3 & ~n3842;
  assign n3844 = ~controllable_ndecide & ~n3416;
  assign n3845 = ~controllable_ndecide & ~n3844;
  assign n3846 = i_hready & ~n3845;
  assign n3847 = ~n3379 & ~n3846;
  assign n3848 = controllable_hgrant4 & ~n3847;
  assign n3849 = ~i_hready & ~n3495;
  assign n3850 = ~controllable_hgrant4 & ~n3849;
  assign n3851 = ~n3848 & ~n3850;
  assign n3852 = ~controllable_hgrant2 & ~n3851;
  assign n3853 = ~n3410 & ~n3852;
  assign n3854 = ~controllable_hmaster0 & ~n3853;
  assign n3855 = ~controllable_hmaster0 & ~n3854;
  assign n3856 = ~controllable_hmaster1 & ~n3855;
  assign n3857 = ~controllable_hmaster1 & ~n3856;
  assign n3858 = i_hbusreq3 & ~n3857;
  assign n3859 = controllable_hgrant2 & ~n3834;
  assign n3860 = i_hbusreq2 & ~n3851;
  assign n3861 = i_hbusreq4 & ~n3847;
  assign n3862 = i_hbusreq0 & ~n3847;
  assign n3863 = ~controllable_ndecide & ~n3438;
  assign n3864 = i_hready & ~n3863;
  assign n3865 = ~n3392 & ~n3864;
  assign n3866 = i_hlock0 & ~n3865;
  assign n3867 = ~i_hlock0 & ~n3847;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = ~i_hbusreq0 & ~n3868;
  assign n3870 = ~n3862 & ~n3869;
  assign n3871 = ~i_hbusreq4 & ~n3870;
  assign n3872 = ~n3861 & ~n3871;
  assign n3873 = controllable_hgrant4 & ~n3872;
  assign n3874 = i_hbusreq4 & ~n3849;
  assign n3875 = i_hbusreq0 & ~n3849;
  assign n3876 = ~i_hready & ~n3511;
  assign n3877 = i_hlock0 & ~n3876;
  assign n3878 = ~i_hlock0 & ~n3849;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = ~i_hbusreq0 & ~n3879;
  assign n3881 = ~n3875 & ~n3880;
  assign n3882 = ~i_hbusreq4 & ~n3881;
  assign n3883 = ~n3874 & ~n3882;
  assign n3884 = ~controllable_hgrant4 & ~n3883;
  assign n3885 = ~n3873 & ~n3884;
  assign n3886 = ~i_hbusreq2 & ~n3885;
  assign n3887 = ~n3860 & ~n3886;
  assign n3888 = ~controllable_hgrant2 & ~n3887;
  assign n3889 = ~n3859 & ~n3888;
  assign n3890 = ~controllable_hmaster0 & ~n3889;
  assign n3891 = ~controllable_hmaster0 & ~n3890;
  assign n3892 = ~controllable_hmaster1 & ~n3891;
  assign n3893 = ~controllable_hmaster1 & ~n3892;
  assign n3894 = ~i_hbusreq3 & ~n3893;
  assign n3895 = ~n3858 & ~n3894;
  assign n3896 = controllable_hmaster2 & ~n3895;
  assign n3897 = controllable_hmaster2 & ~n3896;
  assign n3898 = ~controllable_hgrant3 & ~n3897;
  assign n3899 = ~n3843 & ~n3898;
  assign n3900 = controllable_nhgrant0 & ~n3899;
  assign n3901 = ~controllable_hgrant1 & controllable_locked;
  assign n3902 = ~controllable_hgrant1 & ~n3901;
  assign n3903 = controllable_ndecide & ~n3902;
  assign n3904 = ~i_hready & n3903;
  assign n3905 = ~i_hready & ~n3904;
  assign n3906 = ~controllable_hgrant4 & ~n3905;
  assign n3907 = ~n3411 & ~n3906;
  assign n3908 = ~controllable_hgrant2 & ~n3907;
  assign n3909 = ~n3410 & ~n3908;
  assign n3910 = ~controllable_hmaster0 & ~n3909;
  assign n3911 = ~controllable_hmaster0 & ~n3910;
  assign n3912 = ~controllable_hmaster1 & ~n3911;
  assign n3913 = ~controllable_hmaster1 & ~n3912;
  assign n3914 = i_hbusreq3 & ~n3913;
  assign n3915 = i_hbusreq2 & ~n3907;
  assign n3916 = controllable_hgrant4 & ~n3832;
  assign n3917 = i_hbusreq4 & ~n3905;
  assign n3918 = i_hbusreq0 & ~n3905;
  assign n3919 = ~n3390 & ~n3903;
  assign n3920 = ~i_hready & ~n3919;
  assign n3921 = ~i_hready & ~n3920;
  assign n3922 = i_hlock0 & ~n3921;
  assign n3923 = ~i_hlock0 & ~n3905;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~i_hbusreq0 & ~n3924;
  assign n3926 = ~n3918 & ~n3925;
  assign n3927 = ~i_hbusreq4 & ~n3926;
  assign n3928 = ~n3917 & ~n3927;
  assign n3929 = ~controllable_hgrant4 & ~n3928;
  assign n3930 = ~n3916 & ~n3929;
  assign n3931 = ~i_hbusreq2 & ~n3930;
  assign n3932 = ~n3915 & ~n3931;
  assign n3933 = ~controllable_hgrant2 & ~n3932;
  assign n3934 = ~n3859 & ~n3933;
  assign n3935 = ~controllable_hmaster0 & ~n3934;
  assign n3936 = ~controllable_hmaster0 & ~n3935;
  assign n3937 = ~controllable_hmaster1 & ~n3936;
  assign n3938 = ~controllable_hmaster1 & ~n3937;
  assign n3939 = ~i_hbusreq3 & ~n3938;
  assign n3940 = ~n3914 & ~n3939;
  assign n3941 = controllable_hmaster2 & ~n3940;
  assign n3942 = controllable_hmaster2 & ~n3941;
  assign n3943 = ~controllable_hgrant3 & ~n3942;
  assign n3944 = ~n3843 & ~n3943;
  assign n3945 = ~controllable_nhgrant0 & ~n3944;
  assign n3946 = ~n3900 & ~n3945;
  assign n3947 = ~n3281 & ~n3946;
  assign n3948 = ~n3281 & ~n3947;
  assign n3949 = n3378 & ~n3948;
  assign n3950 = n3281 & ~n3535;
  assign n3951 = i_hbusreq3 & ~n3380;
  assign n3952 = ~n3401 & ~n3835;
  assign n3953 = ~controllable_hmaster1 & ~n3952;
  assign n3954 = ~n3400 & ~n3953;
  assign n3955 = ~i_hbusreq3 & ~n3954;
  assign n3956 = ~n3951 & ~n3955;
  assign n3957 = controllable_hmaster2 & ~n3956;
  assign n3958 = controllable_hmaster2 & ~n3957;
  assign n3959 = controllable_hgrant3 & ~n3958;
  assign n3960 = ~n3502 & ~n3854;
  assign n3961 = ~controllable_hmaster1 & ~n3960;
  assign n3962 = ~n3501 & ~n3961;
  assign n3963 = i_hbusreq3 & ~n3962;
  assign n3964 = ~n3524 & ~n3890;
  assign n3965 = ~controllable_hmaster1 & ~n3964;
  assign n3966 = ~n3523 & ~n3965;
  assign n3967 = ~i_hbusreq3 & ~n3966;
  assign n3968 = ~n3963 & ~n3967;
  assign n3969 = controllable_hmaster2 & ~n3968;
  assign n3970 = controllable_hmaster2 & ~n3969;
  assign n3971 = ~controllable_hgrant3 & ~n3970;
  assign n3972 = ~n3959 & ~n3971;
  assign n3973 = controllable_nhgrant0 & ~n3972;
  assign n3974 = ~n3382 & ~n3910;
  assign n3975 = ~controllable_hmaster1 & ~n3974;
  assign n3976 = ~n3381 & ~n3975;
  assign n3977 = i_hbusreq3 & ~n3976;
  assign n3978 = ~n3401 & ~n3935;
  assign n3979 = ~controllable_hmaster1 & ~n3978;
  assign n3980 = ~n3400 & ~n3979;
  assign n3981 = ~i_hbusreq3 & ~n3980;
  assign n3982 = ~n3977 & ~n3981;
  assign n3983 = controllable_hmaster2 & ~n3982;
  assign n3984 = controllable_hmaster2 & ~n3983;
  assign n3985 = ~controllable_hgrant3 & ~n3984;
  assign n3986 = ~n3959 & ~n3985;
  assign n3987 = ~controllable_nhgrant0 & ~n3986;
  assign n3988 = ~n3973 & ~n3987;
  assign n3989 = ~n3281 & ~n3988;
  assign n3990 = ~n3950 & ~n3989;
  assign n3991 = ~n3378 & ~n3990;
  assign n3992 = ~n3949 & ~n3991;
  assign n3993 = n3492 & ~n3992;
  assign n3994 = ~n3493 & ~n3993;
  assign n3995 = n3485 & ~n3994;
  assign n3996 = ~n3486 & ~n3995;
  assign n3997 = ~n3476 & ~n3996;
  assign n3998 = ~controllable_ndecide & ~n3902;
  assign n3999 = ~controllable_ndecide & ~n3998;
  assign n4000 = i_hready & ~n3999;
  assign n4001 = i_hready & ~n4000;
  assign n4002 = controllable_hgrant4 & ~n4001;
  assign n4003 = controllable_hgrant4 & ~n4002;
  assign n4004 = ~controllable_hgrant2 & ~n4003;
  assign n4005 = ~controllable_hgrant2 & ~n4004;
  assign n4006 = controllable_hmaster1 & ~n4005;
  assign n4007 = controllable_hmaster0 & ~n4005;
  assign n4008 = controllable_locked & ~n3412;
  assign n4009 = ~controllable_hgrant1 & n4008;
  assign n4010 = ~controllable_hgrant1 & ~n4009;
  assign n4011 = ~controllable_ndecide & ~n4010;
  assign n4012 = ~controllable_ndecide & ~n4011;
  assign n4013 = i_hready & ~n4012;
  assign n4014 = ~n3379 & ~n4013;
  assign n4015 = controllable_hgrant4 & ~n4014;
  assign n4016 = ~n3850 & ~n4015;
  assign n4017 = ~controllable_hgrant2 & ~n4016;
  assign n4018 = ~n3410 & ~n4017;
  assign n4019 = ~controllable_hmaster0 & ~n4018;
  assign n4020 = ~n4007 & ~n4019;
  assign n4021 = ~controllable_hmaster1 & ~n4020;
  assign n4022 = ~n4006 & ~n4021;
  assign n4023 = i_hbusreq3 & ~n4022;
  assign n4024 = i_hbusreq2 & ~n4003;
  assign n4025 = i_hbusreq4 & ~n4001;
  assign n4026 = i_hbusreq0 & ~n4001;
  assign n4027 = i_hbusreq1 & ~n3902;
  assign n4028 = i_hbusreq1 & ~n4027;
  assign n4029 = ~controllable_ndecide & ~n4028;
  assign n4030 = ~controllable_ndecide & ~n4029;
  assign n4031 = i_hready & ~n4030;
  assign n4032 = i_hready & ~n4031;
  assign n4033 = i_hlock0 & ~n4032;
  assign n4034 = ~i_hlock0 & ~n4001;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = ~i_hbusreq0 & ~n4035;
  assign n4037 = ~n4026 & ~n4036;
  assign n4038 = ~i_hbusreq4 & ~n4037;
  assign n4039 = ~n4025 & ~n4038;
  assign n4040 = controllable_hgrant4 & ~n4039;
  assign n4041 = controllable_hgrant4 & ~n4040;
  assign n4042 = ~i_hbusreq2 & ~n4041;
  assign n4043 = ~n4024 & ~n4042;
  assign n4044 = ~controllable_hgrant2 & ~n4043;
  assign n4045 = ~controllable_hgrant2 & ~n4044;
  assign n4046 = controllable_hmaster1 & ~n4045;
  assign n4047 = controllable_hmaster0 & ~n4045;
  assign n4048 = i_hbusreq2 & ~n4016;
  assign n4049 = i_hbusreq4 & ~n4014;
  assign n4050 = i_hbusreq0 & ~n4014;
  assign n4051 = i_hbusreq1 & ~n4010;
  assign n4052 = i_hbusreq1 & ~n4051;
  assign n4053 = ~controllable_ndecide & ~n4052;
  assign n4054 = ~controllable_ndecide & ~n4053;
  assign n4055 = i_hready & ~n4054;
  assign n4056 = ~n3392 & ~n4055;
  assign n4057 = i_hlock0 & ~n4056;
  assign n4058 = ~i_hlock0 & ~n4014;
  assign n4059 = ~n4057 & ~n4058;
  assign n4060 = ~i_hbusreq0 & ~n4059;
  assign n4061 = ~n4050 & ~n4060;
  assign n4062 = ~i_hbusreq4 & ~n4061;
  assign n4063 = ~n4049 & ~n4062;
  assign n4064 = controllable_hgrant4 & ~n4063;
  assign n4065 = ~n3884 & ~n4064;
  assign n4066 = ~i_hbusreq2 & ~n4065;
  assign n4067 = ~n4048 & ~n4066;
  assign n4068 = ~controllable_hgrant2 & ~n4067;
  assign n4069 = ~n3859 & ~n4068;
  assign n4070 = ~controllable_hmaster0 & ~n4069;
  assign n4071 = ~n4047 & ~n4070;
  assign n4072 = ~controllable_hmaster1 & ~n4071;
  assign n4073 = ~n4046 & ~n4072;
  assign n4074 = ~i_hbusreq3 & ~n4073;
  assign n4075 = ~n4023 & ~n4074;
  assign n4076 = controllable_hmaster2 & ~n4075;
  assign n4077 = i_hbusreq3 & ~n4005;
  assign n4078 = ~i_hbusreq3 & ~n4045;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~controllable_hmaster2 & ~n4079;
  assign n4081 = ~n4076 & ~n4080;
  assign n4082 = ~controllable_hgrant3 & ~n4081;
  assign n4083 = ~n3843 & ~n4082;
  assign n4084 = controllable_nhgrant0 & ~n4083;
  assign n4085 = ~n3945 & ~n4084;
  assign n4086 = ~n3281 & ~n4085;
  assign n4087 = ~n3281 & ~n4086;
  assign n4088 = n3378 & ~n4087;
  assign n4089 = n3281 & ~n3611;
  assign n4090 = ~n3379 & ~n4000;
  assign n4091 = controllable_hgrant4 & ~n4090;
  assign n4092 = ~n3545 & ~n4091;
  assign n4093 = ~controllable_hgrant2 & ~n4092;
  assign n4094 = ~n3410 & ~n4093;
  assign n4095 = controllable_hmaster1 & ~n4094;
  assign n4096 = controllable_hmaster0 & ~n4094;
  assign n4097 = ~n3545 & ~n4015;
  assign n4098 = ~controllable_hgrant2 & ~n4097;
  assign n4099 = ~n3410 & ~n4098;
  assign n4100 = ~controllable_hmaster0 & ~n4099;
  assign n4101 = ~n4096 & ~n4100;
  assign n4102 = ~controllable_hmaster1 & ~n4101;
  assign n4103 = ~n4095 & ~n4102;
  assign n4104 = i_hbusreq3 & ~n4103;
  assign n4105 = i_hbusreq2 & ~n4092;
  assign n4106 = i_hbusreq4 & ~n4090;
  assign n4107 = i_hbusreq0 & ~n4090;
  assign n4108 = ~n3392 & ~n4031;
  assign n4109 = i_hlock0 & ~n4108;
  assign n4110 = ~n3392 & ~n4000;
  assign n4111 = ~i_hlock0 & ~n4110;
  assign n4112 = ~n4109 & ~n4111;
  assign n4113 = ~i_hbusreq0 & ~n4112;
  assign n4114 = ~n4107 & ~n4113;
  assign n4115 = ~i_hbusreq4 & ~n4114;
  assign n4116 = ~n4106 & ~n4115;
  assign n4117 = controllable_hgrant4 & ~n4116;
  assign n4118 = ~n3574 & ~n4117;
  assign n4119 = ~i_hbusreq2 & ~n4118;
  assign n4120 = ~n4105 & ~n4119;
  assign n4121 = ~controllable_hgrant2 & ~n4120;
  assign n4122 = ~n3431 & ~n4121;
  assign n4123 = controllable_hmaster1 & ~n4122;
  assign n4124 = controllable_hmaster0 & ~n4122;
  assign n4125 = i_hbusreq2 & ~n4097;
  assign n4126 = i_hlock0 & ~n3569;
  assign n4127 = ~n3495 & ~n3568;
  assign n4128 = ~i_hlock0 & ~n4127;
  assign n4129 = ~n4126 & ~n4128;
  assign n4130 = ~i_hbusreq0 & ~n4129;
  assign n4131 = ~n3563 & ~n4130;
  assign n4132 = ~i_hbusreq4 & ~n4131;
  assign n4133 = ~n3562 & ~n4132;
  assign n4134 = ~controllable_hgrant4 & ~n4133;
  assign n4135 = ~n4064 & ~n4134;
  assign n4136 = ~i_hbusreq2 & ~n4135;
  assign n4137 = ~n4125 & ~n4136;
  assign n4138 = ~controllable_hgrant2 & ~n4137;
  assign n4139 = ~n3859 & ~n4138;
  assign n4140 = ~controllable_hmaster0 & ~n4139;
  assign n4141 = ~n4124 & ~n4140;
  assign n4142 = ~controllable_hmaster1 & ~n4141;
  assign n4143 = ~n4123 & ~n4142;
  assign n4144 = ~i_hbusreq3 & ~n4143;
  assign n4145 = ~n4104 & ~n4144;
  assign n4146 = controllable_hmaster2 & ~n4145;
  assign n4147 = ~n3552 & ~n4002;
  assign n4148 = ~controllable_hgrant2 & ~n4147;
  assign n4149 = ~controllable_hgrant2 & ~n4148;
  assign n4150 = i_hbusreq3 & ~n4149;
  assign n4151 = i_hbusreq2 & ~n4147;
  assign n4152 = ~n3590 & ~n4040;
  assign n4153 = ~i_hbusreq2 & ~n4152;
  assign n4154 = ~n4151 & ~n4153;
  assign n4155 = ~controllable_hgrant2 & ~n4154;
  assign n4156 = ~controllable_hgrant2 & ~n4155;
  assign n4157 = ~i_hbusreq3 & ~n4156;
  assign n4158 = ~n4150 & ~n4157;
  assign n4159 = ~controllable_hmaster2 & ~n4158;
  assign n4160 = ~n4146 & ~n4159;
  assign n4161 = ~controllable_hgrant3 & ~n4160;
  assign n4162 = ~n3959 & ~n4161;
  assign n4163 = controllable_nhgrant0 & ~n4162;
  assign n4164 = ~n3987 & ~n4163;
  assign n4165 = ~n3281 & ~n4164;
  assign n4166 = ~n4089 & ~n4165;
  assign n4167 = ~n3378 & ~n4166;
  assign n4168 = ~n4088 & ~n4167;
  assign n4169 = n3492 & ~n4168;
  assign n4170 = ~n3493 & ~n4169;
  assign n4171 = n3485 & ~n4170;
  assign n4172 = ~n3486 & ~n4171;
  assign n4173 = n3476 & ~n4172;
  assign n4174 = ~n3997 & ~n4173;
  assign n4175 = n3374 & ~n4174;
  assign n4176 = ~n3820 & ~n4175;
  assign n4177 = n3655 & ~n4176;
  assign n4178 = controllable_hgrant1 & controllable_locked;
  assign n4179 = controllable_ndecide & n4178;
  assign n4180 = ~i_hready & n4179;
  assign n4181 = ~i_hready & ~n4180;
  assign n4182 = ~controllable_hgrant4 & ~n4181;
  assign n4183 = ~n3848 & ~n4182;
  assign n4184 = ~controllable_hgrant2 & ~n4183;
  assign n4185 = ~n3410 & ~n4184;
  assign n4186 = ~controllable_hmaster0 & ~n4185;
  assign n4187 = ~controllable_hmaster0 & ~n4186;
  assign n4188 = ~controllable_hmaster1 & ~n4187;
  assign n4189 = ~controllable_hmaster1 & ~n4188;
  assign n4190 = i_hbusreq3 & ~n4189;
  assign n4191 = i_hbusreq2 & ~n4183;
  assign n4192 = i_hbusreq4 & ~n4181;
  assign n4193 = i_hbusreq0 & ~n4181;
  assign n4194 = ~n3390 & ~n4179;
  assign n4195 = ~i_hready & ~n4194;
  assign n4196 = ~i_hready & ~n4195;
  assign n4197 = i_hlock0 & ~n4196;
  assign n4198 = ~i_hlock0 & ~n4181;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = ~i_hbusreq0 & ~n4199;
  assign n4201 = ~n4193 & ~n4200;
  assign n4202 = ~i_hbusreq4 & ~n4201;
  assign n4203 = ~n4192 & ~n4202;
  assign n4204 = ~controllable_hgrant4 & ~n4203;
  assign n4205 = ~n3873 & ~n4204;
  assign n4206 = ~i_hbusreq2 & ~n4205;
  assign n4207 = ~n4191 & ~n4206;
  assign n4208 = ~controllable_hgrant2 & ~n4207;
  assign n4209 = ~n3859 & ~n4208;
  assign n4210 = ~controllable_hmaster0 & ~n4209;
  assign n4211 = ~controllable_hmaster0 & ~n4210;
  assign n4212 = ~controllable_hmaster1 & ~n4211;
  assign n4213 = ~controllable_hmaster1 & ~n4212;
  assign n4214 = ~i_hbusreq3 & ~n4213;
  assign n4215 = ~n4190 & ~n4214;
  assign n4216 = controllable_hmaster2 & ~n4215;
  assign n4217 = controllable_hmaster2 & ~n4216;
  assign n4218 = ~controllable_hgrant3 & ~n4217;
  assign n4219 = ~n3843 & ~n4218;
  assign n4220 = controllable_nhgrant0 & ~n4219;
  assign n4221 = ~n3945 & ~n4220;
  assign n4222 = ~n3281 & ~n4221;
  assign n4223 = ~n3281 & ~n4222;
  assign n4224 = n3378 & ~n4223;
  assign n4225 = ~n3502 & ~n4186;
  assign n4226 = ~controllable_hmaster1 & ~n4225;
  assign n4227 = ~n3501 & ~n4226;
  assign n4228 = i_hbusreq3 & ~n4227;
  assign n4229 = ~n3524 & ~n4210;
  assign n4230 = ~controllable_hmaster1 & ~n4229;
  assign n4231 = ~n3523 & ~n4230;
  assign n4232 = ~i_hbusreq3 & ~n4231;
  assign n4233 = ~n4228 & ~n4232;
  assign n4234 = controllable_hmaster2 & ~n4233;
  assign n4235 = controllable_hmaster2 & ~n4234;
  assign n4236 = ~controllable_hgrant3 & ~n4235;
  assign n4237 = ~n3959 & ~n4236;
  assign n4238 = controllable_nhgrant0 & ~n4237;
  assign n4239 = ~n3987 & ~n4238;
  assign n4240 = ~n3281 & ~n4239;
  assign n4241 = ~n3950 & ~n4240;
  assign n4242 = ~n3378 & ~n4241;
  assign n4243 = ~n4224 & ~n4242;
  assign n4244 = n3492 & ~n4243;
  assign n4245 = ~n3493 & ~n4244;
  assign n4246 = n3485 & ~n4245;
  assign n4247 = ~n3486 & ~n4246;
  assign n4248 = ~n3476 & ~n4247;
  assign n4249 = ~n4015 & ~n4182;
  assign n4250 = ~controllable_hgrant2 & ~n4249;
  assign n4251 = ~n3410 & ~n4250;
  assign n4252 = ~controllable_hmaster0 & ~n4251;
  assign n4253 = ~n4007 & ~n4252;
  assign n4254 = ~controllable_hmaster1 & ~n4253;
  assign n4255 = ~n4006 & ~n4254;
  assign n4256 = i_hbusreq3 & ~n4255;
  assign n4257 = i_hbusreq2 & ~n4249;
  assign n4258 = ~n4064 & ~n4204;
  assign n4259 = ~i_hbusreq2 & ~n4258;
  assign n4260 = ~n4257 & ~n4259;
  assign n4261 = ~controllable_hgrant2 & ~n4260;
  assign n4262 = ~n3859 & ~n4261;
  assign n4263 = ~controllable_hmaster0 & ~n4262;
  assign n4264 = ~n4047 & ~n4263;
  assign n4265 = ~controllable_hmaster1 & ~n4264;
  assign n4266 = ~n4046 & ~n4265;
  assign n4267 = ~i_hbusreq3 & ~n4266;
  assign n4268 = ~n4256 & ~n4267;
  assign n4269 = controllable_hmaster2 & ~n4268;
  assign n4270 = ~n4080 & ~n4269;
  assign n4271 = ~controllable_hgrant3 & ~n4270;
  assign n4272 = ~n3843 & ~n4271;
  assign n4273 = controllable_nhgrant0 & ~n4272;
  assign n4274 = ~n3945 & ~n4273;
  assign n4275 = ~n3281 & ~n4274;
  assign n4276 = ~n3281 & ~n4275;
  assign n4277 = n3378 & ~n4276;
  assign n4278 = ~n3543 & ~n4180;
  assign n4279 = ~controllable_hgrant4 & ~n4278;
  assign n4280 = ~n4015 & ~n4279;
  assign n4281 = ~controllable_hgrant2 & ~n4280;
  assign n4282 = ~n3410 & ~n4281;
  assign n4283 = ~controllable_hmaster0 & ~n4282;
  assign n4284 = ~n4096 & ~n4283;
  assign n4285 = ~controllable_hmaster1 & ~n4284;
  assign n4286 = ~n4095 & ~n4285;
  assign n4287 = i_hbusreq3 & ~n4286;
  assign n4288 = i_hbusreq2 & ~n4280;
  assign n4289 = i_hbusreq4 & ~n4278;
  assign n4290 = i_hbusreq0 & ~n4278;
  assign n4291 = ~n3568 & ~n4195;
  assign n4292 = i_hlock0 & ~n4291;
  assign n4293 = ~n3568 & ~n4180;
  assign n4294 = ~i_hlock0 & ~n4293;
  assign n4295 = ~n4292 & ~n4294;
  assign n4296 = ~i_hbusreq0 & ~n4295;
  assign n4297 = ~n4290 & ~n4296;
  assign n4298 = ~i_hbusreq4 & ~n4297;
  assign n4299 = ~n4289 & ~n4298;
  assign n4300 = ~controllable_hgrant4 & ~n4299;
  assign n4301 = ~n4064 & ~n4300;
  assign n4302 = ~i_hbusreq2 & ~n4301;
  assign n4303 = ~n4288 & ~n4302;
  assign n4304 = ~controllable_hgrant2 & ~n4303;
  assign n4305 = ~n3859 & ~n4304;
  assign n4306 = ~controllable_hmaster0 & ~n4305;
  assign n4307 = ~n4124 & ~n4306;
  assign n4308 = ~controllable_hmaster1 & ~n4307;
  assign n4309 = ~n4123 & ~n4308;
  assign n4310 = ~i_hbusreq3 & ~n4309;
  assign n4311 = ~n4287 & ~n4310;
  assign n4312 = controllable_hmaster2 & ~n4311;
  assign n4313 = ~n4159 & ~n4312;
  assign n4314 = ~controllable_hgrant3 & ~n4313;
  assign n4315 = ~n3959 & ~n4314;
  assign n4316 = controllable_nhgrant0 & ~n4315;
  assign n4317 = ~n3987 & ~n4316;
  assign n4318 = ~n3281 & ~n4317;
  assign n4319 = ~n4089 & ~n4318;
  assign n4320 = ~n3378 & ~n4319;
  assign n4321 = ~n4277 & ~n4320;
  assign n4322 = n3492 & ~n4321;
  assign n4323 = ~n3493 & ~n4322;
  assign n4324 = n3485 & ~n4323;
  assign n4325 = ~n3486 & ~n4324;
  assign n4326 = n3476 & ~n4325;
  assign n4327 = ~n4248 & ~n4326;
  assign n4328 = n3374 & ~n4327;
  assign n4329 = ~n3820 & ~n4328;
  assign n4330 = ~n3655 & ~n4329;
  assign n4331 = ~n4177 & ~n4330;
  assign n4332 = n3652 & ~n4331;
  assign n4333 = controllable_hgrant2 & ~n3907;
  assign n4334 = ~n3852 & ~n4333;
  assign n4335 = ~controllable_hmaster0 & ~n4334;
  assign n4336 = ~controllable_hmaster0 & ~n4335;
  assign n4337 = ~controllable_hmaster1 & ~n4336;
  assign n4338 = ~controllable_hmaster1 & ~n4337;
  assign n4339 = i_hbusreq3 & ~n4338;
  assign n4340 = controllable_hgrant2 & ~n3932;
  assign n4341 = ~n3888 & ~n4340;
  assign n4342 = ~controllable_hmaster0 & ~n4341;
  assign n4343 = ~controllable_hmaster0 & ~n4342;
  assign n4344 = ~controllable_hmaster1 & ~n4343;
  assign n4345 = ~controllable_hmaster1 & ~n4344;
  assign n4346 = ~i_hbusreq3 & ~n4345;
  assign n4347 = ~n4339 & ~n4346;
  assign n4348 = controllable_hmaster2 & ~n4347;
  assign n4349 = controllable_hmaster2 & ~n4348;
  assign n4350 = ~controllable_hgrant3 & ~n4349;
  assign n4351 = ~n3843 & ~n4350;
  assign n4352 = controllable_nhgrant0 & ~n4351;
  assign n4353 = ~n3945 & ~n4352;
  assign n4354 = ~n3281 & ~n4353;
  assign n4355 = ~n3281 & ~n4354;
  assign n4356 = n3378 & ~n4355;
  assign n4357 = ~n3502 & ~n4335;
  assign n4358 = ~controllable_hmaster1 & ~n4357;
  assign n4359 = ~n3501 & ~n4358;
  assign n4360 = i_hbusreq3 & ~n4359;
  assign n4361 = ~n3524 & ~n4342;
  assign n4362 = ~controllable_hmaster1 & ~n4361;
  assign n4363 = ~n3523 & ~n4362;
  assign n4364 = ~i_hbusreq3 & ~n4363;
  assign n4365 = ~n4360 & ~n4364;
  assign n4366 = controllable_hmaster2 & ~n4365;
  assign n4367 = controllable_hmaster2 & ~n4366;
  assign n4368 = ~controllable_hgrant3 & ~n4367;
  assign n4369 = ~n3959 & ~n4368;
  assign n4370 = controllable_nhgrant0 & ~n4369;
  assign n4371 = ~n3987 & ~n4370;
  assign n4372 = ~n3281 & ~n4371;
  assign n4373 = ~n3950 & ~n4372;
  assign n4374 = ~n3378 & ~n4373;
  assign n4375 = ~n4356 & ~n4374;
  assign n4376 = n3492 & ~n4375;
  assign n4377 = ~n3493 & ~n4376;
  assign n4378 = n3485 & ~n4377;
  assign n4379 = ~n3486 & ~n4378;
  assign n4380 = ~n3476 & ~n4379;
  assign n4381 = ~n4017 & ~n4333;
  assign n4382 = ~controllable_hmaster0 & ~n4381;
  assign n4383 = ~n4007 & ~n4382;
  assign n4384 = ~controllable_hmaster1 & ~n4383;
  assign n4385 = ~n4006 & ~n4384;
  assign n4386 = i_hbusreq3 & ~n4385;
  assign n4387 = ~n4068 & ~n4340;
  assign n4388 = ~controllable_hmaster0 & ~n4387;
  assign n4389 = ~n4047 & ~n4388;
  assign n4390 = ~controllable_hmaster1 & ~n4389;
  assign n4391 = ~n4046 & ~n4390;
  assign n4392 = ~i_hbusreq3 & ~n4391;
  assign n4393 = ~n4386 & ~n4392;
  assign n4394 = controllable_hmaster2 & ~n4393;
  assign n4395 = ~n4080 & ~n4394;
  assign n4396 = ~controllable_hgrant3 & ~n4395;
  assign n4397 = ~n3843 & ~n4396;
  assign n4398 = controllable_nhgrant0 & ~n4397;
  assign n4399 = ~n3945 & ~n4398;
  assign n4400 = ~n3281 & ~n4399;
  assign n4401 = ~n3281 & ~n4400;
  assign n4402 = n3378 & ~n4401;
  assign n4403 = ~n4098 & ~n4333;
  assign n4404 = ~controllable_hmaster0 & ~n4403;
  assign n4405 = ~n4096 & ~n4404;
  assign n4406 = ~controllable_hmaster1 & ~n4405;
  assign n4407 = ~n4095 & ~n4406;
  assign n4408 = i_hbusreq3 & ~n4407;
  assign n4409 = ~n4138 & ~n4340;
  assign n4410 = ~controllable_hmaster0 & ~n4409;
  assign n4411 = ~n4124 & ~n4410;
  assign n4412 = ~controllable_hmaster1 & ~n4411;
  assign n4413 = ~n4123 & ~n4412;
  assign n4414 = ~i_hbusreq3 & ~n4413;
  assign n4415 = ~n4408 & ~n4414;
  assign n4416 = controllable_hmaster2 & ~n4415;
  assign n4417 = ~n4159 & ~n4416;
  assign n4418 = ~controllable_hgrant3 & ~n4417;
  assign n4419 = ~n3959 & ~n4418;
  assign n4420 = controllable_nhgrant0 & ~n4419;
  assign n4421 = ~n3987 & ~n4420;
  assign n4422 = ~n3281 & ~n4421;
  assign n4423 = ~n4089 & ~n4422;
  assign n4424 = ~n3378 & ~n4423;
  assign n4425 = ~n4402 & ~n4424;
  assign n4426 = n3492 & ~n4425;
  assign n4427 = ~n3493 & ~n4426;
  assign n4428 = n3485 & ~n4427;
  assign n4429 = ~n3486 & ~n4428;
  assign n4430 = n3476 & ~n4429;
  assign n4431 = ~n4380 & ~n4430;
  assign n4432 = n3374 & ~n4431;
  assign n4433 = ~n3820 & ~n4432;
  assign n4434 = n3655 & ~n4433;
  assign n4435 = ~n4184 & ~n4333;
  assign n4436 = ~controllable_hmaster0 & ~n4435;
  assign n4437 = ~controllable_hmaster0 & ~n4436;
  assign n4438 = ~controllable_hmaster1 & ~n4437;
  assign n4439 = ~controllable_hmaster1 & ~n4438;
  assign n4440 = i_hbusreq3 & ~n4439;
  assign n4441 = ~n4208 & ~n4340;
  assign n4442 = ~controllable_hmaster0 & ~n4441;
  assign n4443 = ~controllable_hmaster0 & ~n4442;
  assign n4444 = ~controllable_hmaster1 & ~n4443;
  assign n4445 = ~controllable_hmaster1 & ~n4444;
  assign n4446 = ~i_hbusreq3 & ~n4445;
  assign n4447 = ~n4440 & ~n4446;
  assign n4448 = controllable_hmaster2 & ~n4447;
  assign n4449 = controllable_hmaster2 & ~n4448;
  assign n4450 = ~controllable_hgrant3 & ~n4449;
  assign n4451 = ~n3843 & ~n4450;
  assign n4452 = controllable_nhgrant0 & ~n4451;
  assign n4453 = ~n3945 & ~n4452;
  assign n4454 = ~n3281 & ~n4453;
  assign n4455 = ~n3281 & ~n4454;
  assign n4456 = n3378 & ~n4455;
  assign n4457 = ~n3502 & ~n4436;
  assign n4458 = ~controllable_hmaster1 & ~n4457;
  assign n4459 = ~n3501 & ~n4458;
  assign n4460 = i_hbusreq3 & ~n4459;
  assign n4461 = ~n3524 & ~n4442;
  assign n4462 = ~controllable_hmaster1 & ~n4461;
  assign n4463 = ~n3523 & ~n4462;
  assign n4464 = ~i_hbusreq3 & ~n4463;
  assign n4465 = ~n4460 & ~n4464;
  assign n4466 = controllable_hmaster2 & ~n4465;
  assign n4467 = controllable_hmaster2 & ~n4466;
  assign n4468 = ~controllable_hgrant3 & ~n4467;
  assign n4469 = ~n3959 & ~n4468;
  assign n4470 = controllable_nhgrant0 & ~n4469;
  assign n4471 = ~n3987 & ~n4470;
  assign n4472 = ~n3281 & ~n4471;
  assign n4473 = ~n3950 & ~n4472;
  assign n4474 = ~n3378 & ~n4473;
  assign n4475 = ~n4456 & ~n4474;
  assign n4476 = n3492 & ~n4475;
  assign n4477 = ~n3493 & ~n4476;
  assign n4478 = n3485 & ~n4477;
  assign n4479 = ~n3486 & ~n4478;
  assign n4480 = ~n3476 & ~n4479;
  assign n4481 = ~n4250 & ~n4333;
  assign n4482 = ~controllable_hmaster0 & ~n4481;
  assign n4483 = ~n4007 & ~n4482;
  assign n4484 = ~controllable_hmaster1 & ~n4483;
  assign n4485 = ~n4006 & ~n4484;
  assign n4486 = i_hbusreq3 & ~n4485;
  assign n4487 = ~n4261 & ~n4340;
  assign n4488 = ~controllable_hmaster0 & ~n4487;
  assign n4489 = ~n4047 & ~n4488;
  assign n4490 = ~controllable_hmaster1 & ~n4489;
  assign n4491 = ~n4046 & ~n4490;
  assign n4492 = ~i_hbusreq3 & ~n4491;
  assign n4493 = ~n4486 & ~n4492;
  assign n4494 = controllable_hmaster2 & ~n4493;
  assign n4495 = ~n4080 & ~n4494;
  assign n4496 = ~controllable_hgrant3 & ~n4495;
  assign n4497 = ~n3843 & ~n4496;
  assign n4498 = controllable_nhgrant0 & ~n4497;
  assign n4499 = ~n3945 & ~n4498;
  assign n4500 = ~n3281 & ~n4499;
  assign n4501 = ~n3281 & ~n4500;
  assign n4502 = n3378 & ~n4501;
  assign n4503 = ~n4281 & ~n4333;
  assign n4504 = ~controllable_hmaster0 & ~n4503;
  assign n4505 = ~n4096 & ~n4504;
  assign n4506 = ~controllable_hmaster1 & ~n4505;
  assign n4507 = ~n4095 & ~n4506;
  assign n4508 = i_hbusreq3 & ~n4507;
  assign n4509 = ~n4304 & ~n4340;
  assign n4510 = ~controllable_hmaster0 & ~n4509;
  assign n4511 = ~n4124 & ~n4510;
  assign n4512 = ~controllable_hmaster1 & ~n4511;
  assign n4513 = ~n4123 & ~n4512;
  assign n4514 = ~i_hbusreq3 & ~n4513;
  assign n4515 = ~n4508 & ~n4514;
  assign n4516 = controllable_hmaster2 & ~n4515;
  assign n4517 = ~n4159 & ~n4516;
  assign n4518 = ~controllable_hgrant3 & ~n4517;
  assign n4519 = ~n3959 & ~n4518;
  assign n4520 = controllable_nhgrant0 & ~n4519;
  assign n4521 = ~n3987 & ~n4520;
  assign n4522 = ~n3281 & ~n4521;
  assign n4523 = ~n4089 & ~n4522;
  assign n4524 = ~n3378 & ~n4523;
  assign n4525 = ~n4502 & ~n4524;
  assign n4526 = n3492 & ~n4525;
  assign n4527 = ~n3493 & ~n4526;
  assign n4528 = n3485 & ~n4527;
  assign n4529 = ~n3486 & ~n4528;
  assign n4530 = n3476 & ~n4529;
  assign n4531 = ~n4480 & ~n4530;
  assign n4532 = n3374 & ~n4531;
  assign n4533 = ~n3820 & ~n4532;
  assign n4534 = ~n3655 & ~n4533;
  assign n4535 = ~n4434 & ~n4534;
  assign n4536 = ~n3652 & ~n4535;
  assign n4537 = ~n4332 & ~n4536;
  assign n4538 = ~n3368 & ~n4537;
  assign n4539 = ~i_hbusreq1 & ~controllable_hmastlock;
  assign n4540 = ~i_hbusreq1 & ~n4539;
  assign n4541 = ~controllable_ndecide & n4540;
  assign n4542 = ~controllable_ndecide & ~n4541;
  assign n4543 = ~i_hready & ~n4542;
  assign n4544 = ~i_hready & ~n4543;
  assign n4545 = i_hlock0 & ~n4544;
  assign n4546 = ~n3827 & ~n4545;
  assign n4547 = ~i_hbusreq0 & ~n4546;
  assign n4548 = ~n3389 & ~n4547;
  assign n4549 = ~i_hbusreq4 & ~n4548;
  assign n4550 = ~n3388 & ~n4549;
  assign n4551 = ~i_hbusreq2 & ~n4550;
  assign n4552 = ~n3387 & ~n4551;
  assign n4553 = ~controllable_hmaster0 & ~n4552;
  assign n4554 = ~controllable_hmaster0 & ~n4553;
  assign n4555 = ~controllable_hmaster1 & ~n4554;
  assign n4556 = ~controllable_hmaster1 & ~n4555;
  assign n4557 = ~i_hbusreq3 & ~n4556;
  assign n4558 = ~n3825 & ~n4557;
  assign n4559 = controllable_hmaster2 & ~n4558;
  assign n4560 = controllable_hmaster2 & ~n4559;
  assign n4561 = controllable_hgrant3 & ~n4560;
  assign n4562 = controllable_hgrant2 & ~n4552;
  assign n4563 = ~i_hbusreq1 & ~n3717;
  assign n4564 = ~n3436 & ~n4563;
  assign n4565 = ~controllable_ndecide & ~n4564;
  assign n4566 = ~controllable_ndecide & ~n4565;
  assign n4567 = i_hready & ~n4566;
  assign n4568 = ~n4543 & ~n4567;
  assign n4569 = i_hlock0 & ~n4568;
  assign n4570 = ~n3867 & ~n4569;
  assign n4571 = ~i_hbusreq0 & ~n4570;
  assign n4572 = ~n3862 & ~n4571;
  assign n4573 = ~i_hbusreq4 & ~n4572;
  assign n4574 = ~n3861 & ~n4573;
  assign n4575 = controllable_hgrant4 & ~n4574;
  assign n4576 = ~n3494 & ~n4541;
  assign n4577 = ~i_hready & ~n4576;
  assign n4578 = ~i_hready & ~n4577;
  assign n4579 = i_hlock0 & ~n4578;
  assign n4580 = ~n3878 & ~n4579;
  assign n4581 = ~i_hbusreq0 & ~n4580;
  assign n4582 = ~n3875 & ~n4581;
  assign n4583 = ~i_hbusreq4 & ~n4582;
  assign n4584 = ~n3874 & ~n4583;
  assign n4585 = ~controllable_hgrant4 & ~n4584;
  assign n4586 = ~n4575 & ~n4585;
  assign n4587 = ~i_hbusreq2 & ~n4586;
  assign n4588 = ~n3860 & ~n4587;
  assign n4589 = ~controllable_hgrant2 & ~n4588;
  assign n4590 = ~n4562 & ~n4589;
  assign n4591 = ~controllable_hmaster0 & ~n4590;
  assign n4592 = ~controllable_hmaster0 & ~n4591;
  assign n4593 = ~controllable_hmaster1 & ~n4592;
  assign n4594 = ~controllable_hmaster1 & ~n4593;
  assign n4595 = ~i_hbusreq3 & ~n4594;
  assign n4596 = ~n3858 & ~n4595;
  assign n4597 = controllable_hmaster2 & ~n4596;
  assign n4598 = controllable_hmaster2 & ~n4597;
  assign n4599 = ~controllable_hgrant3 & ~n4598;
  assign n4600 = ~n4561 & ~n4599;
  assign n4601 = controllable_nhgrant0 & ~n4600;
  assign n4602 = ~controllable_hgrant1 & n3412;
  assign n4603 = ~controllable_hgrant1 & ~n4602;
  assign n4604 = controllable_ndecide & ~n4603;
  assign n4605 = ~i_hready & n4604;
  assign n4606 = ~i_hready & ~n4605;
  assign n4607 = ~controllable_hgrant4 & ~n4606;
  assign n4608 = ~n3411 & ~n4607;
  assign n4609 = ~controllable_hgrant2 & ~n4608;
  assign n4610 = ~n3410 & ~n4609;
  assign n4611 = ~controllable_hmaster0 & ~n4610;
  assign n4612 = ~controllable_hmaster0 & ~n4611;
  assign n4613 = ~controllable_hmaster1 & ~n4612;
  assign n4614 = ~controllable_hmaster1 & ~n4613;
  assign n4615 = i_hbusreq3 & ~n4614;
  assign n4616 = i_hbusreq2 & ~n4608;
  assign n4617 = controllable_hgrant4 & ~n4550;
  assign n4618 = i_hbusreq4 & ~n4606;
  assign n4619 = i_hbusreq0 & ~n4606;
  assign n4620 = ~n4541 & ~n4604;
  assign n4621 = ~i_hready & ~n4620;
  assign n4622 = ~i_hready & ~n4621;
  assign n4623 = i_hlock0 & ~n4622;
  assign n4624 = ~i_hlock0 & ~n4606;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~i_hbusreq0 & ~n4625;
  assign n4627 = ~n4619 & ~n4626;
  assign n4628 = ~i_hbusreq4 & ~n4627;
  assign n4629 = ~n4618 & ~n4628;
  assign n4630 = ~controllable_hgrant4 & ~n4629;
  assign n4631 = ~n4617 & ~n4630;
  assign n4632 = ~i_hbusreq2 & ~n4631;
  assign n4633 = ~n4616 & ~n4632;
  assign n4634 = ~controllable_hgrant2 & ~n4633;
  assign n4635 = ~n4562 & ~n4634;
  assign n4636 = ~controllable_hmaster0 & ~n4635;
  assign n4637 = ~controllable_hmaster0 & ~n4636;
  assign n4638 = ~controllable_hmaster1 & ~n4637;
  assign n4639 = ~controllable_hmaster1 & ~n4638;
  assign n4640 = ~i_hbusreq3 & ~n4639;
  assign n4641 = ~n4615 & ~n4640;
  assign n4642 = controllable_hmaster2 & ~n4641;
  assign n4643 = controllable_hmaster2 & ~n4642;
  assign n4644 = ~controllable_hgrant3 & ~n4643;
  assign n4645 = ~n4561 & ~n4644;
  assign n4646 = ~controllable_nhgrant0 & ~n4645;
  assign n4647 = ~n4601 & ~n4646;
  assign n4648 = ~n3281 & ~n4647;
  assign n4649 = ~n3281 & ~n4648;
  assign n4650 = n3492 & ~n4649;
  assign n4651 = n3492 & ~n4650;
  assign n4652 = n3485 & ~n4651;
  assign n4653 = n3485 & ~n4652;
  assign n4654 = ~n3476 & ~n4653;
  assign n4655 = ~i_hbusreq1 & ~n3902;
  assign n4656 = ~n4051 & ~n4655;
  assign n4657 = ~controllable_ndecide & ~n4656;
  assign n4658 = ~controllable_ndecide & ~n4657;
  assign n4659 = i_hready & ~n4658;
  assign n4660 = ~n4543 & ~n4659;
  assign n4661 = i_hlock0 & ~n4660;
  assign n4662 = ~n4058 & ~n4661;
  assign n4663 = ~i_hbusreq0 & ~n4662;
  assign n4664 = ~n4050 & ~n4663;
  assign n4665 = ~i_hbusreq4 & ~n4664;
  assign n4666 = ~n4049 & ~n4665;
  assign n4667 = controllable_hgrant4 & ~n4666;
  assign n4668 = ~n4585 & ~n4667;
  assign n4669 = ~i_hbusreq2 & ~n4668;
  assign n4670 = ~n4048 & ~n4669;
  assign n4671 = ~controllable_hgrant2 & ~n4670;
  assign n4672 = ~n4562 & ~n4671;
  assign n4673 = ~controllable_hmaster0 & ~n4672;
  assign n4674 = ~n4007 & ~n4673;
  assign n4675 = ~controllable_hmaster1 & ~n4674;
  assign n4676 = ~n4006 & ~n4675;
  assign n4677 = ~i_hbusreq3 & ~n4676;
  assign n4678 = ~n4023 & ~n4677;
  assign n4679 = controllable_hmaster2 & ~n4678;
  assign n4680 = ~controllable_hmaster2 & ~n4005;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = ~controllable_hgrant3 & ~n4681;
  assign n4683 = ~n4561 & ~n4682;
  assign n4684 = controllable_nhgrant0 & ~n4683;
  assign n4685 = ~n4646 & ~n4684;
  assign n4686 = ~n3281 & ~n4685;
  assign n4687 = ~n3281 & ~n4686;
  assign n4688 = n3492 & ~n4687;
  assign n4689 = n3492 & ~n4688;
  assign n4690 = n3485 & ~n4689;
  assign n4691 = n3485 & ~n4690;
  assign n4692 = n3476 & ~n4691;
  assign n4693 = ~n4654 & ~n4692;
  assign n4694 = n3374 & ~n4693;
  assign n4695 = n3374 & ~n4694;
  assign n4696 = n3655 & ~n4695;
  assign n4697 = controllable_hgrant1 & n3412;
  assign n4698 = controllable_ndecide & n4697;
  assign n4699 = ~i_hready & n4698;
  assign n4700 = ~i_hready & ~n4699;
  assign n4701 = ~controllable_hgrant4 & ~n4700;
  assign n4702 = ~n3848 & ~n4701;
  assign n4703 = ~controllable_hgrant2 & ~n4702;
  assign n4704 = ~n3410 & ~n4703;
  assign n4705 = ~controllable_hmaster0 & ~n4704;
  assign n4706 = ~controllable_hmaster0 & ~n4705;
  assign n4707 = ~controllable_hmaster1 & ~n4706;
  assign n4708 = ~controllable_hmaster1 & ~n4707;
  assign n4709 = i_hbusreq3 & ~n4708;
  assign n4710 = i_hbusreq2 & ~n4702;
  assign n4711 = i_hbusreq4 & ~n4700;
  assign n4712 = i_hbusreq0 & ~n4700;
  assign n4713 = ~n4541 & ~n4698;
  assign n4714 = ~i_hready & ~n4713;
  assign n4715 = ~i_hready & ~n4714;
  assign n4716 = i_hlock0 & ~n4715;
  assign n4717 = ~i_hlock0 & ~n4700;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~i_hbusreq0 & ~n4718;
  assign n4720 = ~n4712 & ~n4719;
  assign n4721 = ~i_hbusreq4 & ~n4720;
  assign n4722 = ~n4711 & ~n4721;
  assign n4723 = ~controllable_hgrant4 & ~n4722;
  assign n4724 = ~n4575 & ~n4723;
  assign n4725 = ~i_hbusreq2 & ~n4724;
  assign n4726 = ~n4710 & ~n4725;
  assign n4727 = ~controllable_hgrant2 & ~n4726;
  assign n4728 = ~n4562 & ~n4727;
  assign n4729 = ~controllable_hmaster0 & ~n4728;
  assign n4730 = ~controllable_hmaster0 & ~n4729;
  assign n4731 = ~controllable_hmaster1 & ~n4730;
  assign n4732 = ~controllable_hmaster1 & ~n4731;
  assign n4733 = ~i_hbusreq3 & ~n4732;
  assign n4734 = ~n4709 & ~n4733;
  assign n4735 = controllable_hmaster2 & ~n4734;
  assign n4736 = controllable_hmaster2 & ~n4735;
  assign n4737 = ~controllable_hgrant3 & ~n4736;
  assign n4738 = ~n4561 & ~n4737;
  assign n4739 = controllable_nhgrant0 & ~n4738;
  assign n4740 = ~n4646 & ~n4739;
  assign n4741 = ~n3281 & ~n4740;
  assign n4742 = ~n3281 & ~n4741;
  assign n4743 = n3492 & ~n4742;
  assign n4744 = n3492 & ~n4743;
  assign n4745 = n3485 & ~n4744;
  assign n4746 = n3485 & ~n4745;
  assign n4747 = ~n3476 & ~n4746;
  assign n4748 = ~n4015 & ~n4701;
  assign n4749 = ~controllable_hgrant2 & ~n4748;
  assign n4750 = ~n3410 & ~n4749;
  assign n4751 = ~controllable_hmaster0 & ~n4750;
  assign n4752 = ~n4007 & ~n4751;
  assign n4753 = ~controllable_hmaster1 & ~n4752;
  assign n4754 = ~n4006 & ~n4753;
  assign n4755 = i_hbusreq3 & ~n4754;
  assign n4756 = i_hbusreq2 & ~n4748;
  assign n4757 = ~n4667 & ~n4723;
  assign n4758 = ~i_hbusreq2 & ~n4757;
  assign n4759 = ~n4756 & ~n4758;
  assign n4760 = ~controllable_hgrant2 & ~n4759;
  assign n4761 = ~n4562 & ~n4760;
  assign n4762 = ~controllable_hmaster0 & ~n4761;
  assign n4763 = ~n4007 & ~n4762;
  assign n4764 = ~controllable_hmaster1 & ~n4763;
  assign n4765 = ~n4006 & ~n4764;
  assign n4766 = ~i_hbusreq3 & ~n4765;
  assign n4767 = ~n4755 & ~n4766;
  assign n4768 = controllable_hmaster2 & ~n4767;
  assign n4769 = ~n4680 & ~n4768;
  assign n4770 = ~controllable_hgrant3 & ~n4769;
  assign n4771 = ~n4561 & ~n4770;
  assign n4772 = controllable_nhgrant0 & ~n4771;
  assign n4773 = ~n4646 & ~n4772;
  assign n4774 = ~n3281 & ~n4773;
  assign n4775 = ~n3281 & ~n4774;
  assign n4776 = n3492 & ~n4775;
  assign n4777 = n3492 & ~n4776;
  assign n4778 = n3485 & ~n4777;
  assign n4779 = n3485 & ~n4778;
  assign n4780 = n3476 & ~n4779;
  assign n4781 = ~n4747 & ~n4780;
  assign n4782 = n3374 & ~n4781;
  assign n4783 = n3374 & ~n4782;
  assign n4784 = ~n3655 & ~n4783;
  assign n4785 = ~n4696 & ~n4784;
  assign n4786 = n3652 & ~n4785;
  assign n4787 = controllable_hgrant2 & ~n4608;
  assign n4788 = ~n3852 & ~n4787;
  assign n4789 = ~controllable_hmaster0 & ~n4788;
  assign n4790 = ~controllable_hmaster0 & ~n4789;
  assign n4791 = ~controllable_hmaster1 & ~n4790;
  assign n4792 = ~controllable_hmaster1 & ~n4791;
  assign n4793 = i_hbusreq3 & ~n4792;
  assign n4794 = controllable_hgrant2 & ~n4633;
  assign n4795 = ~n4589 & ~n4794;
  assign n4796 = ~controllable_hmaster0 & ~n4795;
  assign n4797 = ~controllable_hmaster0 & ~n4796;
  assign n4798 = ~controllable_hmaster1 & ~n4797;
  assign n4799 = ~controllable_hmaster1 & ~n4798;
  assign n4800 = ~i_hbusreq3 & ~n4799;
  assign n4801 = ~n4793 & ~n4800;
  assign n4802 = controllable_hmaster2 & ~n4801;
  assign n4803 = controllable_hmaster2 & ~n4802;
  assign n4804 = ~controllable_hgrant3 & ~n4803;
  assign n4805 = ~n4561 & ~n4804;
  assign n4806 = controllable_nhgrant0 & ~n4805;
  assign n4807 = ~n4646 & ~n4806;
  assign n4808 = ~n3281 & ~n4807;
  assign n4809 = ~n3281 & ~n4808;
  assign n4810 = n3492 & ~n4809;
  assign n4811 = n3492 & ~n4810;
  assign n4812 = n3485 & ~n4811;
  assign n4813 = n3485 & ~n4812;
  assign n4814 = ~n3476 & ~n4813;
  assign n4815 = ~n4017 & ~n4787;
  assign n4816 = ~controllable_hmaster0 & ~n4815;
  assign n4817 = ~n4007 & ~n4816;
  assign n4818 = ~controllable_hmaster1 & ~n4817;
  assign n4819 = ~n4006 & ~n4818;
  assign n4820 = i_hbusreq3 & ~n4819;
  assign n4821 = ~n4671 & ~n4794;
  assign n4822 = ~controllable_hmaster0 & ~n4821;
  assign n4823 = ~n4007 & ~n4822;
  assign n4824 = ~controllable_hmaster1 & ~n4823;
  assign n4825 = ~n4006 & ~n4824;
  assign n4826 = ~i_hbusreq3 & ~n4825;
  assign n4827 = ~n4820 & ~n4826;
  assign n4828 = controllable_hmaster2 & ~n4827;
  assign n4829 = ~n4680 & ~n4828;
  assign n4830 = ~controllable_hgrant3 & ~n4829;
  assign n4831 = ~n4561 & ~n4830;
  assign n4832 = controllable_nhgrant0 & ~n4831;
  assign n4833 = ~n4646 & ~n4832;
  assign n4834 = ~n3281 & ~n4833;
  assign n4835 = ~n3281 & ~n4834;
  assign n4836 = n3492 & ~n4835;
  assign n4837 = n3492 & ~n4836;
  assign n4838 = n3485 & ~n4837;
  assign n4839 = n3485 & ~n4838;
  assign n4840 = n3476 & ~n4839;
  assign n4841 = ~n4814 & ~n4840;
  assign n4842 = n3374 & ~n4841;
  assign n4843 = n3374 & ~n4842;
  assign n4844 = n3655 & ~n4843;
  assign n4845 = ~n4703 & ~n4787;
  assign n4846 = ~controllable_hmaster0 & ~n4845;
  assign n4847 = ~controllable_hmaster0 & ~n4846;
  assign n4848 = ~controllable_hmaster1 & ~n4847;
  assign n4849 = ~controllable_hmaster1 & ~n4848;
  assign n4850 = i_hbusreq3 & ~n4849;
  assign n4851 = ~n4727 & ~n4794;
  assign n4852 = ~controllable_hmaster0 & ~n4851;
  assign n4853 = ~controllable_hmaster0 & ~n4852;
  assign n4854 = ~controllable_hmaster1 & ~n4853;
  assign n4855 = ~controllable_hmaster1 & ~n4854;
  assign n4856 = ~i_hbusreq3 & ~n4855;
  assign n4857 = ~n4850 & ~n4856;
  assign n4858 = controllable_hmaster2 & ~n4857;
  assign n4859 = controllable_hmaster2 & ~n4858;
  assign n4860 = ~controllable_hgrant3 & ~n4859;
  assign n4861 = ~n4561 & ~n4860;
  assign n4862 = controllable_nhgrant0 & ~n4861;
  assign n4863 = ~n4646 & ~n4862;
  assign n4864 = ~n3281 & ~n4863;
  assign n4865 = ~n3281 & ~n4864;
  assign n4866 = n3492 & ~n4865;
  assign n4867 = n3492 & ~n4866;
  assign n4868 = n3485 & ~n4867;
  assign n4869 = n3485 & ~n4868;
  assign n4870 = ~n3476 & ~n4869;
  assign n4871 = ~n4749 & ~n4787;
  assign n4872 = ~controllable_hmaster0 & ~n4871;
  assign n4873 = ~n4007 & ~n4872;
  assign n4874 = ~controllable_hmaster1 & ~n4873;
  assign n4875 = ~n4006 & ~n4874;
  assign n4876 = i_hbusreq3 & ~n4875;
  assign n4877 = ~n4760 & ~n4794;
  assign n4878 = ~controllable_hmaster0 & ~n4877;
  assign n4879 = ~n4007 & ~n4878;
  assign n4880 = ~controllable_hmaster1 & ~n4879;
  assign n4881 = ~n4006 & ~n4880;
  assign n4882 = ~i_hbusreq3 & ~n4881;
  assign n4883 = ~n4876 & ~n4882;
  assign n4884 = controllable_hmaster2 & ~n4883;
  assign n4885 = ~n4680 & ~n4884;
  assign n4886 = ~controllable_hgrant3 & ~n4885;
  assign n4887 = ~n4561 & ~n4886;
  assign n4888 = controllable_nhgrant0 & ~n4887;
  assign n4889 = ~n4646 & ~n4888;
  assign n4890 = ~n3281 & ~n4889;
  assign n4891 = ~n3281 & ~n4890;
  assign n4892 = n3492 & ~n4891;
  assign n4893 = n3492 & ~n4892;
  assign n4894 = n3485 & ~n4893;
  assign n4895 = n3485 & ~n4894;
  assign n4896 = n3476 & ~n4895;
  assign n4897 = ~n4870 & ~n4896;
  assign n4898 = n3374 & ~n4897;
  assign n4899 = n3374 & ~n4898;
  assign n4900 = ~n3655 & ~n4899;
  assign n4901 = ~n4844 & ~n4900;
  assign n4902 = ~n3652 & ~n4901;
  assign n4903 = ~n4786 & ~n4902;
  assign n4904 = n3368 & ~n4903;
  assign n4905 = ~n4538 & ~n4904;
  assign n4906 = ~n3362 & ~n4905;
  assign n4907 = ~n3362 & ~n4906;
  assign n4908 = ~n3359 & ~n4907;
  assign n4909 = ~n3359 & ~n4908;
  assign n4910 = n3356 & ~n4909;
  assign n4911 = n3378 & ~n3813;
  assign n4912 = controllable_hmaster1 & ~n3834;
  assign n4913 = controllable_hmaster0 & ~n3834;
  assign n4914 = ~n3697 & ~n4913;
  assign n4915 = ~controllable_hmaster1 & ~n4914;
  assign n4916 = ~n4912 & ~n4915;
  assign n4917 = ~i_hbusreq3 & ~n4916;
  assign n4918 = ~n3787 & ~n4917;
  assign n4919 = controllable_hmaster2 & ~n4918;
  assign n4920 = controllable_hgrant2 & ~n3659;
  assign n4921 = controllable_hgrant4 & ~n3659;
  assign n4922 = ~controllable_hgrant4 & ~n3712;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~controllable_hgrant2 & ~n4923;
  assign n4925 = ~n4920 & ~n4924;
  assign n4926 = controllable_hmaster0 & ~n4925;
  assign n4927 = i_hlock2 & ~n3659;
  assign n4928 = ~i_hlock2 & ~n3664;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~controllable_hmaster0 & ~n4929;
  assign n4931 = ~n4926 & ~n4930;
  assign n4932 = controllable_hmaster1 & ~n4931;
  assign n4933 = i_hlock1 & controllable_hmastlock;
  assign n4934 = ~i_hlock1 & ~controllable_hmastlock;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = ~controllable_ndecide & n4935;
  assign n4937 = ~controllable_ndecide & ~n4936;
  assign n4938 = ~i_hready & ~n4937;
  assign n4939 = ~i_hready & ~n4938;
  assign n4940 = controllable_hmaster0 & ~n4939;
  assign n4941 = i_hlock0 & ~n3659;
  assign n4942 = ~i_hlock0 & ~n3664;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~controllable_hmaster0 & ~n4943;
  assign n4945 = ~n4940 & ~n4944;
  assign n4946 = ~controllable_hmaster1 & ~n4945;
  assign n4947 = ~n4932 & ~n4946;
  assign n4948 = i_hlock3 & ~n4947;
  assign n4949 = controllable_hgrant2 & ~n3664;
  assign n4950 = controllable_hgrant4 & ~n3664;
  assign n4951 = ~controllable_hgrant4 & ~n3721;
  assign n4952 = ~n4950 & ~n4951;
  assign n4953 = ~controllable_hgrant2 & ~n4952;
  assign n4954 = ~n4949 & ~n4953;
  assign n4955 = controllable_hmaster0 & ~n4954;
  assign n4956 = ~n4930 & ~n4955;
  assign n4957 = controllable_hmaster1 & ~n4956;
  assign n4958 = ~n4946 & ~n4957;
  assign n4959 = ~i_hlock3 & ~n4958;
  assign n4960 = ~n4948 & ~n4959;
  assign n4961 = i_hbusreq3 & ~n4960;
  assign n4962 = i_hbusreq2 & ~n3659;
  assign n4963 = i_hbusreq4 & ~n3659;
  assign n4964 = ~i_hbusreq4 & ~n3681;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = ~i_hbusreq2 & ~n4965;
  assign n4967 = ~n4962 & ~n4966;
  assign n4968 = controllable_hgrant2 & ~n4967;
  assign n4969 = i_hbusreq2 & ~n4923;
  assign n4970 = controllable_hgrant4 & ~n4965;
  assign n4971 = i_hbusreq4 & ~n3712;
  assign n4972 = ~i_hbusreq4 & ~n3745;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = ~controllable_hgrant4 & ~n4973;
  assign n4975 = ~n4970 & ~n4974;
  assign n4976 = ~i_hbusreq2 & ~n4975;
  assign n4977 = ~n4969 & ~n4976;
  assign n4978 = ~controllable_hgrant2 & ~n4977;
  assign n4979 = ~n4968 & ~n4978;
  assign n4980 = controllable_hmaster0 & ~n4979;
  assign n4981 = i_hbusreq2 & ~n4929;
  assign n4982 = i_hlock2 & ~n4965;
  assign n4983 = i_hbusreq4 & ~n3664;
  assign n4984 = ~i_hbusreq4 & ~n3690;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = ~i_hlock2 & ~n4985;
  assign n4987 = ~n4982 & ~n4986;
  assign n4988 = ~i_hbusreq2 & ~n4987;
  assign n4989 = ~n4981 & ~n4988;
  assign n4990 = ~controllable_hmaster0 & ~n4989;
  assign n4991 = ~n4980 & ~n4990;
  assign n4992 = controllable_hmaster1 & ~n4991;
  assign n4993 = i_hbusreq2 & ~n4939;
  assign n4994 = i_hbusreq4 & ~n4939;
  assign n4995 = i_hbusreq0 & ~n4939;
  assign n4996 = i_hbusreq1 & ~n4935;
  assign n4997 = ~controllable_ndecide & ~n4996;
  assign n4998 = ~controllable_ndecide & ~n4997;
  assign n4999 = ~i_hready & ~n4998;
  assign n5000 = ~i_hready & ~n4999;
  assign n5001 = ~i_hbusreq0 & ~n5000;
  assign n5002 = ~n4995 & ~n5001;
  assign n5003 = ~i_hbusreq4 & ~n5002;
  assign n5004 = ~n4994 & ~n5003;
  assign n5005 = ~i_hbusreq2 & ~n5004;
  assign n5006 = ~n4993 & ~n5005;
  assign n5007 = controllable_hmaster0 & ~n5006;
  assign n5008 = ~n4944 & ~n5007;
  assign n5009 = ~controllable_hmaster1 & ~n5008;
  assign n5010 = ~n4992 & ~n5009;
  assign n5011 = i_hlock3 & ~n5010;
  assign n5012 = i_hbusreq2 & ~n3664;
  assign n5013 = ~i_hbusreq2 & ~n4985;
  assign n5014 = ~n5012 & ~n5013;
  assign n5015 = controllable_hgrant2 & ~n5014;
  assign n5016 = i_hbusreq2 & ~n4952;
  assign n5017 = controllable_hgrant4 & ~n4985;
  assign n5018 = i_hbusreq4 & ~n3721;
  assign n5019 = ~i_hbusreq4 & ~n3755;
  assign n5020 = ~n5018 & ~n5019;
  assign n5021 = ~controllable_hgrant4 & ~n5020;
  assign n5022 = ~n5017 & ~n5021;
  assign n5023 = ~i_hbusreq2 & ~n5022;
  assign n5024 = ~n5016 & ~n5023;
  assign n5025 = ~controllable_hgrant2 & ~n5024;
  assign n5026 = ~n5015 & ~n5025;
  assign n5027 = controllable_hmaster0 & ~n5026;
  assign n5028 = ~n4990 & ~n5027;
  assign n5029 = controllable_hmaster1 & ~n5028;
  assign n5030 = ~n5009 & ~n5029;
  assign n5031 = ~i_hlock3 & ~n5030;
  assign n5032 = ~n5011 & ~n5031;
  assign n5033 = ~i_hbusreq3 & ~n5032;
  assign n5034 = ~n4961 & ~n5033;
  assign n5035 = ~controllable_hmaster2 & ~n5034;
  assign n5036 = ~n4919 & ~n5035;
  assign n5037 = controllable_hgrant3 & ~n5036;
  assign n5038 = controllable_ndecide & ~n4010;
  assign n5039 = ~i_hready & n5038;
  assign n5040 = ~n3417 & ~n5039;
  assign n5041 = ~controllable_hgrant4 & ~n5040;
  assign n5042 = ~n3411 & ~n5041;
  assign n5043 = ~controllable_hgrant2 & ~n5042;
  assign n5044 = ~n3410 & ~n5043;
  assign n5045 = controllable_hmaster1 & ~n5044;
  assign n5046 = controllable_hmaster0 & ~n5044;
  assign n5047 = ~n3729 & ~n5046;
  assign n5048 = ~controllable_hmaster1 & ~n5047;
  assign n5049 = ~n5045 & ~n5048;
  assign n5050 = i_hbusreq3 & ~n5049;
  assign n5051 = i_hbusreq2 & ~n5042;
  assign n5052 = i_hbusreq4 & ~n5040;
  assign n5053 = i_hbusreq0 & ~n5040;
  assign n5054 = ~n3390 & ~n5038;
  assign n5055 = ~i_hready & ~n5054;
  assign n5056 = ~n3440 & ~n5055;
  assign n5057 = i_hlock0 & ~n5056;
  assign n5058 = ~i_hlock0 & ~n5040;
  assign n5059 = ~n5057 & ~n5058;
  assign n5060 = ~i_hbusreq0 & ~n5059;
  assign n5061 = ~n5053 & ~n5060;
  assign n5062 = ~i_hbusreq4 & ~n5061;
  assign n5063 = ~n5052 & ~n5062;
  assign n5064 = ~controllable_hgrant4 & ~n5063;
  assign n5065 = ~n3916 & ~n5064;
  assign n5066 = ~i_hbusreq2 & ~n5065;
  assign n5067 = ~n5051 & ~n5066;
  assign n5068 = ~controllable_hgrant2 & ~n5067;
  assign n5069 = ~n3859 & ~n5068;
  assign n5070 = controllable_hmaster1 & ~n5069;
  assign n5071 = controllable_hmaster0 & ~n5069;
  assign n5072 = ~n3767 & ~n5071;
  assign n5073 = ~controllable_hmaster1 & ~n5072;
  assign n5074 = ~n5070 & ~n5073;
  assign n5075 = ~i_hbusreq3 & ~n5074;
  assign n5076 = ~n5050 & ~n5075;
  assign n5077 = controllable_hmaster2 & ~n5076;
  assign n5078 = controllable_hmaster0 & ~n3659;
  assign n5079 = i_hlock2 & ~n4923;
  assign n5080 = ~i_hlock2 & ~n4952;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = controllable_hgrant2 & ~n5081;
  assign n5083 = ~controllable_hgrant2 & ~n4929;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = ~controllable_hmaster0 & ~n5084;
  assign n5086 = ~n5078 & ~n5085;
  assign n5087 = controllable_hmaster1 & ~n5086;
  assign n5088 = controllable_hgrant2 & ~n4939;
  assign n5089 = controllable_hgrant4 & ~n4939;
  assign n5090 = i_hlock1 & n4697;
  assign n5091 = controllable_hgrant1 & ~n3715;
  assign n5092 = controllable_hgrant1 & ~n5091;
  assign n5093 = ~i_hlock1 & n5092;
  assign n5094 = ~n5090 & ~n5093;
  assign n5095 = ~controllable_ndecide & n5094;
  assign n5096 = ~controllable_ndecide & ~n5095;
  assign n5097 = i_hready & ~n5096;
  assign n5098 = ~n4938 & ~n5097;
  assign n5099 = ~controllable_hgrant4 & ~n5098;
  assign n5100 = ~n5089 & ~n5099;
  assign n5101 = ~controllable_hgrant2 & ~n5100;
  assign n5102 = ~n5088 & ~n5101;
  assign n5103 = controllable_hmaster0 & ~n5102;
  assign n5104 = ~n4944 & ~n5103;
  assign n5105 = ~controllable_hmaster1 & ~n5104;
  assign n5106 = ~n5087 & ~n5105;
  assign n5107 = i_hlock3 & ~n5106;
  assign n5108 = controllable_hmaster0 & ~n3664;
  assign n5109 = ~n5085 & ~n5108;
  assign n5110 = controllable_hmaster1 & ~n5109;
  assign n5111 = ~n5105 & ~n5110;
  assign n5112 = ~i_hlock3 & ~n5111;
  assign n5113 = ~n5107 & ~n5112;
  assign n5114 = i_hbusreq3 & ~n5113;
  assign n5115 = controllable_hmaster0 & ~n4967;
  assign n5116 = i_hbusreq2 & ~n5081;
  assign n5117 = i_hlock2 & ~n4975;
  assign n5118 = ~i_hlock2 & ~n5022;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = ~i_hbusreq2 & ~n5119;
  assign n5121 = ~n5116 & ~n5120;
  assign n5122 = controllable_hgrant2 & ~n5121;
  assign n5123 = ~controllable_hgrant2 & ~n4989;
  assign n5124 = ~n5122 & ~n5123;
  assign n5125 = ~controllable_hmaster0 & ~n5124;
  assign n5126 = ~n5115 & ~n5125;
  assign n5127 = controllable_hmaster1 & ~n5126;
  assign n5128 = controllable_hgrant2 & ~n5006;
  assign n5129 = i_hbusreq2 & ~n5100;
  assign n5130 = controllable_hgrant4 & ~n5004;
  assign n5131 = i_hbusreq4 & ~n5098;
  assign n5132 = i_hbusreq0 & ~n5098;
  assign n5133 = i_hbusreq1 & ~n5094;
  assign n5134 = ~controllable_ndecide & ~n5133;
  assign n5135 = ~controllable_ndecide & ~n5134;
  assign n5136 = i_hready & ~n5135;
  assign n5137 = ~n4999 & ~n5136;
  assign n5138 = ~i_hbusreq0 & ~n5137;
  assign n5139 = ~n5132 & ~n5138;
  assign n5140 = ~i_hbusreq4 & ~n5139;
  assign n5141 = ~n5131 & ~n5140;
  assign n5142 = ~controllable_hgrant4 & ~n5141;
  assign n5143 = ~n5130 & ~n5142;
  assign n5144 = ~i_hbusreq2 & ~n5143;
  assign n5145 = ~n5129 & ~n5144;
  assign n5146 = ~controllable_hgrant2 & ~n5145;
  assign n5147 = ~n5128 & ~n5146;
  assign n5148 = controllable_hmaster0 & ~n5147;
  assign n5149 = ~n4944 & ~n5148;
  assign n5150 = ~controllable_hmaster1 & ~n5149;
  assign n5151 = ~n5127 & ~n5150;
  assign n5152 = i_hlock3 & ~n5151;
  assign n5153 = controllable_hmaster0 & ~n5014;
  assign n5154 = ~n5125 & ~n5153;
  assign n5155 = controllable_hmaster1 & ~n5154;
  assign n5156 = ~n5150 & ~n5155;
  assign n5157 = ~i_hlock3 & ~n5156;
  assign n5158 = ~n5152 & ~n5157;
  assign n5159 = ~i_hbusreq3 & ~n5158;
  assign n5160 = ~n5114 & ~n5159;
  assign n5161 = ~controllable_hmaster2 & ~n5160;
  assign n5162 = ~n5077 & ~n5161;
  assign n5163 = ~controllable_hgrant3 & ~n5162;
  assign n5164 = ~n5037 & ~n5163;
  assign n5165 = controllable_nhgrant0 & ~n5164;
  assign n5166 = ~n4930 & ~n5078;
  assign n5167 = controllable_hmaster1 & ~n5166;
  assign n5168 = ~n4946 & ~n5167;
  assign n5169 = i_hlock3 & ~n5168;
  assign n5170 = ~n4930 & ~n5108;
  assign n5171 = controllable_hmaster1 & ~n5170;
  assign n5172 = ~n4946 & ~n5171;
  assign n5173 = ~i_hlock3 & ~n5172;
  assign n5174 = ~n5169 & ~n5173;
  assign n5175 = i_hbusreq3 & ~n5174;
  assign n5176 = ~n4990 & ~n5115;
  assign n5177 = controllable_hmaster1 & ~n5176;
  assign n5178 = ~n5009 & ~n5177;
  assign n5179 = i_hlock3 & ~n5178;
  assign n5180 = ~n4990 & ~n5153;
  assign n5181 = controllable_hmaster1 & ~n5180;
  assign n5182 = ~n5009 & ~n5181;
  assign n5183 = ~i_hlock3 & ~n5182;
  assign n5184 = ~n5179 & ~n5183;
  assign n5185 = ~i_hbusreq3 & ~n5184;
  assign n5186 = ~n5175 & ~n5185;
  assign n5187 = ~controllable_hmaster2 & ~n5186;
  assign n5188 = ~n4919 & ~n5187;
  assign n5189 = controllable_hgrant3 & ~n5188;
  assign n5190 = controllable_hmaster1 & ~n3909;
  assign n5191 = controllable_hmaster0 & ~n3909;
  assign n5192 = ~n3667 & ~n5191;
  assign n5193 = ~controllable_hmaster1 & ~n5192;
  assign n5194 = ~n5190 & ~n5193;
  assign n5195 = i_hbusreq3 & ~n5194;
  assign n5196 = controllable_hmaster1 & ~n3934;
  assign n5197 = controllable_hmaster0 & ~n3934;
  assign n5198 = ~n3697 & ~n5197;
  assign n5199 = ~controllable_hmaster1 & ~n5198;
  assign n5200 = ~n5196 & ~n5199;
  assign n5201 = ~i_hbusreq3 & ~n5200;
  assign n5202 = ~n5195 & ~n5201;
  assign n5203 = controllable_hmaster2 & ~n5202;
  assign n5204 = controllable_hgrant2 & ~n4943;
  assign n5205 = controllable_hgrant4 & ~n4943;
  assign n5206 = ~n3418 & ~n3709;
  assign n5207 = i_hready & ~n5206;
  assign n5208 = ~n3418 & ~n3656;
  assign n5209 = ~i_hready & ~n5208;
  assign n5210 = ~n5207 & ~n5209;
  assign n5211 = i_hlock0 & ~n5210;
  assign n5212 = ~n3418 & ~n3718;
  assign n5213 = i_hready & ~n5212;
  assign n5214 = ~n3418 & ~n3661;
  assign n5215 = ~i_hready & ~n5214;
  assign n5216 = ~n5213 & ~n5215;
  assign n5217 = ~i_hlock0 & ~n5216;
  assign n5218 = ~n5211 & ~n5217;
  assign n5219 = ~controllable_hgrant4 & ~n5218;
  assign n5220 = ~n5205 & ~n5219;
  assign n5221 = ~controllable_hgrant2 & ~n5220;
  assign n5222 = ~n5204 & ~n5221;
  assign n5223 = ~controllable_hmaster0 & ~n5222;
  assign n5224 = ~n4940 & ~n5223;
  assign n5225 = ~controllable_hmaster1 & ~n5224;
  assign n5226 = ~n5167 & ~n5225;
  assign n5227 = i_hlock3 & ~n5226;
  assign n5228 = ~n5171 & ~n5225;
  assign n5229 = ~i_hlock3 & ~n5228;
  assign n5230 = ~n5227 & ~n5229;
  assign n5231 = i_hbusreq3 & ~n5230;
  assign n5232 = ~n5007 & ~n5223;
  assign n5233 = ~controllable_hmaster1 & ~n5232;
  assign n5234 = ~n5177 & ~n5233;
  assign n5235 = i_hlock3 & ~n5234;
  assign n5236 = ~n5181 & ~n5233;
  assign n5237 = ~i_hlock3 & ~n5236;
  assign n5238 = ~n5235 & ~n5237;
  assign n5239 = ~i_hbusreq3 & ~n5238;
  assign n5240 = ~n5231 & ~n5239;
  assign n5241 = ~controllable_hmaster2 & ~n5240;
  assign n5242 = ~n5203 & ~n5241;
  assign n5243 = ~controllable_hgrant3 & ~n5242;
  assign n5244 = ~n5189 & ~n5243;
  assign n5245 = ~controllable_nhgrant0 & ~n5244;
  assign n5246 = ~n5165 & ~n5245;
  assign n5247 = ~n3281 & ~n5246;
  assign n5248 = ~n3783 & ~n5247;
  assign n5249 = ~n3378 & ~n5248;
  assign n5250 = ~n4911 & ~n5249;
  assign n5251 = n3492 & ~n5250;
  assign n5252 = ~n3631 & ~n5251;
  assign n5253 = n3485 & ~n5252;
  assign n5254 = ~n3630 & ~n5253;
  assign n5255 = ~n3374 & ~n5254;
  assign n5256 = ~controllable_hgrant4 & ~n3847;
  assign n5257 = ~n3411 & ~n5256;
  assign n5258 = ~controllable_hgrant2 & ~n5257;
  assign n5259 = ~n3410 & ~n5258;
  assign n5260 = controllable_hmaster0 & ~n5259;
  assign n5261 = ~n3821 & ~n5260;
  assign n5262 = controllable_hmaster1 & ~n5261;
  assign n5263 = ~controllable_hmaster1 & ~n3380;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = i_hbusreq3 & ~n5264;
  assign n5266 = i_hbusreq2 & ~n5257;
  assign n5267 = ~i_hbusreq0 & ~n3865;
  assign n5268 = ~n3862 & ~n5267;
  assign n5269 = ~i_hbusreq4 & ~n5268;
  assign n5270 = ~n3861 & ~n5269;
  assign n5271 = ~controllable_hgrant4 & ~n5270;
  assign n5272 = ~n3433 & ~n5271;
  assign n5273 = ~i_hbusreq2 & ~n5272;
  assign n5274 = ~n5266 & ~n5273;
  assign n5275 = ~controllable_hgrant2 & ~n5274;
  assign n5276 = ~n3431 & ~n5275;
  assign n5277 = controllable_hmaster0 & ~n5276;
  assign n5278 = ~controllable_hmaster0 & ~n3399;
  assign n5279 = ~n5277 & ~n5278;
  assign n5280 = controllable_hmaster1 & ~n5279;
  assign n5281 = ~controllable_hmaster1 & ~n3399;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~i_hbusreq3 & ~n5282;
  assign n5284 = ~n5265 & ~n5283;
  assign n5285 = ~controllable_hmaster2 & ~n5284;
  assign n5286 = ~n3957 & ~n5285;
  assign n5287 = controllable_hgrant3 & ~n5286;
  assign n5288 = controllable_hgrant2 & ~n5257;
  assign n5289 = ~controllable_hgrant2 & ~n3380;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~controllable_hmaster0 & ~n5290;
  assign n5292 = ~n3382 & ~n5291;
  assign n5293 = controllable_hmaster1 & ~n5292;
  assign n5294 = controllable_hgrant1 & ~n3414;
  assign n5295 = ~controllable_ndecide & ~n5294;
  assign n5296 = ~controllable_ndecide & ~n5295;
  assign n5297 = i_hready & ~n5296;
  assign n5298 = ~n3379 & ~n5297;
  assign n5299 = ~controllable_hgrant4 & ~n5298;
  assign n5300 = ~n3411 & ~n5299;
  assign n5301 = ~controllable_hgrant2 & ~n5300;
  assign n5302 = ~n3410 & ~n5301;
  assign n5303 = controllable_hmaster0 & ~n5302;
  assign n5304 = ~n3821 & ~n5303;
  assign n5305 = ~controllable_hmaster1 & ~n5304;
  assign n5306 = ~n5293 & ~n5305;
  assign n5307 = i_hbusreq3 & ~n5306;
  assign n5308 = controllable_hgrant2 & ~n5274;
  assign n5309 = ~controllable_hgrant2 & ~n3399;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = ~controllable_hmaster0 & ~n5310;
  assign n5312 = ~n3401 & ~n5311;
  assign n5313 = controllable_hmaster1 & ~n5312;
  assign n5314 = i_hbusreq2 & ~n5300;
  assign n5315 = i_hbusreq4 & ~n5298;
  assign n5316 = i_hbusreq0 & ~n5298;
  assign n5317 = i_hbusreq1 & n5294;
  assign n5318 = ~controllable_ndecide & ~n5317;
  assign n5319 = ~controllable_ndecide & ~n5318;
  assign n5320 = i_hready & ~n5319;
  assign n5321 = ~n3392 & ~n5320;
  assign n5322 = ~i_hbusreq0 & ~n5321;
  assign n5323 = ~n5316 & ~n5322;
  assign n5324 = ~i_hbusreq4 & ~n5323;
  assign n5325 = ~n5315 & ~n5324;
  assign n5326 = ~controllable_hgrant4 & ~n5325;
  assign n5327 = ~n3433 & ~n5326;
  assign n5328 = ~i_hbusreq2 & ~n5327;
  assign n5329 = ~n5314 & ~n5328;
  assign n5330 = ~controllable_hgrant2 & ~n5329;
  assign n5331 = ~n3431 & ~n5330;
  assign n5332 = controllable_hmaster0 & ~n5331;
  assign n5333 = ~n5278 & ~n5332;
  assign n5334 = ~controllable_hmaster1 & ~n5333;
  assign n5335 = ~n5313 & ~n5334;
  assign n5336 = ~i_hbusreq3 & ~n5335;
  assign n5337 = ~n5307 & ~n5336;
  assign n5338 = ~controllable_hmaster2 & ~n5337;
  assign n5339 = ~n3969 & ~n5338;
  assign n5340 = ~controllable_hgrant3 & ~n5339;
  assign n5341 = ~n5287 & ~n5340;
  assign n5342 = controllable_nhgrant0 & ~n5341;
  assign n5343 = ~i_hbusreq3 & ~n3399;
  assign n5344 = ~n3951 & ~n5343;
  assign n5345 = ~controllable_hmaster2 & ~n5344;
  assign n5346 = ~n3957 & ~n5345;
  assign n5347 = controllable_hgrant3 & ~n5346;
  assign n5348 = ~controllable_hmaster0 & ~n5259;
  assign n5349 = ~n3382 & ~n5348;
  assign n5350 = ~controllable_hmaster1 & ~n5349;
  assign n5351 = ~n3381 & ~n5350;
  assign n5352 = i_hbusreq3 & ~n5351;
  assign n5353 = ~controllable_hmaster0 & ~n5276;
  assign n5354 = ~n3401 & ~n5353;
  assign n5355 = ~controllable_hmaster1 & ~n5354;
  assign n5356 = ~n3400 & ~n5355;
  assign n5357 = ~i_hbusreq3 & ~n5356;
  assign n5358 = ~n5352 & ~n5357;
  assign n5359 = ~controllable_hmaster2 & ~n5358;
  assign n5360 = ~n3983 & ~n5359;
  assign n5361 = ~controllable_hgrant3 & ~n5360;
  assign n5362 = ~n5347 & ~n5361;
  assign n5363 = ~controllable_nhgrant0 & ~n5362;
  assign n5364 = ~n5342 & ~n5363;
  assign n5365 = ~n3281 & ~n5364;
  assign n5366 = ~n3950 & ~n5365;
  assign n5367 = n3378 & ~n5366;
  assign n5368 = ~i_hbusreq3 & ~n3834;
  assign n5369 = ~n3951 & ~n5368;
  assign n5370 = controllable_hmaster2 & ~n5369;
  assign n5371 = ~controllable_hgrant4 & ~n3872;
  assign n5372 = ~n3916 & ~n5371;
  assign n5373 = ~i_hbusreq2 & ~n5372;
  assign n5374 = ~n5266 & ~n5373;
  assign n5375 = ~controllable_hgrant2 & ~n5374;
  assign n5376 = ~n3859 & ~n5375;
  assign n5377 = controllable_hmaster0 & ~n5376;
  assign n5378 = ~n3835 & ~n5377;
  assign n5379 = controllable_hmaster1 & ~n5378;
  assign n5380 = ~i_hbusreq1 & controllable_hmastlock;
  assign n5381 = ~i_hbusreq1 & ~n5380;
  assign n5382 = ~controllable_ndecide & n5381;
  assign n5383 = ~controllable_ndecide & ~n5382;
  assign n5384 = ~i_hready & ~n5383;
  assign n5385 = ~i_hready & ~n5384;
  assign n5386 = i_hlock0 & ~n5385;
  assign n5387 = ~n3827 & ~n5386;
  assign n5388 = ~i_hbusreq0 & ~n5387;
  assign n5389 = ~n3389 & ~n5388;
  assign n5390 = ~i_hbusreq4 & ~n5389;
  assign n5391 = ~n3388 & ~n5390;
  assign n5392 = ~i_hbusreq2 & ~n5391;
  assign n5393 = ~n3387 & ~n5392;
  assign n5394 = ~controllable_hmaster0 & ~n5393;
  assign n5395 = ~n4913 & ~n5394;
  assign n5396 = ~controllable_hmaster1 & ~n5395;
  assign n5397 = ~n5379 & ~n5396;
  assign n5398 = ~i_hbusreq3 & ~n5397;
  assign n5399 = ~n5265 & ~n5398;
  assign n5400 = ~controllable_hmaster2 & ~n5399;
  assign n5401 = ~n5370 & ~n5400;
  assign n5402 = controllable_hgrant3 & ~n5401;
  assign n5403 = i_hlock0 & ~n3512;
  assign n5404 = ~i_hlock0 & ~n3496;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~i_hbusreq0 & ~n5405;
  assign n5407 = ~n3509 & ~n5406;
  assign n5408 = ~i_hbusreq4 & ~n5407;
  assign n5409 = ~n3508 & ~n5408;
  assign n5410 = ~controllable_hgrant4 & ~n5409;
  assign n5411 = ~n3916 & ~n5410;
  assign n5412 = ~i_hbusreq2 & ~n5411;
  assign n5413 = ~n3507 & ~n5412;
  assign n5414 = ~controllable_hgrant2 & ~n5413;
  assign n5415 = ~n3859 & ~n5414;
  assign n5416 = controllable_hmaster1 & ~n5415;
  assign n5417 = controllable_hmaster0 & ~n5415;
  assign n5418 = ~n3890 & ~n5417;
  assign n5419 = ~controllable_hmaster1 & ~n5418;
  assign n5420 = ~n5416 & ~n5419;
  assign n5421 = ~i_hbusreq3 & ~n5420;
  assign n5422 = ~n3963 & ~n5421;
  assign n5423 = controllable_hmaster2 & ~n5422;
  assign n5424 = ~n3908 & ~n5288;
  assign n5425 = ~controllable_hmaster0 & ~n5424;
  assign n5426 = ~n5191 & ~n5425;
  assign n5427 = controllable_hmaster1 & ~n5426;
  assign n5428 = ~n3904 & ~n5297;
  assign n5429 = ~controllable_hgrant4 & ~n5428;
  assign n5430 = ~n3411 & ~n5429;
  assign n5431 = ~controllable_hgrant2 & ~n5430;
  assign n5432 = ~n3410 & ~n5431;
  assign n5433 = controllable_hmaster0 & ~n5432;
  assign n5434 = ~n3910 & ~n5433;
  assign n5435 = ~controllable_hmaster1 & ~n5434;
  assign n5436 = ~n5427 & ~n5435;
  assign n5437 = i_hbusreq3 & ~n5436;
  assign n5438 = controllable_hgrant2 & ~n5374;
  assign n5439 = ~n3933 & ~n5438;
  assign n5440 = ~controllable_hmaster0 & ~n5439;
  assign n5441 = ~n5197 & ~n5440;
  assign n5442 = controllable_hmaster1 & ~n5441;
  assign n5443 = i_hbusreq2 & ~n5430;
  assign n5444 = i_hbusreq4 & ~n5428;
  assign n5445 = i_hbusreq0 & ~n5428;
  assign n5446 = ~n3920 & ~n5320;
  assign n5447 = i_hlock0 & ~n5446;
  assign n5448 = ~i_hlock0 & ~n5428;
  assign n5449 = ~n5447 & ~n5448;
  assign n5450 = ~i_hbusreq0 & ~n5449;
  assign n5451 = ~n5445 & ~n5450;
  assign n5452 = ~i_hbusreq4 & ~n5451;
  assign n5453 = ~n5444 & ~n5452;
  assign n5454 = ~controllable_hgrant4 & ~n5453;
  assign n5455 = ~n3916 & ~n5454;
  assign n5456 = ~i_hbusreq2 & ~n5455;
  assign n5457 = ~n5443 & ~n5456;
  assign n5458 = ~controllable_hgrant2 & ~n5457;
  assign n5459 = ~n3859 & ~n5458;
  assign n5460 = controllable_hmaster0 & ~n5459;
  assign n5461 = controllable_hgrant2 & ~n5393;
  assign n5462 = controllable_hgrant4 & ~n5391;
  assign n5463 = ~n3903 & ~n5382;
  assign n5464 = ~i_hready & ~n5463;
  assign n5465 = ~i_hready & ~n5464;
  assign n5466 = i_hlock0 & ~n5465;
  assign n5467 = ~n3923 & ~n5466;
  assign n5468 = ~i_hbusreq0 & ~n5467;
  assign n5469 = ~n3918 & ~n5468;
  assign n5470 = ~i_hbusreq4 & ~n5469;
  assign n5471 = ~n3917 & ~n5470;
  assign n5472 = ~controllable_hgrant4 & ~n5471;
  assign n5473 = ~n5462 & ~n5472;
  assign n5474 = ~i_hbusreq2 & ~n5473;
  assign n5475 = ~n3915 & ~n5474;
  assign n5476 = ~controllable_hgrant2 & ~n5475;
  assign n5477 = ~n5461 & ~n5476;
  assign n5478 = ~controllable_hmaster0 & ~n5477;
  assign n5479 = ~n5460 & ~n5478;
  assign n5480 = ~controllable_hmaster1 & ~n5479;
  assign n5481 = ~n5442 & ~n5480;
  assign n5482 = ~i_hbusreq3 & ~n5481;
  assign n5483 = ~n5437 & ~n5482;
  assign n5484 = ~controllable_hmaster2 & ~n5483;
  assign n5485 = ~n5423 & ~n5484;
  assign n5486 = ~controllable_hgrant3 & ~n5485;
  assign n5487 = ~n5402 & ~n5486;
  assign n5488 = controllable_nhgrant0 & ~n5487;
  assign n5489 = ~n4912 & ~n5396;
  assign n5490 = ~i_hbusreq3 & ~n5489;
  assign n5491 = ~n3951 & ~n5490;
  assign n5492 = ~controllable_hmaster2 & ~n5491;
  assign n5493 = ~n5370 & ~n5492;
  assign n5494 = controllable_hgrant3 & ~n5493;
  assign n5495 = i_hbusreq3 & ~n3909;
  assign n5496 = ~i_hbusreq3 & ~n3934;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = controllable_hmaster2 & ~n5497;
  assign n5499 = ~controllable_hmaster0 & ~n5044;
  assign n5500 = ~n5191 & ~n5499;
  assign n5501 = ~controllable_hmaster1 & ~n5500;
  assign n5502 = ~n5190 & ~n5501;
  assign n5503 = i_hbusreq3 & ~n5502;
  assign n5504 = ~i_hbusreq1 & ~n3708;
  assign n5505 = ~n3436 & ~n5504;
  assign n5506 = ~controllable_ndecide & ~n5505;
  assign n5507 = ~n3418 & ~n5506;
  assign n5508 = i_hready & ~n5507;
  assign n5509 = ~n5038 & ~n5382;
  assign n5510 = ~i_hready & ~n5509;
  assign n5511 = ~n5508 & ~n5510;
  assign n5512 = i_hlock0 & ~n5511;
  assign n5513 = ~n5058 & ~n5512;
  assign n5514 = ~i_hbusreq0 & ~n5513;
  assign n5515 = ~n5053 & ~n5514;
  assign n5516 = ~i_hbusreq4 & ~n5515;
  assign n5517 = ~n5052 & ~n5516;
  assign n5518 = ~controllable_hgrant4 & ~n5517;
  assign n5519 = ~n5462 & ~n5518;
  assign n5520 = ~i_hbusreq2 & ~n5519;
  assign n5521 = ~n5051 & ~n5520;
  assign n5522 = ~controllable_hgrant2 & ~n5521;
  assign n5523 = ~n5461 & ~n5522;
  assign n5524 = ~controllable_hmaster0 & ~n5523;
  assign n5525 = ~n5197 & ~n5524;
  assign n5526 = ~controllable_hmaster1 & ~n5525;
  assign n5527 = ~n5196 & ~n5526;
  assign n5528 = ~i_hbusreq3 & ~n5527;
  assign n5529 = ~n5503 & ~n5528;
  assign n5530 = ~controllable_hmaster2 & ~n5529;
  assign n5531 = ~n5498 & ~n5530;
  assign n5532 = ~controllable_hgrant3 & ~n5531;
  assign n5533 = ~n5494 & ~n5532;
  assign n5534 = ~controllable_nhgrant0 & ~n5533;
  assign n5535 = ~n5488 & ~n5534;
  assign n5536 = ~n3281 & ~n5535;
  assign n5537 = ~n3950 & ~n5536;
  assign n5538 = ~n3378 & ~n5537;
  assign n5539 = ~n5367 & ~n5538;
  assign n5540 = n3492 & ~n5539;
  assign n5541 = ~n3631 & ~n5540;
  assign n5542 = n3485 & ~n5541;
  assign n5543 = ~n3630 & ~n5542;
  assign n5544 = ~n3476 & ~n5543;
  assign n5545 = ~controllable_hgrant4 & ~n4090;
  assign n5546 = ~n3411 & ~n5545;
  assign n5547 = ~controllable_hgrant2 & ~n5546;
  assign n5548 = ~n3410 & ~n5547;
  assign n5549 = i_hbusreq3 & ~n5548;
  assign n5550 = i_hbusreq2 & ~n5546;
  assign n5551 = ~i_hbusreq0 & ~n4108;
  assign n5552 = ~n4107 & ~n5551;
  assign n5553 = ~i_hbusreq4 & ~n5552;
  assign n5554 = ~n4106 & ~n5553;
  assign n5555 = ~controllable_hgrant4 & ~n5554;
  assign n5556 = ~n3433 & ~n5555;
  assign n5557 = ~i_hbusreq2 & ~n5556;
  assign n5558 = ~n5550 & ~n5557;
  assign n5559 = ~controllable_hgrant2 & ~n5558;
  assign n5560 = ~n3431 & ~n5559;
  assign n5561 = controllable_hmaster1 & ~n5560;
  assign n5562 = controllable_hmaster0 & ~n5560;
  assign n5563 = ~n3379 & ~n4031;
  assign n5564 = ~i_hlock0 & ~n5563;
  assign n5565 = ~n4109 & ~n5564;
  assign n5566 = ~i_hbusreq0 & ~n5565;
  assign n5567 = ~n4107 & ~n5566;
  assign n5568 = ~i_hbusreq4 & ~n5567;
  assign n5569 = ~n4106 & ~n5568;
  assign n5570 = ~controllable_hgrant4 & ~n5569;
  assign n5571 = ~n3916 & ~n5570;
  assign n5572 = ~i_hbusreq2 & ~n5571;
  assign n5573 = ~n5550 & ~n5572;
  assign n5574 = ~controllable_hgrant2 & ~n5573;
  assign n5575 = ~n3859 & ~n5574;
  assign n5576 = ~controllable_hmaster0 & ~n5575;
  assign n5577 = ~n5562 & ~n5576;
  assign n5578 = ~controllable_hmaster1 & ~n5577;
  assign n5579 = ~n5561 & ~n5578;
  assign n5580 = ~i_hbusreq3 & ~n5579;
  assign n5581 = ~n5549 & ~n5580;
  assign n5582 = controllable_hmaster2 & ~n5581;
  assign n5583 = ~controllable_hgrant4 & ~n4014;
  assign n5584 = ~n3411 & ~n5583;
  assign n5585 = ~controllable_hgrant2 & ~n5584;
  assign n5586 = ~n3410 & ~n5585;
  assign n5587 = controllable_hmaster0 & ~n5586;
  assign n5588 = ~controllable_hmaster0 & ~n5548;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = controllable_hmaster1 & ~n5589;
  assign n5591 = ~controllable_hmaster1 & ~n5548;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = i_hbusreq3 & ~n5592;
  assign n5594 = i_hbusreq2 & ~n5584;
  assign n5595 = ~i_hbusreq0 & ~n4056;
  assign n5596 = ~n4050 & ~n5595;
  assign n5597 = ~i_hbusreq4 & ~n5596;
  assign n5598 = ~n4049 & ~n5597;
  assign n5599 = ~controllable_hgrant4 & ~n5598;
  assign n5600 = ~n3433 & ~n5599;
  assign n5601 = ~i_hbusreq2 & ~n5600;
  assign n5602 = ~n5594 & ~n5601;
  assign n5603 = ~controllable_hgrant2 & ~n5602;
  assign n5604 = ~n3431 & ~n5603;
  assign n5605 = controllable_hmaster0 & ~n5604;
  assign n5606 = ~controllable_hmaster0 & ~n5560;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = controllable_hmaster1 & ~n5607;
  assign n5609 = ~controllable_hmaster1 & ~n5560;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = ~i_hbusreq3 & ~n5610;
  assign n5612 = ~n5593 & ~n5611;
  assign n5613 = ~controllable_hmaster2 & ~n5612;
  assign n5614 = ~n5582 & ~n5613;
  assign n5615 = controllable_hgrant3 & ~n5614;
  assign n5616 = controllable_hgrant2 & ~n5546;
  assign n5617 = ~controllable_ndecide & n4178;
  assign n5618 = ~n3494 & ~n5617;
  assign n5619 = i_hready & ~n5618;
  assign n5620 = ~n3495 & ~n5619;
  assign n5621 = ~controllable_hgrant4 & ~n5620;
  assign n5622 = ~n4091 & ~n5621;
  assign n5623 = ~controllable_hgrant2 & ~n5622;
  assign n5624 = ~n5616 & ~n5623;
  assign n5625 = controllable_hmaster1 & ~n5624;
  assign n5626 = controllable_hmaster0 & ~n5624;
  assign n5627 = ~n4015 & ~n5621;
  assign n5628 = ~controllable_hgrant2 & ~n5627;
  assign n5629 = ~n5616 & ~n5628;
  assign n5630 = ~controllable_hmaster0 & ~n5629;
  assign n5631 = ~n5626 & ~n5630;
  assign n5632 = ~controllable_hmaster1 & ~n5631;
  assign n5633 = ~n5625 & ~n5632;
  assign n5634 = i_hbusreq3 & ~n5633;
  assign n5635 = controllable_hgrant2 & ~n5558;
  assign n5636 = i_hbusreq2 & ~n5622;
  assign n5637 = i_hbusreq4 & ~n5620;
  assign n5638 = i_hbusreq0 & ~n5620;
  assign n5639 = i_hbusreq1 & n4178;
  assign n5640 = i_hbusreq1 & ~n5639;
  assign n5641 = ~controllable_ndecide & ~n5640;
  assign n5642 = ~n3494 & ~n5641;
  assign n5643 = i_hready & ~n5642;
  assign n5644 = ~n3511 & ~n5643;
  assign n5645 = ~i_hbusreq0 & ~n5644;
  assign n5646 = ~n5638 & ~n5645;
  assign n5647 = ~i_hbusreq4 & ~n5646;
  assign n5648 = ~n5637 & ~n5647;
  assign n5649 = ~controllable_hgrant4 & ~n5648;
  assign n5650 = ~n4117 & ~n5649;
  assign n5651 = ~i_hbusreq2 & ~n5650;
  assign n5652 = ~n5636 & ~n5651;
  assign n5653 = ~controllable_hgrant2 & ~n5652;
  assign n5654 = ~n5635 & ~n5653;
  assign n5655 = controllable_hmaster1 & ~n5654;
  assign n5656 = controllable_hmaster0 & ~n5654;
  assign n5657 = controllable_hgrant2 & ~n5573;
  assign n5658 = i_hbusreq2 & ~n5627;
  assign n5659 = i_hlock0 & ~n5644;
  assign n5660 = ~n3495 & ~n5643;
  assign n5661 = ~i_hlock0 & ~n5660;
  assign n5662 = ~n5659 & ~n5661;
  assign n5663 = ~i_hbusreq0 & ~n5662;
  assign n5664 = ~n5638 & ~n5663;
  assign n5665 = ~i_hbusreq4 & ~n5664;
  assign n5666 = ~n5637 & ~n5665;
  assign n5667 = ~controllable_hgrant4 & ~n5666;
  assign n5668 = ~n4064 & ~n5667;
  assign n5669 = ~i_hbusreq2 & ~n5668;
  assign n5670 = ~n5658 & ~n5669;
  assign n5671 = ~controllable_hgrant2 & ~n5670;
  assign n5672 = ~n5657 & ~n5671;
  assign n5673 = ~controllable_hmaster0 & ~n5672;
  assign n5674 = ~n5656 & ~n5673;
  assign n5675 = ~controllable_hmaster1 & ~n5674;
  assign n5676 = ~n5655 & ~n5675;
  assign n5677 = ~i_hbusreq3 & ~n5676;
  assign n5678 = ~n5634 & ~n5677;
  assign n5679 = controllable_hmaster2 & ~n5678;
  assign n5680 = ~n3379 & ~n5619;
  assign n5681 = ~controllable_hgrant4 & ~n5680;
  assign n5682 = ~n4091 & ~n5681;
  assign n5683 = ~controllable_hgrant2 & ~n5682;
  assign n5684 = ~n5616 & ~n5683;
  assign n5685 = controllable_hmaster0 & ~n5684;
  assign n5686 = controllable_hgrant2 & ~n5584;
  assign n5687 = ~n5683 & ~n5686;
  assign n5688 = ~controllable_hmaster0 & ~n5687;
  assign n5689 = ~n5685 & ~n5688;
  assign n5690 = controllable_hmaster1 & ~n5689;
  assign n5691 = controllable_hgrant1 & ~n4008;
  assign n5692 = controllable_hgrant1 & ~n5691;
  assign n5693 = ~controllable_ndecide & n5692;
  assign n5694 = ~n3494 & ~n5693;
  assign n5695 = i_hready & ~n5694;
  assign n5696 = ~n3379 & ~n5695;
  assign n5697 = ~controllable_hgrant4 & ~n5696;
  assign n5698 = ~n4091 & ~n5697;
  assign n5699 = ~controllable_hgrant2 & ~n5698;
  assign n5700 = ~n5616 & ~n5699;
  assign n5701 = controllable_hmaster0 & ~n5700;
  assign n5702 = ~controllable_hmaster0 & ~n5684;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = ~controllable_hmaster1 & ~n5703;
  assign n5705 = ~n5690 & ~n5704;
  assign n5706 = i_hbusreq3 & ~n5705;
  assign n5707 = i_hbusreq2 & ~n5682;
  assign n5708 = i_hbusreq4 & ~n5680;
  assign n5709 = i_hbusreq0 & ~n5680;
  assign n5710 = ~n3392 & ~n5643;
  assign n5711 = ~i_hbusreq0 & ~n5710;
  assign n5712 = ~n5709 & ~n5711;
  assign n5713 = ~i_hbusreq4 & ~n5712;
  assign n5714 = ~n5708 & ~n5713;
  assign n5715 = ~controllable_hgrant4 & ~n5714;
  assign n5716 = ~n4117 & ~n5715;
  assign n5717 = ~i_hbusreq2 & ~n5716;
  assign n5718 = ~n5707 & ~n5717;
  assign n5719 = ~controllable_hgrant2 & ~n5718;
  assign n5720 = ~n5635 & ~n5719;
  assign n5721 = controllable_hmaster0 & ~n5720;
  assign n5722 = controllable_hgrant2 & ~n5602;
  assign n5723 = ~n5719 & ~n5722;
  assign n5724 = ~controllable_hmaster0 & ~n5723;
  assign n5725 = ~n5721 & ~n5724;
  assign n5726 = controllable_hmaster1 & ~n5725;
  assign n5727 = i_hbusreq2 & ~n5698;
  assign n5728 = i_hbusreq4 & ~n5696;
  assign n5729 = i_hbusreq0 & ~n5696;
  assign n5730 = i_hbusreq1 & ~n5692;
  assign n5731 = ~controllable_ndecide & ~n5730;
  assign n5732 = ~n3494 & ~n5731;
  assign n5733 = i_hready & ~n5732;
  assign n5734 = ~n3392 & ~n5733;
  assign n5735 = ~i_hbusreq0 & ~n5734;
  assign n5736 = ~n5729 & ~n5735;
  assign n5737 = ~i_hbusreq4 & ~n5736;
  assign n5738 = ~n5728 & ~n5737;
  assign n5739 = ~controllable_hgrant4 & ~n5738;
  assign n5740 = ~n4117 & ~n5739;
  assign n5741 = ~i_hbusreq2 & ~n5740;
  assign n5742 = ~n5727 & ~n5741;
  assign n5743 = ~controllable_hgrant2 & ~n5742;
  assign n5744 = ~n5635 & ~n5743;
  assign n5745 = controllable_hmaster0 & ~n5744;
  assign n5746 = ~controllable_hmaster0 & ~n5720;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~controllable_hmaster1 & ~n5747;
  assign n5749 = ~n5726 & ~n5748;
  assign n5750 = ~i_hbusreq3 & ~n5749;
  assign n5751 = ~n5706 & ~n5750;
  assign n5752 = ~controllable_hmaster2 & ~n5751;
  assign n5753 = ~n5679 & ~n5752;
  assign n5754 = ~controllable_hgrant3 & ~n5753;
  assign n5755 = ~n5615 & ~n5754;
  assign n5756 = controllable_nhgrant0 & ~n5755;
  assign n5757 = controllable_hmaster1 & ~n5548;
  assign n5758 = controllable_hmaster0 & ~n5548;
  assign n5759 = ~n3904 & ~n4000;
  assign n5760 = ~controllable_hgrant4 & ~n5759;
  assign n5761 = ~n3411 & ~n5760;
  assign n5762 = ~controllable_hgrant2 & ~n5761;
  assign n5763 = ~n3410 & ~n5762;
  assign n5764 = ~controllable_hmaster0 & ~n5763;
  assign n5765 = ~n5758 & ~n5764;
  assign n5766 = ~controllable_hmaster1 & ~n5765;
  assign n5767 = ~n5757 & ~n5766;
  assign n5768 = i_hbusreq3 & ~n5767;
  assign n5769 = i_hbusreq2 & ~n5761;
  assign n5770 = i_hbusreq4 & ~n5759;
  assign n5771 = i_hbusreq0 & ~n5759;
  assign n5772 = ~n3920 & ~n4031;
  assign n5773 = i_hlock0 & ~n5772;
  assign n5774 = ~n3904 & ~n4031;
  assign n5775 = ~i_hlock0 & ~n5774;
  assign n5776 = ~n5773 & ~n5775;
  assign n5777 = ~i_hbusreq0 & ~n5776;
  assign n5778 = ~n5771 & ~n5777;
  assign n5779 = ~i_hbusreq4 & ~n5778;
  assign n5780 = ~n5770 & ~n5779;
  assign n5781 = ~controllable_hgrant4 & ~n5780;
  assign n5782 = ~n3916 & ~n5781;
  assign n5783 = ~i_hbusreq2 & ~n5782;
  assign n5784 = ~n5769 & ~n5783;
  assign n5785 = ~controllable_hgrant2 & ~n5784;
  assign n5786 = ~n3859 & ~n5785;
  assign n5787 = ~controllable_hmaster0 & ~n5786;
  assign n5788 = ~n5562 & ~n5787;
  assign n5789 = ~controllable_hmaster1 & ~n5788;
  assign n5790 = ~n5561 & ~n5789;
  assign n5791 = ~i_hbusreq3 & ~n5790;
  assign n5792 = ~n5768 & ~n5791;
  assign n5793 = controllable_hmaster2 & ~n5792;
  assign n5794 = ~controllable_hmaster0 & ~n5586;
  assign n5795 = ~n5758 & ~n5794;
  assign n5796 = ~controllable_hmaster1 & ~n5795;
  assign n5797 = ~n5757 & ~n5796;
  assign n5798 = i_hbusreq3 & ~n5797;
  assign n5799 = ~controllable_hmaster0 & ~n5604;
  assign n5800 = ~n5562 & ~n5799;
  assign n5801 = ~controllable_hmaster1 & ~n5800;
  assign n5802 = ~n5561 & ~n5801;
  assign n5803 = ~i_hbusreq3 & ~n5802;
  assign n5804 = ~n5798 & ~n5803;
  assign n5805 = ~controllable_hmaster2 & ~n5804;
  assign n5806 = ~n5793 & ~n5805;
  assign n5807 = ~controllable_hgrant3 & ~n5806;
  assign n5808 = ~n5347 & ~n5807;
  assign n5809 = ~controllable_nhgrant0 & ~n5808;
  assign n5810 = ~n5756 & ~n5809;
  assign n5811 = ~n3281 & ~n5810;
  assign n5812 = ~n4089 & ~n5811;
  assign n5813 = n3378 & ~n5812;
  assign n5814 = ~i_hlock0 & ~n4090;
  assign n5815 = ~n4109 & ~n5814;
  assign n5816 = ~i_hbusreq0 & ~n5815;
  assign n5817 = ~n4107 & ~n5816;
  assign n5818 = ~i_hbusreq4 & ~n5817;
  assign n5819 = ~n4106 & ~n5818;
  assign n5820 = ~controllable_hgrant4 & ~n5819;
  assign n5821 = ~n3916 & ~n5820;
  assign n5822 = ~i_hbusreq2 & ~n5821;
  assign n5823 = ~n5550 & ~n5822;
  assign n5824 = ~controllable_hgrant2 & ~n5823;
  assign n5825 = ~n3859 & ~n5824;
  assign n5826 = ~i_hbusreq3 & ~n5825;
  assign n5827 = ~n5549 & ~n5826;
  assign n5828 = controllable_hmaster2 & ~n5827;
  assign n5829 = ~controllable_hgrant4 & ~n4063;
  assign n5830 = ~n3916 & ~n5829;
  assign n5831 = ~i_hbusreq2 & ~n5830;
  assign n5832 = ~n5594 & ~n5831;
  assign n5833 = ~controllable_hgrant2 & ~n5832;
  assign n5834 = ~n3859 & ~n5833;
  assign n5835 = controllable_hmaster0 & ~n5834;
  assign n5836 = ~controllable_hmaster0 & ~n5825;
  assign n5837 = ~n5835 & ~n5836;
  assign n5838 = controllable_hmaster1 & ~n5837;
  assign n5839 = controllable_hmaster0 & ~n5825;
  assign n5840 = ~n4031 & ~n5384;
  assign n5841 = i_hlock0 & ~n5840;
  assign n5842 = ~n5814 & ~n5841;
  assign n5843 = ~i_hbusreq0 & ~n5842;
  assign n5844 = ~n4107 & ~n5843;
  assign n5845 = ~i_hbusreq4 & ~n5844;
  assign n5846 = ~n4106 & ~n5845;
  assign n5847 = ~controllable_hgrant4 & ~n5846;
  assign n5848 = ~n5462 & ~n5847;
  assign n5849 = ~i_hbusreq2 & ~n5848;
  assign n5850 = ~n5550 & ~n5849;
  assign n5851 = ~controllable_hgrant2 & ~n5850;
  assign n5852 = ~n5461 & ~n5851;
  assign n5853 = ~controllable_hmaster0 & ~n5852;
  assign n5854 = ~n5839 & ~n5853;
  assign n5855 = ~controllable_hmaster1 & ~n5854;
  assign n5856 = ~n5838 & ~n5855;
  assign n5857 = ~i_hbusreq3 & ~n5856;
  assign n5858 = ~n5593 & ~n5857;
  assign n5859 = ~controllable_hmaster2 & ~n5858;
  assign n5860 = ~n5828 & ~n5859;
  assign n5861 = controllable_hgrant3 & ~n5860;
  assign n5862 = controllable_hgrant2 & ~n5823;
  assign n5863 = controllable_hgrant4 & ~n5819;
  assign n5864 = ~n4009 & ~n4178;
  assign n5865 = ~i_hbusreq1 & ~n5864;
  assign n5866 = ~n5639 & ~n5865;
  assign n5867 = ~controllable_ndecide & ~n5866;
  assign n5868 = ~n3494 & ~n5867;
  assign n5869 = i_hready & ~n5868;
  assign n5870 = ~n3495 & ~n5869;
  assign n5871 = ~i_hlock0 & ~n5870;
  assign n5872 = ~n5659 & ~n5871;
  assign n5873 = ~i_hbusreq0 & ~n5872;
  assign n5874 = ~n5638 & ~n5873;
  assign n5875 = ~i_hbusreq4 & ~n5874;
  assign n5876 = ~n5637 & ~n5875;
  assign n5877 = ~controllable_hgrant4 & ~n5876;
  assign n5878 = ~n5863 & ~n5877;
  assign n5879 = ~i_hbusreq2 & ~n5878;
  assign n5880 = ~n5636 & ~n5879;
  assign n5881 = ~controllable_hgrant2 & ~n5880;
  assign n5882 = ~n5862 & ~n5881;
  assign n5883 = controllable_hmaster1 & ~n5882;
  assign n5884 = controllable_hmaster0 & ~n5882;
  assign n5885 = ~i_hbusreq1 & controllable_locked;
  assign n5886 = ~n5639 & ~n5885;
  assign n5887 = ~controllable_ndecide & ~n5886;
  assign n5888 = ~n3494 & ~n5887;
  assign n5889 = i_hready & ~n5888;
  assign n5890 = ~n3495 & ~n5889;
  assign n5891 = ~i_hlock0 & ~n5890;
  assign n5892 = ~n5659 & ~n5891;
  assign n5893 = ~i_hbusreq0 & ~n5892;
  assign n5894 = ~n5638 & ~n5893;
  assign n5895 = ~i_hbusreq4 & ~n5894;
  assign n5896 = ~n5637 & ~n5895;
  assign n5897 = ~controllable_hgrant4 & ~n5896;
  assign n5898 = ~n4064 & ~n5897;
  assign n5899 = ~i_hbusreq2 & ~n5898;
  assign n5900 = ~n5658 & ~n5899;
  assign n5901 = ~controllable_hgrant2 & ~n5900;
  assign n5902 = ~n5862 & ~n5901;
  assign n5903 = ~controllable_hmaster0 & ~n5902;
  assign n5904 = ~n5884 & ~n5903;
  assign n5905 = ~controllable_hmaster1 & ~n5904;
  assign n5906 = ~n5883 & ~n5905;
  assign n5907 = ~i_hbusreq3 & ~n5906;
  assign n5908 = ~n5634 & ~n5907;
  assign n5909 = controllable_hmaster2 & ~n5908;
  assign n5910 = ~n3904 & ~n5619;
  assign n5911 = ~controllable_hgrant4 & ~n5910;
  assign n5912 = ~n4091 & ~n5911;
  assign n5913 = ~controllable_hgrant2 & ~n5912;
  assign n5914 = ~n5616 & ~n5913;
  assign n5915 = controllable_hmaster0 & ~n5914;
  assign n5916 = ~n5686 & ~n5913;
  assign n5917 = ~controllable_hmaster0 & ~n5916;
  assign n5918 = ~n5915 & ~n5917;
  assign n5919 = controllable_hmaster1 & ~n5918;
  assign n5920 = ~n3904 & ~n5695;
  assign n5921 = ~controllable_hgrant4 & ~n5920;
  assign n5922 = ~n4091 & ~n5921;
  assign n5923 = ~controllable_hgrant2 & ~n5922;
  assign n5924 = ~n5616 & ~n5923;
  assign n5925 = controllable_hmaster0 & ~n5924;
  assign n5926 = ~controllable_hmaster0 & ~n5914;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~controllable_hmaster1 & ~n5927;
  assign n5929 = ~n5919 & ~n5928;
  assign n5930 = i_hbusreq3 & ~n5929;
  assign n5931 = i_hbusreq2 & ~n5912;
  assign n5932 = i_hbusreq4 & ~n5910;
  assign n5933 = i_hbusreq0 & ~n5910;
  assign n5934 = ~n3920 & ~n5643;
  assign n5935 = i_hlock0 & ~n5934;
  assign n5936 = ~n3904 & ~n5889;
  assign n5937 = ~i_hlock0 & ~n5936;
  assign n5938 = ~n5935 & ~n5937;
  assign n5939 = ~i_hbusreq0 & ~n5938;
  assign n5940 = ~n5933 & ~n5939;
  assign n5941 = ~i_hbusreq4 & ~n5940;
  assign n5942 = ~n5932 & ~n5941;
  assign n5943 = ~controllable_hgrant4 & ~n5942;
  assign n5944 = ~n5863 & ~n5943;
  assign n5945 = ~i_hbusreq2 & ~n5944;
  assign n5946 = ~n5931 & ~n5945;
  assign n5947 = ~controllable_hgrant2 & ~n5946;
  assign n5948 = ~n5862 & ~n5947;
  assign n5949 = controllable_hmaster0 & ~n5948;
  assign n5950 = controllable_hgrant2 & ~n5832;
  assign n5951 = ~n5947 & ~n5950;
  assign n5952 = ~controllable_hmaster0 & ~n5951;
  assign n5953 = ~n5949 & ~n5952;
  assign n5954 = controllable_hmaster1 & ~n5953;
  assign n5955 = i_hbusreq2 & ~n5922;
  assign n5956 = i_hbusreq4 & ~n5920;
  assign n5957 = i_hbusreq0 & ~n5920;
  assign n5958 = ~n3920 & ~n5733;
  assign n5959 = i_hlock0 & ~n5958;
  assign n5960 = ~controllable_hgrant1 & ~controllable_locked;
  assign n5961 = ~n5691 & ~n5960;
  assign n5962 = ~i_hbusreq1 & ~n5961;
  assign n5963 = ~n5730 & ~n5962;
  assign n5964 = ~controllable_ndecide & n5963;
  assign n5965 = ~n3494 & ~n5964;
  assign n5966 = i_hready & ~n5965;
  assign n5967 = ~n3904 & ~n5966;
  assign n5968 = ~i_hlock0 & ~n5967;
  assign n5969 = ~n5959 & ~n5968;
  assign n5970 = ~i_hbusreq0 & ~n5969;
  assign n5971 = ~n5957 & ~n5970;
  assign n5972 = ~i_hbusreq4 & ~n5971;
  assign n5973 = ~n5956 & ~n5972;
  assign n5974 = ~controllable_hgrant4 & ~n5973;
  assign n5975 = ~n5863 & ~n5974;
  assign n5976 = ~i_hbusreq2 & ~n5975;
  assign n5977 = ~n5955 & ~n5976;
  assign n5978 = ~controllable_hgrant2 & ~n5977;
  assign n5979 = ~n5862 & ~n5978;
  assign n5980 = controllable_hmaster0 & ~n5979;
  assign n5981 = controllable_hgrant2 & ~n5850;
  assign n5982 = controllable_hgrant4 & ~n5846;
  assign n5983 = ~n5464 & ~n5643;
  assign n5984 = i_hlock0 & ~n5983;
  assign n5985 = ~n5937 & ~n5984;
  assign n5986 = ~i_hbusreq0 & ~n5985;
  assign n5987 = ~n5933 & ~n5986;
  assign n5988 = ~i_hbusreq4 & ~n5987;
  assign n5989 = ~n5932 & ~n5988;
  assign n5990 = ~controllable_hgrant4 & ~n5989;
  assign n5991 = ~n5982 & ~n5990;
  assign n5992 = ~i_hbusreq2 & ~n5991;
  assign n5993 = ~n5931 & ~n5992;
  assign n5994 = ~controllable_hgrant2 & ~n5993;
  assign n5995 = ~n5981 & ~n5994;
  assign n5996 = ~controllable_hmaster0 & ~n5995;
  assign n5997 = ~n5980 & ~n5996;
  assign n5998 = ~controllable_hmaster1 & ~n5997;
  assign n5999 = ~n5954 & ~n5998;
  assign n6000 = ~i_hbusreq3 & ~n5999;
  assign n6001 = ~n5930 & ~n6000;
  assign n6002 = ~controllable_hmaster2 & ~n6001;
  assign n6003 = ~n5909 & ~n6002;
  assign n6004 = ~controllable_hgrant3 & ~n6003;
  assign n6005 = ~n5861 & ~n6004;
  assign n6006 = controllable_nhgrant0 & ~n6005;
  assign n6007 = i_hready & ~n3902;
  assign n6008 = ~n3904 & ~n6007;
  assign n6009 = ~controllable_hgrant4 & ~n6008;
  assign n6010 = ~n3411 & ~n6009;
  assign n6011 = ~controllable_hgrant2 & ~n6010;
  assign n6012 = ~n3410 & ~n6011;
  assign n6013 = i_hbusreq3 & ~n6012;
  assign n6014 = i_hbusreq2 & ~n6010;
  assign n6015 = i_hbusreq4 & ~n6008;
  assign n6016 = i_hbusreq0 & ~n6008;
  assign n6017 = ~n3903 & ~n4029;
  assign n6018 = i_hready & ~n6017;
  assign n6019 = ~n3920 & ~n6018;
  assign n6020 = i_hlock0 & ~n6019;
  assign n6021 = ~i_hlock0 & ~n6008;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = ~i_hbusreq0 & ~n6022;
  assign n6024 = ~n6016 & ~n6023;
  assign n6025 = ~i_hbusreq4 & ~n6024;
  assign n6026 = ~n6015 & ~n6025;
  assign n6027 = ~controllable_hgrant4 & ~n6026;
  assign n6028 = ~n3916 & ~n6027;
  assign n6029 = ~i_hbusreq2 & ~n6028;
  assign n6030 = ~n6014 & ~n6029;
  assign n6031 = ~controllable_hgrant2 & ~n6030;
  assign n6032 = ~n3859 & ~n6031;
  assign n6033 = ~i_hbusreq3 & ~n6032;
  assign n6034 = ~n6013 & ~n6033;
  assign n6035 = controllable_hmaster2 & ~n6034;
  assign n6036 = controllable_hmaster1 & ~n6012;
  assign n6037 = controllable_hmaster0 & ~n6012;
  assign n6038 = i_hready & ~n4010;
  assign n6039 = ~n5039 & ~n6038;
  assign n6040 = ~controllable_hgrant4 & ~n6039;
  assign n6041 = ~n3411 & ~n6040;
  assign n6042 = ~controllable_hgrant2 & ~n6041;
  assign n6043 = ~n3410 & ~n6042;
  assign n6044 = ~controllable_hmaster0 & ~n6043;
  assign n6045 = ~n6037 & ~n6044;
  assign n6046 = ~controllable_hmaster1 & ~n6045;
  assign n6047 = ~n6036 & ~n6046;
  assign n6048 = i_hbusreq3 & ~n6047;
  assign n6049 = controllable_hmaster1 & ~n6032;
  assign n6050 = controllable_hmaster0 & ~n6032;
  assign n6051 = i_hbusreq2 & ~n6041;
  assign n6052 = i_hbusreq4 & ~n6039;
  assign n6053 = i_hbusreq0 & ~n6039;
  assign n6054 = ~n4051 & ~n5504;
  assign n6055 = ~controllable_ndecide & ~n6054;
  assign n6056 = ~n5038 & ~n6055;
  assign n6057 = i_hready & ~n6056;
  assign n6058 = ~n5510 & ~n6057;
  assign n6059 = i_hlock0 & ~n6058;
  assign n6060 = ~i_hlock0 & ~n6039;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~i_hbusreq0 & ~n6061;
  assign n6063 = ~n6053 & ~n6062;
  assign n6064 = ~i_hbusreq4 & ~n6063;
  assign n6065 = ~n6052 & ~n6064;
  assign n6066 = ~controllable_hgrant4 & ~n6065;
  assign n6067 = ~n5462 & ~n6066;
  assign n6068 = ~i_hbusreq2 & ~n6067;
  assign n6069 = ~n6051 & ~n6068;
  assign n6070 = ~controllable_hgrant2 & ~n6069;
  assign n6071 = ~n5461 & ~n6070;
  assign n6072 = ~controllable_hmaster0 & ~n6071;
  assign n6073 = ~n6050 & ~n6072;
  assign n6074 = ~controllable_hmaster1 & ~n6073;
  assign n6075 = ~n6049 & ~n6074;
  assign n6076 = ~i_hbusreq3 & ~n6075;
  assign n6077 = ~n6048 & ~n6076;
  assign n6078 = ~controllable_hmaster2 & ~n6077;
  assign n6079 = ~n6035 & ~n6078;
  assign n6080 = ~controllable_hgrant3 & ~n6079;
  assign n6081 = ~n5494 & ~n6080;
  assign n6082 = ~controllable_nhgrant0 & ~n6081;
  assign n6083 = ~n6006 & ~n6082;
  assign n6084 = ~n3281 & ~n6083;
  assign n6085 = ~n4089 & ~n6084;
  assign n6086 = ~n3378 & ~n6085;
  assign n6087 = ~n5813 & ~n6086;
  assign n6088 = n3492 & ~n6087;
  assign n6089 = ~n3631 & ~n6088;
  assign n6090 = n3485 & ~n6089;
  assign n6091 = ~n3630 & ~n6090;
  assign n6092 = n3476 & ~n6091;
  assign n6093 = ~n5544 & ~n6092;
  assign n6094 = n3374 & ~n6093;
  assign n6095 = ~n5255 & ~n6094;
  assign n6096 = n3655 & ~n6095;
  assign n6097 = controllable_ndecide & ~n5864;
  assign n6098 = ~i_hready & n6097;
  assign n6099 = ~n3417 & ~n6098;
  assign n6100 = ~controllable_hgrant4 & ~n6099;
  assign n6101 = ~n3411 & ~n6100;
  assign n6102 = ~controllable_hgrant2 & ~n6101;
  assign n6103 = ~n3410 & ~n6102;
  assign n6104 = controllable_hmaster1 & ~n6103;
  assign n6105 = controllable_hmaster0 & ~n6103;
  assign n6106 = ~n3729 & ~n6105;
  assign n6107 = ~controllable_hmaster1 & ~n6106;
  assign n6108 = ~n6104 & ~n6107;
  assign n6109 = i_hbusreq3 & ~n6108;
  assign n6110 = i_hbusreq2 & ~n6101;
  assign n6111 = i_hbusreq4 & ~n6099;
  assign n6112 = i_hbusreq0 & ~n6099;
  assign n6113 = ~n3390 & ~n6097;
  assign n6114 = ~i_hready & ~n6113;
  assign n6115 = ~n3440 & ~n6114;
  assign n6116 = i_hlock0 & ~n6115;
  assign n6117 = ~i_hlock0 & ~n6099;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = ~i_hbusreq0 & ~n6118;
  assign n6120 = ~n6112 & ~n6119;
  assign n6121 = ~i_hbusreq4 & ~n6120;
  assign n6122 = ~n6111 & ~n6121;
  assign n6123 = ~controllable_hgrant4 & ~n6122;
  assign n6124 = ~n3916 & ~n6123;
  assign n6125 = ~i_hbusreq2 & ~n6124;
  assign n6126 = ~n6110 & ~n6125;
  assign n6127 = ~controllable_hgrant2 & ~n6126;
  assign n6128 = ~n3859 & ~n6127;
  assign n6129 = controllable_hmaster1 & ~n6128;
  assign n6130 = controllable_hmaster0 & ~n6128;
  assign n6131 = ~n3767 & ~n6130;
  assign n6132 = ~controllable_hmaster1 & ~n6131;
  assign n6133 = ~n6129 & ~n6132;
  assign n6134 = ~i_hbusreq3 & ~n6133;
  assign n6135 = ~n6109 & ~n6134;
  assign n6136 = controllable_hmaster2 & ~n6135;
  assign n6137 = controllable_ndecide & n5294;
  assign n6138 = ~controllable_ndecide & ~n5094;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = i_hready & ~n6139;
  assign n6141 = ~controllable_ndecide & ~n4935;
  assign n6142 = ~n6137 & ~n6141;
  assign n6143 = ~i_hready & ~n6142;
  assign n6144 = ~n6140 & ~n6143;
  assign n6145 = ~controllable_hgrant4 & n6144;
  assign n6146 = ~n5089 & ~n6145;
  assign n6147 = ~controllable_hgrant2 & ~n6146;
  assign n6148 = ~n5088 & ~n6147;
  assign n6149 = controllable_hmaster0 & ~n6148;
  assign n6150 = ~n4944 & ~n6149;
  assign n6151 = ~controllable_hmaster1 & ~n6150;
  assign n6152 = ~n5087 & ~n6151;
  assign n6153 = i_hlock3 & ~n6152;
  assign n6154 = ~n5110 & ~n6151;
  assign n6155 = ~i_hlock3 & ~n6154;
  assign n6156 = ~n6153 & ~n6155;
  assign n6157 = i_hbusreq3 & ~n6156;
  assign n6158 = i_hbusreq2 & ~n6146;
  assign n6159 = i_hbusreq4 & ~n6144;
  assign n6160 = i_hbusreq0 & ~n6144;
  assign n6161 = ~controllable_ndecide & n5133;
  assign n6162 = ~n6137 & ~n6161;
  assign n6163 = i_hready & ~n6162;
  assign n6164 = ~controllable_ndecide & n4996;
  assign n6165 = ~n6137 & ~n6164;
  assign n6166 = ~i_hready & ~n6165;
  assign n6167 = ~n6163 & ~n6166;
  assign n6168 = ~i_hbusreq0 & ~n6167;
  assign n6169 = ~n6160 & ~n6168;
  assign n6170 = ~i_hbusreq4 & ~n6169;
  assign n6171 = ~n6159 & ~n6170;
  assign n6172 = ~controllable_hgrant4 & n6171;
  assign n6173 = ~n5130 & ~n6172;
  assign n6174 = ~i_hbusreq2 & ~n6173;
  assign n6175 = ~n6158 & ~n6174;
  assign n6176 = ~controllable_hgrant2 & ~n6175;
  assign n6177 = ~n5128 & ~n6176;
  assign n6178 = controllable_hmaster0 & ~n6177;
  assign n6179 = ~n4944 & ~n6178;
  assign n6180 = ~controllable_hmaster1 & ~n6179;
  assign n6181 = ~n5127 & ~n6180;
  assign n6182 = i_hlock3 & ~n6181;
  assign n6183 = ~n5155 & ~n6180;
  assign n6184 = ~i_hlock3 & ~n6183;
  assign n6185 = ~n6182 & ~n6184;
  assign n6186 = ~i_hbusreq3 & ~n6185;
  assign n6187 = ~n6157 & ~n6186;
  assign n6188 = ~controllable_hmaster2 & ~n6187;
  assign n6189 = ~n6136 & ~n6188;
  assign n6190 = ~controllable_hgrant3 & ~n6189;
  assign n6191 = ~n5037 & ~n6190;
  assign n6192 = controllable_nhgrant0 & ~n6191;
  assign n6193 = ~n5245 & ~n6192;
  assign n6194 = ~n3281 & ~n6193;
  assign n6195 = ~n3783 & ~n6194;
  assign n6196 = ~n3378 & ~n6195;
  assign n6197 = ~n4911 & ~n6196;
  assign n6198 = n3492 & ~n6197;
  assign n6199 = ~n3631 & ~n6198;
  assign n6200 = n3485 & ~n6199;
  assign n6201 = ~n3630 & ~n6200;
  assign n6202 = ~n3374 & ~n6201;
  assign n6203 = ~n4234 & ~n5338;
  assign n6204 = ~controllable_hgrant3 & ~n6203;
  assign n6205 = ~n5287 & ~n6204;
  assign n6206 = controllable_nhgrant0 & ~n6205;
  assign n6207 = ~n5363 & ~n6206;
  assign n6208 = ~n3281 & ~n6207;
  assign n6209 = ~n3950 & ~n6208;
  assign n6210 = n3378 & ~n6209;
  assign n6211 = ~n3417 & ~n4180;
  assign n6212 = ~controllable_hgrant4 & ~n6211;
  assign n6213 = ~n3411 & ~n6212;
  assign n6214 = ~controllable_hgrant2 & ~n6213;
  assign n6215 = ~n3410 & ~n6214;
  assign n6216 = controllable_hmaster1 & ~n6215;
  assign n6217 = controllable_hmaster0 & ~n6215;
  assign n6218 = ~n4186 & ~n6217;
  assign n6219 = ~controllable_hmaster1 & ~n6218;
  assign n6220 = ~n6216 & ~n6219;
  assign n6221 = i_hbusreq3 & ~n6220;
  assign n6222 = i_hbusreq2 & ~n6213;
  assign n6223 = i_hbusreq4 & ~n6211;
  assign n6224 = i_hbusreq0 & ~n6211;
  assign n6225 = ~n3440 & ~n4195;
  assign n6226 = i_hlock0 & ~n6225;
  assign n6227 = ~i_hlock0 & ~n6211;
  assign n6228 = ~n6226 & ~n6227;
  assign n6229 = ~i_hbusreq0 & ~n6228;
  assign n6230 = ~n6224 & ~n6229;
  assign n6231 = ~i_hbusreq4 & ~n6230;
  assign n6232 = ~n6223 & ~n6231;
  assign n6233 = ~controllable_hgrant4 & ~n6232;
  assign n6234 = ~n3916 & ~n6233;
  assign n6235 = ~i_hbusreq2 & ~n6234;
  assign n6236 = ~n6222 & ~n6235;
  assign n6237 = ~controllable_hgrant2 & ~n6236;
  assign n6238 = ~n3859 & ~n6237;
  assign n6239 = controllable_hmaster1 & ~n6238;
  assign n6240 = controllable_hmaster0 & ~n6238;
  assign n6241 = ~n4210 & ~n6240;
  assign n6242 = ~controllable_hmaster1 & ~n6241;
  assign n6243 = ~n6239 & ~n6242;
  assign n6244 = ~i_hbusreq3 & ~n6243;
  assign n6245 = ~n6221 & ~n6244;
  assign n6246 = controllable_hmaster2 & ~n6245;
  assign n6247 = controllable_locked & controllable_ndecide;
  assign n6248 = ~i_hready & n6247;
  assign n6249 = ~i_hready & ~n6248;
  assign n6250 = ~controllable_hgrant4 & ~n6249;
  assign n6251 = ~n3411 & ~n6250;
  assign n6252 = ~controllable_hgrant2 & ~n6251;
  assign n6253 = ~n3410 & ~n6252;
  assign n6254 = controllable_hmaster0 & ~n6253;
  assign n6255 = ~n5288 & ~n6252;
  assign n6256 = ~controllable_hmaster0 & ~n6255;
  assign n6257 = ~n6254 & ~n6256;
  assign n6258 = controllable_hmaster1 & ~n6257;
  assign n6259 = i_hready & n5294;
  assign n6260 = controllable_ndecide & ~n5961;
  assign n6261 = controllable_ndecide & ~n6260;
  assign n6262 = ~i_hready & ~n6261;
  assign n6263 = ~n6259 & ~n6262;
  assign n6264 = ~controllable_hgrant4 & n6263;
  assign n6265 = ~n3411 & ~n6264;
  assign n6266 = ~controllable_hgrant2 & ~n6265;
  assign n6267 = ~n3410 & ~n6266;
  assign n6268 = controllable_hmaster0 & ~n6267;
  assign n6269 = ~controllable_hmaster0 & ~n6253;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = ~controllable_hmaster1 & ~n6270;
  assign n6272 = ~n6258 & ~n6271;
  assign n6273 = i_hbusreq3 & ~n6272;
  assign n6274 = i_hbusreq2 & ~n6251;
  assign n6275 = i_hbusreq4 & ~n6249;
  assign n6276 = i_hbusreq0 & ~n6249;
  assign n6277 = ~n3390 & ~n6247;
  assign n6278 = ~i_hready & ~n6277;
  assign n6279 = ~i_hready & ~n6278;
  assign n6280 = i_hlock0 & ~n6279;
  assign n6281 = ~i_hlock0 & ~n6249;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = ~i_hbusreq0 & ~n6282;
  assign n6284 = ~n6276 & ~n6283;
  assign n6285 = ~i_hbusreq4 & ~n6284;
  assign n6286 = ~n6275 & ~n6285;
  assign n6287 = ~controllable_hgrant4 & ~n6286;
  assign n6288 = ~n3916 & ~n6287;
  assign n6289 = ~i_hbusreq2 & ~n6288;
  assign n6290 = ~n6274 & ~n6289;
  assign n6291 = ~controllable_hgrant2 & ~n6290;
  assign n6292 = ~n3859 & ~n6291;
  assign n6293 = controllable_hmaster0 & ~n6292;
  assign n6294 = ~n5438 & ~n6291;
  assign n6295 = ~controllable_hmaster0 & ~n6294;
  assign n6296 = ~n6293 & ~n6295;
  assign n6297 = controllable_hmaster1 & ~n6296;
  assign n6298 = i_hbusreq2 & ~n6265;
  assign n6299 = i_hbusreq4 & ~n6263;
  assign n6300 = i_hbusreq0 & ~n6263;
  assign n6301 = ~controllable_ndecide & n5317;
  assign n6302 = ~n6137 & ~n6301;
  assign n6303 = i_hready & ~n6302;
  assign n6304 = i_hbusreq1 & ~controllable_ndecide;
  assign n6305 = ~n6260 & ~n6304;
  assign n6306 = ~i_hready & ~n6305;
  assign n6307 = ~n6303 & ~n6306;
  assign n6308 = i_hlock0 & ~n6307;
  assign n6309 = ~i_hlock0 & ~n6263;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~i_hbusreq0 & ~n6310;
  assign n6312 = ~n6300 & ~n6311;
  assign n6313 = ~i_hbusreq4 & ~n6312;
  assign n6314 = ~n6299 & ~n6313;
  assign n6315 = ~controllable_hgrant4 & n6314;
  assign n6316 = ~n3916 & ~n6315;
  assign n6317 = ~i_hbusreq2 & ~n6316;
  assign n6318 = ~n6298 & ~n6317;
  assign n6319 = ~controllable_hgrant2 & ~n6318;
  assign n6320 = ~n3859 & ~n6319;
  assign n6321 = controllable_hmaster0 & ~n6320;
  assign n6322 = ~n5382 & ~n6247;
  assign n6323 = ~i_hready & ~n6322;
  assign n6324 = ~i_hready & ~n6323;
  assign n6325 = i_hlock0 & ~n6324;
  assign n6326 = ~n6281 & ~n6325;
  assign n6327 = ~i_hbusreq0 & ~n6326;
  assign n6328 = ~n6276 & ~n6327;
  assign n6329 = ~i_hbusreq4 & ~n6328;
  assign n6330 = ~n6275 & ~n6329;
  assign n6331 = ~controllable_hgrant4 & ~n6330;
  assign n6332 = ~n5462 & ~n6331;
  assign n6333 = ~i_hbusreq2 & ~n6332;
  assign n6334 = ~n6274 & ~n6333;
  assign n6335 = ~controllable_hgrant2 & ~n6334;
  assign n6336 = ~n5461 & ~n6335;
  assign n6337 = ~controllable_hmaster0 & ~n6336;
  assign n6338 = ~n6321 & ~n6337;
  assign n6339 = ~controllable_hmaster1 & ~n6338;
  assign n6340 = ~n6297 & ~n6339;
  assign n6341 = ~i_hbusreq3 & ~n6340;
  assign n6342 = ~n6273 & ~n6341;
  assign n6343 = ~controllable_hmaster2 & ~n6342;
  assign n6344 = ~n6246 & ~n6343;
  assign n6345 = ~controllable_hgrant3 & ~n6344;
  assign n6346 = ~n5402 & ~n6345;
  assign n6347 = controllable_nhgrant0 & ~n6346;
  assign n6348 = ~n5534 & ~n6347;
  assign n6349 = ~n3281 & ~n6348;
  assign n6350 = ~n3950 & ~n6349;
  assign n6351 = ~n3378 & ~n6350;
  assign n6352 = ~n6210 & ~n6351;
  assign n6353 = n3492 & ~n6352;
  assign n6354 = ~n3631 & ~n6353;
  assign n6355 = n3485 & ~n6354;
  assign n6356 = ~n3630 & ~n6355;
  assign n6357 = ~n3476 & ~n6356;
  assign n6358 = ~n4180 & ~n5619;
  assign n6359 = ~controllable_hgrant4 & ~n6358;
  assign n6360 = ~n4015 & ~n6359;
  assign n6361 = ~controllable_hgrant2 & ~n6360;
  assign n6362 = ~n5616 & ~n6361;
  assign n6363 = ~controllable_hmaster0 & ~n6362;
  assign n6364 = ~n5626 & ~n6363;
  assign n6365 = ~controllable_hmaster1 & ~n6364;
  assign n6366 = ~n5625 & ~n6365;
  assign n6367 = i_hbusreq3 & ~n6366;
  assign n6368 = i_hbusreq2 & ~n6360;
  assign n6369 = i_hbusreq4 & ~n6358;
  assign n6370 = i_hbusreq0 & ~n6358;
  assign n6371 = ~n4195 & ~n5643;
  assign n6372 = i_hlock0 & ~n6371;
  assign n6373 = ~n4180 & ~n5643;
  assign n6374 = ~i_hlock0 & ~n6373;
  assign n6375 = ~n6372 & ~n6374;
  assign n6376 = ~i_hbusreq0 & ~n6375;
  assign n6377 = ~n6370 & ~n6376;
  assign n6378 = ~i_hbusreq4 & ~n6377;
  assign n6379 = ~n6369 & ~n6378;
  assign n6380 = ~controllable_hgrant4 & ~n6379;
  assign n6381 = ~n4064 & ~n6380;
  assign n6382 = ~i_hbusreq2 & ~n6381;
  assign n6383 = ~n6368 & ~n6382;
  assign n6384 = ~controllable_hgrant2 & ~n6383;
  assign n6385 = ~n5657 & ~n6384;
  assign n6386 = ~controllable_hmaster0 & ~n6385;
  assign n6387 = ~n5656 & ~n6386;
  assign n6388 = ~controllable_hmaster1 & ~n6387;
  assign n6389 = ~n5655 & ~n6388;
  assign n6390 = ~i_hbusreq3 & ~n6389;
  assign n6391 = ~n6367 & ~n6390;
  assign n6392 = controllable_hmaster2 & ~n6391;
  assign n6393 = ~n5752 & ~n6392;
  assign n6394 = ~controllable_hgrant3 & ~n6393;
  assign n6395 = ~n5615 & ~n6394;
  assign n6396 = controllable_nhgrant0 & ~n6395;
  assign n6397 = ~n5809 & ~n6396;
  assign n6398 = ~n3281 & ~n6397;
  assign n6399 = ~n4089 & ~n6398;
  assign n6400 = n3378 & ~n6399;
  assign n6401 = i_hready & n4178;
  assign n6402 = ~n4180 & ~n6401;
  assign n6403 = ~controllable_hgrant4 & ~n6402;
  assign n6404 = ~n4091 & ~n6403;
  assign n6405 = ~controllable_hgrant2 & ~n6404;
  assign n6406 = ~n5616 & ~n6405;
  assign n6407 = controllable_hmaster1 & ~n6406;
  assign n6408 = controllable_hmaster0 & ~n6406;
  assign n6409 = ~n4015 & ~n6403;
  assign n6410 = ~controllable_hgrant2 & ~n6409;
  assign n6411 = ~n5616 & ~n6410;
  assign n6412 = ~controllable_hmaster0 & ~n6411;
  assign n6413 = ~n6408 & ~n6412;
  assign n6414 = ~controllable_hmaster1 & ~n6413;
  assign n6415 = ~n6407 & ~n6414;
  assign n6416 = i_hbusreq3 & ~n6415;
  assign n6417 = i_hbusreq2 & ~n6404;
  assign n6418 = i_hbusreq4 & ~n6402;
  assign n6419 = i_hbusreq0 & ~n6402;
  assign n6420 = ~n4179 & ~n5641;
  assign n6421 = i_hready & ~n6420;
  assign n6422 = ~n4195 & ~n6421;
  assign n6423 = i_hlock0 & ~n6422;
  assign n6424 = ~n4179 & ~n5867;
  assign n6425 = i_hready & ~n6424;
  assign n6426 = ~n4180 & ~n6425;
  assign n6427 = ~i_hlock0 & ~n6426;
  assign n6428 = ~n6423 & ~n6427;
  assign n6429 = ~i_hbusreq0 & ~n6428;
  assign n6430 = ~n6419 & ~n6429;
  assign n6431 = ~i_hbusreq4 & ~n6430;
  assign n6432 = ~n6418 & ~n6431;
  assign n6433 = ~controllable_hgrant4 & ~n6432;
  assign n6434 = ~n5863 & ~n6433;
  assign n6435 = ~i_hbusreq2 & ~n6434;
  assign n6436 = ~n6417 & ~n6435;
  assign n6437 = ~controllable_hgrant2 & ~n6436;
  assign n6438 = ~n5862 & ~n6437;
  assign n6439 = controllable_hmaster1 & ~n6438;
  assign n6440 = controllable_hmaster0 & ~n6438;
  assign n6441 = i_hbusreq2 & ~n6409;
  assign n6442 = ~n4179 & ~n5887;
  assign n6443 = i_hready & ~n6442;
  assign n6444 = ~n4180 & ~n6443;
  assign n6445 = ~i_hlock0 & ~n6444;
  assign n6446 = ~n6423 & ~n6445;
  assign n6447 = ~i_hbusreq0 & ~n6446;
  assign n6448 = ~n6419 & ~n6447;
  assign n6449 = ~i_hbusreq4 & ~n6448;
  assign n6450 = ~n6418 & ~n6449;
  assign n6451 = ~controllable_hgrant4 & ~n6450;
  assign n6452 = ~n4064 & ~n6451;
  assign n6453 = ~i_hbusreq2 & ~n6452;
  assign n6454 = ~n6441 & ~n6453;
  assign n6455 = ~controllable_hgrant2 & ~n6454;
  assign n6456 = ~n5862 & ~n6455;
  assign n6457 = ~controllable_hmaster0 & ~n6456;
  assign n6458 = ~n6440 & ~n6457;
  assign n6459 = ~controllable_hmaster1 & ~n6458;
  assign n6460 = ~n6439 & ~n6459;
  assign n6461 = ~i_hbusreq3 & ~n6460;
  assign n6462 = ~n6416 & ~n6461;
  assign n6463 = controllable_hmaster2 & ~n6462;
  assign n6464 = ~n6248 & ~n6401;
  assign n6465 = ~controllable_hgrant4 & ~n6464;
  assign n6466 = ~n4091 & ~n6465;
  assign n6467 = ~controllable_hgrant2 & ~n6466;
  assign n6468 = ~n5616 & ~n6467;
  assign n6469 = controllable_hmaster0 & ~n6468;
  assign n6470 = ~n5686 & ~n6467;
  assign n6471 = ~controllable_hmaster0 & ~n6470;
  assign n6472 = ~n6469 & ~n6471;
  assign n6473 = controllable_hmaster1 & ~n6472;
  assign n6474 = i_hready & ~n5692;
  assign n6475 = ~n6262 & ~n6474;
  assign n6476 = ~controllable_hgrant4 & n6475;
  assign n6477 = ~n4091 & ~n6476;
  assign n6478 = ~controllable_hgrant2 & ~n6477;
  assign n6479 = ~n5616 & ~n6478;
  assign n6480 = controllable_hmaster0 & ~n6479;
  assign n6481 = ~controllable_hmaster0 & ~n6468;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = ~controllable_hmaster1 & ~n6482;
  assign n6484 = ~n6473 & ~n6483;
  assign n6485 = i_hbusreq3 & ~n6484;
  assign n6486 = i_hbusreq2 & ~n6466;
  assign n6487 = i_hbusreq4 & ~n6464;
  assign n6488 = i_hbusreq0 & ~n6464;
  assign n6489 = ~n6278 & ~n6421;
  assign n6490 = i_hlock0 & ~n6489;
  assign n6491 = ~n6248 & ~n6443;
  assign n6492 = ~i_hlock0 & ~n6491;
  assign n6493 = ~n6490 & ~n6492;
  assign n6494 = ~i_hbusreq0 & ~n6493;
  assign n6495 = ~n6488 & ~n6494;
  assign n6496 = ~i_hbusreq4 & ~n6495;
  assign n6497 = ~n6487 & ~n6496;
  assign n6498 = ~controllable_hgrant4 & ~n6497;
  assign n6499 = ~n5863 & ~n6498;
  assign n6500 = ~i_hbusreq2 & ~n6499;
  assign n6501 = ~n6486 & ~n6500;
  assign n6502 = ~controllable_hgrant2 & ~n6501;
  assign n6503 = ~n5862 & ~n6502;
  assign n6504 = controllable_hmaster0 & ~n6503;
  assign n6505 = ~n5950 & ~n6502;
  assign n6506 = ~controllable_hmaster0 & ~n6505;
  assign n6507 = ~n6504 & ~n6506;
  assign n6508 = controllable_hmaster1 & ~n6507;
  assign n6509 = i_hbusreq2 & ~n6477;
  assign n6510 = i_hbusreq4 & ~n6475;
  assign n6511 = i_hbusreq0 & ~n6475;
  assign n6512 = controllable_ndecide & ~n5692;
  assign n6513 = ~controllable_ndecide & n5730;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = i_hready & ~n6514;
  assign n6516 = ~n6306 & ~n6515;
  assign n6517 = i_hlock0 & ~n6516;
  assign n6518 = ~controllable_ndecide & ~n5963;
  assign n6519 = ~n6512 & ~n6518;
  assign n6520 = i_hready & ~n6519;
  assign n6521 = ~n6262 & ~n6520;
  assign n6522 = ~i_hlock0 & ~n6521;
  assign n6523 = ~n6517 & ~n6522;
  assign n6524 = ~i_hbusreq0 & ~n6523;
  assign n6525 = ~n6511 & ~n6524;
  assign n6526 = ~i_hbusreq4 & ~n6525;
  assign n6527 = ~n6510 & ~n6526;
  assign n6528 = ~controllable_hgrant4 & n6527;
  assign n6529 = ~n5863 & ~n6528;
  assign n6530 = ~i_hbusreq2 & ~n6529;
  assign n6531 = ~n6509 & ~n6530;
  assign n6532 = ~controllable_hgrant2 & ~n6531;
  assign n6533 = ~n5862 & ~n6532;
  assign n6534 = controllable_hmaster0 & ~n6533;
  assign n6535 = ~n6323 & ~n6421;
  assign n6536 = i_hlock0 & ~n6535;
  assign n6537 = ~n6492 & ~n6536;
  assign n6538 = ~i_hbusreq0 & ~n6537;
  assign n6539 = ~n6488 & ~n6538;
  assign n6540 = ~i_hbusreq4 & ~n6539;
  assign n6541 = ~n6487 & ~n6540;
  assign n6542 = ~controllable_hgrant4 & ~n6541;
  assign n6543 = ~n5982 & ~n6542;
  assign n6544 = ~i_hbusreq2 & ~n6543;
  assign n6545 = ~n6486 & ~n6544;
  assign n6546 = ~controllable_hgrant2 & ~n6545;
  assign n6547 = ~n5981 & ~n6546;
  assign n6548 = ~controllable_hmaster0 & ~n6547;
  assign n6549 = ~n6534 & ~n6548;
  assign n6550 = ~controllable_hmaster1 & ~n6549;
  assign n6551 = ~n6508 & ~n6550;
  assign n6552 = ~i_hbusreq3 & ~n6551;
  assign n6553 = ~n6485 & ~n6552;
  assign n6554 = ~controllable_hmaster2 & ~n6553;
  assign n6555 = ~n6463 & ~n6554;
  assign n6556 = ~controllable_hgrant3 & ~n6555;
  assign n6557 = ~n5861 & ~n6556;
  assign n6558 = controllable_nhgrant0 & ~n6557;
  assign n6559 = ~n6082 & ~n6558;
  assign n6560 = ~n3281 & ~n6559;
  assign n6561 = ~n4089 & ~n6560;
  assign n6562 = ~n3378 & ~n6561;
  assign n6563 = ~n6400 & ~n6562;
  assign n6564 = n3492 & ~n6563;
  assign n6565 = ~n3631 & ~n6564;
  assign n6566 = n3485 & ~n6565;
  assign n6567 = ~n3630 & ~n6566;
  assign n6568 = n3476 & ~n6567;
  assign n6569 = ~n6357 & ~n6568;
  assign n6570 = n3374 & ~n6569;
  assign n6571 = ~n6202 & ~n6570;
  assign n6572 = ~n3655 & ~n6571;
  assign n6573 = ~n6096 & ~n6572;
  assign n6574 = n3652 & ~n6573;
  assign n6575 = ~n4333 & ~n5043;
  assign n6576 = controllable_hmaster1 & ~n6575;
  assign n6577 = controllable_hmaster0 & ~n6575;
  assign n6578 = ~n3729 & ~n6577;
  assign n6579 = ~controllable_hmaster1 & ~n6578;
  assign n6580 = ~n6576 & ~n6579;
  assign n6581 = i_hbusreq3 & ~n6580;
  assign n6582 = ~n4340 & ~n5068;
  assign n6583 = controllable_hmaster1 & ~n6582;
  assign n6584 = controllable_hmaster0 & ~n6582;
  assign n6585 = ~n3767 & ~n6584;
  assign n6586 = ~controllable_hmaster1 & ~n6585;
  assign n6587 = ~n6583 & ~n6586;
  assign n6588 = ~i_hbusreq3 & ~n6587;
  assign n6589 = ~n6581 & ~n6588;
  assign n6590 = controllable_hmaster2 & ~n6589;
  assign n6591 = ~controllable_hgrant4 & ~n5210;
  assign n6592 = ~n4921 & ~n6591;
  assign n6593 = i_hlock2 & ~n6592;
  assign n6594 = ~controllable_hgrant4 & ~n5216;
  assign n6595 = ~n4950 & ~n6594;
  assign n6596 = ~i_hlock2 & ~n6595;
  assign n6597 = ~n6593 & ~n6596;
  assign n6598 = controllable_hgrant2 & ~n6597;
  assign n6599 = ~n5083 & ~n6598;
  assign n6600 = ~controllable_hmaster0 & ~n6599;
  assign n6601 = ~n5078 & ~n6600;
  assign n6602 = controllable_hmaster1 & ~n6601;
  assign n6603 = ~n5105 & ~n6602;
  assign n6604 = i_hlock3 & ~n6603;
  assign n6605 = ~n5108 & ~n6600;
  assign n6606 = controllable_hmaster1 & ~n6605;
  assign n6607 = ~n5105 & ~n6606;
  assign n6608 = ~i_hlock3 & ~n6607;
  assign n6609 = ~n6604 & ~n6608;
  assign n6610 = i_hbusreq3 & ~n6609;
  assign n6611 = i_hbusreq2 & ~n6597;
  assign n6612 = i_hbusreq4 & ~n5210;
  assign n6613 = i_hbusreq0 & ~n5210;
  assign n6614 = ~n3418 & ~n3740;
  assign n6615 = i_hready & ~n6614;
  assign n6616 = ~n3418 & ~n3676;
  assign n6617 = ~i_hready & ~n6616;
  assign n6618 = ~n6615 & ~n6617;
  assign n6619 = ~i_hbusreq0 & ~n6618;
  assign n6620 = ~n6613 & ~n6619;
  assign n6621 = ~i_hbusreq4 & ~n6620;
  assign n6622 = ~n6612 & ~n6621;
  assign n6623 = ~controllable_hgrant4 & ~n6622;
  assign n6624 = ~n4970 & ~n6623;
  assign n6625 = i_hlock2 & ~n6624;
  assign n6626 = i_hbusreq4 & ~n5216;
  assign n6627 = i_hbusreq0 & ~n5216;
  assign n6628 = ~n3418 & ~n3750;
  assign n6629 = i_hready & ~n6628;
  assign n6630 = ~n3418 & ~n3685;
  assign n6631 = ~i_hready & ~n6630;
  assign n6632 = ~n6629 & ~n6631;
  assign n6633 = ~i_hbusreq0 & ~n6632;
  assign n6634 = ~n6627 & ~n6633;
  assign n6635 = ~i_hbusreq4 & ~n6634;
  assign n6636 = ~n6626 & ~n6635;
  assign n6637 = ~controllable_hgrant4 & ~n6636;
  assign n6638 = ~n5017 & ~n6637;
  assign n6639 = ~i_hlock2 & ~n6638;
  assign n6640 = ~n6625 & ~n6639;
  assign n6641 = ~i_hbusreq2 & ~n6640;
  assign n6642 = ~n6611 & ~n6641;
  assign n6643 = controllable_hgrant2 & ~n6642;
  assign n6644 = ~n5123 & ~n6643;
  assign n6645 = ~controllable_hmaster0 & ~n6644;
  assign n6646 = ~n5115 & ~n6645;
  assign n6647 = controllable_hmaster1 & ~n6646;
  assign n6648 = ~n5150 & ~n6647;
  assign n6649 = i_hlock3 & ~n6648;
  assign n6650 = ~n5153 & ~n6645;
  assign n6651 = controllable_hmaster1 & ~n6650;
  assign n6652 = ~n5150 & ~n6651;
  assign n6653 = ~i_hlock3 & ~n6652;
  assign n6654 = ~n6649 & ~n6653;
  assign n6655 = ~i_hbusreq3 & ~n6654;
  assign n6656 = ~n6610 & ~n6655;
  assign n6657 = ~controllable_hmaster2 & ~n6656;
  assign n6658 = ~n6590 & ~n6657;
  assign n6659 = ~controllable_hgrant3 & ~n6658;
  assign n6660 = ~n5037 & ~n6659;
  assign n6661 = controllable_nhgrant0 & ~n6660;
  assign n6662 = ~n5245 & ~n6661;
  assign n6663 = ~n3281 & ~n6662;
  assign n6664 = ~n3783 & ~n6663;
  assign n6665 = ~n3378 & ~n6664;
  assign n6666 = ~n4911 & ~n6665;
  assign n6667 = n3492 & ~n6666;
  assign n6668 = ~n3631 & ~n6667;
  assign n6669 = n3485 & ~n6668;
  assign n6670 = ~n3630 & ~n6669;
  assign n6671 = ~n3374 & ~n6670;
  assign n6672 = ~n4366 & ~n5338;
  assign n6673 = ~controllable_hgrant3 & ~n6672;
  assign n6674 = ~n5287 & ~n6673;
  assign n6675 = controllable_nhgrant0 & ~n6674;
  assign n6676 = ~n5363 & ~n6675;
  assign n6677 = ~n3281 & ~n6676;
  assign n6678 = ~n3950 & ~n6677;
  assign n6679 = n3378 & ~n6678;
  assign n6680 = ~n3499 & ~n4333;
  assign n6681 = controllable_hmaster1 & ~n6680;
  assign n6682 = controllable_hmaster0 & ~n6680;
  assign n6683 = ~n4335 & ~n6682;
  assign n6684 = ~controllable_hmaster1 & ~n6683;
  assign n6685 = ~n6681 & ~n6684;
  assign n6686 = i_hbusreq3 & ~n6685;
  assign n6687 = ~n4340 & ~n5414;
  assign n6688 = controllable_hmaster1 & ~n6687;
  assign n6689 = controllable_hmaster0 & ~n6687;
  assign n6690 = ~n4342 & ~n6689;
  assign n6691 = ~controllable_hmaster1 & ~n6690;
  assign n6692 = ~n6688 & ~n6691;
  assign n6693 = ~i_hbusreq3 & ~n6692;
  assign n6694 = ~n6686 & ~n6693;
  assign n6695 = controllable_hmaster2 & ~n6694;
  assign n6696 = controllable_hmaster0 & ~n3907;
  assign n6697 = controllable_hgrant2 & ~n5042;
  assign n6698 = ~n3908 & ~n6697;
  assign n6699 = ~controllable_hmaster0 & ~n6698;
  assign n6700 = ~n6696 & ~n6699;
  assign n6701 = controllable_hmaster1 & ~n6700;
  assign n6702 = ~n4333 & ~n5431;
  assign n6703 = controllable_hmaster0 & ~n6702;
  assign n6704 = ~controllable_hmaster0 & ~n3907;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = ~controllable_hmaster1 & ~n6705;
  assign n6707 = ~n6701 & ~n6706;
  assign n6708 = i_hbusreq3 & ~n6707;
  assign n6709 = controllable_hmaster0 & ~n3932;
  assign n6710 = controllable_hgrant2 & ~n5067;
  assign n6711 = ~n3933 & ~n6710;
  assign n6712 = ~controllable_hmaster0 & ~n6711;
  assign n6713 = ~n6709 & ~n6712;
  assign n6714 = controllable_hmaster1 & ~n6713;
  assign n6715 = ~n4340 & ~n5458;
  assign n6716 = controllable_hmaster0 & ~n6715;
  assign n6717 = ~controllable_hmaster0 & ~n5475;
  assign n6718 = ~n6716 & ~n6717;
  assign n6719 = ~controllable_hmaster1 & ~n6718;
  assign n6720 = ~n6714 & ~n6719;
  assign n6721 = ~i_hbusreq3 & ~n6720;
  assign n6722 = ~n6708 & ~n6721;
  assign n6723 = ~controllable_hmaster2 & ~n6722;
  assign n6724 = ~n6695 & ~n6723;
  assign n6725 = ~controllable_hgrant3 & ~n6724;
  assign n6726 = ~n5402 & ~n6725;
  assign n6727 = controllable_nhgrant0 & ~n6726;
  assign n6728 = ~n5534 & ~n6727;
  assign n6729 = ~n3281 & ~n6728;
  assign n6730 = ~n3950 & ~n6729;
  assign n6731 = ~n3378 & ~n6730;
  assign n6732 = ~n6679 & ~n6731;
  assign n6733 = n3492 & ~n6732;
  assign n6734 = ~n3631 & ~n6733;
  assign n6735 = n3485 & ~n6734;
  assign n6736 = ~n3630 & ~n6735;
  assign n6737 = ~n3476 & ~n6736;
  assign n6738 = controllable_hgrant2 & ~n5761;
  assign n6739 = ~n5628 & ~n6738;
  assign n6740 = ~controllable_hmaster0 & ~n6739;
  assign n6741 = ~n5626 & ~n6740;
  assign n6742 = ~controllable_hmaster1 & ~n6741;
  assign n6743 = ~n5625 & ~n6742;
  assign n6744 = i_hbusreq3 & ~n6743;
  assign n6745 = controllable_hgrant2 & ~n5784;
  assign n6746 = ~n5671 & ~n6745;
  assign n6747 = ~controllable_hmaster0 & ~n6746;
  assign n6748 = ~n5656 & ~n6747;
  assign n6749 = ~controllable_hmaster1 & ~n6748;
  assign n6750 = ~n5655 & ~n6749;
  assign n6751 = ~i_hbusreq3 & ~n6750;
  assign n6752 = ~n6744 & ~n6751;
  assign n6753 = controllable_hmaster2 & ~n6752;
  assign n6754 = ~n5752 & ~n6753;
  assign n6755 = ~controllable_hgrant3 & ~n6754;
  assign n6756 = ~n5615 & ~n6755;
  assign n6757 = controllable_nhgrant0 & ~n6756;
  assign n6758 = ~n5809 & ~n6757;
  assign n6759 = ~n3281 & ~n6758;
  assign n6760 = ~n4089 & ~n6759;
  assign n6761 = n3378 & ~n6760;
  assign n6762 = controllable_hgrant2 & ~n6010;
  assign n6763 = ~n5623 & ~n6762;
  assign n6764 = controllable_hmaster1 & ~n6763;
  assign n6765 = controllable_hmaster0 & ~n6763;
  assign n6766 = ~n5628 & ~n6762;
  assign n6767 = ~controllable_hmaster0 & ~n6766;
  assign n6768 = ~n6765 & ~n6767;
  assign n6769 = ~controllable_hmaster1 & ~n6768;
  assign n6770 = ~n6764 & ~n6769;
  assign n6771 = i_hbusreq3 & ~n6770;
  assign n6772 = controllable_hgrant2 & ~n6030;
  assign n6773 = ~n5881 & ~n6772;
  assign n6774 = controllable_hmaster1 & ~n6773;
  assign n6775 = controllable_hmaster0 & ~n6773;
  assign n6776 = ~n5901 & ~n6772;
  assign n6777 = ~controllable_hmaster0 & ~n6776;
  assign n6778 = ~n6775 & ~n6777;
  assign n6779 = ~controllable_hmaster1 & ~n6778;
  assign n6780 = ~n6774 & ~n6779;
  assign n6781 = ~i_hbusreq3 & ~n6780;
  assign n6782 = ~n6771 & ~n6781;
  assign n6783 = controllable_hmaster2 & ~n6782;
  assign n6784 = ~n5913 & ~n6762;
  assign n6785 = controllable_hmaster0 & ~n6784;
  assign n6786 = controllable_hgrant2 & ~n6041;
  assign n6787 = ~n5913 & ~n6786;
  assign n6788 = ~controllable_hmaster0 & ~n6787;
  assign n6789 = ~n6785 & ~n6788;
  assign n6790 = controllable_hmaster1 & ~n6789;
  assign n6791 = ~n5923 & ~n6762;
  assign n6792 = controllable_hmaster0 & ~n6791;
  assign n6793 = ~controllable_hmaster0 & ~n6784;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = ~controllable_hmaster1 & ~n6794;
  assign n6796 = ~n6790 & ~n6795;
  assign n6797 = i_hbusreq3 & ~n6796;
  assign n6798 = ~n5947 & ~n6772;
  assign n6799 = controllable_hmaster0 & ~n6798;
  assign n6800 = ~n4053 & ~n5038;
  assign n6801 = i_hready & ~n6800;
  assign n6802 = ~n5055 & ~n6801;
  assign n6803 = i_hlock0 & ~n6802;
  assign n6804 = ~n6060 & ~n6803;
  assign n6805 = ~i_hbusreq0 & ~n6804;
  assign n6806 = ~n6053 & ~n6805;
  assign n6807 = ~i_hbusreq4 & ~n6806;
  assign n6808 = ~n6052 & ~n6807;
  assign n6809 = ~controllable_hgrant4 & ~n6808;
  assign n6810 = ~n3916 & ~n6809;
  assign n6811 = ~i_hbusreq2 & ~n6810;
  assign n6812 = ~n6051 & ~n6811;
  assign n6813 = controllable_hgrant2 & ~n6812;
  assign n6814 = ~n5947 & ~n6813;
  assign n6815 = ~controllable_hmaster0 & ~n6814;
  assign n6816 = ~n6799 & ~n6815;
  assign n6817 = controllable_hmaster1 & ~n6816;
  assign n6818 = ~n5978 & ~n6772;
  assign n6819 = controllable_hmaster0 & ~n6818;
  assign n6820 = ~n5464 & ~n6018;
  assign n6821 = i_hlock0 & ~n6820;
  assign n6822 = ~n6021 & ~n6821;
  assign n6823 = ~i_hbusreq0 & ~n6822;
  assign n6824 = ~n6016 & ~n6823;
  assign n6825 = ~i_hbusreq4 & ~n6824;
  assign n6826 = ~n6015 & ~n6825;
  assign n6827 = ~controllable_hgrant4 & ~n6826;
  assign n6828 = ~n5462 & ~n6827;
  assign n6829 = ~i_hbusreq2 & ~n6828;
  assign n6830 = ~n6014 & ~n6829;
  assign n6831 = controllable_hgrant2 & ~n6830;
  assign n6832 = ~n5994 & ~n6831;
  assign n6833 = ~controllable_hmaster0 & ~n6832;
  assign n6834 = ~n6819 & ~n6833;
  assign n6835 = ~controllable_hmaster1 & ~n6834;
  assign n6836 = ~n6817 & ~n6835;
  assign n6837 = ~i_hbusreq3 & ~n6836;
  assign n6838 = ~n6797 & ~n6837;
  assign n6839 = ~controllable_hmaster2 & ~n6838;
  assign n6840 = ~n6783 & ~n6839;
  assign n6841 = ~controllable_hgrant3 & ~n6840;
  assign n6842 = ~n5861 & ~n6841;
  assign n6843 = controllable_nhgrant0 & ~n6842;
  assign n6844 = ~n6082 & ~n6843;
  assign n6845 = ~n3281 & ~n6844;
  assign n6846 = ~n4089 & ~n6845;
  assign n6847 = ~n3378 & ~n6846;
  assign n6848 = ~n6761 & ~n6847;
  assign n6849 = n3492 & ~n6848;
  assign n6850 = ~n3631 & ~n6849;
  assign n6851 = n3485 & ~n6850;
  assign n6852 = ~n3630 & ~n6851;
  assign n6853 = n3476 & ~n6852;
  assign n6854 = ~n6737 & ~n6853;
  assign n6855 = n3374 & ~n6854;
  assign n6856 = ~n6671 & ~n6855;
  assign n6857 = n3655 & ~n6856;
  assign n6858 = ~n4333 & ~n6102;
  assign n6859 = controllable_hmaster1 & ~n6858;
  assign n6860 = controllable_hmaster0 & ~n6858;
  assign n6861 = ~n3729 & ~n6860;
  assign n6862 = ~controllable_hmaster1 & ~n6861;
  assign n6863 = ~n6859 & ~n6862;
  assign n6864 = i_hbusreq3 & ~n6863;
  assign n6865 = ~n4340 & ~n6127;
  assign n6866 = controllable_hmaster1 & ~n6865;
  assign n6867 = controllable_hmaster0 & ~n6865;
  assign n6868 = ~n3767 & ~n6867;
  assign n6869 = ~controllable_hmaster1 & ~n6868;
  assign n6870 = ~n6866 & ~n6869;
  assign n6871 = ~i_hbusreq3 & ~n6870;
  assign n6872 = ~n6864 & ~n6871;
  assign n6873 = controllable_hmaster2 & ~n6872;
  assign n6874 = ~n6151 & ~n6602;
  assign n6875 = i_hlock3 & ~n6874;
  assign n6876 = ~n6151 & ~n6606;
  assign n6877 = ~i_hlock3 & ~n6876;
  assign n6878 = ~n6875 & ~n6877;
  assign n6879 = i_hbusreq3 & ~n6878;
  assign n6880 = ~n6180 & ~n6647;
  assign n6881 = i_hlock3 & ~n6880;
  assign n6882 = ~n6180 & ~n6651;
  assign n6883 = ~i_hlock3 & ~n6882;
  assign n6884 = ~n6881 & ~n6883;
  assign n6885 = ~i_hbusreq3 & ~n6884;
  assign n6886 = ~n6879 & ~n6885;
  assign n6887 = ~controllable_hmaster2 & ~n6886;
  assign n6888 = ~n6873 & ~n6887;
  assign n6889 = ~controllable_hgrant3 & ~n6888;
  assign n6890 = ~n5037 & ~n6889;
  assign n6891 = controllable_nhgrant0 & ~n6890;
  assign n6892 = ~n5245 & ~n6891;
  assign n6893 = ~n3281 & ~n6892;
  assign n6894 = ~n3783 & ~n6893;
  assign n6895 = ~n3378 & ~n6894;
  assign n6896 = ~n4911 & ~n6895;
  assign n6897 = n3492 & ~n6896;
  assign n6898 = ~n3631 & ~n6897;
  assign n6899 = n3485 & ~n6898;
  assign n6900 = ~n3630 & ~n6899;
  assign n6901 = ~n3374 & ~n6900;
  assign n6902 = ~n4466 & ~n5338;
  assign n6903 = ~controllable_hgrant3 & ~n6902;
  assign n6904 = ~n5287 & ~n6903;
  assign n6905 = controllable_nhgrant0 & ~n6904;
  assign n6906 = ~n5363 & ~n6905;
  assign n6907 = ~n3281 & ~n6906;
  assign n6908 = ~n3950 & ~n6907;
  assign n6909 = n3378 & ~n6908;
  assign n6910 = ~n4333 & ~n6214;
  assign n6911 = controllable_hmaster1 & ~n6910;
  assign n6912 = controllable_hmaster0 & ~n6910;
  assign n6913 = ~n4436 & ~n6912;
  assign n6914 = ~controllable_hmaster1 & ~n6913;
  assign n6915 = ~n6911 & ~n6914;
  assign n6916 = i_hbusreq3 & ~n6915;
  assign n6917 = ~n4340 & ~n6237;
  assign n6918 = controllable_hmaster1 & ~n6917;
  assign n6919 = controllable_hmaster0 & ~n6917;
  assign n6920 = ~n4442 & ~n6919;
  assign n6921 = ~controllable_hmaster1 & ~n6920;
  assign n6922 = ~n6918 & ~n6921;
  assign n6923 = ~i_hbusreq3 & ~n6922;
  assign n6924 = ~n6916 & ~n6923;
  assign n6925 = controllable_hmaster2 & ~n6924;
  assign n6926 = ~n4333 & ~n6252;
  assign n6927 = controllable_hmaster0 & ~n6926;
  assign n6928 = ~n6252 & ~n6697;
  assign n6929 = ~controllable_hmaster0 & ~n6928;
  assign n6930 = ~n6927 & ~n6929;
  assign n6931 = controllable_hmaster1 & ~n6930;
  assign n6932 = ~n4333 & ~n6266;
  assign n6933 = controllable_hmaster0 & ~n6932;
  assign n6934 = ~controllable_hmaster0 & ~n6926;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = ~controllable_hmaster1 & ~n6935;
  assign n6937 = ~n6931 & ~n6936;
  assign n6938 = i_hbusreq3 & ~n6937;
  assign n6939 = ~n4340 & ~n6291;
  assign n6940 = controllable_hmaster0 & ~n6939;
  assign n6941 = ~n6291 & ~n6710;
  assign n6942 = ~controllable_hmaster0 & ~n6941;
  assign n6943 = ~n6940 & ~n6942;
  assign n6944 = controllable_hmaster1 & ~n6943;
  assign n6945 = ~n4340 & ~n6319;
  assign n6946 = controllable_hmaster0 & ~n6945;
  assign n6947 = controllable_hgrant2 & ~n5475;
  assign n6948 = ~n6335 & ~n6947;
  assign n6949 = ~controllable_hmaster0 & ~n6948;
  assign n6950 = ~n6946 & ~n6949;
  assign n6951 = ~controllable_hmaster1 & ~n6950;
  assign n6952 = ~n6944 & ~n6951;
  assign n6953 = ~i_hbusreq3 & ~n6952;
  assign n6954 = ~n6938 & ~n6953;
  assign n6955 = ~controllable_hmaster2 & ~n6954;
  assign n6956 = ~n6925 & ~n6955;
  assign n6957 = ~controllable_hgrant3 & ~n6956;
  assign n6958 = ~n5402 & ~n6957;
  assign n6959 = controllable_nhgrant0 & ~n6958;
  assign n6960 = ~n5534 & ~n6959;
  assign n6961 = ~n3281 & ~n6960;
  assign n6962 = ~n3950 & ~n6961;
  assign n6963 = ~n3378 & ~n6962;
  assign n6964 = ~n6909 & ~n6963;
  assign n6965 = n3492 & ~n6964;
  assign n6966 = ~n3631 & ~n6965;
  assign n6967 = n3485 & ~n6966;
  assign n6968 = ~n3630 & ~n6967;
  assign n6969 = ~n3476 & ~n6968;
  assign n6970 = ~n6361 & ~n6738;
  assign n6971 = ~controllable_hmaster0 & ~n6970;
  assign n6972 = ~n5626 & ~n6971;
  assign n6973 = ~controllable_hmaster1 & ~n6972;
  assign n6974 = ~n5625 & ~n6973;
  assign n6975 = i_hbusreq3 & ~n6974;
  assign n6976 = ~n6384 & ~n6745;
  assign n6977 = ~controllable_hmaster0 & ~n6976;
  assign n6978 = ~n5656 & ~n6977;
  assign n6979 = ~controllable_hmaster1 & ~n6978;
  assign n6980 = ~n5655 & ~n6979;
  assign n6981 = ~i_hbusreq3 & ~n6980;
  assign n6982 = ~n6975 & ~n6981;
  assign n6983 = controllable_hmaster2 & ~n6982;
  assign n6984 = ~n5752 & ~n6983;
  assign n6985 = ~controllable_hgrant3 & ~n6984;
  assign n6986 = ~n5615 & ~n6985;
  assign n6987 = controllable_nhgrant0 & ~n6986;
  assign n6988 = ~n5809 & ~n6987;
  assign n6989 = ~n3281 & ~n6988;
  assign n6990 = ~n4089 & ~n6989;
  assign n6991 = n3378 & ~n6990;
  assign n6992 = ~n6405 & ~n6762;
  assign n6993 = controllable_hmaster1 & ~n6992;
  assign n6994 = controllable_hmaster0 & ~n6992;
  assign n6995 = ~n6410 & ~n6762;
  assign n6996 = ~controllable_hmaster0 & ~n6995;
  assign n6997 = ~n6994 & ~n6996;
  assign n6998 = ~controllable_hmaster1 & ~n6997;
  assign n6999 = ~n6993 & ~n6998;
  assign n7000 = i_hbusreq3 & ~n6999;
  assign n7001 = ~n6437 & ~n6772;
  assign n7002 = controllable_hmaster1 & ~n7001;
  assign n7003 = controllable_hmaster0 & ~n7001;
  assign n7004 = ~n6455 & ~n6772;
  assign n7005 = ~controllable_hmaster0 & ~n7004;
  assign n7006 = ~n7003 & ~n7005;
  assign n7007 = ~controllable_hmaster1 & ~n7006;
  assign n7008 = ~n7002 & ~n7007;
  assign n7009 = ~i_hbusreq3 & ~n7008;
  assign n7010 = ~n7000 & ~n7009;
  assign n7011 = controllable_hmaster2 & ~n7010;
  assign n7012 = ~n6467 & ~n6762;
  assign n7013 = controllable_hmaster0 & ~n7012;
  assign n7014 = ~n6467 & ~n6786;
  assign n7015 = ~controllable_hmaster0 & ~n7014;
  assign n7016 = ~n7013 & ~n7015;
  assign n7017 = controllable_hmaster1 & ~n7016;
  assign n7018 = ~n6478 & ~n6762;
  assign n7019 = controllable_hmaster0 & ~n7018;
  assign n7020 = ~controllable_hmaster0 & ~n7012;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = ~controllable_hmaster1 & ~n7021;
  assign n7023 = ~n7017 & ~n7022;
  assign n7024 = i_hbusreq3 & ~n7023;
  assign n7025 = ~n6502 & ~n6772;
  assign n7026 = controllable_hmaster0 & ~n7025;
  assign n7027 = ~n6502 & ~n6813;
  assign n7028 = ~controllable_hmaster0 & ~n7027;
  assign n7029 = ~n7026 & ~n7028;
  assign n7030 = controllable_hmaster1 & ~n7029;
  assign n7031 = ~n6532 & ~n6772;
  assign n7032 = controllable_hmaster0 & ~n7031;
  assign n7033 = ~n6546 & ~n6831;
  assign n7034 = ~controllable_hmaster0 & ~n7033;
  assign n7035 = ~n7032 & ~n7034;
  assign n7036 = ~controllable_hmaster1 & ~n7035;
  assign n7037 = ~n7030 & ~n7036;
  assign n7038 = ~i_hbusreq3 & ~n7037;
  assign n7039 = ~n7024 & ~n7038;
  assign n7040 = ~controllable_hmaster2 & ~n7039;
  assign n7041 = ~n7011 & ~n7040;
  assign n7042 = ~controllable_hgrant3 & ~n7041;
  assign n7043 = ~n5861 & ~n7042;
  assign n7044 = controllable_nhgrant0 & ~n7043;
  assign n7045 = ~n6082 & ~n7044;
  assign n7046 = ~n3281 & ~n7045;
  assign n7047 = ~n4089 & ~n7046;
  assign n7048 = ~n3378 & ~n7047;
  assign n7049 = ~n6991 & ~n7048;
  assign n7050 = n3492 & ~n7049;
  assign n7051 = ~n3631 & ~n7050;
  assign n7052 = n3485 & ~n7051;
  assign n7053 = ~n3630 & ~n7052;
  assign n7054 = n3476 & ~n7053;
  assign n7055 = ~n6969 & ~n7054;
  assign n7056 = n3374 & ~n7055;
  assign n7057 = ~n6901 & ~n7056;
  assign n7058 = ~n3655 & ~n7057;
  assign n7059 = ~n6857 & ~n7058;
  assign n7060 = ~n3652 & ~n7059;
  assign n7061 = ~n6574 & ~n7060;
  assign n7062 = ~n3368 & ~n7061;
  assign n7063 = controllable_hmaster1 & ~n5259;
  assign n7064 = controllable_hmaster0 & ~n5260;
  assign n7065 = ~controllable_hmaster1 & ~n7064;
  assign n7066 = ~n7063 & ~n7065;
  assign n7067 = i_hbusreq3 & ~n7066;
  assign n7068 = controllable_hmaster1 & ~n5276;
  assign n7069 = controllable_hmaster0 & ~n5277;
  assign n7070 = ~controllable_hmaster1 & ~n7069;
  assign n7071 = ~n7068 & ~n7070;
  assign n7072 = ~i_hbusreq3 & ~n7071;
  assign n7073 = ~n7067 & ~n7072;
  assign n7074 = controllable_hmaster2 & ~n7073;
  assign n7075 = controllable_hmaster2 & ~n7074;
  assign n7076 = ~controllable_hgrant3 & ~n7075;
  assign n7077 = ~n3409 & ~n7076;
  assign n7078 = controllable_nhgrant0 & ~n7077;
  assign n7079 = ~n3466 & ~n7078;
  assign n7080 = ~n3281 & ~n7079;
  assign n7081 = ~n3281 & ~n7080;
  assign n7082 = n3378 & ~n7081;
  assign n7083 = controllable_hmaster0 & ~n4913;
  assign n7084 = ~controllable_hmaster1 & ~n7083;
  assign n7085 = ~n4912 & ~n7084;
  assign n7086 = ~i_hbusreq3 & ~n7085;
  assign n7087 = ~n3386 & ~n7086;
  assign n7088 = controllable_hmaster2 & ~n7087;
  assign n7089 = controllable_hmaster2 & ~n7088;
  assign n7090 = controllable_hgrant3 & ~n7089;
  assign n7091 = controllable_hmaster0 & ~n5046;
  assign n7092 = ~controllable_hmaster1 & ~n7091;
  assign n7093 = ~n5045 & ~n7092;
  assign n7094 = i_hbusreq3 & ~n7093;
  assign n7095 = controllable_hmaster0 & ~n5071;
  assign n7096 = ~controllable_hmaster1 & ~n7095;
  assign n7097 = ~n5070 & ~n7096;
  assign n7098 = ~i_hbusreq3 & ~n7097;
  assign n7099 = ~n7094 & ~n7098;
  assign n7100 = controllable_hmaster2 & ~n7099;
  assign n7101 = controllable_hmaster2 & ~n7100;
  assign n7102 = ~controllable_hgrant3 & ~n7101;
  assign n7103 = ~n7090 & ~n7102;
  assign n7104 = controllable_nhgrant0 & ~n7103;
  assign n7105 = controllable_hmaster0 & ~n5191;
  assign n7106 = ~controllable_hmaster1 & ~n7105;
  assign n7107 = ~n5190 & ~n7106;
  assign n7108 = i_hbusreq3 & ~n7107;
  assign n7109 = controllable_hmaster0 & ~n5197;
  assign n7110 = ~controllable_hmaster1 & ~n7109;
  assign n7111 = ~n5196 & ~n7110;
  assign n7112 = ~i_hbusreq3 & ~n7111;
  assign n7113 = ~n7108 & ~n7112;
  assign n7114 = controllable_hmaster2 & ~n7113;
  assign n7115 = controllable_hmaster2 & ~n7114;
  assign n7116 = ~controllable_hgrant3 & ~n7115;
  assign n7117 = ~n7090 & ~n7116;
  assign n7118 = ~controllable_nhgrant0 & ~n7117;
  assign n7119 = ~n7104 & ~n7118;
  assign n7120 = ~n3281 & ~n7119;
  assign n7121 = ~n3281 & ~n7120;
  assign n7122 = ~n3378 & ~n7121;
  assign n7123 = ~n7082 & ~n7122;
  assign n7124 = n3492 & ~n7123;
  assign n7125 = n3492 & ~n7124;
  assign n7126 = n3485 & ~n7125;
  assign n7127 = n3485 & ~n7126;
  assign n7128 = ~n3374 & ~n7127;
  assign n7129 = ~n3401 & ~n4553;
  assign n7130 = ~controllable_hmaster1 & ~n7129;
  assign n7131 = ~n3400 & ~n7130;
  assign n7132 = ~i_hbusreq3 & ~n7131;
  assign n7133 = ~n3951 & ~n7132;
  assign n7134 = controllable_hmaster2 & ~n7133;
  assign n7135 = ~n5285 & ~n7134;
  assign n7136 = controllable_hgrant3 & ~n7135;
  assign n7137 = ~n3854 & ~n5260;
  assign n7138 = ~controllable_hmaster1 & ~n7137;
  assign n7139 = ~n7063 & ~n7138;
  assign n7140 = i_hbusreq3 & ~n7139;
  assign n7141 = ~n4591 & ~n5277;
  assign n7142 = ~controllable_hmaster1 & ~n7141;
  assign n7143 = ~n7068 & ~n7142;
  assign n7144 = ~i_hbusreq3 & ~n7143;
  assign n7145 = ~n7140 & ~n7144;
  assign n7146 = controllable_hmaster2 & ~n7145;
  assign n7147 = ~n5338 & ~n7146;
  assign n7148 = ~controllable_hgrant3 & ~n7147;
  assign n7149 = ~n7136 & ~n7148;
  assign n7150 = controllable_nhgrant0 & ~n7149;
  assign n7151 = ~n5345 & ~n7134;
  assign n7152 = controllable_hgrant3 & ~n7151;
  assign n7153 = ~n3382 & ~n4611;
  assign n7154 = ~controllable_hmaster1 & ~n7153;
  assign n7155 = ~n3381 & ~n7154;
  assign n7156 = i_hbusreq3 & ~n7155;
  assign n7157 = ~n3401 & ~n4636;
  assign n7158 = ~controllable_hmaster1 & ~n7157;
  assign n7159 = ~n3400 & ~n7158;
  assign n7160 = ~i_hbusreq3 & ~n7159;
  assign n7161 = ~n7156 & ~n7160;
  assign n7162 = controllable_hmaster2 & ~n7161;
  assign n7163 = ~n5359 & ~n7162;
  assign n7164 = ~controllable_hgrant3 & ~n7163;
  assign n7165 = ~n7152 & ~n7164;
  assign n7166 = ~controllable_nhgrant0 & ~n7165;
  assign n7167 = ~n7150 & ~n7166;
  assign n7168 = ~n3281 & ~n7167;
  assign n7169 = ~n3281 & ~n7168;
  assign n7170 = n3378 & ~n7169;
  assign n7171 = ~n4553 & ~n4913;
  assign n7172 = ~controllable_hmaster1 & ~n7171;
  assign n7173 = ~n4912 & ~n7172;
  assign n7174 = ~i_hbusreq3 & ~n7173;
  assign n7175 = ~n3951 & ~n7174;
  assign n7176 = controllable_hmaster2 & ~n7175;
  assign n7177 = ~n5400 & ~n7176;
  assign n7178 = controllable_hgrant3 & ~n7177;
  assign n7179 = ~n3854 & ~n5046;
  assign n7180 = ~controllable_hmaster1 & ~n7179;
  assign n7181 = ~n5045 & ~n7180;
  assign n7182 = i_hbusreq3 & ~n7181;
  assign n7183 = ~n4591 & ~n5071;
  assign n7184 = ~controllable_hmaster1 & ~n7183;
  assign n7185 = ~n5070 & ~n7184;
  assign n7186 = ~i_hbusreq3 & ~n7185;
  assign n7187 = ~n7182 & ~n7186;
  assign n7188 = controllable_hmaster2 & ~n7187;
  assign n7189 = ~n5484 & ~n7188;
  assign n7190 = ~controllable_hgrant3 & ~n7189;
  assign n7191 = ~n7178 & ~n7190;
  assign n7192 = controllable_nhgrant0 & ~n7191;
  assign n7193 = ~n5492 & ~n7176;
  assign n7194 = controllable_hgrant3 & ~n7193;
  assign n7195 = ~n4611 & ~n5191;
  assign n7196 = ~controllable_hmaster1 & ~n7195;
  assign n7197 = ~n5190 & ~n7196;
  assign n7198 = i_hbusreq3 & ~n7197;
  assign n7199 = ~n4636 & ~n5197;
  assign n7200 = ~controllable_hmaster1 & ~n7199;
  assign n7201 = ~n5196 & ~n7200;
  assign n7202 = ~i_hbusreq3 & ~n7201;
  assign n7203 = ~n7198 & ~n7202;
  assign n7204 = controllable_hmaster2 & ~n7203;
  assign n7205 = ~n5530 & ~n7204;
  assign n7206 = ~controllable_hgrant3 & ~n7205;
  assign n7207 = ~n7194 & ~n7206;
  assign n7208 = ~controllable_nhgrant0 & ~n7207;
  assign n7209 = ~n7192 & ~n7208;
  assign n7210 = ~n3281 & ~n7209;
  assign n7211 = ~n3281 & ~n7210;
  assign n7212 = ~n3378 & ~n7211;
  assign n7213 = ~n7170 & ~n7212;
  assign n7214 = n3492 & ~n7213;
  assign n7215 = n3492 & ~n7214;
  assign n7216 = n3485 & ~n7215;
  assign n7217 = n3485 & ~n7216;
  assign n7218 = ~n3476 & ~n7217;
  assign n7219 = ~n4031 & ~n4543;
  assign n7220 = i_hlock0 & ~n7219;
  assign n7221 = ~n5564 & ~n7220;
  assign n7222 = ~i_hbusreq0 & ~n7221;
  assign n7223 = ~n4107 & ~n7222;
  assign n7224 = ~i_hbusreq4 & ~n7223;
  assign n7225 = ~n4106 & ~n7224;
  assign n7226 = ~controllable_hgrant4 & ~n7225;
  assign n7227 = ~n4617 & ~n7226;
  assign n7228 = ~i_hbusreq2 & ~n7227;
  assign n7229 = ~n5550 & ~n7228;
  assign n7230 = ~controllable_hgrant2 & ~n7229;
  assign n7231 = ~n4562 & ~n7230;
  assign n7232 = ~controllable_hmaster0 & ~n7231;
  assign n7233 = ~n5562 & ~n7232;
  assign n7234 = ~controllable_hmaster1 & ~n7233;
  assign n7235 = ~n5561 & ~n7234;
  assign n7236 = ~i_hbusreq3 & ~n7235;
  assign n7237 = ~n5549 & ~n7236;
  assign n7238 = controllable_hmaster2 & ~n7237;
  assign n7239 = ~n5613 & ~n7238;
  assign n7240 = controllable_hgrant3 & ~n7239;
  assign n7241 = ~controllable_ndecide & ~n5864;
  assign n7242 = ~controllable_ndecide & ~n7241;
  assign n7243 = i_hready & ~n7242;
  assign n7244 = ~n3379 & ~n7243;
  assign n7245 = ~controllable_hgrant4 & ~n7244;
  assign n7246 = ~n4091 & ~n7245;
  assign n7247 = ~controllable_hgrant2 & ~n7246;
  assign n7248 = ~n5616 & ~n7247;
  assign n7249 = controllable_hmaster1 & ~n7248;
  assign n7250 = controllable_hmaster0 & ~n7248;
  assign n7251 = controllable_locked & ~controllable_ndecide;
  assign n7252 = ~controllable_ndecide & ~n7251;
  assign n7253 = i_hready & ~n7252;
  assign n7254 = ~n3495 & ~n7253;
  assign n7255 = ~controllable_hgrant4 & ~n7254;
  assign n7256 = ~n4015 & ~n7255;
  assign n7257 = ~controllable_hgrant2 & ~n7256;
  assign n7258 = ~n5616 & ~n7257;
  assign n7259 = ~controllable_hmaster0 & ~n7258;
  assign n7260 = ~n7250 & ~n7259;
  assign n7261 = ~controllable_hmaster1 & ~n7260;
  assign n7262 = ~n7249 & ~n7261;
  assign n7263 = i_hbusreq3 & ~n7262;
  assign n7264 = i_hbusreq2 & ~n7246;
  assign n7265 = ~i_hbusreq0 & ~n4110;
  assign n7266 = ~n4107 & ~n7265;
  assign n7267 = ~i_hbusreq4 & ~n7266;
  assign n7268 = ~n4106 & ~n7267;
  assign n7269 = controllable_hgrant4 & ~n7268;
  assign n7270 = i_hbusreq4 & ~n7244;
  assign n7271 = i_hbusreq0 & ~n7244;
  assign n7272 = i_hbusreq1 & ~n5864;
  assign n7273 = i_hbusreq1 & ~n7272;
  assign n7274 = ~controllable_ndecide & ~n7273;
  assign n7275 = ~controllable_ndecide & ~n7274;
  assign n7276 = i_hready & ~n7275;
  assign n7277 = ~n3392 & ~n7276;
  assign n7278 = ~i_hbusreq0 & ~n7277;
  assign n7279 = ~n7271 & ~n7278;
  assign n7280 = ~i_hbusreq4 & ~n7279;
  assign n7281 = ~n7270 & ~n7280;
  assign n7282 = ~controllable_hgrant4 & ~n7281;
  assign n7283 = ~n7269 & ~n7282;
  assign n7284 = ~i_hbusreq2 & ~n7283;
  assign n7285 = ~n7264 & ~n7284;
  assign n7286 = ~controllable_hgrant2 & ~n7285;
  assign n7287 = ~n5635 & ~n7286;
  assign n7288 = controllable_hmaster1 & ~n7287;
  assign n7289 = controllable_hmaster0 & ~n7287;
  assign n7290 = controllable_hgrant2 & ~n7229;
  assign n7291 = i_hbusreq2 & ~n7256;
  assign n7292 = i_hbusreq4 & ~n7254;
  assign n7293 = i_hbusreq0 & ~n7254;
  assign n7294 = i_hbusreq1 & controllable_locked;
  assign n7295 = i_hbusreq1 & ~n7294;
  assign n7296 = ~controllable_ndecide & ~n7295;
  assign n7297 = ~controllable_ndecide & ~n7296;
  assign n7298 = i_hready & ~n7297;
  assign n7299 = ~n4577 & ~n7298;
  assign n7300 = i_hlock0 & ~n7299;
  assign n7301 = ~n3495 & ~n7298;
  assign n7302 = ~i_hlock0 & ~n7301;
  assign n7303 = ~n7300 & ~n7302;
  assign n7304 = ~i_hbusreq0 & ~n7303;
  assign n7305 = ~n7293 & ~n7304;
  assign n7306 = ~i_hbusreq4 & ~n7305;
  assign n7307 = ~n7292 & ~n7306;
  assign n7308 = ~controllable_hgrant4 & ~n7307;
  assign n7309 = ~n4667 & ~n7308;
  assign n7310 = ~i_hbusreq2 & ~n7309;
  assign n7311 = ~n7291 & ~n7310;
  assign n7312 = ~controllable_hgrant2 & ~n7311;
  assign n7313 = ~n7290 & ~n7312;
  assign n7314 = ~controllable_hmaster0 & ~n7313;
  assign n7315 = ~n7289 & ~n7314;
  assign n7316 = ~controllable_hmaster1 & ~n7315;
  assign n7317 = ~n7288 & ~n7316;
  assign n7318 = ~i_hbusreq3 & ~n7317;
  assign n7319 = ~n7263 & ~n7318;
  assign n7320 = controllable_hmaster2 & ~n7319;
  assign n7321 = ~n3379 & ~n7253;
  assign n7322 = ~controllable_hgrant4 & ~n7321;
  assign n7323 = ~n4091 & ~n7322;
  assign n7324 = ~controllable_hgrant2 & ~n7323;
  assign n7325 = ~n5616 & ~n7324;
  assign n7326 = controllable_hmaster0 & ~n7325;
  assign n7327 = ~n5686 & ~n7324;
  assign n7328 = ~controllable_hmaster0 & ~n7327;
  assign n7329 = ~n7326 & ~n7328;
  assign n7330 = controllable_hmaster1 & ~n7329;
  assign n7331 = ~controllable_ndecide & n5961;
  assign n7332 = ~controllable_ndecide & ~n7331;
  assign n7333 = i_hready & ~n7332;
  assign n7334 = ~n3379 & ~n7333;
  assign n7335 = ~controllable_hgrant4 & ~n7334;
  assign n7336 = ~n4091 & ~n7335;
  assign n7337 = ~controllable_hgrant2 & ~n7336;
  assign n7338 = ~n5616 & ~n7337;
  assign n7339 = controllable_hmaster0 & ~n7338;
  assign n7340 = ~controllable_hmaster0 & ~n7325;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = ~controllable_hmaster1 & ~n7341;
  assign n7343 = ~n7330 & ~n7342;
  assign n7344 = i_hbusreq3 & ~n7343;
  assign n7345 = i_hbusreq2 & ~n7323;
  assign n7346 = i_hbusreq4 & ~n7321;
  assign n7347 = i_hbusreq0 & ~n7321;
  assign n7348 = ~n3392 & ~n7298;
  assign n7349 = ~i_hbusreq0 & ~n7348;
  assign n7350 = ~n7347 & ~n7349;
  assign n7351 = ~i_hbusreq4 & ~n7350;
  assign n7352 = ~n7346 & ~n7351;
  assign n7353 = ~controllable_hgrant4 & ~n7352;
  assign n7354 = ~n7269 & ~n7353;
  assign n7355 = ~i_hbusreq2 & ~n7354;
  assign n7356 = ~n7345 & ~n7355;
  assign n7357 = ~controllable_hgrant2 & ~n7356;
  assign n7358 = ~n5635 & ~n7357;
  assign n7359 = controllable_hmaster0 & ~n7358;
  assign n7360 = ~n5722 & ~n7357;
  assign n7361 = ~controllable_hmaster0 & ~n7360;
  assign n7362 = ~n7359 & ~n7361;
  assign n7363 = controllable_hmaster1 & ~n7362;
  assign n7364 = i_hbusreq2 & ~n7336;
  assign n7365 = i_hbusreq4 & ~n7334;
  assign n7366 = i_hbusreq0 & ~n7334;
  assign n7367 = i_hbusreq1 & ~n5961;
  assign n7368 = ~controllable_ndecide & ~n7367;
  assign n7369 = ~controllable_ndecide & ~n7368;
  assign n7370 = i_hready & ~n7369;
  assign n7371 = ~n3392 & ~n7370;
  assign n7372 = ~i_hbusreq0 & ~n7371;
  assign n7373 = ~n7366 & ~n7372;
  assign n7374 = ~i_hbusreq4 & ~n7373;
  assign n7375 = ~n7365 & ~n7374;
  assign n7376 = ~controllable_hgrant4 & ~n7375;
  assign n7377 = ~n7269 & ~n7376;
  assign n7378 = ~i_hbusreq2 & ~n7377;
  assign n7379 = ~n7364 & ~n7378;
  assign n7380 = ~controllable_hgrant2 & ~n7379;
  assign n7381 = ~n5635 & ~n7380;
  assign n7382 = controllable_hmaster0 & ~n7381;
  assign n7383 = ~controllable_hmaster0 & ~n7358;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = ~controllable_hmaster1 & ~n7384;
  assign n7386 = ~n7363 & ~n7385;
  assign n7387 = ~i_hbusreq3 & ~n7386;
  assign n7388 = ~n7344 & ~n7387;
  assign n7389 = ~controllable_hmaster2 & ~n7388;
  assign n7390 = ~n7320 & ~n7389;
  assign n7391 = ~controllable_hgrant3 & ~n7390;
  assign n7392 = ~n7240 & ~n7391;
  assign n7393 = controllable_nhgrant0 & ~n7392;
  assign n7394 = ~n4000 & ~n4605;
  assign n7395 = ~controllable_hgrant4 & ~n7394;
  assign n7396 = ~n3411 & ~n7395;
  assign n7397 = ~controllable_hgrant2 & ~n7396;
  assign n7398 = ~n3410 & ~n7397;
  assign n7399 = ~controllable_hmaster0 & ~n7398;
  assign n7400 = ~n5758 & ~n7399;
  assign n7401 = ~controllable_hmaster1 & ~n7400;
  assign n7402 = ~n5757 & ~n7401;
  assign n7403 = i_hbusreq3 & ~n7402;
  assign n7404 = i_hbusreq2 & ~n7396;
  assign n7405 = i_hbusreq4 & ~n7394;
  assign n7406 = i_hbusreq0 & ~n7394;
  assign n7407 = ~n4031 & ~n4621;
  assign n7408 = i_hlock0 & ~n7407;
  assign n7409 = ~n4031 & ~n4605;
  assign n7410 = ~i_hlock0 & ~n7409;
  assign n7411 = ~n7408 & ~n7410;
  assign n7412 = ~i_hbusreq0 & ~n7411;
  assign n7413 = ~n7406 & ~n7412;
  assign n7414 = ~i_hbusreq4 & ~n7413;
  assign n7415 = ~n7405 & ~n7414;
  assign n7416 = ~controllable_hgrant4 & ~n7415;
  assign n7417 = ~n4617 & ~n7416;
  assign n7418 = ~i_hbusreq2 & ~n7417;
  assign n7419 = ~n7404 & ~n7418;
  assign n7420 = ~controllable_hgrant2 & ~n7419;
  assign n7421 = ~n4562 & ~n7420;
  assign n7422 = ~controllable_hmaster0 & ~n7421;
  assign n7423 = ~n5562 & ~n7422;
  assign n7424 = ~controllable_hmaster1 & ~n7423;
  assign n7425 = ~n5561 & ~n7424;
  assign n7426 = ~i_hbusreq3 & ~n7425;
  assign n7427 = ~n7403 & ~n7426;
  assign n7428 = controllable_hmaster2 & ~n7427;
  assign n7429 = ~n5805 & ~n7428;
  assign n7430 = ~controllable_hgrant3 & ~n7429;
  assign n7431 = ~n7152 & ~n7430;
  assign n7432 = ~controllable_nhgrant0 & ~n7431;
  assign n7433 = ~n7393 & ~n7432;
  assign n7434 = ~n3281 & ~n7433;
  assign n7435 = ~n3281 & ~n7434;
  assign n7436 = n3378 & ~n7435;
  assign n7437 = controllable_hmaster1 & ~n5825;
  assign n7438 = ~n5814 & ~n7220;
  assign n7439 = ~i_hbusreq0 & ~n7438;
  assign n7440 = ~n4107 & ~n7439;
  assign n7441 = ~i_hbusreq4 & ~n7440;
  assign n7442 = ~n4106 & ~n7441;
  assign n7443 = ~controllable_hgrant4 & ~n7442;
  assign n7444 = ~n4617 & ~n7443;
  assign n7445 = ~i_hbusreq2 & ~n7444;
  assign n7446 = ~n5550 & ~n7445;
  assign n7447 = ~controllable_hgrant2 & ~n7446;
  assign n7448 = ~n4562 & ~n7447;
  assign n7449 = ~controllable_hmaster0 & ~n7448;
  assign n7450 = ~n5839 & ~n7449;
  assign n7451 = ~controllable_hmaster1 & ~n7450;
  assign n7452 = ~n7437 & ~n7451;
  assign n7453 = ~i_hbusreq3 & ~n7452;
  assign n7454 = ~n5549 & ~n7453;
  assign n7455 = controllable_hmaster2 & ~n7454;
  assign n7456 = ~n5859 & ~n7455;
  assign n7457 = controllable_hgrant3 & ~n7456;
  assign n7458 = ~n5038 & ~n7241;
  assign n7459 = i_hready & ~n7458;
  assign n7460 = ~n5039 & ~n7459;
  assign n7461 = ~controllable_hgrant4 & ~n7460;
  assign n7462 = ~n4091 & ~n7461;
  assign n7463 = ~controllable_hgrant2 & ~n7462;
  assign n7464 = ~n5616 & ~n7463;
  assign n7465 = controllable_hmaster1 & ~n7464;
  assign n7466 = controllable_hmaster0 & ~n7464;
  assign n7467 = ~n3903 & ~n7251;
  assign n7468 = i_hready & ~n7467;
  assign n7469 = ~n3495 & ~n7468;
  assign n7470 = ~controllable_hgrant4 & ~n7469;
  assign n7471 = ~n4015 & ~n7470;
  assign n7472 = ~controllable_hgrant2 & ~n7471;
  assign n7473 = ~n5616 & ~n7472;
  assign n7474 = ~controllable_hmaster0 & ~n7473;
  assign n7475 = ~n7466 & ~n7474;
  assign n7476 = ~controllable_hmaster1 & ~n7475;
  assign n7477 = ~n7465 & ~n7476;
  assign n7478 = i_hbusreq3 & ~n7477;
  assign n7479 = i_hbusreq2 & ~n7462;
  assign n7480 = i_hlock0 & ~n4110;
  assign n7481 = ~n5814 & ~n7480;
  assign n7482 = ~i_hbusreq0 & ~n7481;
  assign n7483 = ~n4107 & ~n7482;
  assign n7484 = ~i_hbusreq4 & ~n7483;
  assign n7485 = ~n4106 & ~n7484;
  assign n7486 = controllable_hgrant4 & ~n7485;
  assign n7487 = i_hbusreq4 & ~n7460;
  assign n7488 = i_hbusreq0 & ~n7460;
  assign n7489 = ~n5038 & ~n7274;
  assign n7490 = i_hready & ~n7489;
  assign n7491 = ~n5055 & ~n7490;
  assign n7492 = i_hlock0 & ~n7491;
  assign n7493 = ~i_hlock0 & ~n7460;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~i_hbusreq0 & ~n7494;
  assign n7496 = ~n7488 & ~n7495;
  assign n7497 = ~i_hbusreq4 & ~n7496;
  assign n7498 = ~n7487 & ~n7497;
  assign n7499 = ~controllable_hgrant4 & ~n7498;
  assign n7500 = ~n7486 & ~n7499;
  assign n7501 = ~i_hbusreq2 & ~n7500;
  assign n7502 = ~n7479 & ~n7501;
  assign n7503 = ~controllable_hgrant2 & ~n7502;
  assign n7504 = ~n5862 & ~n7503;
  assign n7505 = controllable_hmaster1 & ~n7504;
  assign n7506 = controllable_hmaster0 & ~n7504;
  assign n7507 = controllable_hgrant2 & ~n7446;
  assign n7508 = i_hbusreq2 & ~n7471;
  assign n7509 = i_hbusreq4 & ~n7469;
  assign n7510 = i_hbusreq0 & ~n7469;
  assign n7511 = ~n3903 & ~n7296;
  assign n7512 = i_hready & ~n7511;
  assign n7513 = ~n4577 & ~n7512;
  assign n7514 = i_hlock0 & ~n7513;
  assign n7515 = ~i_hlock0 & ~n7469;
  assign n7516 = ~n7514 & ~n7515;
  assign n7517 = ~i_hbusreq0 & ~n7516;
  assign n7518 = ~n7510 & ~n7517;
  assign n7519 = ~i_hbusreq4 & ~n7518;
  assign n7520 = ~n7509 & ~n7519;
  assign n7521 = ~controllable_hgrant4 & ~n7520;
  assign n7522 = ~n4667 & ~n7521;
  assign n7523 = ~i_hbusreq2 & ~n7522;
  assign n7524 = ~n7508 & ~n7523;
  assign n7525 = ~controllable_hgrant2 & ~n7524;
  assign n7526 = ~n7507 & ~n7525;
  assign n7527 = ~controllable_hmaster0 & ~n7526;
  assign n7528 = ~n7506 & ~n7527;
  assign n7529 = ~controllable_hmaster1 & ~n7528;
  assign n7530 = ~n7505 & ~n7529;
  assign n7531 = ~i_hbusreq3 & ~n7530;
  assign n7532 = ~n7478 & ~n7531;
  assign n7533 = controllable_hmaster2 & ~n7532;
  assign n7534 = ~n3904 & ~n7468;
  assign n7535 = ~controllable_hgrant4 & ~n7534;
  assign n7536 = ~n4091 & ~n7535;
  assign n7537 = ~controllable_hgrant2 & ~n7536;
  assign n7538 = ~n5616 & ~n7537;
  assign n7539 = controllable_hmaster0 & ~n7538;
  assign n7540 = ~n5686 & ~n7537;
  assign n7541 = ~controllable_hmaster0 & ~n7540;
  assign n7542 = ~n7539 & ~n7541;
  assign n7543 = controllable_hmaster1 & ~n7542;
  assign n7544 = ~n3903 & ~n7331;
  assign n7545 = i_hready & ~n7544;
  assign n7546 = ~n3904 & ~n7545;
  assign n7547 = ~controllable_hgrant4 & ~n7546;
  assign n7548 = ~n4091 & ~n7547;
  assign n7549 = ~controllable_hgrant2 & ~n7548;
  assign n7550 = ~n5616 & ~n7549;
  assign n7551 = controllable_hmaster0 & ~n7550;
  assign n7552 = ~controllable_hmaster0 & ~n7538;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~controllable_hmaster1 & ~n7553;
  assign n7555 = ~n7543 & ~n7554;
  assign n7556 = i_hbusreq3 & ~n7555;
  assign n7557 = i_hbusreq2 & ~n7536;
  assign n7558 = i_hbusreq4 & ~n7534;
  assign n7559 = i_hbusreq0 & ~n7534;
  assign n7560 = ~n3920 & ~n7512;
  assign n7561 = i_hlock0 & ~n7560;
  assign n7562 = ~i_hlock0 & ~n7534;
  assign n7563 = ~n7561 & ~n7562;
  assign n7564 = ~i_hbusreq0 & ~n7563;
  assign n7565 = ~n7559 & ~n7564;
  assign n7566 = ~i_hbusreq4 & ~n7565;
  assign n7567 = ~n7558 & ~n7566;
  assign n7568 = ~controllable_hgrant4 & ~n7567;
  assign n7569 = ~n7486 & ~n7568;
  assign n7570 = ~i_hbusreq2 & ~n7569;
  assign n7571 = ~n7557 & ~n7570;
  assign n7572 = ~controllable_hgrant2 & ~n7571;
  assign n7573 = ~n5862 & ~n7572;
  assign n7574 = controllable_hmaster0 & ~n7573;
  assign n7575 = ~n5950 & ~n7572;
  assign n7576 = ~controllable_hmaster0 & ~n7575;
  assign n7577 = ~n7574 & ~n7576;
  assign n7578 = controllable_hmaster1 & ~n7577;
  assign n7579 = i_hbusreq2 & ~n7548;
  assign n7580 = i_hbusreq4 & ~n7546;
  assign n7581 = i_hbusreq0 & ~n7546;
  assign n7582 = ~n3903 & ~n7368;
  assign n7583 = i_hready & ~n7582;
  assign n7584 = ~n3920 & ~n7583;
  assign n7585 = i_hlock0 & ~n7584;
  assign n7586 = ~i_hlock0 & ~n7546;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = ~i_hbusreq0 & ~n7587;
  assign n7589 = ~n7581 & ~n7588;
  assign n7590 = ~i_hbusreq4 & ~n7589;
  assign n7591 = ~n7580 & ~n7590;
  assign n7592 = ~controllable_hgrant4 & ~n7591;
  assign n7593 = ~n7486 & ~n7592;
  assign n7594 = ~i_hbusreq2 & ~n7593;
  assign n7595 = ~n7579 & ~n7594;
  assign n7596 = ~controllable_hgrant2 & ~n7595;
  assign n7597 = ~n5862 & ~n7596;
  assign n7598 = controllable_hmaster0 & ~n7597;
  assign n7599 = ~n4000 & ~n5384;
  assign n7600 = i_hlock0 & ~n7599;
  assign n7601 = ~n5814 & ~n7600;
  assign n7602 = ~i_hbusreq0 & ~n7601;
  assign n7603 = ~n4107 & ~n7602;
  assign n7604 = ~i_hbusreq4 & ~n7603;
  assign n7605 = ~n4106 & ~n7604;
  assign n7606 = controllable_hgrant4 & ~n7605;
  assign n7607 = ~n5464 & ~n7512;
  assign n7608 = i_hlock0 & ~n7607;
  assign n7609 = ~n7562 & ~n7608;
  assign n7610 = ~i_hbusreq0 & ~n7609;
  assign n7611 = ~n7559 & ~n7610;
  assign n7612 = ~i_hbusreq4 & ~n7611;
  assign n7613 = ~n7558 & ~n7612;
  assign n7614 = ~controllable_hgrant4 & ~n7613;
  assign n7615 = ~n7606 & ~n7614;
  assign n7616 = ~i_hbusreq2 & ~n7615;
  assign n7617 = ~n7557 & ~n7616;
  assign n7618 = ~controllable_hgrant2 & ~n7617;
  assign n7619 = ~n5981 & ~n7618;
  assign n7620 = ~controllable_hmaster0 & ~n7619;
  assign n7621 = ~n7598 & ~n7620;
  assign n7622 = ~controllable_hmaster1 & ~n7621;
  assign n7623 = ~n7578 & ~n7622;
  assign n7624 = ~i_hbusreq3 & ~n7623;
  assign n7625 = ~n7556 & ~n7624;
  assign n7626 = ~controllable_hmaster2 & ~n7625;
  assign n7627 = ~n7533 & ~n7626;
  assign n7628 = ~controllable_hgrant3 & ~n7627;
  assign n7629 = ~n7457 & ~n7628;
  assign n7630 = controllable_nhgrant0 & ~n7629;
  assign n7631 = ~n4605 & ~n6007;
  assign n7632 = ~controllable_hgrant4 & ~n7631;
  assign n7633 = ~n3411 & ~n7632;
  assign n7634 = ~controllable_hgrant2 & ~n7633;
  assign n7635 = ~n3410 & ~n7634;
  assign n7636 = ~controllable_hmaster0 & ~n7635;
  assign n7637 = ~n6037 & ~n7636;
  assign n7638 = ~controllable_hmaster1 & ~n7637;
  assign n7639 = ~n6036 & ~n7638;
  assign n7640 = i_hbusreq3 & ~n7639;
  assign n7641 = i_hbusreq2 & ~n7633;
  assign n7642 = i_hbusreq4 & ~n7631;
  assign n7643 = i_hbusreq0 & ~n7631;
  assign n7644 = ~n4621 & ~n6018;
  assign n7645 = i_hlock0 & ~n7644;
  assign n7646 = ~i_hlock0 & ~n7631;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = ~i_hbusreq0 & ~n7647;
  assign n7649 = ~n7643 & ~n7648;
  assign n7650 = ~i_hbusreq4 & ~n7649;
  assign n7651 = ~n7642 & ~n7650;
  assign n7652 = ~controllable_hgrant4 & ~n7651;
  assign n7653 = ~n4617 & ~n7652;
  assign n7654 = ~i_hbusreq2 & ~n7653;
  assign n7655 = ~n7641 & ~n7654;
  assign n7656 = ~controllable_hgrant2 & ~n7655;
  assign n7657 = ~n4562 & ~n7656;
  assign n7658 = ~controllable_hmaster0 & ~n7657;
  assign n7659 = ~n6050 & ~n7658;
  assign n7660 = ~controllable_hmaster1 & ~n7659;
  assign n7661 = ~n6049 & ~n7660;
  assign n7662 = ~i_hbusreq3 & ~n7661;
  assign n7663 = ~n7640 & ~n7662;
  assign n7664 = controllable_hmaster2 & ~n7663;
  assign n7665 = ~n6078 & ~n7664;
  assign n7666 = ~controllable_hgrant3 & ~n7665;
  assign n7667 = ~n7194 & ~n7666;
  assign n7668 = ~controllable_nhgrant0 & ~n7667;
  assign n7669 = ~n7630 & ~n7668;
  assign n7670 = ~n3281 & ~n7669;
  assign n7671 = ~n3281 & ~n7670;
  assign n7672 = ~n3378 & ~n7671;
  assign n7673 = ~n7436 & ~n7672;
  assign n7674 = n3492 & ~n7673;
  assign n7675 = n3492 & ~n7674;
  assign n7676 = n3485 & ~n7675;
  assign n7677 = n3485 & ~n7676;
  assign n7678 = n3476 & ~n7677;
  assign n7679 = ~n7218 & ~n7678;
  assign n7680 = n3374 & ~n7679;
  assign n7681 = ~n7128 & ~n7680;
  assign n7682 = n3655 & ~n7681;
  assign n7683 = controllable_hmaster0 & ~n6105;
  assign n7684 = ~controllable_hmaster1 & ~n7683;
  assign n7685 = ~n6104 & ~n7684;
  assign n7686 = i_hbusreq3 & ~n7685;
  assign n7687 = controllable_hmaster0 & ~n6130;
  assign n7688 = ~controllable_hmaster1 & ~n7687;
  assign n7689 = ~n6129 & ~n7688;
  assign n7690 = ~i_hbusreq3 & ~n7689;
  assign n7691 = ~n7686 & ~n7690;
  assign n7692 = controllable_hmaster2 & ~n7691;
  assign n7693 = controllable_hmaster2 & ~n7692;
  assign n7694 = ~controllable_hgrant3 & ~n7693;
  assign n7695 = ~n7090 & ~n7694;
  assign n7696 = controllable_nhgrant0 & ~n7695;
  assign n7697 = ~n7118 & ~n7696;
  assign n7698 = ~n3281 & ~n7697;
  assign n7699 = ~n3281 & ~n7698;
  assign n7700 = ~n3378 & ~n7699;
  assign n7701 = ~n7082 & ~n7700;
  assign n7702 = n3492 & ~n7701;
  assign n7703 = n3492 & ~n7702;
  assign n7704 = n3485 & ~n7703;
  assign n7705 = n3485 & ~n7704;
  assign n7706 = ~n3374 & ~n7705;
  assign n7707 = ~n4705 & ~n5260;
  assign n7708 = ~controllable_hmaster1 & ~n7707;
  assign n7709 = ~n7063 & ~n7708;
  assign n7710 = i_hbusreq3 & ~n7709;
  assign n7711 = ~n4729 & ~n5277;
  assign n7712 = ~controllable_hmaster1 & ~n7711;
  assign n7713 = ~n7068 & ~n7712;
  assign n7714 = ~i_hbusreq3 & ~n7713;
  assign n7715 = ~n7710 & ~n7714;
  assign n7716 = controllable_hmaster2 & ~n7715;
  assign n7717 = ~n5338 & ~n7716;
  assign n7718 = ~controllable_hgrant3 & ~n7717;
  assign n7719 = ~n7136 & ~n7718;
  assign n7720 = controllable_nhgrant0 & ~n7719;
  assign n7721 = ~n7166 & ~n7720;
  assign n7722 = ~n3281 & ~n7721;
  assign n7723 = ~n3281 & ~n7722;
  assign n7724 = n3378 & ~n7723;
  assign n7725 = ~n4705 & ~n6105;
  assign n7726 = ~controllable_hmaster1 & ~n7725;
  assign n7727 = ~n6104 & ~n7726;
  assign n7728 = i_hbusreq3 & ~n7727;
  assign n7729 = ~n4729 & ~n6130;
  assign n7730 = ~controllable_hmaster1 & ~n7729;
  assign n7731 = ~n6129 & ~n7730;
  assign n7732 = ~i_hbusreq3 & ~n7731;
  assign n7733 = ~n7728 & ~n7732;
  assign n7734 = controllable_hmaster2 & ~n7733;
  assign n7735 = ~n6343 & ~n7734;
  assign n7736 = ~controllable_hgrant3 & ~n7735;
  assign n7737 = ~n7178 & ~n7736;
  assign n7738 = controllable_nhgrant0 & ~n7737;
  assign n7739 = ~n7208 & ~n7738;
  assign n7740 = ~n3281 & ~n7739;
  assign n7741 = ~n3281 & ~n7740;
  assign n7742 = ~n3378 & ~n7741;
  assign n7743 = ~n7724 & ~n7742;
  assign n7744 = n3492 & ~n7743;
  assign n7745 = n3492 & ~n7744;
  assign n7746 = n3485 & ~n7745;
  assign n7747 = n3485 & ~n7746;
  assign n7748 = ~n3476 & ~n7747;
  assign n7749 = ~n4699 & ~n7253;
  assign n7750 = ~controllable_hgrant4 & ~n7749;
  assign n7751 = ~n4015 & ~n7750;
  assign n7752 = ~controllable_hgrant2 & ~n7751;
  assign n7753 = ~n5616 & ~n7752;
  assign n7754 = ~controllable_hmaster0 & ~n7753;
  assign n7755 = ~n7250 & ~n7754;
  assign n7756 = ~controllable_hmaster1 & ~n7755;
  assign n7757 = ~n7249 & ~n7756;
  assign n7758 = i_hbusreq3 & ~n7757;
  assign n7759 = i_hbusreq2 & ~n7751;
  assign n7760 = i_hbusreq4 & ~n7749;
  assign n7761 = i_hbusreq0 & ~n7749;
  assign n7762 = ~n4714 & ~n7298;
  assign n7763 = i_hlock0 & ~n7762;
  assign n7764 = ~n4699 & ~n7298;
  assign n7765 = ~i_hlock0 & ~n7764;
  assign n7766 = ~n7763 & ~n7765;
  assign n7767 = ~i_hbusreq0 & ~n7766;
  assign n7768 = ~n7761 & ~n7767;
  assign n7769 = ~i_hbusreq4 & ~n7768;
  assign n7770 = ~n7760 & ~n7769;
  assign n7771 = ~controllable_hgrant4 & ~n7770;
  assign n7772 = ~n4667 & ~n7771;
  assign n7773 = ~i_hbusreq2 & ~n7772;
  assign n7774 = ~n7759 & ~n7773;
  assign n7775 = ~controllable_hgrant2 & ~n7774;
  assign n7776 = ~n7290 & ~n7775;
  assign n7777 = ~controllable_hmaster0 & ~n7776;
  assign n7778 = ~n7289 & ~n7777;
  assign n7779 = ~controllable_hmaster1 & ~n7778;
  assign n7780 = ~n7288 & ~n7779;
  assign n7781 = ~i_hbusreq3 & ~n7780;
  assign n7782 = ~n7758 & ~n7781;
  assign n7783 = controllable_hmaster2 & ~n7782;
  assign n7784 = ~n7389 & ~n7783;
  assign n7785 = ~controllable_hgrant3 & ~n7784;
  assign n7786 = ~n7240 & ~n7785;
  assign n7787 = controllable_nhgrant0 & ~n7786;
  assign n7788 = ~n7432 & ~n7787;
  assign n7789 = ~n3281 & ~n7788;
  assign n7790 = ~n3281 & ~n7789;
  assign n7791 = n3378 & ~n7790;
  assign n7792 = i_hready & ~n5864;
  assign n7793 = ~n6098 & ~n7792;
  assign n7794 = ~controllable_hgrant4 & ~n7793;
  assign n7795 = ~n4091 & ~n7794;
  assign n7796 = ~controllable_hgrant2 & ~n7795;
  assign n7797 = ~n5616 & ~n7796;
  assign n7798 = controllable_hmaster1 & ~n7797;
  assign n7799 = controllable_hmaster0 & ~n7797;
  assign n7800 = i_hready & controllable_locked;
  assign n7801 = ~n4699 & ~n7800;
  assign n7802 = ~controllable_hgrant4 & ~n7801;
  assign n7803 = ~n4015 & ~n7802;
  assign n7804 = ~controllable_hgrant2 & ~n7803;
  assign n7805 = ~n5616 & ~n7804;
  assign n7806 = ~controllable_hmaster0 & ~n7805;
  assign n7807 = ~n7799 & ~n7806;
  assign n7808 = ~controllable_hmaster1 & ~n7807;
  assign n7809 = ~n7798 & ~n7808;
  assign n7810 = i_hbusreq3 & ~n7809;
  assign n7811 = i_hbusreq2 & ~n7795;
  assign n7812 = i_hbusreq4 & ~n7793;
  assign n7813 = i_hbusreq0 & ~n7793;
  assign n7814 = ~n6097 & ~n7274;
  assign n7815 = i_hready & ~n7814;
  assign n7816 = ~n6114 & ~n7815;
  assign n7817 = i_hlock0 & ~n7816;
  assign n7818 = ~i_hlock0 & ~n7793;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = ~i_hbusreq0 & ~n7819;
  assign n7821 = ~n7813 & ~n7820;
  assign n7822 = ~i_hbusreq4 & ~n7821;
  assign n7823 = ~n7812 & ~n7822;
  assign n7824 = ~controllable_hgrant4 & ~n7823;
  assign n7825 = ~n7486 & ~n7824;
  assign n7826 = ~i_hbusreq2 & ~n7825;
  assign n7827 = ~n7811 & ~n7826;
  assign n7828 = ~controllable_hgrant2 & ~n7827;
  assign n7829 = ~n5862 & ~n7828;
  assign n7830 = controllable_hmaster1 & ~n7829;
  assign n7831 = controllable_hmaster0 & ~n7829;
  assign n7832 = i_hbusreq2 & ~n7803;
  assign n7833 = i_hbusreq4 & ~n7801;
  assign n7834 = i_hbusreq0 & ~n7801;
  assign n7835 = ~n6247 & ~n7296;
  assign n7836 = i_hready & ~n7835;
  assign n7837 = ~n4714 & ~n7836;
  assign n7838 = i_hlock0 & ~n7837;
  assign n7839 = ~i_hlock0 & ~n7801;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = ~i_hbusreq0 & ~n7840;
  assign n7842 = ~n7834 & ~n7841;
  assign n7843 = ~i_hbusreq4 & ~n7842;
  assign n7844 = ~n7833 & ~n7843;
  assign n7845 = ~controllable_hgrant4 & ~n7844;
  assign n7846 = ~n4667 & ~n7845;
  assign n7847 = ~i_hbusreq2 & ~n7846;
  assign n7848 = ~n7832 & ~n7847;
  assign n7849 = ~controllable_hgrant2 & ~n7848;
  assign n7850 = ~n7507 & ~n7849;
  assign n7851 = ~controllable_hmaster0 & ~n7850;
  assign n7852 = ~n7831 & ~n7851;
  assign n7853 = ~controllable_hmaster1 & ~n7852;
  assign n7854 = ~n7830 & ~n7853;
  assign n7855 = ~i_hbusreq3 & ~n7854;
  assign n7856 = ~n7810 & ~n7855;
  assign n7857 = controllable_hmaster2 & ~n7856;
  assign n7858 = ~n6248 & ~n7800;
  assign n7859 = ~controllable_hgrant4 & ~n7858;
  assign n7860 = ~n4091 & ~n7859;
  assign n7861 = ~controllable_hgrant2 & ~n7860;
  assign n7862 = ~n5616 & ~n7861;
  assign n7863 = controllable_hmaster0 & ~n7862;
  assign n7864 = ~n5686 & ~n7861;
  assign n7865 = ~controllable_hmaster0 & ~n7864;
  assign n7866 = ~n7863 & ~n7865;
  assign n7867 = controllable_hmaster1 & ~n7866;
  assign n7868 = i_hready & ~n5961;
  assign n7869 = ~n6262 & ~n7868;
  assign n7870 = ~controllable_hgrant4 & n7869;
  assign n7871 = ~n4091 & ~n7870;
  assign n7872 = ~controllable_hgrant2 & ~n7871;
  assign n7873 = ~n5616 & ~n7872;
  assign n7874 = controllable_hmaster0 & ~n7873;
  assign n7875 = ~controllable_hmaster0 & ~n7862;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = ~controllable_hmaster1 & ~n7876;
  assign n7878 = ~n7867 & ~n7877;
  assign n7879 = i_hbusreq3 & ~n7878;
  assign n7880 = i_hbusreq2 & ~n7860;
  assign n7881 = i_hbusreq4 & ~n7858;
  assign n7882 = i_hbusreq0 & ~n7858;
  assign n7883 = ~n6278 & ~n7836;
  assign n7884 = i_hlock0 & ~n7883;
  assign n7885 = ~i_hlock0 & ~n7858;
  assign n7886 = ~n7884 & ~n7885;
  assign n7887 = ~i_hbusreq0 & ~n7886;
  assign n7888 = ~n7882 & ~n7887;
  assign n7889 = ~i_hbusreq4 & ~n7888;
  assign n7890 = ~n7881 & ~n7889;
  assign n7891 = ~controllable_hgrant4 & ~n7890;
  assign n7892 = ~n7486 & ~n7891;
  assign n7893 = ~i_hbusreq2 & ~n7892;
  assign n7894 = ~n7880 & ~n7893;
  assign n7895 = ~controllable_hgrant2 & ~n7894;
  assign n7896 = ~n5862 & ~n7895;
  assign n7897 = controllable_hmaster0 & ~n7896;
  assign n7898 = ~n5950 & ~n7895;
  assign n7899 = ~controllable_hmaster0 & ~n7898;
  assign n7900 = ~n7897 & ~n7899;
  assign n7901 = controllable_hmaster1 & ~n7900;
  assign n7902 = i_hbusreq2 & ~n7871;
  assign n7903 = i_hbusreq4 & ~n7869;
  assign n7904 = i_hbusreq0 & ~n7869;
  assign n7905 = ~controllable_ndecide & n7367;
  assign n7906 = ~n6260 & ~n7905;
  assign n7907 = i_hready & ~n7906;
  assign n7908 = ~n6306 & ~n7907;
  assign n7909 = i_hlock0 & ~n7908;
  assign n7910 = ~i_hlock0 & ~n7869;
  assign n7911 = ~n7909 & ~n7910;
  assign n7912 = ~i_hbusreq0 & ~n7911;
  assign n7913 = ~n7904 & ~n7912;
  assign n7914 = ~i_hbusreq4 & ~n7913;
  assign n7915 = ~n7903 & ~n7914;
  assign n7916 = ~controllable_hgrant4 & n7915;
  assign n7917 = ~n7486 & ~n7916;
  assign n7918 = ~i_hbusreq2 & ~n7917;
  assign n7919 = ~n7902 & ~n7918;
  assign n7920 = ~controllable_hgrant2 & ~n7919;
  assign n7921 = ~n5862 & ~n7920;
  assign n7922 = controllable_hmaster0 & ~n7921;
  assign n7923 = ~n6323 & ~n7836;
  assign n7924 = i_hlock0 & ~n7923;
  assign n7925 = ~n7885 & ~n7924;
  assign n7926 = ~i_hbusreq0 & ~n7925;
  assign n7927 = ~n7882 & ~n7926;
  assign n7928 = ~i_hbusreq4 & ~n7927;
  assign n7929 = ~n7881 & ~n7928;
  assign n7930 = ~controllable_hgrant4 & ~n7929;
  assign n7931 = ~n7606 & ~n7930;
  assign n7932 = ~i_hbusreq2 & ~n7931;
  assign n7933 = ~n7880 & ~n7932;
  assign n7934 = ~controllable_hgrant2 & ~n7933;
  assign n7935 = ~n5981 & ~n7934;
  assign n7936 = ~controllable_hmaster0 & ~n7935;
  assign n7937 = ~n7922 & ~n7936;
  assign n7938 = ~controllable_hmaster1 & ~n7937;
  assign n7939 = ~n7901 & ~n7938;
  assign n7940 = ~i_hbusreq3 & ~n7939;
  assign n7941 = ~n7879 & ~n7940;
  assign n7942 = ~controllable_hmaster2 & ~n7941;
  assign n7943 = ~n7857 & ~n7942;
  assign n7944 = ~controllable_hgrant3 & ~n7943;
  assign n7945 = ~n7457 & ~n7944;
  assign n7946 = controllable_nhgrant0 & ~n7945;
  assign n7947 = ~n7668 & ~n7946;
  assign n7948 = ~n3281 & ~n7947;
  assign n7949 = ~n3281 & ~n7948;
  assign n7950 = ~n3378 & ~n7949;
  assign n7951 = ~n7791 & ~n7950;
  assign n7952 = n3492 & ~n7951;
  assign n7953 = n3492 & ~n7952;
  assign n7954 = n3485 & ~n7953;
  assign n7955 = n3485 & ~n7954;
  assign n7956 = n3476 & ~n7955;
  assign n7957 = ~n7748 & ~n7956;
  assign n7958 = n3374 & ~n7957;
  assign n7959 = ~n7706 & ~n7958;
  assign n7960 = ~n3655 & ~n7959;
  assign n7961 = ~n7682 & ~n7960;
  assign n7962 = n3652 & ~n7961;
  assign n7963 = controllable_hmaster0 & ~n6577;
  assign n7964 = ~controllable_hmaster1 & ~n7963;
  assign n7965 = ~n6576 & ~n7964;
  assign n7966 = i_hbusreq3 & ~n7965;
  assign n7967 = controllable_hmaster0 & ~n6584;
  assign n7968 = ~controllable_hmaster1 & ~n7967;
  assign n7969 = ~n6583 & ~n7968;
  assign n7970 = ~i_hbusreq3 & ~n7969;
  assign n7971 = ~n7966 & ~n7970;
  assign n7972 = controllable_hmaster2 & ~n7971;
  assign n7973 = controllable_hmaster2 & ~n7972;
  assign n7974 = ~controllable_hgrant3 & ~n7973;
  assign n7975 = ~n7090 & ~n7974;
  assign n7976 = controllable_nhgrant0 & ~n7975;
  assign n7977 = ~n7118 & ~n7976;
  assign n7978 = ~n3281 & ~n7977;
  assign n7979 = ~n3281 & ~n7978;
  assign n7980 = ~n3378 & ~n7979;
  assign n7981 = ~n7082 & ~n7980;
  assign n7982 = n3492 & ~n7981;
  assign n7983 = n3492 & ~n7982;
  assign n7984 = n3485 & ~n7983;
  assign n7985 = n3485 & ~n7984;
  assign n7986 = ~n3374 & ~n7985;
  assign n7987 = ~n4789 & ~n5260;
  assign n7988 = ~controllable_hmaster1 & ~n7987;
  assign n7989 = ~n7063 & ~n7988;
  assign n7990 = i_hbusreq3 & ~n7989;
  assign n7991 = ~n4796 & ~n5277;
  assign n7992 = ~controllable_hmaster1 & ~n7991;
  assign n7993 = ~n7068 & ~n7992;
  assign n7994 = ~i_hbusreq3 & ~n7993;
  assign n7995 = ~n7990 & ~n7994;
  assign n7996 = controllable_hmaster2 & ~n7995;
  assign n7997 = ~n5338 & ~n7996;
  assign n7998 = ~controllable_hgrant3 & ~n7997;
  assign n7999 = ~n7136 & ~n7998;
  assign n8000 = controllable_nhgrant0 & ~n7999;
  assign n8001 = ~n7166 & ~n8000;
  assign n8002 = ~n3281 & ~n8001;
  assign n8003 = ~n3281 & ~n8002;
  assign n8004 = n3378 & ~n8003;
  assign n8005 = ~n4789 & ~n6577;
  assign n8006 = ~controllable_hmaster1 & ~n8005;
  assign n8007 = ~n6576 & ~n8006;
  assign n8008 = i_hbusreq3 & ~n8007;
  assign n8009 = ~n4796 & ~n6584;
  assign n8010 = ~controllable_hmaster1 & ~n8009;
  assign n8011 = ~n6583 & ~n8010;
  assign n8012 = ~i_hbusreq3 & ~n8011;
  assign n8013 = ~n8008 & ~n8012;
  assign n8014 = controllable_hmaster2 & ~n8013;
  assign n8015 = ~n6723 & ~n8014;
  assign n8016 = ~controllable_hgrant3 & ~n8015;
  assign n8017 = ~n7178 & ~n8016;
  assign n8018 = controllable_nhgrant0 & ~n8017;
  assign n8019 = ~n7208 & ~n8018;
  assign n8020 = ~n3281 & ~n8019;
  assign n8021 = ~n3281 & ~n8020;
  assign n8022 = ~n3378 & ~n8021;
  assign n8023 = ~n8004 & ~n8022;
  assign n8024 = n3492 & ~n8023;
  assign n8025 = n3492 & ~n8024;
  assign n8026 = n3485 & ~n8025;
  assign n8027 = n3485 & ~n8026;
  assign n8028 = ~n3476 & ~n8027;
  assign n8029 = controllable_hgrant2 & ~n7396;
  assign n8030 = ~n7257 & ~n8029;
  assign n8031 = ~controllable_hmaster0 & ~n8030;
  assign n8032 = ~n7250 & ~n8031;
  assign n8033 = ~controllable_hmaster1 & ~n8032;
  assign n8034 = ~n7249 & ~n8033;
  assign n8035 = i_hbusreq3 & ~n8034;
  assign n8036 = controllable_hgrant2 & ~n7419;
  assign n8037 = ~n7312 & ~n8036;
  assign n8038 = ~controllable_hmaster0 & ~n8037;
  assign n8039 = ~n7289 & ~n8038;
  assign n8040 = ~controllable_hmaster1 & ~n8039;
  assign n8041 = ~n7288 & ~n8040;
  assign n8042 = ~i_hbusreq3 & ~n8041;
  assign n8043 = ~n8035 & ~n8042;
  assign n8044 = controllable_hmaster2 & ~n8043;
  assign n8045 = ~n7389 & ~n8044;
  assign n8046 = ~controllable_hgrant3 & ~n8045;
  assign n8047 = ~n7240 & ~n8046;
  assign n8048 = controllable_nhgrant0 & ~n8047;
  assign n8049 = ~n7432 & ~n8048;
  assign n8050 = ~n3281 & ~n8049;
  assign n8051 = ~n3281 & ~n8050;
  assign n8052 = n3378 & ~n8051;
  assign n8053 = ~n6762 & ~n7463;
  assign n8054 = controllable_hmaster1 & ~n8053;
  assign n8055 = controllable_hmaster0 & ~n8053;
  assign n8056 = controllable_hgrant2 & ~n7633;
  assign n8057 = ~n7472 & ~n8056;
  assign n8058 = ~controllable_hmaster0 & ~n8057;
  assign n8059 = ~n8055 & ~n8058;
  assign n8060 = ~controllable_hmaster1 & ~n8059;
  assign n8061 = ~n8054 & ~n8060;
  assign n8062 = i_hbusreq3 & ~n8061;
  assign n8063 = ~n6772 & ~n7503;
  assign n8064 = controllable_hmaster1 & ~n8063;
  assign n8065 = controllable_hmaster0 & ~n8063;
  assign n8066 = controllable_hgrant2 & ~n7655;
  assign n8067 = ~n7525 & ~n8066;
  assign n8068 = ~controllable_hmaster0 & ~n8067;
  assign n8069 = ~n8065 & ~n8068;
  assign n8070 = ~controllable_hmaster1 & ~n8069;
  assign n8071 = ~n8064 & ~n8070;
  assign n8072 = ~i_hbusreq3 & ~n8071;
  assign n8073 = ~n8062 & ~n8072;
  assign n8074 = controllable_hmaster2 & ~n8073;
  assign n8075 = ~n6762 & ~n7537;
  assign n8076 = controllable_hmaster0 & ~n8075;
  assign n8077 = ~n6786 & ~n7537;
  assign n8078 = ~controllable_hmaster0 & ~n8077;
  assign n8079 = ~n8076 & ~n8078;
  assign n8080 = controllable_hmaster1 & ~n8079;
  assign n8081 = ~n6762 & ~n7549;
  assign n8082 = controllable_hmaster0 & ~n8081;
  assign n8083 = ~controllable_hmaster0 & ~n8075;
  assign n8084 = ~n8082 & ~n8083;
  assign n8085 = ~controllable_hmaster1 & ~n8084;
  assign n8086 = ~n8080 & ~n8085;
  assign n8087 = i_hbusreq3 & ~n8086;
  assign n8088 = ~n6772 & ~n7572;
  assign n8089 = controllable_hmaster0 & ~n8088;
  assign n8090 = ~n6813 & ~n7572;
  assign n8091 = ~controllable_hmaster0 & ~n8090;
  assign n8092 = ~n8089 & ~n8091;
  assign n8093 = controllable_hmaster1 & ~n8092;
  assign n8094 = ~n6772 & ~n7596;
  assign n8095 = controllable_hmaster0 & ~n8094;
  assign n8096 = ~n6831 & ~n7618;
  assign n8097 = ~controllable_hmaster0 & ~n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = ~controllable_hmaster1 & ~n8098;
  assign n8100 = ~n8093 & ~n8099;
  assign n8101 = ~i_hbusreq3 & ~n8100;
  assign n8102 = ~n8087 & ~n8101;
  assign n8103 = ~controllable_hmaster2 & ~n8102;
  assign n8104 = ~n8074 & ~n8103;
  assign n8105 = ~controllable_hgrant3 & ~n8104;
  assign n8106 = ~n7457 & ~n8105;
  assign n8107 = controllable_nhgrant0 & ~n8106;
  assign n8108 = ~n7668 & ~n8107;
  assign n8109 = ~n3281 & ~n8108;
  assign n8110 = ~n3281 & ~n8109;
  assign n8111 = ~n3378 & ~n8110;
  assign n8112 = ~n8052 & ~n8111;
  assign n8113 = n3492 & ~n8112;
  assign n8114 = n3492 & ~n8113;
  assign n8115 = n3485 & ~n8114;
  assign n8116 = n3485 & ~n8115;
  assign n8117 = n3476 & ~n8116;
  assign n8118 = ~n8028 & ~n8117;
  assign n8119 = n3374 & ~n8118;
  assign n8120 = ~n7986 & ~n8119;
  assign n8121 = n3655 & ~n8120;
  assign n8122 = controllable_hmaster0 & ~n6860;
  assign n8123 = ~controllable_hmaster1 & ~n8122;
  assign n8124 = ~n6859 & ~n8123;
  assign n8125 = i_hbusreq3 & ~n8124;
  assign n8126 = controllable_hmaster0 & ~n6867;
  assign n8127 = ~controllable_hmaster1 & ~n8126;
  assign n8128 = ~n6866 & ~n8127;
  assign n8129 = ~i_hbusreq3 & ~n8128;
  assign n8130 = ~n8125 & ~n8129;
  assign n8131 = controllable_hmaster2 & ~n8130;
  assign n8132 = controllable_hmaster2 & ~n8131;
  assign n8133 = ~controllable_hgrant3 & ~n8132;
  assign n8134 = ~n7090 & ~n8133;
  assign n8135 = controllable_nhgrant0 & ~n8134;
  assign n8136 = ~n7118 & ~n8135;
  assign n8137 = ~n3281 & ~n8136;
  assign n8138 = ~n3281 & ~n8137;
  assign n8139 = ~n3378 & ~n8138;
  assign n8140 = ~n7082 & ~n8139;
  assign n8141 = n3492 & ~n8140;
  assign n8142 = n3492 & ~n8141;
  assign n8143 = n3485 & ~n8142;
  assign n8144 = n3485 & ~n8143;
  assign n8145 = ~n3374 & ~n8144;
  assign n8146 = ~n4846 & ~n5260;
  assign n8147 = ~controllable_hmaster1 & ~n8146;
  assign n8148 = ~n7063 & ~n8147;
  assign n8149 = i_hbusreq3 & ~n8148;
  assign n8150 = ~n4852 & ~n5277;
  assign n8151 = ~controllable_hmaster1 & ~n8150;
  assign n8152 = ~n7068 & ~n8151;
  assign n8153 = ~i_hbusreq3 & ~n8152;
  assign n8154 = ~n8149 & ~n8153;
  assign n8155 = controllable_hmaster2 & ~n8154;
  assign n8156 = ~n5338 & ~n8155;
  assign n8157 = ~controllable_hgrant3 & ~n8156;
  assign n8158 = ~n7136 & ~n8157;
  assign n8159 = controllable_nhgrant0 & ~n8158;
  assign n8160 = ~n7166 & ~n8159;
  assign n8161 = ~n3281 & ~n8160;
  assign n8162 = ~n3281 & ~n8161;
  assign n8163 = n3378 & ~n8162;
  assign n8164 = ~n4846 & ~n6860;
  assign n8165 = ~controllable_hmaster1 & ~n8164;
  assign n8166 = ~n6859 & ~n8165;
  assign n8167 = i_hbusreq3 & ~n8166;
  assign n8168 = ~n4852 & ~n6867;
  assign n8169 = ~controllable_hmaster1 & ~n8168;
  assign n8170 = ~n6866 & ~n8169;
  assign n8171 = ~i_hbusreq3 & ~n8170;
  assign n8172 = ~n8167 & ~n8171;
  assign n8173 = controllable_hmaster2 & ~n8172;
  assign n8174 = ~n6955 & ~n8173;
  assign n8175 = ~controllable_hgrant3 & ~n8174;
  assign n8176 = ~n7178 & ~n8175;
  assign n8177 = controllable_nhgrant0 & ~n8176;
  assign n8178 = ~n7208 & ~n8177;
  assign n8179 = ~n3281 & ~n8178;
  assign n8180 = ~n3281 & ~n8179;
  assign n8181 = ~n3378 & ~n8180;
  assign n8182 = ~n8163 & ~n8181;
  assign n8183 = n3492 & ~n8182;
  assign n8184 = n3492 & ~n8183;
  assign n8185 = n3485 & ~n8184;
  assign n8186 = n3485 & ~n8185;
  assign n8187 = ~n3476 & ~n8186;
  assign n8188 = ~n7752 & ~n8029;
  assign n8189 = ~controllable_hmaster0 & ~n8188;
  assign n8190 = ~n7250 & ~n8189;
  assign n8191 = ~controllable_hmaster1 & ~n8190;
  assign n8192 = ~n7249 & ~n8191;
  assign n8193 = i_hbusreq3 & ~n8192;
  assign n8194 = ~n7775 & ~n8036;
  assign n8195 = ~controllable_hmaster0 & ~n8194;
  assign n8196 = ~n7289 & ~n8195;
  assign n8197 = ~controllable_hmaster1 & ~n8196;
  assign n8198 = ~n7288 & ~n8197;
  assign n8199 = ~i_hbusreq3 & ~n8198;
  assign n8200 = ~n8193 & ~n8199;
  assign n8201 = controllable_hmaster2 & ~n8200;
  assign n8202 = ~n7389 & ~n8201;
  assign n8203 = ~controllable_hgrant3 & ~n8202;
  assign n8204 = ~n7240 & ~n8203;
  assign n8205 = controllable_nhgrant0 & ~n8204;
  assign n8206 = ~n7432 & ~n8205;
  assign n8207 = ~n3281 & ~n8206;
  assign n8208 = ~n3281 & ~n8207;
  assign n8209 = n3378 & ~n8208;
  assign n8210 = ~n6762 & ~n7796;
  assign n8211 = controllable_hmaster1 & ~n8210;
  assign n8212 = controllable_hmaster0 & ~n8210;
  assign n8213 = ~n7804 & ~n8056;
  assign n8214 = ~controllable_hmaster0 & ~n8213;
  assign n8215 = ~n8212 & ~n8214;
  assign n8216 = ~controllable_hmaster1 & ~n8215;
  assign n8217 = ~n8211 & ~n8216;
  assign n8218 = i_hbusreq3 & ~n8217;
  assign n8219 = ~n6772 & ~n7828;
  assign n8220 = controllable_hmaster1 & ~n8219;
  assign n8221 = controllable_hmaster0 & ~n8219;
  assign n8222 = ~n7849 & ~n8066;
  assign n8223 = ~controllable_hmaster0 & ~n8222;
  assign n8224 = ~n8221 & ~n8223;
  assign n8225 = ~controllable_hmaster1 & ~n8224;
  assign n8226 = ~n8220 & ~n8225;
  assign n8227 = ~i_hbusreq3 & ~n8226;
  assign n8228 = ~n8218 & ~n8227;
  assign n8229 = controllable_hmaster2 & ~n8228;
  assign n8230 = ~n6762 & ~n7861;
  assign n8231 = controllable_hmaster0 & ~n8230;
  assign n8232 = ~n6786 & ~n7861;
  assign n8233 = ~controllable_hmaster0 & ~n8232;
  assign n8234 = ~n8231 & ~n8233;
  assign n8235 = controllable_hmaster1 & ~n8234;
  assign n8236 = ~n6762 & ~n7872;
  assign n8237 = controllable_hmaster0 & ~n8236;
  assign n8238 = ~controllable_hmaster0 & ~n8230;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = ~controllable_hmaster1 & ~n8239;
  assign n8241 = ~n8235 & ~n8240;
  assign n8242 = i_hbusreq3 & ~n8241;
  assign n8243 = ~n6772 & ~n7895;
  assign n8244 = controllable_hmaster0 & ~n8243;
  assign n8245 = ~n6813 & ~n7895;
  assign n8246 = ~controllable_hmaster0 & ~n8245;
  assign n8247 = ~n8244 & ~n8246;
  assign n8248 = controllable_hmaster1 & ~n8247;
  assign n8249 = ~n6772 & ~n7920;
  assign n8250 = controllable_hmaster0 & ~n8249;
  assign n8251 = ~n6831 & ~n7934;
  assign n8252 = ~controllable_hmaster0 & ~n8251;
  assign n8253 = ~n8250 & ~n8252;
  assign n8254 = ~controllable_hmaster1 & ~n8253;
  assign n8255 = ~n8248 & ~n8254;
  assign n8256 = ~i_hbusreq3 & ~n8255;
  assign n8257 = ~n8242 & ~n8256;
  assign n8258 = ~controllable_hmaster2 & ~n8257;
  assign n8259 = ~n8229 & ~n8258;
  assign n8260 = ~controllable_hgrant3 & ~n8259;
  assign n8261 = ~n7457 & ~n8260;
  assign n8262 = controllable_nhgrant0 & ~n8261;
  assign n8263 = ~n7668 & ~n8262;
  assign n8264 = ~n3281 & ~n8263;
  assign n8265 = ~n3281 & ~n8264;
  assign n8266 = ~n3378 & ~n8265;
  assign n8267 = ~n8209 & ~n8266;
  assign n8268 = n3492 & ~n8267;
  assign n8269 = n3492 & ~n8268;
  assign n8270 = n3485 & ~n8269;
  assign n8271 = n3485 & ~n8270;
  assign n8272 = n3476 & ~n8271;
  assign n8273 = ~n8187 & ~n8272;
  assign n8274 = n3374 & ~n8273;
  assign n8275 = ~n8145 & ~n8274;
  assign n8276 = ~n3655 & ~n8275;
  assign n8277 = ~n8121 & ~n8276;
  assign n8278 = ~n3652 & ~n8277;
  assign n8279 = ~n7962 & ~n8278;
  assign n8280 = n3368 & ~n8279;
  assign n8281 = ~n7062 & ~n8280;
  assign n8282 = n3362 & ~n8281;
  assign n8283 = n3492 & ~n5248;
  assign n8284 = ~n3631 & ~n8283;
  assign n8285 = n3485 & ~n8284;
  assign n8286 = ~n3630 & ~n8285;
  assign n8287 = ~n3476 & ~n8286;
  assign n8288 = ~controllable_hmaster0 & ~n4944;
  assign n8289 = ~controllable_hmaster1 & ~n8288;
  assign n8290 = ~controllable_hmaster1 & ~n8289;
  assign n8291 = ~controllable_hmaster2 & ~n8290;
  assign n8292 = ~n3407 & ~n8291;
  assign n8293 = controllable_hgrant3 & ~n8292;
  assign n8294 = ~n3461 & ~n8291;
  assign n8295 = ~controllable_hgrant3 & ~n8294;
  assign n8296 = ~n8293 & ~n8295;
  assign n8297 = controllable_nhgrant0 & ~n8296;
  assign n8298 = ~controllable_hmaster0 & ~n5223;
  assign n8299 = ~controllable_hmaster1 & ~n8298;
  assign n8300 = ~controllable_hmaster1 & ~n8299;
  assign n8301 = ~controllable_hmaster2 & ~n8300;
  assign n8302 = ~n3407 & ~n8301;
  assign n8303 = ~controllable_hgrant3 & ~n8302;
  assign n8304 = ~n8293 & ~n8303;
  assign n8305 = ~controllable_nhgrant0 & ~n8304;
  assign n8306 = ~n8297 & ~n8305;
  assign n8307 = ~n3281 & ~n8306;
  assign n8308 = ~n3783 & ~n8307;
  assign n8309 = ~n3492 & ~n8308;
  assign n8310 = ~n3467 & n3492;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = ~n3485 & ~n8311;
  assign n8313 = ~n8285 & ~n8312;
  assign n8314 = n3476 & ~n8313;
  assign n8315 = ~n8287 & ~n8314;
  assign n8316 = ~n3374 & ~n8315;
  assign n8317 = n3492 & ~n5537;
  assign n8318 = ~n3631 & ~n8317;
  assign n8319 = n3485 & ~n8318;
  assign n8320 = ~n3630 & ~n8319;
  assign n8321 = ~n3476 & ~n8320;
  assign n8322 = n3492 & ~n6085;
  assign n8323 = ~n3631 & ~n8322;
  assign n8324 = n3485 & ~n8323;
  assign n8325 = ~n8312 & ~n8324;
  assign n8326 = n3476 & ~n8325;
  assign n8327 = ~n8321 & ~n8326;
  assign n8328 = n3374 & ~n8327;
  assign n8329 = ~n8316 & ~n8328;
  assign n8330 = n3655 & ~n8329;
  assign n8331 = n3492 & ~n6195;
  assign n8332 = ~n3631 & ~n8331;
  assign n8333 = n3485 & ~n8332;
  assign n8334 = ~n3630 & ~n8333;
  assign n8335 = ~n3476 & ~n8334;
  assign n8336 = ~controllable_hmaster1 & ~n4946;
  assign n8337 = i_hbusreq3 & ~n8336;
  assign n8338 = ~controllable_hmaster1 & ~n5009;
  assign n8339 = ~i_hbusreq3 & ~n8338;
  assign n8340 = ~n8337 & ~n8339;
  assign n8341 = ~controllable_hmaster2 & ~n8340;
  assign n8342 = ~n3407 & ~n8341;
  assign n8343 = controllable_hgrant3 & ~n8342;
  assign n8344 = ~controllable_hmaster1 & ~n6151;
  assign n8345 = i_hbusreq3 & ~n8344;
  assign n8346 = ~controllable_hmaster1 & ~n6180;
  assign n8347 = ~i_hbusreq3 & ~n8346;
  assign n8348 = ~n8345 & ~n8347;
  assign n8349 = ~controllable_hmaster2 & ~n8348;
  assign n8350 = ~n3461 & ~n8349;
  assign n8351 = ~controllable_hgrant3 & ~n8350;
  assign n8352 = ~n8343 & ~n8351;
  assign n8353 = controllable_nhgrant0 & ~n8352;
  assign n8354 = ~controllable_hmaster1 & ~n5225;
  assign n8355 = i_hbusreq3 & ~n8354;
  assign n8356 = ~controllable_hmaster1 & ~n5233;
  assign n8357 = ~i_hbusreq3 & ~n8356;
  assign n8358 = ~n8355 & ~n8357;
  assign n8359 = ~controllable_hmaster2 & ~n8358;
  assign n8360 = ~n3407 & ~n8359;
  assign n8361 = ~controllable_hgrant3 & ~n8360;
  assign n8362 = ~n8343 & ~n8361;
  assign n8363 = ~controllable_nhgrant0 & ~n8362;
  assign n8364 = ~n8353 & ~n8363;
  assign n8365 = ~n3281 & ~n8364;
  assign n8366 = ~n3783 & ~n8365;
  assign n8367 = ~n3492 & ~n8366;
  assign n8368 = ~n8310 & ~n8367;
  assign n8369 = ~n3485 & ~n8368;
  assign n8370 = ~n8333 & ~n8369;
  assign n8371 = n3476 & ~n8370;
  assign n8372 = ~n8335 & ~n8371;
  assign n8373 = ~n3374 & ~n8372;
  assign n8374 = n3492 & ~n6350;
  assign n8375 = ~n3631 & ~n8374;
  assign n8376 = n3485 & ~n8375;
  assign n8377 = ~n3630 & ~n8376;
  assign n8378 = ~n3476 & ~n8377;
  assign n8379 = n3492 & ~n6561;
  assign n8380 = ~n3631 & ~n8379;
  assign n8381 = n3485 & ~n8380;
  assign n8382 = ~n8369 & ~n8381;
  assign n8383 = n3476 & ~n8382;
  assign n8384 = ~n8378 & ~n8383;
  assign n8385 = n3374 & ~n8384;
  assign n8386 = ~n8373 & ~n8385;
  assign n8387 = ~n3655 & ~n8386;
  assign n8388 = ~n8330 & ~n8387;
  assign n8389 = n3652 & ~n8388;
  assign n8390 = n3492 & ~n6664;
  assign n8391 = ~n3631 & ~n8390;
  assign n8392 = n3485 & ~n8391;
  assign n8393 = ~n3630 & ~n8392;
  assign n8394 = ~n3476 & ~n8393;
  assign n8395 = ~controllable_hmaster0 & ~n4930;
  assign n8396 = controllable_hmaster1 & ~n8395;
  assign n8397 = ~n8289 & ~n8396;
  assign n8398 = i_hbusreq3 & ~n8397;
  assign n8399 = ~controllable_hmaster0 & ~n4990;
  assign n8400 = controllable_hmaster1 & ~n8399;
  assign n8401 = ~n8289 & ~n8400;
  assign n8402 = ~i_hbusreq3 & ~n8401;
  assign n8403 = ~n8398 & ~n8402;
  assign n8404 = ~controllable_hmaster2 & ~n8403;
  assign n8405 = ~n3407 & ~n8404;
  assign n8406 = controllable_hgrant3 & ~n8405;
  assign n8407 = ~controllable_hmaster0 & ~n6600;
  assign n8408 = controllable_hmaster1 & ~n8407;
  assign n8409 = ~n8289 & ~n8408;
  assign n8410 = i_hbusreq3 & ~n8409;
  assign n8411 = ~controllable_hmaster0 & ~n6645;
  assign n8412 = controllable_hmaster1 & ~n8411;
  assign n8413 = ~n8289 & ~n8412;
  assign n8414 = ~i_hbusreq3 & ~n8413;
  assign n8415 = ~n8410 & ~n8414;
  assign n8416 = ~controllable_hmaster2 & ~n8415;
  assign n8417 = ~n3461 & ~n8416;
  assign n8418 = ~controllable_hgrant3 & ~n8417;
  assign n8419 = ~n8406 & ~n8418;
  assign n8420 = controllable_nhgrant0 & ~n8419;
  assign n8421 = ~n8299 & ~n8396;
  assign n8422 = i_hbusreq3 & ~n8421;
  assign n8423 = ~n8299 & ~n8400;
  assign n8424 = ~i_hbusreq3 & ~n8423;
  assign n8425 = ~n8422 & ~n8424;
  assign n8426 = ~controllable_hmaster2 & ~n8425;
  assign n8427 = ~n3407 & ~n8426;
  assign n8428 = ~controllable_hgrant3 & ~n8427;
  assign n8429 = ~n8406 & ~n8428;
  assign n8430 = ~controllable_nhgrant0 & ~n8429;
  assign n8431 = ~n8420 & ~n8430;
  assign n8432 = ~n3281 & ~n8431;
  assign n8433 = ~n3783 & ~n8432;
  assign n8434 = ~n3492 & ~n8433;
  assign n8435 = ~n8310 & ~n8434;
  assign n8436 = ~n3485 & ~n8435;
  assign n8437 = ~n8392 & ~n8436;
  assign n8438 = n3476 & ~n8437;
  assign n8439 = ~n8394 & ~n8438;
  assign n8440 = ~n3374 & ~n8439;
  assign n8441 = n3492 & ~n6730;
  assign n8442 = ~n3631 & ~n8441;
  assign n8443 = n3485 & ~n8442;
  assign n8444 = ~n3630 & ~n8443;
  assign n8445 = ~n3476 & ~n8444;
  assign n8446 = n3492 & ~n6846;
  assign n8447 = ~n3631 & ~n8446;
  assign n8448 = n3485 & ~n8447;
  assign n8449 = ~n8436 & ~n8448;
  assign n8450 = n3476 & ~n8449;
  assign n8451 = ~n8445 & ~n8450;
  assign n8452 = n3374 & ~n8451;
  assign n8453 = ~n8440 & ~n8452;
  assign n8454 = n3655 & ~n8453;
  assign n8455 = n3492 & ~n6894;
  assign n8456 = ~n3631 & ~n8455;
  assign n8457 = n3485 & ~n8456;
  assign n8458 = ~n3630 & ~n8457;
  assign n8459 = ~n3476 & ~n8458;
  assign n8460 = ~n4946 & ~n8396;
  assign n8461 = i_hbusreq3 & ~n8460;
  assign n8462 = ~n5009 & ~n8400;
  assign n8463 = ~i_hbusreq3 & ~n8462;
  assign n8464 = ~n8461 & ~n8463;
  assign n8465 = ~controllable_hmaster2 & ~n8464;
  assign n8466 = ~n3407 & ~n8465;
  assign n8467 = controllable_hgrant3 & ~n8466;
  assign n8468 = ~n6151 & ~n8408;
  assign n8469 = i_hbusreq3 & ~n8468;
  assign n8470 = ~n6180 & ~n8412;
  assign n8471 = ~i_hbusreq3 & ~n8470;
  assign n8472 = ~n8469 & ~n8471;
  assign n8473 = ~controllable_hmaster2 & ~n8472;
  assign n8474 = ~n3461 & ~n8473;
  assign n8475 = ~controllable_hgrant3 & ~n8474;
  assign n8476 = ~n8467 & ~n8475;
  assign n8477 = controllable_nhgrant0 & ~n8476;
  assign n8478 = ~n5225 & ~n8396;
  assign n8479 = i_hbusreq3 & ~n8478;
  assign n8480 = ~n5233 & ~n8400;
  assign n8481 = ~i_hbusreq3 & ~n8480;
  assign n8482 = ~n8479 & ~n8481;
  assign n8483 = ~controllable_hmaster2 & ~n8482;
  assign n8484 = ~n3407 & ~n8483;
  assign n8485 = ~controllable_hgrant3 & ~n8484;
  assign n8486 = ~n8467 & ~n8485;
  assign n8487 = ~controllable_nhgrant0 & ~n8486;
  assign n8488 = ~n8477 & ~n8487;
  assign n8489 = ~n3281 & ~n8488;
  assign n8490 = ~n3783 & ~n8489;
  assign n8491 = ~n3492 & ~n8490;
  assign n8492 = ~n8310 & ~n8491;
  assign n8493 = ~n3485 & ~n8492;
  assign n8494 = ~n8457 & ~n8493;
  assign n8495 = n3476 & ~n8494;
  assign n8496 = ~n8459 & ~n8495;
  assign n8497 = ~n3374 & ~n8496;
  assign n8498 = n3492 & ~n6962;
  assign n8499 = ~n3631 & ~n8498;
  assign n8500 = n3485 & ~n8499;
  assign n8501 = ~n3630 & ~n8500;
  assign n8502 = ~n3476 & ~n8501;
  assign n8503 = n3492 & ~n7047;
  assign n8504 = ~n3631 & ~n8503;
  assign n8505 = n3485 & ~n8504;
  assign n8506 = ~n8493 & ~n8505;
  assign n8507 = n3476 & ~n8506;
  assign n8508 = ~n8502 & ~n8507;
  assign n8509 = n3374 & ~n8508;
  assign n8510 = ~n8497 & ~n8509;
  assign n8511 = ~n3655 & ~n8510;
  assign n8512 = ~n8454 & ~n8511;
  assign n8513 = ~n3652 & ~n8512;
  assign n8514 = ~n8389 & ~n8513;
  assign n8515 = ~n3368 & ~n8514;
  assign n8516 = n3492 & ~n7121;
  assign n8517 = n3492 & ~n8516;
  assign n8518 = n3485 & ~n8517;
  assign n8519 = n3485 & ~n8518;
  assign n8520 = ~n3476 & ~n8519;
  assign n8521 = ~n3281 & ~n3467;
  assign n8522 = ~n3281 & ~n8521;
  assign n8523 = ~n3492 & ~n8522;
  assign n8524 = ~n3492 & ~n8523;
  assign n8525 = ~n3485 & ~n8524;
  assign n8526 = ~n8518 & ~n8525;
  assign n8527 = n3476 & ~n8526;
  assign n8528 = ~n8520 & ~n8527;
  assign n8529 = ~n3374 & ~n8528;
  assign n8530 = n3492 & ~n7211;
  assign n8531 = n3492 & ~n8530;
  assign n8532 = n3485 & ~n8531;
  assign n8533 = n3485 & ~n8532;
  assign n8534 = ~n3476 & ~n8533;
  assign n8535 = ~n3281 & ~n8307;
  assign n8536 = ~n3492 & ~n8535;
  assign n8537 = ~n3492 & ~n8536;
  assign n8538 = ~n3485 & ~n8537;
  assign n8539 = n3492 & ~n7671;
  assign n8540 = n3492 & ~n8539;
  assign n8541 = n3485 & ~n8540;
  assign n8542 = ~n8538 & ~n8541;
  assign n8543 = n3476 & ~n8542;
  assign n8544 = ~n8534 & ~n8543;
  assign n8545 = n3374 & ~n8544;
  assign n8546 = ~n8529 & ~n8545;
  assign n8547 = n3655 & ~n8546;
  assign n8548 = n3492 & ~n7699;
  assign n8549 = n3492 & ~n8548;
  assign n8550 = n3485 & ~n8549;
  assign n8551 = n3485 & ~n8550;
  assign n8552 = ~n3476 & ~n8551;
  assign n8553 = ~n8525 & ~n8550;
  assign n8554 = n3476 & ~n8553;
  assign n8555 = ~n8552 & ~n8554;
  assign n8556 = ~n3374 & ~n8555;
  assign n8557 = n3492 & ~n7741;
  assign n8558 = n3492 & ~n8557;
  assign n8559 = n3485 & ~n8558;
  assign n8560 = n3485 & ~n8559;
  assign n8561 = ~n3476 & ~n8560;
  assign n8562 = ~n3281 & ~n8365;
  assign n8563 = ~n3492 & ~n8562;
  assign n8564 = ~n3492 & ~n8563;
  assign n8565 = ~n3485 & ~n8564;
  assign n8566 = n3492 & ~n7949;
  assign n8567 = n3492 & ~n8566;
  assign n8568 = n3485 & ~n8567;
  assign n8569 = ~n8565 & ~n8568;
  assign n8570 = n3476 & ~n8569;
  assign n8571 = ~n8561 & ~n8570;
  assign n8572 = n3374 & ~n8571;
  assign n8573 = ~n8556 & ~n8572;
  assign n8574 = ~n3655 & ~n8573;
  assign n8575 = ~n8547 & ~n8574;
  assign n8576 = n3652 & ~n8575;
  assign n8577 = n3492 & ~n7979;
  assign n8578 = n3492 & ~n8577;
  assign n8579 = n3485 & ~n8578;
  assign n8580 = n3485 & ~n8579;
  assign n8581 = ~n3476 & ~n8580;
  assign n8582 = ~n8525 & ~n8579;
  assign n8583 = n3476 & ~n8582;
  assign n8584 = ~n8581 & ~n8583;
  assign n8585 = ~n3374 & ~n8584;
  assign n8586 = n3492 & ~n8021;
  assign n8587 = n3492 & ~n8586;
  assign n8588 = n3485 & ~n8587;
  assign n8589 = n3485 & ~n8588;
  assign n8590 = ~n3476 & ~n8589;
  assign n8591 = ~n3281 & ~n8432;
  assign n8592 = ~n3492 & ~n8591;
  assign n8593 = ~n3492 & ~n8592;
  assign n8594 = ~n3485 & ~n8593;
  assign n8595 = n3492 & ~n8110;
  assign n8596 = n3492 & ~n8595;
  assign n8597 = n3485 & ~n8596;
  assign n8598 = ~n8594 & ~n8597;
  assign n8599 = n3476 & ~n8598;
  assign n8600 = ~n8590 & ~n8599;
  assign n8601 = n3374 & ~n8600;
  assign n8602 = ~n8585 & ~n8601;
  assign n8603 = n3655 & ~n8602;
  assign n8604 = n3492 & ~n8138;
  assign n8605 = n3492 & ~n8604;
  assign n8606 = n3485 & ~n8605;
  assign n8607 = n3485 & ~n8606;
  assign n8608 = ~n3476 & ~n8607;
  assign n8609 = ~n8525 & ~n8606;
  assign n8610 = n3476 & ~n8609;
  assign n8611 = ~n8608 & ~n8610;
  assign n8612 = ~n3374 & ~n8611;
  assign n8613 = n3492 & ~n8180;
  assign n8614 = n3492 & ~n8613;
  assign n8615 = n3485 & ~n8614;
  assign n8616 = n3485 & ~n8615;
  assign n8617 = ~n3476 & ~n8616;
  assign n8618 = ~n3281 & ~n8489;
  assign n8619 = ~n3492 & ~n8618;
  assign n8620 = ~n3492 & ~n8619;
  assign n8621 = ~n3485 & ~n8620;
  assign n8622 = n3492 & ~n8265;
  assign n8623 = n3492 & ~n8622;
  assign n8624 = n3485 & ~n8623;
  assign n8625 = ~n8621 & ~n8624;
  assign n8626 = n3476 & ~n8625;
  assign n8627 = ~n8617 & ~n8626;
  assign n8628 = n3374 & ~n8627;
  assign n8629 = ~n8612 & ~n8628;
  assign n8630 = ~n3655 & ~n8629;
  assign n8631 = ~n8603 & ~n8630;
  assign n8632 = ~n3652 & ~n8631;
  assign n8633 = ~n8576 & ~n8632;
  assign n8634 = n3368 & ~n8633;
  assign n8635 = ~n8515 & ~n8634;
  assign n8636 = ~n3362 & ~n8635;
  assign n8637 = ~n8282 & ~n8636;
  assign n8638 = n3359 & ~n8637;
  assign n8639 = ~n3485 & ~n8308;
  assign n8640 = ~n8285 & ~n8639;
  assign n8641 = n3476 & ~n8640;
  assign n8642 = ~n8287 & ~n8641;
  assign n8643 = ~n3374 & ~n8642;
  assign n8644 = ~n8324 & ~n8639;
  assign n8645 = n3476 & ~n8644;
  assign n8646 = ~n8321 & ~n8645;
  assign n8647 = n3374 & ~n8646;
  assign n8648 = ~n8643 & ~n8647;
  assign n8649 = n3655 & ~n8648;
  assign n8650 = ~n3485 & ~n8366;
  assign n8651 = ~n8333 & ~n8650;
  assign n8652 = n3476 & ~n8651;
  assign n8653 = ~n8335 & ~n8652;
  assign n8654 = ~n3374 & ~n8653;
  assign n8655 = ~n8381 & ~n8650;
  assign n8656 = n3476 & ~n8655;
  assign n8657 = ~n8378 & ~n8656;
  assign n8658 = n3374 & ~n8657;
  assign n8659 = ~n8654 & ~n8658;
  assign n8660 = ~n3655 & ~n8659;
  assign n8661 = ~n8649 & ~n8660;
  assign n8662 = n3652 & ~n8661;
  assign n8663 = ~n3485 & ~n8433;
  assign n8664 = ~n8392 & ~n8663;
  assign n8665 = n3476 & ~n8664;
  assign n8666 = ~n8394 & ~n8665;
  assign n8667 = ~n3374 & ~n8666;
  assign n8668 = ~n8448 & ~n8663;
  assign n8669 = n3476 & ~n8668;
  assign n8670 = ~n8445 & ~n8669;
  assign n8671 = n3374 & ~n8670;
  assign n8672 = ~n8667 & ~n8671;
  assign n8673 = n3655 & ~n8672;
  assign n8674 = ~n3485 & ~n8490;
  assign n8675 = ~n8457 & ~n8674;
  assign n8676 = n3476 & ~n8675;
  assign n8677 = ~n8459 & ~n8676;
  assign n8678 = ~n3374 & ~n8677;
  assign n8679 = ~n8505 & ~n8674;
  assign n8680 = n3476 & ~n8679;
  assign n8681 = ~n8502 & ~n8680;
  assign n8682 = n3374 & ~n8681;
  assign n8683 = ~n8678 & ~n8682;
  assign n8684 = ~n3655 & ~n8683;
  assign n8685 = ~n8673 & ~n8684;
  assign n8686 = ~n3652 & ~n8685;
  assign n8687 = ~n8662 & ~n8686;
  assign n8688 = ~n3368 & ~n8687;
  assign n8689 = ~n3485 & ~n8522;
  assign n8690 = ~n8518 & ~n8689;
  assign n8691 = n3476 & ~n8690;
  assign n8692 = ~n8520 & ~n8691;
  assign n8693 = ~n3374 & ~n8692;
  assign n8694 = ~n3485 & ~n8535;
  assign n8695 = ~n8541 & ~n8694;
  assign n8696 = n3476 & ~n8695;
  assign n8697 = ~n8534 & ~n8696;
  assign n8698 = n3374 & ~n8697;
  assign n8699 = ~n8693 & ~n8698;
  assign n8700 = n3655 & ~n8699;
  assign n8701 = ~n8550 & ~n8689;
  assign n8702 = n3476 & ~n8701;
  assign n8703 = ~n8552 & ~n8702;
  assign n8704 = ~n3374 & ~n8703;
  assign n8705 = ~n3485 & ~n8562;
  assign n8706 = ~n8568 & ~n8705;
  assign n8707 = n3476 & ~n8706;
  assign n8708 = ~n8561 & ~n8707;
  assign n8709 = n3374 & ~n8708;
  assign n8710 = ~n8704 & ~n8709;
  assign n8711 = ~n3655 & ~n8710;
  assign n8712 = ~n8700 & ~n8711;
  assign n8713 = n3652 & ~n8712;
  assign n8714 = ~n8579 & ~n8689;
  assign n8715 = n3476 & ~n8714;
  assign n8716 = ~n8581 & ~n8715;
  assign n8717 = ~n3374 & ~n8716;
  assign n8718 = ~n3485 & ~n8591;
  assign n8719 = ~n8597 & ~n8718;
  assign n8720 = n3476 & ~n8719;
  assign n8721 = ~n8590 & ~n8720;
  assign n8722 = n3374 & ~n8721;
  assign n8723 = ~n8717 & ~n8722;
  assign n8724 = n3655 & ~n8723;
  assign n8725 = ~n8606 & ~n8689;
  assign n8726 = n3476 & ~n8725;
  assign n8727 = ~n8608 & ~n8726;
  assign n8728 = ~n3374 & ~n8727;
  assign n8729 = ~n3485 & ~n8618;
  assign n8730 = ~n8624 & ~n8729;
  assign n8731 = n3476 & ~n8730;
  assign n8732 = ~n8617 & ~n8731;
  assign n8733 = n3374 & ~n8732;
  assign n8734 = ~n8728 & ~n8733;
  assign n8735 = ~n3655 & ~n8734;
  assign n8736 = ~n8724 & ~n8735;
  assign n8737 = ~n3652 & ~n8736;
  assign n8738 = ~n8713 & ~n8737;
  assign n8739 = n3368 & ~n8738;
  assign n8740 = ~n8688 & ~n8739;
  assign n8741 = n3362 & ~n8740;
  assign n8742 = n3378 & ~n5248;
  assign n8743 = ~n3382 & ~n3697;
  assign n8744 = ~controllable_hmaster1 & ~n8743;
  assign n8745 = ~n3381 & ~n8744;
  assign n8746 = ~i_hbusreq3 & ~n8745;
  assign n8747 = ~n3787 & ~n8746;
  assign n8748 = controllable_hmaster2 & ~n8747;
  assign n8749 = ~n5035 & ~n8748;
  assign n8750 = controllable_hgrant3 & ~n8749;
  assign n8751 = ~n3502 & ~n3729;
  assign n8752 = ~controllable_hmaster1 & ~n8751;
  assign n8753 = ~n3501 & ~n8752;
  assign n8754 = i_hbusreq3 & ~n8753;
  assign n8755 = ~n3502 & ~n3767;
  assign n8756 = ~controllable_hmaster1 & ~n8755;
  assign n8757 = ~n3501 & ~n8756;
  assign n8758 = ~i_hbusreq3 & ~n8757;
  assign n8759 = ~n8754 & ~n8758;
  assign n8760 = controllable_hmaster2 & ~n8759;
  assign n8761 = ~n5161 & ~n8760;
  assign n8762 = ~controllable_hgrant3 & ~n8761;
  assign n8763 = ~n8750 & ~n8762;
  assign n8764 = controllable_nhgrant0 & ~n8763;
  assign n8765 = ~n5187 & ~n8748;
  assign n8766 = controllable_hgrant3 & ~n8765;
  assign n8767 = ~n3411 & ~n3850;
  assign n8768 = ~controllable_hgrant2 & ~n8767;
  assign n8769 = ~n3410 & ~n8768;
  assign n8770 = controllable_hmaster1 & ~n8769;
  assign n8771 = controllable_hmaster0 & ~n8769;
  assign n8772 = ~n3667 & ~n8771;
  assign n8773 = ~controllable_hmaster1 & ~n8772;
  assign n8774 = ~n8770 & ~n8773;
  assign n8775 = i_hbusreq3 & ~n8774;
  assign n8776 = ~n3697 & ~n8771;
  assign n8777 = ~controllable_hmaster1 & ~n8776;
  assign n8778 = ~n8770 & ~n8777;
  assign n8779 = ~i_hbusreq3 & ~n8778;
  assign n8780 = ~n8775 & ~n8779;
  assign n8781 = controllable_hmaster2 & ~n8780;
  assign n8782 = ~n5241 & ~n8781;
  assign n8783 = ~controllable_hgrant3 & ~n8782;
  assign n8784 = ~n8766 & ~n8783;
  assign n8785 = ~controllable_nhgrant0 & ~n8784;
  assign n8786 = ~n8764 & ~n8785;
  assign n8787 = ~n3281 & ~n8786;
  assign n8788 = ~n3783 & ~n8787;
  assign n8789 = ~n3378 & ~n8788;
  assign n8790 = ~n8742 & ~n8789;
  assign n8791 = n3492 & ~n8790;
  assign n8792 = ~n3631 & ~n8791;
  assign n8793 = n3485 & ~n8792;
  assign n8794 = ~n3630 & ~n8793;
  assign n8795 = ~n3476 & ~n8794;
  assign n8796 = ~n8309 & ~n8791;
  assign n8797 = n3485 & ~n8796;
  assign n8798 = ~n8639 & ~n8797;
  assign n8799 = n3476 & ~n8798;
  assign n8800 = ~n8795 & ~n8799;
  assign n8801 = ~n3374 & ~n8800;
  assign n8802 = n3378 & ~n5537;
  assign n8803 = ~n3382 & ~n3835;
  assign n8804 = ~controllable_hmaster1 & ~n8803;
  assign n8805 = ~n3381 & ~n8804;
  assign n8806 = ~i_hbusreq3 & ~n8805;
  assign n8807 = ~n3951 & ~n8806;
  assign n8808 = controllable_hmaster2 & ~n8807;
  assign n8809 = ~n5400 & ~n8808;
  assign n8810 = controllable_hgrant3 & ~n8809;
  assign n8811 = ~n3502 & ~n3890;
  assign n8812 = ~controllable_hmaster1 & ~n8811;
  assign n8813 = ~n3501 & ~n8812;
  assign n8814 = ~i_hbusreq3 & ~n8813;
  assign n8815 = ~n3963 & ~n8814;
  assign n8816 = controllable_hmaster2 & ~n8815;
  assign n8817 = ~n5288 & ~n8768;
  assign n8818 = ~controllable_hmaster0 & ~n8817;
  assign n8819 = ~n8771 & ~n8818;
  assign n8820 = controllable_hmaster1 & ~n8819;
  assign n8821 = ~n3495 & ~n5297;
  assign n8822 = ~controllable_hgrant4 & ~n8821;
  assign n8823 = ~n3411 & ~n8822;
  assign n8824 = ~controllable_hgrant2 & ~n8823;
  assign n8825 = ~n3410 & ~n8824;
  assign n8826 = controllable_hmaster0 & ~n8825;
  assign n8827 = ~controllable_hmaster0 & ~n8769;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = ~controllable_hmaster1 & ~n8828;
  assign n8830 = ~n8820 & ~n8829;
  assign n8831 = i_hbusreq3 & ~n8830;
  assign n8832 = i_hbusreq2 & ~n8767;
  assign n8833 = ~n3884 & ~n3916;
  assign n8834 = ~i_hbusreq2 & ~n8833;
  assign n8835 = ~n8832 & ~n8834;
  assign n8836 = ~controllable_hgrant2 & ~n8835;
  assign n8837 = ~n3859 & ~n8836;
  assign n8838 = controllable_hmaster0 & ~n8837;
  assign n8839 = ~n5438 & ~n8836;
  assign n8840 = ~controllable_hmaster0 & ~n8839;
  assign n8841 = ~n8838 & ~n8840;
  assign n8842 = controllable_hmaster1 & ~n8841;
  assign n8843 = i_hbusreq2 & ~n8823;
  assign n8844 = i_hbusreq4 & ~n8821;
  assign n8845 = i_hbusreq0 & ~n8821;
  assign n8846 = ~n3511 & ~n5320;
  assign n8847 = i_hlock0 & ~n8846;
  assign n8848 = ~i_hlock0 & ~n8821;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~i_hbusreq0 & ~n8849;
  assign n8851 = ~n8845 & ~n8850;
  assign n8852 = ~i_hbusreq4 & ~n8851;
  assign n8853 = ~n8844 & ~n8852;
  assign n8854 = ~controllable_hgrant4 & ~n8853;
  assign n8855 = ~n3916 & ~n8854;
  assign n8856 = ~i_hbusreq2 & ~n8855;
  assign n8857 = ~n8843 & ~n8856;
  assign n8858 = ~controllable_hgrant2 & ~n8857;
  assign n8859 = ~n3859 & ~n8858;
  assign n8860 = controllable_hmaster0 & ~n8859;
  assign n8861 = ~n3494 & ~n5382;
  assign n8862 = ~i_hready & ~n8861;
  assign n8863 = ~i_hready & ~n8862;
  assign n8864 = i_hlock0 & ~n8863;
  assign n8865 = ~n3878 & ~n8864;
  assign n8866 = ~i_hbusreq0 & ~n8865;
  assign n8867 = ~n3875 & ~n8866;
  assign n8868 = ~i_hbusreq4 & ~n8867;
  assign n8869 = ~n3874 & ~n8868;
  assign n8870 = ~controllable_hgrant4 & ~n8869;
  assign n8871 = ~n5462 & ~n8870;
  assign n8872 = ~i_hbusreq2 & ~n8871;
  assign n8873 = ~n8832 & ~n8872;
  assign n8874 = ~controllable_hgrant2 & ~n8873;
  assign n8875 = ~n5461 & ~n8874;
  assign n8876 = ~controllable_hmaster0 & ~n8875;
  assign n8877 = ~n8860 & ~n8876;
  assign n8878 = ~controllable_hmaster1 & ~n8877;
  assign n8879 = ~n8842 & ~n8878;
  assign n8880 = ~i_hbusreq3 & ~n8879;
  assign n8881 = ~n8831 & ~n8880;
  assign n8882 = ~controllable_hmaster2 & ~n8881;
  assign n8883 = ~n8816 & ~n8882;
  assign n8884 = ~controllable_hgrant3 & ~n8883;
  assign n8885 = ~n8810 & ~n8884;
  assign n8886 = controllable_nhgrant0 & ~n8885;
  assign n8887 = ~n5492 & ~n8808;
  assign n8888 = controllable_hgrant3 & ~n8887;
  assign n8889 = ~n3910 & ~n8771;
  assign n8890 = ~controllable_hmaster1 & ~n8889;
  assign n8891 = ~n8770 & ~n8890;
  assign n8892 = i_hbusreq3 & ~n8891;
  assign n8893 = ~n3935 & ~n8771;
  assign n8894 = ~controllable_hmaster1 & ~n8893;
  assign n8895 = ~n8770 & ~n8894;
  assign n8896 = ~i_hbusreq3 & ~n8895;
  assign n8897 = ~n8892 & ~n8896;
  assign n8898 = controllable_hmaster2 & ~n8897;
  assign n8899 = ~n5530 & ~n8898;
  assign n8900 = ~controllable_hgrant3 & ~n8899;
  assign n8901 = ~n8888 & ~n8900;
  assign n8902 = ~controllable_nhgrant0 & ~n8901;
  assign n8903 = ~n8886 & ~n8902;
  assign n8904 = ~n3281 & ~n8903;
  assign n8905 = ~n3950 & ~n8904;
  assign n8906 = ~n3378 & ~n8905;
  assign n8907 = ~n8802 & ~n8906;
  assign n8908 = n3492 & ~n8907;
  assign n8909 = ~n3631 & ~n8908;
  assign n8910 = n3485 & ~n8909;
  assign n8911 = ~n3630 & ~n8910;
  assign n8912 = ~n3476 & ~n8911;
  assign n8913 = n3378 & ~n6085;
  assign n8914 = i_hlock0 & ~n5563;
  assign n8915 = ~n5814 & ~n8914;
  assign n8916 = ~i_hbusreq0 & ~n8915;
  assign n8917 = ~n4107 & ~n8916;
  assign n8918 = ~i_hbusreq4 & ~n8917;
  assign n8919 = ~n4106 & ~n8918;
  assign n8920 = ~controllable_hgrant4 & ~n8919;
  assign n8921 = ~n3411 & ~n8920;
  assign n8922 = ~i_hbusreq2 & ~n8921;
  assign n8923 = ~n5550 & ~n8922;
  assign n8924 = ~controllable_hgrant2 & ~n8923;
  assign n8925 = ~n3410 & ~n8924;
  assign n8926 = controllable_hmaster1 & ~n8925;
  assign n8927 = controllable_hmaster0 & ~n8925;
  assign n8928 = ~n5836 & ~n8927;
  assign n8929 = ~controllable_hmaster1 & ~n8928;
  assign n8930 = ~n8926 & ~n8929;
  assign n8931 = ~i_hbusreq3 & ~n8930;
  assign n8932 = ~n5549 & ~n8931;
  assign n8933 = controllable_hmaster2 & ~n8932;
  assign n8934 = ~n5859 & ~n8933;
  assign n8935 = controllable_hgrant3 & ~n8934;
  assign n8936 = controllable_hgrant2 & ~n8923;
  assign n8937 = controllable_hgrant4 & ~n8919;
  assign n8938 = ~i_hbusreq1 & ~n4010;
  assign n8939 = ~n5639 & ~n8938;
  assign n8940 = ~controllable_ndecide & ~n8939;
  assign n8941 = ~n3494 & ~n8940;
  assign n8942 = i_hready & ~n8941;
  assign n8943 = ~n3495 & ~n8942;
  assign n8944 = i_hlock0 & ~n8943;
  assign n8945 = ~n5871 & ~n8944;
  assign n8946 = ~i_hbusreq0 & ~n8945;
  assign n8947 = ~n5638 & ~n8946;
  assign n8948 = ~i_hbusreq4 & ~n8947;
  assign n8949 = ~n5637 & ~n8948;
  assign n8950 = ~controllable_hgrant4 & ~n8949;
  assign n8951 = ~n8937 & ~n8950;
  assign n8952 = ~i_hbusreq2 & ~n8951;
  assign n8953 = ~n5636 & ~n8952;
  assign n8954 = ~controllable_hgrant2 & ~n8953;
  assign n8955 = ~n8936 & ~n8954;
  assign n8956 = controllable_hmaster1 & ~n8955;
  assign n8957 = controllable_hmaster0 & ~n8955;
  assign n8958 = ~n4655 & ~n5639;
  assign n8959 = ~controllable_ndecide & ~n8958;
  assign n8960 = ~n3494 & ~n8959;
  assign n8961 = i_hready & ~n8960;
  assign n8962 = ~n3511 & ~n8961;
  assign n8963 = i_hlock0 & ~n8962;
  assign n8964 = ~n5891 & ~n8963;
  assign n8965 = ~i_hbusreq0 & ~n8964;
  assign n8966 = ~n5638 & ~n8965;
  assign n8967 = ~i_hbusreq4 & ~n8966;
  assign n8968 = ~n5637 & ~n8967;
  assign n8969 = ~controllable_hgrant4 & ~n8968;
  assign n8970 = ~n4064 & ~n8969;
  assign n8971 = ~i_hbusreq2 & ~n8970;
  assign n8972 = ~n5658 & ~n8971;
  assign n8973 = ~controllable_hgrant2 & ~n8972;
  assign n8974 = ~n5862 & ~n8973;
  assign n8975 = ~controllable_hmaster0 & ~n8974;
  assign n8976 = ~n8957 & ~n8975;
  assign n8977 = ~controllable_hmaster1 & ~n8976;
  assign n8978 = ~n8956 & ~n8977;
  assign n8979 = ~i_hbusreq3 & ~n8978;
  assign n8980 = ~n5634 & ~n8979;
  assign n8981 = controllable_hmaster2 & ~n8980;
  assign n8982 = ~n5623 & ~n5686;
  assign n8983 = ~controllable_hmaster0 & ~n8982;
  assign n8984 = ~n5626 & ~n8983;
  assign n8985 = controllable_hmaster1 & ~n8984;
  assign n8986 = ~n3495 & ~n5695;
  assign n8987 = ~controllable_hgrant4 & ~n8986;
  assign n8988 = ~n4091 & ~n8987;
  assign n8989 = ~controllable_hgrant2 & ~n8988;
  assign n8990 = ~n5616 & ~n8989;
  assign n8991 = controllable_hmaster0 & ~n8990;
  assign n8992 = ~controllable_hmaster0 & ~n5624;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = ~controllable_hmaster1 & ~n8993;
  assign n8995 = ~n8985 & ~n8994;
  assign n8996 = i_hbusreq3 & ~n8995;
  assign n8997 = ~n5863 & ~n8969;
  assign n8998 = ~i_hbusreq2 & ~n8997;
  assign n8999 = ~n5636 & ~n8998;
  assign n9000 = ~controllable_hgrant2 & ~n8999;
  assign n9001 = ~n5862 & ~n9000;
  assign n9002 = controllable_hmaster0 & ~n9001;
  assign n9003 = ~n5950 & ~n9000;
  assign n9004 = ~controllable_hmaster0 & ~n9003;
  assign n9005 = ~n9002 & ~n9004;
  assign n9006 = controllable_hmaster1 & ~n9005;
  assign n9007 = i_hbusreq2 & ~n8988;
  assign n9008 = i_hbusreq4 & ~n8986;
  assign n9009 = i_hbusreq0 & ~n8986;
  assign n9010 = ~i_hbusreq1 & n3902;
  assign n9011 = ~n5730 & ~n9010;
  assign n9012 = ~controllable_ndecide & n9011;
  assign n9013 = ~n3494 & ~n9012;
  assign n9014 = i_hready & ~n9013;
  assign n9015 = ~n3511 & ~n9014;
  assign n9016 = i_hlock0 & ~n9015;
  assign n9017 = ~n3495 & ~n5966;
  assign n9018 = ~i_hlock0 & ~n9017;
  assign n9019 = ~n9016 & ~n9018;
  assign n9020 = ~i_hbusreq0 & ~n9019;
  assign n9021 = ~n9009 & ~n9020;
  assign n9022 = ~i_hbusreq4 & ~n9021;
  assign n9023 = ~n9008 & ~n9022;
  assign n9024 = ~controllable_hgrant4 & ~n9023;
  assign n9025 = ~n5863 & ~n9024;
  assign n9026 = ~i_hbusreq2 & ~n9025;
  assign n9027 = ~n9007 & ~n9026;
  assign n9028 = ~controllable_hgrant2 & ~n9027;
  assign n9029 = ~n5862 & ~n9028;
  assign n9030 = controllable_hmaster0 & ~n9029;
  assign n9031 = ~n8862 & ~n8961;
  assign n9032 = i_hlock0 & ~n9031;
  assign n9033 = ~n5891 & ~n9032;
  assign n9034 = ~i_hbusreq0 & ~n9033;
  assign n9035 = ~n5638 & ~n9034;
  assign n9036 = ~i_hbusreq4 & ~n9035;
  assign n9037 = ~n5637 & ~n9036;
  assign n9038 = ~controllable_hgrant4 & ~n9037;
  assign n9039 = ~n5982 & ~n9038;
  assign n9040 = ~i_hbusreq2 & ~n9039;
  assign n9041 = ~n5636 & ~n9040;
  assign n9042 = ~controllable_hgrant2 & ~n9041;
  assign n9043 = ~n5981 & ~n9042;
  assign n9044 = ~controllable_hmaster0 & ~n9043;
  assign n9045 = ~n9030 & ~n9044;
  assign n9046 = ~controllable_hmaster1 & ~n9045;
  assign n9047 = ~n9006 & ~n9046;
  assign n9048 = ~i_hbusreq3 & ~n9047;
  assign n9049 = ~n8996 & ~n9048;
  assign n9050 = ~controllable_hmaster2 & ~n9049;
  assign n9051 = ~n8981 & ~n9050;
  assign n9052 = ~controllable_hgrant3 & ~n9051;
  assign n9053 = ~n8935 & ~n9052;
  assign n9054 = controllable_nhgrant0 & ~n9053;
  assign n9055 = ~n3495 & ~n6007;
  assign n9056 = ~controllable_hgrant4 & ~n9055;
  assign n9057 = ~n3411 & ~n9056;
  assign n9058 = ~controllable_hgrant2 & ~n9057;
  assign n9059 = ~n3410 & ~n9058;
  assign n9060 = controllable_hmaster1 & ~n9059;
  assign n9061 = controllable_hmaster0 & ~n9059;
  assign n9062 = ~controllable_hmaster0 & ~n6012;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = ~controllable_hmaster1 & ~n9063;
  assign n9065 = ~n9060 & ~n9064;
  assign n9066 = i_hbusreq3 & ~n9065;
  assign n9067 = i_hbusreq2 & ~n9057;
  assign n9068 = i_hbusreq4 & ~n9055;
  assign n9069 = i_hbusreq0 & ~n9055;
  assign n9070 = ~n3495 & ~n6018;
  assign n9071 = i_hlock0 & ~n9070;
  assign n9072 = ~i_hlock0 & ~n9055;
  assign n9073 = ~n9071 & ~n9072;
  assign n9074 = ~i_hbusreq0 & ~n9073;
  assign n9075 = ~n9069 & ~n9074;
  assign n9076 = ~i_hbusreq4 & ~n9075;
  assign n9077 = ~n9068 & ~n9076;
  assign n9078 = ~controllable_hgrant4 & ~n9077;
  assign n9079 = ~n3411 & ~n9078;
  assign n9080 = ~i_hbusreq2 & ~n9079;
  assign n9081 = ~n9067 & ~n9080;
  assign n9082 = ~controllable_hgrant2 & ~n9081;
  assign n9083 = ~n3410 & ~n9082;
  assign n9084 = controllable_hmaster1 & ~n9083;
  assign n9085 = controllable_hmaster0 & ~n9083;
  assign n9086 = ~controllable_hmaster0 & ~n6032;
  assign n9087 = ~n9085 & ~n9086;
  assign n9088 = ~controllable_hmaster1 & ~n9087;
  assign n9089 = ~n9084 & ~n9088;
  assign n9090 = ~i_hbusreq3 & ~n9089;
  assign n9091 = ~n9066 & ~n9090;
  assign n9092 = controllable_hmaster2 & ~n9091;
  assign n9093 = ~n6078 & ~n9092;
  assign n9094 = ~controllable_hgrant3 & ~n9093;
  assign n9095 = ~n8888 & ~n9094;
  assign n9096 = ~controllable_nhgrant0 & ~n9095;
  assign n9097 = ~n9054 & ~n9096;
  assign n9098 = ~n3281 & ~n9097;
  assign n9099 = ~n4089 & ~n9098;
  assign n9100 = ~n3378 & ~n9099;
  assign n9101 = ~n8913 & ~n9100;
  assign n9102 = n3492 & ~n9101;
  assign n9103 = ~n8309 & ~n9102;
  assign n9104 = n3485 & ~n9103;
  assign n9105 = ~n8639 & ~n9104;
  assign n9106 = n3476 & ~n9105;
  assign n9107 = ~n8912 & ~n9106;
  assign n9108 = n3374 & ~n9107;
  assign n9109 = ~n8801 & ~n9108;
  assign n9110 = n3655 & ~n9109;
  assign n9111 = n3378 & ~n6195;
  assign n9112 = ~controllable_hgrant4 & n3417;
  assign n9113 = ~n3411 & ~n9112;
  assign n9114 = ~controllable_hgrant2 & ~n9113;
  assign n9115 = ~n3410 & ~n9114;
  assign n9116 = controllable_hmaster1 & ~n9115;
  assign n9117 = controllable_hmaster0 & ~n9115;
  assign n9118 = ~n3729 & ~n9117;
  assign n9119 = ~controllable_hmaster1 & ~n9118;
  assign n9120 = ~n9116 & ~n9119;
  assign n9121 = i_hbusreq3 & ~n9120;
  assign n9122 = ~n3767 & ~n9117;
  assign n9123 = ~controllable_hmaster1 & ~n9122;
  assign n9124 = ~n9116 & ~n9123;
  assign n9125 = ~i_hbusreq3 & ~n9124;
  assign n9126 = ~n9121 & ~n9125;
  assign n9127 = controllable_hmaster2 & ~n9126;
  assign n9128 = ~n6188 & ~n9127;
  assign n9129 = ~controllable_hgrant3 & ~n9128;
  assign n9130 = ~n8750 & ~n9129;
  assign n9131 = controllable_nhgrant0 & ~n9130;
  assign n9132 = ~n8785 & ~n9131;
  assign n9133 = ~n3281 & ~n9132;
  assign n9134 = ~n3783 & ~n9133;
  assign n9135 = ~n3378 & ~n9134;
  assign n9136 = ~n9111 & ~n9135;
  assign n9137 = n3492 & ~n9136;
  assign n9138 = ~n3631 & ~n9137;
  assign n9139 = n3485 & ~n9138;
  assign n9140 = ~n3630 & ~n9139;
  assign n9141 = ~n3476 & ~n9140;
  assign n9142 = ~n8367 & ~n9137;
  assign n9143 = n3485 & ~n9142;
  assign n9144 = ~n8650 & ~n9143;
  assign n9145 = n3476 & ~n9144;
  assign n9146 = ~n9141 & ~n9145;
  assign n9147 = ~n3374 & ~n9146;
  assign n9148 = n3378 & ~n6350;
  assign n9149 = ~n4186 & ~n9117;
  assign n9150 = ~controllable_hmaster1 & ~n9149;
  assign n9151 = ~n9116 & ~n9150;
  assign n9152 = i_hbusreq3 & ~n9151;
  assign n9153 = ~n4210 & ~n9117;
  assign n9154 = ~controllable_hmaster1 & ~n9153;
  assign n9155 = ~n9116 & ~n9154;
  assign n9156 = ~i_hbusreq3 & ~n9155;
  assign n9157 = ~n9152 & ~n9156;
  assign n9158 = controllable_hmaster2 & ~n9157;
  assign n9159 = ~n3411 & ~n4182;
  assign n9160 = ~controllable_hgrant2 & ~n9159;
  assign n9161 = ~n3410 & ~n9160;
  assign n9162 = controllable_hmaster0 & ~n9161;
  assign n9163 = ~n5288 & ~n9160;
  assign n9164 = ~controllable_hmaster0 & ~n9163;
  assign n9165 = ~n9162 & ~n9164;
  assign n9166 = controllable_hmaster1 & ~n9165;
  assign n9167 = controllable_ndecide & ~n6512;
  assign n9168 = ~i_hready & ~n9167;
  assign n9169 = ~n6259 & ~n9168;
  assign n9170 = ~controllable_hgrant4 & n9169;
  assign n9171 = ~n3411 & ~n9170;
  assign n9172 = ~controllable_hgrant2 & ~n9171;
  assign n9173 = ~n3410 & ~n9172;
  assign n9174 = controllable_hmaster0 & ~n9173;
  assign n9175 = ~controllable_hmaster0 & ~n9161;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = ~controllable_hmaster1 & ~n9176;
  assign n9178 = ~n9166 & ~n9177;
  assign n9179 = i_hbusreq3 & ~n9178;
  assign n9180 = i_hbusreq2 & ~n9159;
  assign n9181 = ~n3916 & ~n4204;
  assign n9182 = ~i_hbusreq2 & ~n9181;
  assign n9183 = ~n9180 & ~n9182;
  assign n9184 = ~controllable_hgrant2 & ~n9183;
  assign n9185 = ~n3859 & ~n9184;
  assign n9186 = controllable_hmaster0 & ~n9185;
  assign n9187 = ~n5438 & ~n9184;
  assign n9188 = ~controllable_hmaster0 & ~n9187;
  assign n9189 = ~n9186 & ~n9188;
  assign n9190 = controllable_hmaster1 & ~n9189;
  assign n9191 = i_hbusreq2 & ~n9171;
  assign n9192 = i_hbusreq4 & ~n9169;
  assign n9193 = i_hbusreq0 & ~n9169;
  assign n9194 = ~n6304 & ~n6512;
  assign n9195 = ~i_hready & ~n9194;
  assign n9196 = ~n6303 & ~n9195;
  assign n9197 = i_hlock0 & ~n9196;
  assign n9198 = ~i_hlock0 & ~n9169;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = ~i_hbusreq0 & ~n9199;
  assign n9201 = ~n9193 & ~n9200;
  assign n9202 = ~i_hbusreq4 & ~n9201;
  assign n9203 = ~n9192 & ~n9202;
  assign n9204 = ~controllable_hgrant4 & n9203;
  assign n9205 = ~n3916 & ~n9204;
  assign n9206 = ~i_hbusreq2 & ~n9205;
  assign n9207 = ~n9191 & ~n9206;
  assign n9208 = ~controllable_hgrant2 & ~n9207;
  assign n9209 = ~n3859 & ~n9208;
  assign n9210 = controllable_hmaster0 & ~n9209;
  assign n9211 = ~n4179 & ~n5382;
  assign n9212 = ~i_hready & ~n9211;
  assign n9213 = ~i_hready & ~n9212;
  assign n9214 = i_hlock0 & ~n9213;
  assign n9215 = ~n4198 & ~n9214;
  assign n9216 = ~i_hbusreq0 & ~n9215;
  assign n9217 = ~n4193 & ~n9216;
  assign n9218 = ~i_hbusreq4 & ~n9217;
  assign n9219 = ~n4192 & ~n9218;
  assign n9220 = ~controllable_hgrant4 & ~n9219;
  assign n9221 = ~n5462 & ~n9220;
  assign n9222 = ~i_hbusreq2 & ~n9221;
  assign n9223 = ~n9180 & ~n9222;
  assign n9224 = ~controllable_hgrant2 & ~n9223;
  assign n9225 = ~n5461 & ~n9224;
  assign n9226 = ~controllable_hmaster0 & ~n9225;
  assign n9227 = ~n9210 & ~n9226;
  assign n9228 = ~controllable_hmaster1 & ~n9227;
  assign n9229 = ~n9190 & ~n9228;
  assign n9230 = ~i_hbusreq3 & ~n9229;
  assign n9231 = ~n9179 & ~n9230;
  assign n9232 = ~controllable_hmaster2 & ~n9231;
  assign n9233 = ~n9158 & ~n9232;
  assign n9234 = ~controllable_hgrant3 & ~n9233;
  assign n9235 = ~n8810 & ~n9234;
  assign n9236 = controllable_nhgrant0 & ~n9235;
  assign n9237 = ~n8902 & ~n9236;
  assign n9238 = ~n3281 & ~n9237;
  assign n9239 = ~n3950 & ~n9238;
  assign n9240 = ~n3378 & ~n9239;
  assign n9241 = ~n9148 & ~n9240;
  assign n9242 = n3492 & ~n9241;
  assign n9243 = ~n3631 & ~n9242;
  assign n9244 = n3485 & ~n9243;
  assign n9245 = ~n3630 & ~n9244;
  assign n9246 = ~n3476 & ~n9245;
  assign n9247 = n3378 & ~n6561;
  assign n9248 = ~controllable_hgrant4 & n6401;
  assign n9249 = ~n4091 & ~n9248;
  assign n9250 = ~controllable_hgrant2 & ~n9249;
  assign n9251 = ~n5616 & ~n9250;
  assign n9252 = controllable_hmaster1 & ~n9251;
  assign n9253 = controllable_hmaster0 & ~n9251;
  assign n9254 = ~n6412 & ~n9253;
  assign n9255 = ~controllable_hmaster1 & ~n9254;
  assign n9256 = ~n9252 & ~n9255;
  assign n9257 = i_hbusreq3 & ~n9256;
  assign n9258 = i_hbusreq2 & ~n9249;
  assign n9259 = i_hbusreq4 & n6401;
  assign n9260 = i_hbusreq0 & n6401;
  assign n9261 = ~n4179 & ~n8940;
  assign n9262 = i_hready & ~n9261;
  assign n9263 = i_hlock0 & n9262;
  assign n9264 = ~i_hlock0 & n6425;
  assign n9265 = ~n9263 & ~n9264;
  assign n9266 = ~i_hbusreq0 & ~n9265;
  assign n9267 = ~n9260 & ~n9266;
  assign n9268 = ~i_hbusreq4 & ~n9267;
  assign n9269 = ~n9259 & ~n9268;
  assign n9270 = ~controllable_hgrant4 & ~n9269;
  assign n9271 = ~n8937 & ~n9270;
  assign n9272 = ~i_hbusreq2 & ~n9271;
  assign n9273 = ~n9258 & ~n9272;
  assign n9274 = ~controllable_hgrant2 & ~n9273;
  assign n9275 = ~n8936 & ~n9274;
  assign n9276 = controllable_hmaster1 & ~n9275;
  assign n9277 = controllable_hmaster0 & ~n9275;
  assign n9278 = ~n4179 & ~n8959;
  assign n9279 = i_hready & ~n9278;
  assign n9280 = ~n4195 & ~n9279;
  assign n9281 = i_hlock0 & ~n9280;
  assign n9282 = ~n6445 & ~n9281;
  assign n9283 = ~i_hbusreq0 & ~n9282;
  assign n9284 = ~n6419 & ~n9283;
  assign n9285 = ~i_hbusreq4 & ~n9284;
  assign n9286 = ~n6418 & ~n9285;
  assign n9287 = ~controllable_hgrant4 & ~n9286;
  assign n9288 = ~n4064 & ~n9287;
  assign n9289 = ~i_hbusreq2 & ~n9288;
  assign n9290 = ~n6441 & ~n9289;
  assign n9291 = ~controllable_hgrant2 & ~n9290;
  assign n9292 = ~n5862 & ~n9291;
  assign n9293 = ~controllable_hmaster0 & ~n9292;
  assign n9294 = ~n9277 & ~n9293;
  assign n9295 = ~controllable_hmaster1 & ~n9294;
  assign n9296 = ~n9276 & ~n9295;
  assign n9297 = ~i_hbusreq3 & ~n9296;
  assign n9298 = ~n9257 & ~n9297;
  assign n9299 = controllable_hmaster2 & ~n9298;
  assign n9300 = ~n5686 & ~n6405;
  assign n9301 = ~controllable_hmaster0 & ~n9300;
  assign n9302 = ~n6408 & ~n9301;
  assign n9303 = controllable_hmaster1 & ~n9302;
  assign n9304 = ~n6474 & ~n9168;
  assign n9305 = ~controllable_hgrant4 & n9304;
  assign n9306 = ~n4091 & ~n9305;
  assign n9307 = ~controllable_hgrant2 & ~n9306;
  assign n9308 = ~n5616 & ~n9307;
  assign n9309 = controllable_hmaster0 & ~n9308;
  assign n9310 = ~controllable_hmaster0 & ~n6406;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = ~controllable_hmaster1 & ~n9311;
  assign n9313 = ~n9303 & ~n9312;
  assign n9314 = i_hbusreq3 & ~n9313;
  assign n9315 = ~n5863 & ~n9287;
  assign n9316 = ~i_hbusreq2 & ~n9315;
  assign n9317 = ~n6417 & ~n9316;
  assign n9318 = ~controllable_hgrant2 & ~n9317;
  assign n9319 = ~n5862 & ~n9318;
  assign n9320 = controllable_hmaster0 & ~n9319;
  assign n9321 = ~n5950 & ~n9318;
  assign n9322 = ~controllable_hmaster0 & ~n9321;
  assign n9323 = ~n9320 & ~n9322;
  assign n9324 = controllable_hmaster1 & ~n9323;
  assign n9325 = i_hbusreq2 & ~n9306;
  assign n9326 = i_hbusreq4 & ~n9304;
  assign n9327 = i_hbusreq0 & ~n9304;
  assign n9328 = ~controllable_ndecide & ~n9011;
  assign n9329 = ~n6512 & ~n9328;
  assign n9330 = i_hready & ~n9329;
  assign n9331 = ~n9195 & ~n9330;
  assign n9332 = i_hlock0 & ~n9331;
  assign n9333 = ~n6520 & ~n9168;
  assign n9334 = ~i_hlock0 & ~n9333;
  assign n9335 = ~n9332 & ~n9334;
  assign n9336 = ~i_hbusreq0 & ~n9335;
  assign n9337 = ~n9327 & ~n9336;
  assign n9338 = ~i_hbusreq4 & ~n9337;
  assign n9339 = ~n9326 & ~n9338;
  assign n9340 = ~controllable_hgrant4 & n9339;
  assign n9341 = ~n5863 & ~n9340;
  assign n9342 = ~i_hbusreq2 & ~n9341;
  assign n9343 = ~n9325 & ~n9342;
  assign n9344 = ~controllable_hgrant2 & ~n9343;
  assign n9345 = ~n5862 & ~n9344;
  assign n9346 = controllable_hmaster0 & ~n9345;
  assign n9347 = ~n9212 & ~n9279;
  assign n9348 = i_hlock0 & ~n9347;
  assign n9349 = ~n6445 & ~n9348;
  assign n9350 = ~i_hbusreq0 & ~n9349;
  assign n9351 = ~n6419 & ~n9350;
  assign n9352 = ~i_hbusreq4 & ~n9351;
  assign n9353 = ~n6418 & ~n9352;
  assign n9354 = ~controllable_hgrant4 & ~n9353;
  assign n9355 = ~n5982 & ~n9354;
  assign n9356 = ~i_hbusreq2 & ~n9355;
  assign n9357 = ~n6417 & ~n9356;
  assign n9358 = ~controllable_hgrant2 & ~n9357;
  assign n9359 = ~n5981 & ~n9358;
  assign n9360 = ~controllable_hmaster0 & ~n9359;
  assign n9361 = ~n9346 & ~n9360;
  assign n9362 = ~controllable_hmaster1 & ~n9361;
  assign n9363 = ~n9324 & ~n9362;
  assign n9364 = ~i_hbusreq3 & ~n9363;
  assign n9365 = ~n9314 & ~n9364;
  assign n9366 = ~controllable_hmaster2 & ~n9365;
  assign n9367 = ~n9299 & ~n9366;
  assign n9368 = ~controllable_hgrant3 & ~n9367;
  assign n9369 = ~n8935 & ~n9368;
  assign n9370 = controllable_nhgrant0 & ~n9369;
  assign n9371 = ~n9096 & ~n9370;
  assign n9372 = ~n3281 & ~n9371;
  assign n9373 = ~n4089 & ~n9372;
  assign n9374 = ~n3378 & ~n9373;
  assign n9375 = ~n9247 & ~n9374;
  assign n9376 = n3492 & ~n9375;
  assign n9377 = ~n8367 & ~n9376;
  assign n9378 = n3485 & ~n9377;
  assign n9379 = ~n8650 & ~n9378;
  assign n9380 = n3476 & ~n9379;
  assign n9381 = ~n9246 & ~n9380;
  assign n9382 = n3374 & ~n9381;
  assign n9383 = ~n9147 & ~n9382;
  assign n9384 = ~n3655 & ~n9383;
  assign n9385 = ~n9110 & ~n9384;
  assign n9386 = n3652 & ~n9385;
  assign n9387 = n3378 & ~n6664;
  assign n9388 = controllable_hgrant2 & ~n8767;
  assign n9389 = ~n3499 & ~n9388;
  assign n9390 = controllable_hmaster1 & ~n9389;
  assign n9391 = controllable_hmaster0 & ~n9389;
  assign n9392 = ~n3729 & ~n9391;
  assign n9393 = ~controllable_hmaster1 & ~n9392;
  assign n9394 = ~n9390 & ~n9393;
  assign n9395 = i_hbusreq3 & ~n9394;
  assign n9396 = ~n3767 & ~n9391;
  assign n9397 = ~controllable_hmaster1 & ~n9396;
  assign n9398 = ~n9390 & ~n9397;
  assign n9399 = ~i_hbusreq3 & ~n9398;
  assign n9400 = ~n9395 & ~n9399;
  assign n9401 = controllable_hmaster2 & ~n9400;
  assign n9402 = ~n6657 & ~n9401;
  assign n9403 = ~controllable_hgrant3 & ~n9402;
  assign n9404 = ~n8750 & ~n9403;
  assign n9405 = controllable_nhgrant0 & ~n9404;
  assign n9406 = ~n8785 & ~n9405;
  assign n9407 = ~n3281 & ~n9406;
  assign n9408 = ~n3783 & ~n9407;
  assign n9409 = ~n3378 & ~n9408;
  assign n9410 = ~n9387 & ~n9409;
  assign n9411 = n3492 & ~n9410;
  assign n9412 = ~n3631 & ~n9411;
  assign n9413 = n3485 & ~n9412;
  assign n9414 = ~n3630 & ~n9413;
  assign n9415 = ~n3476 & ~n9414;
  assign n9416 = ~n8434 & ~n9411;
  assign n9417 = n3485 & ~n9416;
  assign n9418 = ~n8663 & ~n9417;
  assign n9419 = n3476 & ~n9418;
  assign n9420 = ~n9415 & ~n9419;
  assign n9421 = ~n3374 & ~n9420;
  assign n9422 = n3378 & ~n6730;
  assign n9423 = ~n4335 & ~n9391;
  assign n9424 = ~controllable_hmaster1 & ~n9423;
  assign n9425 = ~n9390 & ~n9424;
  assign n9426 = i_hbusreq3 & ~n9425;
  assign n9427 = ~n4342 & ~n9391;
  assign n9428 = ~controllable_hmaster1 & ~n9427;
  assign n9429 = ~n9390 & ~n9428;
  assign n9430 = ~i_hbusreq3 & ~n9429;
  assign n9431 = ~n9426 & ~n9430;
  assign n9432 = controllable_hmaster2 & ~n9431;
  assign n9433 = ~n4333 & ~n8768;
  assign n9434 = controllable_hmaster0 & ~n9433;
  assign n9435 = ~n6697 & ~n8768;
  assign n9436 = ~controllable_hmaster0 & ~n9435;
  assign n9437 = ~n9434 & ~n9436;
  assign n9438 = controllable_hmaster1 & ~n9437;
  assign n9439 = ~n4333 & ~n8824;
  assign n9440 = controllable_hmaster0 & ~n9439;
  assign n9441 = ~controllable_hmaster0 & ~n9433;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = ~controllable_hmaster1 & ~n9442;
  assign n9444 = ~n9438 & ~n9443;
  assign n9445 = i_hbusreq3 & ~n9444;
  assign n9446 = ~n4340 & ~n8836;
  assign n9447 = controllable_hmaster0 & ~n9446;
  assign n9448 = ~n6710 & ~n8836;
  assign n9449 = ~controllable_hmaster0 & ~n9448;
  assign n9450 = ~n9447 & ~n9449;
  assign n9451 = controllable_hmaster1 & ~n9450;
  assign n9452 = ~n4340 & ~n8858;
  assign n9453 = controllable_hmaster0 & ~n9452;
  assign n9454 = ~n6947 & ~n8874;
  assign n9455 = ~controllable_hmaster0 & ~n9454;
  assign n9456 = ~n9453 & ~n9455;
  assign n9457 = ~controllable_hmaster1 & ~n9456;
  assign n9458 = ~n9451 & ~n9457;
  assign n9459 = ~i_hbusreq3 & ~n9458;
  assign n9460 = ~n9445 & ~n9459;
  assign n9461 = ~controllable_hmaster2 & ~n9460;
  assign n9462 = ~n9432 & ~n9461;
  assign n9463 = ~controllable_hgrant3 & ~n9462;
  assign n9464 = ~n8810 & ~n9463;
  assign n9465 = controllable_nhgrant0 & ~n9464;
  assign n9466 = ~n8902 & ~n9465;
  assign n9467 = ~n3281 & ~n9466;
  assign n9468 = ~n3950 & ~n9467;
  assign n9469 = ~n3378 & ~n9468;
  assign n9470 = ~n9422 & ~n9469;
  assign n9471 = n3492 & ~n9470;
  assign n9472 = ~n3631 & ~n9471;
  assign n9473 = n3485 & ~n9472;
  assign n9474 = ~n3630 & ~n9473;
  assign n9475 = ~n3476 & ~n9474;
  assign n9476 = n3378 & ~n6846;
  assign n9477 = controllable_hgrant2 & ~n9057;
  assign n9478 = ~n5623 & ~n9477;
  assign n9479 = controllable_hmaster1 & ~n9478;
  assign n9480 = controllable_hmaster0 & ~n9478;
  assign n9481 = ~n6767 & ~n9480;
  assign n9482 = ~controllable_hmaster1 & ~n9481;
  assign n9483 = ~n9479 & ~n9482;
  assign n9484 = i_hbusreq3 & ~n9483;
  assign n9485 = controllable_hgrant2 & ~n9081;
  assign n9486 = ~n8954 & ~n9485;
  assign n9487 = controllable_hmaster1 & ~n9486;
  assign n9488 = controllable_hmaster0 & ~n9486;
  assign n9489 = ~n6772 & ~n8973;
  assign n9490 = ~controllable_hmaster0 & ~n9489;
  assign n9491 = ~n9488 & ~n9490;
  assign n9492 = ~controllable_hmaster1 & ~n9491;
  assign n9493 = ~n9487 & ~n9492;
  assign n9494 = ~i_hbusreq3 & ~n9493;
  assign n9495 = ~n9484 & ~n9494;
  assign n9496 = controllable_hmaster2 & ~n9495;
  assign n9497 = ~n5623 & ~n6786;
  assign n9498 = ~controllable_hmaster0 & ~n9497;
  assign n9499 = ~n6765 & ~n9498;
  assign n9500 = controllable_hmaster1 & ~n9499;
  assign n9501 = ~n6762 & ~n8989;
  assign n9502 = controllable_hmaster0 & ~n9501;
  assign n9503 = ~controllable_hmaster0 & ~n6763;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = ~controllable_hmaster1 & ~n9504;
  assign n9506 = ~n9500 & ~n9505;
  assign n9507 = i_hbusreq3 & ~n9506;
  assign n9508 = ~n6772 & ~n9000;
  assign n9509 = controllable_hmaster0 & ~n9508;
  assign n9510 = ~n6813 & ~n9000;
  assign n9511 = ~controllable_hmaster0 & ~n9510;
  assign n9512 = ~n9509 & ~n9511;
  assign n9513 = controllable_hmaster1 & ~n9512;
  assign n9514 = ~n6772 & ~n9028;
  assign n9515 = controllable_hmaster0 & ~n9514;
  assign n9516 = ~n6831 & ~n9042;
  assign n9517 = ~controllable_hmaster0 & ~n9516;
  assign n9518 = ~n9515 & ~n9517;
  assign n9519 = ~controllable_hmaster1 & ~n9518;
  assign n9520 = ~n9513 & ~n9519;
  assign n9521 = ~i_hbusreq3 & ~n9520;
  assign n9522 = ~n9507 & ~n9521;
  assign n9523 = ~controllable_hmaster2 & ~n9522;
  assign n9524 = ~n9496 & ~n9523;
  assign n9525 = ~controllable_hgrant3 & ~n9524;
  assign n9526 = ~n8935 & ~n9525;
  assign n9527 = controllable_nhgrant0 & ~n9526;
  assign n9528 = ~n9096 & ~n9527;
  assign n9529 = ~n3281 & ~n9528;
  assign n9530 = ~n4089 & ~n9529;
  assign n9531 = ~n3378 & ~n9530;
  assign n9532 = ~n9476 & ~n9531;
  assign n9533 = n3492 & ~n9532;
  assign n9534 = ~n8434 & ~n9533;
  assign n9535 = n3485 & ~n9534;
  assign n9536 = ~n8663 & ~n9535;
  assign n9537 = n3476 & ~n9536;
  assign n9538 = ~n9475 & ~n9537;
  assign n9539 = n3374 & ~n9538;
  assign n9540 = ~n9421 & ~n9539;
  assign n9541 = n3655 & ~n9540;
  assign n9542 = n3378 & ~n6894;
  assign n9543 = ~n9114 & ~n9388;
  assign n9544 = controllable_hmaster1 & ~n9543;
  assign n9545 = controllable_hmaster0 & ~n9543;
  assign n9546 = ~n3729 & ~n9545;
  assign n9547 = ~controllable_hmaster1 & ~n9546;
  assign n9548 = ~n9544 & ~n9547;
  assign n9549 = i_hbusreq3 & ~n9548;
  assign n9550 = ~n3767 & ~n9545;
  assign n9551 = ~controllable_hmaster1 & ~n9550;
  assign n9552 = ~n9544 & ~n9551;
  assign n9553 = ~i_hbusreq3 & ~n9552;
  assign n9554 = ~n9549 & ~n9553;
  assign n9555 = controllable_hmaster2 & ~n9554;
  assign n9556 = ~n6887 & ~n9555;
  assign n9557 = ~controllable_hgrant3 & ~n9556;
  assign n9558 = ~n8750 & ~n9557;
  assign n9559 = controllable_nhgrant0 & ~n9558;
  assign n9560 = ~n8785 & ~n9559;
  assign n9561 = ~n3281 & ~n9560;
  assign n9562 = ~n3783 & ~n9561;
  assign n9563 = ~n3378 & ~n9562;
  assign n9564 = ~n9542 & ~n9563;
  assign n9565 = n3492 & ~n9564;
  assign n9566 = ~n3631 & ~n9565;
  assign n9567 = n3485 & ~n9566;
  assign n9568 = ~n3630 & ~n9567;
  assign n9569 = ~n3476 & ~n9568;
  assign n9570 = ~n8491 & ~n9565;
  assign n9571 = n3485 & ~n9570;
  assign n9572 = ~n8674 & ~n9571;
  assign n9573 = n3476 & ~n9572;
  assign n9574 = ~n9569 & ~n9573;
  assign n9575 = ~n3374 & ~n9574;
  assign n9576 = n3378 & ~n6962;
  assign n9577 = ~n4436 & ~n9545;
  assign n9578 = ~controllable_hmaster1 & ~n9577;
  assign n9579 = ~n9544 & ~n9578;
  assign n9580 = i_hbusreq3 & ~n9579;
  assign n9581 = ~n4442 & ~n9545;
  assign n9582 = ~controllable_hmaster1 & ~n9581;
  assign n9583 = ~n9544 & ~n9582;
  assign n9584 = ~i_hbusreq3 & ~n9583;
  assign n9585 = ~n9580 & ~n9584;
  assign n9586 = controllable_hmaster2 & ~n9585;
  assign n9587 = ~n4333 & ~n9160;
  assign n9588 = controllable_hmaster0 & ~n9587;
  assign n9589 = ~n6697 & ~n9160;
  assign n9590 = ~controllable_hmaster0 & ~n9589;
  assign n9591 = ~n9588 & ~n9590;
  assign n9592 = controllable_hmaster1 & ~n9591;
  assign n9593 = ~n4333 & ~n9172;
  assign n9594 = controllable_hmaster0 & ~n9593;
  assign n9595 = ~controllable_hmaster0 & ~n9587;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = ~controllable_hmaster1 & ~n9596;
  assign n9598 = ~n9592 & ~n9597;
  assign n9599 = i_hbusreq3 & ~n9598;
  assign n9600 = ~n4340 & ~n9184;
  assign n9601 = controllable_hmaster0 & ~n9600;
  assign n9602 = ~n6710 & ~n9184;
  assign n9603 = ~controllable_hmaster0 & ~n9602;
  assign n9604 = ~n9601 & ~n9603;
  assign n9605 = controllable_hmaster1 & ~n9604;
  assign n9606 = ~n4340 & ~n9208;
  assign n9607 = controllable_hmaster0 & ~n9606;
  assign n9608 = ~n6947 & ~n9224;
  assign n9609 = ~controllable_hmaster0 & ~n9608;
  assign n9610 = ~n9607 & ~n9609;
  assign n9611 = ~controllable_hmaster1 & ~n9610;
  assign n9612 = ~n9605 & ~n9611;
  assign n9613 = ~i_hbusreq3 & ~n9612;
  assign n9614 = ~n9599 & ~n9613;
  assign n9615 = ~controllable_hmaster2 & ~n9614;
  assign n9616 = ~n9586 & ~n9615;
  assign n9617 = ~controllable_hgrant3 & ~n9616;
  assign n9618 = ~n8810 & ~n9617;
  assign n9619 = controllable_nhgrant0 & ~n9618;
  assign n9620 = ~n8902 & ~n9619;
  assign n9621 = ~n3281 & ~n9620;
  assign n9622 = ~n3950 & ~n9621;
  assign n9623 = ~n3378 & ~n9622;
  assign n9624 = ~n9576 & ~n9623;
  assign n9625 = n3492 & ~n9624;
  assign n9626 = ~n3631 & ~n9625;
  assign n9627 = n3485 & ~n9626;
  assign n9628 = ~n3630 & ~n9627;
  assign n9629 = ~n3476 & ~n9628;
  assign n9630 = n3378 & ~n7047;
  assign n9631 = ~n9250 & ~n9477;
  assign n9632 = controllable_hmaster1 & ~n9631;
  assign n9633 = controllable_hmaster0 & ~n9631;
  assign n9634 = ~n6996 & ~n9633;
  assign n9635 = ~controllable_hmaster1 & ~n9634;
  assign n9636 = ~n9632 & ~n9635;
  assign n9637 = i_hbusreq3 & ~n9636;
  assign n9638 = ~n9274 & ~n9485;
  assign n9639 = controllable_hmaster1 & ~n9638;
  assign n9640 = controllable_hmaster0 & ~n9638;
  assign n9641 = ~n6772 & ~n9291;
  assign n9642 = ~controllable_hmaster0 & ~n9641;
  assign n9643 = ~n9640 & ~n9642;
  assign n9644 = ~controllable_hmaster1 & ~n9643;
  assign n9645 = ~n9639 & ~n9644;
  assign n9646 = ~i_hbusreq3 & ~n9645;
  assign n9647 = ~n9637 & ~n9646;
  assign n9648 = controllable_hmaster2 & ~n9647;
  assign n9649 = ~n6405 & ~n6786;
  assign n9650 = ~controllable_hmaster0 & ~n9649;
  assign n9651 = ~n6994 & ~n9650;
  assign n9652 = controllable_hmaster1 & ~n9651;
  assign n9653 = ~n6762 & ~n9307;
  assign n9654 = controllable_hmaster0 & ~n9653;
  assign n9655 = ~controllable_hmaster0 & ~n6992;
  assign n9656 = ~n9654 & ~n9655;
  assign n9657 = ~controllable_hmaster1 & ~n9656;
  assign n9658 = ~n9652 & ~n9657;
  assign n9659 = i_hbusreq3 & ~n9658;
  assign n9660 = ~n6772 & ~n9318;
  assign n9661 = controllable_hmaster0 & ~n9660;
  assign n9662 = ~n6813 & ~n9318;
  assign n9663 = ~controllable_hmaster0 & ~n9662;
  assign n9664 = ~n9661 & ~n9663;
  assign n9665 = controllable_hmaster1 & ~n9664;
  assign n9666 = ~n6772 & ~n9344;
  assign n9667 = controllable_hmaster0 & ~n9666;
  assign n9668 = ~n6831 & ~n9358;
  assign n9669 = ~controllable_hmaster0 & ~n9668;
  assign n9670 = ~n9667 & ~n9669;
  assign n9671 = ~controllable_hmaster1 & ~n9670;
  assign n9672 = ~n9665 & ~n9671;
  assign n9673 = ~i_hbusreq3 & ~n9672;
  assign n9674 = ~n9659 & ~n9673;
  assign n9675 = ~controllable_hmaster2 & ~n9674;
  assign n9676 = ~n9648 & ~n9675;
  assign n9677 = ~controllable_hgrant3 & ~n9676;
  assign n9678 = ~n8935 & ~n9677;
  assign n9679 = controllable_nhgrant0 & ~n9678;
  assign n9680 = ~n9096 & ~n9679;
  assign n9681 = ~n3281 & ~n9680;
  assign n9682 = ~n4089 & ~n9681;
  assign n9683 = ~n3378 & ~n9682;
  assign n9684 = ~n9630 & ~n9683;
  assign n9685 = n3492 & ~n9684;
  assign n9686 = ~n8491 & ~n9685;
  assign n9687 = n3485 & ~n9686;
  assign n9688 = ~n8674 & ~n9687;
  assign n9689 = n3476 & ~n9688;
  assign n9690 = ~n9629 & ~n9689;
  assign n9691 = n3374 & ~n9690;
  assign n9692 = ~n9575 & ~n9691;
  assign n9693 = ~n3655 & ~n9692;
  assign n9694 = ~n9541 & ~n9693;
  assign n9695 = ~n3652 & ~n9694;
  assign n9696 = ~n9386 & ~n9695;
  assign n9697 = ~n3368 & ~n9696;
  assign n9698 = n3378 & ~n7121;
  assign n9699 = controllable_hmaster1 & ~n4552;
  assign n9700 = controllable_hmaster0 & ~n4552;
  assign n9701 = controllable_hmaster0 & ~n9700;
  assign n9702 = ~controllable_hmaster1 & ~n9701;
  assign n9703 = ~n9699 & ~n9702;
  assign n9704 = ~i_hbusreq3 & ~n9703;
  assign n9705 = ~n3386 & ~n9704;
  assign n9706 = controllable_hmaster2 & ~n9705;
  assign n9707 = controllable_hmaster2 & ~n9706;
  assign n9708 = controllable_hgrant3 & ~n9707;
  assign n9709 = ~n3418 & ~n4565;
  assign n9710 = i_hready & ~n9709;
  assign n9711 = ~n4577 & ~n9710;
  assign n9712 = i_hlock0 & ~n9711;
  assign n9713 = ~n5404 & ~n9712;
  assign n9714 = ~i_hbusreq0 & ~n9713;
  assign n9715 = ~n3509 & ~n9714;
  assign n9716 = ~i_hbusreq4 & ~n9715;
  assign n9717 = ~n3508 & ~n9716;
  assign n9718 = ~controllable_hgrant4 & ~n9717;
  assign n9719 = ~n4617 & ~n9718;
  assign n9720 = ~i_hbusreq2 & ~n9719;
  assign n9721 = ~n3507 & ~n9720;
  assign n9722 = ~controllable_hgrant2 & ~n9721;
  assign n9723 = ~n4562 & ~n9722;
  assign n9724 = controllable_hmaster1 & ~n9723;
  assign n9725 = controllable_hmaster0 & ~n9723;
  assign n9726 = controllable_hmaster0 & ~n9725;
  assign n9727 = ~controllable_hmaster1 & ~n9726;
  assign n9728 = ~n9724 & ~n9727;
  assign n9729 = ~i_hbusreq3 & ~n9728;
  assign n9730 = ~n3506 & ~n9729;
  assign n9731 = controllable_hmaster2 & ~n9730;
  assign n9732 = controllable_hmaster2 & ~n9731;
  assign n9733 = ~controllable_hgrant3 & ~n9732;
  assign n9734 = ~n9708 & ~n9733;
  assign n9735 = controllable_nhgrant0 & ~n9734;
  assign n9736 = controllable_hmaster1 & ~n4610;
  assign n9737 = controllable_hmaster0 & ~n4610;
  assign n9738 = controllable_hmaster0 & ~n9737;
  assign n9739 = ~controllable_hmaster1 & ~n9738;
  assign n9740 = ~n9736 & ~n9739;
  assign n9741 = i_hbusreq3 & ~n9740;
  assign n9742 = controllable_hmaster1 & ~n4635;
  assign n9743 = controllable_hmaster0 & ~n4635;
  assign n9744 = controllable_hmaster0 & ~n9743;
  assign n9745 = ~controllable_hmaster1 & ~n9744;
  assign n9746 = ~n9742 & ~n9745;
  assign n9747 = ~i_hbusreq3 & ~n9746;
  assign n9748 = ~n9741 & ~n9747;
  assign n9749 = controllable_hmaster2 & ~n9748;
  assign n9750 = controllable_hmaster2 & ~n9749;
  assign n9751 = ~controllable_hgrant3 & ~n9750;
  assign n9752 = ~n9708 & ~n9751;
  assign n9753 = ~controllable_nhgrant0 & ~n9752;
  assign n9754 = ~n9735 & ~n9753;
  assign n9755 = ~n3281 & ~n9754;
  assign n9756 = ~n3281 & ~n9755;
  assign n9757 = ~n3378 & ~n9756;
  assign n9758 = ~n9698 & ~n9757;
  assign n9759 = n3492 & ~n9758;
  assign n9760 = n3492 & ~n9759;
  assign n9761 = n3485 & ~n9760;
  assign n9762 = n3485 & ~n9761;
  assign n9763 = ~n3476 & ~n9762;
  assign n9764 = ~n8523 & ~n9759;
  assign n9765 = n3485 & ~n9764;
  assign n9766 = ~n8689 & ~n9765;
  assign n9767 = n3476 & ~n9766;
  assign n9768 = ~n9763 & ~n9767;
  assign n9769 = ~n3374 & ~n9768;
  assign n9770 = n3378 & ~n7211;
  assign n9771 = ~i_hbusreq3 & ~n4552;
  assign n9772 = ~n3951 & ~n9771;
  assign n9773 = controllable_hmaster2 & ~n9772;
  assign n9774 = ~controllable_hgrant4 & ~n4574;
  assign n9775 = ~n4617 & ~n9774;
  assign n9776 = ~i_hbusreq2 & ~n9775;
  assign n9777 = ~n5266 & ~n9776;
  assign n9778 = ~controllable_hgrant2 & ~n9777;
  assign n9779 = ~n4562 & ~n9778;
  assign n9780 = controllable_hmaster0 & ~n9779;
  assign n9781 = ~n4553 & ~n9780;
  assign n9782 = controllable_hmaster1 & ~n9781;
  assign n9783 = ~n3821 & ~n9700;
  assign n9784 = ~controllable_hmaster1 & ~n9783;
  assign n9785 = ~n9782 & ~n9784;
  assign n9786 = ~i_hbusreq3 & ~n9785;
  assign n9787 = ~n5265 & ~n9786;
  assign n9788 = ~controllable_hmaster2 & ~n9787;
  assign n9789 = ~n9773 & ~n9788;
  assign n9790 = controllable_hgrant3 & ~n9789;
  assign n9791 = ~n4591 & ~n9725;
  assign n9792 = ~controllable_hmaster1 & ~n9791;
  assign n9793 = ~n9724 & ~n9792;
  assign n9794 = ~i_hbusreq3 & ~n9793;
  assign n9795 = ~n3963 & ~n9794;
  assign n9796 = controllable_hmaster2 & ~n9795;
  assign n9797 = ~n4585 & ~n4617;
  assign n9798 = ~i_hbusreq2 & ~n9797;
  assign n9799 = ~n8832 & ~n9798;
  assign n9800 = ~controllable_hgrant2 & ~n9799;
  assign n9801 = ~n4562 & ~n9800;
  assign n9802 = controllable_hmaster0 & ~n9801;
  assign n9803 = controllable_hgrant2 & ~n9777;
  assign n9804 = ~n9800 & ~n9803;
  assign n9805 = ~controllable_hmaster0 & ~n9804;
  assign n9806 = ~n9802 & ~n9805;
  assign n9807 = controllable_hmaster1 & ~n9806;
  assign n9808 = ~i_hbusreq1 & n5092;
  assign n9809 = ~n5317 & ~n9808;
  assign n9810 = ~controllable_ndecide & n9809;
  assign n9811 = ~controllable_ndecide & ~n9810;
  assign n9812 = i_hready & ~n9811;
  assign n9813 = ~n4577 & ~n9812;
  assign n9814 = i_hlock0 & ~n9813;
  assign n9815 = ~n8848 & ~n9814;
  assign n9816 = ~i_hbusreq0 & ~n9815;
  assign n9817 = ~n8845 & ~n9816;
  assign n9818 = ~i_hbusreq4 & ~n9817;
  assign n9819 = ~n8844 & ~n9818;
  assign n9820 = ~controllable_hgrant4 & ~n9819;
  assign n9821 = ~n4617 & ~n9820;
  assign n9822 = ~i_hbusreq2 & ~n9821;
  assign n9823 = ~n8843 & ~n9822;
  assign n9824 = ~controllable_hgrant2 & ~n9823;
  assign n9825 = ~n4562 & ~n9824;
  assign n9826 = controllable_hmaster0 & ~n9825;
  assign n9827 = ~n8827 & ~n9826;
  assign n9828 = ~controllable_hmaster1 & ~n9827;
  assign n9829 = ~n9807 & ~n9828;
  assign n9830 = ~i_hbusreq3 & ~n9829;
  assign n9831 = ~n8831 & ~n9830;
  assign n9832 = ~controllable_hmaster2 & ~n9831;
  assign n9833 = ~n9796 & ~n9832;
  assign n9834 = ~controllable_hgrant3 & ~n9833;
  assign n9835 = ~n9790 & ~n9834;
  assign n9836 = controllable_nhgrant0 & ~n9835;
  assign n9837 = ~n9699 & ~n9784;
  assign n9838 = ~i_hbusreq3 & ~n9837;
  assign n9839 = ~n3951 & ~n9838;
  assign n9840 = ~controllable_hmaster2 & ~n9839;
  assign n9841 = ~n9773 & ~n9840;
  assign n9842 = controllable_hgrant3 & ~n9841;
  assign n9843 = i_hbusreq3 & ~n4610;
  assign n9844 = ~i_hbusreq3 & ~n4635;
  assign n9845 = ~n9843 & ~n9844;
  assign n9846 = controllable_hmaster2 & ~n9845;
  assign n9847 = ~controllable_hmaster0 & ~n3500;
  assign n9848 = ~n9737 & ~n9847;
  assign n9849 = ~controllable_hmaster1 & ~n9848;
  assign n9850 = ~n9736 & ~n9849;
  assign n9851 = i_hbusreq3 & ~n9850;
  assign n9852 = ~n9743 & ~n9847;
  assign n9853 = ~controllable_hmaster1 & ~n9852;
  assign n9854 = ~n9742 & ~n9853;
  assign n9855 = ~i_hbusreq3 & ~n9854;
  assign n9856 = ~n9851 & ~n9855;
  assign n9857 = ~controllable_hmaster2 & ~n9856;
  assign n9858 = ~n9846 & ~n9857;
  assign n9859 = ~controllable_hgrant3 & ~n9858;
  assign n9860 = ~n9842 & ~n9859;
  assign n9861 = ~controllable_nhgrant0 & ~n9860;
  assign n9862 = ~n9836 & ~n9861;
  assign n9863 = ~n3281 & ~n9862;
  assign n9864 = ~n3281 & ~n9863;
  assign n9865 = ~n3378 & ~n9864;
  assign n9866 = ~n9770 & ~n9865;
  assign n9867 = n3492 & ~n9866;
  assign n9868 = n3492 & ~n9867;
  assign n9869 = n3485 & ~n9868;
  assign n9870 = n3485 & ~n9869;
  assign n9871 = ~n3476 & ~n9870;
  assign n9872 = ~n5039 & ~n5619;
  assign n9873 = ~controllable_hgrant4 & ~n9872;
  assign n9874 = ~n4091 & ~n9873;
  assign n9875 = ~controllable_hgrant2 & ~n9874;
  assign n9876 = ~n5616 & ~n9875;
  assign n9877 = controllable_hmaster1 & ~n9876;
  assign n9878 = controllable_hmaster0 & ~n9876;
  assign n9879 = ~n5630 & ~n9878;
  assign n9880 = ~controllable_hmaster1 & ~n9879;
  assign n9881 = ~n9877 & ~n9880;
  assign n9882 = i_hbusreq3 & ~n9881;
  assign n9883 = i_hbusreq2 & ~n9874;
  assign n9884 = i_hbusreq4 & ~n9872;
  assign n9885 = i_hbusreq0 & ~n9872;
  assign n9886 = ~n5055 & ~n5643;
  assign n9887 = i_hlock0 & ~n9886;
  assign n9888 = ~n5039 & ~n5869;
  assign n9889 = ~i_hlock0 & ~n9888;
  assign n9890 = ~n9887 & ~n9889;
  assign n9891 = ~i_hbusreq0 & ~n9890;
  assign n9892 = ~n9885 & ~n9891;
  assign n9893 = ~i_hbusreq4 & ~n9892;
  assign n9894 = ~n9884 & ~n9893;
  assign n9895 = ~controllable_hgrant4 & ~n9894;
  assign n9896 = ~n7486 & ~n9895;
  assign n9897 = ~i_hbusreq2 & ~n9896;
  assign n9898 = ~n9883 & ~n9897;
  assign n9899 = ~controllable_hgrant2 & ~n9898;
  assign n9900 = ~n5862 & ~n9899;
  assign n9901 = controllable_hmaster1 & ~n9900;
  assign n9902 = controllable_hmaster0 & ~n9900;
  assign n9903 = ~n4577 & ~n5643;
  assign n9904 = i_hlock0 & ~n9903;
  assign n9905 = ~n5891 & ~n9904;
  assign n9906 = ~i_hbusreq0 & ~n9905;
  assign n9907 = ~n5638 & ~n9906;
  assign n9908 = ~i_hbusreq4 & ~n9907;
  assign n9909 = ~n5637 & ~n9908;
  assign n9910 = ~controllable_hgrant4 & ~n9909;
  assign n9911 = ~n4667 & ~n9910;
  assign n9912 = ~i_hbusreq2 & ~n9911;
  assign n9913 = ~n5658 & ~n9912;
  assign n9914 = ~controllable_hgrant2 & ~n9913;
  assign n9915 = ~n7507 & ~n9914;
  assign n9916 = ~controllable_hmaster0 & ~n9915;
  assign n9917 = ~n9902 & ~n9916;
  assign n9918 = ~controllable_hmaster1 & ~n9917;
  assign n9919 = ~n9901 & ~n9918;
  assign n9920 = ~i_hbusreq3 & ~n9919;
  assign n9921 = ~n9882 & ~n9920;
  assign n9922 = controllable_hmaster2 & ~n9921;
  assign n9923 = ~n5943 & ~n7486;
  assign n9924 = ~i_hbusreq2 & ~n9923;
  assign n9925 = ~n5931 & ~n9924;
  assign n9926 = ~controllable_hgrant2 & ~n9925;
  assign n9927 = ~n5862 & ~n9926;
  assign n9928 = controllable_hmaster0 & ~n9927;
  assign n9929 = ~n5950 & ~n9926;
  assign n9930 = ~controllable_hmaster0 & ~n9929;
  assign n9931 = ~n9928 & ~n9930;
  assign n9932 = controllable_hmaster1 & ~n9931;
  assign n9933 = ~n5974 & ~n7486;
  assign n9934 = ~i_hbusreq2 & ~n9933;
  assign n9935 = ~n5955 & ~n9934;
  assign n9936 = ~controllable_hgrant2 & ~n9935;
  assign n9937 = ~n5862 & ~n9936;
  assign n9938 = controllable_hmaster0 & ~n9937;
  assign n9939 = ~n5990 & ~n7606;
  assign n9940 = ~i_hbusreq2 & ~n9939;
  assign n9941 = ~n5931 & ~n9940;
  assign n9942 = ~controllable_hgrant2 & ~n9941;
  assign n9943 = ~n5981 & ~n9942;
  assign n9944 = ~controllable_hmaster0 & ~n9943;
  assign n9945 = ~n9938 & ~n9944;
  assign n9946 = ~controllable_hmaster1 & ~n9945;
  assign n9947 = ~n9932 & ~n9946;
  assign n9948 = ~i_hbusreq3 & ~n9947;
  assign n9949 = ~n5930 & ~n9948;
  assign n9950 = ~controllable_hmaster2 & ~n9949;
  assign n9951 = ~n9922 & ~n9950;
  assign n9952 = ~controllable_hgrant3 & ~n9951;
  assign n9953 = ~n7457 & ~n9952;
  assign n9954 = controllable_nhgrant0 & ~n9953;
  assign n9955 = ~n3543 & ~n3904;
  assign n9956 = i_hlock0 & ~n9955;
  assign n9957 = ~n3494 & ~n3998;
  assign n9958 = i_hready & ~n9957;
  assign n9959 = ~n3904 & ~n9958;
  assign n9960 = ~i_hlock0 & ~n9959;
  assign n9961 = ~n9956 & ~n9960;
  assign n9962 = ~controllable_hgrant4 & ~n9961;
  assign n9963 = ~n3411 & ~n9962;
  assign n9964 = ~controllable_hgrant2 & ~n9963;
  assign n9965 = ~n3410 & ~n9964;
  assign n9966 = controllable_hmaster1 & ~n9965;
  assign n9967 = controllable_hmaster0 & ~n9965;
  assign n9968 = ~n3543 & ~n4605;
  assign n9969 = i_hlock0 & ~n9968;
  assign n9970 = ~n4605 & ~n9958;
  assign n9971 = ~i_hlock0 & ~n9970;
  assign n9972 = ~n9969 & ~n9971;
  assign n9973 = ~controllable_hgrant4 & ~n9972;
  assign n9974 = ~n3411 & ~n9973;
  assign n9975 = ~controllable_hgrant2 & ~n9974;
  assign n9976 = ~n3410 & ~n9975;
  assign n9977 = ~controllable_hmaster0 & ~n9976;
  assign n9978 = ~n9967 & ~n9977;
  assign n9979 = ~controllable_hmaster1 & ~n9978;
  assign n9980 = ~n9966 & ~n9979;
  assign n9981 = i_hbusreq3 & ~n9980;
  assign n9982 = i_hbusreq2 & ~n9963;
  assign n9983 = i_hbusreq4 & ~n9961;
  assign n9984 = i_hbusreq0 & ~n9961;
  assign n9985 = ~controllable_hgrant1 & ~n5960;
  assign n9986 = ~i_hbusreq1 & ~n9985;
  assign n9987 = ~n3564 & ~n9986;
  assign n9988 = ~controllable_ndecide & ~n9987;
  assign n9989 = ~n3494 & ~n9988;
  assign n9990 = i_hready & ~n9989;
  assign n9991 = ~n3920 & ~n9990;
  assign n9992 = i_hlock0 & ~n9991;
  assign n9993 = ~n9960 & ~n9992;
  assign n9994 = ~i_hbusreq0 & ~n9993;
  assign n9995 = ~n9984 & ~n9994;
  assign n9996 = ~i_hbusreq4 & ~n9995;
  assign n9997 = ~n9983 & ~n9996;
  assign n9998 = ~controllable_hgrant4 & ~n9997;
  assign n9999 = ~n3916 & ~n9998;
  assign n10000 = ~i_hbusreq2 & ~n9999;
  assign n10001 = ~n9982 & ~n10000;
  assign n10002 = ~controllable_hgrant2 & ~n10001;
  assign n10003 = ~n3859 & ~n10002;
  assign n10004 = controllable_hmaster1 & ~n10003;
  assign n10005 = controllable_hmaster0 & ~n10003;
  assign n10006 = i_hbusreq2 & ~n9974;
  assign n10007 = i_hbusreq4 & ~n9972;
  assign n10008 = i_hbusreq0 & ~n9972;
  assign n10009 = ~n4621 & ~n9990;
  assign n10010 = i_hlock0 & ~n10009;
  assign n10011 = ~n9971 & ~n10010;
  assign n10012 = ~i_hbusreq0 & ~n10011;
  assign n10013 = ~n10008 & ~n10012;
  assign n10014 = ~i_hbusreq4 & ~n10013;
  assign n10015 = ~n10007 & ~n10014;
  assign n10016 = ~controllable_hgrant4 & ~n10015;
  assign n10017 = ~n4617 & ~n10016;
  assign n10018 = ~i_hbusreq2 & ~n10017;
  assign n10019 = ~n10006 & ~n10018;
  assign n10020 = ~controllable_hgrant2 & ~n10019;
  assign n10021 = ~n4562 & ~n10020;
  assign n10022 = ~controllable_hmaster0 & ~n10021;
  assign n10023 = ~n10005 & ~n10022;
  assign n10024 = ~controllable_hmaster1 & ~n10023;
  assign n10025 = ~n10004 & ~n10024;
  assign n10026 = ~i_hbusreq3 & ~n10025;
  assign n10027 = ~n9981 & ~n10026;
  assign n10028 = controllable_hmaster2 & ~n10027;
  assign n10029 = ~n3543 & ~n5039;
  assign n10030 = i_hlock0 & ~n10029;
  assign n10031 = ~n3494 & ~n4011;
  assign n10032 = i_hready & ~n10031;
  assign n10033 = ~n5039 & ~n10032;
  assign n10034 = ~i_hlock0 & ~n10033;
  assign n10035 = ~n10030 & ~n10034;
  assign n10036 = ~controllable_hgrant4 & ~n10035;
  assign n10037 = ~n3411 & ~n10036;
  assign n10038 = ~controllable_hgrant2 & ~n10037;
  assign n10039 = ~n3410 & ~n10038;
  assign n10040 = ~controllable_hmaster0 & ~n10039;
  assign n10041 = ~n9967 & ~n10040;
  assign n10042 = ~controllable_hmaster1 & ~n10041;
  assign n10043 = ~n9966 & ~n10042;
  assign n10044 = i_hbusreq3 & ~n10043;
  assign n10045 = i_hbusreq2 & ~n10037;
  assign n10046 = i_hbusreq4 & ~n10035;
  assign n10047 = i_hbusreq0 & ~n10035;
  assign n10048 = ~n5510 & ~n9990;
  assign n10049 = i_hlock0 & ~n10048;
  assign n10050 = ~n10034 & ~n10049;
  assign n10051 = ~i_hbusreq0 & ~n10050;
  assign n10052 = ~n10047 & ~n10051;
  assign n10053 = ~i_hbusreq4 & ~n10052;
  assign n10054 = ~n10046 & ~n10053;
  assign n10055 = ~controllable_hgrant4 & ~n10054;
  assign n10056 = ~n5462 & ~n10055;
  assign n10057 = ~i_hbusreq2 & ~n10056;
  assign n10058 = ~n10045 & ~n10057;
  assign n10059 = ~controllable_hgrant2 & ~n10058;
  assign n10060 = ~n5461 & ~n10059;
  assign n10061 = ~controllable_hmaster0 & ~n10060;
  assign n10062 = ~n10005 & ~n10061;
  assign n10063 = ~controllable_hmaster1 & ~n10062;
  assign n10064 = ~n10004 & ~n10063;
  assign n10065 = ~i_hbusreq3 & ~n10064;
  assign n10066 = ~n10044 & ~n10065;
  assign n10067 = ~controllable_hmaster2 & ~n10066;
  assign n10068 = ~n10028 & ~n10067;
  assign n10069 = ~controllable_hgrant3 & ~n10068;
  assign n10070 = ~n7194 & ~n10069;
  assign n10071 = ~controllable_nhgrant0 & ~n10070;
  assign n10072 = ~n9954 & ~n10071;
  assign n10073 = ~n3281 & ~n10072;
  assign n10074 = ~n3281 & ~n10073;
  assign n10075 = n3378 & ~n10074;
  assign n10076 = ~n4000 & ~n4543;
  assign n10077 = i_hlock0 & ~n10076;
  assign n10078 = ~n5814 & ~n10077;
  assign n10079 = ~i_hbusreq0 & ~n10078;
  assign n10080 = ~n4107 & ~n10079;
  assign n10081 = ~i_hbusreq4 & ~n10080;
  assign n10082 = ~n4106 & ~n10081;
  assign n10083 = ~controllable_hgrant4 & ~n10082;
  assign n10084 = ~n4617 & ~n10083;
  assign n10085 = ~i_hbusreq2 & ~n10084;
  assign n10086 = ~n5550 & ~n10085;
  assign n10087 = ~controllable_hgrant2 & ~n10086;
  assign n10088 = ~n4562 & ~n10087;
  assign n10089 = ~i_hbusreq3 & ~n10088;
  assign n10090 = ~n5549 & ~n10089;
  assign n10091 = controllable_hmaster2 & ~n10090;
  assign n10092 = ~controllable_hgrant4 & ~n4666;
  assign n10093 = ~n4617 & ~n10092;
  assign n10094 = ~i_hbusreq2 & ~n10093;
  assign n10095 = ~n5594 & ~n10094;
  assign n10096 = ~controllable_hgrant2 & ~n10095;
  assign n10097 = ~n4562 & ~n10096;
  assign n10098 = controllable_hmaster0 & ~n10097;
  assign n10099 = ~controllable_hmaster0 & ~n10088;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = controllable_hmaster1 & ~n10100;
  assign n10102 = controllable_hmaster0 & ~n10088;
  assign n10103 = ~n5588 & ~n10102;
  assign n10104 = ~controllable_hmaster1 & ~n10103;
  assign n10105 = ~n10101 & ~n10104;
  assign n10106 = ~i_hbusreq3 & ~n10105;
  assign n10107 = ~n5593 & ~n10106;
  assign n10108 = ~controllable_hmaster2 & ~n10107;
  assign n10109 = ~n10091 & ~n10108;
  assign n10110 = controllable_hgrant3 & ~n10109;
  assign n10111 = controllable_hgrant2 & ~n10086;
  assign n10112 = controllable_hgrant4 & ~n10082;
  assign n10113 = ~n4577 & ~n5889;
  assign n10114 = i_hlock0 & ~n10113;
  assign n10115 = ~n5871 & ~n10114;
  assign n10116 = ~i_hbusreq0 & ~n10115;
  assign n10117 = ~n5638 & ~n10116;
  assign n10118 = ~i_hbusreq4 & ~n10117;
  assign n10119 = ~n5637 & ~n10118;
  assign n10120 = ~controllable_hgrant4 & ~n10119;
  assign n10121 = ~n10112 & ~n10120;
  assign n10122 = ~i_hbusreq2 & ~n10121;
  assign n10123 = ~n5636 & ~n10122;
  assign n10124 = ~controllable_hgrant2 & ~n10123;
  assign n10125 = ~n10111 & ~n10124;
  assign n10126 = controllable_hmaster1 & ~n10125;
  assign n10127 = controllable_hmaster0 & ~n10125;
  assign n10128 = ~n5891 & ~n10114;
  assign n10129 = ~i_hbusreq0 & ~n10128;
  assign n10130 = ~n5638 & ~n10129;
  assign n10131 = ~i_hbusreq4 & ~n10130;
  assign n10132 = ~n5637 & ~n10131;
  assign n10133 = ~controllable_hgrant4 & ~n10132;
  assign n10134 = ~n4667 & ~n10133;
  assign n10135 = ~i_hbusreq2 & ~n10134;
  assign n10136 = ~n5658 & ~n10135;
  assign n10137 = ~controllable_hgrant2 & ~n10136;
  assign n10138 = ~n10111 & ~n10137;
  assign n10139 = ~controllable_hmaster0 & ~n10138;
  assign n10140 = ~n10127 & ~n10139;
  assign n10141 = ~controllable_hmaster1 & ~n10140;
  assign n10142 = ~n10126 & ~n10141;
  assign n10143 = ~i_hbusreq3 & ~n10142;
  assign n10144 = ~n5634 & ~n10143;
  assign n10145 = controllable_hmaster2 & ~n10144;
  assign n10146 = ~n10112 & ~n10133;
  assign n10147 = ~i_hbusreq2 & ~n10146;
  assign n10148 = ~n5636 & ~n10147;
  assign n10149 = ~controllable_hgrant2 & ~n10148;
  assign n10150 = ~n10111 & ~n10149;
  assign n10151 = controllable_hmaster0 & ~n10150;
  assign n10152 = controllable_hgrant2 & ~n10095;
  assign n10153 = ~n10149 & ~n10152;
  assign n10154 = ~controllable_hmaster0 & ~n10153;
  assign n10155 = ~n10151 & ~n10154;
  assign n10156 = controllable_hmaster1 & ~n10155;
  assign n10157 = ~i_hbusreq1 & ~controllable_locked;
  assign n10158 = ~n5730 & ~n10157;
  assign n10159 = ~controllable_ndecide & n10158;
  assign n10160 = ~n3494 & ~n10159;
  assign n10161 = i_hready & ~n10160;
  assign n10162 = ~n4577 & ~n10161;
  assign n10163 = i_hlock0 & ~n10162;
  assign n10164 = ~n9018 & ~n10163;
  assign n10165 = ~i_hbusreq0 & ~n10164;
  assign n10166 = ~n9009 & ~n10165;
  assign n10167 = ~i_hbusreq4 & ~n10166;
  assign n10168 = ~n9008 & ~n10167;
  assign n10169 = ~controllable_hgrant4 & ~n10168;
  assign n10170 = ~n10112 & ~n10169;
  assign n10171 = ~i_hbusreq2 & ~n10170;
  assign n10172 = ~n9007 & ~n10171;
  assign n10173 = ~controllable_hgrant2 & ~n10172;
  assign n10174 = ~n10111 & ~n10173;
  assign n10175 = controllable_hmaster0 & ~n10174;
  assign n10176 = ~i_hbusreq0 & ~n5890;
  assign n10177 = ~n5638 & ~n10176;
  assign n10178 = ~i_hbusreq4 & ~n10177;
  assign n10179 = ~n5637 & ~n10178;
  assign n10180 = ~controllable_hgrant4 & ~n10179;
  assign n10181 = ~n4091 & ~n10180;
  assign n10182 = ~i_hbusreq2 & ~n10181;
  assign n10183 = ~n5636 & ~n10182;
  assign n10184 = ~controllable_hgrant2 & ~n10183;
  assign n10185 = ~n5616 & ~n10184;
  assign n10186 = ~controllable_hmaster0 & ~n10185;
  assign n10187 = ~n10175 & ~n10186;
  assign n10188 = ~controllable_hmaster1 & ~n10187;
  assign n10189 = ~n10156 & ~n10188;
  assign n10190 = ~i_hbusreq3 & ~n10189;
  assign n10191 = ~n8996 & ~n10190;
  assign n10192 = ~controllable_hmaster2 & ~n10191;
  assign n10193 = ~n10145 & ~n10192;
  assign n10194 = ~controllable_hgrant3 & ~n10193;
  assign n10195 = ~n10110 & ~n10194;
  assign n10196 = controllable_nhgrant0 & ~n10195;
  assign n10197 = i_hbusreq3 & ~n9976;
  assign n10198 = ~n3543 & ~n4621;
  assign n10199 = i_hlock0 & ~n10198;
  assign n10200 = ~n9971 & ~n10199;
  assign n10201 = ~i_hbusreq0 & ~n10200;
  assign n10202 = ~n10008 & ~n10201;
  assign n10203 = ~i_hbusreq4 & ~n10202;
  assign n10204 = ~n10007 & ~n10203;
  assign n10205 = ~controllable_hgrant4 & ~n10204;
  assign n10206 = ~n4617 & ~n10205;
  assign n10207 = ~i_hbusreq2 & ~n10206;
  assign n10208 = ~n10006 & ~n10207;
  assign n10209 = ~controllable_hgrant2 & ~n10208;
  assign n10210 = ~n4562 & ~n10209;
  assign n10211 = ~i_hbusreq3 & ~n10210;
  assign n10212 = ~n10197 & ~n10211;
  assign n10213 = controllable_hmaster2 & ~n10212;
  assign n10214 = controllable_hmaster1 & ~n9976;
  assign n10215 = controllable_hmaster0 & ~n9976;
  assign n10216 = i_hlock0 & ~n3544;
  assign n10217 = ~n3495 & ~n10032;
  assign n10218 = ~i_hlock0 & ~n10217;
  assign n10219 = ~n10216 & ~n10218;
  assign n10220 = ~controllable_hgrant4 & ~n10219;
  assign n10221 = ~n3411 & ~n10220;
  assign n10222 = ~controllable_hgrant2 & ~n10221;
  assign n10223 = ~n3410 & ~n10222;
  assign n10224 = ~controllable_hmaster0 & ~n10223;
  assign n10225 = ~n10215 & ~n10224;
  assign n10226 = ~controllable_hmaster1 & ~n10225;
  assign n10227 = ~n10214 & ~n10226;
  assign n10228 = i_hbusreq3 & ~n10227;
  assign n10229 = controllable_hmaster1 & ~n10210;
  assign n10230 = controllable_hmaster0 & ~n10210;
  assign n10231 = ~n10224 & ~n10230;
  assign n10232 = ~controllable_hmaster1 & ~n10231;
  assign n10233 = ~n10229 & ~n10232;
  assign n10234 = ~i_hbusreq3 & ~n10233;
  assign n10235 = ~n10228 & ~n10234;
  assign n10236 = ~controllable_hmaster2 & ~n10235;
  assign n10237 = ~n10213 & ~n10236;
  assign n10238 = ~controllable_hgrant3 & ~n10237;
  assign n10239 = ~n9842 & ~n10238;
  assign n10240 = ~controllable_nhgrant0 & ~n10239;
  assign n10241 = ~n10196 & ~n10240;
  assign n10242 = ~n3281 & ~n10241;
  assign n10243 = ~n3281 & ~n10242;
  assign n10244 = ~n3378 & ~n10243;
  assign n10245 = ~n10075 & ~n10244;
  assign n10246 = n3492 & ~n10245;
  assign n10247 = ~n8536 & ~n10246;
  assign n10248 = n3485 & ~n10247;
  assign n10249 = ~n8694 & ~n10248;
  assign n10250 = n3476 & ~n10249;
  assign n10251 = ~n9871 & ~n10250;
  assign n10252 = n3374 & ~n10251;
  assign n10253 = ~n9769 & ~n10252;
  assign n10254 = n3655 & ~n10253;
  assign n10255 = n3378 & ~n7699;
  assign n10256 = ~n3417 & ~n4699;
  assign n10257 = ~controllable_hgrant4 & ~n10256;
  assign n10258 = ~n3411 & ~n10257;
  assign n10259 = ~controllable_hgrant2 & ~n10258;
  assign n10260 = ~n3410 & ~n10259;
  assign n10261 = controllable_hmaster1 & ~n10260;
  assign n10262 = controllable_hmaster0 & ~n10260;
  assign n10263 = controllable_hmaster0 & ~n10262;
  assign n10264 = ~controllable_hmaster1 & ~n10263;
  assign n10265 = ~n10261 & ~n10264;
  assign n10266 = i_hbusreq3 & ~n10265;
  assign n10267 = i_hbusreq2 & ~n10258;
  assign n10268 = i_hbusreq4 & ~n10256;
  assign n10269 = i_hbusreq0 & ~n10256;
  assign n10270 = ~n4714 & ~n9710;
  assign n10271 = i_hlock0 & ~n10270;
  assign n10272 = ~i_hlock0 & ~n10256;
  assign n10273 = ~n10271 & ~n10272;
  assign n10274 = ~i_hbusreq0 & ~n10273;
  assign n10275 = ~n10269 & ~n10274;
  assign n10276 = ~i_hbusreq4 & ~n10275;
  assign n10277 = ~n10268 & ~n10276;
  assign n10278 = ~controllable_hgrant4 & ~n10277;
  assign n10279 = ~n4617 & ~n10278;
  assign n10280 = ~i_hbusreq2 & ~n10279;
  assign n10281 = ~n10267 & ~n10280;
  assign n10282 = ~controllable_hgrant2 & ~n10281;
  assign n10283 = ~n4562 & ~n10282;
  assign n10284 = controllable_hmaster1 & ~n10283;
  assign n10285 = controllable_hmaster0 & ~n10283;
  assign n10286 = controllable_hmaster0 & ~n10285;
  assign n10287 = ~controllable_hmaster1 & ~n10286;
  assign n10288 = ~n10284 & ~n10287;
  assign n10289 = ~i_hbusreq3 & ~n10288;
  assign n10290 = ~n10266 & ~n10289;
  assign n10291 = controllable_hmaster2 & ~n10290;
  assign n10292 = controllable_hmaster2 & ~n10291;
  assign n10293 = ~controllable_hgrant3 & ~n10292;
  assign n10294 = ~n9708 & ~n10293;
  assign n10295 = controllable_nhgrant0 & ~n10294;
  assign n10296 = ~n9753 & ~n10295;
  assign n10297 = ~n3281 & ~n10296;
  assign n10298 = ~n3281 & ~n10297;
  assign n10299 = ~n3378 & ~n10298;
  assign n10300 = ~n10255 & ~n10299;
  assign n10301 = n3492 & ~n10300;
  assign n10302 = n3492 & ~n10301;
  assign n10303 = n3485 & ~n10302;
  assign n10304 = n3485 & ~n10303;
  assign n10305 = ~n3476 & ~n10304;
  assign n10306 = ~n8523 & ~n10301;
  assign n10307 = n3485 & ~n10306;
  assign n10308 = ~n8689 & ~n10307;
  assign n10309 = n3476 & ~n10308;
  assign n10310 = ~n10305 & ~n10309;
  assign n10311 = ~n3374 & ~n10310;
  assign n10312 = n3378 & ~n7741;
  assign n10313 = ~n4705 & ~n10262;
  assign n10314 = ~controllable_hmaster1 & ~n10313;
  assign n10315 = ~n10261 & ~n10314;
  assign n10316 = i_hbusreq3 & ~n10315;
  assign n10317 = ~n4729 & ~n10285;
  assign n10318 = ~controllable_hmaster1 & ~n10317;
  assign n10319 = ~n10284 & ~n10318;
  assign n10320 = ~i_hbusreq3 & ~n10319;
  assign n10321 = ~n10316 & ~n10320;
  assign n10322 = controllable_hmaster2 & ~n10321;
  assign n10323 = ~n3411 & ~n4701;
  assign n10324 = ~controllable_hgrant2 & ~n10323;
  assign n10325 = ~n3410 & ~n10324;
  assign n10326 = controllable_hmaster0 & ~n10325;
  assign n10327 = ~n5288 & ~n10324;
  assign n10328 = ~controllable_hmaster0 & ~n10327;
  assign n10329 = ~n10326 & ~n10328;
  assign n10330 = controllable_hmaster1 & ~n10329;
  assign n10331 = i_hready & ~n6259;
  assign n10332 = ~controllable_hgrant4 & n10331;
  assign n10333 = ~n3411 & ~n10332;
  assign n10334 = ~controllable_hgrant2 & ~n10333;
  assign n10335 = ~n3410 & ~n10334;
  assign n10336 = controllable_hmaster0 & ~n10335;
  assign n10337 = ~controllable_hmaster0 & ~n10325;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = ~controllable_hmaster1 & ~n10338;
  assign n10340 = ~n10330 & ~n10339;
  assign n10341 = i_hbusreq3 & ~n10340;
  assign n10342 = i_hbusreq2 & ~n10323;
  assign n10343 = ~n4617 & ~n4723;
  assign n10344 = ~i_hbusreq2 & ~n10343;
  assign n10345 = ~n10342 & ~n10344;
  assign n10346 = ~controllable_hgrant2 & ~n10345;
  assign n10347 = ~n4562 & ~n10346;
  assign n10348 = controllable_hmaster0 & ~n10347;
  assign n10349 = ~n9803 & ~n10346;
  assign n10350 = ~controllable_hmaster0 & ~n10349;
  assign n10351 = ~n10348 & ~n10350;
  assign n10352 = controllable_hmaster1 & ~n10351;
  assign n10353 = i_hbusreq2 & ~n10333;
  assign n10354 = i_hbusreq4 & ~n10331;
  assign n10355 = i_hbusreq0 & ~n10331;
  assign n10356 = ~controllable_ndecide & ~n9809;
  assign n10357 = ~n6137 & ~n10356;
  assign n10358 = i_hready & ~n10357;
  assign n10359 = ~controllable_ndecide & ~n4540;
  assign n10360 = ~controllable_ndecide & ~n10359;
  assign n10361 = ~i_hready & ~n10360;
  assign n10362 = ~n10358 & ~n10361;
  assign n10363 = i_hlock0 & ~n10362;
  assign n10364 = ~i_hlock0 & ~n10331;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = ~i_hbusreq0 & ~n10365;
  assign n10367 = ~n10355 & ~n10366;
  assign n10368 = ~i_hbusreq4 & ~n10367;
  assign n10369 = ~n10354 & ~n10368;
  assign n10370 = ~controllable_hgrant4 & n10369;
  assign n10371 = ~n4617 & ~n10370;
  assign n10372 = ~i_hbusreq2 & ~n10371;
  assign n10373 = ~n10353 & ~n10372;
  assign n10374 = ~controllable_hgrant2 & ~n10373;
  assign n10375 = ~n4562 & ~n10374;
  assign n10376 = controllable_hmaster0 & ~n10375;
  assign n10377 = ~n10337 & ~n10376;
  assign n10378 = ~controllable_hmaster1 & ~n10377;
  assign n10379 = ~n10352 & ~n10378;
  assign n10380 = ~i_hbusreq3 & ~n10379;
  assign n10381 = ~n10341 & ~n10380;
  assign n10382 = ~controllable_hmaster2 & ~n10381;
  assign n10383 = ~n10322 & ~n10382;
  assign n10384 = ~controllable_hgrant3 & ~n10383;
  assign n10385 = ~n9790 & ~n10384;
  assign n10386 = controllable_nhgrant0 & ~n10385;
  assign n10387 = ~n9861 & ~n10386;
  assign n10388 = ~n3281 & ~n10387;
  assign n10389 = ~n3281 & ~n10388;
  assign n10390 = ~n3378 & ~n10389;
  assign n10391 = ~n10312 & ~n10390;
  assign n10392 = n3492 & ~n10391;
  assign n10393 = n3492 & ~n10392;
  assign n10394 = n3485 & ~n10393;
  assign n10395 = n3485 & ~n10394;
  assign n10396 = ~n3476 & ~n10395;
  assign n10397 = ~i_hlock1 & ~n4178;
  assign n10398 = ~i_hlock1 & ~n10397;
  assign n10399 = ~controllable_ndecide & ~n10398;
  assign n10400 = ~controllable_ndecide & ~n10399;
  assign n10401 = i_hready & ~n10400;
  assign n10402 = ~i_hready & ~n6097;
  assign n10403 = ~n10401 & ~n10402;
  assign n10404 = ~controllable_hgrant4 & n10403;
  assign n10405 = ~n4091 & ~n10404;
  assign n10406 = ~controllable_hgrant2 & ~n10405;
  assign n10407 = ~n5616 & ~n10406;
  assign n10408 = controllable_hmaster1 & ~n10407;
  assign n10409 = controllable_hmaster0 & ~n10407;
  assign n10410 = ~i_hready & ~n4698;
  assign n10411 = ~n10401 & ~n10410;
  assign n10412 = ~controllable_hgrant4 & n10411;
  assign n10413 = ~n4015 & ~n10412;
  assign n10414 = ~controllable_hgrant2 & ~n10413;
  assign n10415 = ~n5616 & ~n10414;
  assign n10416 = ~controllable_hmaster0 & ~n10415;
  assign n10417 = ~n10409 & ~n10416;
  assign n10418 = ~controllable_hmaster1 & ~n10417;
  assign n10419 = ~n10408 & ~n10418;
  assign n10420 = i_hbusreq3 & ~n10419;
  assign n10421 = i_hbusreq2 & ~n10405;
  assign n10422 = i_hbusreq4 & ~n10403;
  assign n10423 = i_hbusreq0 & ~n10403;
  assign n10424 = i_hbusreq1 & ~n10398;
  assign n10425 = ~controllable_ndecide & n10424;
  assign n10426 = ~controllable_ndecide & ~n10425;
  assign n10427 = i_hready & ~n10426;
  assign n10428 = ~i_hready & n6113;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = i_hlock0 & ~n10429;
  assign n10431 = ~i_hbusreq1 & n5864;
  assign n10432 = ~n10424 & ~n10431;
  assign n10433 = ~controllable_ndecide & ~n10432;
  assign n10434 = ~controllable_ndecide & ~n10433;
  assign n10435 = i_hready & ~n10434;
  assign n10436 = ~n10402 & ~n10435;
  assign n10437 = ~i_hlock0 & ~n10436;
  assign n10438 = ~n10430 & ~n10437;
  assign n10439 = ~i_hbusreq0 & ~n10438;
  assign n10440 = ~n10423 & ~n10439;
  assign n10441 = ~i_hbusreq4 & ~n10440;
  assign n10442 = ~n10422 & ~n10441;
  assign n10443 = ~controllable_hgrant4 & n10442;
  assign n10444 = ~n7486 & ~n10443;
  assign n10445 = ~i_hbusreq2 & ~n10444;
  assign n10446 = ~n10421 & ~n10445;
  assign n10447 = ~controllable_hgrant2 & ~n10446;
  assign n10448 = ~n5862 & ~n10447;
  assign n10449 = controllable_hmaster1 & ~n10448;
  assign n10450 = controllable_hmaster0 & ~n10448;
  assign n10451 = i_hbusreq2 & ~n10413;
  assign n10452 = i_hbusreq4 & ~n10411;
  assign n10453 = i_hbusreq0 & ~n10411;
  assign n10454 = ~i_hready & n4713;
  assign n10455 = ~n10427 & ~n10454;
  assign n10456 = i_hlock0 & ~n10455;
  assign n10457 = ~n10157 & ~n10424;
  assign n10458 = ~controllable_ndecide & ~n10457;
  assign n10459 = ~controllable_ndecide & ~n10458;
  assign n10460 = i_hready & ~n10459;
  assign n10461 = ~n10410 & ~n10460;
  assign n10462 = ~i_hlock0 & ~n10461;
  assign n10463 = ~n10456 & ~n10462;
  assign n10464 = ~i_hbusreq0 & ~n10463;
  assign n10465 = ~n10453 & ~n10464;
  assign n10466 = ~i_hbusreq4 & ~n10465;
  assign n10467 = ~n10452 & ~n10466;
  assign n10468 = ~controllable_hgrant4 & n10467;
  assign n10469 = ~n4667 & ~n10468;
  assign n10470 = ~i_hbusreq2 & ~n10469;
  assign n10471 = ~n10451 & ~n10470;
  assign n10472 = ~controllable_hgrant2 & ~n10471;
  assign n10473 = ~n7507 & ~n10472;
  assign n10474 = ~controllable_hmaster0 & ~n10473;
  assign n10475 = ~n10450 & ~n10474;
  assign n10476 = ~controllable_hmaster1 & ~n10475;
  assign n10477 = ~n10449 & ~n10476;
  assign n10478 = ~i_hbusreq3 & ~n10477;
  assign n10479 = ~n10420 & ~n10478;
  assign n10480 = controllable_hmaster2 & ~n10479;
  assign n10481 = ~i_hready & ~n6247;
  assign n10482 = ~n10401 & ~n10481;
  assign n10483 = ~controllable_hgrant4 & n10482;
  assign n10484 = ~n4091 & ~n10483;
  assign n10485 = ~controllable_hgrant2 & ~n10484;
  assign n10486 = ~n5616 & ~n10485;
  assign n10487 = controllable_hmaster0 & ~n10486;
  assign n10488 = ~n5686 & ~n10485;
  assign n10489 = ~controllable_hmaster0 & ~n10488;
  assign n10490 = ~n10487 & ~n10489;
  assign n10491 = controllable_hmaster1 & ~n10490;
  assign n10492 = ~i_hlock1 & ~n5692;
  assign n10493 = ~i_hlock1 & ~n10492;
  assign n10494 = ~controllable_ndecide & ~n10493;
  assign n10495 = ~controllable_ndecide & ~n10494;
  assign n10496 = i_hready & ~n10495;
  assign n10497 = ~n6262 & ~n10496;
  assign n10498 = ~controllable_hgrant4 & n10497;
  assign n10499 = ~n4091 & ~n10498;
  assign n10500 = ~controllable_hgrant2 & ~n10499;
  assign n10501 = ~n5616 & ~n10500;
  assign n10502 = controllable_hmaster0 & ~n10501;
  assign n10503 = ~controllable_hmaster0 & ~n10486;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = ~controllable_hmaster1 & ~n10504;
  assign n10506 = ~n10491 & ~n10505;
  assign n10507 = i_hbusreq3 & ~n10506;
  assign n10508 = i_hbusreq2 & ~n10484;
  assign n10509 = i_hbusreq4 & ~n10482;
  assign n10510 = i_hbusreq0 & ~n10482;
  assign n10511 = ~i_hready & n6277;
  assign n10512 = ~n10427 & ~n10511;
  assign n10513 = i_hlock0 & ~n10512;
  assign n10514 = ~n10460 & ~n10481;
  assign n10515 = ~i_hlock0 & ~n10514;
  assign n10516 = ~n10513 & ~n10515;
  assign n10517 = ~i_hbusreq0 & ~n10516;
  assign n10518 = ~n10510 & ~n10517;
  assign n10519 = ~i_hbusreq4 & ~n10518;
  assign n10520 = ~n10509 & ~n10519;
  assign n10521 = ~controllable_hgrant4 & n10520;
  assign n10522 = ~n7486 & ~n10521;
  assign n10523 = ~i_hbusreq2 & ~n10522;
  assign n10524 = ~n10508 & ~n10523;
  assign n10525 = ~controllable_hgrant2 & ~n10524;
  assign n10526 = ~n5862 & ~n10525;
  assign n10527 = controllable_hmaster0 & ~n10526;
  assign n10528 = ~n5950 & ~n10525;
  assign n10529 = ~controllable_hmaster0 & ~n10528;
  assign n10530 = ~n10527 & ~n10529;
  assign n10531 = controllable_hmaster1 & ~n10530;
  assign n10532 = i_hbusreq2 & ~n10499;
  assign n10533 = i_hbusreq4 & ~n10497;
  assign n10534 = i_hbusreq0 & ~n10497;
  assign n10535 = i_hbusreq1 & ~n10493;
  assign n10536 = ~controllable_ndecide & n10535;
  assign n10537 = ~controllable_ndecide & ~n10536;
  assign n10538 = i_hready & ~n10537;
  assign n10539 = ~n6306 & ~n10538;
  assign n10540 = i_hlock0 & ~n10539;
  assign n10541 = ~n5962 & ~n10535;
  assign n10542 = ~controllable_ndecide & ~n10541;
  assign n10543 = ~controllable_ndecide & ~n10542;
  assign n10544 = i_hready & ~n10543;
  assign n10545 = ~n6262 & ~n10544;
  assign n10546 = ~i_hlock0 & ~n10545;
  assign n10547 = ~n10540 & ~n10546;
  assign n10548 = ~i_hbusreq0 & ~n10547;
  assign n10549 = ~n10534 & ~n10548;
  assign n10550 = ~i_hbusreq4 & ~n10549;
  assign n10551 = ~n10533 & ~n10550;
  assign n10552 = ~controllable_hgrant4 & n10551;
  assign n10553 = ~n7486 & ~n10552;
  assign n10554 = ~i_hbusreq2 & ~n10553;
  assign n10555 = ~n10532 & ~n10554;
  assign n10556 = ~controllable_hgrant2 & ~n10555;
  assign n10557 = ~n5862 & ~n10556;
  assign n10558 = controllable_hmaster0 & ~n10557;
  assign n10559 = ~i_hready & n6322;
  assign n10560 = ~n10427 & ~n10559;
  assign n10561 = i_hlock0 & ~n10560;
  assign n10562 = ~n10515 & ~n10561;
  assign n10563 = ~i_hbusreq0 & ~n10562;
  assign n10564 = ~n10510 & ~n10563;
  assign n10565 = ~i_hbusreq4 & ~n10564;
  assign n10566 = ~n10509 & ~n10565;
  assign n10567 = ~controllable_hgrant4 & n10566;
  assign n10568 = ~n7606 & ~n10567;
  assign n10569 = ~i_hbusreq2 & ~n10568;
  assign n10570 = ~n10508 & ~n10569;
  assign n10571 = ~controllable_hgrant2 & ~n10570;
  assign n10572 = ~n5981 & ~n10571;
  assign n10573 = ~controllable_hmaster0 & ~n10572;
  assign n10574 = ~n10558 & ~n10573;
  assign n10575 = ~controllable_hmaster1 & ~n10574;
  assign n10576 = ~n10531 & ~n10575;
  assign n10577 = ~i_hbusreq3 & ~n10576;
  assign n10578 = ~n10507 & ~n10577;
  assign n10579 = ~controllable_hmaster2 & ~n10578;
  assign n10580 = ~n10480 & ~n10579;
  assign n10581 = ~controllable_hgrant3 & ~n10580;
  assign n10582 = ~n7457 & ~n10581;
  assign n10583 = controllable_nhgrant0 & ~n10582;
  assign n10584 = ~n10071 & ~n10583;
  assign n10585 = ~n3281 & ~n10584;
  assign n10586 = ~n3281 & ~n10585;
  assign n10587 = n3378 & ~n10586;
  assign n10588 = ~n4091 & ~n10412;
  assign n10589 = ~controllable_hgrant2 & ~n10588;
  assign n10590 = ~n5616 & ~n10589;
  assign n10591 = controllable_hmaster1 & ~n10590;
  assign n10592 = controllable_hmaster0 & ~n10590;
  assign n10593 = ~n10416 & ~n10592;
  assign n10594 = ~controllable_hmaster1 & ~n10593;
  assign n10595 = ~n10591 & ~n10594;
  assign n10596 = i_hbusreq3 & ~n10595;
  assign n10597 = i_hbusreq2 & ~n10588;
  assign n10598 = ~n10454 & ~n10460;
  assign n10599 = i_hlock0 & ~n10598;
  assign n10600 = ~n10410 & ~n10435;
  assign n10601 = ~i_hlock0 & ~n10600;
  assign n10602 = ~n10599 & ~n10601;
  assign n10603 = ~i_hbusreq0 & ~n10602;
  assign n10604 = ~n10453 & ~n10603;
  assign n10605 = ~i_hbusreq4 & ~n10604;
  assign n10606 = ~n10452 & ~n10605;
  assign n10607 = ~controllable_hgrant4 & n10606;
  assign n10608 = ~n10112 & ~n10607;
  assign n10609 = ~i_hbusreq2 & ~n10608;
  assign n10610 = ~n10597 & ~n10609;
  assign n10611 = ~controllable_hgrant2 & ~n10610;
  assign n10612 = ~n10111 & ~n10611;
  assign n10613 = controllable_hmaster1 & ~n10612;
  assign n10614 = controllable_hmaster0 & ~n10612;
  assign n10615 = ~n10462 & ~n10599;
  assign n10616 = ~i_hbusreq0 & ~n10615;
  assign n10617 = ~n10453 & ~n10616;
  assign n10618 = ~i_hbusreq4 & ~n10617;
  assign n10619 = ~n10452 & ~n10618;
  assign n10620 = ~controllable_hgrant4 & n10619;
  assign n10621 = ~n4667 & ~n10620;
  assign n10622 = ~i_hbusreq2 & ~n10621;
  assign n10623 = ~n10451 & ~n10622;
  assign n10624 = ~controllable_hgrant2 & ~n10623;
  assign n10625 = ~n10111 & ~n10624;
  assign n10626 = ~controllable_hmaster0 & ~n10625;
  assign n10627 = ~n10614 & ~n10626;
  assign n10628 = ~controllable_hmaster1 & ~n10627;
  assign n10629 = ~n10613 & ~n10628;
  assign n10630 = ~i_hbusreq3 & ~n10629;
  assign n10631 = ~n10596 & ~n10630;
  assign n10632 = controllable_hmaster2 & ~n10631;
  assign n10633 = ~n5686 & ~n10589;
  assign n10634 = ~controllable_hmaster0 & ~n10633;
  assign n10635 = ~n10592 & ~n10634;
  assign n10636 = controllable_hmaster1 & ~n10635;
  assign n10637 = i_hready & ~n10496;
  assign n10638 = ~controllable_hgrant4 & n10637;
  assign n10639 = ~n4091 & ~n10638;
  assign n10640 = ~controllable_hgrant2 & ~n10639;
  assign n10641 = ~n5616 & ~n10640;
  assign n10642 = controllable_hmaster0 & ~n10641;
  assign n10643 = ~controllable_hmaster0 & ~n10590;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = ~controllable_hmaster1 & ~n10644;
  assign n10646 = ~n10636 & ~n10645;
  assign n10647 = i_hbusreq3 & ~n10646;
  assign n10648 = ~n10112 & ~n10620;
  assign n10649 = ~i_hbusreq2 & ~n10648;
  assign n10650 = ~n10597 & ~n10649;
  assign n10651 = ~controllable_hgrant2 & ~n10650;
  assign n10652 = ~n10111 & ~n10651;
  assign n10653 = controllable_hmaster0 & ~n10652;
  assign n10654 = ~n10152 & ~n10651;
  assign n10655 = ~controllable_hmaster0 & ~n10654;
  assign n10656 = ~n10653 & ~n10655;
  assign n10657 = controllable_hmaster1 & ~n10656;
  assign n10658 = i_hbusreq2 & ~n10639;
  assign n10659 = i_hbusreq4 & ~n10637;
  assign n10660 = i_hbusreq0 & ~n10637;
  assign n10661 = ~n10157 & ~n10535;
  assign n10662 = ~controllable_ndecide & ~n10661;
  assign n10663 = ~controllable_ndecide & ~n10662;
  assign n10664 = i_hready & ~n10663;
  assign n10665 = ~n10361 & ~n10664;
  assign n10666 = i_hlock0 & ~n10665;
  assign n10667 = i_hready & ~n10544;
  assign n10668 = ~i_hlock0 & ~n10667;
  assign n10669 = ~n10666 & ~n10668;
  assign n10670 = ~i_hbusreq0 & ~n10669;
  assign n10671 = ~n10660 & ~n10670;
  assign n10672 = ~i_hbusreq4 & ~n10671;
  assign n10673 = ~n10659 & ~n10672;
  assign n10674 = ~controllable_hgrant4 & n10673;
  assign n10675 = ~n10112 & ~n10674;
  assign n10676 = ~i_hbusreq2 & ~n10675;
  assign n10677 = ~n10658 & ~n10676;
  assign n10678 = ~controllable_hgrant2 & ~n10677;
  assign n10679 = ~n10111 & ~n10678;
  assign n10680 = controllable_hmaster0 & ~n10679;
  assign n10681 = ~i_hbusreq0 & ~n10461;
  assign n10682 = ~n10453 & ~n10681;
  assign n10683 = ~i_hbusreq4 & ~n10682;
  assign n10684 = ~n10452 & ~n10683;
  assign n10685 = ~controllable_hgrant4 & n10684;
  assign n10686 = ~n4091 & ~n10685;
  assign n10687 = ~i_hbusreq2 & ~n10686;
  assign n10688 = ~n10597 & ~n10687;
  assign n10689 = ~controllable_hgrant2 & ~n10688;
  assign n10690 = ~n5616 & ~n10689;
  assign n10691 = ~controllable_hmaster0 & ~n10690;
  assign n10692 = ~n10680 & ~n10691;
  assign n10693 = ~controllable_hmaster1 & ~n10692;
  assign n10694 = ~n10657 & ~n10693;
  assign n10695 = ~i_hbusreq3 & ~n10694;
  assign n10696 = ~n10647 & ~n10695;
  assign n10697 = ~controllable_hmaster2 & ~n10696;
  assign n10698 = ~n10632 & ~n10697;
  assign n10699 = ~controllable_hgrant3 & ~n10698;
  assign n10700 = ~n10110 & ~n10699;
  assign n10701 = controllable_nhgrant0 & ~n10700;
  assign n10702 = ~n10240 & ~n10701;
  assign n10703 = ~n3281 & ~n10702;
  assign n10704 = ~n3281 & ~n10703;
  assign n10705 = ~n3378 & ~n10704;
  assign n10706 = ~n10587 & ~n10705;
  assign n10707 = n3492 & ~n10706;
  assign n10708 = ~n8563 & ~n10707;
  assign n10709 = n3485 & ~n10708;
  assign n10710 = ~n8705 & ~n10709;
  assign n10711 = n3476 & ~n10710;
  assign n10712 = ~n10396 & ~n10711;
  assign n10713 = n3374 & ~n10712;
  assign n10714 = ~n10311 & ~n10713;
  assign n10715 = ~n3655 & ~n10714;
  assign n10716 = ~n10254 & ~n10715;
  assign n10717 = n3652 & ~n10716;
  assign n10718 = n3378 & ~n7979;
  assign n10719 = ~n3499 & ~n4787;
  assign n10720 = controllable_hmaster1 & ~n10719;
  assign n10721 = controllable_hmaster0 & ~n10719;
  assign n10722 = controllable_hmaster0 & ~n10721;
  assign n10723 = ~controllable_hmaster1 & ~n10722;
  assign n10724 = ~n10720 & ~n10723;
  assign n10725 = i_hbusreq3 & ~n10724;
  assign n10726 = ~n4794 & ~n9722;
  assign n10727 = controllable_hmaster1 & ~n10726;
  assign n10728 = controllable_hmaster0 & ~n10726;
  assign n10729 = controllable_hmaster0 & ~n10728;
  assign n10730 = ~controllable_hmaster1 & ~n10729;
  assign n10731 = ~n10727 & ~n10730;
  assign n10732 = ~i_hbusreq3 & ~n10731;
  assign n10733 = ~n10725 & ~n10732;
  assign n10734 = controllable_hmaster2 & ~n10733;
  assign n10735 = controllable_hmaster2 & ~n10734;
  assign n10736 = ~controllable_hgrant3 & ~n10735;
  assign n10737 = ~n9708 & ~n10736;
  assign n10738 = controllable_nhgrant0 & ~n10737;
  assign n10739 = ~n9753 & ~n10738;
  assign n10740 = ~n3281 & ~n10739;
  assign n10741 = ~n3281 & ~n10740;
  assign n10742 = ~n3378 & ~n10741;
  assign n10743 = ~n10718 & ~n10742;
  assign n10744 = n3492 & ~n10743;
  assign n10745 = n3492 & ~n10744;
  assign n10746 = n3485 & ~n10745;
  assign n10747 = n3485 & ~n10746;
  assign n10748 = ~n3476 & ~n10747;
  assign n10749 = ~n8523 & ~n10744;
  assign n10750 = n3485 & ~n10749;
  assign n10751 = ~n8689 & ~n10750;
  assign n10752 = n3476 & ~n10751;
  assign n10753 = ~n10748 & ~n10752;
  assign n10754 = ~n3374 & ~n10753;
  assign n10755 = n3378 & ~n8021;
  assign n10756 = ~n4789 & ~n10721;
  assign n10757 = ~controllable_hmaster1 & ~n10756;
  assign n10758 = ~n10720 & ~n10757;
  assign n10759 = i_hbusreq3 & ~n10758;
  assign n10760 = ~n4796 & ~n10728;
  assign n10761 = ~controllable_hmaster1 & ~n10760;
  assign n10762 = ~n10727 & ~n10761;
  assign n10763 = ~i_hbusreq3 & ~n10762;
  assign n10764 = ~n10759 & ~n10763;
  assign n10765 = controllable_hmaster2 & ~n10764;
  assign n10766 = ~n4787 & ~n8768;
  assign n10767 = controllable_hmaster0 & ~n10766;
  assign n10768 = controllable_hgrant2 & ~n3498;
  assign n10769 = ~n8768 & ~n10768;
  assign n10770 = ~controllable_hmaster0 & ~n10769;
  assign n10771 = ~n10767 & ~n10770;
  assign n10772 = controllable_hmaster1 & ~n10771;
  assign n10773 = ~n4787 & ~n8824;
  assign n10774 = controllable_hmaster0 & ~n10773;
  assign n10775 = ~controllable_hmaster0 & ~n10766;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = ~controllable_hmaster1 & ~n10776;
  assign n10778 = ~n10772 & ~n10777;
  assign n10779 = i_hbusreq3 & ~n10778;
  assign n10780 = ~n4794 & ~n9800;
  assign n10781 = controllable_hmaster0 & ~n10780;
  assign n10782 = controllable_hgrant2 & ~n9721;
  assign n10783 = ~n9800 & ~n10782;
  assign n10784 = ~controllable_hmaster0 & ~n10783;
  assign n10785 = ~n10781 & ~n10784;
  assign n10786 = controllable_hmaster1 & ~n10785;
  assign n10787 = ~n4794 & ~n9824;
  assign n10788 = controllable_hmaster0 & ~n10787;
  assign n10789 = ~n10775 & ~n10788;
  assign n10790 = ~controllable_hmaster1 & ~n10789;
  assign n10791 = ~n10786 & ~n10790;
  assign n10792 = ~i_hbusreq3 & ~n10791;
  assign n10793 = ~n10779 & ~n10792;
  assign n10794 = ~controllable_hmaster2 & ~n10793;
  assign n10795 = ~n10765 & ~n10794;
  assign n10796 = ~controllable_hgrant3 & ~n10795;
  assign n10797 = ~n9790 & ~n10796;
  assign n10798 = controllable_nhgrant0 & ~n10797;
  assign n10799 = ~n9861 & ~n10798;
  assign n10800 = ~n3281 & ~n10799;
  assign n10801 = ~n3281 & ~n10800;
  assign n10802 = ~n3378 & ~n10801;
  assign n10803 = ~n10755 & ~n10802;
  assign n10804 = n3492 & ~n10803;
  assign n10805 = n3492 & ~n10804;
  assign n10806 = n3485 & ~n10805;
  assign n10807 = n3485 & ~n10806;
  assign n10808 = ~n3476 & ~n10807;
  assign n10809 = ~controllable_hgrant4 & ~n9955;
  assign n10810 = ~n3411 & ~n10809;
  assign n10811 = i_hlock2 & ~n10810;
  assign n10812 = ~controllable_hgrant4 & ~n9959;
  assign n10813 = ~n3411 & ~n10812;
  assign n10814 = ~i_hlock2 & ~n10813;
  assign n10815 = ~n10811 & ~n10814;
  assign n10816 = controllable_hgrant2 & ~n10815;
  assign n10817 = ~n9875 & ~n10816;
  assign n10818 = controllable_hmaster1 & ~n10817;
  assign n10819 = controllable_hmaster0 & ~n10817;
  assign n10820 = ~controllable_hgrant4 & ~n9968;
  assign n10821 = ~n3411 & ~n10820;
  assign n10822 = i_hlock2 & ~n10821;
  assign n10823 = ~controllable_hgrant4 & ~n9970;
  assign n10824 = ~n3411 & ~n10823;
  assign n10825 = ~i_hlock2 & ~n10824;
  assign n10826 = ~n10822 & ~n10825;
  assign n10827 = controllable_hgrant2 & ~n10826;
  assign n10828 = ~n5628 & ~n10827;
  assign n10829 = ~controllable_hmaster0 & ~n10828;
  assign n10830 = ~n10819 & ~n10829;
  assign n10831 = ~controllable_hmaster1 & ~n10830;
  assign n10832 = ~n10818 & ~n10831;
  assign n10833 = i_hbusreq3 & ~n10832;
  assign n10834 = i_hbusreq2 & ~n10815;
  assign n10835 = i_hbusreq4 & ~n9955;
  assign n10836 = i_hbusreq0 & ~n9955;
  assign n10837 = ~n3568 & ~n3920;
  assign n10838 = i_hlock0 & ~n10837;
  assign n10839 = ~n3564 & ~n4655;
  assign n10840 = ~controllable_ndecide & ~n10839;
  assign n10841 = ~n3494 & ~n10840;
  assign n10842 = i_hready & ~n10841;
  assign n10843 = ~n3904 & ~n10842;
  assign n10844 = ~i_hlock0 & ~n10843;
  assign n10845 = ~n10838 & ~n10844;
  assign n10846 = ~i_hbusreq0 & ~n10845;
  assign n10847 = ~n10836 & ~n10846;
  assign n10848 = ~i_hbusreq4 & ~n10847;
  assign n10849 = ~n10835 & ~n10848;
  assign n10850 = ~controllable_hgrant4 & ~n10849;
  assign n10851 = ~n3916 & ~n10850;
  assign n10852 = i_hlock2 & ~n10851;
  assign n10853 = i_hbusreq4 & ~n9959;
  assign n10854 = i_hbusreq0 & ~n9959;
  assign n10855 = ~n3494 & ~n4029;
  assign n10856 = i_hready & ~n10855;
  assign n10857 = ~n3920 & ~n10856;
  assign n10858 = i_hlock0 & ~n10857;
  assign n10859 = ~n9960 & ~n10858;
  assign n10860 = ~i_hbusreq0 & ~n10859;
  assign n10861 = ~n10854 & ~n10860;
  assign n10862 = ~i_hbusreq4 & ~n10861;
  assign n10863 = ~n10853 & ~n10862;
  assign n10864 = ~controllable_hgrant4 & ~n10863;
  assign n10865 = ~n3916 & ~n10864;
  assign n10866 = ~i_hlock2 & ~n10865;
  assign n10867 = ~n10852 & ~n10866;
  assign n10868 = ~i_hbusreq2 & ~n10867;
  assign n10869 = ~n10834 & ~n10868;
  assign n10870 = controllable_hgrant2 & ~n10869;
  assign n10871 = ~n9899 & ~n10870;
  assign n10872 = controllable_hmaster1 & ~n10871;
  assign n10873 = controllable_hmaster0 & ~n10871;
  assign n10874 = i_hbusreq2 & ~n10826;
  assign n10875 = i_hbusreq4 & ~n9968;
  assign n10876 = i_hbusreq0 & ~n9968;
  assign n10877 = ~n3568 & ~n4621;
  assign n10878 = i_hlock0 & ~n10877;
  assign n10879 = ~n4605 & ~n10842;
  assign n10880 = ~i_hlock0 & ~n10879;
  assign n10881 = ~n10878 & ~n10880;
  assign n10882 = ~i_hbusreq0 & ~n10881;
  assign n10883 = ~n10876 & ~n10882;
  assign n10884 = ~i_hbusreq4 & ~n10883;
  assign n10885 = ~n10875 & ~n10884;
  assign n10886 = ~controllable_hgrant4 & ~n10885;
  assign n10887 = ~n4617 & ~n10886;
  assign n10888 = i_hlock2 & ~n10887;
  assign n10889 = i_hbusreq4 & ~n9970;
  assign n10890 = i_hbusreq0 & ~n9970;
  assign n10891 = ~n4621 & ~n10856;
  assign n10892 = i_hlock0 & ~n10891;
  assign n10893 = ~n9971 & ~n10892;
  assign n10894 = ~i_hbusreq0 & ~n10893;
  assign n10895 = ~n10890 & ~n10894;
  assign n10896 = ~i_hbusreq4 & ~n10895;
  assign n10897 = ~n10889 & ~n10896;
  assign n10898 = ~controllable_hgrant4 & ~n10897;
  assign n10899 = ~n4617 & ~n10898;
  assign n10900 = ~i_hlock2 & ~n10899;
  assign n10901 = ~n10888 & ~n10900;
  assign n10902 = ~i_hbusreq2 & ~n10901;
  assign n10903 = ~n10874 & ~n10902;
  assign n10904 = controllable_hgrant2 & ~n10903;
  assign n10905 = ~n9914 & ~n10904;
  assign n10906 = ~controllable_hmaster0 & ~n10905;
  assign n10907 = ~n10873 & ~n10906;
  assign n10908 = ~controllable_hmaster1 & ~n10907;
  assign n10909 = ~n10872 & ~n10908;
  assign n10910 = ~i_hbusreq3 & ~n10909;
  assign n10911 = ~n10833 & ~n10910;
  assign n10912 = controllable_hmaster2 & ~n10911;
  assign n10913 = ~n5913 & ~n10816;
  assign n10914 = controllable_hmaster0 & ~n10913;
  assign n10915 = ~controllable_hgrant4 & ~n10029;
  assign n10916 = ~n3411 & ~n10915;
  assign n10917 = i_hlock2 & ~n10916;
  assign n10918 = ~controllable_hgrant4 & ~n10033;
  assign n10919 = ~n3411 & ~n10918;
  assign n10920 = ~i_hlock2 & ~n10919;
  assign n10921 = ~n10917 & ~n10920;
  assign n10922 = controllable_hgrant2 & ~n10921;
  assign n10923 = ~n5913 & ~n10922;
  assign n10924 = ~controllable_hmaster0 & ~n10923;
  assign n10925 = ~n10914 & ~n10924;
  assign n10926 = controllable_hmaster1 & ~n10925;
  assign n10927 = ~n5923 & ~n10816;
  assign n10928 = controllable_hmaster0 & ~n10927;
  assign n10929 = ~controllable_hmaster0 & ~n10913;
  assign n10930 = ~n10928 & ~n10929;
  assign n10931 = ~controllable_hmaster1 & ~n10930;
  assign n10932 = ~n10926 & ~n10931;
  assign n10933 = i_hbusreq3 & ~n10932;
  assign n10934 = ~n9926 & ~n10870;
  assign n10935 = controllable_hmaster0 & ~n10934;
  assign n10936 = i_hbusreq2 & ~n10921;
  assign n10937 = i_hbusreq4 & ~n10029;
  assign n10938 = i_hbusreq0 & ~n10029;
  assign n10939 = ~n3568 & ~n5055;
  assign n10940 = i_hlock0 & ~n10939;
  assign n10941 = ~n3564 & ~n8938;
  assign n10942 = ~controllable_ndecide & ~n10941;
  assign n10943 = ~n3494 & ~n10942;
  assign n10944 = i_hready & ~n10943;
  assign n10945 = ~n5039 & ~n10944;
  assign n10946 = ~i_hlock0 & ~n10945;
  assign n10947 = ~n10940 & ~n10946;
  assign n10948 = ~i_hbusreq0 & ~n10947;
  assign n10949 = ~n10938 & ~n10948;
  assign n10950 = ~i_hbusreq4 & ~n10949;
  assign n10951 = ~n10937 & ~n10950;
  assign n10952 = ~controllable_hgrant4 & ~n10951;
  assign n10953 = ~n3916 & ~n10952;
  assign n10954 = i_hlock2 & ~n10953;
  assign n10955 = i_hbusreq4 & ~n10033;
  assign n10956 = i_hbusreq0 & ~n10033;
  assign n10957 = ~n3494 & ~n4053;
  assign n10958 = i_hready & ~n10957;
  assign n10959 = ~n5055 & ~n10958;
  assign n10960 = i_hlock0 & ~n10959;
  assign n10961 = ~n10034 & ~n10960;
  assign n10962 = ~i_hbusreq0 & ~n10961;
  assign n10963 = ~n10956 & ~n10962;
  assign n10964 = ~i_hbusreq4 & ~n10963;
  assign n10965 = ~n10955 & ~n10964;
  assign n10966 = ~controllable_hgrant4 & ~n10965;
  assign n10967 = ~n3916 & ~n10966;
  assign n10968 = ~i_hlock2 & ~n10967;
  assign n10969 = ~n10954 & ~n10968;
  assign n10970 = ~i_hbusreq2 & ~n10969;
  assign n10971 = ~n10936 & ~n10970;
  assign n10972 = controllable_hgrant2 & ~n10971;
  assign n10973 = ~n9926 & ~n10972;
  assign n10974 = ~controllable_hmaster0 & ~n10973;
  assign n10975 = ~n10935 & ~n10974;
  assign n10976 = controllable_hmaster1 & ~n10975;
  assign n10977 = ~n9936 & ~n10870;
  assign n10978 = controllable_hmaster0 & ~n10977;
  assign n10979 = ~n3568 & ~n5464;
  assign n10980 = i_hlock0 & ~n10979;
  assign n10981 = ~n10844 & ~n10980;
  assign n10982 = ~i_hbusreq0 & ~n10981;
  assign n10983 = ~n10836 & ~n10982;
  assign n10984 = ~i_hbusreq4 & ~n10983;
  assign n10985 = ~n10835 & ~n10984;
  assign n10986 = ~controllable_hgrant4 & ~n10985;
  assign n10987 = ~n5462 & ~n10986;
  assign n10988 = i_hlock2 & ~n10987;
  assign n10989 = ~n5464 & ~n10856;
  assign n10990 = i_hlock0 & ~n10989;
  assign n10991 = ~n9960 & ~n10990;
  assign n10992 = ~i_hbusreq0 & ~n10991;
  assign n10993 = ~n10854 & ~n10992;
  assign n10994 = ~i_hbusreq4 & ~n10993;
  assign n10995 = ~n10853 & ~n10994;
  assign n10996 = ~controllable_hgrant4 & ~n10995;
  assign n10997 = ~n5462 & ~n10996;
  assign n10998 = ~i_hlock2 & ~n10997;
  assign n10999 = ~n10988 & ~n10998;
  assign n11000 = ~i_hbusreq2 & ~n10999;
  assign n11001 = ~n10834 & ~n11000;
  assign n11002 = controllable_hgrant2 & ~n11001;
  assign n11003 = ~n9942 & ~n11002;
  assign n11004 = ~controllable_hmaster0 & ~n11003;
  assign n11005 = ~n10978 & ~n11004;
  assign n11006 = ~controllable_hmaster1 & ~n11005;
  assign n11007 = ~n10976 & ~n11006;
  assign n11008 = ~i_hbusreq3 & ~n11007;
  assign n11009 = ~n10933 & ~n11008;
  assign n11010 = ~controllable_hmaster2 & ~n11009;
  assign n11011 = ~n10912 & ~n11010;
  assign n11012 = ~controllable_hgrant3 & ~n11011;
  assign n11013 = ~n7457 & ~n11012;
  assign n11014 = controllable_nhgrant0 & ~n11013;
  assign n11015 = ~n10071 & ~n11014;
  assign n11016 = ~n3281 & ~n11015;
  assign n11017 = ~n3281 & ~n11016;
  assign n11018 = n3378 & ~n11017;
  assign n11019 = ~n5623 & ~n10827;
  assign n11020 = controllable_hmaster1 & ~n11019;
  assign n11021 = controllable_hmaster0 & ~n11019;
  assign n11022 = ~n10829 & ~n11021;
  assign n11023 = ~controllable_hmaster1 & ~n11022;
  assign n11024 = ~n11020 & ~n11023;
  assign n11025 = i_hbusreq3 & ~n11024;
  assign n11026 = ~n4621 & ~n10842;
  assign n11027 = i_hlock0 & ~n11026;
  assign n11028 = ~n10880 & ~n11027;
  assign n11029 = ~i_hbusreq0 & ~n11028;
  assign n11030 = ~n10876 & ~n11029;
  assign n11031 = ~i_hbusreq4 & ~n11030;
  assign n11032 = ~n10875 & ~n11031;
  assign n11033 = ~controllable_hgrant4 & ~n11032;
  assign n11034 = ~n4617 & ~n11033;
  assign n11035 = i_hlock2 & ~n11034;
  assign n11036 = ~n4621 & ~n9958;
  assign n11037 = i_hlock0 & ~n11036;
  assign n11038 = ~n9971 & ~n11037;
  assign n11039 = ~i_hbusreq0 & ~n11038;
  assign n11040 = ~n10890 & ~n11039;
  assign n11041 = ~i_hbusreq4 & ~n11040;
  assign n11042 = ~n10889 & ~n11041;
  assign n11043 = ~controllable_hgrant4 & ~n11042;
  assign n11044 = ~n4617 & ~n11043;
  assign n11045 = ~i_hlock2 & ~n11044;
  assign n11046 = ~n11035 & ~n11045;
  assign n11047 = ~i_hbusreq2 & ~n11046;
  assign n11048 = ~n10874 & ~n11047;
  assign n11049 = controllable_hgrant2 & ~n11048;
  assign n11050 = ~n10124 & ~n11049;
  assign n11051 = controllable_hmaster1 & ~n11050;
  assign n11052 = controllable_hmaster0 & ~n11050;
  assign n11053 = ~n10137 & ~n11049;
  assign n11054 = ~controllable_hmaster0 & ~n11053;
  assign n11055 = ~n11052 & ~n11054;
  assign n11056 = ~controllable_hmaster1 & ~n11055;
  assign n11057 = ~n11051 & ~n11056;
  assign n11058 = ~i_hbusreq3 & ~n11057;
  assign n11059 = ~n11025 & ~n11058;
  assign n11060 = controllable_hmaster2 & ~n11059;
  assign n11061 = i_hlock2 & ~n3546;
  assign n11062 = ~controllable_hgrant4 & ~n10217;
  assign n11063 = ~n3411 & ~n11062;
  assign n11064 = ~i_hlock2 & ~n11063;
  assign n11065 = ~n11061 & ~n11064;
  assign n11066 = controllable_hgrant2 & ~n11065;
  assign n11067 = ~n5623 & ~n11066;
  assign n11068 = ~controllable_hmaster0 & ~n11067;
  assign n11069 = ~n11021 & ~n11068;
  assign n11070 = controllable_hmaster1 & ~n11069;
  assign n11071 = ~n8989 & ~n10827;
  assign n11072 = controllable_hmaster0 & ~n11071;
  assign n11073 = ~controllable_hmaster0 & ~n11019;
  assign n11074 = ~n11072 & ~n11073;
  assign n11075 = ~controllable_hmaster1 & ~n11074;
  assign n11076 = ~n11070 & ~n11075;
  assign n11077 = i_hbusreq3 & ~n11076;
  assign n11078 = ~n10149 & ~n11049;
  assign n11079 = controllable_hmaster0 & ~n11078;
  assign n11080 = i_hbusreq2 & ~n11065;
  assign n11081 = ~n4577 & ~n10842;
  assign n11082 = i_hlock0 & ~n11081;
  assign n11083 = ~n3495 & ~n10944;
  assign n11084 = ~i_hlock0 & ~n11083;
  assign n11085 = ~n11082 & ~n11084;
  assign n11086 = ~i_hbusreq0 & ~n11085;
  assign n11087 = ~n3563 & ~n11086;
  assign n11088 = ~i_hbusreq4 & ~n11087;
  assign n11089 = ~n3562 & ~n11088;
  assign n11090 = ~controllable_hgrant4 & ~n11089;
  assign n11091 = ~n4617 & ~n11090;
  assign n11092 = i_hlock2 & ~n11091;
  assign n11093 = i_hbusreq4 & ~n10217;
  assign n11094 = i_hbusreq0 & ~n10217;
  assign n11095 = ~n3494 & ~n4657;
  assign n11096 = i_hready & ~n11095;
  assign n11097 = ~n4577 & ~n11096;
  assign n11098 = i_hlock0 & ~n11097;
  assign n11099 = ~n10218 & ~n11098;
  assign n11100 = ~i_hbusreq0 & ~n11099;
  assign n11101 = ~n11094 & ~n11100;
  assign n11102 = ~i_hbusreq4 & ~n11101;
  assign n11103 = ~n11093 & ~n11102;
  assign n11104 = ~controllable_hgrant4 & ~n11103;
  assign n11105 = ~n4617 & ~n11104;
  assign n11106 = ~i_hlock2 & ~n11105;
  assign n11107 = ~n11092 & ~n11106;
  assign n11108 = ~i_hbusreq2 & ~n11107;
  assign n11109 = ~n11080 & ~n11108;
  assign n11110 = controllable_hgrant2 & ~n11109;
  assign n11111 = ~n10149 & ~n11110;
  assign n11112 = ~controllable_hmaster0 & ~n11111;
  assign n11113 = ~n11079 & ~n11112;
  assign n11114 = controllable_hmaster1 & ~n11113;
  assign n11115 = ~n10173 & ~n11049;
  assign n11116 = controllable_hmaster0 & ~n11115;
  assign n11117 = ~i_hbusreq0 & ~n10879;
  assign n11118 = ~n10876 & ~n11117;
  assign n11119 = ~i_hbusreq4 & ~n11118;
  assign n11120 = ~n10875 & ~n11119;
  assign n11121 = ~controllable_hgrant4 & ~n11120;
  assign n11122 = ~n3411 & ~n11121;
  assign n11123 = i_hlock2 & ~n11122;
  assign n11124 = ~n10825 & ~n11123;
  assign n11125 = ~i_hbusreq2 & ~n11124;
  assign n11126 = ~n10874 & ~n11125;
  assign n11127 = controllable_hgrant2 & ~n11126;
  assign n11128 = ~n10184 & ~n11127;
  assign n11129 = ~controllable_hmaster0 & ~n11128;
  assign n11130 = ~n11116 & ~n11129;
  assign n11131 = ~controllable_hmaster1 & ~n11130;
  assign n11132 = ~n11114 & ~n11131;
  assign n11133 = ~i_hbusreq3 & ~n11132;
  assign n11134 = ~n11077 & ~n11133;
  assign n11135 = ~controllable_hmaster2 & ~n11134;
  assign n11136 = ~n11060 & ~n11135;
  assign n11137 = ~controllable_hgrant3 & ~n11136;
  assign n11138 = ~n10110 & ~n11137;
  assign n11139 = controllable_nhgrant0 & ~n11138;
  assign n11140 = ~n10240 & ~n11139;
  assign n11141 = ~n3281 & ~n11140;
  assign n11142 = ~n3281 & ~n11141;
  assign n11143 = ~n3378 & ~n11142;
  assign n11144 = ~n11018 & ~n11143;
  assign n11145 = n3492 & ~n11144;
  assign n11146 = ~n8592 & ~n11145;
  assign n11147 = n3485 & ~n11146;
  assign n11148 = ~n8718 & ~n11147;
  assign n11149 = n3476 & ~n11148;
  assign n11150 = ~n10808 & ~n11149;
  assign n11151 = n3374 & ~n11150;
  assign n11152 = ~n10754 & ~n11151;
  assign n11153 = n3655 & ~n11152;
  assign n11154 = n3378 & ~n8138;
  assign n11155 = ~n4787 & ~n10259;
  assign n11156 = controllable_hmaster1 & ~n11155;
  assign n11157 = controllable_hmaster0 & ~n11155;
  assign n11158 = controllable_hmaster0 & ~n11157;
  assign n11159 = ~controllable_hmaster1 & ~n11158;
  assign n11160 = ~n11156 & ~n11159;
  assign n11161 = i_hbusreq3 & ~n11160;
  assign n11162 = ~n4794 & ~n10282;
  assign n11163 = controllable_hmaster1 & ~n11162;
  assign n11164 = controllable_hmaster0 & ~n11162;
  assign n11165 = controllable_hmaster0 & ~n11164;
  assign n11166 = ~controllable_hmaster1 & ~n11165;
  assign n11167 = ~n11163 & ~n11166;
  assign n11168 = ~i_hbusreq3 & ~n11167;
  assign n11169 = ~n11161 & ~n11168;
  assign n11170 = controllable_hmaster2 & ~n11169;
  assign n11171 = controllable_hmaster2 & ~n11170;
  assign n11172 = ~controllable_hgrant3 & ~n11171;
  assign n11173 = ~n9708 & ~n11172;
  assign n11174 = controllable_nhgrant0 & ~n11173;
  assign n11175 = ~n9753 & ~n11174;
  assign n11176 = ~n3281 & ~n11175;
  assign n11177 = ~n3281 & ~n11176;
  assign n11178 = ~n3378 & ~n11177;
  assign n11179 = ~n11154 & ~n11178;
  assign n11180 = n3492 & ~n11179;
  assign n11181 = n3492 & ~n11180;
  assign n11182 = n3485 & ~n11181;
  assign n11183 = n3485 & ~n11182;
  assign n11184 = ~n3476 & ~n11183;
  assign n11185 = ~n8523 & ~n11180;
  assign n11186 = n3485 & ~n11185;
  assign n11187 = ~n8689 & ~n11186;
  assign n11188 = n3476 & ~n11187;
  assign n11189 = ~n11184 & ~n11188;
  assign n11190 = ~n3374 & ~n11189;
  assign n11191 = n3378 & ~n8180;
  assign n11192 = ~n4846 & ~n11157;
  assign n11193 = ~controllable_hmaster1 & ~n11192;
  assign n11194 = ~n11156 & ~n11193;
  assign n11195 = i_hbusreq3 & ~n11194;
  assign n11196 = ~n4852 & ~n11164;
  assign n11197 = ~controllable_hmaster1 & ~n11196;
  assign n11198 = ~n11163 & ~n11197;
  assign n11199 = ~i_hbusreq3 & ~n11198;
  assign n11200 = ~n11195 & ~n11199;
  assign n11201 = controllable_hmaster2 & ~n11200;
  assign n11202 = ~n4787 & ~n10324;
  assign n11203 = controllable_hmaster0 & ~n11202;
  assign n11204 = ~n10324 & ~n10768;
  assign n11205 = ~controllable_hmaster0 & ~n11204;
  assign n11206 = ~n11203 & ~n11205;
  assign n11207 = controllable_hmaster1 & ~n11206;
  assign n11208 = ~n4787 & ~n10334;
  assign n11209 = controllable_hmaster0 & ~n11208;
  assign n11210 = ~controllable_hmaster0 & ~n11202;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = ~controllable_hmaster1 & ~n11211;
  assign n11213 = ~n11207 & ~n11212;
  assign n11214 = i_hbusreq3 & ~n11213;
  assign n11215 = ~n4794 & ~n10346;
  assign n11216 = controllable_hmaster0 & ~n11215;
  assign n11217 = ~n10346 & ~n10782;
  assign n11218 = ~controllable_hmaster0 & ~n11217;
  assign n11219 = ~n11216 & ~n11218;
  assign n11220 = controllable_hmaster1 & ~n11219;
  assign n11221 = ~n4794 & ~n10374;
  assign n11222 = controllable_hmaster0 & ~n11221;
  assign n11223 = ~n11210 & ~n11222;
  assign n11224 = ~controllable_hmaster1 & ~n11223;
  assign n11225 = ~n11220 & ~n11224;
  assign n11226 = ~i_hbusreq3 & ~n11225;
  assign n11227 = ~n11214 & ~n11226;
  assign n11228 = ~controllable_hmaster2 & ~n11227;
  assign n11229 = ~n11201 & ~n11228;
  assign n11230 = ~controllable_hgrant3 & ~n11229;
  assign n11231 = ~n9790 & ~n11230;
  assign n11232 = controllable_nhgrant0 & ~n11231;
  assign n11233 = ~n9861 & ~n11232;
  assign n11234 = ~n3281 & ~n11233;
  assign n11235 = ~n3281 & ~n11234;
  assign n11236 = ~n3378 & ~n11235;
  assign n11237 = ~n11191 & ~n11236;
  assign n11238 = n3492 & ~n11237;
  assign n11239 = n3492 & ~n11238;
  assign n11240 = n3485 & ~n11239;
  assign n11241 = n3485 & ~n11240;
  assign n11242 = ~n3476 & ~n11241;
  assign n11243 = ~n10406 & ~n10816;
  assign n11244 = controllable_hmaster1 & ~n11243;
  assign n11245 = controllable_hmaster0 & ~n11243;
  assign n11246 = ~n10414 & ~n10827;
  assign n11247 = ~controllable_hmaster0 & ~n11246;
  assign n11248 = ~n11245 & ~n11247;
  assign n11249 = ~controllable_hmaster1 & ~n11248;
  assign n11250 = ~n11244 & ~n11249;
  assign n11251 = i_hbusreq3 & ~n11250;
  assign n11252 = ~n10447 & ~n10870;
  assign n11253 = controllable_hmaster1 & ~n11252;
  assign n11254 = controllable_hmaster0 & ~n11252;
  assign n11255 = ~n10472 & ~n10904;
  assign n11256 = ~controllable_hmaster0 & ~n11255;
  assign n11257 = ~n11254 & ~n11256;
  assign n11258 = ~controllable_hmaster1 & ~n11257;
  assign n11259 = ~n11253 & ~n11258;
  assign n11260 = ~i_hbusreq3 & ~n11259;
  assign n11261 = ~n11251 & ~n11260;
  assign n11262 = controllable_hmaster2 & ~n11261;
  assign n11263 = ~n10485 & ~n10816;
  assign n11264 = controllable_hmaster0 & ~n11263;
  assign n11265 = ~n10485 & ~n10922;
  assign n11266 = ~controllable_hmaster0 & ~n11265;
  assign n11267 = ~n11264 & ~n11266;
  assign n11268 = controllable_hmaster1 & ~n11267;
  assign n11269 = ~n10500 & ~n10816;
  assign n11270 = controllable_hmaster0 & ~n11269;
  assign n11271 = ~controllable_hmaster0 & ~n11263;
  assign n11272 = ~n11270 & ~n11271;
  assign n11273 = ~controllable_hmaster1 & ~n11272;
  assign n11274 = ~n11268 & ~n11273;
  assign n11275 = i_hbusreq3 & ~n11274;
  assign n11276 = ~n10525 & ~n10870;
  assign n11277 = controllable_hmaster0 & ~n11276;
  assign n11278 = ~n10525 & ~n10972;
  assign n11279 = ~controllable_hmaster0 & ~n11278;
  assign n11280 = ~n11277 & ~n11279;
  assign n11281 = controllable_hmaster1 & ~n11280;
  assign n11282 = ~n10556 & ~n10870;
  assign n11283 = controllable_hmaster0 & ~n11282;
  assign n11284 = ~n10571 & ~n11002;
  assign n11285 = ~controllable_hmaster0 & ~n11284;
  assign n11286 = ~n11283 & ~n11285;
  assign n11287 = ~controllable_hmaster1 & ~n11286;
  assign n11288 = ~n11281 & ~n11287;
  assign n11289 = ~i_hbusreq3 & ~n11288;
  assign n11290 = ~n11275 & ~n11289;
  assign n11291 = ~controllable_hmaster2 & ~n11290;
  assign n11292 = ~n11262 & ~n11291;
  assign n11293 = ~controllable_hgrant3 & ~n11292;
  assign n11294 = ~n7457 & ~n11293;
  assign n11295 = controllable_nhgrant0 & ~n11294;
  assign n11296 = ~n10071 & ~n11295;
  assign n11297 = ~n3281 & ~n11296;
  assign n11298 = ~n3281 & ~n11297;
  assign n11299 = n3378 & ~n11298;
  assign n11300 = ~n10589 & ~n10827;
  assign n11301 = controllable_hmaster1 & ~n11300;
  assign n11302 = controllable_hmaster0 & ~n11300;
  assign n11303 = ~n11247 & ~n11302;
  assign n11304 = ~controllable_hmaster1 & ~n11303;
  assign n11305 = ~n11301 & ~n11304;
  assign n11306 = i_hbusreq3 & ~n11305;
  assign n11307 = ~n10611 & ~n11049;
  assign n11308 = controllable_hmaster1 & ~n11307;
  assign n11309 = controllable_hmaster0 & ~n11307;
  assign n11310 = ~n10624 & ~n11049;
  assign n11311 = ~controllable_hmaster0 & ~n11310;
  assign n11312 = ~n11309 & ~n11311;
  assign n11313 = ~controllable_hmaster1 & ~n11312;
  assign n11314 = ~n11308 & ~n11313;
  assign n11315 = ~i_hbusreq3 & ~n11314;
  assign n11316 = ~n11306 & ~n11315;
  assign n11317 = controllable_hmaster2 & ~n11316;
  assign n11318 = ~n10589 & ~n11066;
  assign n11319 = ~controllable_hmaster0 & ~n11318;
  assign n11320 = ~n11302 & ~n11319;
  assign n11321 = controllable_hmaster1 & ~n11320;
  assign n11322 = ~n10640 & ~n10827;
  assign n11323 = controllable_hmaster0 & ~n11322;
  assign n11324 = ~controllable_hmaster0 & ~n11300;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = ~controllable_hmaster1 & ~n11325;
  assign n11327 = ~n11321 & ~n11326;
  assign n11328 = i_hbusreq3 & ~n11327;
  assign n11329 = ~n10651 & ~n11049;
  assign n11330 = controllable_hmaster0 & ~n11329;
  assign n11331 = ~n10651 & ~n11110;
  assign n11332 = ~controllable_hmaster0 & ~n11331;
  assign n11333 = ~n11330 & ~n11332;
  assign n11334 = controllable_hmaster1 & ~n11333;
  assign n11335 = ~n10678 & ~n11049;
  assign n11336 = controllable_hmaster0 & ~n11335;
  assign n11337 = ~n10689 & ~n11127;
  assign n11338 = ~controllable_hmaster0 & ~n11337;
  assign n11339 = ~n11336 & ~n11338;
  assign n11340 = ~controllable_hmaster1 & ~n11339;
  assign n11341 = ~n11334 & ~n11340;
  assign n11342 = ~i_hbusreq3 & ~n11341;
  assign n11343 = ~n11328 & ~n11342;
  assign n11344 = ~controllable_hmaster2 & ~n11343;
  assign n11345 = ~n11317 & ~n11344;
  assign n11346 = ~controllable_hgrant3 & ~n11345;
  assign n11347 = ~n10110 & ~n11346;
  assign n11348 = controllable_nhgrant0 & ~n11347;
  assign n11349 = ~n10240 & ~n11348;
  assign n11350 = ~n3281 & ~n11349;
  assign n11351 = ~n3281 & ~n11350;
  assign n11352 = ~n3378 & ~n11351;
  assign n11353 = ~n11299 & ~n11352;
  assign n11354 = n3492 & ~n11353;
  assign n11355 = ~n8619 & ~n11354;
  assign n11356 = n3485 & ~n11355;
  assign n11357 = ~n8729 & ~n11356;
  assign n11358 = n3476 & ~n11357;
  assign n11359 = ~n11242 & ~n11358;
  assign n11360 = n3374 & ~n11359;
  assign n11361 = ~n11190 & ~n11360;
  assign n11362 = ~n3655 & ~n11361;
  assign n11363 = ~n11153 & ~n11362;
  assign n11364 = ~n3652 & ~n11363;
  assign n11365 = ~n10717 & ~n11364;
  assign n11366 = n3368 & ~n11365;
  assign n11367 = ~n9697 & ~n11366;
  assign n11368 = ~n3362 & ~n11367;
  assign n11369 = ~n8741 & ~n11368;
  assign n11370 = ~n3359 & ~n11369;
  assign n11371 = ~n8638 & ~n11370;
  assign n11372 = ~n3356 & ~n11371;
  assign n11373 = ~n4910 & ~n11372;
  assign n11374 = n3345 & ~n11373;
  assign n11375 = ~n3649 & ~n11374;
  assign n11376 = ~n3341 & ~n11375;
  assign n11377 = controllable_hmaster0 & ~n4926;
  assign n11378 = controllable_hmaster1 & ~n11377;
  assign n11379 = controllable_hmaster1 & ~n11378;
  assign n11380 = i_hlock3 & ~n11379;
  assign n11381 = controllable_hmaster0 & ~n4955;
  assign n11382 = controllable_hmaster1 & ~n11381;
  assign n11383 = controllable_hmaster1 & ~n11382;
  assign n11384 = ~i_hlock3 & ~n11383;
  assign n11385 = ~n11380 & ~n11384;
  assign n11386 = i_hbusreq3 & ~n11385;
  assign n11387 = controllable_hmaster0 & ~n4980;
  assign n11388 = controllable_hmaster1 & ~n11387;
  assign n11389 = controllable_hmaster1 & ~n11388;
  assign n11390 = i_hlock3 & ~n11389;
  assign n11391 = controllable_hmaster0 & ~n5027;
  assign n11392 = controllable_hmaster1 & ~n11391;
  assign n11393 = controllable_hmaster1 & ~n11392;
  assign n11394 = ~i_hlock3 & ~n11393;
  assign n11395 = ~n11390 & ~n11394;
  assign n11396 = ~i_hbusreq3 & ~n11395;
  assign n11397 = ~n11386 & ~n11396;
  assign n11398 = ~controllable_hmaster2 & ~n11397;
  assign n11399 = ~controllable_hmaster2 & ~n11398;
  assign n11400 = controllable_hgrant3 & ~n11399;
  assign n11401 = controllable_hmaster0 & ~n5078;
  assign n11402 = controllable_hmaster1 & ~n11401;
  assign n11403 = controllable_hmaster1 & ~n11402;
  assign n11404 = i_hlock3 & ~n11403;
  assign n11405 = controllable_hmaster0 & ~n5108;
  assign n11406 = controllable_hmaster1 & ~n11405;
  assign n11407 = controllable_hmaster1 & ~n11406;
  assign n11408 = ~i_hlock3 & ~n11407;
  assign n11409 = ~n11404 & ~n11408;
  assign n11410 = i_hbusreq3 & ~n11409;
  assign n11411 = controllable_hmaster0 & ~n5115;
  assign n11412 = controllable_hmaster1 & ~n11411;
  assign n11413 = controllable_hmaster1 & ~n11412;
  assign n11414 = i_hlock3 & ~n11413;
  assign n11415 = controllable_hmaster0 & ~n5153;
  assign n11416 = controllable_hmaster1 & ~n11415;
  assign n11417 = controllable_hmaster1 & ~n11416;
  assign n11418 = ~i_hlock3 & ~n11417;
  assign n11419 = ~n11414 & ~n11418;
  assign n11420 = ~i_hbusreq3 & ~n11419;
  assign n11421 = ~n11410 & ~n11420;
  assign n11422 = ~controllable_hmaster2 & ~n11421;
  assign n11423 = ~controllable_hmaster2 & ~n11422;
  assign n11424 = ~controllable_hgrant3 & ~n11423;
  assign n11425 = ~n11400 & ~n11424;
  assign n11426 = controllable_nhgrant0 & ~n11425;
  assign n11427 = ~controllable_nhgrant0 & ~n11423;
  assign n11428 = ~n11426 & ~n11427;
  assign n11429 = ~n3281 & ~n11428;
  assign n11430 = ~n3281 & ~n11429;
  assign n11431 = n3378 & ~n11430;
  assign n11432 = ~n3407 & ~n11398;
  assign n11433 = controllable_hgrant3 & ~n11432;
  assign n11434 = ~n3461 & ~n11422;
  assign n11435 = ~controllable_hgrant3 & ~n11434;
  assign n11436 = ~n11433 & ~n11435;
  assign n11437 = controllable_nhgrant0 & ~n11436;
  assign n11438 = ~n3407 & ~n11422;
  assign n11439 = ~controllable_nhgrant0 & ~n11438;
  assign n11440 = ~n11437 & ~n11439;
  assign n11441 = ~n3281 & ~n11440;
  assign n11442 = ~n3783 & ~n11441;
  assign n11443 = ~n3378 & ~n11442;
  assign n11444 = ~n11431 & ~n11443;
  assign n11445 = n3492 & ~n11444;
  assign n11446 = ~n3493 & ~n11445;
  assign n11447 = n3485 & ~n11446;
  assign n11448 = ~n3486 & ~n11447;
  assign n11449 = ~n3374 & ~n11448;
  assign n11450 = controllable_hmaster1 & ~n7064;
  assign n11451 = controllable_hmaster1 & ~n11450;
  assign n11452 = i_hbusreq3 & ~n11451;
  assign n11453 = controllable_hmaster0 & ~n5377;
  assign n11454 = controllable_hmaster1 & ~n11453;
  assign n11455 = controllable_hmaster1 & ~n11454;
  assign n11456 = ~i_hbusreq3 & ~n11455;
  assign n11457 = ~n11452 & ~n11456;
  assign n11458 = ~controllable_hmaster2 & ~n11457;
  assign n11459 = ~controllable_hmaster2 & ~n11458;
  assign n11460 = controllable_hgrant3 & ~n11459;
  assign n11461 = controllable_hmaster0 & ~n8771;
  assign n11462 = controllable_hmaster1 & ~n11461;
  assign n11463 = controllable_hmaster1 & ~n11462;
  assign n11464 = i_hbusreq3 & ~n11463;
  assign n11465 = controllable_hmaster0 & ~n8838;
  assign n11466 = controllable_hmaster1 & ~n11465;
  assign n11467 = controllable_hmaster1 & ~n11466;
  assign n11468 = ~i_hbusreq3 & ~n11467;
  assign n11469 = ~n11464 & ~n11468;
  assign n11470 = ~controllable_hmaster2 & ~n11469;
  assign n11471 = ~controllable_hmaster2 & ~n11470;
  assign n11472 = ~controllable_hgrant3 & ~n11471;
  assign n11473 = ~n11460 & ~n11472;
  assign n11474 = controllable_nhgrant0 & ~n11473;
  assign n11475 = controllable_hmaster1 & ~n3383;
  assign n11476 = controllable_hmaster1 & ~n11475;
  assign n11477 = i_hbusreq3 & ~n11476;
  assign n11478 = controllable_hmaster1 & ~n7083;
  assign n11479 = controllable_hmaster1 & ~n11478;
  assign n11480 = ~i_hbusreq3 & ~n11479;
  assign n11481 = ~n11477 & ~n11480;
  assign n11482 = ~controllable_hmaster2 & ~n11481;
  assign n11483 = ~controllable_hmaster2 & ~n11482;
  assign n11484 = controllable_hgrant3 & ~n11483;
  assign n11485 = controllable_hmaster1 & ~n7105;
  assign n11486 = controllable_hmaster1 & ~n11485;
  assign n11487 = i_hbusreq3 & ~n11486;
  assign n11488 = controllable_hmaster1 & ~n7109;
  assign n11489 = controllable_hmaster1 & ~n11488;
  assign n11490 = ~i_hbusreq3 & ~n11489;
  assign n11491 = ~n11487 & ~n11490;
  assign n11492 = ~controllable_hmaster2 & ~n11491;
  assign n11493 = ~controllable_hmaster2 & ~n11492;
  assign n11494 = ~controllable_hgrant3 & ~n11493;
  assign n11495 = ~n11484 & ~n11494;
  assign n11496 = ~controllable_nhgrant0 & ~n11495;
  assign n11497 = ~n11474 & ~n11496;
  assign n11498 = ~n3281 & ~n11497;
  assign n11499 = ~n3281 & ~n11498;
  assign n11500 = n3378 & ~n11499;
  assign n11501 = ~n3407 & ~n11458;
  assign n11502 = controllable_hgrant3 & ~n11501;
  assign n11503 = ~n3530 & ~n11470;
  assign n11504 = ~controllable_hgrant3 & ~n11503;
  assign n11505 = ~n11502 & ~n11504;
  assign n11506 = controllable_nhgrant0 & ~n11505;
  assign n11507 = ~n3407 & ~n11482;
  assign n11508 = controllable_hgrant3 & ~n11507;
  assign n11509 = ~n3407 & ~n11492;
  assign n11510 = ~controllable_hgrant3 & ~n11509;
  assign n11511 = ~n11508 & ~n11510;
  assign n11512 = ~controllable_nhgrant0 & ~n11511;
  assign n11513 = ~n11506 & ~n11512;
  assign n11514 = ~n3281 & ~n11513;
  assign n11515 = ~n3950 & ~n11514;
  assign n11516 = ~n3378 & ~n11515;
  assign n11517 = ~n11500 & ~n11516;
  assign n11518 = n3492 & ~n11517;
  assign n11519 = ~n3493 & ~n11518;
  assign n11520 = n3485 & ~n11519;
  assign n11521 = ~n3486 & ~n11520;
  assign n11522 = ~n3476 & ~n11521;
  assign n11523 = ~controllable_hgrant4 & ~n4001;
  assign n11524 = ~controllable_hgrant4 & ~n11523;
  assign n11525 = ~controllable_hgrant2 & ~n11524;
  assign n11526 = ~controllable_hgrant2 & ~n11525;
  assign n11527 = i_hbusreq3 & ~n11526;
  assign n11528 = i_hbusreq2 & ~n11524;
  assign n11529 = ~controllable_hgrant4 & ~n4039;
  assign n11530 = ~controllable_hgrant4 & ~n11529;
  assign n11531 = ~i_hbusreq2 & ~n11530;
  assign n11532 = ~n11528 & ~n11531;
  assign n11533 = ~controllable_hgrant2 & ~n11532;
  assign n11534 = ~controllable_hgrant2 & ~n11533;
  assign n11535 = ~i_hbusreq3 & ~n11534;
  assign n11536 = ~n11527 & ~n11535;
  assign n11537 = controllable_hmaster2 & ~n11536;
  assign n11538 = ~controllable_hmaster0 & ~n11526;
  assign n11539 = ~n5587 & ~n11538;
  assign n11540 = controllable_hmaster1 & ~n11539;
  assign n11541 = ~controllable_hmaster1 & ~n11526;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = i_hbusreq3 & ~n11542;
  assign n11544 = ~controllable_hmaster0 & ~n11534;
  assign n11545 = ~n5835 & ~n11544;
  assign n11546 = controllable_hmaster1 & ~n11545;
  assign n11547 = ~controllable_hmaster1 & ~n11534;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = ~i_hbusreq3 & ~n11548;
  assign n11550 = ~n11543 & ~n11549;
  assign n11551 = ~controllable_hmaster2 & ~n11550;
  assign n11552 = ~n11537 & ~n11551;
  assign n11553 = controllable_hgrant3 & ~n11552;
  assign n11554 = ~n11472 & ~n11553;
  assign n11555 = controllable_nhgrant0 & ~n11554;
  assign n11556 = ~n11496 & ~n11555;
  assign n11557 = ~n3281 & ~n11556;
  assign n11558 = ~n3281 & ~n11557;
  assign n11559 = n3378 & ~n11558;
  assign n11560 = ~n5758 & ~n11538;
  assign n11561 = ~controllable_hmaster1 & ~n11560;
  assign n11562 = ~n5757 & ~n11561;
  assign n11563 = i_hbusreq3 & ~n11562;
  assign n11564 = ~controllable_hgrant4 & ~n4116;
  assign n11565 = ~n3433 & ~n11564;
  assign n11566 = ~i_hbusreq2 & ~n11565;
  assign n11567 = ~n5550 & ~n11566;
  assign n11568 = ~controllable_hgrant2 & ~n11567;
  assign n11569 = ~n3431 & ~n11568;
  assign n11570 = controllable_hmaster1 & ~n11569;
  assign n11571 = controllable_hmaster0 & ~n11569;
  assign n11572 = ~n11544 & ~n11571;
  assign n11573 = ~controllable_hmaster1 & ~n11572;
  assign n11574 = ~n11570 & ~n11573;
  assign n11575 = ~i_hbusreq3 & ~n11574;
  assign n11576 = ~n11563 & ~n11575;
  assign n11577 = controllable_hmaster2 & ~n11576;
  assign n11578 = ~n11551 & ~n11577;
  assign n11579 = controllable_hgrant3 & ~n11578;
  assign n11580 = controllable_hmaster1 & ~n3557;
  assign n11581 = ~controllable_hmaster1 & ~n3555;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = i_hbusreq3 & ~n11582;
  assign n11584 = ~n3916 & ~n4134;
  assign n11585 = ~i_hbusreq2 & ~n11584;
  assign n11586 = ~n3561 & ~n11585;
  assign n11587 = ~controllable_hgrant2 & ~n11586;
  assign n11588 = ~n3859 & ~n11587;
  assign n11589 = controllable_hmaster0 & ~n11588;
  assign n11590 = ~n3596 & ~n11589;
  assign n11591 = controllable_hmaster1 & ~n11590;
  assign n11592 = ~controllable_hmaster1 & ~n3595;
  assign n11593 = ~n11591 & ~n11592;
  assign n11594 = ~i_hbusreq3 & ~n11593;
  assign n11595 = ~n11583 & ~n11594;
  assign n11596 = ~controllable_hmaster2 & ~n11595;
  assign n11597 = ~n3602 & ~n11596;
  assign n11598 = ~controllable_hgrant3 & ~n11597;
  assign n11599 = ~n11579 & ~n11598;
  assign n11600 = controllable_nhgrant0 & ~n11599;
  assign n11601 = ~n11512 & ~n11600;
  assign n11602 = ~n3281 & ~n11601;
  assign n11603 = ~n4089 & ~n11602;
  assign n11604 = ~n3378 & ~n11603;
  assign n11605 = ~n11559 & ~n11604;
  assign n11606 = n3492 & ~n11605;
  assign n11607 = ~n3493 & ~n11606;
  assign n11608 = n3485 & ~n11607;
  assign n11609 = ~n3486 & ~n11608;
  assign n11610 = n3476 & ~n11609;
  assign n11611 = ~n11522 & ~n11610;
  assign n11612 = n3374 & ~n11611;
  assign n11613 = ~n11449 & ~n11612;
  assign n11614 = n3655 & ~n11613;
  assign n11615 = controllable_hmaster0 & ~n9162;
  assign n11616 = controllable_hmaster1 & ~n11615;
  assign n11617 = controllable_hmaster1 & ~n11616;
  assign n11618 = i_hbusreq3 & ~n11617;
  assign n11619 = controllable_hmaster0 & ~n9186;
  assign n11620 = controllable_hmaster1 & ~n11619;
  assign n11621 = controllable_hmaster1 & ~n11620;
  assign n11622 = ~i_hbusreq3 & ~n11621;
  assign n11623 = ~n11618 & ~n11622;
  assign n11624 = ~controllable_hmaster2 & ~n11623;
  assign n11625 = ~controllable_hmaster2 & ~n11624;
  assign n11626 = ~controllable_hgrant3 & ~n11625;
  assign n11627 = ~n11460 & ~n11626;
  assign n11628 = controllable_nhgrant0 & ~n11627;
  assign n11629 = ~n11496 & ~n11628;
  assign n11630 = ~n3281 & ~n11629;
  assign n11631 = ~n3281 & ~n11630;
  assign n11632 = n3378 & ~n11631;
  assign n11633 = ~n3530 & ~n11624;
  assign n11634 = ~controllable_hgrant3 & ~n11633;
  assign n11635 = ~n11502 & ~n11634;
  assign n11636 = controllable_nhgrant0 & ~n11635;
  assign n11637 = ~n11512 & ~n11636;
  assign n11638 = ~n3281 & ~n11637;
  assign n11639 = ~n3950 & ~n11638;
  assign n11640 = ~n3378 & ~n11639;
  assign n11641 = ~n11632 & ~n11640;
  assign n11642 = n3492 & ~n11641;
  assign n11643 = ~n3493 & ~n11642;
  assign n11644 = n3485 & ~n11643;
  assign n11645 = ~n3486 & ~n11644;
  assign n11646 = ~n3476 & ~n11645;
  assign n11647 = ~n11553 & ~n11626;
  assign n11648 = controllable_nhgrant0 & ~n11647;
  assign n11649 = ~n11496 & ~n11648;
  assign n11650 = ~n3281 & ~n11649;
  assign n11651 = ~n3281 & ~n11650;
  assign n11652 = n3378 & ~n11651;
  assign n11653 = ~n3411 & ~n4279;
  assign n11654 = ~controllable_hgrant2 & ~n11653;
  assign n11655 = ~n3410 & ~n11654;
  assign n11656 = controllable_hmaster0 & ~n11655;
  assign n11657 = ~n3556 & ~n11656;
  assign n11658 = controllable_hmaster1 & ~n11657;
  assign n11659 = ~n11581 & ~n11658;
  assign n11660 = i_hbusreq3 & ~n11659;
  assign n11661 = i_hbusreq2 & ~n11653;
  assign n11662 = ~n3916 & ~n4300;
  assign n11663 = ~i_hbusreq2 & ~n11662;
  assign n11664 = ~n11661 & ~n11663;
  assign n11665 = ~controllable_hgrant2 & ~n11664;
  assign n11666 = ~n3859 & ~n11665;
  assign n11667 = controllable_hmaster0 & ~n11666;
  assign n11668 = ~n3596 & ~n11667;
  assign n11669 = controllable_hmaster1 & ~n11668;
  assign n11670 = ~n11592 & ~n11669;
  assign n11671 = ~i_hbusreq3 & ~n11670;
  assign n11672 = ~n11660 & ~n11671;
  assign n11673 = ~controllable_hmaster2 & ~n11672;
  assign n11674 = ~n3602 & ~n11673;
  assign n11675 = ~controllable_hgrant3 & ~n11674;
  assign n11676 = ~n11579 & ~n11675;
  assign n11677 = controllable_nhgrant0 & ~n11676;
  assign n11678 = ~n11512 & ~n11677;
  assign n11679 = ~n3281 & ~n11678;
  assign n11680 = ~n4089 & ~n11679;
  assign n11681 = ~n3378 & ~n11680;
  assign n11682 = ~n11652 & ~n11681;
  assign n11683 = n3492 & ~n11682;
  assign n11684 = ~n3493 & ~n11683;
  assign n11685 = n3485 & ~n11684;
  assign n11686 = ~n3486 & ~n11685;
  assign n11687 = n3476 & ~n11686;
  assign n11688 = ~n11646 & ~n11687;
  assign n11689 = n3374 & ~n11688;
  assign n11690 = ~n11449 & ~n11689;
  assign n11691 = ~n3655 & ~n11690;
  assign n11692 = ~n11614 & ~n11691;
  assign n11693 = n3652 & ~n11692;
  assign n11694 = controllable_hmaster0 & ~n9434;
  assign n11695 = controllable_hmaster1 & ~n11694;
  assign n11696 = controllable_hmaster1 & ~n11695;
  assign n11697 = i_hbusreq3 & ~n11696;
  assign n11698 = controllable_hmaster0 & ~n9447;
  assign n11699 = controllable_hmaster1 & ~n11698;
  assign n11700 = controllable_hmaster1 & ~n11699;
  assign n11701 = ~i_hbusreq3 & ~n11700;
  assign n11702 = ~n11697 & ~n11701;
  assign n11703 = ~controllable_hmaster2 & ~n11702;
  assign n11704 = ~controllable_hmaster2 & ~n11703;
  assign n11705 = ~controllable_hgrant3 & ~n11704;
  assign n11706 = ~n11460 & ~n11705;
  assign n11707 = controllable_nhgrant0 & ~n11706;
  assign n11708 = ~n11496 & ~n11707;
  assign n11709 = ~n3281 & ~n11708;
  assign n11710 = ~n3281 & ~n11709;
  assign n11711 = n3378 & ~n11710;
  assign n11712 = ~n3530 & ~n11703;
  assign n11713 = ~controllable_hgrant3 & ~n11712;
  assign n11714 = ~n11502 & ~n11713;
  assign n11715 = controllable_nhgrant0 & ~n11714;
  assign n11716 = ~n11512 & ~n11715;
  assign n11717 = ~n3281 & ~n11716;
  assign n11718 = ~n3950 & ~n11717;
  assign n11719 = ~n3378 & ~n11718;
  assign n11720 = ~n11711 & ~n11719;
  assign n11721 = n3492 & ~n11720;
  assign n11722 = ~n3493 & ~n11721;
  assign n11723 = n3485 & ~n11722;
  assign n11724 = ~n3486 & ~n11723;
  assign n11725 = ~n3476 & ~n11724;
  assign n11726 = ~n11553 & ~n11705;
  assign n11727 = controllable_nhgrant0 & ~n11726;
  assign n11728 = ~n11496 & ~n11727;
  assign n11729 = ~n3281 & ~n11728;
  assign n11730 = ~n3281 & ~n11729;
  assign n11731 = n3378 & ~n11730;
  assign n11732 = ~n3547 & ~n4333;
  assign n11733 = controllable_hmaster0 & ~n11732;
  assign n11734 = ~n3556 & ~n11733;
  assign n11735 = controllable_hmaster1 & ~n11734;
  assign n11736 = ~n11581 & ~n11735;
  assign n11737 = i_hbusreq3 & ~n11736;
  assign n11738 = ~n4340 & ~n11587;
  assign n11739 = controllable_hmaster0 & ~n11738;
  assign n11740 = ~n3596 & ~n11739;
  assign n11741 = controllable_hmaster1 & ~n11740;
  assign n11742 = ~n11592 & ~n11741;
  assign n11743 = ~i_hbusreq3 & ~n11742;
  assign n11744 = ~n11737 & ~n11743;
  assign n11745 = ~controllable_hmaster2 & ~n11744;
  assign n11746 = ~n3602 & ~n11745;
  assign n11747 = ~controllable_hgrant3 & ~n11746;
  assign n11748 = ~n11579 & ~n11747;
  assign n11749 = controllable_nhgrant0 & ~n11748;
  assign n11750 = ~n11512 & ~n11749;
  assign n11751 = ~n3281 & ~n11750;
  assign n11752 = ~n4089 & ~n11751;
  assign n11753 = ~n3378 & ~n11752;
  assign n11754 = ~n11731 & ~n11753;
  assign n11755 = n3492 & ~n11754;
  assign n11756 = ~n3493 & ~n11755;
  assign n11757 = n3485 & ~n11756;
  assign n11758 = ~n3486 & ~n11757;
  assign n11759 = n3476 & ~n11758;
  assign n11760 = ~n11725 & ~n11759;
  assign n11761 = n3374 & ~n11760;
  assign n11762 = ~n11449 & ~n11761;
  assign n11763 = n3655 & ~n11762;
  assign n11764 = controllable_hmaster0 & ~n9588;
  assign n11765 = controllable_hmaster1 & ~n11764;
  assign n11766 = controllable_hmaster1 & ~n11765;
  assign n11767 = i_hbusreq3 & ~n11766;
  assign n11768 = controllable_hmaster0 & ~n9601;
  assign n11769 = controllable_hmaster1 & ~n11768;
  assign n11770 = controllable_hmaster1 & ~n11769;
  assign n11771 = ~i_hbusreq3 & ~n11770;
  assign n11772 = ~n11767 & ~n11771;
  assign n11773 = ~controllable_hmaster2 & ~n11772;
  assign n11774 = ~controllable_hmaster2 & ~n11773;
  assign n11775 = ~controllable_hgrant3 & ~n11774;
  assign n11776 = ~n11460 & ~n11775;
  assign n11777 = controllable_nhgrant0 & ~n11776;
  assign n11778 = ~n11496 & ~n11777;
  assign n11779 = ~n3281 & ~n11778;
  assign n11780 = ~n3281 & ~n11779;
  assign n11781 = n3378 & ~n11780;
  assign n11782 = ~n3530 & ~n11773;
  assign n11783 = ~controllable_hgrant3 & ~n11782;
  assign n11784 = ~n11502 & ~n11783;
  assign n11785 = controllable_nhgrant0 & ~n11784;
  assign n11786 = ~n11512 & ~n11785;
  assign n11787 = ~n3281 & ~n11786;
  assign n11788 = ~n3950 & ~n11787;
  assign n11789 = ~n3378 & ~n11788;
  assign n11790 = ~n11781 & ~n11789;
  assign n11791 = n3492 & ~n11790;
  assign n11792 = ~n3493 & ~n11791;
  assign n11793 = n3485 & ~n11792;
  assign n11794 = ~n3486 & ~n11793;
  assign n11795 = ~n3476 & ~n11794;
  assign n11796 = ~n11553 & ~n11775;
  assign n11797 = controllable_nhgrant0 & ~n11796;
  assign n11798 = ~n11496 & ~n11797;
  assign n11799 = ~n3281 & ~n11798;
  assign n11800 = ~n3281 & ~n11799;
  assign n11801 = n3378 & ~n11800;
  assign n11802 = ~n4333 & ~n11654;
  assign n11803 = controllable_hmaster0 & ~n11802;
  assign n11804 = ~n3556 & ~n11803;
  assign n11805 = controllable_hmaster1 & ~n11804;
  assign n11806 = ~n11581 & ~n11805;
  assign n11807 = i_hbusreq3 & ~n11806;
  assign n11808 = ~n4340 & ~n11665;
  assign n11809 = controllable_hmaster0 & ~n11808;
  assign n11810 = ~n3596 & ~n11809;
  assign n11811 = controllable_hmaster1 & ~n11810;
  assign n11812 = ~n11592 & ~n11811;
  assign n11813 = ~i_hbusreq3 & ~n11812;
  assign n11814 = ~n11807 & ~n11813;
  assign n11815 = ~controllable_hmaster2 & ~n11814;
  assign n11816 = ~n3602 & ~n11815;
  assign n11817 = ~controllable_hgrant3 & ~n11816;
  assign n11818 = ~n11579 & ~n11817;
  assign n11819 = controllable_nhgrant0 & ~n11818;
  assign n11820 = ~n11512 & ~n11819;
  assign n11821 = ~n3281 & ~n11820;
  assign n11822 = ~n4089 & ~n11821;
  assign n11823 = ~n3378 & ~n11822;
  assign n11824 = ~n11801 & ~n11823;
  assign n11825 = n3492 & ~n11824;
  assign n11826 = ~n3493 & ~n11825;
  assign n11827 = n3485 & ~n11826;
  assign n11828 = ~n3486 & ~n11827;
  assign n11829 = n3476 & ~n11828;
  assign n11830 = ~n11795 & ~n11829;
  assign n11831 = n3374 & ~n11830;
  assign n11832 = ~n11449 & ~n11831;
  assign n11833 = ~n3655 & ~n11832;
  assign n11834 = ~n11763 & ~n11833;
  assign n11835 = ~n3652 & ~n11834;
  assign n11836 = ~n11693 & ~n11835;
  assign n11837 = ~n3368 & ~n11836;
  assign n11838 = controllable_hmaster0 & ~n9780;
  assign n11839 = controllable_hmaster1 & ~n11838;
  assign n11840 = controllable_hmaster1 & ~n11839;
  assign n11841 = ~i_hbusreq3 & ~n11840;
  assign n11842 = ~n11452 & ~n11841;
  assign n11843 = ~controllable_hmaster2 & ~n11842;
  assign n11844 = ~controllable_hmaster2 & ~n11843;
  assign n11845 = controllable_hgrant3 & ~n11844;
  assign n11846 = controllable_hmaster0 & ~n9802;
  assign n11847 = controllable_hmaster1 & ~n11846;
  assign n11848 = controllable_hmaster1 & ~n11847;
  assign n11849 = ~i_hbusreq3 & ~n11848;
  assign n11850 = ~n11464 & ~n11849;
  assign n11851 = ~controllable_hmaster2 & ~n11850;
  assign n11852 = ~controllable_hmaster2 & ~n11851;
  assign n11853 = ~controllable_hgrant3 & ~n11852;
  assign n11854 = ~n11845 & ~n11853;
  assign n11855 = controllable_nhgrant0 & ~n11854;
  assign n11856 = controllable_hmaster1 & ~n9701;
  assign n11857 = controllable_hmaster1 & ~n11856;
  assign n11858 = ~i_hbusreq3 & ~n11857;
  assign n11859 = ~n11477 & ~n11858;
  assign n11860 = ~controllable_hmaster2 & ~n11859;
  assign n11861 = ~controllable_hmaster2 & ~n11860;
  assign n11862 = controllable_hgrant3 & ~n11861;
  assign n11863 = controllable_hmaster1 & ~n9738;
  assign n11864 = controllable_hmaster1 & ~n11863;
  assign n11865 = i_hbusreq3 & ~n11864;
  assign n11866 = controllable_hmaster1 & ~n9744;
  assign n11867 = controllable_hmaster1 & ~n11866;
  assign n11868 = ~i_hbusreq3 & ~n11867;
  assign n11869 = ~n11865 & ~n11868;
  assign n11870 = ~controllable_hmaster2 & ~n11869;
  assign n11871 = ~controllable_hmaster2 & ~n11870;
  assign n11872 = ~controllable_hgrant3 & ~n11871;
  assign n11873 = ~n11862 & ~n11872;
  assign n11874 = ~controllable_nhgrant0 & ~n11873;
  assign n11875 = ~n11855 & ~n11874;
  assign n11876 = ~n3281 & ~n11875;
  assign n11877 = ~n3281 & ~n11876;
  assign n11878 = n3492 & ~n11877;
  assign n11879 = n3492 & ~n11878;
  assign n11880 = n3485 & ~n11879;
  assign n11881 = n3485 & ~n11880;
  assign n11882 = ~n3476 & ~n11881;
  assign n11883 = controllable_hmaster2 & ~n11526;
  assign n11884 = ~n10098 & ~n11538;
  assign n11885 = controllable_hmaster1 & ~n11884;
  assign n11886 = ~n11541 & ~n11885;
  assign n11887 = ~i_hbusreq3 & ~n11886;
  assign n11888 = ~n11543 & ~n11887;
  assign n11889 = ~controllable_hmaster2 & ~n11888;
  assign n11890 = ~n11883 & ~n11889;
  assign n11891 = controllable_hgrant3 & ~n11890;
  assign n11892 = ~n11853 & ~n11891;
  assign n11893 = controllable_nhgrant0 & ~n11892;
  assign n11894 = ~n11874 & ~n11893;
  assign n11895 = ~n3281 & ~n11894;
  assign n11896 = ~n3281 & ~n11895;
  assign n11897 = n3492 & ~n11896;
  assign n11898 = n3492 & ~n11897;
  assign n11899 = n3485 & ~n11898;
  assign n11900 = n3485 & ~n11899;
  assign n11901 = n3476 & ~n11900;
  assign n11902 = ~n11882 & ~n11901;
  assign n11903 = n3374 & ~n11902;
  assign n11904 = n3374 & ~n11903;
  assign n11905 = n3655 & ~n11904;
  assign n11906 = controllable_hmaster0 & ~n10326;
  assign n11907 = controllable_hmaster1 & ~n11906;
  assign n11908 = controllable_hmaster1 & ~n11907;
  assign n11909 = i_hbusreq3 & ~n11908;
  assign n11910 = controllable_hmaster0 & ~n10348;
  assign n11911 = controllable_hmaster1 & ~n11910;
  assign n11912 = controllable_hmaster1 & ~n11911;
  assign n11913 = ~i_hbusreq3 & ~n11912;
  assign n11914 = ~n11909 & ~n11913;
  assign n11915 = ~controllable_hmaster2 & ~n11914;
  assign n11916 = ~controllable_hmaster2 & ~n11915;
  assign n11917 = ~controllable_hgrant3 & ~n11916;
  assign n11918 = ~n11845 & ~n11917;
  assign n11919 = controllable_nhgrant0 & ~n11918;
  assign n11920 = ~n11874 & ~n11919;
  assign n11921 = ~n3281 & ~n11920;
  assign n11922 = ~n3281 & ~n11921;
  assign n11923 = n3492 & ~n11922;
  assign n11924 = n3492 & ~n11923;
  assign n11925 = n3485 & ~n11924;
  assign n11926 = n3485 & ~n11925;
  assign n11927 = ~n3476 & ~n11926;
  assign n11928 = ~n11891 & ~n11917;
  assign n11929 = controllable_nhgrant0 & ~n11928;
  assign n11930 = ~n11874 & ~n11929;
  assign n11931 = ~n3281 & ~n11930;
  assign n11932 = ~n3281 & ~n11931;
  assign n11933 = n3492 & ~n11932;
  assign n11934 = n3492 & ~n11933;
  assign n11935 = n3485 & ~n11934;
  assign n11936 = n3485 & ~n11935;
  assign n11937 = n3476 & ~n11936;
  assign n11938 = ~n11927 & ~n11937;
  assign n11939 = n3374 & ~n11938;
  assign n11940 = n3374 & ~n11939;
  assign n11941 = ~n3655 & ~n11940;
  assign n11942 = ~n11905 & ~n11941;
  assign n11943 = n3652 & ~n11942;
  assign n11944 = controllable_hmaster0 & ~n10767;
  assign n11945 = controllable_hmaster1 & ~n11944;
  assign n11946 = controllable_hmaster1 & ~n11945;
  assign n11947 = i_hbusreq3 & ~n11946;
  assign n11948 = controllable_hmaster0 & ~n10781;
  assign n11949 = controllable_hmaster1 & ~n11948;
  assign n11950 = controllable_hmaster1 & ~n11949;
  assign n11951 = ~i_hbusreq3 & ~n11950;
  assign n11952 = ~n11947 & ~n11951;
  assign n11953 = ~controllable_hmaster2 & ~n11952;
  assign n11954 = ~controllable_hmaster2 & ~n11953;
  assign n11955 = ~controllable_hgrant3 & ~n11954;
  assign n11956 = ~n11845 & ~n11955;
  assign n11957 = controllable_nhgrant0 & ~n11956;
  assign n11958 = ~n11874 & ~n11957;
  assign n11959 = ~n3281 & ~n11958;
  assign n11960 = ~n3281 & ~n11959;
  assign n11961 = n3492 & ~n11960;
  assign n11962 = n3492 & ~n11961;
  assign n11963 = n3485 & ~n11962;
  assign n11964 = n3485 & ~n11963;
  assign n11965 = ~n3476 & ~n11964;
  assign n11966 = ~n11891 & ~n11955;
  assign n11967 = controllable_nhgrant0 & ~n11966;
  assign n11968 = ~n11874 & ~n11967;
  assign n11969 = ~n3281 & ~n11968;
  assign n11970 = ~n3281 & ~n11969;
  assign n11971 = n3492 & ~n11970;
  assign n11972 = n3492 & ~n11971;
  assign n11973 = n3485 & ~n11972;
  assign n11974 = n3485 & ~n11973;
  assign n11975 = n3476 & ~n11974;
  assign n11976 = ~n11965 & ~n11975;
  assign n11977 = n3374 & ~n11976;
  assign n11978 = n3374 & ~n11977;
  assign n11979 = n3655 & ~n11978;
  assign n11980 = controllable_hmaster0 & ~n11203;
  assign n11981 = controllable_hmaster1 & ~n11980;
  assign n11982 = controllable_hmaster1 & ~n11981;
  assign n11983 = i_hbusreq3 & ~n11982;
  assign n11984 = controllable_hmaster0 & ~n11216;
  assign n11985 = controllable_hmaster1 & ~n11984;
  assign n11986 = controllable_hmaster1 & ~n11985;
  assign n11987 = ~i_hbusreq3 & ~n11986;
  assign n11988 = ~n11983 & ~n11987;
  assign n11989 = ~controllable_hmaster2 & ~n11988;
  assign n11990 = ~controllable_hmaster2 & ~n11989;
  assign n11991 = ~controllable_hgrant3 & ~n11990;
  assign n11992 = ~n11845 & ~n11991;
  assign n11993 = controllable_nhgrant0 & ~n11992;
  assign n11994 = ~n11874 & ~n11993;
  assign n11995 = ~n3281 & ~n11994;
  assign n11996 = ~n3281 & ~n11995;
  assign n11997 = n3492 & ~n11996;
  assign n11998 = n3492 & ~n11997;
  assign n11999 = n3485 & ~n11998;
  assign n12000 = n3485 & ~n11999;
  assign n12001 = ~n3476 & ~n12000;
  assign n12002 = ~n11891 & ~n11991;
  assign n12003 = controllable_nhgrant0 & ~n12002;
  assign n12004 = ~n11874 & ~n12003;
  assign n12005 = ~n3281 & ~n12004;
  assign n12006 = ~n3281 & ~n12005;
  assign n12007 = n3492 & ~n12006;
  assign n12008 = n3492 & ~n12007;
  assign n12009 = n3485 & ~n12008;
  assign n12010 = n3485 & ~n12009;
  assign n12011 = n3476 & ~n12010;
  assign n12012 = ~n12001 & ~n12011;
  assign n12013 = n3374 & ~n12012;
  assign n12014 = n3374 & ~n12013;
  assign n12015 = ~n3655 & ~n12014;
  assign n12016 = ~n11979 & ~n12015;
  assign n12017 = ~n3652 & ~n12016;
  assign n12018 = ~n11943 & ~n12017;
  assign n12019 = n3368 & ~n12018;
  assign n12020 = ~n11837 & ~n12019;
  assign n12021 = ~n3362 & ~n12020;
  assign n12022 = ~n3362 & ~n12021;
  assign n12023 = ~n3359 & ~n12022;
  assign n12024 = ~n3359 & ~n12023;
  assign n12025 = n3356 & ~n12024;
  assign n12026 = n3378 & ~n11442;
  assign n12027 = ~n5249 & ~n12026;
  assign n12028 = n3492 & ~n12027;
  assign n12029 = ~n3631 & ~n12028;
  assign n12030 = n3485 & ~n12029;
  assign n12031 = ~n3630 & ~n12030;
  assign n12032 = ~n3374 & ~n12031;
  assign n12033 = controllable_hmaster2 & ~n5344;
  assign n12034 = ~n5278 & ~n5377;
  assign n12035 = controllable_hmaster1 & ~n12034;
  assign n12036 = ~n5281 & ~n12035;
  assign n12037 = ~i_hbusreq3 & ~n12036;
  assign n12038 = ~n5265 & ~n12037;
  assign n12039 = ~controllable_hmaster2 & ~n12038;
  assign n12040 = ~n12033 & ~n12039;
  assign n12041 = controllable_hgrant3 & ~n12040;
  assign n12042 = ~controllable_hgrant4 & ~n3380;
  assign n12043 = ~n3848 & ~n12042;
  assign n12044 = ~controllable_hgrant2 & ~n12043;
  assign n12045 = ~n3410 & ~n12044;
  assign n12046 = ~controllable_hmaster0 & ~n12045;
  assign n12047 = ~n3502 & ~n12046;
  assign n12048 = ~controllable_hmaster1 & ~n12047;
  assign n12049 = ~n3501 & ~n12048;
  assign n12050 = i_hbusreq3 & ~n12049;
  assign n12051 = i_hbusreq2 & ~n12043;
  assign n12052 = controllable_hgrant4 & ~n5270;
  assign n12053 = ~controllable_hgrant4 & ~n3397;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = ~i_hbusreq2 & ~n12054;
  assign n12056 = ~n12051 & ~n12055;
  assign n12057 = ~controllable_hgrant2 & ~n12056;
  assign n12058 = ~n3431 & ~n12057;
  assign n12059 = ~controllable_hmaster0 & ~n12058;
  assign n12060 = ~n3524 & ~n12059;
  assign n12061 = ~controllable_hmaster1 & ~n12060;
  assign n12062 = ~n3523 & ~n12061;
  assign n12063 = ~i_hbusreq3 & ~n12062;
  assign n12064 = ~n12050 & ~n12063;
  assign n12065 = controllable_hmaster2 & ~n12064;
  assign n12066 = ~n5291 & ~n8771;
  assign n12067 = controllable_hmaster1 & ~n12066;
  assign n12068 = ~n5305 & ~n12067;
  assign n12069 = i_hbusreq3 & ~n12068;
  assign n12070 = ~n5311 & ~n8838;
  assign n12071 = controllable_hmaster1 & ~n12070;
  assign n12072 = ~n5334 & ~n12071;
  assign n12073 = ~i_hbusreq3 & ~n12072;
  assign n12074 = ~n12069 & ~n12073;
  assign n12075 = ~controllable_hmaster2 & ~n12074;
  assign n12076 = ~n12065 & ~n12075;
  assign n12077 = ~controllable_hgrant3 & ~n12076;
  assign n12078 = ~n12041 & ~n12077;
  assign n12079 = controllable_nhgrant0 & ~n12078;
  assign n12080 = ~n4913 & ~n5278;
  assign n12081 = controllable_hmaster1 & ~n12080;
  assign n12082 = ~n5281 & ~n12081;
  assign n12083 = ~i_hbusreq3 & ~n12082;
  assign n12084 = ~n3951 & ~n12083;
  assign n12085 = ~controllable_hmaster2 & ~n12084;
  assign n12086 = ~n12033 & ~n12085;
  assign n12087 = controllable_hgrant3 & ~n12086;
  assign n12088 = ~n3821 & ~n5191;
  assign n12089 = controllable_hmaster1 & ~n12088;
  assign n12090 = ~n5350 & ~n12089;
  assign n12091 = i_hbusreq3 & ~n12090;
  assign n12092 = ~n5197 & ~n5278;
  assign n12093 = controllable_hmaster1 & ~n12092;
  assign n12094 = ~n5355 & ~n12093;
  assign n12095 = ~i_hbusreq3 & ~n12094;
  assign n12096 = ~n12091 & ~n12095;
  assign n12097 = ~controllable_hmaster2 & ~n12096;
  assign n12098 = ~n12033 & ~n12097;
  assign n12099 = ~controllable_hgrant3 & ~n12098;
  assign n12100 = ~n12087 & ~n12099;
  assign n12101 = ~controllable_nhgrant0 & ~n12100;
  assign n12102 = ~n12079 & ~n12101;
  assign n12103 = ~n3281 & ~n12102;
  assign n12104 = ~n3950 & ~n12103;
  assign n12105 = n3378 & ~n12104;
  assign n12106 = ~n3848 & ~n3906;
  assign n12107 = ~controllable_hgrant2 & ~n12106;
  assign n12108 = ~n3410 & ~n12107;
  assign n12109 = ~controllable_hmaster0 & ~n12108;
  assign n12110 = ~n3502 & ~n12109;
  assign n12111 = ~controllable_hmaster1 & ~n12110;
  assign n12112 = ~n3501 & ~n12111;
  assign n12113 = i_hbusreq3 & ~n12112;
  assign n12114 = i_hbusreq2 & ~n12106;
  assign n12115 = ~n3873 & ~n3929;
  assign n12116 = ~i_hbusreq2 & ~n12115;
  assign n12117 = ~n12114 & ~n12116;
  assign n12118 = ~controllable_hgrant2 & ~n12117;
  assign n12119 = ~n3859 & ~n12118;
  assign n12120 = ~controllable_hmaster0 & ~n12119;
  assign n12121 = ~n5417 & ~n12120;
  assign n12122 = ~controllable_hmaster1 & ~n12121;
  assign n12123 = ~n5416 & ~n12122;
  assign n12124 = ~i_hbusreq3 & ~n12123;
  assign n12125 = ~n12113 & ~n12124;
  assign n12126 = controllable_hmaster2 & ~n12125;
  assign n12127 = ~n5425 & ~n8771;
  assign n12128 = controllable_hmaster1 & ~n12127;
  assign n12129 = ~n5435 & ~n12128;
  assign n12130 = i_hbusreq3 & ~n12129;
  assign n12131 = ~n5440 & ~n8838;
  assign n12132 = controllable_hmaster1 & ~n12131;
  assign n12133 = ~n5480 & ~n12132;
  assign n12134 = ~i_hbusreq3 & ~n12133;
  assign n12135 = ~n12130 & ~n12134;
  assign n12136 = ~controllable_hmaster2 & ~n12135;
  assign n12137 = ~n12126 & ~n12136;
  assign n12138 = ~controllable_hgrant3 & ~n12137;
  assign n12139 = ~n5402 & ~n12138;
  assign n12140 = controllable_nhgrant0 & ~n12139;
  assign n12141 = ~n5534 & ~n12140;
  assign n12142 = ~n3281 & ~n12141;
  assign n12143 = ~n3950 & ~n12142;
  assign n12144 = ~n3378 & ~n12143;
  assign n12145 = ~n12105 & ~n12144;
  assign n12146 = n3492 & ~n12145;
  assign n12147 = ~n3631 & ~n12146;
  assign n12148 = n3485 & ~n12147;
  assign n12149 = ~n3630 & ~n12148;
  assign n12150 = ~n3476 & ~n12149;
  assign n12151 = ~i_hbusreq3 & ~n11569;
  assign n12152 = ~n5549 & ~n12151;
  assign n12153 = controllable_hmaster2 & ~n12152;
  assign n12154 = ~controllable_hmaster0 & ~n11569;
  assign n12155 = ~n5835 & ~n12154;
  assign n12156 = controllable_hmaster1 & ~n12155;
  assign n12157 = ~controllable_hmaster1 & ~n11569;
  assign n12158 = ~n12156 & ~n12157;
  assign n12159 = ~i_hbusreq3 & ~n12158;
  assign n12160 = ~n5593 & ~n12159;
  assign n12161 = ~controllable_hmaster2 & ~n12160;
  assign n12162 = ~n12153 & ~n12161;
  assign n12163 = controllable_hgrant3 & ~n12162;
  assign n12164 = ~n4015 & ~n5681;
  assign n12165 = ~controllable_hgrant2 & ~n12164;
  assign n12166 = ~n5616 & ~n12165;
  assign n12167 = ~controllable_hmaster0 & ~n12166;
  assign n12168 = ~n5626 & ~n12167;
  assign n12169 = ~controllable_hmaster1 & ~n12168;
  assign n12170 = ~n5625 & ~n12169;
  assign n12171 = i_hbusreq3 & ~n12170;
  assign n12172 = controllable_hgrant4 & ~n5554;
  assign n12173 = ~n5649 & ~n12172;
  assign n12174 = ~i_hbusreq2 & ~n12173;
  assign n12175 = ~n5636 & ~n12174;
  assign n12176 = ~controllable_hgrant2 & ~n12175;
  assign n12177 = ~n5635 & ~n12176;
  assign n12178 = controllable_hmaster1 & ~n12177;
  assign n12179 = controllable_hmaster0 & ~n12177;
  assign n12180 = i_hbusreq2 & ~n12164;
  assign n12181 = controllable_hgrant4 & ~n5598;
  assign n12182 = ~n5715 & ~n12181;
  assign n12183 = ~i_hbusreq2 & ~n12182;
  assign n12184 = ~n12180 & ~n12183;
  assign n12185 = ~controllable_hgrant2 & ~n12184;
  assign n12186 = ~n5635 & ~n12185;
  assign n12187 = ~controllable_hmaster0 & ~n12186;
  assign n12188 = ~n12179 & ~n12187;
  assign n12189 = ~controllable_hmaster1 & ~n12188;
  assign n12190 = ~n12178 & ~n12189;
  assign n12191 = ~i_hbusreq3 & ~n12190;
  assign n12192 = ~n12171 & ~n12191;
  assign n12193 = controllable_hmaster2 & ~n12192;
  assign n12194 = ~n5626 & ~n5688;
  assign n12195 = controllable_hmaster1 & ~n12194;
  assign n12196 = ~n5704 & ~n12195;
  assign n12197 = i_hbusreq3 & ~n12196;
  assign n12198 = controllable_hgrant4 & ~n5569;
  assign n12199 = ~n5667 & ~n12198;
  assign n12200 = ~i_hbusreq2 & ~n12199;
  assign n12201 = ~n5636 & ~n12200;
  assign n12202 = ~controllable_hgrant2 & ~n12201;
  assign n12203 = ~n5657 & ~n12202;
  assign n12204 = controllable_hmaster0 & ~n12203;
  assign n12205 = ~n5715 & ~n12172;
  assign n12206 = ~i_hbusreq2 & ~n12205;
  assign n12207 = ~n5707 & ~n12206;
  assign n12208 = ~controllable_hgrant2 & ~n12207;
  assign n12209 = ~n5722 & ~n12208;
  assign n12210 = ~controllable_hmaster0 & ~n12209;
  assign n12211 = ~n12204 & ~n12210;
  assign n12212 = controllable_hmaster1 & ~n12211;
  assign n12213 = ~n5739 & ~n12172;
  assign n12214 = ~i_hbusreq2 & ~n12213;
  assign n12215 = ~n5727 & ~n12214;
  assign n12216 = ~controllable_hgrant2 & ~n12215;
  assign n12217 = ~n5635 & ~n12216;
  assign n12218 = controllable_hmaster0 & ~n12217;
  assign n12219 = ~n5635 & ~n12208;
  assign n12220 = ~controllable_hmaster0 & ~n12219;
  assign n12221 = ~n12218 & ~n12220;
  assign n12222 = ~controllable_hmaster1 & ~n12221;
  assign n12223 = ~n12212 & ~n12222;
  assign n12224 = ~i_hbusreq3 & ~n12223;
  assign n12225 = ~n12197 & ~n12224;
  assign n12226 = ~controllable_hmaster2 & ~n12225;
  assign n12227 = ~n12193 & ~n12226;
  assign n12228 = ~controllable_hgrant3 & ~n12227;
  assign n12229 = ~n12163 & ~n12228;
  assign n12230 = controllable_nhgrant0 & ~n12229;
  assign n12231 = ~i_hbusreq3 & ~n5560;
  assign n12232 = ~n5549 & ~n12231;
  assign n12233 = controllable_hmaster2 & ~n12232;
  assign n12234 = controllable_hmaster0 & ~n5763;
  assign n12235 = ~n5588 & ~n12234;
  assign n12236 = controllable_hmaster1 & ~n12235;
  assign n12237 = ~n5796 & ~n12236;
  assign n12238 = i_hbusreq3 & ~n12237;
  assign n12239 = controllable_hmaster0 & ~n5786;
  assign n12240 = ~n5606 & ~n12239;
  assign n12241 = controllable_hmaster1 & ~n12240;
  assign n12242 = ~n5801 & ~n12241;
  assign n12243 = ~i_hbusreq3 & ~n12242;
  assign n12244 = ~n12238 & ~n12243;
  assign n12245 = ~controllable_hmaster2 & ~n12244;
  assign n12246 = ~n12233 & ~n12245;
  assign n12247 = ~controllable_hgrant3 & ~n12246;
  assign n12248 = ~n12087 & ~n12247;
  assign n12249 = ~controllable_nhgrant0 & ~n12248;
  assign n12250 = ~n12230 & ~n12249;
  assign n12251 = ~n3281 & ~n12250;
  assign n12252 = ~n4089 & ~n12251;
  assign n12253 = n3378 & ~n12252;
  assign n12254 = ~n4015 & ~n5911;
  assign n12255 = ~controllable_hgrant2 & ~n12254;
  assign n12256 = ~n5616 & ~n12255;
  assign n12257 = ~controllable_hmaster0 & ~n12256;
  assign n12258 = ~n5626 & ~n12257;
  assign n12259 = ~controllable_hmaster1 & ~n12258;
  assign n12260 = ~n5625 & ~n12259;
  assign n12261 = i_hbusreq3 & ~n12260;
  assign n12262 = i_hbusreq2 & ~n12254;
  assign n12263 = ~n4064 & ~n5943;
  assign n12264 = ~i_hbusreq2 & ~n12263;
  assign n12265 = ~n12262 & ~n12264;
  assign n12266 = ~controllable_hgrant2 & ~n12265;
  assign n12267 = ~n5862 & ~n12266;
  assign n12268 = ~controllable_hmaster0 & ~n12267;
  assign n12269 = ~n5884 & ~n12268;
  assign n12270 = ~controllable_hmaster1 & ~n12269;
  assign n12271 = ~n5883 & ~n12270;
  assign n12272 = ~i_hbusreq3 & ~n12271;
  assign n12273 = ~n12261 & ~n12272;
  assign n12274 = controllable_hmaster2 & ~n12273;
  assign n12275 = ~n5626 & ~n5917;
  assign n12276 = controllable_hmaster1 & ~n12275;
  assign n12277 = ~n5928 & ~n12276;
  assign n12278 = i_hbusreq3 & ~n12277;
  assign n12279 = ~n5863 & ~n5897;
  assign n12280 = ~i_hbusreq2 & ~n12279;
  assign n12281 = ~n5636 & ~n12280;
  assign n12282 = ~controllable_hgrant2 & ~n12281;
  assign n12283 = ~n5862 & ~n12282;
  assign n12284 = controllable_hmaster0 & ~n12283;
  assign n12285 = ~n5952 & ~n12284;
  assign n12286 = controllable_hmaster1 & ~n12285;
  assign n12287 = ~n5998 & ~n12286;
  assign n12288 = ~i_hbusreq3 & ~n12287;
  assign n12289 = ~n12278 & ~n12288;
  assign n12290 = ~controllable_hmaster2 & ~n12289;
  assign n12291 = ~n12274 & ~n12290;
  assign n12292 = ~controllable_hgrant3 & ~n12291;
  assign n12293 = ~n5861 & ~n12292;
  assign n12294 = controllable_nhgrant0 & ~n12293;
  assign n12295 = ~n6082 & ~n12294;
  assign n12296 = ~n3281 & ~n12295;
  assign n12297 = ~n4089 & ~n12296;
  assign n12298 = ~n3378 & ~n12297;
  assign n12299 = ~n12253 & ~n12298;
  assign n12300 = n3492 & ~n12299;
  assign n12301 = ~n3631 & ~n12300;
  assign n12302 = n3485 & ~n12301;
  assign n12303 = ~n3630 & ~n12302;
  assign n12304 = n3476 & ~n12303;
  assign n12305 = ~n12150 & ~n12304;
  assign n12306 = n3374 & ~n12305;
  assign n12307 = ~n12032 & ~n12306;
  assign n12308 = n3655 & ~n12307;
  assign n12309 = ~n6196 & ~n12026;
  assign n12310 = n3492 & ~n12309;
  assign n12311 = ~n3631 & ~n12310;
  assign n12312 = n3485 & ~n12311;
  assign n12313 = ~n3630 & ~n12312;
  assign n12314 = ~n3374 & ~n12313;
  assign n12315 = ~n5291 & ~n9162;
  assign n12316 = controllable_hmaster1 & ~n12315;
  assign n12317 = ~n5305 & ~n12316;
  assign n12318 = i_hbusreq3 & ~n12317;
  assign n12319 = ~n5311 & ~n9186;
  assign n12320 = controllable_hmaster1 & ~n12319;
  assign n12321 = ~n5334 & ~n12320;
  assign n12322 = ~i_hbusreq3 & ~n12321;
  assign n12323 = ~n12318 & ~n12322;
  assign n12324 = ~controllable_hmaster2 & ~n12323;
  assign n12325 = ~n12065 & ~n12324;
  assign n12326 = ~controllable_hgrant3 & ~n12325;
  assign n12327 = ~n12041 & ~n12326;
  assign n12328 = controllable_nhgrant0 & ~n12327;
  assign n12329 = ~n12101 & ~n12328;
  assign n12330 = ~n3281 & ~n12329;
  assign n12331 = ~n3950 & ~n12330;
  assign n12332 = n3378 & ~n12331;
  assign n12333 = ~n3848 & ~n6250;
  assign n12334 = ~controllable_hgrant2 & ~n12333;
  assign n12335 = ~n3410 & ~n12334;
  assign n12336 = ~controllable_hmaster0 & ~n12335;
  assign n12337 = ~n6217 & ~n12336;
  assign n12338 = ~controllable_hmaster1 & ~n12337;
  assign n12339 = ~n6216 & ~n12338;
  assign n12340 = i_hbusreq3 & ~n12339;
  assign n12341 = i_hbusreq2 & ~n12333;
  assign n12342 = ~n3873 & ~n6287;
  assign n12343 = ~i_hbusreq2 & ~n12342;
  assign n12344 = ~n12341 & ~n12343;
  assign n12345 = ~controllable_hgrant2 & ~n12344;
  assign n12346 = ~n3859 & ~n12345;
  assign n12347 = ~controllable_hmaster0 & ~n12346;
  assign n12348 = ~n6240 & ~n12347;
  assign n12349 = ~controllable_hmaster1 & ~n12348;
  assign n12350 = ~n6239 & ~n12349;
  assign n12351 = ~i_hbusreq3 & ~n12350;
  assign n12352 = ~n12340 & ~n12351;
  assign n12353 = controllable_hmaster2 & ~n12352;
  assign n12354 = ~n6256 & ~n9162;
  assign n12355 = controllable_hmaster1 & ~n12354;
  assign n12356 = ~n6271 & ~n12355;
  assign n12357 = i_hbusreq3 & ~n12356;
  assign n12358 = ~n6295 & ~n9186;
  assign n12359 = controllable_hmaster1 & ~n12358;
  assign n12360 = ~n6339 & ~n12359;
  assign n12361 = ~i_hbusreq3 & ~n12360;
  assign n12362 = ~n12357 & ~n12361;
  assign n12363 = ~controllable_hmaster2 & ~n12362;
  assign n12364 = ~n12353 & ~n12363;
  assign n12365 = ~controllable_hgrant3 & ~n12364;
  assign n12366 = ~n5402 & ~n12365;
  assign n12367 = controllable_nhgrant0 & ~n12366;
  assign n12368 = ~n5534 & ~n12367;
  assign n12369 = ~n3281 & ~n12368;
  assign n12370 = ~n3950 & ~n12369;
  assign n12371 = ~n3378 & ~n12370;
  assign n12372 = ~n12332 & ~n12371;
  assign n12373 = n3492 & ~n12372;
  assign n12374 = ~n3631 & ~n12373;
  assign n12375 = n3485 & ~n12374;
  assign n12376 = ~n3630 & ~n12375;
  assign n12377 = ~n3476 & ~n12376;
  assign n12378 = ~n4091 & ~n6359;
  assign n12379 = ~controllable_hgrant2 & ~n12378;
  assign n12380 = ~n5616 & ~n12379;
  assign n12381 = controllable_hmaster0 & ~n12380;
  assign n12382 = ~n5688 & ~n12381;
  assign n12383 = controllable_hmaster1 & ~n12382;
  assign n12384 = ~n5704 & ~n12383;
  assign n12385 = i_hbusreq3 & ~n12384;
  assign n12386 = i_hbusreq2 & ~n12378;
  assign n12387 = ~n6380 & ~n12198;
  assign n12388 = ~i_hbusreq2 & ~n12387;
  assign n12389 = ~n12386 & ~n12388;
  assign n12390 = ~controllable_hgrant2 & ~n12389;
  assign n12391 = ~n5657 & ~n12390;
  assign n12392 = controllable_hmaster0 & ~n12391;
  assign n12393 = ~n12210 & ~n12392;
  assign n12394 = controllable_hmaster1 & ~n12393;
  assign n12395 = ~n12222 & ~n12394;
  assign n12396 = ~i_hbusreq3 & ~n12395;
  assign n12397 = ~n12385 & ~n12396;
  assign n12398 = ~controllable_hmaster2 & ~n12397;
  assign n12399 = ~n12193 & ~n12398;
  assign n12400 = ~controllable_hgrant3 & ~n12399;
  assign n12401 = ~n12163 & ~n12400;
  assign n12402 = controllable_nhgrant0 & ~n12401;
  assign n12403 = ~n12249 & ~n12402;
  assign n12404 = ~n3281 & ~n12403;
  assign n12405 = ~n4089 & ~n12404;
  assign n12406 = n3378 & ~n12405;
  assign n12407 = ~n4015 & ~n6465;
  assign n12408 = ~controllable_hgrant2 & ~n12407;
  assign n12409 = ~n5616 & ~n12408;
  assign n12410 = ~controllable_hmaster0 & ~n12409;
  assign n12411 = ~n6408 & ~n12410;
  assign n12412 = ~controllable_hmaster1 & ~n12411;
  assign n12413 = ~n6407 & ~n12412;
  assign n12414 = i_hbusreq3 & ~n12413;
  assign n12415 = i_hbusreq2 & ~n12407;
  assign n12416 = ~n4064 & ~n6498;
  assign n12417 = ~i_hbusreq2 & ~n12416;
  assign n12418 = ~n12415 & ~n12417;
  assign n12419 = ~controllable_hgrant2 & ~n12418;
  assign n12420 = ~n5862 & ~n12419;
  assign n12421 = ~controllable_hmaster0 & ~n12420;
  assign n12422 = ~n6440 & ~n12421;
  assign n12423 = ~controllable_hmaster1 & ~n12422;
  assign n12424 = ~n6439 & ~n12423;
  assign n12425 = ~i_hbusreq3 & ~n12424;
  assign n12426 = ~n12414 & ~n12425;
  assign n12427 = controllable_hmaster2 & ~n12426;
  assign n12428 = ~n6408 & ~n6471;
  assign n12429 = controllable_hmaster1 & ~n12428;
  assign n12430 = ~n6483 & ~n12429;
  assign n12431 = i_hbusreq3 & ~n12430;
  assign n12432 = ~n5863 & ~n6451;
  assign n12433 = ~i_hbusreq2 & ~n12432;
  assign n12434 = ~n6417 & ~n12433;
  assign n12435 = ~controllable_hgrant2 & ~n12434;
  assign n12436 = ~n5862 & ~n12435;
  assign n12437 = controllable_hmaster0 & ~n12436;
  assign n12438 = ~n6506 & ~n12437;
  assign n12439 = controllable_hmaster1 & ~n12438;
  assign n12440 = ~n6550 & ~n12439;
  assign n12441 = ~i_hbusreq3 & ~n12440;
  assign n12442 = ~n12431 & ~n12441;
  assign n12443 = ~controllable_hmaster2 & ~n12442;
  assign n12444 = ~n12427 & ~n12443;
  assign n12445 = ~controllable_hgrant3 & ~n12444;
  assign n12446 = ~n5861 & ~n12445;
  assign n12447 = controllable_nhgrant0 & ~n12446;
  assign n12448 = ~n6082 & ~n12447;
  assign n12449 = ~n3281 & ~n12448;
  assign n12450 = ~n4089 & ~n12449;
  assign n12451 = ~n3378 & ~n12450;
  assign n12452 = ~n12406 & ~n12451;
  assign n12453 = n3492 & ~n12452;
  assign n12454 = ~n3631 & ~n12453;
  assign n12455 = n3485 & ~n12454;
  assign n12456 = ~n3630 & ~n12455;
  assign n12457 = n3476 & ~n12456;
  assign n12458 = ~n12377 & ~n12457;
  assign n12459 = n3374 & ~n12458;
  assign n12460 = ~n12314 & ~n12459;
  assign n12461 = ~n3655 & ~n12460;
  assign n12462 = ~n12308 & ~n12461;
  assign n12463 = n3652 & ~n12462;
  assign n12464 = ~n6665 & ~n12026;
  assign n12465 = n3492 & ~n12464;
  assign n12466 = ~n3631 & ~n12465;
  assign n12467 = n3485 & ~n12466;
  assign n12468 = ~n3630 & ~n12467;
  assign n12469 = ~n3374 & ~n12468;
  assign n12470 = ~n5291 & ~n9434;
  assign n12471 = controllable_hmaster1 & ~n12470;
  assign n12472 = ~n5305 & ~n12471;
  assign n12473 = i_hbusreq3 & ~n12472;
  assign n12474 = ~n5311 & ~n9447;
  assign n12475 = controllable_hmaster1 & ~n12474;
  assign n12476 = ~n5334 & ~n12475;
  assign n12477 = ~i_hbusreq3 & ~n12476;
  assign n12478 = ~n12473 & ~n12477;
  assign n12479 = ~controllable_hmaster2 & ~n12478;
  assign n12480 = ~n12065 & ~n12479;
  assign n12481 = ~controllable_hgrant3 & ~n12480;
  assign n12482 = ~n12041 & ~n12481;
  assign n12483 = controllable_nhgrant0 & ~n12482;
  assign n12484 = ~n12101 & ~n12483;
  assign n12485 = ~n3281 & ~n12484;
  assign n12486 = ~n3950 & ~n12485;
  assign n12487 = n3378 & ~n12486;
  assign n12488 = ~n4333 & ~n12107;
  assign n12489 = ~controllable_hmaster0 & ~n12488;
  assign n12490 = ~n6682 & ~n12489;
  assign n12491 = ~controllable_hmaster1 & ~n12490;
  assign n12492 = ~n6681 & ~n12491;
  assign n12493 = i_hbusreq3 & ~n12492;
  assign n12494 = ~n4340 & ~n12118;
  assign n12495 = ~controllable_hmaster0 & ~n12494;
  assign n12496 = ~n6689 & ~n12495;
  assign n12497 = ~controllable_hmaster1 & ~n12496;
  assign n12498 = ~n6688 & ~n12497;
  assign n12499 = ~i_hbusreq3 & ~n12498;
  assign n12500 = ~n12493 & ~n12499;
  assign n12501 = controllable_hmaster2 & ~n12500;
  assign n12502 = ~n6699 & ~n9434;
  assign n12503 = controllable_hmaster1 & ~n12502;
  assign n12504 = ~n6706 & ~n12503;
  assign n12505 = i_hbusreq3 & ~n12504;
  assign n12506 = ~n6712 & ~n9447;
  assign n12507 = controllable_hmaster1 & ~n12506;
  assign n12508 = ~n6719 & ~n12507;
  assign n12509 = ~i_hbusreq3 & ~n12508;
  assign n12510 = ~n12505 & ~n12509;
  assign n12511 = ~controllable_hmaster2 & ~n12510;
  assign n12512 = ~n12501 & ~n12511;
  assign n12513 = ~controllable_hgrant3 & ~n12512;
  assign n12514 = ~n5402 & ~n12513;
  assign n12515 = controllable_nhgrant0 & ~n12514;
  assign n12516 = ~n5534 & ~n12515;
  assign n12517 = ~n3281 & ~n12516;
  assign n12518 = ~n3950 & ~n12517;
  assign n12519 = ~n3378 & ~n12518;
  assign n12520 = ~n12487 & ~n12519;
  assign n12521 = n3492 & ~n12520;
  assign n12522 = ~n3631 & ~n12521;
  assign n12523 = n3485 & ~n12522;
  assign n12524 = ~n3630 & ~n12523;
  assign n12525 = ~n3476 & ~n12524;
  assign n12526 = ~n5623 & ~n6738;
  assign n12527 = controllable_hmaster0 & ~n12526;
  assign n12528 = ~n5688 & ~n12527;
  assign n12529 = controllable_hmaster1 & ~n12528;
  assign n12530 = ~n5704 & ~n12529;
  assign n12531 = i_hbusreq3 & ~n12530;
  assign n12532 = ~n6745 & ~n12202;
  assign n12533 = controllable_hmaster0 & ~n12532;
  assign n12534 = ~n12210 & ~n12533;
  assign n12535 = controllable_hmaster1 & ~n12534;
  assign n12536 = ~n12222 & ~n12535;
  assign n12537 = ~i_hbusreq3 & ~n12536;
  assign n12538 = ~n12531 & ~n12537;
  assign n12539 = ~controllable_hmaster2 & ~n12538;
  assign n12540 = ~n12193 & ~n12539;
  assign n12541 = ~controllable_hgrant3 & ~n12540;
  assign n12542 = ~n12163 & ~n12541;
  assign n12543 = controllable_nhgrant0 & ~n12542;
  assign n12544 = ~n12249 & ~n12543;
  assign n12545 = ~n3281 & ~n12544;
  assign n12546 = ~n4089 & ~n12545;
  assign n12547 = n3378 & ~n12546;
  assign n12548 = ~n6762 & ~n12255;
  assign n12549 = ~controllable_hmaster0 & ~n12548;
  assign n12550 = ~n6765 & ~n12549;
  assign n12551 = ~controllable_hmaster1 & ~n12550;
  assign n12552 = ~n6764 & ~n12551;
  assign n12553 = i_hbusreq3 & ~n12552;
  assign n12554 = ~n6772 & ~n12266;
  assign n12555 = ~controllable_hmaster0 & ~n12554;
  assign n12556 = ~n6775 & ~n12555;
  assign n12557 = ~controllable_hmaster1 & ~n12556;
  assign n12558 = ~n6774 & ~n12557;
  assign n12559 = ~i_hbusreq3 & ~n12558;
  assign n12560 = ~n12553 & ~n12559;
  assign n12561 = controllable_hmaster2 & ~n12560;
  assign n12562 = ~n6765 & ~n6788;
  assign n12563 = controllable_hmaster1 & ~n12562;
  assign n12564 = ~n6795 & ~n12563;
  assign n12565 = i_hbusreq3 & ~n12564;
  assign n12566 = ~n6772 & ~n12282;
  assign n12567 = controllable_hmaster0 & ~n12566;
  assign n12568 = ~n6815 & ~n12567;
  assign n12569 = controllable_hmaster1 & ~n12568;
  assign n12570 = ~n6835 & ~n12569;
  assign n12571 = ~i_hbusreq3 & ~n12570;
  assign n12572 = ~n12565 & ~n12571;
  assign n12573 = ~controllable_hmaster2 & ~n12572;
  assign n12574 = ~n12561 & ~n12573;
  assign n12575 = ~controllable_hgrant3 & ~n12574;
  assign n12576 = ~n5861 & ~n12575;
  assign n12577 = controllable_nhgrant0 & ~n12576;
  assign n12578 = ~n6082 & ~n12577;
  assign n12579 = ~n3281 & ~n12578;
  assign n12580 = ~n4089 & ~n12579;
  assign n12581 = ~n3378 & ~n12580;
  assign n12582 = ~n12547 & ~n12581;
  assign n12583 = n3492 & ~n12582;
  assign n12584 = ~n3631 & ~n12583;
  assign n12585 = n3485 & ~n12584;
  assign n12586 = ~n3630 & ~n12585;
  assign n12587 = n3476 & ~n12586;
  assign n12588 = ~n12525 & ~n12587;
  assign n12589 = n3374 & ~n12588;
  assign n12590 = ~n12469 & ~n12589;
  assign n12591 = n3655 & ~n12590;
  assign n12592 = ~n6895 & ~n12026;
  assign n12593 = n3492 & ~n12592;
  assign n12594 = ~n3631 & ~n12593;
  assign n12595 = n3485 & ~n12594;
  assign n12596 = ~n3630 & ~n12595;
  assign n12597 = ~n3374 & ~n12596;
  assign n12598 = ~n5291 & ~n9588;
  assign n12599 = controllable_hmaster1 & ~n12598;
  assign n12600 = ~n5305 & ~n12599;
  assign n12601 = i_hbusreq3 & ~n12600;
  assign n12602 = ~n5311 & ~n9601;
  assign n12603 = controllable_hmaster1 & ~n12602;
  assign n12604 = ~n5334 & ~n12603;
  assign n12605 = ~i_hbusreq3 & ~n12604;
  assign n12606 = ~n12601 & ~n12605;
  assign n12607 = ~controllable_hmaster2 & ~n12606;
  assign n12608 = ~n12065 & ~n12607;
  assign n12609 = ~controllable_hgrant3 & ~n12608;
  assign n12610 = ~n12041 & ~n12609;
  assign n12611 = controllable_nhgrant0 & ~n12610;
  assign n12612 = ~n12101 & ~n12611;
  assign n12613 = ~n3281 & ~n12612;
  assign n12614 = ~n3950 & ~n12613;
  assign n12615 = n3378 & ~n12614;
  assign n12616 = ~n4333 & ~n12334;
  assign n12617 = ~controllable_hmaster0 & ~n12616;
  assign n12618 = ~n6912 & ~n12617;
  assign n12619 = ~controllable_hmaster1 & ~n12618;
  assign n12620 = ~n6911 & ~n12619;
  assign n12621 = i_hbusreq3 & ~n12620;
  assign n12622 = ~n4340 & ~n12345;
  assign n12623 = ~controllable_hmaster0 & ~n12622;
  assign n12624 = ~n6919 & ~n12623;
  assign n12625 = ~controllable_hmaster1 & ~n12624;
  assign n12626 = ~n6918 & ~n12625;
  assign n12627 = ~i_hbusreq3 & ~n12626;
  assign n12628 = ~n12621 & ~n12627;
  assign n12629 = controllable_hmaster2 & ~n12628;
  assign n12630 = ~n6929 & ~n9588;
  assign n12631 = controllable_hmaster1 & ~n12630;
  assign n12632 = ~n6936 & ~n12631;
  assign n12633 = i_hbusreq3 & ~n12632;
  assign n12634 = ~n6942 & ~n9601;
  assign n12635 = controllable_hmaster1 & ~n12634;
  assign n12636 = ~n6951 & ~n12635;
  assign n12637 = ~i_hbusreq3 & ~n12636;
  assign n12638 = ~n12633 & ~n12637;
  assign n12639 = ~controllable_hmaster2 & ~n12638;
  assign n12640 = ~n12629 & ~n12639;
  assign n12641 = ~controllable_hgrant3 & ~n12640;
  assign n12642 = ~n5402 & ~n12641;
  assign n12643 = controllable_nhgrant0 & ~n12642;
  assign n12644 = ~n5534 & ~n12643;
  assign n12645 = ~n3281 & ~n12644;
  assign n12646 = ~n3950 & ~n12645;
  assign n12647 = ~n3378 & ~n12646;
  assign n12648 = ~n12615 & ~n12647;
  assign n12649 = n3492 & ~n12648;
  assign n12650 = ~n3631 & ~n12649;
  assign n12651 = n3485 & ~n12650;
  assign n12652 = ~n3630 & ~n12651;
  assign n12653 = ~n3476 & ~n12652;
  assign n12654 = ~n6738 & ~n12379;
  assign n12655 = controllable_hmaster0 & ~n12654;
  assign n12656 = ~n5688 & ~n12655;
  assign n12657 = controllable_hmaster1 & ~n12656;
  assign n12658 = ~n5704 & ~n12657;
  assign n12659 = i_hbusreq3 & ~n12658;
  assign n12660 = ~n6745 & ~n12390;
  assign n12661 = controllable_hmaster0 & ~n12660;
  assign n12662 = ~n12210 & ~n12661;
  assign n12663 = controllable_hmaster1 & ~n12662;
  assign n12664 = ~n12222 & ~n12663;
  assign n12665 = ~i_hbusreq3 & ~n12664;
  assign n12666 = ~n12659 & ~n12665;
  assign n12667 = ~controllable_hmaster2 & ~n12666;
  assign n12668 = ~n12193 & ~n12667;
  assign n12669 = ~controllable_hgrant3 & ~n12668;
  assign n12670 = ~n12163 & ~n12669;
  assign n12671 = controllable_nhgrant0 & ~n12670;
  assign n12672 = ~n12249 & ~n12671;
  assign n12673 = ~n3281 & ~n12672;
  assign n12674 = ~n4089 & ~n12673;
  assign n12675 = n3378 & ~n12674;
  assign n12676 = ~n6762 & ~n12408;
  assign n12677 = ~controllable_hmaster0 & ~n12676;
  assign n12678 = ~n6994 & ~n12677;
  assign n12679 = ~controllable_hmaster1 & ~n12678;
  assign n12680 = ~n6993 & ~n12679;
  assign n12681 = i_hbusreq3 & ~n12680;
  assign n12682 = ~n6772 & ~n12419;
  assign n12683 = ~controllable_hmaster0 & ~n12682;
  assign n12684 = ~n7003 & ~n12683;
  assign n12685 = ~controllable_hmaster1 & ~n12684;
  assign n12686 = ~n7002 & ~n12685;
  assign n12687 = ~i_hbusreq3 & ~n12686;
  assign n12688 = ~n12681 & ~n12687;
  assign n12689 = controllable_hmaster2 & ~n12688;
  assign n12690 = ~n6994 & ~n7015;
  assign n12691 = controllable_hmaster1 & ~n12690;
  assign n12692 = ~n7022 & ~n12691;
  assign n12693 = i_hbusreq3 & ~n12692;
  assign n12694 = ~n6772 & ~n12435;
  assign n12695 = controllable_hmaster0 & ~n12694;
  assign n12696 = ~n7028 & ~n12695;
  assign n12697 = controllable_hmaster1 & ~n12696;
  assign n12698 = ~n7036 & ~n12697;
  assign n12699 = ~i_hbusreq3 & ~n12698;
  assign n12700 = ~n12693 & ~n12699;
  assign n12701 = ~controllable_hmaster2 & ~n12700;
  assign n12702 = ~n12689 & ~n12701;
  assign n12703 = ~controllable_hgrant3 & ~n12702;
  assign n12704 = ~n5861 & ~n12703;
  assign n12705 = controllable_nhgrant0 & ~n12704;
  assign n12706 = ~n6082 & ~n12705;
  assign n12707 = ~n3281 & ~n12706;
  assign n12708 = ~n4089 & ~n12707;
  assign n12709 = ~n3378 & ~n12708;
  assign n12710 = ~n12675 & ~n12709;
  assign n12711 = n3492 & ~n12710;
  assign n12712 = ~n3631 & ~n12711;
  assign n12713 = n3485 & ~n12712;
  assign n12714 = ~n3630 & ~n12713;
  assign n12715 = n3476 & ~n12714;
  assign n12716 = ~n12653 & ~n12715;
  assign n12717 = n3374 & ~n12716;
  assign n12718 = ~n12597 & ~n12717;
  assign n12719 = ~n3655 & ~n12718;
  assign n12720 = ~n12591 & ~n12719;
  assign n12721 = ~n3652 & ~n12720;
  assign n12722 = ~n12463 & ~n12721;
  assign n12723 = ~n3368 & ~n12722;
  assign n12724 = ~n5278 & ~n9780;
  assign n12725 = controllable_hmaster1 & ~n12724;
  assign n12726 = ~n5281 & ~n12725;
  assign n12727 = ~i_hbusreq3 & ~n12726;
  assign n12728 = ~n5265 & ~n12727;
  assign n12729 = ~controllable_hmaster2 & ~n12728;
  assign n12730 = ~n12033 & ~n12729;
  assign n12731 = controllable_hgrant3 & ~n12730;
  assign n12732 = ~n5260 & ~n12046;
  assign n12733 = ~controllable_hmaster1 & ~n12732;
  assign n12734 = ~n7063 & ~n12733;
  assign n12735 = i_hbusreq3 & ~n12734;
  assign n12736 = ~n5277 & ~n12059;
  assign n12737 = ~controllable_hmaster1 & ~n12736;
  assign n12738 = ~n7068 & ~n12737;
  assign n12739 = ~i_hbusreq3 & ~n12738;
  assign n12740 = ~n12735 & ~n12739;
  assign n12741 = controllable_hmaster2 & ~n12740;
  assign n12742 = ~n5311 & ~n9802;
  assign n12743 = controllable_hmaster1 & ~n12742;
  assign n12744 = ~n5334 & ~n12743;
  assign n12745 = ~i_hbusreq3 & ~n12744;
  assign n12746 = ~n12069 & ~n12745;
  assign n12747 = ~controllable_hmaster2 & ~n12746;
  assign n12748 = ~n12741 & ~n12747;
  assign n12749 = ~controllable_hgrant3 & ~n12748;
  assign n12750 = ~n12731 & ~n12749;
  assign n12751 = controllable_nhgrant0 & ~n12750;
  assign n12752 = ~n5278 & ~n9700;
  assign n12753 = controllable_hmaster1 & ~n12752;
  assign n12754 = ~n5281 & ~n12753;
  assign n12755 = ~i_hbusreq3 & ~n12754;
  assign n12756 = ~n3951 & ~n12755;
  assign n12757 = ~controllable_hmaster2 & ~n12756;
  assign n12758 = ~n12033 & ~n12757;
  assign n12759 = controllable_hgrant3 & ~n12758;
  assign n12760 = ~n3821 & ~n9737;
  assign n12761 = controllable_hmaster1 & ~n12760;
  assign n12762 = ~n5350 & ~n12761;
  assign n12763 = i_hbusreq3 & ~n12762;
  assign n12764 = ~n5278 & ~n9743;
  assign n12765 = controllable_hmaster1 & ~n12764;
  assign n12766 = ~n5355 & ~n12765;
  assign n12767 = ~i_hbusreq3 & ~n12766;
  assign n12768 = ~n12763 & ~n12767;
  assign n12769 = ~controllable_hmaster2 & ~n12768;
  assign n12770 = ~n12033 & ~n12769;
  assign n12771 = ~controllable_hgrant3 & ~n12770;
  assign n12772 = ~n12759 & ~n12771;
  assign n12773 = ~controllable_nhgrant0 & ~n12772;
  assign n12774 = ~n12751 & ~n12773;
  assign n12775 = ~n3281 & ~n12774;
  assign n12776 = ~n3281 & ~n12775;
  assign n12777 = n3378 & ~n12776;
  assign n12778 = ~n3835 & ~n9780;
  assign n12779 = controllable_hmaster1 & ~n12778;
  assign n12780 = ~n5396 & ~n12779;
  assign n12781 = ~i_hbusreq3 & ~n12780;
  assign n12782 = ~n5265 & ~n12781;
  assign n12783 = ~controllable_hmaster2 & ~n12782;
  assign n12784 = ~n5370 & ~n12783;
  assign n12785 = controllable_hgrant3 & ~n12784;
  assign n12786 = ~n5046 & ~n12109;
  assign n12787 = ~controllable_hmaster1 & ~n12786;
  assign n12788 = ~n5045 & ~n12787;
  assign n12789 = i_hbusreq3 & ~n12788;
  assign n12790 = ~n5071 & ~n12120;
  assign n12791 = ~controllable_hmaster1 & ~n12790;
  assign n12792 = ~n5070 & ~n12791;
  assign n12793 = ~i_hbusreq3 & ~n12792;
  assign n12794 = ~n12789 & ~n12793;
  assign n12795 = controllable_hmaster2 & ~n12794;
  assign n12796 = ~n5440 & ~n9802;
  assign n12797 = controllable_hmaster1 & ~n12796;
  assign n12798 = ~n5480 & ~n12797;
  assign n12799 = ~i_hbusreq3 & ~n12798;
  assign n12800 = ~n12130 & ~n12799;
  assign n12801 = ~controllable_hmaster2 & ~n12800;
  assign n12802 = ~n12795 & ~n12801;
  assign n12803 = ~controllable_hgrant3 & ~n12802;
  assign n12804 = ~n12785 & ~n12803;
  assign n12805 = controllable_nhgrant0 & ~n12804;
  assign n12806 = ~n3835 & ~n9700;
  assign n12807 = controllable_hmaster1 & ~n12806;
  assign n12808 = ~n5396 & ~n12807;
  assign n12809 = ~i_hbusreq3 & ~n12808;
  assign n12810 = ~n3951 & ~n12809;
  assign n12811 = ~controllable_hmaster2 & ~n12810;
  assign n12812 = ~n5370 & ~n12811;
  assign n12813 = controllable_hgrant3 & ~n12812;
  assign n12814 = ~n3910 & ~n9737;
  assign n12815 = controllable_hmaster1 & ~n12814;
  assign n12816 = ~n5501 & ~n12815;
  assign n12817 = i_hbusreq3 & ~n12816;
  assign n12818 = ~n3935 & ~n9743;
  assign n12819 = controllable_hmaster1 & ~n12818;
  assign n12820 = ~n5526 & ~n12819;
  assign n12821 = ~i_hbusreq3 & ~n12820;
  assign n12822 = ~n12817 & ~n12821;
  assign n12823 = ~controllable_hmaster2 & ~n12822;
  assign n12824 = ~n5498 & ~n12823;
  assign n12825 = ~controllable_hgrant3 & ~n12824;
  assign n12826 = ~n12813 & ~n12825;
  assign n12827 = ~controllable_nhgrant0 & ~n12826;
  assign n12828 = ~n12805 & ~n12827;
  assign n12829 = ~n3281 & ~n12828;
  assign n12830 = ~n3281 & ~n12829;
  assign n12831 = ~n3378 & ~n12830;
  assign n12832 = ~n12777 & ~n12831;
  assign n12833 = n3492 & ~n12832;
  assign n12834 = n3492 & ~n12833;
  assign n12835 = n3485 & ~n12834;
  assign n12836 = n3485 & ~n12835;
  assign n12837 = ~n3476 & ~n12836;
  assign n12838 = ~controllable_hgrant4 & ~n7268;
  assign n12839 = ~n3433 & ~n12838;
  assign n12840 = ~i_hbusreq2 & ~n12839;
  assign n12841 = ~n5550 & ~n12840;
  assign n12842 = ~controllable_hgrant2 & ~n12841;
  assign n12843 = ~n3431 & ~n12842;
  assign n12844 = ~i_hbusreq3 & ~n12843;
  assign n12845 = ~n5549 & ~n12844;
  assign n12846 = controllable_hmaster2 & ~n12845;
  assign n12847 = ~controllable_hmaster0 & ~n12843;
  assign n12848 = ~n10098 & ~n12847;
  assign n12849 = controllable_hmaster1 & ~n12848;
  assign n12850 = ~controllable_hmaster1 & ~n12843;
  assign n12851 = ~n12849 & ~n12850;
  assign n12852 = ~i_hbusreq3 & ~n12851;
  assign n12853 = ~n5593 & ~n12852;
  assign n12854 = ~controllable_hmaster2 & ~n12853;
  assign n12855 = ~n12846 & ~n12854;
  assign n12856 = controllable_hgrant3 & ~n12855;
  assign n12857 = ~n4015 & ~n7322;
  assign n12858 = ~controllable_hgrant2 & ~n12857;
  assign n12859 = ~n5616 & ~n12858;
  assign n12860 = ~controllable_hmaster0 & ~n12859;
  assign n12861 = ~n7250 & ~n12860;
  assign n12862 = ~controllable_hmaster1 & ~n12861;
  assign n12863 = ~n7249 & ~n12862;
  assign n12864 = i_hbusreq3 & ~n12863;
  assign n12865 = ~n7282 & ~n12172;
  assign n12866 = ~i_hbusreq2 & ~n12865;
  assign n12867 = ~n7264 & ~n12866;
  assign n12868 = ~controllable_hgrant2 & ~n12867;
  assign n12869 = ~n5635 & ~n12868;
  assign n12870 = controllable_hmaster1 & ~n12869;
  assign n12871 = controllable_hmaster0 & ~n12869;
  assign n12872 = i_hbusreq2 & ~n12857;
  assign n12873 = ~n7353 & ~n12181;
  assign n12874 = ~i_hbusreq2 & ~n12873;
  assign n12875 = ~n12872 & ~n12874;
  assign n12876 = ~controllable_hgrant2 & ~n12875;
  assign n12877 = ~n5635 & ~n12876;
  assign n12878 = ~controllable_hmaster0 & ~n12877;
  assign n12879 = ~n12871 & ~n12878;
  assign n12880 = ~controllable_hmaster1 & ~n12879;
  assign n12881 = ~n12870 & ~n12880;
  assign n12882 = ~i_hbusreq3 & ~n12881;
  assign n12883 = ~n12864 & ~n12882;
  assign n12884 = controllable_hmaster2 & ~n12883;
  assign n12885 = ~n4091 & ~n7255;
  assign n12886 = ~controllable_hgrant2 & ~n12885;
  assign n12887 = ~n5616 & ~n12886;
  assign n12888 = controllable_hmaster0 & ~n12887;
  assign n12889 = ~n7328 & ~n12888;
  assign n12890 = controllable_hmaster1 & ~n12889;
  assign n12891 = ~n7342 & ~n12890;
  assign n12892 = i_hbusreq3 & ~n12891;
  assign n12893 = i_hbusreq2 & ~n12885;
  assign n12894 = controllable_hgrant4 & ~n7225;
  assign n12895 = ~n7308 & ~n12894;
  assign n12896 = ~i_hbusreq2 & ~n12895;
  assign n12897 = ~n12893 & ~n12896;
  assign n12898 = ~controllable_hgrant2 & ~n12897;
  assign n12899 = ~n7290 & ~n12898;
  assign n12900 = controllable_hmaster0 & ~n12899;
  assign n12901 = ~n7353 & ~n12172;
  assign n12902 = ~i_hbusreq2 & ~n12901;
  assign n12903 = ~n7345 & ~n12902;
  assign n12904 = ~controllable_hgrant2 & ~n12903;
  assign n12905 = ~n5722 & ~n12904;
  assign n12906 = ~controllable_hmaster0 & ~n12905;
  assign n12907 = ~n12900 & ~n12906;
  assign n12908 = controllable_hmaster1 & ~n12907;
  assign n12909 = ~n7376 & ~n12172;
  assign n12910 = ~i_hbusreq2 & ~n12909;
  assign n12911 = ~n7364 & ~n12910;
  assign n12912 = ~controllable_hgrant2 & ~n12911;
  assign n12913 = ~n5635 & ~n12912;
  assign n12914 = controllable_hmaster0 & ~n12913;
  assign n12915 = ~n5635 & ~n12904;
  assign n12916 = ~controllable_hmaster0 & ~n12915;
  assign n12917 = ~n12914 & ~n12916;
  assign n12918 = ~controllable_hmaster1 & ~n12917;
  assign n12919 = ~n12908 & ~n12918;
  assign n12920 = ~i_hbusreq3 & ~n12919;
  assign n12921 = ~n12892 & ~n12920;
  assign n12922 = ~controllable_hmaster2 & ~n12921;
  assign n12923 = ~n12884 & ~n12922;
  assign n12924 = ~controllable_hgrant3 & ~n12923;
  assign n12925 = ~n12856 & ~n12924;
  assign n12926 = controllable_nhgrant0 & ~n12925;
  assign n12927 = controllable_hmaster0 & ~n7398;
  assign n12928 = ~n5588 & ~n12927;
  assign n12929 = controllable_hmaster1 & ~n12928;
  assign n12930 = ~n5796 & ~n12929;
  assign n12931 = i_hbusreq3 & ~n12930;
  assign n12932 = controllable_hmaster0 & ~n7421;
  assign n12933 = ~n5606 & ~n12932;
  assign n12934 = controllable_hmaster1 & ~n12933;
  assign n12935 = ~n5801 & ~n12934;
  assign n12936 = ~i_hbusreq3 & ~n12935;
  assign n12937 = ~n12931 & ~n12936;
  assign n12938 = ~controllable_hmaster2 & ~n12937;
  assign n12939 = ~n12233 & ~n12938;
  assign n12940 = ~controllable_hgrant3 & ~n12939;
  assign n12941 = ~n12759 & ~n12940;
  assign n12942 = ~controllable_nhgrant0 & ~n12941;
  assign n12943 = ~n12926 & ~n12942;
  assign n12944 = ~n3281 & ~n12943;
  assign n12945 = ~n3281 & ~n12944;
  assign n12946 = n3378 & ~n12945;
  assign n12947 = ~controllable_hgrant4 & ~n7485;
  assign n12948 = ~n3916 & ~n12947;
  assign n12949 = ~i_hbusreq2 & ~n12948;
  assign n12950 = ~n5550 & ~n12949;
  assign n12951 = ~controllable_hgrant2 & ~n12950;
  assign n12952 = ~n3859 & ~n12951;
  assign n12953 = ~i_hbusreq3 & ~n12952;
  assign n12954 = ~n5549 & ~n12953;
  assign n12955 = controllable_hmaster2 & ~n12954;
  assign n12956 = ~controllable_hmaster0 & ~n12952;
  assign n12957 = ~n10098 & ~n12956;
  assign n12958 = controllable_hmaster1 & ~n12957;
  assign n12959 = controllable_hmaster0 & ~n12952;
  assign n12960 = ~controllable_hgrant4 & ~n7605;
  assign n12961 = ~n5462 & ~n12960;
  assign n12962 = ~i_hbusreq2 & ~n12961;
  assign n12963 = ~n5550 & ~n12962;
  assign n12964 = ~controllable_hgrant2 & ~n12963;
  assign n12965 = ~n5461 & ~n12964;
  assign n12966 = ~controllable_hmaster0 & ~n12965;
  assign n12967 = ~n12959 & ~n12966;
  assign n12968 = ~controllable_hmaster1 & ~n12967;
  assign n12969 = ~n12958 & ~n12968;
  assign n12970 = ~i_hbusreq3 & ~n12969;
  assign n12971 = ~n5593 & ~n12970;
  assign n12972 = ~controllable_hmaster2 & ~n12971;
  assign n12973 = ~n12955 & ~n12972;
  assign n12974 = controllable_hgrant3 & ~n12973;
  assign n12975 = ~n4015 & ~n7535;
  assign n12976 = ~controllable_hgrant2 & ~n12975;
  assign n12977 = ~n5616 & ~n12976;
  assign n12978 = ~controllable_hmaster0 & ~n12977;
  assign n12979 = ~n7466 & ~n12978;
  assign n12980 = ~controllable_hmaster1 & ~n12979;
  assign n12981 = ~n7465 & ~n12980;
  assign n12982 = i_hbusreq3 & ~n12981;
  assign n12983 = ~n5863 & ~n7499;
  assign n12984 = ~i_hbusreq2 & ~n12983;
  assign n12985 = ~n7479 & ~n12984;
  assign n12986 = ~controllable_hgrant2 & ~n12985;
  assign n12987 = ~n5862 & ~n12986;
  assign n12988 = controllable_hmaster1 & ~n12987;
  assign n12989 = controllable_hmaster0 & ~n12987;
  assign n12990 = i_hbusreq2 & ~n12975;
  assign n12991 = ~n4064 & ~n7568;
  assign n12992 = ~i_hbusreq2 & ~n12991;
  assign n12993 = ~n12990 & ~n12992;
  assign n12994 = ~controllable_hgrant2 & ~n12993;
  assign n12995 = ~n5862 & ~n12994;
  assign n12996 = ~controllable_hmaster0 & ~n12995;
  assign n12997 = ~n12989 & ~n12996;
  assign n12998 = ~controllable_hmaster1 & ~n12997;
  assign n12999 = ~n12988 & ~n12998;
  assign n13000 = ~i_hbusreq3 & ~n12999;
  assign n13001 = ~n12982 & ~n13000;
  assign n13002 = controllable_hmaster2 & ~n13001;
  assign n13003 = ~n4091 & ~n7470;
  assign n13004 = ~controllable_hgrant2 & ~n13003;
  assign n13005 = ~n5616 & ~n13004;
  assign n13006 = controllable_hmaster0 & ~n13005;
  assign n13007 = ~n7541 & ~n13006;
  assign n13008 = controllable_hmaster1 & ~n13007;
  assign n13009 = ~n7554 & ~n13008;
  assign n13010 = i_hbusreq3 & ~n13009;
  assign n13011 = i_hbusreq2 & ~n13003;
  assign n13012 = controllable_hgrant4 & ~n7442;
  assign n13013 = ~n7521 & ~n13012;
  assign n13014 = ~i_hbusreq2 & ~n13013;
  assign n13015 = ~n13011 & ~n13014;
  assign n13016 = ~controllable_hgrant2 & ~n13015;
  assign n13017 = ~n7507 & ~n13016;
  assign n13018 = controllable_hmaster0 & ~n13017;
  assign n13019 = ~n5863 & ~n7568;
  assign n13020 = ~i_hbusreq2 & ~n13019;
  assign n13021 = ~n7557 & ~n13020;
  assign n13022 = ~controllable_hgrant2 & ~n13021;
  assign n13023 = ~n5950 & ~n13022;
  assign n13024 = ~controllable_hmaster0 & ~n13023;
  assign n13025 = ~n13018 & ~n13024;
  assign n13026 = controllable_hmaster1 & ~n13025;
  assign n13027 = ~n5863 & ~n7592;
  assign n13028 = ~i_hbusreq2 & ~n13027;
  assign n13029 = ~n7579 & ~n13028;
  assign n13030 = ~controllable_hgrant2 & ~n13029;
  assign n13031 = ~n5862 & ~n13030;
  assign n13032 = controllable_hmaster0 & ~n13031;
  assign n13033 = ~n5982 & ~n7614;
  assign n13034 = ~i_hbusreq2 & ~n13033;
  assign n13035 = ~n7557 & ~n13034;
  assign n13036 = ~controllable_hgrant2 & ~n13035;
  assign n13037 = ~n5981 & ~n13036;
  assign n13038 = ~controllable_hmaster0 & ~n13037;
  assign n13039 = ~n13032 & ~n13038;
  assign n13040 = ~controllable_hmaster1 & ~n13039;
  assign n13041 = ~n13026 & ~n13040;
  assign n13042 = ~i_hbusreq3 & ~n13041;
  assign n13043 = ~n13010 & ~n13042;
  assign n13044 = ~controllable_hmaster2 & ~n13043;
  assign n13045 = ~n13002 & ~n13044;
  assign n13046 = ~controllable_hgrant3 & ~n13045;
  assign n13047 = ~n12974 & ~n13046;
  assign n13048 = controllable_nhgrant0 & ~n13047;
  assign n13049 = controllable_hmaster0 & ~n7635;
  assign n13050 = ~n9062 & ~n13049;
  assign n13051 = controllable_hmaster1 & ~n13050;
  assign n13052 = ~n6046 & ~n13051;
  assign n13053 = i_hbusreq3 & ~n13052;
  assign n13054 = controllable_hmaster0 & ~n7657;
  assign n13055 = ~n9086 & ~n13054;
  assign n13056 = controllable_hmaster1 & ~n13055;
  assign n13057 = ~n6074 & ~n13056;
  assign n13058 = ~i_hbusreq3 & ~n13057;
  assign n13059 = ~n13053 & ~n13058;
  assign n13060 = ~controllable_hmaster2 & ~n13059;
  assign n13061 = ~n6035 & ~n13060;
  assign n13062 = ~controllable_hgrant3 & ~n13061;
  assign n13063 = ~n12813 & ~n13062;
  assign n13064 = ~controllable_nhgrant0 & ~n13063;
  assign n13065 = ~n13048 & ~n13064;
  assign n13066 = ~n3281 & ~n13065;
  assign n13067 = ~n3281 & ~n13066;
  assign n13068 = ~n3378 & ~n13067;
  assign n13069 = ~n12946 & ~n13068;
  assign n13070 = n3492 & ~n13069;
  assign n13071 = n3492 & ~n13070;
  assign n13072 = n3485 & ~n13071;
  assign n13073 = n3485 & ~n13072;
  assign n13074 = n3476 & ~n13073;
  assign n13075 = ~n12837 & ~n13074;
  assign n13076 = n3374 & ~n13075;
  assign n13077 = ~n7128 & ~n13076;
  assign n13078 = n3655 & ~n13077;
  assign n13079 = ~n5291 & ~n10326;
  assign n13080 = controllable_hmaster1 & ~n13079;
  assign n13081 = ~n5305 & ~n13080;
  assign n13082 = i_hbusreq3 & ~n13081;
  assign n13083 = ~n5311 & ~n10348;
  assign n13084 = controllable_hmaster1 & ~n13083;
  assign n13085 = ~n5334 & ~n13084;
  assign n13086 = ~i_hbusreq3 & ~n13085;
  assign n13087 = ~n13082 & ~n13086;
  assign n13088 = ~controllable_hmaster2 & ~n13087;
  assign n13089 = ~n12741 & ~n13088;
  assign n13090 = ~controllable_hgrant3 & ~n13089;
  assign n13091 = ~n12731 & ~n13090;
  assign n13092 = controllable_nhgrant0 & ~n13091;
  assign n13093 = ~n12773 & ~n13092;
  assign n13094 = ~n3281 & ~n13093;
  assign n13095 = ~n3281 & ~n13094;
  assign n13096 = n3378 & ~n13095;
  assign n13097 = ~n6105 & ~n12336;
  assign n13098 = ~controllable_hmaster1 & ~n13097;
  assign n13099 = ~n6104 & ~n13098;
  assign n13100 = i_hbusreq3 & ~n13099;
  assign n13101 = ~n6130 & ~n12347;
  assign n13102 = ~controllable_hmaster1 & ~n13101;
  assign n13103 = ~n6129 & ~n13102;
  assign n13104 = ~i_hbusreq3 & ~n13103;
  assign n13105 = ~n13100 & ~n13104;
  assign n13106 = controllable_hmaster2 & ~n13105;
  assign n13107 = ~n6256 & ~n10326;
  assign n13108 = controllable_hmaster1 & ~n13107;
  assign n13109 = ~n6271 & ~n13108;
  assign n13110 = i_hbusreq3 & ~n13109;
  assign n13111 = ~n6295 & ~n10348;
  assign n13112 = controllable_hmaster1 & ~n13111;
  assign n13113 = ~n6339 & ~n13112;
  assign n13114 = ~i_hbusreq3 & ~n13113;
  assign n13115 = ~n13110 & ~n13114;
  assign n13116 = ~controllable_hmaster2 & ~n13115;
  assign n13117 = ~n13106 & ~n13116;
  assign n13118 = ~controllable_hgrant3 & ~n13117;
  assign n13119 = ~n12785 & ~n13118;
  assign n13120 = controllable_nhgrant0 & ~n13119;
  assign n13121 = ~n12827 & ~n13120;
  assign n13122 = ~n3281 & ~n13121;
  assign n13123 = ~n3281 & ~n13122;
  assign n13124 = ~n3378 & ~n13123;
  assign n13125 = ~n13096 & ~n13124;
  assign n13126 = n3492 & ~n13125;
  assign n13127 = n3492 & ~n13126;
  assign n13128 = n3485 & ~n13127;
  assign n13129 = n3485 & ~n13128;
  assign n13130 = ~n3476 & ~n13129;
  assign n13131 = ~n4091 & ~n7750;
  assign n13132 = ~controllable_hgrant2 & ~n13131;
  assign n13133 = ~n5616 & ~n13132;
  assign n13134 = controllable_hmaster0 & ~n13133;
  assign n13135 = ~n7328 & ~n13134;
  assign n13136 = controllable_hmaster1 & ~n13135;
  assign n13137 = ~n7342 & ~n13136;
  assign n13138 = i_hbusreq3 & ~n13137;
  assign n13139 = i_hbusreq2 & ~n13131;
  assign n13140 = ~n7771 & ~n12894;
  assign n13141 = ~i_hbusreq2 & ~n13140;
  assign n13142 = ~n13139 & ~n13141;
  assign n13143 = ~controllable_hgrant2 & ~n13142;
  assign n13144 = ~n7290 & ~n13143;
  assign n13145 = controllable_hmaster0 & ~n13144;
  assign n13146 = ~n12906 & ~n13145;
  assign n13147 = controllable_hmaster1 & ~n13146;
  assign n13148 = ~n12918 & ~n13147;
  assign n13149 = ~i_hbusreq3 & ~n13148;
  assign n13150 = ~n13138 & ~n13149;
  assign n13151 = ~controllable_hmaster2 & ~n13150;
  assign n13152 = ~n12884 & ~n13151;
  assign n13153 = ~controllable_hgrant3 & ~n13152;
  assign n13154 = ~n12856 & ~n13153;
  assign n13155 = controllable_nhgrant0 & ~n13154;
  assign n13156 = ~n12942 & ~n13155;
  assign n13157 = ~n3281 & ~n13156;
  assign n13158 = ~n3281 & ~n13157;
  assign n13159 = n3378 & ~n13158;
  assign n13160 = ~n4015 & ~n7859;
  assign n13161 = ~controllable_hgrant2 & ~n13160;
  assign n13162 = ~n5616 & ~n13161;
  assign n13163 = ~controllable_hmaster0 & ~n13162;
  assign n13164 = ~n7799 & ~n13163;
  assign n13165 = ~controllable_hmaster1 & ~n13164;
  assign n13166 = ~n7798 & ~n13165;
  assign n13167 = i_hbusreq3 & ~n13166;
  assign n13168 = ~n5863 & ~n7824;
  assign n13169 = ~i_hbusreq2 & ~n13168;
  assign n13170 = ~n7811 & ~n13169;
  assign n13171 = ~controllable_hgrant2 & ~n13170;
  assign n13172 = ~n5862 & ~n13171;
  assign n13173 = controllable_hmaster1 & ~n13172;
  assign n13174 = controllable_hmaster0 & ~n13172;
  assign n13175 = i_hbusreq2 & ~n13160;
  assign n13176 = ~n4064 & ~n7891;
  assign n13177 = ~i_hbusreq2 & ~n13176;
  assign n13178 = ~n13175 & ~n13177;
  assign n13179 = ~controllable_hgrant2 & ~n13178;
  assign n13180 = ~n5862 & ~n13179;
  assign n13181 = ~controllable_hmaster0 & ~n13180;
  assign n13182 = ~n13174 & ~n13181;
  assign n13183 = ~controllable_hmaster1 & ~n13182;
  assign n13184 = ~n13173 & ~n13183;
  assign n13185 = ~i_hbusreq3 & ~n13184;
  assign n13186 = ~n13167 & ~n13185;
  assign n13187 = controllable_hmaster2 & ~n13186;
  assign n13188 = ~n4091 & ~n7802;
  assign n13189 = ~controllable_hgrant2 & ~n13188;
  assign n13190 = ~n5616 & ~n13189;
  assign n13191 = controllable_hmaster0 & ~n13190;
  assign n13192 = ~n7865 & ~n13191;
  assign n13193 = controllable_hmaster1 & ~n13192;
  assign n13194 = ~n7877 & ~n13193;
  assign n13195 = i_hbusreq3 & ~n13194;
  assign n13196 = i_hbusreq2 & ~n13188;
  assign n13197 = ~n7845 & ~n13012;
  assign n13198 = ~i_hbusreq2 & ~n13197;
  assign n13199 = ~n13196 & ~n13198;
  assign n13200 = ~controllable_hgrant2 & ~n13199;
  assign n13201 = ~n7507 & ~n13200;
  assign n13202 = controllable_hmaster0 & ~n13201;
  assign n13203 = ~n5863 & ~n7891;
  assign n13204 = ~i_hbusreq2 & ~n13203;
  assign n13205 = ~n7880 & ~n13204;
  assign n13206 = ~controllable_hgrant2 & ~n13205;
  assign n13207 = ~n5950 & ~n13206;
  assign n13208 = ~controllable_hmaster0 & ~n13207;
  assign n13209 = ~n13202 & ~n13208;
  assign n13210 = controllable_hmaster1 & ~n13209;
  assign n13211 = ~n5863 & ~n7916;
  assign n13212 = ~i_hbusreq2 & ~n13211;
  assign n13213 = ~n7902 & ~n13212;
  assign n13214 = ~controllable_hgrant2 & ~n13213;
  assign n13215 = ~n5862 & ~n13214;
  assign n13216 = controllable_hmaster0 & ~n13215;
  assign n13217 = ~n5982 & ~n7930;
  assign n13218 = ~i_hbusreq2 & ~n13217;
  assign n13219 = ~n7880 & ~n13218;
  assign n13220 = ~controllable_hgrant2 & ~n13219;
  assign n13221 = ~n5981 & ~n13220;
  assign n13222 = ~controllable_hmaster0 & ~n13221;
  assign n13223 = ~n13216 & ~n13222;
  assign n13224 = ~controllable_hmaster1 & ~n13223;
  assign n13225 = ~n13210 & ~n13224;
  assign n13226 = ~i_hbusreq3 & ~n13225;
  assign n13227 = ~n13195 & ~n13226;
  assign n13228 = ~controllable_hmaster2 & ~n13227;
  assign n13229 = ~n13187 & ~n13228;
  assign n13230 = ~controllable_hgrant3 & ~n13229;
  assign n13231 = ~n12974 & ~n13230;
  assign n13232 = controllable_nhgrant0 & ~n13231;
  assign n13233 = ~n13064 & ~n13232;
  assign n13234 = ~n3281 & ~n13233;
  assign n13235 = ~n3281 & ~n13234;
  assign n13236 = ~n3378 & ~n13235;
  assign n13237 = ~n13159 & ~n13236;
  assign n13238 = n3492 & ~n13237;
  assign n13239 = n3492 & ~n13238;
  assign n13240 = n3485 & ~n13239;
  assign n13241 = n3485 & ~n13240;
  assign n13242 = n3476 & ~n13241;
  assign n13243 = ~n13130 & ~n13242;
  assign n13244 = n3374 & ~n13243;
  assign n13245 = ~n7706 & ~n13244;
  assign n13246 = ~n3655 & ~n13245;
  assign n13247 = ~n13078 & ~n13246;
  assign n13248 = n3652 & ~n13247;
  assign n13249 = ~n5291 & ~n10767;
  assign n13250 = controllable_hmaster1 & ~n13249;
  assign n13251 = ~n5305 & ~n13250;
  assign n13252 = i_hbusreq3 & ~n13251;
  assign n13253 = ~n5311 & ~n10781;
  assign n13254 = controllable_hmaster1 & ~n13253;
  assign n13255 = ~n5334 & ~n13254;
  assign n13256 = ~i_hbusreq3 & ~n13255;
  assign n13257 = ~n13252 & ~n13256;
  assign n13258 = ~controllable_hmaster2 & ~n13257;
  assign n13259 = ~n12741 & ~n13258;
  assign n13260 = ~controllable_hgrant3 & ~n13259;
  assign n13261 = ~n12731 & ~n13260;
  assign n13262 = controllable_nhgrant0 & ~n13261;
  assign n13263 = ~n12773 & ~n13262;
  assign n13264 = ~n3281 & ~n13263;
  assign n13265 = ~n3281 & ~n13264;
  assign n13266 = n3378 & ~n13265;
  assign n13267 = ~n6577 & ~n12489;
  assign n13268 = ~controllable_hmaster1 & ~n13267;
  assign n13269 = ~n6576 & ~n13268;
  assign n13270 = i_hbusreq3 & ~n13269;
  assign n13271 = ~n6584 & ~n12495;
  assign n13272 = ~controllable_hmaster1 & ~n13271;
  assign n13273 = ~n6583 & ~n13272;
  assign n13274 = ~i_hbusreq3 & ~n13273;
  assign n13275 = ~n13270 & ~n13274;
  assign n13276 = controllable_hmaster2 & ~n13275;
  assign n13277 = ~n6699 & ~n10767;
  assign n13278 = controllable_hmaster1 & ~n13277;
  assign n13279 = ~n6706 & ~n13278;
  assign n13280 = i_hbusreq3 & ~n13279;
  assign n13281 = ~n6712 & ~n10781;
  assign n13282 = controllable_hmaster1 & ~n13281;
  assign n13283 = ~n6719 & ~n13282;
  assign n13284 = ~i_hbusreq3 & ~n13283;
  assign n13285 = ~n13280 & ~n13284;
  assign n13286 = ~controllable_hmaster2 & ~n13285;
  assign n13287 = ~n13276 & ~n13286;
  assign n13288 = ~controllable_hgrant3 & ~n13287;
  assign n13289 = ~n12785 & ~n13288;
  assign n13290 = controllable_nhgrant0 & ~n13289;
  assign n13291 = ~n12827 & ~n13290;
  assign n13292 = ~n3281 & ~n13291;
  assign n13293 = ~n3281 & ~n13292;
  assign n13294 = ~n3378 & ~n13293;
  assign n13295 = ~n13266 & ~n13294;
  assign n13296 = n3492 & ~n13295;
  assign n13297 = n3492 & ~n13296;
  assign n13298 = n3485 & ~n13297;
  assign n13299 = n3485 & ~n13298;
  assign n13300 = ~n3476 & ~n13299;
  assign n13301 = ~n8029 & ~n12886;
  assign n13302 = controllable_hmaster0 & ~n13301;
  assign n13303 = ~n7328 & ~n13302;
  assign n13304 = controllable_hmaster1 & ~n13303;
  assign n13305 = ~n7342 & ~n13304;
  assign n13306 = i_hbusreq3 & ~n13305;
  assign n13307 = ~n8036 & ~n12898;
  assign n13308 = controllable_hmaster0 & ~n13307;
  assign n13309 = ~n12906 & ~n13308;
  assign n13310 = controllable_hmaster1 & ~n13309;
  assign n13311 = ~n12918 & ~n13310;
  assign n13312 = ~i_hbusreq3 & ~n13311;
  assign n13313 = ~n13306 & ~n13312;
  assign n13314 = ~controllable_hmaster2 & ~n13313;
  assign n13315 = ~n12884 & ~n13314;
  assign n13316 = ~controllable_hgrant3 & ~n13315;
  assign n13317 = ~n12856 & ~n13316;
  assign n13318 = controllable_nhgrant0 & ~n13317;
  assign n13319 = ~n12942 & ~n13318;
  assign n13320 = ~n3281 & ~n13319;
  assign n13321 = ~n3281 & ~n13320;
  assign n13322 = n3378 & ~n13321;
  assign n13323 = ~n6762 & ~n12976;
  assign n13324 = ~controllable_hmaster0 & ~n13323;
  assign n13325 = ~n8055 & ~n13324;
  assign n13326 = ~controllable_hmaster1 & ~n13325;
  assign n13327 = ~n8054 & ~n13326;
  assign n13328 = i_hbusreq3 & ~n13327;
  assign n13329 = ~n6772 & ~n12986;
  assign n13330 = controllable_hmaster1 & ~n13329;
  assign n13331 = controllable_hmaster0 & ~n13329;
  assign n13332 = ~n6772 & ~n12994;
  assign n13333 = ~controllable_hmaster0 & ~n13332;
  assign n13334 = ~n13331 & ~n13333;
  assign n13335 = ~controllable_hmaster1 & ~n13334;
  assign n13336 = ~n13330 & ~n13335;
  assign n13337 = ~i_hbusreq3 & ~n13336;
  assign n13338 = ~n13328 & ~n13337;
  assign n13339 = controllable_hmaster2 & ~n13338;
  assign n13340 = ~n8056 & ~n13004;
  assign n13341 = controllable_hmaster0 & ~n13340;
  assign n13342 = ~n8078 & ~n13341;
  assign n13343 = controllable_hmaster1 & ~n13342;
  assign n13344 = ~n8085 & ~n13343;
  assign n13345 = i_hbusreq3 & ~n13344;
  assign n13346 = ~n8066 & ~n13016;
  assign n13347 = controllable_hmaster0 & ~n13346;
  assign n13348 = ~n6813 & ~n13022;
  assign n13349 = ~controllable_hmaster0 & ~n13348;
  assign n13350 = ~n13347 & ~n13349;
  assign n13351 = controllable_hmaster1 & ~n13350;
  assign n13352 = ~n6772 & ~n13030;
  assign n13353 = controllable_hmaster0 & ~n13352;
  assign n13354 = ~n6831 & ~n13036;
  assign n13355 = ~controllable_hmaster0 & ~n13354;
  assign n13356 = ~n13353 & ~n13355;
  assign n13357 = ~controllable_hmaster1 & ~n13356;
  assign n13358 = ~n13351 & ~n13357;
  assign n13359 = ~i_hbusreq3 & ~n13358;
  assign n13360 = ~n13345 & ~n13359;
  assign n13361 = ~controllable_hmaster2 & ~n13360;
  assign n13362 = ~n13339 & ~n13361;
  assign n13363 = ~controllable_hgrant3 & ~n13362;
  assign n13364 = ~n12974 & ~n13363;
  assign n13365 = controllable_nhgrant0 & ~n13364;
  assign n13366 = ~n13064 & ~n13365;
  assign n13367 = ~n3281 & ~n13366;
  assign n13368 = ~n3281 & ~n13367;
  assign n13369 = ~n3378 & ~n13368;
  assign n13370 = ~n13322 & ~n13369;
  assign n13371 = n3492 & ~n13370;
  assign n13372 = n3492 & ~n13371;
  assign n13373 = n3485 & ~n13372;
  assign n13374 = n3485 & ~n13373;
  assign n13375 = n3476 & ~n13374;
  assign n13376 = ~n13300 & ~n13375;
  assign n13377 = n3374 & ~n13376;
  assign n13378 = ~n7986 & ~n13377;
  assign n13379 = n3655 & ~n13378;
  assign n13380 = ~n5291 & ~n11203;
  assign n13381 = controllable_hmaster1 & ~n13380;
  assign n13382 = ~n5305 & ~n13381;
  assign n13383 = i_hbusreq3 & ~n13382;
  assign n13384 = ~n5311 & ~n11216;
  assign n13385 = controllable_hmaster1 & ~n13384;
  assign n13386 = ~n5334 & ~n13385;
  assign n13387 = ~i_hbusreq3 & ~n13386;
  assign n13388 = ~n13383 & ~n13387;
  assign n13389 = ~controllable_hmaster2 & ~n13388;
  assign n13390 = ~n12741 & ~n13389;
  assign n13391 = ~controllable_hgrant3 & ~n13390;
  assign n13392 = ~n12731 & ~n13391;
  assign n13393 = controllable_nhgrant0 & ~n13392;
  assign n13394 = ~n12773 & ~n13393;
  assign n13395 = ~n3281 & ~n13394;
  assign n13396 = ~n3281 & ~n13395;
  assign n13397 = n3378 & ~n13396;
  assign n13398 = ~n6860 & ~n12617;
  assign n13399 = ~controllable_hmaster1 & ~n13398;
  assign n13400 = ~n6859 & ~n13399;
  assign n13401 = i_hbusreq3 & ~n13400;
  assign n13402 = ~n6867 & ~n12623;
  assign n13403 = ~controllable_hmaster1 & ~n13402;
  assign n13404 = ~n6866 & ~n13403;
  assign n13405 = ~i_hbusreq3 & ~n13404;
  assign n13406 = ~n13401 & ~n13405;
  assign n13407 = controllable_hmaster2 & ~n13406;
  assign n13408 = ~n6929 & ~n11203;
  assign n13409 = controllable_hmaster1 & ~n13408;
  assign n13410 = ~n6936 & ~n13409;
  assign n13411 = i_hbusreq3 & ~n13410;
  assign n13412 = ~n6942 & ~n11216;
  assign n13413 = controllable_hmaster1 & ~n13412;
  assign n13414 = ~n6951 & ~n13413;
  assign n13415 = ~i_hbusreq3 & ~n13414;
  assign n13416 = ~n13411 & ~n13415;
  assign n13417 = ~controllable_hmaster2 & ~n13416;
  assign n13418 = ~n13407 & ~n13417;
  assign n13419 = ~controllable_hgrant3 & ~n13418;
  assign n13420 = ~n12785 & ~n13419;
  assign n13421 = controllable_nhgrant0 & ~n13420;
  assign n13422 = ~n12827 & ~n13421;
  assign n13423 = ~n3281 & ~n13422;
  assign n13424 = ~n3281 & ~n13423;
  assign n13425 = ~n3378 & ~n13424;
  assign n13426 = ~n13397 & ~n13425;
  assign n13427 = n3492 & ~n13426;
  assign n13428 = n3492 & ~n13427;
  assign n13429 = n3485 & ~n13428;
  assign n13430 = n3485 & ~n13429;
  assign n13431 = ~n3476 & ~n13430;
  assign n13432 = ~n8029 & ~n13132;
  assign n13433 = controllable_hmaster0 & ~n13432;
  assign n13434 = ~n7328 & ~n13433;
  assign n13435 = controllable_hmaster1 & ~n13434;
  assign n13436 = ~n7342 & ~n13435;
  assign n13437 = i_hbusreq3 & ~n13436;
  assign n13438 = ~n8036 & ~n13143;
  assign n13439 = controllable_hmaster0 & ~n13438;
  assign n13440 = ~n12906 & ~n13439;
  assign n13441 = controllable_hmaster1 & ~n13440;
  assign n13442 = ~n12918 & ~n13441;
  assign n13443 = ~i_hbusreq3 & ~n13442;
  assign n13444 = ~n13437 & ~n13443;
  assign n13445 = ~controllable_hmaster2 & ~n13444;
  assign n13446 = ~n12884 & ~n13445;
  assign n13447 = ~controllable_hgrant3 & ~n13446;
  assign n13448 = ~n12856 & ~n13447;
  assign n13449 = controllable_nhgrant0 & ~n13448;
  assign n13450 = ~n12942 & ~n13449;
  assign n13451 = ~n3281 & ~n13450;
  assign n13452 = ~n3281 & ~n13451;
  assign n13453 = n3378 & ~n13452;
  assign n13454 = ~n6762 & ~n13161;
  assign n13455 = ~controllable_hmaster0 & ~n13454;
  assign n13456 = ~n8212 & ~n13455;
  assign n13457 = ~controllable_hmaster1 & ~n13456;
  assign n13458 = ~n8211 & ~n13457;
  assign n13459 = i_hbusreq3 & ~n13458;
  assign n13460 = ~n6772 & ~n13171;
  assign n13461 = controllable_hmaster1 & ~n13460;
  assign n13462 = controllable_hmaster0 & ~n13460;
  assign n13463 = ~n6772 & ~n13179;
  assign n13464 = ~controllable_hmaster0 & ~n13463;
  assign n13465 = ~n13462 & ~n13464;
  assign n13466 = ~controllable_hmaster1 & ~n13465;
  assign n13467 = ~n13461 & ~n13466;
  assign n13468 = ~i_hbusreq3 & ~n13467;
  assign n13469 = ~n13459 & ~n13468;
  assign n13470 = controllable_hmaster2 & ~n13469;
  assign n13471 = ~n8056 & ~n13189;
  assign n13472 = controllable_hmaster0 & ~n13471;
  assign n13473 = ~n8233 & ~n13472;
  assign n13474 = controllable_hmaster1 & ~n13473;
  assign n13475 = ~n8240 & ~n13474;
  assign n13476 = i_hbusreq3 & ~n13475;
  assign n13477 = ~n8066 & ~n13200;
  assign n13478 = controllable_hmaster0 & ~n13477;
  assign n13479 = ~n6813 & ~n13206;
  assign n13480 = ~controllable_hmaster0 & ~n13479;
  assign n13481 = ~n13478 & ~n13480;
  assign n13482 = controllable_hmaster1 & ~n13481;
  assign n13483 = ~n6772 & ~n13214;
  assign n13484 = controllable_hmaster0 & ~n13483;
  assign n13485 = ~n6831 & ~n13220;
  assign n13486 = ~controllable_hmaster0 & ~n13485;
  assign n13487 = ~n13484 & ~n13486;
  assign n13488 = ~controllable_hmaster1 & ~n13487;
  assign n13489 = ~n13482 & ~n13488;
  assign n13490 = ~i_hbusreq3 & ~n13489;
  assign n13491 = ~n13476 & ~n13490;
  assign n13492 = ~controllable_hmaster2 & ~n13491;
  assign n13493 = ~n13470 & ~n13492;
  assign n13494 = ~controllable_hgrant3 & ~n13493;
  assign n13495 = ~n12974 & ~n13494;
  assign n13496 = controllable_nhgrant0 & ~n13495;
  assign n13497 = ~n13064 & ~n13496;
  assign n13498 = ~n3281 & ~n13497;
  assign n13499 = ~n3281 & ~n13498;
  assign n13500 = ~n3378 & ~n13499;
  assign n13501 = ~n13453 & ~n13500;
  assign n13502 = n3492 & ~n13501;
  assign n13503 = n3492 & ~n13502;
  assign n13504 = n3485 & ~n13503;
  assign n13505 = n3485 & ~n13504;
  assign n13506 = n3476 & ~n13505;
  assign n13507 = ~n13431 & ~n13506;
  assign n13508 = n3374 & ~n13507;
  assign n13509 = ~n8145 & ~n13508;
  assign n13510 = ~n3655 & ~n13509;
  assign n13511 = ~n13379 & ~n13510;
  assign n13512 = ~n3652 & ~n13511;
  assign n13513 = ~n13248 & ~n13512;
  assign n13514 = n3368 & ~n13513;
  assign n13515 = ~n12723 & ~n13514;
  assign n13516 = n3362 & ~n13515;
  assign n13517 = n3492 & ~n12143;
  assign n13518 = ~n3631 & ~n13517;
  assign n13519 = n3485 & ~n13518;
  assign n13520 = ~n3630 & ~n13519;
  assign n13521 = ~n3476 & ~n13520;
  assign n13522 = n3492 & ~n12297;
  assign n13523 = ~n3631 & ~n13522;
  assign n13524 = n3485 & ~n13523;
  assign n13525 = ~n8312 & ~n13524;
  assign n13526 = n3476 & ~n13525;
  assign n13527 = ~n13521 & ~n13526;
  assign n13528 = n3374 & ~n13527;
  assign n13529 = ~n8316 & ~n13528;
  assign n13530 = n3655 & ~n13529;
  assign n13531 = n3492 & ~n12370;
  assign n13532 = ~n3631 & ~n13531;
  assign n13533 = n3485 & ~n13532;
  assign n13534 = ~n3630 & ~n13533;
  assign n13535 = ~n3476 & ~n13534;
  assign n13536 = n3492 & ~n12450;
  assign n13537 = ~n3631 & ~n13536;
  assign n13538 = n3485 & ~n13537;
  assign n13539 = ~n8369 & ~n13538;
  assign n13540 = n3476 & ~n13539;
  assign n13541 = ~n13535 & ~n13540;
  assign n13542 = n3374 & ~n13541;
  assign n13543 = ~n8373 & ~n13542;
  assign n13544 = ~n3655 & ~n13543;
  assign n13545 = ~n13530 & ~n13544;
  assign n13546 = n3652 & ~n13545;
  assign n13547 = n3492 & ~n12518;
  assign n13548 = ~n3631 & ~n13547;
  assign n13549 = n3485 & ~n13548;
  assign n13550 = ~n3630 & ~n13549;
  assign n13551 = ~n3476 & ~n13550;
  assign n13552 = n3492 & ~n12580;
  assign n13553 = ~n3631 & ~n13552;
  assign n13554 = n3485 & ~n13553;
  assign n13555 = ~n8436 & ~n13554;
  assign n13556 = n3476 & ~n13555;
  assign n13557 = ~n13551 & ~n13556;
  assign n13558 = n3374 & ~n13557;
  assign n13559 = ~n8440 & ~n13558;
  assign n13560 = n3655 & ~n13559;
  assign n13561 = n3492 & ~n12646;
  assign n13562 = ~n3631 & ~n13561;
  assign n13563 = n3485 & ~n13562;
  assign n13564 = ~n3630 & ~n13563;
  assign n13565 = ~n3476 & ~n13564;
  assign n13566 = n3492 & ~n12708;
  assign n13567 = ~n3631 & ~n13566;
  assign n13568 = n3485 & ~n13567;
  assign n13569 = ~n8493 & ~n13568;
  assign n13570 = n3476 & ~n13569;
  assign n13571 = ~n13565 & ~n13570;
  assign n13572 = n3374 & ~n13571;
  assign n13573 = ~n8497 & ~n13572;
  assign n13574 = ~n3655 & ~n13573;
  assign n13575 = ~n13560 & ~n13574;
  assign n13576 = ~n3652 & ~n13575;
  assign n13577 = ~n13546 & ~n13576;
  assign n13578 = ~n3368 & ~n13577;
  assign n13579 = n3492 & ~n12830;
  assign n13580 = n3492 & ~n13579;
  assign n13581 = n3485 & ~n13580;
  assign n13582 = n3485 & ~n13581;
  assign n13583 = ~n3476 & ~n13582;
  assign n13584 = n3492 & ~n13067;
  assign n13585 = n3492 & ~n13584;
  assign n13586 = n3485 & ~n13585;
  assign n13587 = ~n8538 & ~n13586;
  assign n13588 = n3476 & ~n13587;
  assign n13589 = ~n13583 & ~n13588;
  assign n13590 = n3374 & ~n13589;
  assign n13591 = ~n8529 & ~n13590;
  assign n13592 = n3655 & ~n13591;
  assign n13593 = n3492 & ~n13123;
  assign n13594 = n3492 & ~n13593;
  assign n13595 = n3485 & ~n13594;
  assign n13596 = n3485 & ~n13595;
  assign n13597 = ~n3476 & ~n13596;
  assign n13598 = n3492 & ~n13235;
  assign n13599 = n3492 & ~n13598;
  assign n13600 = n3485 & ~n13599;
  assign n13601 = ~n8565 & ~n13600;
  assign n13602 = n3476 & ~n13601;
  assign n13603 = ~n13597 & ~n13602;
  assign n13604 = n3374 & ~n13603;
  assign n13605 = ~n8556 & ~n13604;
  assign n13606 = ~n3655 & ~n13605;
  assign n13607 = ~n13592 & ~n13606;
  assign n13608 = n3652 & ~n13607;
  assign n13609 = n3492 & ~n13293;
  assign n13610 = n3492 & ~n13609;
  assign n13611 = n3485 & ~n13610;
  assign n13612 = n3485 & ~n13611;
  assign n13613 = ~n3476 & ~n13612;
  assign n13614 = n3492 & ~n13368;
  assign n13615 = n3492 & ~n13614;
  assign n13616 = n3485 & ~n13615;
  assign n13617 = ~n8594 & ~n13616;
  assign n13618 = n3476 & ~n13617;
  assign n13619 = ~n13613 & ~n13618;
  assign n13620 = n3374 & ~n13619;
  assign n13621 = ~n8585 & ~n13620;
  assign n13622 = n3655 & ~n13621;
  assign n13623 = n3492 & ~n13424;
  assign n13624 = n3492 & ~n13623;
  assign n13625 = n3485 & ~n13624;
  assign n13626 = n3485 & ~n13625;
  assign n13627 = ~n3476 & ~n13626;
  assign n13628 = n3492 & ~n13499;
  assign n13629 = n3492 & ~n13628;
  assign n13630 = n3485 & ~n13629;
  assign n13631 = ~n8621 & ~n13630;
  assign n13632 = n3476 & ~n13631;
  assign n13633 = ~n13627 & ~n13632;
  assign n13634 = n3374 & ~n13633;
  assign n13635 = ~n8612 & ~n13634;
  assign n13636 = ~n3655 & ~n13635;
  assign n13637 = ~n13622 & ~n13636;
  assign n13638 = ~n3652 & ~n13637;
  assign n13639 = ~n13608 & ~n13638;
  assign n13640 = n3368 & ~n13639;
  assign n13641 = ~n13578 & ~n13640;
  assign n13642 = ~n3362 & ~n13641;
  assign n13643 = ~n13516 & ~n13642;
  assign n13644 = n3359 & ~n13643;
  assign n13645 = ~n8639 & ~n13524;
  assign n13646 = n3476 & ~n13645;
  assign n13647 = ~n13521 & ~n13646;
  assign n13648 = n3374 & ~n13647;
  assign n13649 = ~n8643 & ~n13648;
  assign n13650 = n3655 & ~n13649;
  assign n13651 = ~n8650 & ~n13538;
  assign n13652 = n3476 & ~n13651;
  assign n13653 = ~n13535 & ~n13652;
  assign n13654 = n3374 & ~n13653;
  assign n13655 = ~n8654 & ~n13654;
  assign n13656 = ~n3655 & ~n13655;
  assign n13657 = ~n13650 & ~n13656;
  assign n13658 = n3652 & ~n13657;
  assign n13659 = ~n8663 & ~n13554;
  assign n13660 = n3476 & ~n13659;
  assign n13661 = ~n13551 & ~n13660;
  assign n13662 = n3374 & ~n13661;
  assign n13663 = ~n8667 & ~n13662;
  assign n13664 = n3655 & ~n13663;
  assign n13665 = ~n8674 & ~n13568;
  assign n13666 = n3476 & ~n13665;
  assign n13667 = ~n13565 & ~n13666;
  assign n13668 = n3374 & ~n13667;
  assign n13669 = ~n8678 & ~n13668;
  assign n13670 = ~n3655 & ~n13669;
  assign n13671 = ~n13664 & ~n13670;
  assign n13672 = ~n3652 & ~n13671;
  assign n13673 = ~n13658 & ~n13672;
  assign n13674 = ~n3368 & ~n13673;
  assign n13675 = ~n8694 & ~n13586;
  assign n13676 = n3476 & ~n13675;
  assign n13677 = ~n13583 & ~n13676;
  assign n13678 = n3374 & ~n13677;
  assign n13679 = ~n8693 & ~n13678;
  assign n13680 = n3655 & ~n13679;
  assign n13681 = ~n8705 & ~n13600;
  assign n13682 = n3476 & ~n13681;
  assign n13683 = ~n13597 & ~n13682;
  assign n13684 = n3374 & ~n13683;
  assign n13685 = ~n8704 & ~n13684;
  assign n13686 = ~n3655 & ~n13685;
  assign n13687 = ~n13680 & ~n13686;
  assign n13688 = n3652 & ~n13687;
  assign n13689 = ~n8718 & ~n13616;
  assign n13690 = n3476 & ~n13689;
  assign n13691 = ~n13613 & ~n13690;
  assign n13692 = n3374 & ~n13691;
  assign n13693 = ~n8717 & ~n13692;
  assign n13694 = n3655 & ~n13693;
  assign n13695 = ~n8729 & ~n13630;
  assign n13696 = n3476 & ~n13695;
  assign n13697 = ~n13627 & ~n13696;
  assign n13698 = n3374 & ~n13697;
  assign n13699 = ~n8728 & ~n13698;
  assign n13700 = ~n3655 & ~n13699;
  assign n13701 = ~n13694 & ~n13700;
  assign n13702 = ~n3652 & ~n13701;
  assign n13703 = ~n13688 & ~n13702;
  assign n13704 = n3368 & ~n13703;
  assign n13705 = ~n13674 & ~n13704;
  assign n13706 = n3362 & ~n13705;
  assign n13707 = n3378 & ~n12143;
  assign n13708 = ~n8906 & ~n13707;
  assign n13709 = n3492 & ~n13708;
  assign n13710 = ~n3631 & ~n13709;
  assign n13711 = n3485 & ~n13710;
  assign n13712 = ~n3630 & ~n13711;
  assign n13713 = ~n3476 & ~n13712;
  assign n13714 = n3378 & ~n12297;
  assign n13715 = ~n9100 & ~n13714;
  assign n13716 = n3492 & ~n13715;
  assign n13717 = ~n8309 & ~n13716;
  assign n13718 = n3485 & ~n13717;
  assign n13719 = ~n8639 & ~n13718;
  assign n13720 = n3476 & ~n13719;
  assign n13721 = ~n13713 & ~n13720;
  assign n13722 = n3374 & ~n13721;
  assign n13723 = ~n8801 & ~n13722;
  assign n13724 = n3655 & ~n13723;
  assign n13725 = n3378 & ~n12370;
  assign n13726 = ~n9240 & ~n13725;
  assign n13727 = n3492 & ~n13726;
  assign n13728 = ~n3631 & ~n13727;
  assign n13729 = n3485 & ~n13728;
  assign n13730 = ~n3630 & ~n13729;
  assign n13731 = ~n3476 & ~n13730;
  assign n13732 = n3378 & ~n12450;
  assign n13733 = ~n9374 & ~n13732;
  assign n13734 = n3492 & ~n13733;
  assign n13735 = ~n8367 & ~n13734;
  assign n13736 = n3485 & ~n13735;
  assign n13737 = ~n8650 & ~n13736;
  assign n13738 = n3476 & ~n13737;
  assign n13739 = ~n13731 & ~n13738;
  assign n13740 = n3374 & ~n13739;
  assign n13741 = ~n9147 & ~n13740;
  assign n13742 = ~n3655 & ~n13741;
  assign n13743 = ~n13724 & ~n13742;
  assign n13744 = n3652 & ~n13743;
  assign n13745 = n3378 & ~n12518;
  assign n13746 = ~n9469 & ~n13745;
  assign n13747 = n3492 & ~n13746;
  assign n13748 = ~n3631 & ~n13747;
  assign n13749 = n3485 & ~n13748;
  assign n13750 = ~n3630 & ~n13749;
  assign n13751 = ~n3476 & ~n13750;
  assign n13752 = n3378 & ~n12580;
  assign n13753 = ~n9531 & ~n13752;
  assign n13754 = n3492 & ~n13753;
  assign n13755 = ~n8434 & ~n13754;
  assign n13756 = n3485 & ~n13755;
  assign n13757 = ~n8663 & ~n13756;
  assign n13758 = n3476 & ~n13757;
  assign n13759 = ~n13751 & ~n13758;
  assign n13760 = n3374 & ~n13759;
  assign n13761 = ~n9421 & ~n13760;
  assign n13762 = n3655 & ~n13761;
  assign n13763 = n3378 & ~n12646;
  assign n13764 = ~n9623 & ~n13763;
  assign n13765 = n3492 & ~n13764;
  assign n13766 = ~n3631 & ~n13765;
  assign n13767 = n3485 & ~n13766;
  assign n13768 = ~n3630 & ~n13767;
  assign n13769 = ~n3476 & ~n13768;
  assign n13770 = n3378 & ~n12708;
  assign n13771 = ~n9683 & ~n13770;
  assign n13772 = n3492 & ~n13771;
  assign n13773 = ~n8491 & ~n13772;
  assign n13774 = n3485 & ~n13773;
  assign n13775 = ~n8674 & ~n13774;
  assign n13776 = n3476 & ~n13775;
  assign n13777 = ~n13769 & ~n13776;
  assign n13778 = n3374 & ~n13777;
  assign n13779 = ~n9575 & ~n13778;
  assign n13780 = ~n3655 & ~n13779;
  assign n13781 = ~n13762 & ~n13780;
  assign n13782 = ~n3652 & ~n13781;
  assign n13783 = ~n13744 & ~n13782;
  assign n13784 = ~n3368 & ~n13783;
  assign n13785 = n3378 & ~n12830;
  assign n13786 = ~n9865 & ~n13785;
  assign n13787 = n3492 & ~n13786;
  assign n13788 = n3492 & ~n13787;
  assign n13789 = n3485 & ~n13788;
  assign n13790 = n3485 & ~n13789;
  assign n13791 = ~n3476 & ~n13790;
  assign n13792 = ~n9878 & ~n12257;
  assign n13793 = ~controllable_hmaster1 & ~n13792;
  assign n13794 = ~n9877 & ~n13793;
  assign n13795 = i_hbusreq3 & ~n13794;
  assign n13796 = ~n5863 & ~n9895;
  assign n13797 = ~i_hbusreq2 & ~n13796;
  assign n13798 = ~n9883 & ~n13797;
  assign n13799 = ~controllable_hgrant2 & ~n13798;
  assign n13800 = ~n5862 & ~n13799;
  assign n13801 = controllable_hmaster1 & ~n13800;
  assign n13802 = controllable_hmaster0 & ~n13800;
  assign n13803 = ~n12268 & ~n13802;
  assign n13804 = ~controllable_hmaster1 & ~n13803;
  assign n13805 = ~n13801 & ~n13804;
  assign n13806 = ~i_hbusreq3 & ~n13805;
  assign n13807 = ~n13795 & ~n13806;
  assign n13808 = controllable_hmaster2 & ~n13807;
  assign n13809 = ~n9910 & ~n13012;
  assign n13810 = ~i_hbusreq2 & ~n13809;
  assign n13811 = ~n5636 & ~n13810;
  assign n13812 = ~controllable_hgrant2 & ~n13811;
  assign n13813 = ~n7507 & ~n13812;
  assign n13814 = controllable_hmaster0 & ~n13813;
  assign n13815 = ~n5952 & ~n13814;
  assign n13816 = controllable_hmaster1 & ~n13815;
  assign n13817 = ~n5998 & ~n13816;
  assign n13818 = ~i_hbusreq3 & ~n13817;
  assign n13819 = ~n12278 & ~n13818;
  assign n13820 = ~controllable_hmaster2 & ~n13819;
  assign n13821 = ~n13808 & ~n13820;
  assign n13822 = ~controllable_hgrant3 & ~n13821;
  assign n13823 = ~n12974 & ~n13822;
  assign n13824 = controllable_nhgrant0 & ~n13823;
  assign n13825 = i_hbusreq3 & ~n9965;
  assign n13826 = ~i_hbusreq3 & ~n10003;
  assign n13827 = ~n13825 & ~n13826;
  assign n13828 = controllable_hmaster2 & ~n13827;
  assign n13829 = ~controllable_hmaster0 & ~n9965;
  assign n13830 = ~n10215 & ~n13829;
  assign n13831 = controllable_hmaster1 & ~n13830;
  assign n13832 = ~n10042 & ~n13831;
  assign n13833 = i_hbusreq3 & ~n13832;
  assign n13834 = controllable_hmaster0 & ~n10021;
  assign n13835 = ~controllable_hmaster0 & ~n10003;
  assign n13836 = ~n13834 & ~n13835;
  assign n13837 = controllable_hmaster1 & ~n13836;
  assign n13838 = ~n10063 & ~n13837;
  assign n13839 = ~i_hbusreq3 & ~n13838;
  assign n13840 = ~n13833 & ~n13839;
  assign n13841 = ~controllable_hmaster2 & ~n13840;
  assign n13842 = ~n13828 & ~n13841;
  assign n13843 = ~controllable_hgrant3 & ~n13842;
  assign n13844 = ~n12813 & ~n13843;
  assign n13845 = ~controllable_nhgrant0 & ~n13844;
  assign n13846 = ~n13824 & ~n13845;
  assign n13847 = ~n3281 & ~n13846;
  assign n13848 = ~n3281 & ~n13847;
  assign n13849 = n3378 & ~n13848;
  assign n13850 = ~n10244 & ~n13849;
  assign n13851 = n3492 & ~n13850;
  assign n13852 = ~n8536 & ~n13851;
  assign n13853 = n3485 & ~n13852;
  assign n13854 = ~n8694 & ~n13853;
  assign n13855 = n3476 & ~n13854;
  assign n13856 = ~n13791 & ~n13855;
  assign n13857 = n3374 & ~n13856;
  assign n13858 = ~n9769 & ~n13857;
  assign n13859 = n3655 & ~n13858;
  assign n13860 = n3378 & ~n13123;
  assign n13861 = ~n10390 & ~n13860;
  assign n13862 = n3492 & ~n13861;
  assign n13863 = n3492 & ~n13862;
  assign n13864 = n3485 & ~n13863;
  assign n13865 = n3485 & ~n13864;
  assign n13866 = ~n3476 & ~n13865;
  assign n13867 = ~n4015 & ~n10483;
  assign n13868 = ~controllable_hgrant2 & ~n13867;
  assign n13869 = ~n5616 & ~n13868;
  assign n13870 = ~controllable_hmaster0 & ~n13869;
  assign n13871 = ~n10409 & ~n13870;
  assign n13872 = ~controllable_hmaster1 & ~n13871;
  assign n13873 = ~n10408 & ~n13872;
  assign n13874 = i_hbusreq3 & ~n13873;
  assign n13875 = ~n5863 & ~n10443;
  assign n13876 = ~i_hbusreq2 & ~n13875;
  assign n13877 = ~n10421 & ~n13876;
  assign n13878 = ~controllable_hgrant2 & ~n13877;
  assign n13879 = ~n5862 & ~n13878;
  assign n13880 = controllable_hmaster1 & ~n13879;
  assign n13881 = controllable_hmaster0 & ~n13879;
  assign n13882 = i_hbusreq2 & ~n13867;
  assign n13883 = ~n4064 & ~n10521;
  assign n13884 = ~i_hbusreq2 & ~n13883;
  assign n13885 = ~n13882 & ~n13884;
  assign n13886 = ~controllable_hgrant2 & ~n13885;
  assign n13887 = ~n5862 & ~n13886;
  assign n13888 = ~controllable_hmaster0 & ~n13887;
  assign n13889 = ~n13881 & ~n13888;
  assign n13890 = ~controllable_hmaster1 & ~n13889;
  assign n13891 = ~n13880 & ~n13890;
  assign n13892 = ~i_hbusreq3 & ~n13891;
  assign n13893 = ~n13874 & ~n13892;
  assign n13894 = controllable_hmaster2 & ~n13893;
  assign n13895 = ~n10489 & ~n10592;
  assign n13896 = controllable_hmaster1 & ~n13895;
  assign n13897 = ~n10505 & ~n13896;
  assign n13898 = i_hbusreq3 & ~n13897;
  assign n13899 = ~n10468 & ~n13012;
  assign n13900 = ~i_hbusreq2 & ~n13899;
  assign n13901 = ~n10597 & ~n13900;
  assign n13902 = ~controllable_hgrant2 & ~n13901;
  assign n13903 = ~n7507 & ~n13902;
  assign n13904 = controllable_hmaster0 & ~n13903;
  assign n13905 = ~n5863 & ~n10521;
  assign n13906 = ~i_hbusreq2 & ~n13905;
  assign n13907 = ~n10508 & ~n13906;
  assign n13908 = ~controllable_hgrant2 & ~n13907;
  assign n13909 = ~n5950 & ~n13908;
  assign n13910 = ~controllable_hmaster0 & ~n13909;
  assign n13911 = ~n13904 & ~n13910;
  assign n13912 = controllable_hmaster1 & ~n13911;
  assign n13913 = ~n5863 & ~n10552;
  assign n13914 = ~i_hbusreq2 & ~n13913;
  assign n13915 = ~n10532 & ~n13914;
  assign n13916 = ~controllable_hgrant2 & ~n13915;
  assign n13917 = ~n5862 & ~n13916;
  assign n13918 = controllable_hmaster0 & ~n13917;
  assign n13919 = ~n5982 & ~n10567;
  assign n13920 = ~i_hbusreq2 & ~n13919;
  assign n13921 = ~n10508 & ~n13920;
  assign n13922 = ~controllable_hgrant2 & ~n13921;
  assign n13923 = ~n5981 & ~n13922;
  assign n13924 = ~controllable_hmaster0 & ~n13923;
  assign n13925 = ~n13918 & ~n13924;
  assign n13926 = ~controllable_hmaster1 & ~n13925;
  assign n13927 = ~n13912 & ~n13926;
  assign n13928 = ~i_hbusreq3 & ~n13927;
  assign n13929 = ~n13898 & ~n13928;
  assign n13930 = ~controllable_hmaster2 & ~n13929;
  assign n13931 = ~n13894 & ~n13930;
  assign n13932 = ~controllable_hgrant3 & ~n13931;
  assign n13933 = ~n12974 & ~n13932;
  assign n13934 = controllable_nhgrant0 & ~n13933;
  assign n13935 = ~n13845 & ~n13934;
  assign n13936 = ~n3281 & ~n13935;
  assign n13937 = ~n3281 & ~n13936;
  assign n13938 = n3378 & ~n13937;
  assign n13939 = ~n10705 & ~n13938;
  assign n13940 = n3492 & ~n13939;
  assign n13941 = ~n8563 & ~n13940;
  assign n13942 = n3485 & ~n13941;
  assign n13943 = ~n8705 & ~n13942;
  assign n13944 = n3476 & ~n13943;
  assign n13945 = ~n13866 & ~n13944;
  assign n13946 = n3374 & ~n13945;
  assign n13947 = ~n10311 & ~n13946;
  assign n13948 = ~n3655 & ~n13947;
  assign n13949 = ~n13859 & ~n13948;
  assign n13950 = n3652 & ~n13949;
  assign n13951 = n3378 & ~n13293;
  assign n13952 = ~n10802 & ~n13951;
  assign n13953 = n3492 & ~n13952;
  assign n13954 = n3492 & ~n13953;
  assign n13955 = n3485 & ~n13954;
  assign n13956 = n3485 & ~n13955;
  assign n13957 = ~n3476 & ~n13956;
  assign n13958 = ~n10816 & ~n12255;
  assign n13959 = ~controllable_hmaster0 & ~n13958;
  assign n13960 = ~n10819 & ~n13959;
  assign n13961 = ~controllable_hmaster1 & ~n13960;
  assign n13962 = ~n10818 & ~n13961;
  assign n13963 = i_hbusreq3 & ~n13962;
  assign n13964 = ~n10870 & ~n13799;
  assign n13965 = controllable_hmaster1 & ~n13964;
  assign n13966 = controllable_hmaster0 & ~n13964;
  assign n13967 = ~n10870 & ~n12266;
  assign n13968 = ~controllable_hmaster0 & ~n13967;
  assign n13969 = ~n13966 & ~n13968;
  assign n13970 = ~controllable_hmaster1 & ~n13969;
  assign n13971 = ~n13965 & ~n13970;
  assign n13972 = ~i_hbusreq3 & ~n13971;
  assign n13973 = ~n13963 & ~n13972;
  assign n13974 = controllable_hmaster2 & ~n13973;
  assign n13975 = ~n10924 & ~n11021;
  assign n13976 = controllable_hmaster1 & ~n13975;
  assign n13977 = ~n10931 & ~n13976;
  assign n13978 = i_hbusreq3 & ~n13977;
  assign n13979 = ~n10904 & ~n13812;
  assign n13980 = controllable_hmaster0 & ~n13979;
  assign n13981 = ~n5947 & ~n10972;
  assign n13982 = ~controllable_hmaster0 & ~n13981;
  assign n13983 = ~n13980 & ~n13982;
  assign n13984 = controllable_hmaster1 & ~n13983;
  assign n13985 = ~n5978 & ~n10870;
  assign n13986 = controllable_hmaster0 & ~n13985;
  assign n13987 = ~n5994 & ~n11002;
  assign n13988 = ~controllable_hmaster0 & ~n13987;
  assign n13989 = ~n13986 & ~n13988;
  assign n13990 = ~controllable_hmaster1 & ~n13989;
  assign n13991 = ~n13984 & ~n13990;
  assign n13992 = ~i_hbusreq3 & ~n13991;
  assign n13993 = ~n13978 & ~n13992;
  assign n13994 = ~controllable_hmaster2 & ~n13993;
  assign n13995 = ~n13974 & ~n13994;
  assign n13996 = ~controllable_hgrant3 & ~n13995;
  assign n13997 = ~n12974 & ~n13996;
  assign n13998 = controllable_nhgrant0 & ~n13997;
  assign n13999 = ~n13845 & ~n13998;
  assign n14000 = ~n3281 & ~n13999;
  assign n14001 = ~n3281 & ~n14000;
  assign n14002 = n3378 & ~n14001;
  assign n14003 = ~n11143 & ~n14002;
  assign n14004 = n3492 & ~n14003;
  assign n14005 = ~n8592 & ~n14004;
  assign n14006 = n3485 & ~n14005;
  assign n14007 = ~n8718 & ~n14006;
  assign n14008 = n3476 & ~n14007;
  assign n14009 = ~n13957 & ~n14008;
  assign n14010 = n3374 & ~n14009;
  assign n14011 = ~n10754 & ~n14010;
  assign n14012 = n3655 & ~n14011;
  assign n14013 = n3378 & ~n13424;
  assign n14014 = ~n11236 & ~n14013;
  assign n14015 = n3492 & ~n14014;
  assign n14016 = n3492 & ~n14015;
  assign n14017 = n3485 & ~n14016;
  assign n14018 = n3485 & ~n14017;
  assign n14019 = ~n3476 & ~n14018;
  assign n14020 = ~n10816 & ~n13868;
  assign n14021 = ~controllable_hmaster0 & ~n14020;
  assign n14022 = ~n11245 & ~n14021;
  assign n14023 = ~controllable_hmaster1 & ~n14022;
  assign n14024 = ~n11244 & ~n14023;
  assign n14025 = i_hbusreq3 & ~n14024;
  assign n14026 = ~n10870 & ~n13878;
  assign n14027 = controllable_hmaster1 & ~n14026;
  assign n14028 = controllable_hmaster0 & ~n14026;
  assign n14029 = ~n10870 & ~n13886;
  assign n14030 = ~controllable_hmaster0 & ~n14029;
  assign n14031 = ~n14028 & ~n14030;
  assign n14032 = ~controllable_hmaster1 & ~n14031;
  assign n14033 = ~n14027 & ~n14032;
  assign n14034 = ~i_hbusreq3 & ~n14033;
  assign n14035 = ~n14025 & ~n14034;
  assign n14036 = controllable_hmaster2 & ~n14035;
  assign n14037 = ~n11266 & ~n11302;
  assign n14038 = controllable_hmaster1 & ~n14037;
  assign n14039 = ~n11273 & ~n14038;
  assign n14040 = i_hbusreq3 & ~n14039;
  assign n14041 = ~n10904 & ~n13902;
  assign n14042 = controllable_hmaster0 & ~n14041;
  assign n14043 = ~n10972 & ~n13908;
  assign n14044 = ~controllable_hmaster0 & ~n14043;
  assign n14045 = ~n14042 & ~n14044;
  assign n14046 = controllable_hmaster1 & ~n14045;
  assign n14047 = ~n10870 & ~n13916;
  assign n14048 = controllable_hmaster0 & ~n14047;
  assign n14049 = ~n11002 & ~n13922;
  assign n14050 = ~controllable_hmaster0 & ~n14049;
  assign n14051 = ~n14048 & ~n14050;
  assign n14052 = ~controllable_hmaster1 & ~n14051;
  assign n14053 = ~n14046 & ~n14052;
  assign n14054 = ~i_hbusreq3 & ~n14053;
  assign n14055 = ~n14040 & ~n14054;
  assign n14056 = ~controllable_hmaster2 & ~n14055;
  assign n14057 = ~n14036 & ~n14056;
  assign n14058 = ~controllable_hgrant3 & ~n14057;
  assign n14059 = ~n12974 & ~n14058;
  assign n14060 = controllable_nhgrant0 & ~n14059;
  assign n14061 = ~n13845 & ~n14060;
  assign n14062 = ~n3281 & ~n14061;
  assign n14063 = ~n3281 & ~n14062;
  assign n14064 = n3378 & ~n14063;
  assign n14065 = ~n11352 & ~n14064;
  assign n14066 = n3492 & ~n14065;
  assign n14067 = ~n8619 & ~n14066;
  assign n14068 = n3485 & ~n14067;
  assign n14069 = ~n8729 & ~n14068;
  assign n14070 = n3476 & ~n14069;
  assign n14071 = ~n14019 & ~n14070;
  assign n14072 = n3374 & ~n14071;
  assign n14073 = ~n11190 & ~n14072;
  assign n14074 = ~n3655 & ~n14073;
  assign n14075 = ~n14012 & ~n14074;
  assign n14076 = ~n3652 & ~n14075;
  assign n14077 = ~n13950 & ~n14076;
  assign n14078 = n3368 & ~n14077;
  assign n14079 = ~n13784 & ~n14078;
  assign n14080 = ~n3362 & ~n14079;
  assign n14081 = ~n13706 & ~n14080;
  assign n14082 = ~n3359 & ~n14081;
  assign n14083 = ~n13644 & ~n14082;
  assign n14084 = ~n3356 & ~n14083;
  assign n14085 = ~n12025 & ~n14084;
  assign n14086 = ~n3345 & ~n14085;
  assign n14087 = controllable_hmaster1 & ~n8396;
  assign n14088 = i_hbusreq3 & ~n14087;
  assign n14089 = controllable_hmaster1 & ~n8400;
  assign n14090 = ~i_hbusreq3 & ~n14089;
  assign n14091 = ~n14088 & ~n14090;
  assign n14092 = ~controllable_hmaster2 & ~n14091;
  assign n14093 = ~controllable_hmaster2 & ~n14092;
  assign n14094 = controllable_hgrant3 & ~n14093;
  assign n14095 = ~controllable_hmaster0 & ~n5085;
  assign n14096 = controllable_hmaster1 & ~n14095;
  assign n14097 = controllable_hmaster1 & ~n14096;
  assign n14098 = i_hbusreq3 & ~n14097;
  assign n14099 = ~controllable_hmaster0 & ~n5125;
  assign n14100 = controllable_hmaster1 & ~n14099;
  assign n14101 = controllable_hmaster1 & ~n14100;
  assign n14102 = ~i_hbusreq3 & ~n14101;
  assign n14103 = ~n14098 & ~n14102;
  assign n14104 = ~controllable_hmaster2 & ~n14103;
  assign n14105 = ~controllable_hmaster2 & ~n14104;
  assign n14106 = ~controllable_hgrant3 & ~n14105;
  assign n14107 = ~n14094 & ~n14106;
  assign n14108 = controllable_nhgrant0 & ~n14107;
  assign n14109 = ~controllable_nhgrant0 & ~n14093;
  assign n14110 = ~n14108 & ~n14109;
  assign n14111 = ~n3281 & ~n14110;
  assign n14112 = ~n3281 & ~n14111;
  assign n14113 = n3378 & ~n14112;
  assign n14114 = ~n3407 & ~n14092;
  assign n14115 = controllable_hgrant3 & ~n14114;
  assign n14116 = ~n3461 & ~n14104;
  assign n14117 = ~controllable_hgrant3 & ~n14116;
  assign n14118 = ~n14115 & ~n14117;
  assign n14119 = controllable_nhgrant0 & ~n14118;
  assign n14120 = ~controllable_nhgrant0 & ~n14114;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = ~n3281 & ~n14121;
  assign n14123 = ~n3783 & ~n14122;
  assign n14124 = ~n3378 & ~n14123;
  assign n14125 = ~n14113 & ~n14124;
  assign n14126 = n3492 & ~n14125;
  assign n14127 = ~n3493 & ~n14126;
  assign n14128 = n3485 & ~n14127;
  assign n14129 = ~n3486 & ~n14128;
  assign n14130 = ~n3374 & ~n14129;
  assign n14131 = controllable_hmaster1 & ~n3822;
  assign n14132 = controllable_hmaster1 & ~n14131;
  assign n14133 = i_hbusreq3 & ~n14132;
  assign n14134 = controllable_hmaster1 & ~n3836;
  assign n14135 = controllable_hmaster1 & ~n14134;
  assign n14136 = ~i_hbusreq3 & ~n14135;
  assign n14137 = ~n14133 & ~n14136;
  assign n14138 = ~controllable_hmaster2 & ~n14137;
  assign n14139 = ~controllable_hmaster2 & ~n14138;
  assign n14140 = controllable_hgrant3 & ~n14139;
  assign n14141 = ~controllable_hmaster0 & ~n8818;
  assign n14142 = controllable_hmaster1 & ~n14141;
  assign n14143 = controllable_hmaster1 & ~n14142;
  assign n14144 = i_hbusreq3 & ~n14143;
  assign n14145 = ~controllable_hmaster0 & ~n8840;
  assign n14146 = controllable_hmaster1 & ~n14145;
  assign n14147 = controllable_hmaster1 & ~n14146;
  assign n14148 = ~i_hbusreq3 & ~n14147;
  assign n14149 = ~n14144 & ~n14148;
  assign n14150 = ~controllable_hmaster2 & ~n14149;
  assign n14151 = ~controllable_hmaster2 & ~n14150;
  assign n14152 = ~controllable_hgrant3 & ~n14151;
  assign n14153 = ~n14140 & ~n14152;
  assign n14154 = controllable_nhgrant0 & ~n14153;
  assign n14155 = controllable_hmaster1 & ~n3911;
  assign n14156 = controllable_hmaster1 & ~n14155;
  assign n14157 = i_hbusreq3 & ~n14156;
  assign n14158 = controllable_hmaster1 & ~n3936;
  assign n14159 = controllable_hmaster1 & ~n14158;
  assign n14160 = ~i_hbusreq3 & ~n14159;
  assign n14161 = ~n14157 & ~n14160;
  assign n14162 = ~controllable_hmaster2 & ~n14161;
  assign n14163 = ~controllable_hmaster2 & ~n14162;
  assign n14164 = ~controllable_hgrant3 & ~n14163;
  assign n14165 = ~n14140 & ~n14164;
  assign n14166 = ~controllable_nhgrant0 & ~n14165;
  assign n14167 = ~n14154 & ~n14166;
  assign n14168 = ~n3281 & ~n14167;
  assign n14169 = ~n3281 & ~n14168;
  assign n14170 = n3378 & ~n14169;
  assign n14171 = ~n3407 & ~n14138;
  assign n14172 = controllable_hgrant3 & ~n14171;
  assign n14173 = ~n3530 & ~n14150;
  assign n14174 = ~controllable_hgrant3 & ~n14173;
  assign n14175 = ~n14172 & ~n14174;
  assign n14176 = controllable_nhgrant0 & ~n14175;
  assign n14177 = ~n3407 & ~n14162;
  assign n14178 = ~controllable_hgrant3 & ~n14177;
  assign n14179 = ~n14172 & ~n14178;
  assign n14180 = ~controllable_nhgrant0 & ~n14179;
  assign n14181 = ~n14176 & ~n14180;
  assign n14182 = ~n3281 & ~n14181;
  assign n14183 = ~n3950 & ~n14182;
  assign n14184 = ~n3378 & ~n14183;
  assign n14185 = ~n14170 & ~n14184;
  assign n14186 = n3492 & ~n14185;
  assign n14187 = ~n3493 & ~n14186;
  assign n14188 = n3485 & ~n14187;
  assign n14189 = ~n3486 & ~n14188;
  assign n14190 = ~n3476 & ~n14189;
  assign n14191 = controllable_hgrant2 & ~n11524;
  assign n14192 = controllable_hgrant2 & ~n14191;
  assign n14193 = i_hbusreq3 & ~n14192;
  assign n14194 = controllable_hgrant2 & ~n11532;
  assign n14195 = controllable_hgrant2 & ~n14194;
  assign n14196 = ~i_hbusreq3 & ~n14195;
  assign n14197 = ~n14193 & ~n14196;
  assign n14198 = controllable_hmaster2 & ~n14197;
  assign n14199 = controllable_hmaster0 & ~n14192;
  assign n14200 = ~n5686 & ~n8768;
  assign n14201 = ~controllable_hmaster0 & ~n14200;
  assign n14202 = ~n14199 & ~n14201;
  assign n14203 = controllable_hmaster1 & ~n14202;
  assign n14204 = ~controllable_hmaster1 & ~n14192;
  assign n14205 = ~n14203 & ~n14204;
  assign n14206 = i_hbusreq3 & ~n14205;
  assign n14207 = controllable_hmaster0 & ~n14195;
  assign n14208 = ~n5950 & ~n8836;
  assign n14209 = ~controllable_hmaster0 & ~n14208;
  assign n14210 = ~n14207 & ~n14209;
  assign n14211 = controllable_hmaster1 & ~n14210;
  assign n14212 = ~controllable_hmaster1 & ~n14195;
  assign n14213 = ~n14211 & ~n14212;
  assign n14214 = ~i_hbusreq3 & ~n14213;
  assign n14215 = ~n14206 & ~n14214;
  assign n14216 = ~controllable_hmaster2 & ~n14215;
  assign n14217 = ~n14198 & ~n14216;
  assign n14218 = ~controllable_hgrant3 & ~n14217;
  assign n14219 = ~n14140 & ~n14218;
  assign n14220 = controllable_nhgrant0 & ~n14219;
  assign n14221 = ~n14166 & ~n14220;
  assign n14222 = ~n3281 & ~n14221;
  assign n14223 = ~n3281 & ~n14222;
  assign n14224 = n3378 & ~n14223;
  assign n14225 = ~n3547 & ~n5616;
  assign n14226 = controllable_hmaster1 & ~n14225;
  assign n14227 = controllable_hmaster0 & ~n14225;
  assign n14228 = ~n3554 & ~n14191;
  assign n14229 = ~controllable_hmaster0 & ~n14228;
  assign n14230 = ~n14227 & ~n14229;
  assign n14231 = ~controllable_hmaster1 & ~n14230;
  assign n14232 = ~n14226 & ~n14231;
  assign n14233 = i_hbusreq3 & ~n14232;
  assign n14234 = controllable_hgrant2 & ~n11567;
  assign n14235 = ~n3578 & ~n14234;
  assign n14236 = controllable_hmaster1 & ~n14235;
  assign n14237 = controllable_hmaster0 & ~n14235;
  assign n14238 = ~n3594 & ~n14194;
  assign n14239 = ~controllable_hmaster0 & ~n14238;
  assign n14240 = ~n14237 & ~n14239;
  assign n14241 = ~controllable_hmaster1 & ~n14240;
  assign n14242 = ~n14236 & ~n14241;
  assign n14243 = ~i_hbusreq3 & ~n14242;
  assign n14244 = ~n14233 & ~n14243;
  assign n14245 = controllable_hmaster2 & ~n14244;
  assign n14246 = controllable_hmaster0 & ~n14228;
  assign n14247 = ~n3547 & ~n5686;
  assign n14248 = ~controllable_hmaster0 & ~n14247;
  assign n14249 = ~n14246 & ~n14248;
  assign n14250 = controllable_hmaster1 & ~n14249;
  assign n14251 = ~controllable_hmaster1 & ~n14228;
  assign n14252 = ~n14250 & ~n14251;
  assign n14253 = i_hbusreq3 & ~n14252;
  assign n14254 = controllable_hmaster0 & ~n14238;
  assign n14255 = ~n5950 & ~n11587;
  assign n14256 = ~controllable_hmaster0 & ~n14255;
  assign n14257 = ~n14254 & ~n14256;
  assign n14258 = controllable_hmaster1 & ~n14257;
  assign n14259 = ~controllable_hmaster1 & ~n14238;
  assign n14260 = ~n14258 & ~n14259;
  assign n14261 = ~i_hbusreq3 & ~n14260;
  assign n14262 = ~n14253 & ~n14261;
  assign n14263 = ~controllable_hmaster2 & ~n14262;
  assign n14264 = ~n14245 & ~n14263;
  assign n14265 = ~controllable_hgrant3 & ~n14264;
  assign n14266 = ~n14172 & ~n14265;
  assign n14267 = controllable_nhgrant0 & ~n14266;
  assign n14268 = ~n14180 & ~n14267;
  assign n14269 = ~n3281 & ~n14268;
  assign n14270 = ~n4089 & ~n14269;
  assign n14271 = ~n3378 & ~n14270;
  assign n14272 = ~n14224 & ~n14271;
  assign n14273 = n3492 & ~n14272;
  assign n14274 = ~n3493 & ~n14273;
  assign n14275 = n3485 & ~n14274;
  assign n14276 = ~n3486 & ~n14275;
  assign n14277 = n3476 & ~n14276;
  assign n14278 = ~n14190 & ~n14277;
  assign n14279 = n3374 & ~n14278;
  assign n14280 = ~n14130 & ~n14279;
  assign n14281 = n3655 & ~n14280;
  assign n14282 = ~controllable_hmaster0 & ~n9164;
  assign n14283 = controllable_hmaster1 & ~n14282;
  assign n14284 = controllable_hmaster1 & ~n14283;
  assign n14285 = i_hbusreq3 & ~n14284;
  assign n14286 = ~controllable_hmaster0 & ~n9188;
  assign n14287 = controllable_hmaster1 & ~n14286;
  assign n14288 = controllable_hmaster1 & ~n14287;
  assign n14289 = ~i_hbusreq3 & ~n14288;
  assign n14290 = ~n14285 & ~n14289;
  assign n14291 = ~controllable_hmaster2 & ~n14290;
  assign n14292 = ~controllable_hmaster2 & ~n14291;
  assign n14293 = ~controllable_hgrant3 & ~n14292;
  assign n14294 = ~n14140 & ~n14293;
  assign n14295 = controllable_nhgrant0 & ~n14294;
  assign n14296 = ~n14166 & ~n14295;
  assign n14297 = ~n3281 & ~n14296;
  assign n14298 = ~n3281 & ~n14297;
  assign n14299 = n3378 & ~n14298;
  assign n14300 = ~n3530 & ~n14291;
  assign n14301 = ~controllable_hgrant3 & ~n14300;
  assign n14302 = ~n14172 & ~n14301;
  assign n14303 = controllable_nhgrant0 & ~n14302;
  assign n14304 = ~n14180 & ~n14303;
  assign n14305 = ~n3281 & ~n14304;
  assign n14306 = ~n3950 & ~n14305;
  assign n14307 = ~n3378 & ~n14306;
  assign n14308 = ~n14299 & ~n14307;
  assign n14309 = n3492 & ~n14308;
  assign n14310 = ~n3493 & ~n14309;
  assign n14311 = n3485 & ~n14310;
  assign n14312 = ~n3486 & ~n14311;
  assign n14313 = ~n3476 & ~n14312;
  assign n14314 = ~n5686 & ~n9160;
  assign n14315 = ~controllable_hmaster0 & ~n14314;
  assign n14316 = ~n14199 & ~n14315;
  assign n14317 = controllable_hmaster1 & ~n14316;
  assign n14318 = ~n14204 & ~n14317;
  assign n14319 = i_hbusreq3 & ~n14318;
  assign n14320 = ~n5950 & ~n9184;
  assign n14321 = ~controllable_hmaster0 & ~n14320;
  assign n14322 = ~n14207 & ~n14321;
  assign n14323 = controllable_hmaster1 & ~n14322;
  assign n14324 = ~n14212 & ~n14323;
  assign n14325 = ~i_hbusreq3 & ~n14324;
  assign n14326 = ~n14319 & ~n14325;
  assign n14327 = ~controllable_hmaster2 & ~n14326;
  assign n14328 = ~n14198 & ~n14327;
  assign n14329 = ~controllable_hgrant3 & ~n14328;
  assign n14330 = ~n14140 & ~n14329;
  assign n14331 = controllable_nhgrant0 & ~n14330;
  assign n14332 = ~n14166 & ~n14331;
  assign n14333 = ~n3281 & ~n14332;
  assign n14334 = ~n3281 & ~n14333;
  assign n14335 = n3378 & ~n14334;
  assign n14336 = ~n5686 & ~n11654;
  assign n14337 = ~controllable_hmaster0 & ~n14336;
  assign n14338 = ~n14246 & ~n14337;
  assign n14339 = controllable_hmaster1 & ~n14338;
  assign n14340 = ~n14251 & ~n14339;
  assign n14341 = i_hbusreq3 & ~n14340;
  assign n14342 = ~n5950 & ~n11665;
  assign n14343 = ~controllable_hmaster0 & ~n14342;
  assign n14344 = ~n14254 & ~n14343;
  assign n14345 = controllable_hmaster1 & ~n14344;
  assign n14346 = ~n14259 & ~n14345;
  assign n14347 = ~i_hbusreq3 & ~n14346;
  assign n14348 = ~n14341 & ~n14347;
  assign n14349 = ~controllable_hmaster2 & ~n14348;
  assign n14350 = ~n14245 & ~n14349;
  assign n14351 = ~controllable_hgrant3 & ~n14350;
  assign n14352 = ~n14172 & ~n14351;
  assign n14353 = controllable_nhgrant0 & ~n14352;
  assign n14354 = ~n14180 & ~n14353;
  assign n14355 = ~n3281 & ~n14354;
  assign n14356 = ~n4089 & ~n14355;
  assign n14357 = ~n3378 & ~n14356;
  assign n14358 = ~n14335 & ~n14357;
  assign n14359 = n3492 & ~n14358;
  assign n14360 = ~n3493 & ~n14359;
  assign n14361 = n3485 & ~n14360;
  assign n14362 = ~n3486 & ~n14361;
  assign n14363 = n3476 & ~n14362;
  assign n14364 = ~n14313 & ~n14363;
  assign n14365 = n3374 & ~n14364;
  assign n14366 = ~n14130 & ~n14365;
  assign n14367 = ~n3655 & ~n14366;
  assign n14368 = ~n14281 & ~n14367;
  assign n14369 = n3652 & ~n14368;
  assign n14370 = controllable_hmaster1 & ~n8408;
  assign n14371 = i_hbusreq3 & ~n14370;
  assign n14372 = controllable_hmaster1 & ~n8412;
  assign n14373 = ~i_hbusreq3 & ~n14372;
  assign n14374 = ~n14371 & ~n14373;
  assign n14375 = ~controllable_hmaster2 & ~n14374;
  assign n14376 = ~controllable_hmaster2 & ~n14375;
  assign n14377 = ~controllable_hgrant3 & ~n14376;
  assign n14378 = ~n14094 & ~n14377;
  assign n14379 = controllable_nhgrant0 & ~n14378;
  assign n14380 = ~n14109 & ~n14379;
  assign n14381 = ~n3281 & ~n14380;
  assign n14382 = ~n3281 & ~n14381;
  assign n14383 = n3378 & ~n14382;
  assign n14384 = ~n3423 & ~n9388;
  assign n14385 = controllable_hmaster1 & ~n14384;
  assign n14386 = controllable_hmaster0 & ~n14384;
  assign n14387 = controllable_hmaster0 & ~n14386;
  assign n14388 = ~controllable_hmaster1 & ~n14387;
  assign n14389 = ~n14385 & ~n14388;
  assign n14390 = i_hbusreq3 & ~n14389;
  assign n14391 = ~i_hbusreq0 & ~n3876;
  assign n14392 = ~n3875 & ~n14391;
  assign n14393 = ~i_hbusreq4 & ~n14392;
  assign n14394 = ~n3874 & ~n14393;
  assign n14395 = ~controllable_hgrant4 & ~n14394;
  assign n14396 = ~n3433 & ~n14395;
  assign n14397 = ~i_hbusreq2 & ~n14396;
  assign n14398 = ~n8832 & ~n14397;
  assign n14399 = controllable_hgrant2 & ~n14398;
  assign n14400 = ~n3452 & ~n14399;
  assign n14401 = controllable_hmaster1 & ~n14400;
  assign n14402 = controllable_hmaster0 & ~n14400;
  assign n14403 = controllable_hmaster0 & ~n14402;
  assign n14404 = ~controllable_hmaster1 & ~n14403;
  assign n14405 = ~n14401 & ~n14404;
  assign n14406 = ~i_hbusreq3 & ~n14405;
  assign n14407 = ~n14390 & ~n14406;
  assign n14408 = controllable_hmaster2 & ~n14407;
  assign n14409 = ~n14375 & ~n14408;
  assign n14410 = ~controllable_hgrant3 & ~n14409;
  assign n14411 = ~n14115 & ~n14410;
  assign n14412 = controllable_nhgrant0 & ~n14411;
  assign n14413 = ~n14120 & ~n14412;
  assign n14414 = ~n3281 & ~n14413;
  assign n14415 = ~n3783 & ~n14414;
  assign n14416 = ~n3378 & ~n14415;
  assign n14417 = ~n14383 & ~n14416;
  assign n14418 = n3492 & ~n14417;
  assign n14419 = ~n3493 & ~n14418;
  assign n14420 = n3485 & ~n14419;
  assign n14421 = ~n3486 & ~n14420;
  assign n14422 = ~n3476 & ~n14421;
  assign n14423 = ~n3461 & ~n14375;
  assign n14424 = ~controllable_hgrant3 & ~n14423;
  assign n14425 = ~n14115 & ~n14424;
  assign n14426 = controllable_nhgrant0 & ~n14425;
  assign n14427 = ~n14120 & ~n14426;
  assign n14428 = ~n3281 & ~n14427;
  assign n14429 = ~n3783 & ~n14428;
  assign n14430 = ~n3378 & ~n14429;
  assign n14431 = ~n14383 & ~n14430;
  assign n14432 = ~n3485 & ~n14431;
  assign n14433 = ~n3492 & ~n14431;
  assign n14434 = ~n14418 & ~n14433;
  assign n14435 = n3485 & ~n14434;
  assign n14436 = ~n14432 & ~n14435;
  assign n14437 = n3476 & ~n14436;
  assign n14438 = ~n14422 & ~n14437;
  assign n14439 = ~n3374 & ~n14438;
  assign n14440 = ~controllable_hmaster0 & ~n9436;
  assign n14441 = controllable_hmaster1 & ~n14440;
  assign n14442 = controllable_hmaster1 & ~n14441;
  assign n14443 = i_hbusreq3 & ~n14442;
  assign n14444 = ~controllable_hmaster0 & ~n9449;
  assign n14445 = controllable_hmaster1 & ~n14444;
  assign n14446 = controllable_hmaster1 & ~n14445;
  assign n14447 = ~i_hbusreq3 & ~n14446;
  assign n14448 = ~n14443 & ~n14447;
  assign n14449 = ~controllable_hmaster2 & ~n14448;
  assign n14450 = ~controllable_hmaster2 & ~n14449;
  assign n14451 = ~controllable_hgrant3 & ~n14450;
  assign n14452 = ~n14140 & ~n14451;
  assign n14453 = controllable_nhgrant0 & ~n14452;
  assign n14454 = ~n14166 & ~n14453;
  assign n14455 = ~n3281 & ~n14454;
  assign n14456 = ~n3281 & ~n14455;
  assign n14457 = n3378 & ~n14456;
  assign n14458 = controllable_hmaster0 & ~n9391;
  assign n14459 = ~controllable_hmaster1 & ~n14458;
  assign n14460 = ~n9390 & ~n14459;
  assign n14461 = i_hbusreq3 & ~n14460;
  assign n14462 = ~n3521 & ~n14399;
  assign n14463 = controllable_hmaster1 & ~n14462;
  assign n14464 = controllable_hmaster0 & ~n14462;
  assign n14465 = controllable_hmaster0 & ~n14464;
  assign n14466 = ~controllable_hmaster1 & ~n14465;
  assign n14467 = ~n14463 & ~n14466;
  assign n14468 = ~i_hbusreq3 & ~n14467;
  assign n14469 = ~n14461 & ~n14468;
  assign n14470 = controllable_hmaster2 & ~n14469;
  assign n14471 = ~n14449 & ~n14470;
  assign n14472 = ~controllable_hgrant3 & ~n14471;
  assign n14473 = ~n14172 & ~n14472;
  assign n14474 = controllable_nhgrant0 & ~n14473;
  assign n14475 = ~n14180 & ~n14474;
  assign n14476 = ~n3281 & ~n14475;
  assign n14477 = ~n3950 & ~n14476;
  assign n14478 = ~n3378 & ~n14477;
  assign n14479 = ~n14457 & ~n14478;
  assign n14480 = n3492 & ~n14479;
  assign n14481 = ~n3493 & ~n14480;
  assign n14482 = n3485 & ~n14481;
  assign n14483 = ~n3486 & ~n14482;
  assign n14484 = ~n3476 & ~n14483;
  assign n14485 = i_hready & ~n6007;
  assign n14486 = ~controllable_hgrant4 & ~n14485;
  assign n14487 = ~controllable_hgrant4 & ~n14486;
  assign n14488 = controllable_hgrant2 & ~n14487;
  assign n14489 = controllable_hgrant2 & ~n14488;
  assign n14490 = i_hbusreq3 & ~n14489;
  assign n14491 = i_hbusreq2 & ~n14487;
  assign n14492 = i_hbusreq4 & ~n14485;
  assign n14493 = i_hbusreq0 & ~n14485;
  assign n14494 = i_hready & ~n6018;
  assign n14495 = i_hlock0 & ~n14494;
  assign n14496 = ~i_hlock0 & ~n14485;
  assign n14497 = ~n14495 & ~n14496;
  assign n14498 = ~i_hbusreq0 & ~n14497;
  assign n14499 = ~n14493 & ~n14498;
  assign n14500 = ~i_hbusreq4 & ~n14499;
  assign n14501 = ~n14492 & ~n14500;
  assign n14502 = ~controllable_hgrant4 & ~n14501;
  assign n14503 = ~controllable_hgrant4 & ~n14502;
  assign n14504 = ~i_hbusreq2 & ~n14503;
  assign n14505 = ~n14491 & ~n14504;
  assign n14506 = controllable_hgrant2 & ~n14505;
  assign n14507 = controllable_hgrant2 & ~n14506;
  assign n14508 = ~i_hbusreq3 & ~n14507;
  assign n14509 = ~n14490 & ~n14508;
  assign n14510 = controllable_hmaster2 & ~n14509;
  assign n14511 = controllable_hmaster0 & ~n14489;
  assign n14512 = ~n6786 & ~n8768;
  assign n14513 = ~controllable_hmaster0 & ~n14512;
  assign n14514 = ~n14511 & ~n14513;
  assign n14515 = controllable_hmaster1 & ~n14514;
  assign n14516 = ~controllable_hmaster1 & ~n14489;
  assign n14517 = ~n14515 & ~n14516;
  assign n14518 = i_hbusreq3 & ~n14517;
  assign n14519 = controllable_hmaster0 & ~n14507;
  assign n14520 = ~n6813 & ~n8836;
  assign n14521 = ~controllable_hmaster0 & ~n14520;
  assign n14522 = ~n14519 & ~n14521;
  assign n14523 = controllable_hmaster1 & ~n14522;
  assign n14524 = ~controllable_hmaster1 & ~n14507;
  assign n14525 = ~n14523 & ~n14524;
  assign n14526 = ~i_hbusreq3 & ~n14525;
  assign n14527 = ~n14518 & ~n14526;
  assign n14528 = ~controllable_hmaster2 & ~n14527;
  assign n14529 = ~n14510 & ~n14528;
  assign n14530 = ~controllable_hgrant3 & ~n14529;
  assign n14531 = ~n14140 & ~n14530;
  assign n14532 = controllable_nhgrant0 & ~n14531;
  assign n14533 = ~n14166 & ~n14532;
  assign n14534 = ~n3281 & ~n14533;
  assign n14535 = ~n3281 & ~n14534;
  assign n14536 = n3378 & ~n14535;
  assign n14537 = ~n3547 & ~n9477;
  assign n14538 = controllable_hmaster1 & ~n14537;
  assign n14539 = controllable_hmaster0 & ~n14537;
  assign n14540 = ~n3554 & ~n14488;
  assign n14541 = ~controllable_hmaster0 & ~n14540;
  assign n14542 = ~n14539 & ~n14541;
  assign n14543 = ~controllable_hmaster1 & ~n14542;
  assign n14544 = ~n14538 & ~n14543;
  assign n14545 = i_hbusreq3 & ~n14544;
  assign n14546 = ~n3511 & ~n6018;
  assign n14547 = i_hlock0 & ~n14546;
  assign n14548 = ~n3511 & ~n6007;
  assign n14549 = ~i_hlock0 & ~n14548;
  assign n14550 = ~n14547 & ~n14549;
  assign n14551 = ~i_hbusreq0 & ~n14550;
  assign n14552 = ~n9069 & ~n14551;
  assign n14553 = ~i_hbusreq4 & ~n14552;
  assign n14554 = ~n9068 & ~n14553;
  assign n14555 = ~controllable_hgrant4 & ~n14554;
  assign n14556 = ~n3433 & ~n14555;
  assign n14557 = ~i_hbusreq2 & ~n14556;
  assign n14558 = ~n9067 & ~n14557;
  assign n14559 = controllable_hgrant2 & ~n14558;
  assign n14560 = ~n3578 & ~n14559;
  assign n14561 = controllable_hmaster1 & ~n14560;
  assign n14562 = controllable_hmaster0 & ~n14560;
  assign n14563 = ~n3594 & ~n14506;
  assign n14564 = ~controllable_hmaster0 & ~n14563;
  assign n14565 = ~n14562 & ~n14564;
  assign n14566 = ~controllable_hmaster1 & ~n14565;
  assign n14567 = ~n14561 & ~n14566;
  assign n14568 = ~i_hbusreq3 & ~n14567;
  assign n14569 = ~n14545 & ~n14568;
  assign n14570 = controllable_hmaster2 & ~n14569;
  assign n14571 = controllable_hmaster0 & ~n14540;
  assign n14572 = ~n3547 & ~n6786;
  assign n14573 = ~controllable_hmaster0 & ~n14572;
  assign n14574 = ~n14571 & ~n14573;
  assign n14575 = controllable_hmaster1 & ~n14574;
  assign n14576 = ~controllable_hmaster1 & ~n14540;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = i_hbusreq3 & ~n14577;
  assign n14579 = controllable_hmaster0 & ~n14563;
  assign n14580 = ~n6813 & ~n11587;
  assign n14581 = ~controllable_hmaster0 & ~n14580;
  assign n14582 = ~n14579 & ~n14581;
  assign n14583 = controllable_hmaster1 & ~n14582;
  assign n14584 = ~controllable_hmaster1 & ~n14563;
  assign n14585 = ~n14583 & ~n14584;
  assign n14586 = ~i_hbusreq3 & ~n14585;
  assign n14587 = ~n14578 & ~n14586;
  assign n14588 = ~controllable_hmaster2 & ~n14587;
  assign n14589 = ~n14570 & ~n14588;
  assign n14590 = ~controllable_hgrant3 & ~n14589;
  assign n14591 = ~n14172 & ~n14590;
  assign n14592 = controllable_nhgrant0 & ~n14591;
  assign n14593 = ~n14180 & ~n14592;
  assign n14594 = ~n3281 & ~n14593;
  assign n14595 = ~n4089 & ~n14594;
  assign n14596 = ~n3378 & ~n14595;
  assign n14597 = ~n14536 & ~n14596;
  assign n14598 = n3492 & ~n14597;
  assign n14599 = ~n14433 & ~n14598;
  assign n14600 = n3485 & ~n14599;
  assign n14601 = ~n14432 & ~n14600;
  assign n14602 = n3476 & ~n14601;
  assign n14603 = ~n14484 & ~n14602;
  assign n14604 = n3374 & ~n14603;
  assign n14605 = ~n14439 & ~n14604;
  assign n14606 = n3655 & ~n14605;
  assign n14607 = ~controllable_hmaster0 & ~n9590;
  assign n14608 = controllable_hmaster1 & ~n14607;
  assign n14609 = controllable_hmaster1 & ~n14608;
  assign n14610 = i_hbusreq3 & ~n14609;
  assign n14611 = ~controllable_hmaster0 & ~n9603;
  assign n14612 = controllable_hmaster1 & ~n14611;
  assign n14613 = controllable_hmaster1 & ~n14612;
  assign n14614 = ~i_hbusreq3 & ~n14613;
  assign n14615 = ~n14610 & ~n14614;
  assign n14616 = ~controllable_hmaster2 & ~n14615;
  assign n14617 = ~controllable_hmaster2 & ~n14616;
  assign n14618 = ~controllable_hgrant3 & ~n14617;
  assign n14619 = ~n14140 & ~n14618;
  assign n14620 = controllable_nhgrant0 & ~n14619;
  assign n14621 = ~n14166 & ~n14620;
  assign n14622 = ~n3281 & ~n14621;
  assign n14623 = ~n3281 & ~n14622;
  assign n14624 = n3378 & ~n14623;
  assign n14625 = ~n14470 & ~n14616;
  assign n14626 = ~controllable_hgrant3 & ~n14625;
  assign n14627 = ~n14172 & ~n14626;
  assign n14628 = controllable_nhgrant0 & ~n14627;
  assign n14629 = ~n14180 & ~n14628;
  assign n14630 = ~n3281 & ~n14629;
  assign n14631 = ~n3950 & ~n14630;
  assign n14632 = ~n3378 & ~n14631;
  assign n14633 = ~n14624 & ~n14632;
  assign n14634 = n3492 & ~n14633;
  assign n14635 = ~n3493 & ~n14634;
  assign n14636 = n3485 & ~n14635;
  assign n14637 = ~n3486 & ~n14636;
  assign n14638 = ~n3476 & ~n14637;
  assign n14639 = ~n6786 & ~n9160;
  assign n14640 = ~controllable_hmaster0 & ~n14639;
  assign n14641 = ~n14511 & ~n14640;
  assign n14642 = controllable_hmaster1 & ~n14641;
  assign n14643 = ~n14516 & ~n14642;
  assign n14644 = i_hbusreq3 & ~n14643;
  assign n14645 = ~n6813 & ~n9184;
  assign n14646 = ~controllable_hmaster0 & ~n14645;
  assign n14647 = ~n14519 & ~n14646;
  assign n14648 = controllable_hmaster1 & ~n14647;
  assign n14649 = ~n14524 & ~n14648;
  assign n14650 = ~i_hbusreq3 & ~n14649;
  assign n14651 = ~n14644 & ~n14650;
  assign n14652 = ~controllable_hmaster2 & ~n14651;
  assign n14653 = ~n14510 & ~n14652;
  assign n14654 = ~controllable_hgrant3 & ~n14653;
  assign n14655 = ~n14140 & ~n14654;
  assign n14656 = controllable_nhgrant0 & ~n14655;
  assign n14657 = ~n14166 & ~n14656;
  assign n14658 = ~n3281 & ~n14657;
  assign n14659 = ~n3281 & ~n14658;
  assign n14660 = n3378 & ~n14659;
  assign n14661 = ~n6786 & ~n11654;
  assign n14662 = ~controllable_hmaster0 & ~n14661;
  assign n14663 = ~n14571 & ~n14662;
  assign n14664 = controllable_hmaster1 & ~n14663;
  assign n14665 = ~n14576 & ~n14664;
  assign n14666 = i_hbusreq3 & ~n14665;
  assign n14667 = ~n6813 & ~n11665;
  assign n14668 = ~controllable_hmaster0 & ~n14667;
  assign n14669 = ~n14579 & ~n14668;
  assign n14670 = controllable_hmaster1 & ~n14669;
  assign n14671 = ~n14584 & ~n14670;
  assign n14672 = ~i_hbusreq3 & ~n14671;
  assign n14673 = ~n14666 & ~n14672;
  assign n14674 = ~controllable_hmaster2 & ~n14673;
  assign n14675 = ~n14570 & ~n14674;
  assign n14676 = ~controllable_hgrant3 & ~n14675;
  assign n14677 = ~n14172 & ~n14676;
  assign n14678 = controllable_nhgrant0 & ~n14677;
  assign n14679 = ~n14180 & ~n14678;
  assign n14680 = ~n3281 & ~n14679;
  assign n14681 = ~n4089 & ~n14680;
  assign n14682 = ~n3378 & ~n14681;
  assign n14683 = ~n14660 & ~n14682;
  assign n14684 = n3492 & ~n14683;
  assign n14685 = ~n14433 & ~n14684;
  assign n14686 = n3485 & ~n14685;
  assign n14687 = ~n14432 & ~n14686;
  assign n14688 = n3476 & ~n14687;
  assign n14689 = ~n14638 & ~n14688;
  assign n14690 = n3374 & ~n14689;
  assign n14691 = ~n14439 & ~n14690;
  assign n14692 = ~n3655 & ~n14691;
  assign n14693 = ~n14606 & ~n14692;
  assign n14694 = ~n3652 & ~n14693;
  assign n14695 = ~n14369 & ~n14694;
  assign n14696 = ~n3368 & ~n14695;
  assign n14697 = controllable_hmaster1 & ~n4554;
  assign n14698 = controllable_hmaster1 & ~n14697;
  assign n14699 = ~i_hbusreq3 & ~n14698;
  assign n14700 = ~n14133 & ~n14699;
  assign n14701 = ~controllable_hmaster2 & ~n14700;
  assign n14702 = ~controllable_hmaster2 & ~n14701;
  assign n14703 = controllable_hgrant3 & ~n14702;
  assign n14704 = ~controllable_hmaster0 & ~n9805;
  assign n14705 = controllable_hmaster1 & ~n14704;
  assign n14706 = controllable_hmaster1 & ~n14705;
  assign n14707 = ~i_hbusreq3 & ~n14706;
  assign n14708 = ~n14144 & ~n14707;
  assign n14709 = ~controllable_hmaster2 & ~n14708;
  assign n14710 = ~controllable_hmaster2 & ~n14709;
  assign n14711 = ~controllable_hgrant3 & ~n14710;
  assign n14712 = ~n14703 & ~n14711;
  assign n14713 = controllable_nhgrant0 & ~n14712;
  assign n14714 = controllable_hmaster1 & ~n4612;
  assign n14715 = controllable_hmaster1 & ~n14714;
  assign n14716 = i_hbusreq3 & ~n14715;
  assign n14717 = controllable_hmaster1 & ~n4637;
  assign n14718 = controllable_hmaster1 & ~n14717;
  assign n14719 = ~i_hbusreq3 & ~n14718;
  assign n14720 = ~n14716 & ~n14719;
  assign n14721 = ~controllable_hmaster2 & ~n14720;
  assign n14722 = ~controllable_hmaster2 & ~n14721;
  assign n14723 = ~controllable_hgrant3 & ~n14722;
  assign n14724 = ~n14703 & ~n14723;
  assign n14725 = ~controllable_nhgrant0 & ~n14724;
  assign n14726 = ~n14713 & ~n14725;
  assign n14727 = ~n3281 & ~n14726;
  assign n14728 = ~n3281 & ~n14727;
  assign n14729 = n3492 & ~n14728;
  assign n14730 = n3492 & ~n14729;
  assign n14731 = n3485 & ~n14730;
  assign n14732 = n3485 & ~n14731;
  assign n14733 = ~n3476 & ~n14732;
  assign n14734 = controllable_hmaster2 & ~n14192;
  assign n14735 = ~n9800 & ~n10152;
  assign n14736 = ~controllable_hmaster0 & ~n14735;
  assign n14737 = ~n14199 & ~n14736;
  assign n14738 = controllable_hmaster1 & ~n14737;
  assign n14739 = ~n14204 & ~n14738;
  assign n14740 = ~i_hbusreq3 & ~n14739;
  assign n14741 = ~n14206 & ~n14740;
  assign n14742 = ~controllable_hmaster2 & ~n14741;
  assign n14743 = ~n14734 & ~n14742;
  assign n14744 = ~controllable_hgrant3 & ~n14743;
  assign n14745 = ~n14703 & ~n14744;
  assign n14746 = controllable_nhgrant0 & ~n14745;
  assign n14747 = ~n14725 & ~n14746;
  assign n14748 = ~n3281 & ~n14747;
  assign n14749 = ~n3281 & ~n14748;
  assign n14750 = n3492 & ~n14749;
  assign n14751 = n3492 & ~n14750;
  assign n14752 = n3485 & ~n14751;
  assign n14753 = n3485 & ~n14752;
  assign n14754 = n3476 & ~n14753;
  assign n14755 = ~n14733 & ~n14754;
  assign n14756 = n3374 & ~n14755;
  assign n14757 = n3374 & ~n14756;
  assign n14758 = n3655 & ~n14757;
  assign n14759 = ~controllable_hmaster0 & ~n10328;
  assign n14760 = controllable_hmaster1 & ~n14759;
  assign n14761 = controllable_hmaster1 & ~n14760;
  assign n14762 = i_hbusreq3 & ~n14761;
  assign n14763 = ~controllable_hmaster0 & ~n10350;
  assign n14764 = controllable_hmaster1 & ~n14763;
  assign n14765 = controllable_hmaster1 & ~n14764;
  assign n14766 = ~i_hbusreq3 & ~n14765;
  assign n14767 = ~n14762 & ~n14766;
  assign n14768 = ~controllable_hmaster2 & ~n14767;
  assign n14769 = ~controllable_hmaster2 & ~n14768;
  assign n14770 = ~controllable_hgrant3 & ~n14769;
  assign n14771 = ~n14703 & ~n14770;
  assign n14772 = controllable_nhgrant0 & ~n14771;
  assign n14773 = ~n14725 & ~n14772;
  assign n14774 = ~n3281 & ~n14773;
  assign n14775 = ~n3281 & ~n14774;
  assign n14776 = n3492 & ~n14775;
  assign n14777 = n3492 & ~n14776;
  assign n14778 = n3485 & ~n14777;
  assign n14779 = n3485 & ~n14778;
  assign n14780 = ~n3476 & ~n14779;
  assign n14781 = ~n5686 & ~n10324;
  assign n14782 = ~controllable_hmaster0 & ~n14781;
  assign n14783 = ~n14199 & ~n14782;
  assign n14784 = controllable_hmaster1 & ~n14783;
  assign n14785 = ~n14204 & ~n14784;
  assign n14786 = i_hbusreq3 & ~n14785;
  assign n14787 = ~n10152 & ~n10346;
  assign n14788 = ~controllable_hmaster0 & ~n14787;
  assign n14789 = ~n14199 & ~n14788;
  assign n14790 = controllable_hmaster1 & ~n14789;
  assign n14791 = ~n14204 & ~n14790;
  assign n14792 = ~i_hbusreq3 & ~n14791;
  assign n14793 = ~n14786 & ~n14792;
  assign n14794 = ~controllable_hmaster2 & ~n14793;
  assign n14795 = ~n14734 & ~n14794;
  assign n14796 = ~controllable_hgrant3 & ~n14795;
  assign n14797 = ~n14703 & ~n14796;
  assign n14798 = controllable_nhgrant0 & ~n14797;
  assign n14799 = ~n14725 & ~n14798;
  assign n14800 = ~n3281 & ~n14799;
  assign n14801 = ~n3281 & ~n14800;
  assign n14802 = n3492 & ~n14801;
  assign n14803 = n3492 & ~n14802;
  assign n14804 = n3485 & ~n14803;
  assign n14805 = n3485 & ~n14804;
  assign n14806 = n3476 & ~n14805;
  assign n14807 = ~n14780 & ~n14806;
  assign n14808 = n3374 & ~n14807;
  assign n14809 = n3374 & ~n14808;
  assign n14810 = ~n3655 & ~n14809;
  assign n14811 = ~n14758 & ~n14810;
  assign n14812 = n3652 & ~n14811;
  assign n14813 = ~controllable_hmaster0 & ~n10770;
  assign n14814 = controllable_hmaster1 & ~n14813;
  assign n14815 = controllable_hmaster1 & ~n14814;
  assign n14816 = i_hbusreq3 & ~n14815;
  assign n14817 = ~controllable_hmaster0 & ~n10784;
  assign n14818 = controllable_hmaster1 & ~n14817;
  assign n14819 = controllable_hmaster1 & ~n14818;
  assign n14820 = ~i_hbusreq3 & ~n14819;
  assign n14821 = ~n14816 & ~n14820;
  assign n14822 = ~controllable_hmaster2 & ~n14821;
  assign n14823 = ~controllable_hmaster2 & ~n14822;
  assign n14824 = ~controllable_hgrant3 & ~n14823;
  assign n14825 = ~n14703 & ~n14824;
  assign n14826 = controllable_nhgrant0 & ~n14825;
  assign n14827 = ~n14725 & ~n14826;
  assign n14828 = ~n3281 & ~n14827;
  assign n14829 = ~n3281 & ~n14828;
  assign n14830 = n3492 & ~n14829;
  assign n14831 = n3492 & ~n14830;
  assign n14832 = n3485 & ~n14831;
  assign n14833 = n3485 & ~n14832;
  assign n14834 = ~n3476 & ~n14833;
  assign n14835 = ~n3485 & ~n14382;
  assign n14836 = ~n3492 & ~n14382;
  assign n14837 = i_hlock2 & ~n3553;
  assign n14838 = i_hready & ~n9958;
  assign n14839 = ~controllable_hgrant4 & ~n14838;
  assign n14840 = ~controllable_hgrant4 & ~n14839;
  assign n14841 = ~i_hlock2 & ~n14840;
  assign n14842 = ~n14837 & ~n14841;
  assign n14843 = controllable_hgrant2 & ~n14842;
  assign n14844 = controllable_hgrant2 & ~n14843;
  assign n14845 = i_hbusreq3 & ~n14844;
  assign n14846 = i_hbusreq2 & ~n14842;
  assign n14847 = i_hready & ~n10842;
  assign n14848 = ~i_hbusreq0 & ~n14847;
  assign n14849 = ~n3584 & ~n14848;
  assign n14850 = ~i_hbusreq4 & ~n14849;
  assign n14851 = ~n3583 & ~n14850;
  assign n14852 = ~controllable_hgrant4 & ~n14851;
  assign n14853 = ~controllable_hgrant4 & ~n14852;
  assign n14854 = i_hlock2 & ~n14853;
  assign n14855 = ~n14841 & ~n14854;
  assign n14856 = ~i_hbusreq2 & ~n14855;
  assign n14857 = ~n14846 & ~n14856;
  assign n14858 = controllable_hgrant2 & ~n14857;
  assign n14859 = controllable_hgrant2 & ~n14858;
  assign n14860 = ~i_hbusreq3 & ~n14859;
  assign n14861 = ~n14845 & ~n14860;
  assign n14862 = controllable_hmaster2 & ~n14861;
  assign n14863 = controllable_hmaster0 & ~n14844;
  assign n14864 = ~n8768 & ~n11066;
  assign n14865 = ~controllable_hmaster0 & ~n14864;
  assign n14866 = ~n14863 & ~n14865;
  assign n14867 = controllable_hmaster1 & ~n14866;
  assign n14868 = ~controllable_hmaster1 & ~n14844;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = i_hbusreq3 & ~n14869;
  assign n14871 = controllable_hmaster0 & ~n14859;
  assign n14872 = ~n9800 & ~n11110;
  assign n14873 = ~controllable_hmaster0 & ~n14872;
  assign n14874 = ~n14871 & ~n14873;
  assign n14875 = controllable_hmaster1 & ~n14874;
  assign n14876 = ~controllable_hmaster1 & ~n14859;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = ~i_hbusreq3 & ~n14877;
  assign n14879 = ~n14870 & ~n14878;
  assign n14880 = ~controllable_hmaster2 & ~n14879;
  assign n14881 = ~n14862 & ~n14880;
  assign n14882 = ~controllable_hgrant3 & ~n14881;
  assign n14883 = ~n14703 & ~n14882;
  assign n14884 = controllable_nhgrant0 & ~n14883;
  assign n14885 = ~n14725 & ~n14884;
  assign n14886 = ~n3281 & ~n14885;
  assign n14887 = ~n3281 & ~n14886;
  assign n14888 = n3492 & ~n14887;
  assign n14889 = ~n14836 & ~n14888;
  assign n14890 = n3485 & ~n14889;
  assign n14891 = ~n14835 & ~n14890;
  assign n14892 = n3476 & ~n14891;
  assign n14893 = ~n14834 & ~n14892;
  assign n14894 = n3374 & ~n14893;
  assign n14895 = n3374 & ~n14894;
  assign n14896 = n3655 & ~n14895;
  assign n14897 = ~controllable_hmaster0 & ~n11205;
  assign n14898 = controllable_hmaster1 & ~n14897;
  assign n14899 = controllable_hmaster1 & ~n14898;
  assign n14900 = i_hbusreq3 & ~n14899;
  assign n14901 = ~controllable_hmaster0 & ~n11218;
  assign n14902 = controllable_hmaster1 & ~n14901;
  assign n14903 = controllable_hmaster1 & ~n14902;
  assign n14904 = ~i_hbusreq3 & ~n14903;
  assign n14905 = ~n14900 & ~n14904;
  assign n14906 = ~controllable_hmaster2 & ~n14905;
  assign n14907 = ~controllable_hmaster2 & ~n14906;
  assign n14908 = ~controllable_hgrant3 & ~n14907;
  assign n14909 = ~n14703 & ~n14908;
  assign n14910 = controllable_nhgrant0 & ~n14909;
  assign n14911 = ~n14725 & ~n14910;
  assign n14912 = ~n3281 & ~n14911;
  assign n14913 = ~n3281 & ~n14912;
  assign n14914 = n3492 & ~n14913;
  assign n14915 = n3492 & ~n14914;
  assign n14916 = n3485 & ~n14915;
  assign n14917 = n3485 & ~n14916;
  assign n14918 = ~n3476 & ~n14917;
  assign n14919 = ~n10324 & ~n11066;
  assign n14920 = ~controllable_hmaster0 & ~n14919;
  assign n14921 = ~n14863 & ~n14920;
  assign n14922 = controllable_hmaster1 & ~n14921;
  assign n14923 = ~n14868 & ~n14922;
  assign n14924 = i_hbusreq3 & ~n14923;
  assign n14925 = ~n10346 & ~n11110;
  assign n14926 = ~controllable_hmaster0 & ~n14925;
  assign n14927 = ~n14871 & ~n14926;
  assign n14928 = controllable_hmaster1 & ~n14927;
  assign n14929 = ~n14876 & ~n14928;
  assign n14930 = ~i_hbusreq3 & ~n14929;
  assign n14931 = ~n14924 & ~n14930;
  assign n14932 = ~controllable_hmaster2 & ~n14931;
  assign n14933 = ~n14862 & ~n14932;
  assign n14934 = ~controllable_hgrant3 & ~n14933;
  assign n14935 = ~n14703 & ~n14934;
  assign n14936 = controllable_nhgrant0 & ~n14935;
  assign n14937 = ~n14725 & ~n14936;
  assign n14938 = ~n3281 & ~n14937;
  assign n14939 = ~n3281 & ~n14938;
  assign n14940 = n3492 & ~n14939;
  assign n14941 = ~n14836 & ~n14940;
  assign n14942 = n3485 & ~n14941;
  assign n14943 = ~n14835 & ~n14942;
  assign n14944 = n3476 & ~n14943;
  assign n14945 = ~n14918 & ~n14944;
  assign n14946 = n3374 & ~n14945;
  assign n14947 = n3374 & ~n14946;
  assign n14948 = ~n3655 & ~n14947;
  assign n14949 = ~n14896 & ~n14948;
  assign n14950 = ~n3652 & ~n14949;
  assign n14951 = ~n14812 & ~n14950;
  assign n14952 = n3368 & ~n14951;
  assign n14953 = ~n14696 & ~n14952;
  assign n14954 = ~n3362 & ~n14953;
  assign n14955 = ~n3362 & ~n14954;
  assign n14956 = ~n3359 & ~n14955;
  assign n14957 = ~n3359 & ~n14956;
  assign n14958 = n3356 & ~n14957;
  assign n14959 = n3378 & ~n14123;
  assign n14960 = ~n5249 & ~n14959;
  assign n14961 = n3492 & ~n14960;
  assign n14962 = ~n3631 & ~n14961;
  assign n14963 = n3485 & ~n14962;
  assign n14964 = ~n3630 & ~n14963;
  assign n14965 = ~n3374 & ~n14964;
  assign n14966 = ~n3835 & ~n5277;
  assign n14967 = controllable_hmaster1 & ~n14966;
  assign n14968 = ~n5281 & ~n14967;
  assign n14969 = ~i_hbusreq3 & ~n14968;
  assign n14970 = ~n5265 & ~n14969;
  assign n14971 = ~controllable_hmaster2 & ~n14970;
  assign n14972 = ~n12033 & ~n14971;
  assign n14973 = controllable_hgrant3 & ~n14972;
  assign n14974 = ~n3382 & ~n8818;
  assign n14975 = controllable_hmaster1 & ~n14974;
  assign n14976 = ~n5305 & ~n14975;
  assign n14977 = i_hbusreq3 & ~n14976;
  assign n14978 = ~n3401 & ~n8840;
  assign n14979 = controllable_hmaster1 & ~n14978;
  assign n14980 = ~n5334 & ~n14979;
  assign n14981 = ~i_hbusreq3 & ~n14980;
  assign n14982 = ~n14977 & ~n14981;
  assign n14983 = ~controllable_hmaster2 & ~n14982;
  assign n14984 = ~n12065 & ~n14983;
  assign n14985 = ~controllable_hgrant3 & ~n14984;
  assign n14986 = ~n14973 & ~n14985;
  assign n14987 = controllable_nhgrant0 & ~n14986;
  assign n14988 = controllable_hmaster1 & ~n3952;
  assign n14989 = ~n5281 & ~n14988;
  assign n14990 = ~i_hbusreq3 & ~n14989;
  assign n14991 = ~n3951 & ~n14990;
  assign n14992 = ~controllable_hmaster2 & ~n14991;
  assign n14993 = ~n12033 & ~n14992;
  assign n14994 = controllable_hgrant3 & ~n14993;
  assign n14995 = controllable_hmaster1 & ~n3974;
  assign n14996 = ~n5350 & ~n14995;
  assign n14997 = i_hbusreq3 & ~n14996;
  assign n14998 = controllable_hmaster1 & ~n3978;
  assign n14999 = ~n5355 & ~n14998;
  assign n15000 = ~i_hbusreq3 & ~n14999;
  assign n15001 = ~n14997 & ~n15000;
  assign n15002 = ~controllable_hmaster2 & ~n15001;
  assign n15003 = ~n12033 & ~n15002;
  assign n15004 = ~controllable_hgrant3 & ~n15003;
  assign n15005 = ~n14994 & ~n15004;
  assign n15006 = ~controllable_nhgrant0 & ~n15005;
  assign n15007 = ~n14987 & ~n15006;
  assign n15008 = ~n3281 & ~n15007;
  assign n15009 = ~n3950 & ~n15008;
  assign n15010 = n3378 & ~n15009;
  assign n15011 = ~n5191 & ~n8818;
  assign n15012 = controllable_hmaster1 & ~n15011;
  assign n15013 = ~n5435 & ~n15012;
  assign n15014 = i_hbusreq3 & ~n15013;
  assign n15015 = ~n5197 & ~n8840;
  assign n15016 = controllable_hmaster1 & ~n15015;
  assign n15017 = ~n5480 & ~n15016;
  assign n15018 = ~i_hbusreq3 & ~n15017;
  assign n15019 = ~n15014 & ~n15018;
  assign n15020 = ~controllable_hmaster2 & ~n15019;
  assign n15021 = ~n12126 & ~n15020;
  assign n15022 = ~controllable_hgrant3 & ~n15021;
  assign n15023 = ~n5402 & ~n15022;
  assign n15024 = controllable_nhgrant0 & ~n15023;
  assign n15025 = ~n5534 & ~n15024;
  assign n15026 = ~n3281 & ~n15025;
  assign n15027 = ~n3950 & ~n15026;
  assign n15028 = ~n3378 & ~n15027;
  assign n15029 = ~n15010 & ~n15028;
  assign n15030 = n3492 & ~n15029;
  assign n15031 = ~n3631 & ~n15030;
  assign n15032 = n3485 & ~n15031;
  assign n15033 = ~n3630 & ~n15032;
  assign n15034 = ~n3476 & ~n15033;
  assign n15035 = ~n5576 & ~n5605;
  assign n15036 = controllable_hmaster1 & ~n15035;
  assign n15037 = ~n5609 & ~n15036;
  assign n15038 = ~i_hbusreq3 & ~n15037;
  assign n15039 = ~n5593 & ~n15038;
  assign n15040 = ~controllable_hmaster2 & ~n15039;
  assign n15041 = ~n12233 & ~n15040;
  assign n15042 = controllable_hgrant3 & ~n15041;
  assign n15043 = ~n12176 & ~n14234;
  assign n15044 = controllable_hmaster1 & ~n15043;
  assign n15045 = controllable_hmaster0 & ~n15043;
  assign n15046 = ~n12185 & ~n14234;
  assign n15047 = ~controllable_hmaster0 & ~n15046;
  assign n15048 = ~n15045 & ~n15047;
  assign n15049 = ~controllable_hmaster1 & ~n15048;
  assign n15050 = ~n15044 & ~n15049;
  assign n15051 = ~i_hbusreq3 & ~n15050;
  assign n15052 = ~n12171 & ~n15051;
  assign n15053 = controllable_hmaster2 & ~n15052;
  assign n15054 = ~n5685 & ~n8983;
  assign n15055 = controllable_hmaster1 & ~n15054;
  assign n15056 = ~n5704 & ~n15055;
  assign n15057 = i_hbusreq3 & ~n15056;
  assign n15058 = ~n12208 & ~n14234;
  assign n15059 = controllable_hmaster0 & ~n15058;
  assign n15060 = ~n5950 & ~n12202;
  assign n15061 = ~controllable_hmaster0 & ~n15060;
  assign n15062 = ~n15059 & ~n15061;
  assign n15063 = controllable_hmaster1 & ~n15062;
  assign n15064 = ~n12216 & ~n14234;
  assign n15065 = controllable_hmaster0 & ~n15064;
  assign n15066 = ~controllable_hmaster0 & ~n15058;
  assign n15067 = ~n15065 & ~n15066;
  assign n15068 = ~controllable_hmaster1 & ~n15067;
  assign n15069 = ~n15063 & ~n15068;
  assign n15070 = ~i_hbusreq3 & ~n15069;
  assign n15071 = ~n15057 & ~n15070;
  assign n15072 = ~controllable_hmaster2 & ~n15071;
  assign n15073 = ~n15053 & ~n15072;
  assign n15074 = ~controllable_hgrant3 & ~n15073;
  assign n15075 = ~n15042 & ~n15074;
  assign n15076 = controllable_nhgrant0 & ~n15075;
  assign n15077 = controllable_hmaster1 & ~n5765;
  assign n15078 = ~n5796 & ~n15077;
  assign n15079 = i_hbusreq3 & ~n15078;
  assign n15080 = controllable_hmaster1 & ~n5788;
  assign n15081 = ~n5801 & ~n15080;
  assign n15082 = ~i_hbusreq3 & ~n15081;
  assign n15083 = ~n15079 & ~n15082;
  assign n15084 = ~controllable_hmaster2 & ~n15083;
  assign n15085 = ~n12233 & ~n15084;
  assign n15086 = ~controllable_hgrant3 & ~n15085;
  assign n15087 = ~n14994 & ~n15086;
  assign n15088 = ~controllable_nhgrant0 & ~n15087;
  assign n15089 = ~n15076 & ~n15088;
  assign n15090 = ~n3281 & ~n15089;
  assign n15091 = ~n4089 & ~n15090;
  assign n15092 = n3378 & ~n15091;
  assign n15093 = ~n5915 & ~n8983;
  assign n15094 = controllable_hmaster1 & ~n15093;
  assign n15095 = ~n5928 & ~n15094;
  assign n15096 = i_hbusreq3 & ~n15095;
  assign n15097 = ~n5950 & ~n12282;
  assign n15098 = ~controllable_hmaster0 & ~n15097;
  assign n15099 = ~n5949 & ~n15098;
  assign n15100 = controllable_hmaster1 & ~n15099;
  assign n15101 = ~n5998 & ~n15100;
  assign n15102 = ~i_hbusreq3 & ~n15101;
  assign n15103 = ~n15096 & ~n15102;
  assign n15104 = ~controllable_hmaster2 & ~n15103;
  assign n15105 = ~n12274 & ~n15104;
  assign n15106 = ~controllable_hgrant3 & ~n15105;
  assign n15107 = ~n5861 & ~n15106;
  assign n15108 = controllable_nhgrant0 & ~n15107;
  assign n15109 = ~n6082 & ~n15108;
  assign n15110 = ~n3281 & ~n15109;
  assign n15111 = ~n4089 & ~n15110;
  assign n15112 = ~n3378 & ~n15111;
  assign n15113 = ~n15092 & ~n15112;
  assign n15114 = n3492 & ~n15113;
  assign n15115 = ~n3631 & ~n15114;
  assign n15116 = n3485 & ~n15115;
  assign n15117 = ~n3630 & ~n15116;
  assign n15118 = n3476 & ~n15117;
  assign n15119 = ~n15034 & ~n15118;
  assign n15120 = n3374 & ~n15119;
  assign n15121 = ~n14965 & ~n15120;
  assign n15122 = n3655 & ~n15121;
  assign n15123 = ~n6196 & ~n14959;
  assign n15124 = n3492 & ~n15123;
  assign n15125 = ~n3631 & ~n15124;
  assign n15126 = n3485 & ~n15125;
  assign n15127 = ~n3630 & ~n15126;
  assign n15128 = ~n3374 & ~n15127;
  assign n15129 = ~n3382 & ~n9164;
  assign n15130 = controllable_hmaster1 & ~n15129;
  assign n15131 = ~n5305 & ~n15130;
  assign n15132 = i_hbusreq3 & ~n15131;
  assign n15133 = ~n3401 & ~n9188;
  assign n15134 = controllable_hmaster1 & ~n15133;
  assign n15135 = ~n5334 & ~n15134;
  assign n15136 = ~i_hbusreq3 & ~n15135;
  assign n15137 = ~n15132 & ~n15136;
  assign n15138 = ~controllable_hmaster2 & ~n15137;
  assign n15139 = ~n12065 & ~n15138;
  assign n15140 = ~controllable_hgrant3 & ~n15139;
  assign n15141 = ~n14973 & ~n15140;
  assign n15142 = controllable_nhgrant0 & ~n15141;
  assign n15143 = ~n15006 & ~n15142;
  assign n15144 = ~n3281 & ~n15143;
  assign n15145 = ~n3950 & ~n15144;
  assign n15146 = n3378 & ~n15145;
  assign n15147 = ~n6254 & ~n9164;
  assign n15148 = controllable_hmaster1 & ~n15147;
  assign n15149 = ~n6271 & ~n15148;
  assign n15150 = i_hbusreq3 & ~n15149;
  assign n15151 = ~n6293 & ~n9188;
  assign n15152 = controllable_hmaster1 & ~n15151;
  assign n15153 = ~n6339 & ~n15152;
  assign n15154 = ~i_hbusreq3 & ~n15153;
  assign n15155 = ~n15150 & ~n15154;
  assign n15156 = ~controllable_hmaster2 & ~n15155;
  assign n15157 = ~n12353 & ~n15156;
  assign n15158 = ~controllable_hgrant3 & ~n15157;
  assign n15159 = ~n5402 & ~n15158;
  assign n15160 = controllable_nhgrant0 & ~n15159;
  assign n15161 = ~n5534 & ~n15160;
  assign n15162 = ~n3281 & ~n15161;
  assign n15163 = ~n3950 & ~n15162;
  assign n15164 = ~n3378 & ~n15163;
  assign n15165 = ~n15146 & ~n15164;
  assign n15166 = n3492 & ~n15165;
  assign n15167 = ~n3631 & ~n15166;
  assign n15168 = n3485 & ~n15167;
  assign n15169 = ~n3630 & ~n15168;
  assign n15170 = ~n3476 & ~n15169;
  assign n15171 = ~n5686 & ~n12379;
  assign n15172 = ~controllable_hmaster0 & ~n15171;
  assign n15173 = ~n5685 & ~n15172;
  assign n15174 = controllable_hmaster1 & ~n15173;
  assign n15175 = ~n5704 & ~n15174;
  assign n15176 = i_hbusreq3 & ~n15175;
  assign n15177 = ~n5950 & ~n12390;
  assign n15178 = ~controllable_hmaster0 & ~n15177;
  assign n15179 = ~n15059 & ~n15178;
  assign n15180 = controllable_hmaster1 & ~n15179;
  assign n15181 = ~n15068 & ~n15180;
  assign n15182 = ~i_hbusreq3 & ~n15181;
  assign n15183 = ~n15176 & ~n15182;
  assign n15184 = ~controllable_hmaster2 & ~n15183;
  assign n15185 = ~n15053 & ~n15184;
  assign n15186 = ~controllable_hgrant3 & ~n15185;
  assign n15187 = ~n15042 & ~n15186;
  assign n15188 = controllable_nhgrant0 & ~n15187;
  assign n15189 = ~n15088 & ~n15188;
  assign n15190 = ~n3281 & ~n15189;
  assign n15191 = ~n4089 & ~n15190;
  assign n15192 = n3378 & ~n15191;
  assign n15193 = ~n6469 & ~n9301;
  assign n15194 = controllable_hmaster1 & ~n15193;
  assign n15195 = ~n6483 & ~n15194;
  assign n15196 = i_hbusreq3 & ~n15195;
  assign n15197 = ~n5950 & ~n12435;
  assign n15198 = ~controllable_hmaster0 & ~n15197;
  assign n15199 = ~n6504 & ~n15198;
  assign n15200 = controllable_hmaster1 & ~n15199;
  assign n15201 = ~n6550 & ~n15200;
  assign n15202 = ~i_hbusreq3 & ~n15201;
  assign n15203 = ~n15196 & ~n15202;
  assign n15204 = ~controllable_hmaster2 & ~n15203;
  assign n15205 = ~n12427 & ~n15204;
  assign n15206 = ~controllable_hgrant3 & ~n15205;
  assign n15207 = ~n5861 & ~n15206;
  assign n15208 = controllable_nhgrant0 & ~n15207;
  assign n15209 = ~n6082 & ~n15208;
  assign n15210 = ~n3281 & ~n15209;
  assign n15211 = ~n4089 & ~n15210;
  assign n15212 = ~n3378 & ~n15211;
  assign n15213 = ~n15192 & ~n15212;
  assign n15214 = n3492 & ~n15213;
  assign n15215 = ~n3631 & ~n15214;
  assign n15216 = n3485 & ~n15215;
  assign n15217 = ~n3630 & ~n15216;
  assign n15218 = n3476 & ~n15217;
  assign n15219 = ~n15170 & ~n15218;
  assign n15220 = n3374 & ~n15219;
  assign n15221 = ~n15128 & ~n15220;
  assign n15222 = ~n3655 & ~n15221;
  assign n15223 = ~n15122 & ~n15222;
  assign n15224 = n3652 & ~n15223;
  assign n15225 = n3378 & ~n14415;
  assign n15226 = ~n5043 & ~n9388;
  assign n15227 = controllable_hmaster1 & ~n15226;
  assign n15228 = controllable_hmaster0 & ~n15226;
  assign n15229 = ~n3729 & ~n15228;
  assign n15230 = ~controllable_hmaster1 & ~n15229;
  assign n15231 = ~n15227 & ~n15230;
  assign n15232 = i_hbusreq3 & ~n15231;
  assign n15233 = controllable_hgrant2 & ~n8835;
  assign n15234 = ~n5068 & ~n15233;
  assign n15235 = controllable_hmaster1 & ~n15234;
  assign n15236 = controllable_hmaster0 & ~n15234;
  assign n15237 = ~n3767 & ~n15236;
  assign n15238 = ~controllable_hmaster1 & ~n15237;
  assign n15239 = ~n15235 & ~n15238;
  assign n15240 = ~i_hbusreq3 & ~n15239;
  assign n15241 = ~n15232 & ~n15240;
  assign n15242 = controllable_hmaster2 & ~n15241;
  assign n15243 = ~n6657 & ~n15242;
  assign n15244 = ~controllable_hgrant3 & ~n15243;
  assign n15245 = ~n5037 & ~n15244;
  assign n15246 = controllable_nhgrant0 & ~n15245;
  assign n15247 = ~n5245 & ~n15246;
  assign n15248 = ~n3281 & ~n15247;
  assign n15249 = ~n3783 & ~n15248;
  assign n15250 = ~n3378 & ~n15249;
  assign n15251 = ~n15225 & ~n15250;
  assign n15252 = n3492 & ~n15251;
  assign n15253 = ~n3631 & ~n15252;
  assign n15254 = n3485 & ~n15253;
  assign n15255 = ~n3630 & ~n15254;
  assign n15256 = ~n3476 & ~n15255;
  assign n15257 = ~n3485 & ~n14429;
  assign n15258 = ~n3492 & ~n14429;
  assign n15259 = ~n15252 & ~n15258;
  assign n15260 = n3485 & ~n15259;
  assign n15261 = ~n15257 & ~n15260;
  assign n15262 = n3476 & ~n15261;
  assign n15263 = ~n15256 & ~n15262;
  assign n15264 = ~n3374 & ~n15263;
  assign n15265 = ~n4333 & ~n12044;
  assign n15266 = ~controllable_hmaster0 & ~n15265;
  assign n15267 = ~n9391 & ~n15266;
  assign n15268 = ~controllable_hmaster1 & ~n15267;
  assign n15269 = ~n9390 & ~n15268;
  assign n15270 = i_hbusreq3 & ~n15269;
  assign n15271 = ~i_hbusreq0 & ~n3921;
  assign n15272 = ~n3918 & ~n15271;
  assign n15273 = ~i_hbusreq4 & ~n15272;
  assign n15274 = ~n3917 & ~n15273;
  assign n15275 = ~controllable_hgrant4 & ~n15274;
  assign n15276 = ~n3433 & ~n15275;
  assign n15277 = ~i_hbusreq2 & ~n15276;
  assign n15278 = ~n3915 & ~n15277;
  assign n15279 = controllable_hgrant2 & ~n15278;
  assign n15280 = ~n12057 & ~n15279;
  assign n15281 = ~controllable_hmaster0 & ~n15280;
  assign n15282 = ~n14464 & ~n15281;
  assign n15283 = ~controllable_hmaster1 & ~n15282;
  assign n15284 = ~n14463 & ~n15283;
  assign n15285 = ~i_hbusreq3 & ~n15284;
  assign n15286 = ~n15270 & ~n15285;
  assign n15287 = controllable_hmaster2 & ~n15286;
  assign n15288 = ~n4333 & ~n5289;
  assign n15289 = controllable_hmaster0 & ~n15288;
  assign n15290 = ~n9436 & ~n15289;
  assign n15291 = controllable_hmaster1 & ~n15290;
  assign n15292 = ~n4333 & ~n5301;
  assign n15293 = controllable_hmaster0 & ~n15292;
  assign n15294 = ~controllable_hmaster0 & ~n15288;
  assign n15295 = ~n15293 & ~n15294;
  assign n15296 = ~controllable_hmaster1 & ~n15295;
  assign n15297 = ~n15291 & ~n15296;
  assign n15298 = i_hbusreq3 & ~n15297;
  assign n15299 = ~n5309 & ~n15279;
  assign n15300 = controllable_hmaster0 & ~n15299;
  assign n15301 = ~n9449 & ~n15300;
  assign n15302 = controllable_hmaster1 & ~n15301;
  assign n15303 = ~n5330 & ~n15279;
  assign n15304 = controllable_hmaster0 & ~n15303;
  assign n15305 = ~controllable_hmaster0 & ~n15299;
  assign n15306 = ~n15304 & ~n15305;
  assign n15307 = ~controllable_hmaster1 & ~n15306;
  assign n15308 = ~n15302 & ~n15307;
  assign n15309 = ~i_hbusreq3 & ~n15308;
  assign n15310 = ~n15298 & ~n15309;
  assign n15311 = ~controllable_hmaster2 & ~n15310;
  assign n15312 = ~n15287 & ~n15311;
  assign n15313 = ~controllable_hgrant3 & ~n15312;
  assign n15314 = ~n14973 & ~n15313;
  assign n15315 = controllable_nhgrant0 & ~n15314;
  assign n15316 = ~n15006 & ~n15315;
  assign n15317 = ~n3281 & ~n15316;
  assign n15318 = ~n3950 & ~n15317;
  assign n15319 = n3378 & ~n15318;
  assign n15320 = ~n9391 & ~n12489;
  assign n15321 = ~controllable_hmaster1 & ~n15320;
  assign n15322 = ~n9390 & ~n15321;
  assign n15323 = i_hbusreq3 & ~n15322;
  assign n15324 = ~n5414 & ~n15233;
  assign n15325 = controllable_hmaster1 & ~n15324;
  assign n15326 = controllable_hmaster0 & ~n15324;
  assign n15327 = ~n12495 & ~n15326;
  assign n15328 = ~controllable_hmaster1 & ~n15327;
  assign n15329 = ~n15325 & ~n15328;
  assign n15330 = ~i_hbusreq3 & ~n15329;
  assign n15331 = ~n15323 & ~n15330;
  assign n15332 = controllable_hmaster2 & ~n15331;
  assign n15333 = ~n6696 & ~n9436;
  assign n15334 = controllable_hmaster1 & ~n15333;
  assign n15335 = ~n6706 & ~n15334;
  assign n15336 = i_hbusreq3 & ~n15335;
  assign n15337 = ~n6709 & ~n9449;
  assign n15338 = controllable_hmaster1 & ~n15337;
  assign n15339 = ~n6719 & ~n15338;
  assign n15340 = ~i_hbusreq3 & ~n15339;
  assign n15341 = ~n15336 & ~n15340;
  assign n15342 = ~controllable_hmaster2 & ~n15341;
  assign n15343 = ~n15332 & ~n15342;
  assign n15344 = ~controllable_hgrant3 & ~n15343;
  assign n15345 = ~n5402 & ~n15344;
  assign n15346 = controllable_nhgrant0 & ~n15345;
  assign n15347 = ~n5534 & ~n15346;
  assign n15348 = ~n3281 & ~n15347;
  assign n15349 = ~n3950 & ~n15348;
  assign n15350 = ~n3378 & ~n15349;
  assign n15351 = ~n15319 & ~n15350;
  assign n15352 = n3492 & ~n15351;
  assign n15353 = ~n3631 & ~n15352;
  assign n15354 = n3485 & ~n15353;
  assign n15355 = ~n3630 & ~n15354;
  assign n15356 = ~n3476 & ~n15355;
  assign n15357 = ~n6762 & ~n12165;
  assign n15358 = ~controllable_hmaster0 & ~n15357;
  assign n15359 = ~n9480 & ~n15358;
  assign n15360 = ~controllable_hmaster1 & ~n15359;
  assign n15361 = ~n9479 & ~n15360;
  assign n15362 = i_hbusreq3 & ~n15361;
  assign n15363 = ~n12176 & ~n14559;
  assign n15364 = controllable_hmaster1 & ~n15363;
  assign n15365 = controllable_hmaster0 & ~n15363;
  assign n15366 = ~n3920 & ~n6007;
  assign n15367 = ~i_hlock0 & ~n15366;
  assign n15368 = ~n6020 & ~n15367;
  assign n15369 = ~i_hbusreq0 & ~n15368;
  assign n15370 = ~n6016 & ~n15369;
  assign n15371 = ~i_hbusreq4 & ~n15370;
  assign n15372 = ~n6015 & ~n15371;
  assign n15373 = ~controllable_hgrant4 & ~n15372;
  assign n15374 = ~n3433 & ~n15373;
  assign n15375 = ~i_hbusreq2 & ~n15374;
  assign n15376 = ~n6014 & ~n15375;
  assign n15377 = controllable_hgrant2 & ~n15376;
  assign n15378 = ~n12185 & ~n15377;
  assign n15379 = ~controllable_hmaster0 & ~n15378;
  assign n15380 = ~n15365 & ~n15379;
  assign n15381 = ~controllable_hmaster1 & ~n15380;
  assign n15382 = ~n15364 & ~n15381;
  assign n15383 = ~i_hbusreq3 & ~n15382;
  assign n15384 = ~n15362 & ~n15383;
  assign n15385 = controllable_hmaster2 & ~n15384;
  assign n15386 = ~n5683 & ~n6762;
  assign n15387 = controllable_hmaster0 & ~n15386;
  assign n15388 = ~n9498 & ~n15387;
  assign n15389 = controllable_hmaster1 & ~n15388;
  assign n15390 = ~n5699 & ~n6762;
  assign n15391 = controllable_hmaster0 & ~n15390;
  assign n15392 = ~controllable_hmaster0 & ~n15386;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = ~controllable_hmaster1 & ~n15393;
  assign n15395 = ~n15389 & ~n15394;
  assign n15396 = i_hbusreq3 & ~n15395;
  assign n15397 = ~n12208 & ~n15377;
  assign n15398 = controllable_hmaster0 & ~n15397;
  assign n15399 = ~n6813 & ~n12202;
  assign n15400 = ~controllable_hmaster0 & ~n15399;
  assign n15401 = ~n15398 & ~n15400;
  assign n15402 = controllable_hmaster1 & ~n15401;
  assign n15403 = ~n12216 & ~n15377;
  assign n15404 = controllable_hmaster0 & ~n15403;
  assign n15405 = ~controllable_hmaster0 & ~n15397;
  assign n15406 = ~n15404 & ~n15405;
  assign n15407 = ~controllable_hmaster1 & ~n15406;
  assign n15408 = ~n15402 & ~n15407;
  assign n15409 = ~i_hbusreq3 & ~n15408;
  assign n15410 = ~n15396 & ~n15409;
  assign n15411 = ~controllable_hmaster2 & ~n15410;
  assign n15412 = ~n15385 & ~n15411;
  assign n15413 = ~controllable_hgrant3 & ~n15412;
  assign n15414 = ~n15042 & ~n15413;
  assign n15415 = controllable_nhgrant0 & ~n15414;
  assign n15416 = ~n15088 & ~n15415;
  assign n15417 = ~n3281 & ~n15416;
  assign n15418 = ~n4089 & ~n15417;
  assign n15419 = n3378 & ~n15418;
  assign n15420 = ~n9480 & ~n12549;
  assign n15421 = ~controllable_hmaster1 & ~n15420;
  assign n15422 = ~n9479 & ~n15421;
  assign n15423 = i_hbusreq3 & ~n15422;
  assign n15424 = ~n9072 & ~n14547;
  assign n15425 = ~i_hbusreq0 & ~n15424;
  assign n15426 = ~n9069 & ~n15425;
  assign n15427 = ~i_hbusreq4 & ~n15426;
  assign n15428 = ~n9068 & ~n15427;
  assign n15429 = ~controllable_hgrant4 & ~n15428;
  assign n15430 = ~n3916 & ~n15429;
  assign n15431 = ~i_hbusreq2 & ~n15430;
  assign n15432 = ~n9067 & ~n15431;
  assign n15433 = controllable_hgrant2 & ~n15432;
  assign n15434 = ~n5881 & ~n15433;
  assign n15435 = controllable_hmaster1 & ~n15434;
  assign n15436 = controllable_hmaster0 & ~n15434;
  assign n15437 = ~n12555 & ~n15436;
  assign n15438 = ~controllable_hmaster1 & ~n15437;
  assign n15439 = ~n15435 & ~n15438;
  assign n15440 = ~i_hbusreq3 & ~n15439;
  assign n15441 = ~n15423 & ~n15440;
  assign n15442 = controllable_hmaster2 & ~n15441;
  assign n15443 = ~n6785 & ~n9498;
  assign n15444 = controllable_hmaster1 & ~n15443;
  assign n15445 = ~n6795 & ~n15444;
  assign n15446 = i_hbusreq3 & ~n15445;
  assign n15447 = ~n6813 & ~n12282;
  assign n15448 = ~controllable_hmaster0 & ~n15447;
  assign n15449 = ~n6799 & ~n15448;
  assign n15450 = controllable_hmaster1 & ~n15449;
  assign n15451 = ~n6835 & ~n15450;
  assign n15452 = ~i_hbusreq3 & ~n15451;
  assign n15453 = ~n15446 & ~n15452;
  assign n15454 = ~controllable_hmaster2 & ~n15453;
  assign n15455 = ~n15442 & ~n15454;
  assign n15456 = ~controllable_hgrant3 & ~n15455;
  assign n15457 = ~n5861 & ~n15456;
  assign n15458 = controllable_nhgrant0 & ~n15457;
  assign n15459 = ~n6082 & ~n15458;
  assign n15460 = ~n3281 & ~n15459;
  assign n15461 = ~n4089 & ~n15460;
  assign n15462 = ~n3378 & ~n15461;
  assign n15463 = ~n15419 & ~n15462;
  assign n15464 = n3492 & ~n15463;
  assign n15465 = ~n15258 & ~n15464;
  assign n15466 = n3485 & ~n15465;
  assign n15467 = ~n15257 & ~n15466;
  assign n15468 = n3476 & ~n15467;
  assign n15469 = ~n15356 & ~n15468;
  assign n15470 = n3374 & ~n15469;
  assign n15471 = ~n15264 & ~n15470;
  assign n15472 = n3655 & ~n15471;
  assign n15473 = ~n6102 & ~n9388;
  assign n15474 = controllable_hmaster1 & ~n15473;
  assign n15475 = controllable_hmaster0 & ~n15473;
  assign n15476 = ~n3729 & ~n15475;
  assign n15477 = ~controllable_hmaster1 & ~n15476;
  assign n15478 = ~n15474 & ~n15477;
  assign n15479 = i_hbusreq3 & ~n15478;
  assign n15480 = ~n6127 & ~n15233;
  assign n15481 = controllable_hmaster1 & ~n15480;
  assign n15482 = controllable_hmaster0 & ~n15480;
  assign n15483 = ~n3767 & ~n15482;
  assign n15484 = ~controllable_hmaster1 & ~n15483;
  assign n15485 = ~n15481 & ~n15484;
  assign n15486 = ~i_hbusreq3 & ~n15485;
  assign n15487 = ~n15479 & ~n15486;
  assign n15488 = controllable_hmaster2 & ~n15487;
  assign n15489 = ~n6887 & ~n15488;
  assign n15490 = ~controllable_hgrant3 & ~n15489;
  assign n15491 = ~n5037 & ~n15490;
  assign n15492 = controllable_nhgrant0 & ~n15491;
  assign n15493 = ~n5245 & ~n15492;
  assign n15494 = ~n3281 & ~n15493;
  assign n15495 = ~n3783 & ~n15494;
  assign n15496 = ~n3378 & ~n15495;
  assign n15497 = ~n15225 & ~n15496;
  assign n15498 = n3492 & ~n15497;
  assign n15499 = ~n3631 & ~n15498;
  assign n15500 = n3485 & ~n15499;
  assign n15501 = ~n3630 & ~n15500;
  assign n15502 = ~n3476 & ~n15501;
  assign n15503 = ~n15258 & ~n15498;
  assign n15504 = n3485 & ~n15503;
  assign n15505 = ~n15257 & ~n15504;
  assign n15506 = n3476 & ~n15505;
  assign n15507 = ~n15502 & ~n15506;
  assign n15508 = ~n3374 & ~n15507;
  assign n15509 = ~n9590 & ~n15289;
  assign n15510 = controllable_hmaster1 & ~n15509;
  assign n15511 = ~n15296 & ~n15510;
  assign n15512 = i_hbusreq3 & ~n15511;
  assign n15513 = ~n9603 & ~n15300;
  assign n15514 = controllable_hmaster1 & ~n15513;
  assign n15515 = ~n15307 & ~n15514;
  assign n15516 = ~i_hbusreq3 & ~n15515;
  assign n15517 = ~n15512 & ~n15516;
  assign n15518 = ~controllable_hmaster2 & ~n15517;
  assign n15519 = ~n15287 & ~n15518;
  assign n15520 = ~controllable_hgrant3 & ~n15519;
  assign n15521 = ~n14973 & ~n15520;
  assign n15522 = controllable_nhgrant0 & ~n15521;
  assign n15523 = ~n15006 & ~n15522;
  assign n15524 = ~n3281 & ~n15523;
  assign n15525 = ~n3950 & ~n15524;
  assign n15526 = n3378 & ~n15525;
  assign n15527 = ~n6214 & ~n9388;
  assign n15528 = controllable_hmaster1 & ~n15527;
  assign n15529 = controllable_hmaster0 & ~n15527;
  assign n15530 = ~n12617 & ~n15529;
  assign n15531 = ~controllable_hmaster1 & ~n15530;
  assign n15532 = ~n15528 & ~n15531;
  assign n15533 = i_hbusreq3 & ~n15532;
  assign n15534 = ~n6237 & ~n15233;
  assign n15535 = controllable_hmaster1 & ~n15534;
  assign n15536 = controllable_hmaster0 & ~n15534;
  assign n15537 = ~n12623 & ~n15536;
  assign n15538 = ~controllable_hmaster1 & ~n15537;
  assign n15539 = ~n15535 & ~n15538;
  assign n15540 = ~i_hbusreq3 & ~n15539;
  assign n15541 = ~n15533 & ~n15540;
  assign n15542 = controllable_hmaster2 & ~n15541;
  assign n15543 = ~n6927 & ~n9590;
  assign n15544 = controllable_hmaster1 & ~n15543;
  assign n15545 = ~n6936 & ~n15544;
  assign n15546 = i_hbusreq3 & ~n15545;
  assign n15547 = ~n6940 & ~n9603;
  assign n15548 = controllable_hmaster1 & ~n15547;
  assign n15549 = ~n6951 & ~n15548;
  assign n15550 = ~i_hbusreq3 & ~n15549;
  assign n15551 = ~n15546 & ~n15550;
  assign n15552 = ~controllable_hmaster2 & ~n15551;
  assign n15553 = ~n15542 & ~n15552;
  assign n15554 = ~controllable_hgrant3 & ~n15553;
  assign n15555 = ~n5402 & ~n15554;
  assign n15556 = controllable_nhgrant0 & ~n15555;
  assign n15557 = ~n5534 & ~n15556;
  assign n15558 = ~n3281 & ~n15557;
  assign n15559 = ~n3950 & ~n15558;
  assign n15560 = ~n3378 & ~n15559;
  assign n15561 = ~n15526 & ~n15560;
  assign n15562 = n3492 & ~n15561;
  assign n15563 = ~n3631 & ~n15562;
  assign n15564 = n3485 & ~n15563;
  assign n15565 = ~n3630 & ~n15564;
  assign n15566 = ~n3476 & ~n15565;
  assign n15567 = ~n6786 & ~n12379;
  assign n15568 = ~controllable_hmaster0 & ~n15567;
  assign n15569 = ~n15387 & ~n15568;
  assign n15570 = controllable_hmaster1 & ~n15569;
  assign n15571 = ~n15394 & ~n15570;
  assign n15572 = i_hbusreq3 & ~n15571;
  assign n15573 = ~n6813 & ~n12390;
  assign n15574 = ~controllable_hmaster0 & ~n15573;
  assign n15575 = ~n15398 & ~n15574;
  assign n15576 = controllable_hmaster1 & ~n15575;
  assign n15577 = ~n15407 & ~n15576;
  assign n15578 = ~i_hbusreq3 & ~n15577;
  assign n15579 = ~n15572 & ~n15578;
  assign n15580 = ~controllable_hmaster2 & ~n15579;
  assign n15581 = ~n15385 & ~n15580;
  assign n15582 = ~controllable_hgrant3 & ~n15581;
  assign n15583 = ~n15042 & ~n15582;
  assign n15584 = controllable_nhgrant0 & ~n15583;
  assign n15585 = ~n15088 & ~n15584;
  assign n15586 = ~n3281 & ~n15585;
  assign n15587 = ~n4089 & ~n15586;
  assign n15588 = n3378 & ~n15587;
  assign n15589 = ~n6405 & ~n9477;
  assign n15590 = controllable_hmaster1 & ~n15589;
  assign n15591 = controllable_hmaster0 & ~n15589;
  assign n15592 = ~n12677 & ~n15591;
  assign n15593 = ~controllable_hmaster1 & ~n15592;
  assign n15594 = ~n15590 & ~n15593;
  assign n15595 = i_hbusreq3 & ~n15594;
  assign n15596 = ~n6437 & ~n15433;
  assign n15597 = controllable_hmaster1 & ~n15596;
  assign n15598 = controllable_hmaster0 & ~n15596;
  assign n15599 = ~n12683 & ~n15598;
  assign n15600 = ~controllable_hmaster1 & ~n15599;
  assign n15601 = ~n15597 & ~n15600;
  assign n15602 = ~i_hbusreq3 & ~n15601;
  assign n15603 = ~n15595 & ~n15602;
  assign n15604 = controllable_hmaster2 & ~n15603;
  assign n15605 = ~n7013 & ~n9650;
  assign n15606 = controllable_hmaster1 & ~n15605;
  assign n15607 = ~n7022 & ~n15606;
  assign n15608 = i_hbusreq3 & ~n15607;
  assign n15609 = ~n6813 & ~n12435;
  assign n15610 = ~controllable_hmaster0 & ~n15609;
  assign n15611 = ~n7026 & ~n15610;
  assign n15612 = controllable_hmaster1 & ~n15611;
  assign n15613 = ~n7036 & ~n15612;
  assign n15614 = ~i_hbusreq3 & ~n15613;
  assign n15615 = ~n15608 & ~n15614;
  assign n15616 = ~controllable_hmaster2 & ~n15615;
  assign n15617 = ~n15604 & ~n15616;
  assign n15618 = ~controllable_hgrant3 & ~n15617;
  assign n15619 = ~n5861 & ~n15618;
  assign n15620 = controllable_nhgrant0 & ~n15619;
  assign n15621 = ~n6082 & ~n15620;
  assign n15622 = ~n3281 & ~n15621;
  assign n15623 = ~n4089 & ~n15622;
  assign n15624 = ~n3378 & ~n15623;
  assign n15625 = ~n15588 & ~n15624;
  assign n15626 = n3492 & ~n15625;
  assign n15627 = ~n15258 & ~n15626;
  assign n15628 = n3485 & ~n15627;
  assign n15629 = ~n15257 & ~n15628;
  assign n15630 = n3476 & ~n15629;
  assign n15631 = ~n15566 & ~n15630;
  assign n15632 = n3374 & ~n15631;
  assign n15633 = ~n15508 & ~n15632;
  assign n15634 = ~n3655 & ~n15633;
  assign n15635 = ~n15472 & ~n15634;
  assign n15636 = ~n3652 & ~n15635;
  assign n15637 = ~n15224 & ~n15636;
  assign n15638 = ~n3368 & ~n15637;
  assign n15639 = ~n4553 & ~n5277;
  assign n15640 = controllable_hmaster1 & ~n15639;
  assign n15641 = ~n5281 & ~n15640;
  assign n15642 = ~i_hbusreq3 & ~n15641;
  assign n15643 = ~n5265 & ~n15642;
  assign n15644 = ~controllable_hmaster2 & ~n15643;
  assign n15645 = ~n12033 & ~n15644;
  assign n15646 = controllable_hgrant3 & ~n15645;
  assign n15647 = ~n3401 & ~n9805;
  assign n15648 = controllable_hmaster1 & ~n15647;
  assign n15649 = ~n5334 & ~n15648;
  assign n15650 = ~i_hbusreq3 & ~n15649;
  assign n15651 = ~n14977 & ~n15650;
  assign n15652 = ~controllable_hmaster2 & ~n15651;
  assign n15653 = ~n12741 & ~n15652;
  assign n15654 = ~controllable_hgrant3 & ~n15653;
  assign n15655 = ~n15646 & ~n15654;
  assign n15656 = controllable_nhgrant0 & ~n15655;
  assign n15657 = controllable_hmaster1 & ~n7129;
  assign n15658 = ~n5281 & ~n15657;
  assign n15659 = ~i_hbusreq3 & ~n15658;
  assign n15660 = ~n3951 & ~n15659;
  assign n15661 = ~controllable_hmaster2 & ~n15660;
  assign n15662 = ~n12033 & ~n15661;
  assign n15663 = controllable_hgrant3 & ~n15662;
  assign n15664 = controllable_hmaster1 & ~n7153;
  assign n15665 = ~n5350 & ~n15664;
  assign n15666 = i_hbusreq3 & ~n15665;
  assign n15667 = controllable_hmaster1 & ~n7157;
  assign n15668 = ~n5355 & ~n15667;
  assign n15669 = ~i_hbusreq3 & ~n15668;
  assign n15670 = ~n15666 & ~n15669;
  assign n15671 = ~controllable_hmaster2 & ~n15670;
  assign n15672 = ~n12033 & ~n15671;
  assign n15673 = ~controllable_hgrant3 & ~n15672;
  assign n15674 = ~n15663 & ~n15673;
  assign n15675 = ~controllable_nhgrant0 & ~n15674;
  assign n15676 = ~n15656 & ~n15675;
  assign n15677 = ~n3281 & ~n15676;
  assign n15678 = ~n3281 & ~n15677;
  assign n15679 = n3378 & ~n15678;
  assign n15680 = ~n4553 & ~n5377;
  assign n15681 = controllable_hmaster1 & ~n15680;
  assign n15682 = ~n5396 & ~n15681;
  assign n15683 = ~i_hbusreq3 & ~n15682;
  assign n15684 = ~n5265 & ~n15683;
  assign n15685 = ~controllable_hmaster2 & ~n15684;
  assign n15686 = ~n5370 & ~n15685;
  assign n15687 = controllable_hgrant3 & ~n15686;
  assign n15688 = ~n5197 & ~n9805;
  assign n15689 = controllable_hmaster1 & ~n15688;
  assign n15690 = ~n5480 & ~n15689;
  assign n15691 = ~i_hbusreq3 & ~n15690;
  assign n15692 = ~n15014 & ~n15691;
  assign n15693 = ~controllable_hmaster2 & ~n15692;
  assign n15694 = ~n12795 & ~n15693;
  assign n15695 = ~controllable_hgrant3 & ~n15694;
  assign n15696 = ~n15687 & ~n15695;
  assign n15697 = controllable_nhgrant0 & ~n15696;
  assign n15698 = controllable_hmaster1 & ~n7171;
  assign n15699 = ~n5396 & ~n15698;
  assign n15700 = ~i_hbusreq3 & ~n15699;
  assign n15701 = ~n3951 & ~n15700;
  assign n15702 = ~controllable_hmaster2 & ~n15701;
  assign n15703 = ~n5370 & ~n15702;
  assign n15704 = controllable_hgrant3 & ~n15703;
  assign n15705 = controllable_hmaster1 & ~n7195;
  assign n15706 = ~n5501 & ~n15705;
  assign n15707 = i_hbusreq3 & ~n15706;
  assign n15708 = controllable_hmaster1 & ~n7199;
  assign n15709 = ~n5526 & ~n15708;
  assign n15710 = ~i_hbusreq3 & ~n15709;
  assign n15711 = ~n15707 & ~n15710;
  assign n15712 = ~controllable_hmaster2 & ~n15711;
  assign n15713 = ~n5498 & ~n15712;
  assign n15714 = ~controllable_hgrant3 & ~n15713;
  assign n15715 = ~n15704 & ~n15714;
  assign n15716 = ~controllable_nhgrant0 & ~n15715;
  assign n15717 = ~n15697 & ~n15716;
  assign n15718 = ~n3281 & ~n15717;
  assign n15719 = ~n3281 & ~n15718;
  assign n15720 = ~n3378 & ~n15719;
  assign n15721 = ~n15679 & ~n15720;
  assign n15722 = n3492 & ~n15721;
  assign n15723 = n3492 & ~n15722;
  assign n15724 = n3485 & ~n15723;
  assign n15725 = n3485 & ~n15724;
  assign n15726 = ~n3476 & ~n15725;
  assign n15727 = ~n5605 & ~n7232;
  assign n15728 = controllable_hmaster1 & ~n15727;
  assign n15729 = ~n5609 & ~n15728;
  assign n15730 = ~i_hbusreq3 & ~n15729;
  assign n15731 = ~n5593 & ~n15730;
  assign n15732 = ~controllable_hmaster2 & ~n15731;
  assign n15733 = ~n12233 & ~n15732;
  assign n15734 = controllable_hgrant3 & ~n15733;
  assign n15735 = controllable_hgrant2 & ~n12841;
  assign n15736 = ~n12868 & ~n15735;
  assign n15737 = controllable_hmaster1 & ~n15736;
  assign n15738 = controllable_hmaster0 & ~n15736;
  assign n15739 = ~n12876 & ~n15735;
  assign n15740 = ~controllable_hmaster0 & ~n15739;
  assign n15741 = ~n15738 & ~n15740;
  assign n15742 = ~controllable_hmaster1 & ~n15741;
  assign n15743 = ~n15737 & ~n15742;
  assign n15744 = ~i_hbusreq3 & ~n15743;
  assign n15745 = ~n12864 & ~n15744;
  assign n15746 = controllable_hmaster2 & ~n15745;
  assign n15747 = ~n5686 & ~n12886;
  assign n15748 = ~controllable_hmaster0 & ~n15747;
  assign n15749 = ~n7326 & ~n15748;
  assign n15750 = controllable_hmaster1 & ~n15749;
  assign n15751 = ~n7342 & ~n15750;
  assign n15752 = i_hbusreq3 & ~n15751;
  assign n15753 = ~n12904 & ~n15735;
  assign n15754 = controllable_hmaster0 & ~n15753;
  assign n15755 = ~n10152 & ~n12898;
  assign n15756 = ~controllable_hmaster0 & ~n15755;
  assign n15757 = ~n15754 & ~n15756;
  assign n15758 = controllable_hmaster1 & ~n15757;
  assign n15759 = ~n12912 & ~n15735;
  assign n15760 = controllable_hmaster0 & ~n15759;
  assign n15761 = ~controllable_hmaster0 & ~n15753;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = ~controllable_hmaster1 & ~n15762;
  assign n15764 = ~n15758 & ~n15763;
  assign n15765 = ~i_hbusreq3 & ~n15764;
  assign n15766 = ~n15752 & ~n15765;
  assign n15767 = ~controllable_hmaster2 & ~n15766;
  assign n15768 = ~n15746 & ~n15767;
  assign n15769 = ~controllable_hgrant3 & ~n15768;
  assign n15770 = ~n15734 & ~n15769;
  assign n15771 = controllable_nhgrant0 & ~n15770;
  assign n15772 = controllable_hmaster1 & ~n7400;
  assign n15773 = ~n5796 & ~n15772;
  assign n15774 = i_hbusreq3 & ~n15773;
  assign n15775 = controllable_hmaster1 & ~n7423;
  assign n15776 = ~n5801 & ~n15775;
  assign n15777 = ~i_hbusreq3 & ~n15776;
  assign n15778 = ~n15774 & ~n15777;
  assign n15779 = ~controllable_hmaster2 & ~n15778;
  assign n15780 = ~n12233 & ~n15779;
  assign n15781 = ~controllable_hgrant3 & ~n15780;
  assign n15782 = ~n15663 & ~n15781;
  assign n15783 = ~controllable_nhgrant0 & ~n15782;
  assign n15784 = ~n15771 & ~n15783;
  assign n15785 = ~n3281 & ~n15784;
  assign n15786 = ~n3281 & ~n15785;
  assign n15787 = n3378 & ~n15786;
  assign n15788 = ~n5835 & ~n7449;
  assign n15789 = controllable_hmaster1 & ~n15788;
  assign n15790 = ~n5855 & ~n15789;
  assign n15791 = ~i_hbusreq3 & ~n15790;
  assign n15792 = ~n5593 & ~n15791;
  assign n15793 = ~controllable_hmaster2 & ~n15792;
  assign n15794 = ~n5828 & ~n15793;
  assign n15795 = controllable_hgrant3 & ~n15794;
  assign n15796 = controllable_hgrant2 & ~n12950;
  assign n15797 = ~n12986 & ~n15796;
  assign n15798 = controllable_hmaster1 & ~n15797;
  assign n15799 = controllable_hmaster0 & ~n15797;
  assign n15800 = ~n12994 & ~n15796;
  assign n15801 = ~controllable_hmaster0 & ~n15800;
  assign n15802 = ~n15799 & ~n15801;
  assign n15803 = ~controllable_hmaster1 & ~n15802;
  assign n15804 = ~n15798 & ~n15803;
  assign n15805 = ~i_hbusreq3 & ~n15804;
  assign n15806 = ~n12982 & ~n15805;
  assign n15807 = controllable_hmaster2 & ~n15806;
  assign n15808 = ~n5686 & ~n13004;
  assign n15809 = ~controllable_hmaster0 & ~n15808;
  assign n15810 = ~n7539 & ~n15809;
  assign n15811 = controllable_hmaster1 & ~n15810;
  assign n15812 = ~n7554 & ~n15811;
  assign n15813 = i_hbusreq3 & ~n15812;
  assign n15814 = ~n13022 & ~n15796;
  assign n15815 = controllable_hmaster0 & ~n15814;
  assign n15816 = ~n10152 & ~n13016;
  assign n15817 = ~controllable_hmaster0 & ~n15816;
  assign n15818 = ~n15815 & ~n15817;
  assign n15819 = controllable_hmaster1 & ~n15818;
  assign n15820 = ~n13030 & ~n15796;
  assign n15821 = controllable_hmaster0 & ~n15820;
  assign n15822 = controllable_hgrant2 & ~n12963;
  assign n15823 = ~n13036 & ~n15822;
  assign n15824 = ~controllable_hmaster0 & ~n15823;
  assign n15825 = ~n15821 & ~n15824;
  assign n15826 = ~controllable_hmaster1 & ~n15825;
  assign n15827 = ~n15819 & ~n15826;
  assign n15828 = ~i_hbusreq3 & ~n15827;
  assign n15829 = ~n15813 & ~n15828;
  assign n15830 = ~controllable_hmaster2 & ~n15829;
  assign n15831 = ~n15807 & ~n15830;
  assign n15832 = ~controllable_hgrant3 & ~n15831;
  assign n15833 = ~n15795 & ~n15832;
  assign n15834 = controllable_nhgrant0 & ~n15833;
  assign n15835 = controllable_hmaster1 & ~n7637;
  assign n15836 = ~n6046 & ~n15835;
  assign n15837 = i_hbusreq3 & ~n15836;
  assign n15838 = controllable_hmaster1 & ~n7659;
  assign n15839 = ~n6074 & ~n15838;
  assign n15840 = ~i_hbusreq3 & ~n15839;
  assign n15841 = ~n15837 & ~n15840;
  assign n15842 = ~controllable_hmaster2 & ~n15841;
  assign n15843 = ~n6035 & ~n15842;
  assign n15844 = ~controllable_hgrant3 & ~n15843;
  assign n15845 = ~n15704 & ~n15844;
  assign n15846 = ~controllable_nhgrant0 & ~n15845;
  assign n15847 = ~n15834 & ~n15846;
  assign n15848 = ~n3281 & ~n15847;
  assign n15849 = ~n3281 & ~n15848;
  assign n15850 = ~n3378 & ~n15849;
  assign n15851 = ~n15787 & ~n15850;
  assign n15852 = n3492 & ~n15851;
  assign n15853 = n3492 & ~n15852;
  assign n15854 = n3485 & ~n15853;
  assign n15855 = n3485 & ~n15854;
  assign n15856 = n3476 & ~n15855;
  assign n15857 = ~n15726 & ~n15856;
  assign n15858 = n3374 & ~n15857;
  assign n15859 = ~n7128 & ~n15858;
  assign n15860 = n3655 & ~n15859;
  assign n15861 = ~n3382 & ~n10328;
  assign n15862 = controllable_hmaster1 & ~n15861;
  assign n15863 = ~n5305 & ~n15862;
  assign n15864 = i_hbusreq3 & ~n15863;
  assign n15865 = ~n3401 & ~n10350;
  assign n15866 = controllable_hmaster1 & ~n15865;
  assign n15867 = ~n5334 & ~n15866;
  assign n15868 = ~i_hbusreq3 & ~n15867;
  assign n15869 = ~n15864 & ~n15868;
  assign n15870 = ~controllable_hmaster2 & ~n15869;
  assign n15871 = ~n12741 & ~n15870;
  assign n15872 = ~controllable_hgrant3 & ~n15871;
  assign n15873 = ~n15646 & ~n15872;
  assign n15874 = controllable_nhgrant0 & ~n15873;
  assign n15875 = ~n15675 & ~n15874;
  assign n15876 = ~n3281 & ~n15875;
  assign n15877 = ~n3281 & ~n15876;
  assign n15878 = n3378 & ~n15877;
  assign n15879 = ~n6254 & ~n10328;
  assign n15880 = controllable_hmaster1 & ~n15879;
  assign n15881 = ~n6271 & ~n15880;
  assign n15882 = i_hbusreq3 & ~n15881;
  assign n15883 = ~n6293 & ~n10350;
  assign n15884 = controllable_hmaster1 & ~n15883;
  assign n15885 = ~n6339 & ~n15884;
  assign n15886 = ~i_hbusreq3 & ~n15885;
  assign n15887 = ~n15882 & ~n15886;
  assign n15888 = ~controllable_hmaster2 & ~n15887;
  assign n15889 = ~n13106 & ~n15888;
  assign n15890 = ~controllable_hgrant3 & ~n15889;
  assign n15891 = ~n15687 & ~n15890;
  assign n15892 = controllable_nhgrant0 & ~n15891;
  assign n15893 = ~n15716 & ~n15892;
  assign n15894 = ~n3281 & ~n15893;
  assign n15895 = ~n3281 & ~n15894;
  assign n15896 = ~n3378 & ~n15895;
  assign n15897 = ~n15878 & ~n15896;
  assign n15898 = n3492 & ~n15897;
  assign n15899 = n3492 & ~n15898;
  assign n15900 = n3485 & ~n15899;
  assign n15901 = n3485 & ~n15900;
  assign n15902 = ~n3476 & ~n15901;
  assign n15903 = ~n5686 & ~n13132;
  assign n15904 = ~controllable_hmaster0 & ~n15903;
  assign n15905 = ~n7326 & ~n15904;
  assign n15906 = controllable_hmaster1 & ~n15905;
  assign n15907 = ~n7342 & ~n15906;
  assign n15908 = i_hbusreq3 & ~n15907;
  assign n15909 = ~n10152 & ~n13143;
  assign n15910 = ~controllable_hmaster0 & ~n15909;
  assign n15911 = ~n15754 & ~n15910;
  assign n15912 = controllable_hmaster1 & ~n15911;
  assign n15913 = ~n15763 & ~n15912;
  assign n15914 = ~i_hbusreq3 & ~n15913;
  assign n15915 = ~n15908 & ~n15914;
  assign n15916 = ~controllable_hmaster2 & ~n15915;
  assign n15917 = ~n15746 & ~n15916;
  assign n15918 = ~controllable_hgrant3 & ~n15917;
  assign n15919 = ~n15734 & ~n15918;
  assign n15920 = controllable_nhgrant0 & ~n15919;
  assign n15921 = ~n15783 & ~n15920;
  assign n15922 = ~n3281 & ~n15921;
  assign n15923 = ~n3281 & ~n15922;
  assign n15924 = n3378 & ~n15923;
  assign n15925 = ~n13171 & ~n15796;
  assign n15926 = controllable_hmaster1 & ~n15925;
  assign n15927 = controllable_hmaster0 & ~n15925;
  assign n15928 = ~n13179 & ~n15796;
  assign n15929 = ~controllable_hmaster0 & ~n15928;
  assign n15930 = ~n15927 & ~n15929;
  assign n15931 = ~controllable_hmaster1 & ~n15930;
  assign n15932 = ~n15926 & ~n15931;
  assign n15933 = ~i_hbusreq3 & ~n15932;
  assign n15934 = ~n13167 & ~n15933;
  assign n15935 = controllable_hmaster2 & ~n15934;
  assign n15936 = ~n5686 & ~n13189;
  assign n15937 = ~controllable_hmaster0 & ~n15936;
  assign n15938 = ~n7863 & ~n15937;
  assign n15939 = controllable_hmaster1 & ~n15938;
  assign n15940 = ~n7877 & ~n15939;
  assign n15941 = i_hbusreq3 & ~n15940;
  assign n15942 = ~n13206 & ~n15796;
  assign n15943 = controllable_hmaster0 & ~n15942;
  assign n15944 = ~n10152 & ~n13200;
  assign n15945 = ~controllable_hmaster0 & ~n15944;
  assign n15946 = ~n15943 & ~n15945;
  assign n15947 = controllable_hmaster1 & ~n15946;
  assign n15948 = ~n13214 & ~n15796;
  assign n15949 = controllable_hmaster0 & ~n15948;
  assign n15950 = ~n13220 & ~n15822;
  assign n15951 = ~controllable_hmaster0 & ~n15950;
  assign n15952 = ~n15949 & ~n15951;
  assign n15953 = ~controllable_hmaster1 & ~n15952;
  assign n15954 = ~n15947 & ~n15953;
  assign n15955 = ~i_hbusreq3 & ~n15954;
  assign n15956 = ~n15941 & ~n15955;
  assign n15957 = ~controllable_hmaster2 & ~n15956;
  assign n15958 = ~n15935 & ~n15957;
  assign n15959 = ~controllable_hgrant3 & ~n15958;
  assign n15960 = ~n15795 & ~n15959;
  assign n15961 = controllable_nhgrant0 & ~n15960;
  assign n15962 = ~n15846 & ~n15961;
  assign n15963 = ~n3281 & ~n15962;
  assign n15964 = ~n3281 & ~n15963;
  assign n15965 = ~n3378 & ~n15964;
  assign n15966 = ~n15924 & ~n15965;
  assign n15967 = n3492 & ~n15966;
  assign n15968 = n3492 & ~n15967;
  assign n15969 = n3485 & ~n15968;
  assign n15970 = n3485 & ~n15969;
  assign n15971 = n3476 & ~n15970;
  assign n15972 = ~n15902 & ~n15971;
  assign n15973 = n3374 & ~n15972;
  assign n15974 = ~n7706 & ~n15973;
  assign n15975 = ~n3655 & ~n15974;
  assign n15976 = ~n15860 & ~n15975;
  assign n15977 = n3652 & ~n15976;
  assign n15978 = ~n4787 & ~n5258;
  assign n15979 = controllable_hmaster1 & ~n15978;
  assign n15980 = controllable_hmaster0 & ~n15978;
  assign n15981 = controllable_hmaster0 & ~n15980;
  assign n15982 = ~controllable_hmaster1 & ~n15981;
  assign n15983 = ~n15979 & ~n15982;
  assign n15984 = i_hbusreq3 & ~n15983;
  assign n15985 = ~n3390 & ~n4604;
  assign n15986 = ~i_hready & ~n15985;
  assign n15987 = ~i_hready & ~n15986;
  assign n15988 = ~i_hbusreq0 & ~n15987;
  assign n15989 = ~n4619 & ~n15988;
  assign n15990 = ~i_hbusreq4 & ~n15989;
  assign n15991 = ~n4618 & ~n15990;
  assign n15992 = ~controllable_hgrant4 & ~n15991;
  assign n15993 = ~n3433 & ~n15992;
  assign n15994 = ~i_hbusreq2 & ~n15993;
  assign n15995 = ~n4616 & ~n15994;
  assign n15996 = controllable_hgrant2 & ~n15995;
  assign n15997 = ~n5275 & ~n15996;
  assign n15998 = controllable_hmaster1 & ~n15997;
  assign n15999 = controllable_hmaster0 & ~n15997;
  assign n16000 = controllable_hmaster0 & ~n15999;
  assign n16001 = ~controllable_hmaster1 & ~n16000;
  assign n16002 = ~n15998 & ~n16001;
  assign n16003 = ~i_hbusreq3 & ~n16002;
  assign n16004 = ~n15984 & ~n16003;
  assign n16005 = controllable_hmaster2 & ~n16004;
  assign n16006 = controllable_hmaster2 & ~n16005;
  assign n16007 = ~controllable_hgrant3 & ~n16006;
  assign n16008 = ~n3409 & ~n16007;
  assign n16009 = controllable_nhgrant0 & ~n16008;
  assign n16010 = ~n3466 & ~n16009;
  assign n16011 = ~n3281 & ~n16010;
  assign n16012 = ~n3281 & ~n16011;
  assign n16013 = n3378 & ~n16012;
  assign n16014 = ~n4787 & ~n5043;
  assign n16015 = controllable_hmaster1 & ~n16014;
  assign n16016 = controllable_hmaster0 & ~n16014;
  assign n16017 = controllable_hmaster0 & ~n16016;
  assign n16018 = ~controllable_hmaster1 & ~n16017;
  assign n16019 = ~n16015 & ~n16018;
  assign n16020 = i_hbusreq3 & ~n16019;
  assign n16021 = i_hlock0 & ~n15987;
  assign n16022 = ~n4624 & ~n16021;
  assign n16023 = ~i_hbusreq0 & ~n16022;
  assign n16024 = ~n4619 & ~n16023;
  assign n16025 = ~i_hbusreq4 & ~n16024;
  assign n16026 = ~n4618 & ~n16025;
  assign n16027 = ~controllable_hgrant4 & ~n16026;
  assign n16028 = ~n3916 & ~n16027;
  assign n16029 = ~i_hbusreq2 & ~n16028;
  assign n16030 = ~n4616 & ~n16029;
  assign n16031 = controllable_hgrant2 & ~n16030;
  assign n16032 = ~n5068 & ~n16031;
  assign n16033 = controllable_hmaster1 & ~n16032;
  assign n16034 = controllable_hmaster0 & ~n16032;
  assign n16035 = controllable_hmaster0 & ~n16034;
  assign n16036 = ~controllable_hmaster1 & ~n16035;
  assign n16037 = ~n16033 & ~n16036;
  assign n16038 = ~i_hbusreq3 & ~n16037;
  assign n16039 = ~n16020 & ~n16038;
  assign n16040 = controllable_hmaster2 & ~n16039;
  assign n16041 = controllable_hmaster2 & ~n16040;
  assign n16042 = ~controllable_hgrant3 & ~n16041;
  assign n16043 = ~n7090 & ~n16042;
  assign n16044 = controllable_nhgrant0 & ~n16043;
  assign n16045 = ~n7118 & ~n16044;
  assign n16046 = ~n3281 & ~n16045;
  assign n16047 = ~n3281 & ~n16046;
  assign n16048 = ~n3378 & ~n16047;
  assign n16049 = ~n16013 & ~n16048;
  assign n16050 = n3492 & ~n16049;
  assign n16051 = n3492 & ~n16050;
  assign n16052 = n3485 & ~n16051;
  assign n16053 = n3485 & ~n16052;
  assign n16054 = ~n3374 & ~n16053;
  assign n16055 = ~n4787 & ~n12044;
  assign n16056 = ~controllable_hmaster0 & ~n16055;
  assign n16057 = ~n15980 & ~n16056;
  assign n16058 = ~controllable_hmaster1 & ~n16057;
  assign n16059 = ~n15979 & ~n16058;
  assign n16060 = i_hbusreq3 & ~n16059;
  assign n16061 = ~n12057 & ~n15996;
  assign n16062 = ~controllable_hmaster0 & ~n16061;
  assign n16063 = ~n15999 & ~n16062;
  assign n16064 = ~controllable_hmaster1 & ~n16063;
  assign n16065 = ~n15998 & ~n16064;
  assign n16066 = ~i_hbusreq3 & ~n16065;
  assign n16067 = ~n16060 & ~n16066;
  assign n16068 = controllable_hmaster2 & ~n16067;
  assign n16069 = ~n4787 & ~n5289;
  assign n16070 = controllable_hmaster0 & ~n16069;
  assign n16071 = ~n10770 & ~n16070;
  assign n16072 = controllable_hmaster1 & ~n16071;
  assign n16073 = ~n4787 & ~n5301;
  assign n16074 = controllable_hmaster0 & ~n16073;
  assign n16075 = ~controllable_hmaster0 & ~n16069;
  assign n16076 = ~n16074 & ~n16075;
  assign n16077 = ~controllable_hmaster1 & ~n16076;
  assign n16078 = ~n16072 & ~n16077;
  assign n16079 = i_hbusreq3 & ~n16078;
  assign n16080 = ~n5309 & ~n15996;
  assign n16081 = controllable_hmaster0 & ~n16080;
  assign n16082 = ~n10784 & ~n16081;
  assign n16083 = controllable_hmaster1 & ~n16082;
  assign n16084 = ~n5330 & ~n15996;
  assign n16085 = controllable_hmaster0 & ~n16084;
  assign n16086 = ~controllable_hmaster0 & ~n16080;
  assign n16087 = ~n16085 & ~n16086;
  assign n16088 = ~controllable_hmaster1 & ~n16087;
  assign n16089 = ~n16083 & ~n16088;
  assign n16090 = ~i_hbusreq3 & ~n16089;
  assign n16091 = ~n16079 & ~n16090;
  assign n16092 = ~controllable_hmaster2 & ~n16091;
  assign n16093 = ~n16068 & ~n16092;
  assign n16094 = ~controllable_hgrant3 & ~n16093;
  assign n16095 = ~n15646 & ~n16094;
  assign n16096 = controllable_nhgrant0 & ~n16095;
  assign n16097 = ~n15675 & ~n16096;
  assign n16098 = ~n3281 & ~n16097;
  assign n16099 = ~n3281 & ~n16098;
  assign n16100 = n3378 & ~n16099;
  assign n16101 = ~n4787 & ~n12107;
  assign n16102 = ~controllable_hmaster0 & ~n16101;
  assign n16103 = ~n16016 & ~n16102;
  assign n16104 = ~controllable_hmaster1 & ~n16103;
  assign n16105 = ~n16015 & ~n16104;
  assign n16106 = i_hbusreq3 & ~n16105;
  assign n16107 = ~n12118 & ~n16031;
  assign n16108 = ~controllable_hmaster0 & ~n16107;
  assign n16109 = ~n16034 & ~n16108;
  assign n16110 = ~controllable_hmaster1 & ~n16109;
  assign n16111 = ~n16033 & ~n16110;
  assign n16112 = ~i_hbusreq3 & ~n16111;
  assign n16113 = ~n16106 & ~n16112;
  assign n16114 = controllable_hmaster2 & ~n16113;
  assign n16115 = ~n3908 & ~n4787;
  assign n16116 = controllable_hmaster0 & ~n16115;
  assign n16117 = ~n10770 & ~n16116;
  assign n16118 = controllable_hmaster1 & ~n16117;
  assign n16119 = ~n4787 & ~n5431;
  assign n16120 = controllable_hmaster0 & ~n16119;
  assign n16121 = ~controllable_hmaster0 & ~n16115;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = ~controllable_hmaster1 & ~n16122;
  assign n16124 = ~n16118 & ~n16123;
  assign n16125 = i_hbusreq3 & ~n16124;
  assign n16126 = ~n3933 & ~n16031;
  assign n16127 = controllable_hmaster0 & ~n16126;
  assign n16128 = ~n10784 & ~n16127;
  assign n16129 = controllable_hmaster1 & ~n16128;
  assign n16130 = ~n5458 & ~n16031;
  assign n16131 = controllable_hmaster0 & ~n16130;
  assign n16132 = ~n4604 & ~n5382;
  assign n16133 = ~i_hready & ~n16132;
  assign n16134 = ~i_hready & ~n16133;
  assign n16135 = i_hlock0 & ~n16134;
  assign n16136 = ~n4624 & ~n16135;
  assign n16137 = ~i_hbusreq0 & ~n16136;
  assign n16138 = ~n4619 & ~n16137;
  assign n16139 = ~i_hbusreq4 & ~n16138;
  assign n16140 = ~n4618 & ~n16139;
  assign n16141 = ~controllable_hgrant4 & ~n16140;
  assign n16142 = ~n5462 & ~n16141;
  assign n16143 = ~i_hbusreq2 & ~n16142;
  assign n16144 = ~n4616 & ~n16143;
  assign n16145 = controllable_hgrant2 & ~n16144;
  assign n16146 = ~n5476 & ~n16145;
  assign n16147 = ~controllable_hmaster0 & ~n16146;
  assign n16148 = ~n16131 & ~n16147;
  assign n16149 = ~controllable_hmaster1 & ~n16148;
  assign n16150 = ~n16129 & ~n16149;
  assign n16151 = ~i_hbusreq3 & ~n16150;
  assign n16152 = ~n16125 & ~n16151;
  assign n16153 = ~controllable_hmaster2 & ~n16152;
  assign n16154 = ~n16114 & ~n16153;
  assign n16155 = ~controllable_hgrant3 & ~n16154;
  assign n16156 = ~n15687 & ~n16155;
  assign n16157 = controllable_nhgrant0 & ~n16156;
  assign n16158 = ~n15716 & ~n16157;
  assign n16159 = ~n3281 & ~n16158;
  assign n16160 = ~n3281 & ~n16159;
  assign n16161 = ~n3378 & ~n16160;
  assign n16162 = ~n16100 & ~n16161;
  assign n16163 = n3492 & ~n16162;
  assign n16164 = n3492 & ~n16163;
  assign n16165 = n3485 & ~n16164;
  assign n16166 = n3485 & ~n16165;
  assign n16167 = ~n3476 & ~n16166;
  assign n16168 = ~n7247 & ~n10827;
  assign n16169 = controllable_hmaster1 & ~n16168;
  assign n16170 = controllable_hmaster0 & ~n16168;
  assign n16171 = ~n10827 & ~n12858;
  assign n16172 = ~controllable_hmaster0 & ~n16171;
  assign n16173 = ~n16170 & ~n16172;
  assign n16174 = ~controllable_hmaster1 & ~n16173;
  assign n16175 = ~n16169 & ~n16174;
  assign n16176 = i_hbusreq3 & ~n16175;
  assign n16177 = ~n10842 & ~n15986;
  assign n16178 = ~i_hbusreq0 & ~n16177;
  assign n16179 = ~n10876 & ~n16178;
  assign n16180 = ~i_hbusreq4 & ~n16179;
  assign n16181 = ~n10875 & ~n16180;
  assign n16182 = ~controllable_hgrant4 & ~n16181;
  assign n16183 = ~n3433 & ~n16182;
  assign n16184 = i_hlock2 & ~n16183;
  assign n16185 = ~n9958 & ~n15986;
  assign n16186 = ~i_hbusreq0 & ~n16185;
  assign n16187 = ~n10890 & ~n16186;
  assign n16188 = ~i_hbusreq4 & ~n16187;
  assign n16189 = ~n10889 & ~n16188;
  assign n16190 = ~controllable_hgrant4 & ~n16189;
  assign n16191 = ~n3433 & ~n16190;
  assign n16192 = ~i_hlock2 & ~n16191;
  assign n16193 = ~n16184 & ~n16192;
  assign n16194 = ~i_hbusreq2 & ~n16193;
  assign n16195 = ~n10874 & ~n16194;
  assign n16196 = controllable_hgrant2 & ~n16195;
  assign n16197 = ~n12868 & ~n16196;
  assign n16198 = controllable_hmaster1 & ~n16197;
  assign n16199 = controllable_hmaster0 & ~n16197;
  assign n16200 = ~n12876 & ~n16196;
  assign n16201 = ~controllable_hmaster0 & ~n16200;
  assign n16202 = ~n16199 & ~n16201;
  assign n16203 = ~controllable_hmaster1 & ~n16202;
  assign n16204 = ~n16198 & ~n16203;
  assign n16205 = ~i_hbusreq3 & ~n16204;
  assign n16206 = ~n16176 & ~n16205;
  assign n16207 = controllable_hmaster2 & ~n16206;
  assign n16208 = ~n7324 & ~n10827;
  assign n16209 = controllable_hmaster0 & ~n16208;
  assign n16210 = ~n11066 & ~n12886;
  assign n16211 = ~controllable_hmaster0 & ~n16210;
  assign n16212 = ~n16209 & ~n16211;
  assign n16213 = controllable_hmaster1 & ~n16212;
  assign n16214 = ~n7337 & ~n10827;
  assign n16215 = controllable_hmaster0 & ~n16214;
  assign n16216 = ~controllable_hmaster0 & ~n16208;
  assign n16217 = ~n16215 & ~n16216;
  assign n16218 = ~controllable_hmaster1 & ~n16217;
  assign n16219 = ~n16213 & ~n16218;
  assign n16220 = i_hbusreq3 & ~n16219;
  assign n16221 = ~n12904 & ~n16196;
  assign n16222 = controllable_hmaster0 & ~n16221;
  assign n16223 = ~n11110 & ~n12898;
  assign n16224 = ~controllable_hmaster0 & ~n16223;
  assign n16225 = ~n16222 & ~n16224;
  assign n16226 = controllable_hmaster1 & ~n16225;
  assign n16227 = ~n12912 & ~n16196;
  assign n16228 = controllable_hmaster0 & ~n16227;
  assign n16229 = ~controllable_hmaster0 & ~n16221;
  assign n16230 = ~n16228 & ~n16229;
  assign n16231 = ~controllable_hmaster1 & ~n16230;
  assign n16232 = ~n16226 & ~n16231;
  assign n16233 = ~i_hbusreq3 & ~n16232;
  assign n16234 = ~n16220 & ~n16233;
  assign n16235 = ~controllable_hmaster2 & ~n16234;
  assign n16236 = ~n16207 & ~n16235;
  assign n16237 = ~controllable_hgrant3 & ~n16236;
  assign n16238 = ~n15734 & ~n16237;
  assign n16239 = controllable_nhgrant0 & ~n16238;
  assign n16240 = ~n15783 & ~n16239;
  assign n16241 = ~n3281 & ~n16240;
  assign n16242 = ~n3281 & ~n16241;
  assign n16243 = n3378 & ~n16242;
  assign n16244 = ~n7463 & ~n10827;
  assign n16245 = controllable_hmaster1 & ~n16244;
  assign n16246 = controllable_hmaster0 & ~n16244;
  assign n16247 = ~n10827 & ~n12976;
  assign n16248 = ~controllable_hmaster0 & ~n16247;
  assign n16249 = ~n16246 & ~n16248;
  assign n16250 = ~controllable_hmaster1 & ~n16249;
  assign n16251 = ~n16245 & ~n16250;
  assign n16252 = i_hbusreq3 & ~n16251;
  assign n16253 = i_hlock0 & ~n16177;
  assign n16254 = ~n10880 & ~n16253;
  assign n16255 = ~i_hbusreq0 & ~n16254;
  assign n16256 = ~n10876 & ~n16255;
  assign n16257 = ~i_hbusreq4 & ~n16256;
  assign n16258 = ~n10875 & ~n16257;
  assign n16259 = ~controllable_hgrant4 & ~n16258;
  assign n16260 = ~n3916 & ~n16259;
  assign n16261 = i_hlock2 & ~n16260;
  assign n16262 = i_hlock0 & ~n16185;
  assign n16263 = ~n9971 & ~n16262;
  assign n16264 = ~i_hbusreq0 & ~n16263;
  assign n16265 = ~n10890 & ~n16264;
  assign n16266 = ~i_hbusreq4 & ~n16265;
  assign n16267 = ~n10889 & ~n16266;
  assign n16268 = ~controllable_hgrant4 & ~n16267;
  assign n16269 = ~n3916 & ~n16268;
  assign n16270 = ~i_hlock2 & ~n16269;
  assign n16271 = ~n16261 & ~n16270;
  assign n16272 = ~i_hbusreq2 & ~n16271;
  assign n16273 = ~n10874 & ~n16272;
  assign n16274 = controllable_hgrant2 & ~n16273;
  assign n16275 = ~n12986 & ~n16274;
  assign n16276 = controllable_hmaster1 & ~n16275;
  assign n16277 = controllable_hmaster0 & ~n16275;
  assign n16278 = ~n12994 & ~n16274;
  assign n16279 = ~controllable_hmaster0 & ~n16278;
  assign n16280 = ~n16277 & ~n16279;
  assign n16281 = ~controllable_hmaster1 & ~n16280;
  assign n16282 = ~n16276 & ~n16281;
  assign n16283 = ~i_hbusreq3 & ~n16282;
  assign n16284 = ~n16252 & ~n16283;
  assign n16285 = controllable_hmaster2 & ~n16284;
  assign n16286 = ~n7537 & ~n10827;
  assign n16287 = controllable_hmaster0 & ~n16286;
  assign n16288 = ~n11066 & ~n13004;
  assign n16289 = ~controllable_hmaster0 & ~n16288;
  assign n16290 = ~n16287 & ~n16289;
  assign n16291 = controllable_hmaster1 & ~n16290;
  assign n16292 = ~n7549 & ~n10827;
  assign n16293 = controllable_hmaster0 & ~n16292;
  assign n16294 = ~controllable_hmaster0 & ~n16286;
  assign n16295 = ~n16293 & ~n16294;
  assign n16296 = ~controllable_hmaster1 & ~n16295;
  assign n16297 = ~n16291 & ~n16296;
  assign n16298 = i_hbusreq3 & ~n16297;
  assign n16299 = ~n13022 & ~n16274;
  assign n16300 = controllable_hmaster0 & ~n16299;
  assign n16301 = ~n11110 & ~n13016;
  assign n16302 = ~controllable_hmaster0 & ~n16301;
  assign n16303 = ~n16300 & ~n16302;
  assign n16304 = controllable_hmaster1 & ~n16303;
  assign n16305 = ~n13030 & ~n16274;
  assign n16306 = controllable_hmaster0 & ~n16305;
  assign n16307 = ~n10842 & ~n16133;
  assign n16308 = i_hlock0 & ~n16307;
  assign n16309 = ~n10880 & ~n16308;
  assign n16310 = ~i_hbusreq0 & ~n16309;
  assign n16311 = ~n10876 & ~n16310;
  assign n16312 = ~i_hbusreq4 & ~n16311;
  assign n16313 = ~n10875 & ~n16312;
  assign n16314 = ~controllable_hgrant4 & ~n16313;
  assign n16315 = ~n5462 & ~n16314;
  assign n16316 = i_hlock2 & ~n16315;
  assign n16317 = ~n9958 & ~n16133;
  assign n16318 = i_hlock0 & ~n16317;
  assign n16319 = ~n9971 & ~n16318;
  assign n16320 = ~i_hbusreq0 & ~n16319;
  assign n16321 = ~n10890 & ~n16320;
  assign n16322 = ~i_hbusreq4 & ~n16321;
  assign n16323 = ~n10889 & ~n16322;
  assign n16324 = ~controllable_hgrant4 & ~n16323;
  assign n16325 = ~n5462 & ~n16324;
  assign n16326 = ~i_hlock2 & ~n16325;
  assign n16327 = ~n16316 & ~n16326;
  assign n16328 = ~i_hbusreq2 & ~n16327;
  assign n16329 = ~n10874 & ~n16328;
  assign n16330 = controllable_hgrant2 & ~n16329;
  assign n16331 = ~n13036 & ~n16330;
  assign n16332 = ~controllable_hmaster0 & ~n16331;
  assign n16333 = ~n16306 & ~n16332;
  assign n16334 = ~controllable_hmaster1 & ~n16333;
  assign n16335 = ~n16304 & ~n16334;
  assign n16336 = ~i_hbusreq3 & ~n16335;
  assign n16337 = ~n16298 & ~n16336;
  assign n16338 = ~controllable_hmaster2 & ~n16337;
  assign n16339 = ~n16285 & ~n16338;
  assign n16340 = ~controllable_hgrant3 & ~n16339;
  assign n16341 = ~n15795 & ~n16340;
  assign n16342 = controllable_nhgrant0 & ~n16341;
  assign n16343 = ~n15846 & ~n16342;
  assign n16344 = ~n3281 & ~n16343;
  assign n16345 = ~n3281 & ~n16344;
  assign n16346 = ~n3378 & ~n16345;
  assign n16347 = ~n16243 & ~n16346;
  assign n16348 = n3492 & ~n16347;
  assign n16349 = ~n14836 & ~n16348;
  assign n16350 = n3485 & ~n16349;
  assign n16351 = ~n14835 & ~n16350;
  assign n16352 = n3476 & ~n16351;
  assign n16353 = ~n16167 & ~n16352;
  assign n16354 = n3374 & ~n16353;
  assign n16355 = ~n16054 & ~n16354;
  assign n16356 = n3655 & ~n16355;
  assign n16357 = ~n4787 & ~n6102;
  assign n16358 = controllable_hmaster1 & ~n16357;
  assign n16359 = controllable_hmaster0 & ~n16357;
  assign n16360 = controllable_hmaster0 & ~n16359;
  assign n16361 = ~controllable_hmaster1 & ~n16360;
  assign n16362 = ~n16358 & ~n16361;
  assign n16363 = i_hbusreq3 & ~n16362;
  assign n16364 = ~n6127 & ~n16031;
  assign n16365 = controllable_hmaster1 & ~n16364;
  assign n16366 = controllable_hmaster0 & ~n16364;
  assign n16367 = controllable_hmaster0 & ~n16366;
  assign n16368 = ~controllable_hmaster1 & ~n16367;
  assign n16369 = ~n16365 & ~n16368;
  assign n16370 = ~i_hbusreq3 & ~n16369;
  assign n16371 = ~n16363 & ~n16370;
  assign n16372 = controllable_hmaster2 & ~n16371;
  assign n16373 = controllable_hmaster2 & ~n16372;
  assign n16374 = ~controllable_hgrant3 & ~n16373;
  assign n16375 = ~n7090 & ~n16374;
  assign n16376 = controllable_nhgrant0 & ~n16375;
  assign n16377 = ~n7118 & ~n16376;
  assign n16378 = ~n3281 & ~n16377;
  assign n16379 = ~n3281 & ~n16378;
  assign n16380 = ~n3378 & ~n16379;
  assign n16381 = ~n16013 & ~n16380;
  assign n16382 = n3492 & ~n16381;
  assign n16383 = n3492 & ~n16382;
  assign n16384 = n3485 & ~n16383;
  assign n16385 = n3485 & ~n16384;
  assign n16386 = ~n3374 & ~n16385;
  assign n16387 = ~n11205 & ~n16070;
  assign n16388 = controllable_hmaster1 & ~n16387;
  assign n16389 = ~n16077 & ~n16388;
  assign n16390 = i_hbusreq3 & ~n16389;
  assign n16391 = ~n11218 & ~n16081;
  assign n16392 = controllable_hmaster1 & ~n16391;
  assign n16393 = ~n16088 & ~n16392;
  assign n16394 = ~i_hbusreq3 & ~n16393;
  assign n16395 = ~n16390 & ~n16394;
  assign n16396 = ~controllable_hmaster2 & ~n16395;
  assign n16397 = ~n16068 & ~n16396;
  assign n16398 = ~controllable_hgrant3 & ~n16397;
  assign n16399 = ~n15646 & ~n16398;
  assign n16400 = controllable_nhgrant0 & ~n16399;
  assign n16401 = ~n15675 & ~n16400;
  assign n16402 = ~n3281 & ~n16401;
  assign n16403 = ~n3281 & ~n16402;
  assign n16404 = n3378 & ~n16403;
  assign n16405 = ~n4787 & ~n12334;
  assign n16406 = ~controllable_hmaster0 & ~n16405;
  assign n16407 = ~n16359 & ~n16406;
  assign n16408 = ~controllable_hmaster1 & ~n16407;
  assign n16409 = ~n16358 & ~n16408;
  assign n16410 = i_hbusreq3 & ~n16409;
  assign n16411 = ~n12345 & ~n16031;
  assign n16412 = ~controllable_hmaster0 & ~n16411;
  assign n16413 = ~n16366 & ~n16412;
  assign n16414 = ~controllable_hmaster1 & ~n16413;
  assign n16415 = ~n16365 & ~n16414;
  assign n16416 = ~i_hbusreq3 & ~n16415;
  assign n16417 = ~n16410 & ~n16416;
  assign n16418 = controllable_hmaster2 & ~n16417;
  assign n16419 = ~n4787 & ~n6252;
  assign n16420 = controllable_hmaster0 & ~n16419;
  assign n16421 = ~n11205 & ~n16420;
  assign n16422 = controllable_hmaster1 & ~n16421;
  assign n16423 = ~n4787 & ~n6266;
  assign n16424 = controllable_hmaster0 & ~n16423;
  assign n16425 = ~controllable_hmaster0 & ~n16419;
  assign n16426 = ~n16424 & ~n16425;
  assign n16427 = ~controllable_hmaster1 & ~n16426;
  assign n16428 = ~n16422 & ~n16427;
  assign n16429 = i_hbusreq3 & ~n16428;
  assign n16430 = ~n6291 & ~n16031;
  assign n16431 = controllable_hmaster0 & ~n16430;
  assign n16432 = ~n11218 & ~n16431;
  assign n16433 = controllable_hmaster1 & ~n16432;
  assign n16434 = ~n6319 & ~n16031;
  assign n16435 = controllable_hmaster0 & ~n16434;
  assign n16436 = ~n6335 & ~n16145;
  assign n16437 = ~controllable_hmaster0 & ~n16436;
  assign n16438 = ~n16435 & ~n16437;
  assign n16439 = ~controllable_hmaster1 & ~n16438;
  assign n16440 = ~n16433 & ~n16439;
  assign n16441 = ~i_hbusreq3 & ~n16440;
  assign n16442 = ~n16429 & ~n16441;
  assign n16443 = ~controllable_hmaster2 & ~n16442;
  assign n16444 = ~n16418 & ~n16443;
  assign n16445 = ~controllable_hgrant3 & ~n16444;
  assign n16446 = ~n15687 & ~n16445;
  assign n16447 = controllable_nhgrant0 & ~n16446;
  assign n16448 = ~n15716 & ~n16447;
  assign n16449 = ~n3281 & ~n16448;
  assign n16450 = ~n3281 & ~n16449;
  assign n16451 = ~n3378 & ~n16450;
  assign n16452 = ~n16404 & ~n16451;
  assign n16453 = n3492 & ~n16452;
  assign n16454 = n3492 & ~n16453;
  assign n16455 = n3485 & ~n16454;
  assign n16456 = n3485 & ~n16455;
  assign n16457 = ~n3476 & ~n16456;
  assign n16458 = ~n11066 & ~n13132;
  assign n16459 = ~controllable_hmaster0 & ~n16458;
  assign n16460 = ~n16209 & ~n16459;
  assign n16461 = controllable_hmaster1 & ~n16460;
  assign n16462 = ~n16218 & ~n16461;
  assign n16463 = i_hbusreq3 & ~n16462;
  assign n16464 = ~n11110 & ~n13143;
  assign n16465 = ~controllable_hmaster0 & ~n16464;
  assign n16466 = ~n16222 & ~n16465;
  assign n16467 = controllable_hmaster1 & ~n16466;
  assign n16468 = ~n16231 & ~n16467;
  assign n16469 = ~i_hbusreq3 & ~n16468;
  assign n16470 = ~n16463 & ~n16469;
  assign n16471 = ~controllable_hmaster2 & ~n16470;
  assign n16472 = ~n16207 & ~n16471;
  assign n16473 = ~controllable_hgrant3 & ~n16472;
  assign n16474 = ~n15734 & ~n16473;
  assign n16475 = controllable_nhgrant0 & ~n16474;
  assign n16476 = ~n15783 & ~n16475;
  assign n16477 = ~n3281 & ~n16476;
  assign n16478 = ~n3281 & ~n16477;
  assign n16479 = n3378 & ~n16478;
  assign n16480 = ~n7796 & ~n10827;
  assign n16481 = controllable_hmaster1 & ~n16480;
  assign n16482 = controllable_hmaster0 & ~n16480;
  assign n16483 = ~n10827 & ~n13161;
  assign n16484 = ~controllable_hmaster0 & ~n16483;
  assign n16485 = ~n16482 & ~n16484;
  assign n16486 = ~controllable_hmaster1 & ~n16485;
  assign n16487 = ~n16481 & ~n16486;
  assign n16488 = i_hbusreq3 & ~n16487;
  assign n16489 = ~n13171 & ~n16274;
  assign n16490 = controllable_hmaster1 & ~n16489;
  assign n16491 = controllable_hmaster0 & ~n16489;
  assign n16492 = ~n13179 & ~n16274;
  assign n16493 = ~controllable_hmaster0 & ~n16492;
  assign n16494 = ~n16491 & ~n16493;
  assign n16495 = ~controllable_hmaster1 & ~n16494;
  assign n16496 = ~n16490 & ~n16495;
  assign n16497 = ~i_hbusreq3 & ~n16496;
  assign n16498 = ~n16488 & ~n16497;
  assign n16499 = controllable_hmaster2 & ~n16498;
  assign n16500 = ~n7861 & ~n10827;
  assign n16501 = controllable_hmaster0 & ~n16500;
  assign n16502 = ~n11066 & ~n13189;
  assign n16503 = ~controllable_hmaster0 & ~n16502;
  assign n16504 = ~n16501 & ~n16503;
  assign n16505 = controllable_hmaster1 & ~n16504;
  assign n16506 = ~n7872 & ~n10827;
  assign n16507 = controllable_hmaster0 & ~n16506;
  assign n16508 = ~controllable_hmaster0 & ~n16500;
  assign n16509 = ~n16507 & ~n16508;
  assign n16510 = ~controllable_hmaster1 & ~n16509;
  assign n16511 = ~n16505 & ~n16510;
  assign n16512 = i_hbusreq3 & ~n16511;
  assign n16513 = ~n13206 & ~n16274;
  assign n16514 = controllable_hmaster0 & ~n16513;
  assign n16515 = ~n11110 & ~n13200;
  assign n16516 = ~controllable_hmaster0 & ~n16515;
  assign n16517 = ~n16514 & ~n16516;
  assign n16518 = controllable_hmaster1 & ~n16517;
  assign n16519 = ~n13214 & ~n16274;
  assign n16520 = controllable_hmaster0 & ~n16519;
  assign n16521 = ~n13220 & ~n16330;
  assign n16522 = ~controllable_hmaster0 & ~n16521;
  assign n16523 = ~n16520 & ~n16522;
  assign n16524 = ~controllable_hmaster1 & ~n16523;
  assign n16525 = ~n16518 & ~n16524;
  assign n16526 = ~i_hbusreq3 & ~n16525;
  assign n16527 = ~n16512 & ~n16526;
  assign n16528 = ~controllable_hmaster2 & ~n16527;
  assign n16529 = ~n16499 & ~n16528;
  assign n16530 = ~controllable_hgrant3 & ~n16529;
  assign n16531 = ~n15795 & ~n16530;
  assign n16532 = controllable_nhgrant0 & ~n16531;
  assign n16533 = ~n15846 & ~n16532;
  assign n16534 = ~n3281 & ~n16533;
  assign n16535 = ~n3281 & ~n16534;
  assign n16536 = ~n3378 & ~n16535;
  assign n16537 = ~n16479 & ~n16536;
  assign n16538 = n3492 & ~n16537;
  assign n16539 = ~n14836 & ~n16538;
  assign n16540 = n3485 & ~n16539;
  assign n16541 = ~n14835 & ~n16540;
  assign n16542 = n3476 & ~n16541;
  assign n16543 = ~n16457 & ~n16542;
  assign n16544 = n3374 & ~n16543;
  assign n16545 = ~n16386 & ~n16544;
  assign n16546 = ~n3655 & ~n16545;
  assign n16547 = ~n16356 & ~n16546;
  assign n16548 = ~n3652 & ~n16547;
  assign n16549 = ~n15977 & ~n16548;
  assign n16550 = n3368 & ~n16549;
  assign n16551 = ~n15638 & ~n16550;
  assign n16552 = n3362 & ~n16551;
  assign n16553 = n3492 & ~n15027;
  assign n16554 = ~n3631 & ~n16553;
  assign n16555 = n3485 & ~n16554;
  assign n16556 = ~n3630 & ~n16555;
  assign n16557 = ~n3476 & ~n16556;
  assign n16558 = n3492 & ~n15111;
  assign n16559 = ~n3631 & ~n16558;
  assign n16560 = n3485 & ~n16559;
  assign n16561 = ~n8312 & ~n16560;
  assign n16562 = n3476 & ~n16561;
  assign n16563 = ~n16557 & ~n16562;
  assign n16564 = n3374 & ~n16563;
  assign n16565 = ~n8316 & ~n16564;
  assign n16566 = n3655 & ~n16565;
  assign n16567 = n3492 & ~n15163;
  assign n16568 = ~n3631 & ~n16567;
  assign n16569 = n3485 & ~n16568;
  assign n16570 = ~n3630 & ~n16569;
  assign n16571 = ~n3476 & ~n16570;
  assign n16572 = n3492 & ~n15211;
  assign n16573 = ~n3631 & ~n16572;
  assign n16574 = n3485 & ~n16573;
  assign n16575 = ~n8369 & ~n16574;
  assign n16576 = n3476 & ~n16575;
  assign n16577 = ~n16571 & ~n16576;
  assign n16578 = n3374 & ~n16577;
  assign n16579 = ~n8373 & ~n16578;
  assign n16580 = ~n3655 & ~n16579;
  assign n16581 = ~n16566 & ~n16580;
  assign n16582 = n3652 & ~n16581;
  assign n16583 = n3492 & ~n15249;
  assign n16584 = ~n3631 & ~n16583;
  assign n16585 = n3485 & ~n16584;
  assign n16586 = ~n3630 & ~n16585;
  assign n16587 = ~n3476 & ~n16586;
  assign n16588 = n3492 & ~n14429;
  assign n16589 = ~n8434 & ~n16588;
  assign n16590 = ~n3485 & ~n16589;
  assign n16591 = ~n15258 & ~n16583;
  assign n16592 = n3485 & ~n16591;
  assign n16593 = ~n16590 & ~n16592;
  assign n16594 = n3476 & ~n16593;
  assign n16595 = ~n16587 & ~n16594;
  assign n16596 = ~n3374 & ~n16595;
  assign n16597 = n3492 & ~n15349;
  assign n16598 = ~n3631 & ~n16597;
  assign n16599 = n3485 & ~n16598;
  assign n16600 = ~n3630 & ~n16599;
  assign n16601 = ~n3476 & ~n16600;
  assign n16602 = n3492 & ~n15461;
  assign n16603 = ~n15258 & ~n16602;
  assign n16604 = n3485 & ~n16603;
  assign n16605 = ~n16590 & ~n16604;
  assign n16606 = n3476 & ~n16605;
  assign n16607 = ~n16601 & ~n16606;
  assign n16608 = n3374 & ~n16607;
  assign n16609 = ~n16596 & ~n16608;
  assign n16610 = n3655 & ~n16609;
  assign n16611 = n3492 & ~n15495;
  assign n16612 = ~n3631 & ~n16611;
  assign n16613 = n3485 & ~n16612;
  assign n16614 = ~n3630 & ~n16613;
  assign n16615 = ~n3476 & ~n16614;
  assign n16616 = ~n8491 & ~n16588;
  assign n16617 = ~n3485 & ~n16616;
  assign n16618 = ~n15258 & ~n16611;
  assign n16619 = n3485 & ~n16618;
  assign n16620 = ~n16617 & ~n16619;
  assign n16621 = n3476 & ~n16620;
  assign n16622 = ~n16615 & ~n16621;
  assign n16623 = ~n3374 & ~n16622;
  assign n16624 = n3492 & ~n15559;
  assign n16625 = ~n3631 & ~n16624;
  assign n16626 = n3485 & ~n16625;
  assign n16627 = ~n3630 & ~n16626;
  assign n16628 = ~n3476 & ~n16627;
  assign n16629 = n3492 & ~n15623;
  assign n16630 = ~n15258 & ~n16629;
  assign n16631 = n3485 & ~n16630;
  assign n16632 = ~n16617 & ~n16631;
  assign n16633 = n3476 & ~n16632;
  assign n16634 = ~n16628 & ~n16633;
  assign n16635 = n3374 & ~n16634;
  assign n16636 = ~n16623 & ~n16635;
  assign n16637 = ~n3655 & ~n16636;
  assign n16638 = ~n16610 & ~n16637;
  assign n16639 = ~n3652 & ~n16638;
  assign n16640 = ~n16582 & ~n16639;
  assign n16641 = ~n3368 & ~n16640;
  assign n16642 = n3492 & ~n15719;
  assign n16643 = n3492 & ~n16642;
  assign n16644 = n3485 & ~n16643;
  assign n16645 = n3485 & ~n16644;
  assign n16646 = ~n3476 & ~n16645;
  assign n16647 = n3492 & ~n15849;
  assign n16648 = n3492 & ~n16647;
  assign n16649 = n3485 & ~n16648;
  assign n16650 = ~n8538 & ~n16649;
  assign n16651 = n3476 & ~n16650;
  assign n16652 = ~n16646 & ~n16651;
  assign n16653 = n3374 & ~n16652;
  assign n16654 = ~n8529 & ~n16653;
  assign n16655 = n3655 & ~n16654;
  assign n16656 = n3492 & ~n15895;
  assign n16657 = n3492 & ~n16656;
  assign n16658 = n3485 & ~n16657;
  assign n16659 = n3485 & ~n16658;
  assign n16660 = ~n3476 & ~n16659;
  assign n16661 = n3492 & ~n15964;
  assign n16662 = n3492 & ~n16661;
  assign n16663 = n3485 & ~n16662;
  assign n16664 = ~n8565 & ~n16663;
  assign n16665 = n3476 & ~n16664;
  assign n16666 = ~n16660 & ~n16665;
  assign n16667 = n3374 & ~n16666;
  assign n16668 = ~n8556 & ~n16667;
  assign n16669 = ~n3655 & ~n16668;
  assign n16670 = ~n16655 & ~n16669;
  assign n16671 = n3652 & ~n16670;
  assign n16672 = n3492 & ~n16047;
  assign n16673 = n3492 & ~n16672;
  assign n16674 = n3485 & ~n16673;
  assign n16675 = n3485 & ~n16674;
  assign n16676 = ~n3476 & ~n16675;
  assign n16677 = ~n8525 & ~n16674;
  assign n16678 = n3476 & ~n16677;
  assign n16679 = ~n16676 & ~n16678;
  assign n16680 = ~n3374 & ~n16679;
  assign n16681 = n3492 & ~n16160;
  assign n16682 = n3492 & ~n16681;
  assign n16683 = n3485 & ~n16682;
  assign n16684 = n3485 & ~n16683;
  assign n16685 = ~n3476 & ~n16684;
  assign n16686 = n3492 & ~n14382;
  assign n16687 = ~n8592 & ~n16686;
  assign n16688 = ~n3485 & ~n16687;
  assign n16689 = n3492 & ~n16345;
  assign n16690 = ~n14836 & ~n16689;
  assign n16691 = n3485 & ~n16690;
  assign n16692 = ~n16688 & ~n16691;
  assign n16693 = n3476 & ~n16692;
  assign n16694 = ~n16685 & ~n16693;
  assign n16695 = n3374 & ~n16694;
  assign n16696 = ~n16680 & ~n16695;
  assign n16697 = n3655 & ~n16696;
  assign n16698 = n3492 & ~n16379;
  assign n16699 = n3492 & ~n16698;
  assign n16700 = n3485 & ~n16699;
  assign n16701 = n3485 & ~n16700;
  assign n16702 = ~n3476 & ~n16701;
  assign n16703 = ~n8525 & ~n16700;
  assign n16704 = n3476 & ~n16703;
  assign n16705 = ~n16702 & ~n16704;
  assign n16706 = ~n3374 & ~n16705;
  assign n16707 = n3492 & ~n16450;
  assign n16708 = n3492 & ~n16707;
  assign n16709 = n3485 & ~n16708;
  assign n16710 = n3485 & ~n16709;
  assign n16711 = ~n3476 & ~n16710;
  assign n16712 = ~n8619 & ~n16686;
  assign n16713 = ~n3485 & ~n16712;
  assign n16714 = n3492 & ~n16535;
  assign n16715 = ~n14836 & ~n16714;
  assign n16716 = n3485 & ~n16715;
  assign n16717 = ~n16713 & ~n16716;
  assign n16718 = n3476 & ~n16717;
  assign n16719 = ~n16711 & ~n16718;
  assign n16720 = n3374 & ~n16719;
  assign n16721 = ~n16706 & ~n16720;
  assign n16722 = ~n3655 & ~n16721;
  assign n16723 = ~n16697 & ~n16722;
  assign n16724 = ~n3652 & ~n16723;
  assign n16725 = ~n16671 & ~n16724;
  assign n16726 = n3368 & ~n16725;
  assign n16727 = ~n16641 & ~n16726;
  assign n16728 = ~n3362 & ~n16727;
  assign n16729 = ~n16552 & ~n16728;
  assign n16730 = n3359 & ~n16729;
  assign n16731 = ~n8639 & ~n16560;
  assign n16732 = n3476 & ~n16731;
  assign n16733 = ~n16557 & ~n16732;
  assign n16734 = n3374 & ~n16733;
  assign n16735 = ~n8643 & ~n16734;
  assign n16736 = n3655 & ~n16735;
  assign n16737 = ~n8650 & ~n16574;
  assign n16738 = n3476 & ~n16737;
  assign n16739 = ~n16571 & ~n16738;
  assign n16740 = n3374 & ~n16739;
  assign n16741 = ~n8654 & ~n16740;
  assign n16742 = ~n3655 & ~n16741;
  assign n16743 = ~n16736 & ~n16742;
  assign n16744 = n3652 & ~n16743;
  assign n16745 = ~n8663 & ~n16592;
  assign n16746 = n3476 & ~n16745;
  assign n16747 = ~n16587 & ~n16746;
  assign n16748 = ~n3374 & ~n16747;
  assign n16749 = ~n8663 & ~n16604;
  assign n16750 = n3476 & ~n16749;
  assign n16751 = ~n16601 & ~n16750;
  assign n16752 = n3374 & ~n16751;
  assign n16753 = ~n16748 & ~n16752;
  assign n16754 = n3655 & ~n16753;
  assign n16755 = ~n8674 & ~n16619;
  assign n16756 = n3476 & ~n16755;
  assign n16757 = ~n16615 & ~n16756;
  assign n16758 = ~n3374 & ~n16757;
  assign n16759 = ~n8674 & ~n16631;
  assign n16760 = n3476 & ~n16759;
  assign n16761 = ~n16628 & ~n16760;
  assign n16762 = n3374 & ~n16761;
  assign n16763 = ~n16758 & ~n16762;
  assign n16764 = ~n3655 & ~n16763;
  assign n16765 = ~n16754 & ~n16764;
  assign n16766 = ~n3652 & ~n16765;
  assign n16767 = ~n16744 & ~n16766;
  assign n16768 = ~n3368 & ~n16767;
  assign n16769 = ~n8694 & ~n16649;
  assign n16770 = n3476 & ~n16769;
  assign n16771 = ~n16646 & ~n16770;
  assign n16772 = n3374 & ~n16771;
  assign n16773 = ~n8693 & ~n16772;
  assign n16774 = n3655 & ~n16773;
  assign n16775 = ~n8705 & ~n16663;
  assign n16776 = n3476 & ~n16775;
  assign n16777 = ~n16660 & ~n16776;
  assign n16778 = n3374 & ~n16777;
  assign n16779 = ~n8704 & ~n16778;
  assign n16780 = ~n3655 & ~n16779;
  assign n16781 = ~n16774 & ~n16780;
  assign n16782 = n3652 & ~n16781;
  assign n16783 = ~n8689 & ~n16674;
  assign n16784 = n3476 & ~n16783;
  assign n16785 = ~n16676 & ~n16784;
  assign n16786 = ~n3374 & ~n16785;
  assign n16787 = ~n8718 & ~n16691;
  assign n16788 = n3476 & ~n16787;
  assign n16789 = ~n16685 & ~n16788;
  assign n16790 = n3374 & ~n16789;
  assign n16791 = ~n16786 & ~n16790;
  assign n16792 = n3655 & ~n16791;
  assign n16793 = ~n8689 & ~n16700;
  assign n16794 = n3476 & ~n16793;
  assign n16795 = ~n16702 & ~n16794;
  assign n16796 = ~n3374 & ~n16795;
  assign n16797 = ~n8729 & ~n16716;
  assign n16798 = n3476 & ~n16797;
  assign n16799 = ~n16711 & ~n16798;
  assign n16800 = n3374 & ~n16799;
  assign n16801 = ~n16796 & ~n16800;
  assign n16802 = ~n3655 & ~n16801;
  assign n16803 = ~n16792 & ~n16802;
  assign n16804 = ~n3652 & ~n16803;
  assign n16805 = ~n16782 & ~n16804;
  assign n16806 = n3368 & ~n16805;
  assign n16807 = ~n16768 & ~n16806;
  assign n16808 = n3362 & ~n16807;
  assign n16809 = n3378 & ~n15027;
  assign n16810 = ~n8906 & ~n16809;
  assign n16811 = n3492 & ~n16810;
  assign n16812 = ~n3631 & ~n16811;
  assign n16813 = n3485 & ~n16812;
  assign n16814 = ~n3630 & ~n16813;
  assign n16815 = ~n3476 & ~n16814;
  assign n16816 = n3378 & ~n15111;
  assign n16817 = ~n9100 & ~n16816;
  assign n16818 = n3492 & ~n16817;
  assign n16819 = ~n8309 & ~n16818;
  assign n16820 = n3485 & ~n16819;
  assign n16821 = ~n8639 & ~n16820;
  assign n16822 = n3476 & ~n16821;
  assign n16823 = ~n16815 & ~n16822;
  assign n16824 = n3374 & ~n16823;
  assign n16825 = ~n8801 & ~n16824;
  assign n16826 = n3655 & ~n16825;
  assign n16827 = n3378 & ~n15163;
  assign n16828 = ~n9240 & ~n16827;
  assign n16829 = n3492 & ~n16828;
  assign n16830 = ~n3631 & ~n16829;
  assign n16831 = n3485 & ~n16830;
  assign n16832 = ~n3630 & ~n16831;
  assign n16833 = ~n3476 & ~n16832;
  assign n16834 = n3378 & ~n15211;
  assign n16835 = ~n9374 & ~n16834;
  assign n16836 = n3492 & ~n16835;
  assign n16837 = ~n8367 & ~n16836;
  assign n16838 = n3485 & ~n16837;
  assign n16839 = ~n8650 & ~n16838;
  assign n16840 = n3476 & ~n16839;
  assign n16841 = ~n16833 & ~n16840;
  assign n16842 = n3374 & ~n16841;
  assign n16843 = ~n9147 & ~n16842;
  assign n16844 = ~n3655 & ~n16843;
  assign n16845 = ~n16826 & ~n16844;
  assign n16846 = n3652 & ~n16845;
  assign n16847 = n3378 & ~n15249;
  assign n16848 = ~n9409 & ~n16847;
  assign n16849 = n3492 & ~n16848;
  assign n16850 = ~n3631 & ~n16849;
  assign n16851 = n3485 & ~n16850;
  assign n16852 = ~n3630 & ~n16851;
  assign n16853 = ~n3476 & ~n16852;
  assign n16854 = ~n8434 & ~n16849;
  assign n16855 = n3485 & ~n16854;
  assign n16856 = ~n8663 & ~n16855;
  assign n16857 = n3476 & ~n16856;
  assign n16858 = ~n16853 & ~n16857;
  assign n16859 = ~n3374 & ~n16858;
  assign n16860 = n3378 & ~n15349;
  assign n16861 = ~n9469 & ~n16860;
  assign n16862 = n3492 & ~n16861;
  assign n16863 = ~n3631 & ~n16862;
  assign n16864 = n3485 & ~n16863;
  assign n16865 = ~n3630 & ~n16864;
  assign n16866 = ~n3476 & ~n16865;
  assign n16867 = n3378 & ~n15461;
  assign n16868 = ~n9531 & ~n16867;
  assign n16869 = n3492 & ~n16868;
  assign n16870 = ~n8434 & ~n16869;
  assign n16871 = n3485 & ~n16870;
  assign n16872 = ~n8663 & ~n16871;
  assign n16873 = n3476 & ~n16872;
  assign n16874 = ~n16866 & ~n16873;
  assign n16875 = n3374 & ~n16874;
  assign n16876 = ~n16859 & ~n16875;
  assign n16877 = n3655 & ~n16876;
  assign n16878 = n3378 & ~n15495;
  assign n16879 = ~n9563 & ~n16878;
  assign n16880 = n3492 & ~n16879;
  assign n16881 = ~n3631 & ~n16880;
  assign n16882 = n3485 & ~n16881;
  assign n16883 = ~n3630 & ~n16882;
  assign n16884 = ~n3476 & ~n16883;
  assign n16885 = ~n8491 & ~n16880;
  assign n16886 = n3485 & ~n16885;
  assign n16887 = ~n8674 & ~n16886;
  assign n16888 = n3476 & ~n16887;
  assign n16889 = ~n16884 & ~n16888;
  assign n16890 = ~n3374 & ~n16889;
  assign n16891 = n3378 & ~n15559;
  assign n16892 = ~n9623 & ~n16891;
  assign n16893 = n3492 & ~n16892;
  assign n16894 = ~n3631 & ~n16893;
  assign n16895 = n3485 & ~n16894;
  assign n16896 = ~n3630 & ~n16895;
  assign n16897 = ~n3476 & ~n16896;
  assign n16898 = n3378 & ~n15623;
  assign n16899 = ~n9683 & ~n16898;
  assign n16900 = n3492 & ~n16899;
  assign n16901 = ~n8491 & ~n16900;
  assign n16902 = n3485 & ~n16901;
  assign n16903 = ~n8674 & ~n16902;
  assign n16904 = n3476 & ~n16903;
  assign n16905 = ~n16897 & ~n16904;
  assign n16906 = n3374 & ~n16905;
  assign n16907 = ~n16890 & ~n16906;
  assign n16908 = ~n3655 & ~n16907;
  assign n16909 = ~n16877 & ~n16908;
  assign n16910 = ~n3652 & ~n16909;
  assign n16911 = ~n16846 & ~n16910;
  assign n16912 = ~n3368 & ~n16911;
  assign n16913 = n3378 & ~n15719;
  assign n16914 = ~n9865 & ~n16913;
  assign n16915 = n3492 & ~n16914;
  assign n16916 = n3492 & ~n16915;
  assign n16917 = n3485 & ~n16916;
  assign n16918 = n3485 & ~n16917;
  assign n16919 = ~n3476 & ~n16918;
  assign n16920 = ~n13799 & ~n15796;
  assign n16921 = controllable_hmaster1 & ~n16920;
  assign n16922 = controllable_hmaster0 & ~n16920;
  assign n16923 = ~n12266 & ~n15796;
  assign n16924 = ~controllable_hmaster0 & ~n16923;
  assign n16925 = ~n16922 & ~n16924;
  assign n16926 = ~controllable_hmaster1 & ~n16925;
  assign n16927 = ~n16921 & ~n16926;
  assign n16928 = ~i_hbusreq3 & ~n16927;
  assign n16929 = ~n13795 & ~n16928;
  assign n16930 = controllable_hmaster2 & ~n16929;
  assign n16931 = ~n5947 & ~n15796;
  assign n16932 = controllable_hmaster0 & ~n16931;
  assign n16933 = ~n10152 & ~n13812;
  assign n16934 = ~controllable_hmaster0 & ~n16933;
  assign n16935 = ~n16932 & ~n16934;
  assign n16936 = controllable_hmaster1 & ~n16935;
  assign n16937 = ~n5978 & ~n15796;
  assign n16938 = controllable_hmaster0 & ~n16937;
  assign n16939 = ~n5994 & ~n15822;
  assign n16940 = ~controllable_hmaster0 & ~n16939;
  assign n16941 = ~n16938 & ~n16940;
  assign n16942 = ~controllable_hmaster1 & ~n16941;
  assign n16943 = ~n16936 & ~n16942;
  assign n16944 = ~i_hbusreq3 & ~n16943;
  assign n16945 = ~n15096 & ~n16944;
  assign n16946 = ~controllable_hmaster2 & ~n16945;
  assign n16947 = ~n16930 & ~n16946;
  assign n16948 = ~controllable_hgrant3 & ~n16947;
  assign n16949 = ~n15795 & ~n16948;
  assign n16950 = controllable_nhgrant0 & ~n16949;
  assign n16951 = controllable_hmaster1 & ~n9978;
  assign n16952 = ~n10042 & ~n16951;
  assign n16953 = i_hbusreq3 & ~n16952;
  assign n16954 = controllable_hmaster1 & ~n10023;
  assign n16955 = ~n10063 & ~n16954;
  assign n16956 = ~i_hbusreq3 & ~n16955;
  assign n16957 = ~n16953 & ~n16956;
  assign n16958 = ~controllable_hmaster2 & ~n16957;
  assign n16959 = ~n13828 & ~n16958;
  assign n16960 = ~controllable_hgrant3 & ~n16959;
  assign n16961 = ~n15704 & ~n16960;
  assign n16962 = ~controllable_nhgrant0 & ~n16961;
  assign n16963 = ~n16950 & ~n16962;
  assign n16964 = ~n3281 & ~n16963;
  assign n16965 = ~n3281 & ~n16964;
  assign n16966 = n3378 & ~n16965;
  assign n16967 = ~n10244 & ~n16966;
  assign n16968 = n3492 & ~n16967;
  assign n16969 = ~n8536 & ~n16968;
  assign n16970 = n3485 & ~n16969;
  assign n16971 = ~n8694 & ~n16970;
  assign n16972 = n3476 & ~n16971;
  assign n16973 = ~n16919 & ~n16972;
  assign n16974 = n3374 & ~n16973;
  assign n16975 = ~n9769 & ~n16974;
  assign n16976 = n3655 & ~n16975;
  assign n16977 = n3378 & ~n15895;
  assign n16978 = ~n10390 & ~n16977;
  assign n16979 = n3492 & ~n16978;
  assign n16980 = n3492 & ~n16979;
  assign n16981 = n3485 & ~n16980;
  assign n16982 = n3485 & ~n16981;
  assign n16983 = ~n3476 & ~n16982;
  assign n16984 = ~n13878 & ~n15796;
  assign n16985 = controllable_hmaster1 & ~n16984;
  assign n16986 = controllable_hmaster0 & ~n16984;
  assign n16987 = ~n13886 & ~n15796;
  assign n16988 = ~controllable_hmaster0 & ~n16987;
  assign n16989 = ~n16986 & ~n16988;
  assign n16990 = ~controllable_hmaster1 & ~n16989;
  assign n16991 = ~n16985 & ~n16990;
  assign n16992 = ~i_hbusreq3 & ~n16991;
  assign n16993 = ~n13874 & ~n16992;
  assign n16994 = controllable_hmaster2 & ~n16993;
  assign n16995 = ~n10487 & ~n10634;
  assign n16996 = controllable_hmaster1 & ~n16995;
  assign n16997 = ~n10505 & ~n16996;
  assign n16998 = i_hbusreq3 & ~n16997;
  assign n16999 = ~n13908 & ~n15796;
  assign n17000 = controllable_hmaster0 & ~n16999;
  assign n17001 = ~n10152 & ~n13902;
  assign n17002 = ~controllable_hmaster0 & ~n17001;
  assign n17003 = ~n17000 & ~n17002;
  assign n17004 = controllable_hmaster1 & ~n17003;
  assign n17005 = ~n13916 & ~n15796;
  assign n17006 = controllable_hmaster0 & ~n17005;
  assign n17007 = ~n13922 & ~n15822;
  assign n17008 = ~controllable_hmaster0 & ~n17007;
  assign n17009 = ~n17006 & ~n17008;
  assign n17010 = ~controllable_hmaster1 & ~n17009;
  assign n17011 = ~n17004 & ~n17010;
  assign n17012 = ~i_hbusreq3 & ~n17011;
  assign n17013 = ~n16998 & ~n17012;
  assign n17014 = ~controllable_hmaster2 & ~n17013;
  assign n17015 = ~n16994 & ~n17014;
  assign n17016 = ~controllable_hgrant3 & ~n17015;
  assign n17017 = ~n15795 & ~n17016;
  assign n17018 = controllable_nhgrant0 & ~n17017;
  assign n17019 = ~n16962 & ~n17018;
  assign n17020 = ~n3281 & ~n17019;
  assign n17021 = ~n3281 & ~n17020;
  assign n17022 = n3378 & ~n17021;
  assign n17023 = ~n10705 & ~n17022;
  assign n17024 = n3492 & ~n17023;
  assign n17025 = ~n8563 & ~n17024;
  assign n17026 = n3485 & ~n17025;
  assign n17027 = ~n8705 & ~n17026;
  assign n17028 = n3476 & ~n17027;
  assign n17029 = ~n16983 & ~n17028;
  assign n17030 = n3374 & ~n17029;
  assign n17031 = ~n10311 & ~n17030;
  assign n17032 = ~n3655 & ~n17031;
  assign n17033 = ~n16976 & ~n17032;
  assign n17034 = n3652 & ~n17033;
  assign n17035 = n3378 & ~n16047;
  assign n17036 = ~n10742 & ~n17035;
  assign n17037 = n3492 & ~n17036;
  assign n17038 = n3492 & ~n17037;
  assign n17039 = n3485 & ~n17038;
  assign n17040 = n3485 & ~n17039;
  assign n17041 = ~n3476 & ~n17040;
  assign n17042 = ~n8523 & ~n17037;
  assign n17043 = n3485 & ~n17042;
  assign n17044 = ~n8689 & ~n17043;
  assign n17045 = n3476 & ~n17044;
  assign n17046 = ~n17041 & ~n17045;
  assign n17047 = ~n3374 & ~n17046;
  assign n17048 = n3378 & ~n16160;
  assign n17049 = ~n10802 & ~n17048;
  assign n17050 = n3492 & ~n17049;
  assign n17051 = n3492 & ~n17050;
  assign n17052 = n3485 & ~n17051;
  assign n17053 = n3485 & ~n17052;
  assign n17054 = ~n3476 & ~n17053;
  assign n17055 = ~n9875 & ~n10827;
  assign n17056 = controllable_hmaster1 & ~n17055;
  assign n17057 = controllable_hmaster0 & ~n17055;
  assign n17058 = ~n10827 & ~n12255;
  assign n17059 = ~controllable_hmaster0 & ~n17058;
  assign n17060 = ~n17057 & ~n17059;
  assign n17061 = ~controllable_hmaster1 & ~n17060;
  assign n17062 = ~n17056 & ~n17061;
  assign n17063 = i_hbusreq3 & ~n17062;
  assign n17064 = ~n13799 & ~n16274;
  assign n17065 = controllable_hmaster1 & ~n17064;
  assign n17066 = controllable_hmaster0 & ~n17064;
  assign n17067 = ~n12266 & ~n16274;
  assign n17068 = ~controllable_hmaster0 & ~n17067;
  assign n17069 = ~n17066 & ~n17068;
  assign n17070 = ~controllable_hmaster1 & ~n17069;
  assign n17071 = ~n17065 & ~n17070;
  assign n17072 = ~i_hbusreq3 & ~n17071;
  assign n17073 = ~n17063 & ~n17072;
  assign n17074 = controllable_hmaster2 & ~n17073;
  assign n17075 = ~n5913 & ~n10827;
  assign n17076 = controllable_hmaster0 & ~n17075;
  assign n17077 = ~n11068 & ~n17076;
  assign n17078 = controllable_hmaster1 & ~n17077;
  assign n17079 = ~n5923 & ~n10827;
  assign n17080 = controllable_hmaster0 & ~n17079;
  assign n17081 = ~controllable_hmaster0 & ~n17075;
  assign n17082 = ~n17080 & ~n17081;
  assign n17083 = ~controllable_hmaster1 & ~n17082;
  assign n17084 = ~n17078 & ~n17083;
  assign n17085 = i_hbusreq3 & ~n17084;
  assign n17086 = ~n5947 & ~n16274;
  assign n17087 = controllable_hmaster0 & ~n17086;
  assign n17088 = ~n11110 & ~n13812;
  assign n17089 = ~controllable_hmaster0 & ~n17088;
  assign n17090 = ~n17087 & ~n17089;
  assign n17091 = controllable_hmaster1 & ~n17090;
  assign n17092 = ~n5978 & ~n16274;
  assign n17093 = controllable_hmaster0 & ~n17092;
  assign n17094 = ~n5994 & ~n16330;
  assign n17095 = ~controllable_hmaster0 & ~n17094;
  assign n17096 = ~n17093 & ~n17095;
  assign n17097 = ~controllable_hmaster1 & ~n17096;
  assign n17098 = ~n17091 & ~n17097;
  assign n17099 = ~i_hbusreq3 & ~n17098;
  assign n17100 = ~n17085 & ~n17099;
  assign n17101 = ~controllable_hmaster2 & ~n17100;
  assign n17102 = ~n17074 & ~n17101;
  assign n17103 = ~controllable_hgrant3 & ~n17102;
  assign n17104 = ~n15795 & ~n17103;
  assign n17105 = controllable_nhgrant0 & ~n17104;
  assign n17106 = ~n16962 & ~n17105;
  assign n17107 = ~n3281 & ~n17106;
  assign n17108 = ~n3281 & ~n17107;
  assign n17109 = n3378 & ~n17108;
  assign n17110 = ~n11143 & ~n17109;
  assign n17111 = n3492 & ~n17110;
  assign n17112 = ~n8592 & ~n17111;
  assign n17113 = n3485 & ~n17112;
  assign n17114 = ~n8718 & ~n17113;
  assign n17115 = n3476 & ~n17114;
  assign n17116 = ~n17054 & ~n17115;
  assign n17117 = n3374 & ~n17116;
  assign n17118 = ~n17047 & ~n17117;
  assign n17119 = n3655 & ~n17118;
  assign n17120 = n3378 & ~n16379;
  assign n17121 = ~n11178 & ~n17120;
  assign n17122 = n3492 & ~n17121;
  assign n17123 = n3492 & ~n17122;
  assign n17124 = n3485 & ~n17123;
  assign n17125 = n3485 & ~n17124;
  assign n17126 = ~n3476 & ~n17125;
  assign n17127 = ~n8523 & ~n17122;
  assign n17128 = n3485 & ~n17127;
  assign n17129 = ~n8689 & ~n17128;
  assign n17130 = n3476 & ~n17129;
  assign n17131 = ~n17126 & ~n17130;
  assign n17132 = ~n3374 & ~n17131;
  assign n17133 = n3378 & ~n16450;
  assign n17134 = ~n11236 & ~n17133;
  assign n17135 = n3492 & ~n17134;
  assign n17136 = n3492 & ~n17135;
  assign n17137 = n3485 & ~n17136;
  assign n17138 = n3485 & ~n17137;
  assign n17139 = ~n3476 & ~n17138;
  assign n17140 = ~n10406 & ~n10827;
  assign n17141 = controllable_hmaster1 & ~n17140;
  assign n17142 = controllable_hmaster0 & ~n17140;
  assign n17143 = ~n10827 & ~n13868;
  assign n17144 = ~controllable_hmaster0 & ~n17143;
  assign n17145 = ~n17142 & ~n17144;
  assign n17146 = ~controllable_hmaster1 & ~n17145;
  assign n17147 = ~n17141 & ~n17146;
  assign n17148 = i_hbusreq3 & ~n17147;
  assign n17149 = ~n13878 & ~n16274;
  assign n17150 = controllable_hmaster1 & ~n17149;
  assign n17151 = controllable_hmaster0 & ~n17149;
  assign n17152 = ~n13886 & ~n16274;
  assign n17153 = ~controllable_hmaster0 & ~n17152;
  assign n17154 = ~n17151 & ~n17153;
  assign n17155 = ~controllable_hmaster1 & ~n17154;
  assign n17156 = ~n17150 & ~n17155;
  assign n17157 = ~i_hbusreq3 & ~n17156;
  assign n17158 = ~n17148 & ~n17157;
  assign n17159 = controllable_hmaster2 & ~n17158;
  assign n17160 = ~n10485 & ~n10827;
  assign n17161 = controllable_hmaster0 & ~n17160;
  assign n17162 = ~n11319 & ~n17161;
  assign n17163 = controllable_hmaster1 & ~n17162;
  assign n17164 = ~n10500 & ~n10827;
  assign n17165 = controllable_hmaster0 & ~n17164;
  assign n17166 = ~controllable_hmaster0 & ~n17160;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = ~controllable_hmaster1 & ~n17167;
  assign n17169 = ~n17163 & ~n17168;
  assign n17170 = i_hbusreq3 & ~n17169;
  assign n17171 = ~n13908 & ~n16274;
  assign n17172 = controllable_hmaster0 & ~n17171;
  assign n17173 = ~n11110 & ~n13902;
  assign n17174 = ~controllable_hmaster0 & ~n17173;
  assign n17175 = ~n17172 & ~n17174;
  assign n17176 = controllable_hmaster1 & ~n17175;
  assign n17177 = ~n13916 & ~n16274;
  assign n17178 = controllable_hmaster0 & ~n17177;
  assign n17179 = ~n13922 & ~n16330;
  assign n17180 = ~controllable_hmaster0 & ~n17179;
  assign n17181 = ~n17178 & ~n17180;
  assign n17182 = ~controllable_hmaster1 & ~n17181;
  assign n17183 = ~n17176 & ~n17182;
  assign n17184 = ~i_hbusreq3 & ~n17183;
  assign n17185 = ~n17170 & ~n17184;
  assign n17186 = ~controllable_hmaster2 & ~n17185;
  assign n17187 = ~n17159 & ~n17186;
  assign n17188 = ~controllable_hgrant3 & ~n17187;
  assign n17189 = ~n15795 & ~n17188;
  assign n17190 = controllable_nhgrant0 & ~n17189;
  assign n17191 = ~n16962 & ~n17190;
  assign n17192 = ~n3281 & ~n17191;
  assign n17193 = ~n3281 & ~n17192;
  assign n17194 = n3378 & ~n17193;
  assign n17195 = ~n11352 & ~n17194;
  assign n17196 = n3492 & ~n17195;
  assign n17197 = ~n8619 & ~n17196;
  assign n17198 = n3485 & ~n17197;
  assign n17199 = ~n8729 & ~n17198;
  assign n17200 = n3476 & ~n17199;
  assign n17201 = ~n17139 & ~n17200;
  assign n17202 = n3374 & ~n17201;
  assign n17203 = ~n17132 & ~n17202;
  assign n17204 = ~n3655 & ~n17203;
  assign n17205 = ~n17119 & ~n17204;
  assign n17206 = ~n3652 & ~n17205;
  assign n17207 = ~n17034 & ~n17206;
  assign n17208 = n3368 & ~n17207;
  assign n17209 = ~n16912 & ~n17208;
  assign n17210 = ~n3362 & ~n17209;
  assign n17211 = ~n16808 & ~n17210;
  assign n17212 = ~n3359 & ~n17211;
  assign n17213 = ~n16730 & ~n17212;
  assign n17214 = ~n3356 & ~n17213;
  assign n17215 = ~n14958 & ~n17214;
  assign n17216 = n3345 & ~n17215;
  assign n17217 = ~n14086 & ~n17216;
  assign n17218 = n3341 & ~n17217;
  assign n17219 = ~n11376 & ~n17218;
  assign n17220 = ~n3337 & ~n17219;
  assign n17221 = controllable_hmaster0 & ~n4940;
  assign n17222 = ~controllable_hmaster1 & ~n17221;
  assign n17223 = ~controllable_hmaster1 & ~n17222;
  assign n17224 = i_hbusreq3 & ~n17223;
  assign n17225 = controllable_hmaster0 & ~n5007;
  assign n17226 = ~controllable_hmaster1 & ~n17225;
  assign n17227 = ~controllable_hmaster1 & ~n17226;
  assign n17228 = ~i_hbusreq3 & ~n17227;
  assign n17229 = ~n17224 & ~n17228;
  assign n17230 = ~controllable_hmaster2 & ~n17229;
  assign n17231 = ~controllable_hmaster2 & ~n17230;
  assign n17232 = controllable_hgrant3 & ~n17231;
  assign n17233 = controllable_hmaster0 & ~n5103;
  assign n17234 = ~controllable_hmaster1 & ~n17233;
  assign n17235 = ~controllable_hmaster1 & ~n17234;
  assign n17236 = i_hbusreq3 & ~n17235;
  assign n17237 = controllable_hmaster0 & ~n5148;
  assign n17238 = ~controllable_hmaster1 & ~n17237;
  assign n17239 = ~controllable_hmaster1 & ~n17238;
  assign n17240 = ~i_hbusreq3 & ~n17239;
  assign n17241 = ~n17236 & ~n17240;
  assign n17242 = ~controllable_hmaster2 & ~n17241;
  assign n17243 = ~controllable_hmaster2 & ~n17242;
  assign n17244 = ~controllable_hgrant3 & ~n17243;
  assign n17245 = ~n17232 & ~n17244;
  assign n17246 = controllable_nhgrant0 & ~n17245;
  assign n17247 = ~controllable_nhgrant0 & ~n17231;
  assign n17248 = ~n17246 & ~n17247;
  assign n17249 = ~n3281 & ~n17248;
  assign n17250 = ~n3281 & ~n17249;
  assign n17251 = n3378 & ~n17250;
  assign n17252 = ~n3407 & ~n17230;
  assign n17253 = controllable_hgrant3 & ~n17252;
  assign n17254 = ~n3461 & ~n17242;
  assign n17255 = ~controllable_hgrant3 & ~n17254;
  assign n17256 = ~n17253 & ~n17255;
  assign n17257 = controllable_nhgrant0 & ~n17256;
  assign n17258 = ~controllable_nhgrant0 & ~n17252;
  assign n17259 = ~n17257 & ~n17258;
  assign n17260 = ~n3281 & ~n17259;
  assign n17261 = ~n3783 & ~n17260;
  assign n17262 = ~n3378 & ~n17261;
  assign n17263 = ~n17251 & ~n17262;
  assign n17264 = n3492 & ~n17263;
  assign n17265 = ~n3493 & ~n17264;
  assign n17266 = n3485 & ~n17265;
  assign n17267 = ~n3486 & ~n17266;
  assign n17268 = ~n3374 & ~n17267;
  assign n17269 = ~controllable_hmaster1 & ~n3384;
  assign n17270 = i_hbusreq3 & ~n17269;
  assign n17271 = ~controllable_hmaster1 & ~n7084;
  assign n17272 = ~i_hbusreq3 & ~n17271;
  assign n17273 = ~n17270 & ~n17272;
  assign n17274 = ~controllable_hmaster2 & ~n17273;
  assign n17275 = ~controllable_hmaster2 & ~n17274;
  assign n17276 = controllable_hgrant3 & ~n17275;
  assign n17277 = controllable_hmaster0 & ~n8826;
  assign n17278 = ~controllable_hmaster1 & ~n17277;
  assign n17279 = ~controllable_hmaster1 & ~n17278;
  assign n17280 = i_hbusreq3 & ~n17279;
  assign n17281 = controllable_hmaster0 & ~n8860;
  assign n17282 = ~controllable_hmaster1 & ~n17281;
  assign n17283 = ~controllable_hmaster1 & ~n17282;
  assign n17284 = ~i_hbusreq3 & ~n17283;
  assign n17285 = ~n17280 & ~n17284;
  assign n17286 = ~controllable_hmaster2 & ~n17285;
  assign n17287 = ~controllable_hmaster2 & ~n17286;
  assign n17288 = ~controllable_hgrant3 & ~n17287;
  assign n17289 = ~n17276 & ~n17288;
  assign n17290 = controllable_nhgrant0 & ~n17289;
  assign n17291 = ~controllable_hmaster1 & ~n7106;
  assign n17292 = i_hbusreq3 & ~n17291;
  assign n17293 = ~controllable_hmaster1 & ~n7110;
  assign n17294 = ~i_hbusreq3 & ~n17293;
  assign n17295 = ~n17292 & ~n17294;
  assign n17296 = ~controllable_hmaster2 & ~n17295;
  assign n17297 = ~controllable_hmaster2 & ~n17296;
  assign n17298 = ~controllable_hgrant3 & ~n17297;
  assign n17299 = ~n17276 & ~n17298;
  assign n17300 = ~controllable_nhgrant0 & ~n17299;
  assign n17301 = ~n17290 & ~n17300;
  assign n17302 = ~n3281 & ~n17301;
  assign n17303 = ~n3281 & ~n17302;
  assign n17304 = n3378 & ~n17303;
  assign n17305 = ~n3407 & ~n17274;
  assign n17306 = controllable_hgrant3 & ~n17305;
  assign n17307 = ~n3530 & ~n17286;
  assign n17308 = ~controllable_hgrant3 & ~n17307;
  assign n17309 = ~n17306 & ~n17308;
  assign n17310 = controllable_nhgrant0 & ~n17309;
  assign n17311 = ~n3407 & ~n17296;
  assign n17312 = ~controllable_hgrant3 & ~n17311;
  assign n17313 = ~n17306 & ~n17312;
  assign n17314 = ~controllable_nhgrant0 & ~n17313;
  assign n17315 = ~n17310 & ~n17314;
  assign n17316 = ~n3281 & ~n17315;
  assign n17317 = ~n3950 & ~n17316;
  assign n17318 = ~n3378 & ~n17317;
  assign n17319 = ~n17304 & ~n17318;
  assign n17320 = n3492 & ~n17319;
  assign n17321 = ~n3493 & ~n17320;
  assign n17322 = n3485 & ~n17321;
  assign n17323 = ~n3486 & ~n17322;
  assign n17324 = ~n3476 & ~n17323;
  assign n17325 = controllable_hgrant1 & ~n4178;
  assign n17326 = ~controllable_ndecide & ~n17325;
  assign n17327 = ~controllable_ndecide & ~n17326;
  assign n17328 = i_hready & ~n17327;
  assign n17329 = i_hready & ~n17328;
  assign n17330 = ~controllable_hgrant4 & ~n17329;
  assign n17331 = ~controllable_hgrant4 & ~n17330;
  assign n17332 = ~controllable_hgrant2 & ~n17331;
  assign n17333 = ~controllable_hgrant2 & ~n17332;
  assign n17334 = i_hbusreq3 & ~n17333;
  assign n17335 = i_hbusreq2 & ~n17331;
  assign n17336 = i_hbusreq4 & ~n17329;
  assign n17337 = i_hbusreq0 & ~n17329;
  assign n17338 = i_hbusreq1 & ~n17325;
  assign n17339 = i_hbusreq1 & ~n17338;
  assign n17340 = ~controllable_ndecide & ~n17339;
  assign n17341 = ~controllable_ndecide & ~n17340;
  assign n17342 = i_hready & ~n17341;
  assign n17343 = i_hready & ~n17342;
  assign n17344 = i_hlock0 & ~n17343;
  assign n17345 = ~i_hlock0 & ~n17329;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~i_hbusreq0 & ~n17346;
  assign n17348 = ~n17337 & ~n17347;
  assign n17349 = ~i_hbusreq4 & ~n17348;
  assign n17350 = ~n17336 & ~n17349;
  assign n17351 = ~controllable_hgrant4 & ~n17350;
  assign n17352 = ~controllable_hgrant4 & ~n17351;
  assign n17353 = ~i_hbusreq2 & ~n17352;
  assign n17354 = ~n17335 & ~n17353;
  assign n17355 = ~controllable_hgrant2 & ~n17354;
  assign n17356 = ~controllable_hgrant2 & ~n17355;
  assign n17357 = ~i_hbusreq3 & ~n17356;
  assign n17358 = ~n17334 & ~n17357;
  assign n17359 = controllable_hmaster2 & ~n17358;
  assign n17360 = controllable_hmaster1 & ~n17333;
  assign n17361 = ~controllable_ndecide & ~n5691;
  assign n17362 = ~controllable_ndecide & ~n17361;
  assign n17363 = i_hready & ~n17362;
  assign n17364 = ~n3495 & ~n17363;
  assign n17365 = ~controllable_hgrant4 & ~n17364;
  assign n17366 = ~n3411 & ~n17365;
  assign n17367 = ~controllable_hgrant2 & ~n17366;
  assign n17368 = ~n3410 & ~n17367;
  assign n17369 = controllable_hmaster0 & ~n17368;
  assign n17370 = ~controllable_hmaster0 & ~n17333;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = ~controllable_hmaster1 & ~n17371;
  assign n17373 = ~n17360 & ~n17372;
  assign n17374 = i_hbusreq3 & ~n17373;
  assign n17375 = controllable_hmaster1 & ~n17356;
  assign n17376 = i_hbusreq2 & ~n17366;
  assign n17377 = i_hbusreq4 & ~n17364;
  assign n17378 = i_hbusreq0 & ~n17364;
  assign n17379 = i_hbusreq1 & n5691;
  assign n17380 = ~controllable_ndecide & ~n17379;
  assign n17381 = ~controllable_ndecide & ~n17380;
  assign n17382 = i_hready & ~n17381;
  assign n17383 = ~n3511 & ~n17382;
  assign n17384 = i_hlock0 & ~n17383;
  assign n17385 = ~i_hlock0 & ~n17364;
  assign n17386 = ~n17384 & ~n17385;
  assign n17387 = ~i_hbusreq0 & ~n17386;
  assign n17388 = ~n17378 & ~n17387;
  assign n17389 = ~i_hbusreq4 & ~n17388;
  assign n17390 = ~n17377 & ~n17389;
  assign n17391 = ~controllable_hgrant4 & ~n17390;
  assign n17392 = ~n3916 & ~n17391;
  assign n17393 = ~i_hbusreq2 & ~n17392;
  assign n17394 = ~n17376 & ~n17393;
  assign n17395 = ~controllable_hgrant2 & ~n17394;
  assign n17396 = ~n3859 & ~n17395;
  assign n17397 = controllable_hmaster0 & ~n17396;
  assign n17398 = ~controllable_hmaster0 & ~n17356;
  assign n17399 = ~n17397 & ~n17398;
  assign n17400 = ~controllable_hmaster1 & ~n17399;
  assign n17401 = ~n17375 & ~n17400;
  assign n17402 = ~i_hbusreq3 & ~n17401;
  assign n17403 = ~n17374 & ~n17402;
  assign n17404 = ~controllable_hmaster2 & ~n17403;
  assign n17405 = ~n17359 & ~n17404;
  assign n17406 = ~controllable_hgrant3 & ~n17405;
  assign n17407 = ~n17276 & ~n17406;
  assign n17408 = controllable_nhgrant0 & ~n17407;
  assign n17409 = ~n17300 & ~n17408;
  assign n17410 = ~n3281 & ~n17409;
  assign n17411 = ~n3281 & ~n17410;
  assign n17412 = n3378 & ~n17411;
  assign n17413 = ~n3411 & ~n5621;
  assign n17414 = ~controllable_hgrant2 & ~n17413;
  assign n17415 = ~n3410 & ~n17414;
  assign n17416 = controllable_hmaster1 & ~n17415;
  assign n17417 = controllable_hmaster0 & ~n17415;
  assign n17418 = i_hready & ~n5619;
  assign n17419 = ~controllable_hgrant4 & ~n17418;
  assign n17420 = ~controllable_hgrant4 & ~n17419;
  assign n17421 = ~controllable_hgrant2 & ~n17420;
  assign n17422 = ~controllable_hgrant2 & ~n17421;
  assign n17423 = ~controllable_hmaster0 & ~n17422;
  assign n17424 = ~n17417 & ~n17423;
  assign n17425 = ~controllable_hmaster1 & ~n17424;
  assign n17426 = ~n17416 & ~n17425;
  assign n17427 = i_hbusreq3 & ~n17426;
  assign n17428 = i_hbusreq2 & ~n17413;
  assign n17429 = ~i_hbusreq1 & ~n17325;
  assign n17430 = ~n5639 & ~n17429;
  assign n17431 = ~controllable_ndecide & ~n17430;
  assign n17432 = ~n3494 & ~n17431;
  assign n17433 = i_hready & ~n17432;
  assign n17434 = ~n3511 & ~n17433;
  assign n17435 = ~i_hlock0 & ~n17434;
  assign n17436 = ~n5659 & ~n17435;
  assign n17437 = ~i_hbusreq0 & ~n17436;
  assign n17438 = ~n5638 & ~n17437;
  assign n17439 = ~i_hbusreq4 & ~n17438;
  assign n17440 = ~n5637 & ~n17439;
  assign n17441 = ~controllable_hgrant4 & ~n17440;
  assign n17442 = ~n3433 & ~n17441;
  assign n17443 = ~i_hbusreq2 & ~n17442;
  assign n17444 = ~n17428 & ~n17443;
  assign n17445 = ~controllable_hgrant2 & ~n17444;
  assign n17446 = ~n3431 & ~n17445;
  assign n17447 = controllable_hmaster1 & ~n17446;
  assign n17448 = controllable_hmaster0 & ~n17446;
  assign n17449 = i_hbusreq2 & ~n17420;
  assign n17450 = i_hbusreq4 & ~n17418;
  assign n17451 = i_hbusreq0 & ~n17418;
  assign n17452 = i_hready & ~n5643;
  assign n17453 = i_hlock0 & ~n17452;
  assign n17454 = i_hready & ~n17433;
  assign n17455 = ~i_hlock0 & ~n17454;
  assign n17456 = ~n17453 & ~n17455;
  assign n17457 = ~i_hbusreq0 & ~n17456;
  assign n17458 = ~n17451 & ~n17457;
  assign n17459 = ~i_hbusreq4 & ~n17458;
  assign n17460 = ~n17450 & ~n17459;
  assign n17461 = ~controllable_hgrant4 & ~n17460;
  assign n17462 = ~controllable_hgrant4 & ~n17461;
  assign n17463 = ~i_hbusreq2 & ~n17462;
  assign n17464 = ~n17449 & ~n17463;
  assign n17465 = ~controllable_hgrant2 & ~n17464;
  assign n17466 = ~controllable_hgrant2 & ~n17465;
  assign n17467 = ~controllable_hmaster0 & ~n17466;
  assign n17468 = ~n17448 & ~n17467;
  assign n17469 = ~controllable_hmaster1 & ~n17468;
  assign n17470 = ~n17447 & ~n17469;
  assign n17471 = ~i_hbusreq3 & ~n17470;
  assign n17472 = ~n17427 & ~n17471;
  assign n17473 = controllable_hmaster2 & ~n17472;
  assign n17474 = controllable_hmaster1 & ~n17422;
  assign n17475 = ~n3411 & ~n8987;
  assign n17476 = ~controllable_hgrant2 & ~n17475;
  assign n17477 = ~n3410 & ~n17476;
  assign n17478 = controllable_hmaster0 & ~n17477;
  assign n17479 = ~n17423 & ~n17478;
  assign n17480 = ~controllable_hmaster1 & ~n17479;
  assign n17481 = ~n17474 & ~n17480;
  assign n17482 = i_hbusreq3 & ~n17481;
  assign n17483 = controllable_hmaster1 & ~n17466;
  assign n17484 = i_hbusreq2 & ~n17475;
  assign n17485 = ~n3511 & ~n5733;
  assign n17486 = i_hlock0 & ~n17485;
  assign n17487 = ~i_hbusreq1 & n5691;
  assign n17488 = ~n5730 & ~n17487;
  assign n17489 = ~controllable_ndecide & n17488;
  assign n17490 = ~n3494 & ~n17489;
  assign n17491 = i_hready & ~n17490;
  assign n17492 = ~n3495 & ~n17491;
  assign n17493 = ~i_hlock0 & ~n17492;
  assign n17494 = ~n17486 & ~n17493;
  assign n17495 = ~i_hbusreq0 & ~n17494;
  assign n17496 = ~n9009 & ~n17495;
  assign n17497 = ~i_hbusreq4 & ~n17496;
  assign n17498 = ~n9008 & ~n17497;
  assign n17499 = ~controllable_hgrant4 & ~n17498;
  assign n17500 = ~n3916 & ~n17499;
  assign n17501 = ~i_hbusreq2 & ~n17500;
  assign n17502 = ~n17484 & ~n17501;
  assign n17503 = ~controllable_hgrant2 & ~n17502;
  assign n17504 = ~n3859 & ~n17503;
  assign n17505 = controllable_hmaster0 & ~n17504;
  assign n17506 = ~n17467 & ~n17505;
  assign n17507 = ~controllable_hmaster1 & ~n17506;
  assign n17508 = ~n17483 & ~n17507;
  assign n17509 = ~i_hbusreq3 & ~n17508;
  assign n17510 = ~n17482 & ~n17509;
  assign n17511 = ~controllable_hmaster2 & ~n17510;
  assign n17512 = ~n17473 & ~n17511;
  assign n17513 = ~controllable_hgrant3 & ~n17512;
  assign n17514 = ~n17306 & ~n17513;
  assign n17515 = controllable_nhgrant0 & ~n17514;
  assign n17516 = ~n17314 & ~n17515;
  assign n17517 = ~n3281 & ~n17516;
  assign n17518 = ~n4089 & ~n17517;
  assign n17519 = ~n3378 & ~n17518;
  assign n17520 = ~n17412 & ~n17519;
  assign n17521 = n3492 & ~n17520;
  assign n17522 = ~n3493 & ~n17521;
  assign n17523 = n3485 & ~n17522;
  assign n17524 = ~n3486 & ~n17523;
  assign n17525 = n3476 & ~n17524;
  assign n17526 = ~n17324 & ~n17525;
  assign n17527 = n3374 & ~n17526;
  assign n17528 = ~n17268 & ~n17527;
  assign n17529 = n3655 & ~n17528;
  assign n17530 = controllable_hmaster0 & ~n6149;
  assign n17531 = ~controllable_hmaster1 & ~n17530;
  assign n17532 = ~controllable_hmaster1 & ~n17531;
  assign n17533 = i_hbusreq3 & ~n17532;
  assign n17534 = controllable_hmaster0 & ~n6178;
  assign n17535 = ~controllable_hmaster1 & ~n17534;
  assign n17536 = ~controllable_hmaster1 & ~n17535;
  assign n17537 = ~i_hbusreq3 & ~n17536;
  assign n17538 = ~n17533 & ~n17537;
  assign n17539 = ~controllable_hmaster2 & ~n17538;
  assign n17540 = ~controllable_hmaster2 & ~n17539;
  assign n17541 = ~controllable_hgrant3 & ~n17540;
  assign n17542 = ~n17232 & ~n17541;
  assign n17543 = controllable_nhgrant0 & ~n17542;
  assign n17544 = ~n17247 & ~n17543;
  assign n17545 = ~n3281 & ~n17544;
  assign n17546 = ~n3281 & ~n17545;
  assign n17547 = n3378 & ~n17546;
  assign n17548 = ~controllable_hgrant1 & ~n3414;
  assign n17549 = ~controllable_hgrant1 & ~n17548;
  assign n17550 = controllable_ndecide & ~n17549;
  assign n17551 = controllable_ndecide & ~n17550;
  assign n17552 = ~i_hready & n17551;
  assign n17553 = ~n3417 & ~n17552;
  assign n17554 = ~controllable_hgrant4 & ~n17553;
  assign n17555 = ~n3411 & ~n17554;
  assign n17556 = ~controllable_hgrant2 & ~n17555;
  assign n17557 = ~n3410 & ~n17556;
  assign n17558 = controllable_hmaster1 & ~n17557;
  assign n17559 = controllable_hmaster0 & ~n17557;
  assign n17560 = controllable_hmaster0 & ~n17559;
  assign n17561 = ~controllable_hmaster1 & ~n17560;
  assign n17562 = ~n17558 & ~n17561;
  assign n17563 = i_hbusreq3 & ~n17562;
  assign n17564 = i_hbusreq2 & ~n17555;
  assign n17565 = i_hbusreq4 & ~n17553;
  assign n17566 = i_hbusreq0 & ~n17553;
  assign n17567 = ~n6304 & ~n17550;
  assign n17568 = ~i_hready & n17567;
  assign n17569 = ~n3440 & ~n17568;
  assign n17570 = ~i_hbusreq0 & ~n17569;
  assign n17571 = ~n17566 & ~n17570;
  assign n17572 = ~i_hbusreq4 & ~n17571;
  assign n17573 = ~n17565 & ~n17572;
  assign n17574 = ~controllable_hgrant4 & ~n17573;
  assign n17575 = ~n3433 & ~n17574;
  assign n17576 = ~i_hbusreq2 & ~n17575;
  assign n17577 = ~n17564 & ~n17576;
  assign n17578 = ~controllable_hgrant2 & ~n17577;
  assign n17579 = ~n3431 & ~n17578;
  assign n17580 = controllable_hmaster1 & ~n17579;
  assign n17581 = controllable_hmaster0 & ~n17579;
  assign n17582 = controllable_hmaster0 & ~n17581;
  assign n17583 = ~controllable_hmaster1 & ~n17582;
  assign n17584 = ~n17580 & ~n17583;
  assign n17585 = ~i_hbusreq3 & ~n17584;
  assign n17586 = ~n17563 & ~n17585;
  assign n17587 = controllable_hmaster2 & ~n17586;
  assign n17588 = ~n17539 & ~n17587;
  assign n17589 = ~controllable_hgrant3 & ~n17588;
  assign n17590 = ~n17253 & ~n17589;
  assign n17591 = controllable_nhgrant0 & ~n17590;
  assign n17592 = ~n17258 & ~n17591;
  assign n17593 = ~n3281 & ~n17592;
  assign n17594 = ~n3783 & ~n17593;
  assign n17595 = ~n3378 & ~n17594;
  assign n17596 = ~n17547 & ~n17595;
  assign n17597 = n3492 & ~n17596;
  assign n17598 = ~n3493 & ~n17597;
  assign n17599 = n3485 & ~n17598;
  assign n17600 = ~n3486 & ~n17599;
  assign n17601 = ~n3476 & ~n17600;
  assign n17602 = ~n3461 & ~n17539;
  assign n17603 = ~controllable_hgrant3 & ~n17602;
  assign n17604 = ~n17253 & ~n17603;
  assign n17605 = controllable_nhgrant0 & ~n17604;
  assign n17606 = ~n17258 & ~n17605;
  assign n17607 = ~n3281 & ~n17606;
  assign n17608 = ~n3783 & ~n17607;
  assign n17609 = ~n3378 & ~n17608;
  assign n17610 = ~n17547 & ~n17609;
  assign n17611 = ~n3485 & ~n17610;
  assign n17612 = ~n3492 & ~n17610;
  assign n17613 = ~n17597 & ~n17612;
  assign n17614 = n3485 & ~n17613;
  assign n17615 = ~n17611 & ~n17614;
  assign n17616 = n3476 & ~n17615;
  assign n17617 = ~n17601 & ~n17616;
  assign n17618 = ~n3374 & ~n17617;
  assign n17619 = controllable_hmaster0 & ~n9174;
  assign n17620 = ~controllable_hmaster1 & ~n17619;
  assign n17621 = ~controllable_hmaster1 & ~n17620;
  assign n17622 = i_hbusreq3 & ~n17621;
  assign n17623 = controllable_hmaster0 & ~n9210;
  assign n17624 = ~controllable_hmaster1 & ~n17623;
  assign n17625 = ~controllable_hmaster1 & ~n17624;
  assign n17626 = ~i_hbusreq3 & ~n17625;
  assign n17627 = ~n17622 & ~n17626;
  assign n17628 = ~controllable_hmaster2 & ~n17627;
  assign n17629 = ~controllable_hmaster2 & ~n17628;
  assign n17630 = ~controllable_hgrant3 & ~n17629;
  assign n17631 = ~n17276 & ~n17630;
  assign n17632 = controllable_nhgrant0 & ~n17631;
  assign n17633 = ~n17300 & ~n17632;
  assign n17634 = ~n3281 & ~n17633;
  assign n17635 = ~n3281 & ~n17634;
  assign n17636 = n3378 & ~n17635;
  assign n17637 = controllable_hmaster0 & ~n9117;
  assign n17638 = ~controllable_hmaster1 & ~n17637;
  assign n17639 = ~n9116 & ~n17638;
  assign n17640 = i_hbusreq3 & ~n17639;
  assign n17641 = i_hbusreq2 & ~n9113;
  assign n17642 = i_hbusreq4 & n3417;
  assign n17643 = i_hbusreq0 & n3417;
  assign n17644 = ~controllable_ndecide & ~n6304;
  assign n17645 = ~i_hready & n17644;
  assign n17646 = ~n3440 & ~n17645;
  assign n17647 = ~i_hbusreq0 & ~n17646;
  assign n17648 = ~n17643 & ~n17647;
  assign n17649 = ~i_hbusreq4 & ~n17648;
  assign n17650 = ~n17642 & ~n17649;
  assign n17651 = ~controllable_hgrant4 & ~n17650;
  assign n17652 = ~n3433 & ~n17651;
  assign n17653 = ~i_hbusreq2 & ~n17652;
  assign n17654 = ~n17641 & ~n17653;
  assign n17655 = ~controllable_hgrant2 & ~n17654;
  assign n17656 = ~n3431 & ~n17655;
  assign n17657 = controllable_hmaster1 & ~n17656;
  assign n17658 = controllable_hmaster0 & ~n17656;
  assign n17659 = controllable_hmaster0 & ~n17658;
  assign n17660 = ~controllable_hmaster1 & ~n17659;
  assign n17661 = ~n17657 & ~n17660;
  assign n17662 = ~i_hbusreq3 & ~n17661;
  assign n17663 = ~n17640 & ~n17662;
  assign n17664 = controllable_hmaster2 & ~n17663;
  assign n17665 = ~n17628 & ~n17664;
  assign n17666 = ~controllable_hgrant3 & ~n17665;
  assign n17667 = ~n17306 & ~n17666;
  assign n17668 = controllable_nhgrant0 & ~n17667;
  assign n17669 = ~n17314 & ~n17668;
  assign n17670 = ~n3281 & ~n17669;
  assign n17671 = ~n3950 & ~n17670;
  assign n17672 = ~n3378 & ~n17671;
  assign n17673 = ~n17636 & ~n17672;
  assign n17674 = n3492 & ~n17673;
  assign n17675 = ~n3493 & ~n17674;
  assign n17676 = n3485 & ~n17675;
  assign n17677 = ~n3486 & ~n17676;
  assign n17678 = ~n3476 & ~n17677;
  assign n17679 = i_hready & ~n17325;
  assign n17680 = i_hready & ~n17679;
  assign n17681 = ~controllable_hgrant4 & ~n17680;
  assign n17682 = ~controllable_hgrant4 & ~n17681;
  assign n17683 = ~controllable_hgrant2 & ~n17682;
  assign n17684 = ~controllable_hgrant2 & ~n17683;
  assign n17685 = i_hbusreq3 & ~n17684;
  assign n17686 = i_hbusreq2 & ~n17682;
  assign n17687 = i_hbusreq4 & ~n17680;
  assign n17688 = i_hbusreq0 & ~n17680;
  assign n17689 = controllable_ndecide & ~n17325;
  assign n17690 = ~n17340 & ~n17689;
  assign n17691 = i_hready & ~n17690;
  assign n17692 = i_hready & ~n17691;
  assign n17693 = i_hlock0 & ~n17692;
  assign n17694 = ~i_hlock0 & ~n17680;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = ~i_hbusreq0 & ~n17695;
  assign n17697 = ~n17688 & ~n17696;
  assign n17698 = ~i_hbusreq4 & ~n17697;
  assign n17699 = ~n17687 & ~n17698;
  assign n17700 = ~controllable_hgrant4 & ~n17699;
  assign n17701 = ~controllable_hgrant4 & ~n17700;
  assign n17702 = ~i_hbusreq2 & ~n17701;
  assign n17703 = ~n17686 & ~n17702;
  assign n17704 = ~controllable_hgrant2 & ~n17703;
  assign n17705 = ~controllable_hgrant2 & ~n17704;
  assign n17706 = ~i_hbusreq3 & ~n17705;
  assign n17707 = ~n17685 & ~n17706;
  assign n17708 = controllable_hmaster2 & ~n17707;
  assign n17709 = controllable_hmaster1 & ~n17684;
  assign n17710 = i_hready & n5691;
  assign n17711 = ~n9168 & ~n17710;
  assign n17712 = ~controllable_hgrant4 & n17711;
  assign n17713 = ~n3411 & ~n17712;
  assign n17714 = ~controllable_hgrant2 & ~n17713;
  assign n17715 = ~n3410 & ~n17714;
  assign n17716 = controllable_hmaster0 & ~n17715;
  assign n17717 = ~controllable_hmaster0 & ~n17684;
  assign n17718 = ~n17716 & ~n17717;
  assign n17719 = ~controllable_hmaster1 & ~n17718;
  assign n17720 = ~n17709 & ~n17719;
  assign n17721 = i_hbusreq3 & ~n17720;
  assign n17722 = controllable_hmaster1 & ~n17705;
  assign n17723 = i_hbusreq2 & ~n17713;
  assign n17724 = i_hbusreq4 & ~n17711;
  assign n17725 = i_hbusreq0 & ~n17711;
  assign n17726 = controllable_ndecide & n5691;
  assign n17727 = ~controllable_ndecide & n17379;
  assign n17728 = ~n17726 & ~n17727;
  assign n17729 = i_hready & ~n17728;
  assign n17730 = ~n9195 & ~n17729;
  assign n17731 = i_hlock0 & ~n17730;
  assign n17732 = ~i_hlock0 & ~n17711;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = ~i_hbusreq0 & ~n17733;
  assign n17735 = ~n17725 & ~n17734;
  assign n17736 = ~i_hbusreq4 & ~n17735;
  assign n17737 = ~n17724 & ~n17736;
  assign n17738 = ~controllable_hgrant4 & n17737;
  assign n17739 = ~n3916 & ~n17738;
  assign n17740 = ~i_hbusreq2 & ~n17739;
  assign n17741 = ~n17723 & ~n17740;
  assign n17742 = ~controllable_hgrant2 & ~n17741;
  assign n17743 = ~n3859 & ~n17742;
  assign n17744 = controllable_hmaster0 & ~n17743;
  assign n17745 = ~controllable_hmaster0 & ~n17705;
  assign n17746 = ~n17744 & ~n17745;
  assign n17747 = ~controllable_hmaster1 & ~n17746;
  assign n17748 = ~n17722 & ~n17747;
  assign n17749 = ~i_hbusreq3 & ~n17748;
  assign n17750 = ~n17721 & ~n17749;
  assign n17751 = ~controllable_hmaster2 & ~n17750;
  assign n17752 = ~n17708 & ~n17751;
  assign n17753 = ~controllable_hgrant3 & ~n17752;
  assign n17754 = ~n17276 & ~n17753;
  assign n17755 = controllable_nhgrant0 & ~n17754;
  assign n17756 = ~n17300 & ~n17755;
  assign n17757 = ~n3281 & ~n17756;
  assign n17758 = ~n3281 & ~n17757;
  assign n17759 = n3378 & ~n17758;
  assign n17760 = ~n3411 & ~n9248;
  assign n17761 = ~controllable_hgrant2 & ~n17760;
  assign n17762 = ~n3410 & ~n17761;
  assign n17763 = controllable_hmaster1 & ~n17762;
  assign n17764 = controllable_hmaster0 & ~n17762;
  assign n17765 = i_hready & ~n6401;
  assign n17766 = ~controllable_hgrant4 & ~n17765;
  assign n17767 = ~controllable_hgrant4 & ~n17766;
  assign n17768 = ~controllable_hgrant2 & ~n17767;
  assign n17769 = ~controllable_hgrant2 & ~n17768;
  assign n17770 = ~controllable_hmaster0 & ~n17769;
  assign n17771 = ~n17764 & ~n17770;
  assign n17772 = ~controllable_hmaster1 & ~n17771;
  assign n17773 = ~n17763 & ~n17772;
  assign n17774 = i_hbusreq3 & ~n17773;
  assign n17775 = i_hbusreq2 & ~n17760;
  assign n17776 = ~n6421 & ~n17645;
  assign n17777 = i_hlock0 & ~n17776;
  assign n17778 = ~n4179 & ~n17431;
  assign n17779 = i_hready & ~n17778;
  assign n17780 = ~n17645 & ~n17779;
  assign n17781 = ~i_hlock0 & ~n17780;
  assign n17782 = ~n17777 & ~n17781;
  assign n17783 = ~i_hbusreq0 & ~n17782;
  assign n17784 = ~n9260 & ~n17783;
  assign n17785 = ~i_hbusreq4 & ~n17784;
  assign n17786 = ~n9259 & ~n17785;
  assign n17787 = ~controllable_hgrant4 & ~n17786;
  assign n17788 = ~n3433 & ~n17787;
  assign n17789 = ~i_hbusreq2 & ~n17788;
  assign n17790 = ~n17775 & ~n17789;
  assign n17791 = ~controllable_hgrant2 & ~n17790;
  assign n17792 = ~n3431 & ~n17791;
  assign n17793 = controllable_hmaster1 & ~n17792;
  assign n17794 = controllable_hmaster0 & ~n17792;
  assign n17795 = i_hbusreq2 & ~n17767;
  assign n17796 = i_hbusreq4 & ~n17765;
  assign n17797 = i_hbusreq0 & ~n17765;
  assign n17798 = i_hready & ~n6421;
  assign n17799 = i_hlock0 & ~n17798;
  assign n17800 = i_hready & ~n17779;
  assign n17801 = ~i_hlock0 & ~n17800;
  assign n17802 = ~n17799 & ~n17801;
  assign n17803 = ~i_hbusreq0 & ~n17802;
  assign n17804 = ~n17797 & ~n17803;
  assign n17805 = ~i_hbusreq4 & ~n17804;
  assign n17806 = ~n17796 & ~n17805;
  assign n17807 = ~controllable_hgrant4 & ~n17806;
  assign n17808 = ~controllable_hgrant4 & ~n17807;
  assign n17809 = ~i_hbusreq2 & ~n17808;
  assign n17810 = ~n17795 & ~n17809;
  assign n17811 = ~controllable_hgrant2 & ~n17810;
  assign n17812 = ~controllable_hgrant2 & ~n17811;
  assign n17813 = ~controllable_hmaster0 & ~n17812;
  assign n17814 = ~n17794 & ~n17813;
  assign n17815 = ~controllable_hmaster1 & ~n17814;
  assign n17816 = ~n17793 & ~n17815;
  assign n17817 = ~i_hbusreq3 & ~n17816;
  assign n17818 = ~n17774 & ~n17817;
  assign n17819 = controllable_hmaster2 & ~n17818;
  assign n17820 = controllable_hmaster1 & ~n17769;
  assign n17821 = ~n3411 & ~n9305;
  assign n17822 = ~controllable_hgrant2 & ~n17821;
  assign n17823 = ~n3410 & ~n17822;
  assign n17824 = controllable_hmaster0 & ~n17823;
  assign n17825 = ~n17770 & ~n17824;
  assign n17826 = ~controllable_hmaster1 & ~n17825;
  assign n17827 = ~n17820 & ~n17826;
  assign n17828 = i_hbusreq3 & ~n17827;
  assign n17829 = controllable_hmaster1 & ~n17812;
  assign n17830 = i_hbusreq2 & ~n17821;
  assign n17831 = ~n6515 & ~n9195;
  assign n17832 = i_hlock0 & ~n17831;
  assign n17833 = ~controllable_ndecide & ~n17488;
  assign n17834 = ~n6512 & ~n17833;
  assign n17835 = i_hready & ~n17834;
  assign n17836 = ~n9168 & ~n17835;
  assign n17837 = ~i_hlock0 & ~n17836;
  assign n17838 = ~n17832 & ~n17837;
  assign n17839 = ~i_hbusreq0 & ~n17838;
  assign n17840 = ~n9327 & ~n17839;
  assign n17841 = ~i_hbusreq4 & ~n17840;
  assign n17842 = ~n9326 & ~n17841;
  assign n17843 = ~controllable_hgrant4 & n17842;
  assign n17844 = ~n3916 & ~n17843;
  assign n17845 = ~i_hbusreq2 & ~n17844;
  assign n17846 = ~n17830 & ~n17845;
  assign n17847 = ~controllable_hgrant2 & ~n17846;
  assign n17848 = ~n3859 & ~n17847;
  assign n17849 = controllable_hmaster0 & ~n17848;
  assign n17850 = ~n17813 & ~n17849;
  assign n17851 = ~controllable_hmaster1 & ~n17850;
  assign n17852 = ~n17829 & ~n17851;
  assign n17853 = ~i_hbusreq3 & ~n17852;
  assign n17854 = ~n17828 & ~n17853;
  assign n17855 = ~controllable_hmaster2 & ~n17854;
  assign n17856 = ~n17819 & ~n17855;
  assign n17857 = ~controllable_hgrant3 & ~n17856;
  assign n17858 = ~n17306 & ~n17857;
  assign n17859 = controllable_nhgrant0 & ~n17858;
  assign n17860 = ~n17314 & ~n17859;
  assign n17861 = ~n3281 & ~n17860;
  assign n17862 = ~n4089 & ~n17861;
  assign n17863 = ~n3378 & ~n17862;
  assign n17864 = ~n17759 & ~n17863;
  assign n17865 = n3492 & ~n17864;
  assign n17866 = ~n17612 & ~n17865;
  assign n17867 = n3485 & ~n17866;
  assign n17868 = ~n17611 & ~n17867;
  assign n17869 = n3476 & ~n17868;
  assign n17870 = ~n17678 & ~n17869;
  assign n17871 = n3374 & ~n17870;
  assign n17872 = ~n17618 & ~n17871;
  assign n17873 = ~n3655 & ~n17872;
  assign n17874 = ~n17529 & ~n17873;
  assign n17875 = n3652 & ~n17874;
  assign n17876 = controllable_hmaster0 & ~n9440;
  assign n17877 = ~controllable_hmaster1 & ~n17876;
  assign n17878 = ~controllable_hmaster1 & ~n17877;
  assign n17879 = i_hbusreq3 & ~n17878;
  assign n17880 = controllable_hmaster0 & ~n9453;
  assign n17881 = ~controllable_hmaster1 & ~n17880;
  assign n17882 = ~controllable_hmaster1 & ~n17881;
  assign n17883 = ~i_hbusreq3 & ~n17882;
  assign n17884 = ~n17879 & ~n17883;
  assign n17885 = ~controllable_hmaster2 & ~n17884;
  assign n17886 = ~controllable_hmaster2 & ~n17885;
  assign n17887 = ~controllable_hgrant3 & ~n17886;
  assign n17888 = ~n17276 & ~n17887;
  assign n17889 = controllable_nhgrant0 & ~n17888;
  assign n17890 = ~n17300 & ~n17889;
  assign n17891 = ~n3281 & ~n17890;
  assign n17892 = ~n3281 & ~n17891;
  assign n17893 = n3378 & ~n17892;
  assign n17894 = ~n3530 & ~n17885;
  assign n17895 = ~controllable_hgrant3 & ~n17894;
  assign n17896 = ~n17306 & ~n17895;
  assign n17897 = controllable_nhgrant0 & ~n17896;
  assign n17898 = ~n17314 & ~n17897;
  assign n17899 = ~n3281 & ~n17898;
  assign n17900 = ~n3950 & ~n17899;
  assign n17901 = ~n3378 & ~n17900;
  assign n17902 = ~n17893 & ~n17901;
  assign n17903 = n3492 & ~n17902;
  assign n17904 = ~n3493 & ~n17903;
  assign n17905 = n3485 & ~n17904;
  assign n17906 = ~n3486 & ~n17905;
  assign n17907 = ~n3476 & ~n17906;
  assign n17908 = ~n4333 & ~n17367;
  assign n17909 = controllable_hmaster0 & ~n17908;
  assign n17910 = ~n17370 & ~n17909;
  assign n17911 = ~controllable_hmaster1 & ~n17910;
  assign n17912 = ~n17360 & ~n17911;
  assign n17913 = i_hbusreq3 & ~n17912;
  assign n17914 = ~n4340 & ~n17395;
  assign n17915 = controllable_hmaster0 & ~n17914;
  assign n17916 = ~n17398 & ~n17915;
  assign n17917 = ~controllable_hmaster1 & ~n17916;
  assign n17918 = ~n17375 & ~n17917;
  assign n17919 = ~i_hbusreq3 & ~n17918;
  assign n17920 = ~n17913 & ~n17919;
  assign n17921 = ~controllable_hmaster2 & ~n17920;
  assign n17922 = ~n17359 & ~n17921;
  assign n17923 = ~controllable_hgrant3 & ~n17922;
  assign n17924 = ~n17276 & ~n17923;
  assign n17925 = controllable_nhgrant0 & ~n17924;
  assign n17926 = ~n17300 & ~n17925;
  assign n17927 = ~n3281 & ~n17926;
  assign n17928 = ~n3281 & ~n17927;
  assign n17929 = n3378 & ~n17928;
  assign n17930 = ~n4333 & ~n17476;
  assign n17931 = controllable_hmaster0 & ~n17930;
  assign n17932 = ~n17423 & ~n17931;
  assign n17933 = ~controllable_hmaster1 & ~n17932;
  assign n17934 = ~n17474 & ~n17933;
  assign n17935 = i_hbusreq3 & ~n17934;
  assign n17936 = ~n4340 & ~n17503;
  assign n17937 = controllable_hmaster0 & ~n17936;
  assign n17938 = ~n17467 & ~n17937;
  assign n17939 = ~controllable_hmaster1 & ~n17938;
  assign n17940 = ~n17483 & ~n17939;
  assign n17941 = ~i_hbusreq3 & ~n17940;
  assign n17942 = ~n17935 & ~n17941;
  assign n17943 = ~controllable_hmaster2 & ~n17942;
  assign n17944 = ~n17473 & ~n17943;
  assign n17945 = ~controllable_hgrant3 & ~n17944;
  assign n17946 = ~n17306 & ~n17945;
  assign n17947 = controllable_nhgrant0 & ~n17946;
  assign n17948 = ~n17314 & ~n17947;
  assign n17949 = ~n3281 & ~n17948;
  assign n17950 = ~n4089 & ~n17949;
  assign n17951 = ~n3378 & ~n17950;
  assign n17952 = ~n17929 & ~n17951;
  assign n17953 = n3492 & ~n17952;
  assign n17954 = ~n3493 & ~n17953;
  assign n17955 = n3485 & ~n17954;
  assign n17956 = ~n3486 & ~n17955;
  assign n17957 = n3476 & ~n17956;
  assign n17958 = ~n17907 & ~n17957;
  assign n17959 = n3374 & ~n17958;
  assign n17960 = ~n17268 & ~n17959;
  assign n17961 = n3655 & ~n17960;
  assign n17962 = controllable_hmaster0 & ~n9594;
  assign n17963 = ~controllable_hmaster1 & ~n17962;
  assign n17964 = ~controllable_hmaster1 & ~n17963;
  assign n17965 = i_hbusreq3 & ~n17964;
  assign n17966 = controllable_hmaster0 & ~n9607;
  assign n17967 = ~controllable_hmaster1 & ~n17966;
  assign n17968 = ~controllable_hmaster1 & ~n17967;
  assign n17969 = ~i_hbusreq3 & ~n17968;
  assign n17970 = ~n17965 & ~n17969;
  assign n17971 = ~controllable_hmaster2 & ~n17970;
  assign n17972 = ~controllable_hmaster2 & ~n17971;
  assign n17973 = ~controllable_hgrant3 & ~n17972;
  assign n17974 = ~n17276 & ~n17973;
  assign n17975 = controllable_nhgrant0 & ~n17974;
  assign n17976 = ~n17300 & ~n17975;
  assign n17977 = ~n3281 & ~n17976;
  assign n17978 = ~n3281 & ~n17977;
  assign n17979 = n3378 & ~n17978;
  assign n17980 = ~n17664 & ~n17971;
  assign n17981 = ~controllable_hgrant3 & ~n17980;
  assign n17982 = ~n17306 & ~n17981;
  assign n17983 = controllable_nhgrant0 & ~n17982;
  assign n17984 = ~n17314 & ~n17983;
  assign n17985 = ~n3281 & ~n17984;
  assign n17986 = ~n3950 & ~n17985;
  assign n17987 = ~n3378 & ~n17986;
  assign n17988 = ~n17979 & ~n17987;
  assign n17989 = n3492 & ~n17988;
  assign n17990 = ~n3493 & ~n17989;
  assign n17991 = n3485 & ~n17990;
  assign n17992 = ~n3486 & ~n17991;
  assign n17993 = ~n3476 & ~n17992;
  assign n17994 = ~n4333 & ~n17714;
  assign n17995 = controllable_hmaster0 & ~n17994;
  assign n17996 = ~n17717 & ~n17995;
  assign n17997 = ~controllable_hmaster1 & ~n17996;
  assign n17998 = ~n17709 & ~n17997;
  assign n17999 = i_hbusreq3 & ~n17998;
  assign n18000 = ~n4340 & ~n17742;
  assign n18001 = controllable_hmaster0 & ~n18000;
  assign n18002 = ~n17745 & ~n18001;
  assign n18003 = ~controllable_hmaster1 & ~n18002;
  assign n18004 = ~n17722 & ~n18003;
  assign n18005 = ~i_hbusreq3 & ~n18004;
  assign n18006 = ~n17999 & ~n18005;
  assign n18007 = ~controllable_hmaster2 & ~n18006;
  assign n18008 = ~n17708 & ~n18007;
  assign n18009 = ~controllable_hgrant3 & ~n18008;
  assign n18010 = ~n17276 & ~n18009;
  assign n18011 = controllable_nhgrant0 & ~n18010;
  assign n18012 = ~n17300 & ~n18011;
  assign n18013 = ~n3281 & ~n18012;
  assign n18014 = ~n3281 & ~n18013;
  assign n18015 = n3378 & ~n18014;
  assign n18016 = ~n4333 & ~n17822;
  assign n18017 = controllable_hmaster0 & ~n18016;
  assign n18018 = ~n17770 & ~n18017;
  assign n18019 = ~controllable_hmaster1 & ~n18018;
  assign n18020 = ~n17820 & ~n18019;
  assign n18021 = i_hbusreq3 & ~n18020;
  assign n18022 = ~n4340 & ~n17847;
  assign n18023 = controllable_hmaster0 & ~n18022;
  assign n18024 = ~n17813 & ~n18023;
  assign n18025 = ~controllable_hmaster1 & ~n18024;
  assign n18026 = ~n17829 & ~n18025;
  assign n18027 = ~i_hbusreq3 & ~n18026;
  assign n18028 = ~n18021 & ~n18027;
  assign n18029 = ~controllable_hmaster2 & ~n18028;
  assign n18030 = ~n17819 & ~n18029;
  assign n18031 = ~controllable_hgrant3 & ~n18030;
  assign n18032 = ~n17306 & ~n18031;
  assign n18033 = controllable_nhgrant0 & ~n18032;
  assign n18034 = ~n17314 & ~n18033;
  assign n18035 = ~n3281 & ~n18034;
  assign n18036 = ~n4089 & ~n18035;
  assign n18037 = ~n3378 & ~n18036;
  assign n18038 = ~n18015 & ~n18037;
  assign n18039 = n3492 & ~n18038;
  assign n18040 = ~n17612 & ~n18039;
  assign n18041 = n3485 & ~n18040;
  assign n18042 = ~n17611 & ~n18041;
  assign n18043 = n3476 & ~n18042;
  assign n18044 = ~n17993 & ~n18043;
  assign n18045 = n3374 & ~n18044;
  assign n18046 = ~n17618 & ~n18045;
  assign n18047 = ~n3655 & ~n18046;
  assign n18048 = ~n17961 & ~n18047;
  assign n18049 = ~n3652 & ~n18048;
  assign n18050 = ~n17875 & ~n18049;
  assign n18051 = ~n3368 & ~n18050;
  assign n18052 = ~controllable_hmaster1 & ~n9702;
  assign n18053 = ~i_hbusreq3 & ~n18052;
  assign n18054 = ~n17270 & ~n18053;
  assign n18055 = ~controllable_hmaster2 & ~n18054;
  assign n18056 = ~controllable_hmaster2 & ~n18055;
  assign n18057 = controllable_hgrant3 & ~n18056;
  assign n18058 = controllable_hmaster0 & ~n9826;
  assign n18059 = ~controllable_hmaster1 & ~n18058;
  assign n18060 = ~controllable_hmaster1 & ~n18059;
  assign n18061 = ~i_hbusreq3 & ~n18060;
  assign n18062 = ~n17280 & ~n18061;
  assign n18063 = ~controllable_hmaster2 & ~n18062;
  assign n18064 = ~controllable_hmaster2 & ~n18063;
  assign n18065 = ~controllable_hgrant3 & ~n18064;
  assign n18066 = ~n18057 & ~n18065;
  assign n18067 = controllable_nhgrant0 & ~n18066;
  assign n18068 = ~controllable_hmaster1 & ~n9739;
  assign n18069 = i_hbusreq3 & ~n18068;
  assign n18070 = ~controllable_hmaster1 & ~n9745;
  assign n18071 = ~i_hbusreq3 & ~n18070;
  assign n18072 = ~n18069 & ~n18071;
  assign n18073 = ~controllable_hmaster2 & ~n18072;
  assign n18074 = ~controllable_hmaster2 & ~n18073;
  assign n18075 = ~controllable_hgrant3 & ~n18074;
  assign n18076 = ~n18057 & ~n18075;
  assign n18077 = ~controllable_nhgrant0 & ~n18076;
  assign n18078 = ~n18067 & ~n18077;
  assign n18079 = ~n3281 & ~n18078;
  assign n18080 = ~n3281 & ~n18079;
  assign n18081 = n3492 & ~n18080;
  assign n18082 = n3492 & ~n18081;
  assign n18083 = n3485 & ~n18082;
  assign n18084 = n3485 & ~n18083;
  assign n18085 = ~n3476 & ~n18084;
  assign n18086 = controllable_hmaster2 & ~n17333;
  assign n18087 = ~i_hbusreq1 & n17325;
  assign n18088 = ~n17379 & ~n18087;
  assign n18089 = ~controllable_ndecide & n18088;
  assign n18090 = ~controllable_ndecide & ~n18089;
  assign n18091 = i_hready & ~n18090;
  assign n18092 = ~n4577 & ~n18091;
  assign n18093 = i_hlock0 & ~n18092;
  assign n18094 = ~n17385 & ~n18093;
  assign n18095 = ~i_hbusreq0 & ~n18094;
  assign n18096 = ~n17378 & ~n18095;
  assign n18097 = ~i_hbusreq4 & ~n18096;
  assign n18098 = ~n17377 & ~n18097;
  assign n18099 = ~controllable_hgrant4 & ~n18098;
  assign n18100 = ~n4617 & ~n18099;
  assign n18101 = ~i_hbusreq2 & ~n18100;
  assign n18102 = ~n17376 & ~n18101;
  assign n18103 = ~controllable_hgrant2 & ~n18102;
  assign n18104 = ~n4562 & ~n18103;
  assign n18105 = controllable_hmaster0 & ~n18104;
  assign n18106 = ~n17370 & ~n18105;
  assign n18107 = ~controllable_hmaster1 & ~n18106;
  assign n18108 = ~n17360 & ~n18107;
  assign n18109 = ~i_hbusreq3 & ~n18108;
  assign n18110 = ~n17374 & ~n18109;
  assign n18111 = ~controllable_hmaster2 & ~n18110;
  assign n18112 = ~n18086 & ~n18111;
  assign n18113 = ~controllable_hgrant3 & ~n18112;
  assign n18114 = ~n18057 & ~n18113;
  assign n18115 = controllable_nhgrant0 & ~n18114;
  assign n18116 = ~n18077 & ~n18115;
  assign n18117 = ~n3281 & ~n18116;
  assign n18118 = ~n3281 & ~n18117;
  assign n18119 = n3492 & ~n18118;
  assign n18120 = n3492 & ~n18119;
  assign n18121 = n3485 & ~n18120;
  assign n18122 = n3485 & ~n18121;
  assign n18123 = n3476 & ~n18122;
  assign n18124 = ~n18085 & ~n18123;
  assign n18125 = n3374 & ~n18124;
  assign n18126 = n3374 & ~n18125;
  assign n18127 = n3655 & ~n18126;
  assign n18128 = controllable_hmaster0 & ~n10336;
  assign n18129 = ~controllable_hmaster1 & ~n18128;
  assign n18130 = ~controllable_hmaster1 & ~n18129;
  assign n18131 = i_hbusreq3 & ~n18130;
  assign n18132 = controllable_hmaster0 & ~n10376;
  assign n18133 = ~controllable_hmaster1 & ~n18132;
  assign n18134 = ~controllable_hmaster1 & ~n18133;
  assign n18135 = ~i_hbusreq3 & ~n18134;
  assign n18136 = ~n18131 & ~n18135;
  assign n18137 = ~controllable_hmaster2 & ~n18136;
  assign n18138 = ~controllable_hmaster2 & ~n18137;
  assign n18139 = ~controllable_hgrant3 & ~n18138;
  assign n18140 = ~n18057 & ~n18139;
  assign n18141 = controllable_nhgrant0 & ~n18140;
  assign n18142 = ~n18077 & ~n18141;
  assign n18143 = ~n3281 & ~n18142;
  assign n18144 = ~n3281 & ~n18143;
  assign n18145 = n3492 & ~n18144;
  assign n18146 = n3492 & ~n18145;
  assign n18147 = n3485 & ~n18146;
  assign n18148 = n3485 & ~n18147;
  assign n18149 = ~n3476 & ~n18148;
  assign n18150 = ~n3485 & ~n17546;
  assign n18151 = ~n3492 & ~n17546;
  assign n18152 = i_hlock1 & controllable_hgrant1;
  assign n18153 = ~i_hlock1 & n17325;
  assign n18154 = ~n18152 & ~n18153;
  assign n18155 = ~controllable_ndecide & ~n18154;
  assign n18156 = ~n3494 & ~n18155;
  assign n18157 = i_hready & ~n18156;
  assign n18158 = ~controllable_hgrant4 & ~n18157;
  assign n18159 = ~controllable_hgrant4 & ~n18158;
  assign n18160 = ~controllable_hgrant2 & ~n18159;
  assign n18161 = ~controllable_hgrant2 & ~n18160;
  assign n18162 = i_hbusreq3 & ~n18161;
  assign n18163 = i_hbusreq2 & ~n18159;
  assign n18164 = i_hbusreq4 & n18157;
  assign n18165 = i_hbusreq0 & n18157;
  assign n18166 = i_hbusreq1 & ~n18154;
  assign n18167 = ~n18087 & ~n18166;
  assign n18168 = ~controllable_ndecide & ~n18167;
  assign n18169 = ~n3494 & ~n18168;
  assign n18170 = i_hready & ~n18169;
  assign n18171 = ~i_hbusreq0 & n18170;
  assign n18172 = ~n18165 & ~n18171;
  assign n18173 = ~i_hbusreq4 & ~n18172;
  assign n18174 = ~n18164 & ~n18173;
  assign n18175 = ~controllable_hgrant4 & n18174;
  assign n18176 = ~controllable_hgrant4 & ~n18175;
  assign n18177 = ~i_hbusreq2 & ~n18176;
  assign n18178 = ~n18163 & ~n18177;
  assign n18179 = ~controllable_hgrant2 & ~n18178;
  assign n18180 = ~controllable_hgrant2 & ~n18179;
  assign n18181 = ~i_hbusreq3 & ~n18180;
  assign n18182 = ~n18162 & ~n18181;
  assign n18183 = controllable_hmaster2 & ~n18182;
  assign n18184 = controllable_hmaster1 & ~n18161;
  assign n18185 = ~i_hlock1 & n5691;
  assign n18186 = ~n18152 & ~n18185;
  assign n18187 = ~controllable_ndecide & ~n18186;
  assign n18188 = ~n3494 & ~n18187;
  assign n18189 = i_hready & ~n18188;
  assign n18190 = i_hready & ~n18189;
  assign n18191 = ~controllable_hgrant4 & n18190;
  assign n18192 = ~n3411 & ~n18191;
  assign n18193 = ~controllable_hgrant2 & ~n18192;
  assign n18194 = ~n3410 & ~n18193;
  assign n18195 = controllable_hmaster0 & ~n18194;
  assign n18196 = ~controllable_hmaster0 & ~n18161;
  assign n18197 = ~n18195 & ~n18196;
  assign n18198 = ~controllable_hmaster1 & ~n18197;
  assign n18199 = ~n18184 & ~n18198;
  assign n18200 = i_hbusreq3 & ~n18199;
  assign n18201 = controllable_hmaster1 & ~n18180;
  assign n18202 = i_hbusreq2 & ~n18192;
  assign n18203 = i_hbusreq4 & ~n18190;
  assign n18204 = i_hbusreq0 & ~n18190;
  assign n18205 = i_hbusreq1 & ~n18186;
  assign n18206 = ~n18087 & ~n18205;
  assign n18207 = ~controllable_ndecide & ~n18206;
  assign n18208 = ~n3494 & ~n18207;
  assign n18209 = i_hready & ~n18208;
  assign n18210 = ~n10361 & ~n18209;
  assign n18211 = i_hlock0 & ~n18210;
  assign n18212 = ~n17487 & ~n18205;
  assign n18213 = ~controllable_ndecide & ~n18212;
  assign n18214 = ~n3494 & ~n18213;
  assign n18215 = i_hready & ~n18214;
  assign n18216 = i_hready & ~n18215;
  assign n18217 = ~i_hlock0 & ~n18216;
  assign n18218 = ~n18211 & ~n18217;
  assign n18219 = ~i_hbusreq0 & ~n18218;
  assign n18220 = ~n18204 & ~n18219;
  assign n18221 = ~i_hbusreq4 & ~n18220;
  assign n18222 = ~n18203 & ~n18221;
  assign n18223 = ~controllable_hgrant4 & n18222;
  assign n18224 = ~n4617 & ~n18223;
  assign n18225 = ~i_hbusreq2 & ~n18224;
  assign n18226 = ~n18202 & ~n18225;
  assign n18227 = ~controllable_hgrant2 & ~n18226;
  assign n18228 = ~n4562 & ~n18227;
  assign n18229 = controllable_hmaster0 & ~n18228;
  assign n18230 = ~controllable_hmaster0 & ~n18180;
  assign n18231 = ~n18229 & ~n18230;
  assign n18232 = ~controllable_hmaster1 & ~n18231;
  assign n18233 = ~n18201 & ~n18232;
  assign n18234 = ~i_hbusreq3 & ~n18233;
  assign n18235 = ~n18200 & ~n18234;
  assign n18236 = ~controllable_hmaster2 & ~n18235;
  assign n18237 = ~n18183 & ~n18236;
  assign n18238 = ~controllable_hgrant3 & ~n18237;
  assign n18239 = ~n18057 & ~n18238;
  assign n18240 = controllable_nhgrant0 & ~n18239;
  assign n18241 = ~n18077 & ~n18240;
  assign n18242 = ~n3281 & ~n18241;
  assign n18243 = ~n3281 & ~n18242;
  assign n18244 = n3492 & ~n18243;
  assign n18245 = ~n18151 & ~n18244;
  assign n18246 = n3485 & ~n18245;
  assign n18247 = ~n18150 & ~n18246;
  assign n18248 = n3476 & ~n18247;
  assign n18249 = ~n18149 & ~n18248;
  assign n18250 = n3374 & ~n18249;
  assign n18251 = n3374 & ~n18250;
  assign n18252 = ~n3655 & ~n18251;
  assign n18253 = ~n18127 & ~n18252;
  assign n18254 = n3652 & ~n18253;
  assign n18255 = controllable_hmaster0 & ~n10774;
  assign n18256 = ~controllable_hmaster1 & ~n18255;
  assign n18257 = ~controllable_hmaster1 & ~n18256;
  assign n18258 = i_hbusreq3 & ~n18257;
  assign n18259 = controllable_hmaster0 & ~n10788;
  assign n18260 = ~controllable_hmaster1 & ~n18259;
  assign n18261 = ~controllable_hmaster1 & ~n18260;
  assign n18262 = ~i_hbusreq3 & ~n18261;
  assign n18263 = ~n18258 & ~n18262;
  assign n18264 = ~controllable_hmaster2 & ~n18263;
  assign n18265 = ~controllable_hmaster2 & ~n18264;
  assign n18266 = ~controllable_hgrant3 & ~n18265;
  assign n18267 = ~n18057 & ~n18266;
  assign n18268 = controllable_nhgrant0 & ~n18267;
  assign n18269 = ~n18077 & ~n18268;
  assign n18270 = ~n3281 & ~n18269;
  assign n18271 = ~n3281 & ~n18270;
  assign n18272 = n3492 & ~n18271;
  assign n18273 = n3492 & ~n18272;
  assign n18274 = n3485 & ~n18273;
  assign n18275 = n3485 & ~n18274;
  assign n18276 = ~n3476 & ~n18275;
  assign n18277 = ~n4787 & ~n17367;
  assign n18278 = controllable_hmaster0 & ~n18277;
  assign n18279 = ~n17370 & ~n18278;
  assign n18280 = ~controllable_hmaster1 & ~n18279;
  assign n18281 = ~n17360 & ~n18280;
  assign n18282 = i_hbusreq3 & ~n18281;
  assign n18283 = ~n4794 & ~n18103;
  assign n18284 = controllable_hmaster0 & ~n18283;
  assign n18285 = ~n17370 & ~n18284;
  assign n18286 = ~controllable_hmaster1 & ~n18285;
  assign n18287 = ~n17360 & ~n18286;
  assign n18288 = ~i_hbusreq3 & ~n18287;
  assign n18289 = ~n18282 & ~n18288;
  assign n18290 = ~controllable_hmaster2 & ~n18289;
  assign n18291 = ~n18086 & ~n18290;
  assign n18292 = ~controllable_hgrant3 & ~n18291;
  assign n18293 = ~n18057 & ~n18292;
  assign n18294 = controllable_nhgrant0 & ~n18293;
  assign n18295 = ~n18077 & ~n18294;
  assign n18296 = ~n3281 & ~n18295;
  assign n18297 = ~n3281 & ~n18296;
  assign n18298 = n3492 & ~n18297;
  assign n18299 = n3492 & ~n18298;
  assign n18300 = n3485 & ~n18299;
  assign n18301 = n3485 & ~n18300;
  assign n18302 = n3476 & ~n18301;
  assign n18303 = ~n18276 & ~n18302;
  assign n18304 = n3374 & ~n18303;
  assign n18305 = n3374 & ~n18304;
  assign n18306 = n3655 & ~n18305;
  assign n18307 = controllable_hmaster0 & ~n11209;
  assign n18308 = ~controllable_hmaster1 & ~n18307;
  assign n18309 = ~controllable_hmaster1 & ~n18308;
  assign n18310 = i_hbusreq3 & ~n18309;
  assign n18311 = controllable_hmaster0 & ~n11222;
  assign n18312 = ~controllable_hmaster1 & ~n18311;
  assign n18313 = ~controllable_hmaster1 & ~n18312;
  assign n18314 = ~i_hbusreq3 & ~n18313;
  assign n18315 = ~n18310 & ~n18314;
  assign n18316 = ~controllable_hmaster2 & ~n18315;
  assign n18317 = ~controllable_hmaster2 & ~n18316;
  assign n18318 = ~controllable_hgrant3 & ~n18317;
  assign n18319 = ~n18057 & ~n18318;
  assign n18320 = controllable_nhgrant0 & ~n18319;
  assign n18321 = ~n18077 & ~n18320;
  assign n18322 = ~n3281 & ~n18321;
  assign n18323 = ~n3281 & ~n18322;
  assign n18324 = n3492 & ~n18323;
  assign n18325 = n3492 & ~n18324;
  assign n18326 = n3485 & ~n18325;
  assign n18327 = n3485 & ~n18326;
  assign n18328 = ~n3476 & ~n18327;
  assign n18329 = ~n4787 & ~n18193;
  assign n18330 = controllable_hmaster0 & ~n18329;
  assign n18331 = ~n18196 & ~n18330;
  assign n18332 = ~controllable_hmaster1 & ~n18331;
  assign n18333 = ~n18184 & ~n18332;
  assign n18334 = i_hbusreq3 & ~n18333;
  assign n18335 = ~n4794 & ~n18227;
  assign n18336 = controllable_hmaster0 & ~n18335;
  assign n18337 = ~n18230 & ~n18336;
  assign n18338 = ~controllable_hmaster1 & ~n18337;
  assign n18339 = ~n18201 & ~n18338;
  assign n18340 = ~i_hbusreq3 & ~n18339;
  assign n18341 = ~n18334 & ~n18340;
  assign n18342 = ~controllable_hmaster2 & ~n18341;
  assign n18343 = ~n18183 & ~n18342;
  assign n18344 = ~controllable_hgrant3 & ~n18343;
  assign n18345 = ~n18057 & ~n18344;
  assign n18346 = controllable_nhgrant0 & ~n18345;
  assign n18347 = ~n18077 & ~n18346;
  assign n18348 = ~n3281 & ~n18347;
  assign n18349 = ~n3281 & ~n18348;
  assign n18350 = n3492 & ~n18349;
  assign n18351 = ~n18151 & ~n18350;
  assign n18352 = n3485 & ~n18351;
  assign n18353 = ~n18150 & ~n18352;
  assign n18354 = n3476 & ~n18353;
  assign n18355 = ~n18328 & ~n18354;
  assign n18356 = n3374 & ~n18355;
  assign n18357 = n3374 & ~n18356;
  assign n18358 = ~n3655 & ~n18357;
  assign n18359 = ~n18306 & ~n18358;
  assign n18360 = ~n3652 & ~n18359;
  assign n18361 = ~n18254 & ~n18360;
  assign n18362 = n3368 & ~n18361;
  assign n18363 = ~n18051 & ~n18362;
  assign n18364 = ~n3362 & ~n18363;
  assign n18365 = ~n3362 & ~n18364;
  assign n18366 = ~n3359 & ~n18365;
  assign n18367 = ~n3359 & ~n18366;
  assign n18368 = n3356 & ~n18367;
  assign n18369 = n3378 & ~n17261;
  assign n18370 = ~n5249 & ~n18369;
  assign n18371 = n3492 & ~n18370;
  assign n18372 = ~n3631 & ~n18371;
  assign n18373 = n3485 & ~n18372;
  assign n18374 = ~n3630 & ~n18373;
  assign n18375 = ~n3374 & ~n18374;
  assign n18376 = ~controllable_hmaster1 & ~n12080;
  assign n18377 = ~n5280 & ~n18376;
  assign n18378 = ~i_hbusreq3 & ~n18377;
  assign n18379 = ~n5265 & ~n18378;
  assign n18380 = ~controllable_hmaster2 & ~n18379;
  assign n18381 = ~n12033 & ~n18380;
  assign n18382 = controllable_hgrant3 & ~n18381;
  assign n18383 = ~n3821 & ~n8826;
  assign n18384 = ~controllable_hmaster1 & ~n18383;
  assign n18385 = ~n5293 & ~n18384;
  assign n18386 = i_hbusreq3 & ~n18385;
  assign n18387 = ~n5278 & ~n8860;
  assign n18388 = ~controllable_hmaster1 & ~n18387;
  assign n18389 = ~n5313 & ~n18388;
  assign n18390 = ~i_hbusreq3 & ~n18389;
  assign n18391 = ~n18386 & ~n18390;
  assign n18392 = ~controllable_hmaster2 & ~n18391;
  assign n18393 = ~n12065 & ~n18392;
  assign n18394 = ~controllable_hgrant3 & ~n18393;
  assign n18395 = ~n18382 & ~n18394;
  assign n18396 = controllable_nhgrant0 & ~n18395;
  assign n18397 = ~n3400 & ~n18376;
  assign n18398 = ~i_hbusreq3 & ~n18397;
  assign n18399 = ~n3951 & ~n18398;
  assign n18400 = ~controllable_hmaster2 & ~n18399;
  assign n18401 = ~n12033 & ~n18400;
  assign n18402 = controllable_hgrant3 & ~n18401;
  assign n18403 = ~n5191 & ~n5348;
  assign n18404 = ~controllable_hmaster1 & ~n18403;
  assign n18405 = ~n3381 & ~n18404;
  assign n18406 = i_hbusreq3 & ~n18405;
  assign n18407 = ~n5197 & ~n5353;
  assign n18408 = ~controllable_hmaster1 & ~n18407;
  assign n18409 = ~n3400 & ~n18408;
  assign n18410 = ~i_hbusreq3 & ~n18409;
  assign n18411 = ~n18406 & ~n18410;
  assign n18412 = ~controllable_hmaster2 & ~n18411;
  assign n18413 = ~n12033 & ~n18412;
  assign n18414 = ~controllable_hgrant3 & ~n18413;
  assign n18415 = ~n18402 & ~n18414;
  assign n18416 = ~controllable_nhgrant0 & ~n18415;
  assign n18417 = ~n18396 & ~n18416;
  assign n18418 = ~n3281 & ~n18417;
  assign n18419 = ~n3950 & ~n18418;
  assign n18420 = n3378 & ~n18419;
  assign n18421 = ~n3910 & ~n8826;
  assign n18422 = ~controllable_hmaster1 & ~n18421;
  assign n18423 = ~n5427 & ~n18422;
  assign n18424 = i_hbusreq3 & ~n18423;
  assign n18425 = ~n5478 & ~n8860;
  assign n18426 = ~controllable_hmaster1 & ~n18425;
  assign n18427 = ~n5442 & ~n18426;
  assign n18428 = ~i_hbusreq3 & ~n18427;
  assign n18429 = ~n18424 & ~n18428;
  assign n18430 = ~controllable_hmaster2 & ~n18429;
  assign n18431 = ~n12126 & ~n18430;
  assign n18432 = ~controllable_hgrant3 & ~n18431;
  assign n18433 = ~n5402 & ~n18432;
  assign n18434 = controllable_nhgrant0 & ~n18433;
  assign n18435 = ~n5534 & ~n18434;
  assign n18436 = ~n3281 & ~n18435;
  assign n18437 = ~n3950 & ~n18436;
  assign n18438 = ~n3378 & ~n18437;
  assign n18439 = ~n18420 & ~n18438;
  assign n18440 = n3492 & ~n18439;
  assign n18441 = ~n3631 & ~n18440;
  assign n18442 = n3485 & ~n18441;
  assign n18443 = ~n3630 & ~n18442;
  assign n18444 = ~n3476 & ~n18443;
  assign n18445 = controllable_hmaster0 & ~n5575;
  assign n18446 = ~n5606 & ~n18445;
  assign n18447 = ~controllable_hmaster1 & ~n18446;
  assign n18448 = ~n5608 & ~n18447;
  assign n18449 = ~i_hbusreq3 & ~n18448;
  assign n18450 = ~n5593 & ~n18449;
  assign n18451 = ~controllable_hmaster2 & ~n18450;
  assign n18452 = ~n12233 & ~n18451;
  assign n18453 = controllable_hgrant3 & ~n18452;
  assign n18454 = ~n12172 & ~n17441;
  assign n18455 = ~i_hbusreq2 & ~n18454;
  assign n18456 = ~n5636 & ~n18455;
  assign n18457 = ~controllable_hgrant2 & ~n18456;
  assign n18458 = ~n5635 & ~n18457;
  assign n18459 = controllable_hmaster1 & ~n18458;
  assign n18460 = controllable_hmaster0 & ~n18458;
  assign n18461 = i_hlock0 & ~n5710;
  assign n18462 = ~n3392 & ~n17433;
  assign n18463 = ~i_hlock0 & ~n18462;
  assign n18464 = ~n18461 & ~n18463;
  assign n18465 = ~i_hbusreq0 & ~n18464;
  assign n18466 = ~n5709 & ~n18465;
  assign n18467 = ~i_hbusreq4 & ~n18466;
  assign n18468 = ~n5708 & ~n18467;
  assign n18469 = ~controllable_hgrant4 & ~n18468;
  assign n18470 = ~n12181 & ~n18469;
  assign n18471 = ~i_hbusreq2 & ~n18470;
  assign n18472 = ~n12180 & ~n18471;
  assign n18473 = ~controllable_hgrant2 & ~n18472;
  assign n18474 = ~n5635 & ~n18473;
  assign n18475 = ~controllable_hmaster0 & ~n18474;
  assign n18476 = ~n18460 & ~n18475;
  assign n18477 = ~controllable_hmaster1 & ~n18476;
  assign n18478 = ~n18459 & ~n18477;
  assign n18479 = ~i_hbusreq3 & ~n18478;
  assign n18480 = ~n12171 & ~n18479;
  assign n18481 = controllable_hmaster2 & ~n18480;
  assign n18482 = ~n5702 & ~n8991;
  assign n18483 = ~controllable_hmaster1 & ~n18482;
  assign n18484 = ~n5690 & ~n18483;
  assign n18485 = i_hbusreq3 & ~n18484;
  assign n18486 = ~n12172 & ~n18469;
  assign n18487 = ~i_hbusreq2 & ~n18486;
  assign n18488 = ~n5707 & ~n18487;
  assign n18489 = ~controllable_hgrant2 & ~n18488;
  assign n18490 = ~n5635 & ~n18489;
  assign n18491 = controllable_hmaster0 & ~n18490;
  assign n18492 = ~n5722 & ~n18489;
  assign n18493 = ~controllable_hmaster0 & ~n18492;
  assign n18494 = ~n18491 & ~n18493;
  assign n18495 = controllable_hmaster1 & ~n18494;
  assign n18496 = ~n12198 & ~n17499;
  assign n18497 = ~i_hbusreq2 & ~n18496;
  assign n18498 = ~n9007 & ~n18497;
  assign n18499 = ~controllable_hgrant2 & ~n18498;
  assign n18500 = ~n5657 & ~n18499;
  assign n18501 = controllable_hmaster0 & ~n18500;
  assign n18502 = ~controllable_hmaster0 & ~n18490;
  assign n18503 = ~n18501 & ~n18502;
  assign n18504 = ~controllable_hmaster1 & ~n18503;
  assign n18505 = ~n18495 & ~n18504;
  assign n18506 = ~i_hbusreq3 & ~n18505;
  assign n18507 = ~n18485 & ~n18506;
  assign n18508 = ~controllable_hmaster2 & ~n18507;
  assign n18509 = ~n18481 & ~n18508;
  assign n18510 = ~controllable_hgrant3 & ~n18509;
  assign n18511 = ~n18453 & ~n18510;
  assign n18512 = controllable_nhgrant0 & ~n18511;
  assign n18513 = ~n5794 & ~n12234;
  assign n18514 = ~controllable_hmaster1 & ~n18513;
  assign n18515 = ~n5757 & ~n18514;
  assign n18516 = i_hbusreq3 & ~n18515;
  assign n18517 = ~n5799 & ~n12239;
  assign n18518 = ~controllable_hmaster1 & ~n18517;
  assign n18519 = ~n5561 & ~n18518;
  assign n18520 = ~i_hbusreq3 & ~n18519;
  assign n18521 = ~n18516 & ~n18520;
  assign n18522 = ~controllable_hmaster2 & ~n18521;
  assign n18523 = ~n12233 & ~n18522;
  assign n18524 = ~controllable_hgrant3 & ~n18523;
  assign n18525 = ~n18402 & ~n18524;
  assign n18526 = ~controllable_nhgrant0 & ~n18525;
  assign n18527 = ~n18512 & ~n18526;
  assign n18528 = ~n3281 & ~n18527;
  assign n18529 = ~n4089 & ~n18528;
  assign n18530 = n3378 & ~n18529;
  assign n18531 = ~n5926 & ~n8991;
  assign n18532 = ~controllable_hmaster1 & ~n18531;
  assign n18533 = ~n5919 & ~n18532;
  assign n18534 = i_hbusreq3 & ~n18533;
  assign n18535 = ~n9018 & ~n17486;
  assign n18536 = ~i_hbusreq0 & ~n18535;
  assign n18537 = ~n9009 & ~n18536;
  assign n18538 = ~i_hbusreq4 & ~n18537;
  assign n18539 = ~n9008 & ~n18538;
  assign n18540 = ~controllable_hgrant4 & ~n18539;
  assign n18541 = ~n5863 & ~n18540;
  assign n18542 = ~i_hbusreq2 & ~n18541;
  assign n18543 = ~n9007 & ~n18542;
  assign n18544 = ~controllable_hgrant2 & ~n18543;
  assign n18545 = ~n5862 & ~n18544;
  assign n18546 = controllable_hmaster0 & ~n18545;
  assign n18547 = ~n5996 & ~n18546;
  assign n18548 = ~controllable_hmaster1 & ~n18547;
  assign n18549 = ~n5954 & ~n18548;
  assign n18550 = ~i_hbusreq3 & ~n18549;
  assign n18551 = ~n18534 & ~n18550;
  assign n18552 = ~controllable_hmaster2 & ~n18551;
  assign n18553 = ~n12274 & ~n18552;
  assign n18554 = ~controllable_hgrant3 & ~n18553;
  assign n18555 = ~n5861 & ~n18554;
  assign n18556 = controllable_nhgrant0 & ~n18555;
  assign n18557 = ~n6082 & ~n18556;
  assign n18558 = ~n3281 & ~n18557;
  assign n18559 = ~n4089 & ~n18558;
  assign n18560 = ~n3378 & ~n18559;
  assign n18561 = ~n18530 & ~n18560;
  assign n18562 = n3492 & ~n18561;
  assign n18563 = ~n3631 & ~n18562;
  assign n18564 = n3485 & ~n18563;
  assign n18565 = ~n3630 & ~n18564;
  assign n18566 = n3476 & ~n18565;
  assign n18567 = ~n18444 & ~n18566;
  assign n18568 = n3374 & ~n18567;
  assign n18569 = ~n18375 & ~n18568;
  assign n18570 = n3655 & ~n18569;
  assign n18571 = n3378 & ~n17594;
  assign n18572 = ~controllable_hgrant1 & ~n4008;
  assign n18573 = ~controllable_hgrant1 & ~n18572;
  assign n18574 = controllable_ndecide & ~n18573;
  assign n18575 = controllable_ndecide & ~n18574;
  assign n18576 = ~i_hready & n18575;
  assign n18577 = ~n3417 & ~n18576;
  assign n18578 = ~controllable_hgrant4 & ~n18577;
  assign n18579 = ~n3411 & ~n18578;
  assign n18580 = ~controllable_hgrant2 & ~n18579;
  assign n18581 = ~n3410 & ~n18580;
  assign n18582 = controllable_hmaster1 & ~n18581;
  assign n18583 = controllable_hmaster0 & ~n18581;
  assign n18584 = ~n3729 & ~n18583;
  assign n18585 = ~controllable_hmaster1 & ~n18584;
  assign n18586 = ~n18582 & ~n18585;
  assign n18587 = i_hbusreq3 & ~n18586;
  assign n18588 = i_hbusreq2 & ~n18579;
  assign n18589 = i_hbusreq4 & ~n18577;
  assign n18590 = i_hbusreq0 & ~n18577;
  assign n18591 = ~n6304 & ~n18574;
  assign n18592 = ~i_hready & n18591;
  assign n18593 = ~n3440 & ~n18592;
  assign n18594 = i_hlock0 & ~n18593;
  assign n18595 = ~i_hlock0 & ~n18577;
  assign n18596 = ~n18594 & ~n18595;
  assign n18597 = ~i_hbusreq0 & ~n18596;
  assign n18598 = ~n18590 & ~n18597;
  assign n18599 = ~i_hbusreq4 & ~n18598;
  assign n18600 = ~n18589 & ~n18599;
  assign n18601 = ~controllable_hgrant4 & ~n18600;
  assign n18602 = ~n3916 & ~n18601;
  assign n18603 = ~i_hbusreq2 & ~n18602;
  assign n18604 = ~n18588 & ~n18603;
  assign n18605 = ~controllable_hgrant2 & ~n18604;
  assign n18606 = ~n3859 & ~n18605;
  assign n18607 = controllable_hmaster1 & ~n18606;
  assign n18608 = controllable_hmaster0 & ~n18606;
  assign n18609 = ~n3767 & ~n18608;
  assign n18610 = ~controllable_hmaster1 & ~n18609;
  assign n18611 = ~n18607 & ~n18610;
  assign n18612 = ~i_hbusreq3 & ~n18611;
  assign n18613 = ~n18587 & ~n18612;
  assign n18614 = controllable_hmaster2 & ~n18613;
  assign n18615 = ~n6188 & ~n18614;
  assign n18616 = ~controllable_hgrant3 & ~n18615;
  assign n18617 = ~n5037 & ~n18616;
  assign n18618 = controllable_nhgrant0 & ~n18617;
  assign n18619 = ~n5245 & ~n18618;
  assign n18620 = ~n3281 & ~n18619;
  assign n18621 = ~n3783 & ~n18620;
  assign n18622 = ~n3378 & ~n18621;
  assign n18623 = ~n18571 & ~n18622;
  assign n18624 = n3492 & ~n18623;
  assign n18625 = ~n3631 & ~n18624;
  assign n18626 = n3485 & ~n18625;
  assign n18627 = ~n3630 & ~n18626;
  assign n18628 = ~n3476 & ~n18627;
  assign n18629 = ~n3485 & ~n17608;
  assign n18630 = ~n3492 & ~n17608;
  assign n18631 = ~n18624 & ~n18630;
  assign n18632 = n3485 & ~n18631;
  assign n18633 = ~n18629 & ~n18632;
  assign n18634 = n3476 & ~n18633;
  assign n18635 = ~n18628 & ~n18634;
  assign n18636 = ~n3374 & ~n18635;
  assign n18637 = ~i_hready & n17689;
  assign n18638 = ~i_hready & ~n18637;
  assign n18639 = ~controllable_hgrant4 & ~n18638;
  assign n18640 = ~n3848 & ~n18639;
  assign n18641 = ~controllable_hgrant2 & ~n18640;
  assign n18642 = ~n3410 & ~n18641;
  assign n18643 = ~controllable_hmaster0 & ~n18642;
  assign n18644 = ~n9117 & ~n18643;
  assign n18645 = ~controllable_hmaster1 & ~n18644;
  assign n18646 = ~n9116 & ~n18645;
  assign n18647 = i_hbusreq3 & ~n18646;
  assign n18648 = i_hbusreq2 & ~n18640;
  assign n18649 = i_hbusreq4 & ~n18638;
  assign n18650 = i_hbusreq0 & ~n18638;
  assign n18651 = ~n3390 & ~n17689;
  assign n18652 = ~i_hready & ~n18651;
  assign n18653 = ~i_hready & ~n18652;
  assign n18654 = ~i_hbusreq0 & ~n18653;
  assign n18655 = ~n18650 & ~n18654;
  assign n18656 = ~i_hbusreq4 & ~n18655;
  assign n18657 = ~n18649 & ~n18656;
  assign n18658 = ~controllable_hgrant4 & ~n18657;
  assign n18659 = ~n12052 & ~n18658;
  assign n18660 = ~i_hbusreq2 & ~n18659;
  assign n18661 = ~n18648 & ~n18660;
  assign n18662 = ~controllable_hgrant2 & ~n18661;
  assign n18663 = ~n3431 & ~n18662;
  assign n18664 = ~controllable_hmaster0 & ~n18663;
  assign n18665 = ~n17658 & ~n18664;
  assign n18666 = ~controllable_hmaster1 & ~n18665;
  assign n18667 = ~n17657 & ~n18666;
  assign n18668 = ~i_hbusreq3 & ~n18667;
  assign n18669 = ~n18647 & ~n18668;
  assign n18670 = controllable_hmaster2 & ~n18669;
  assign n18671 = ~n3411 & ~n18639;
  assign n18672 = ~controllable_hgrant2 & ~n18671;
  assign n18673 = ~n3410 & ~n18672;
  assign n18674 = controllable_hmaster0 & ~n18673;
  assign n18675 = ~n5288 & ~n18672;
  assign n18676 = ~controllable_hmaster0 & ~n18675;
  assign n18677 = ~n18674 & ~n18676;
  assign n18678 = controllable_hmaster1 & ~n18677;
  assign n18679 = ~controllable_hmaster0 & ~n18673;
  assign n18680 = ~n9174 & ~n18679;
  assign n18681 = ~controllable_hmaster1 & ~n18680;
  assign n18682 = ~n18678 & ~n18681;
  assign n18683 = i_hbusreq3 & ~n18682;
  assign n18684 = i_hbusreq2 & ~n18671;
  assign n18685 = ~n3433 & ~n18658;
  assign n18686 = ~i_hbusreq2 & ~n18685;
  assign n18687 = ~n18684 & ~n18686;
  assign n18688 = ~controllable_hgrant2 & ~n18687;
  assign n18689 = ~n3431 & ~n18688;
  assign n18690 = controllable_hmaster0 & ~n18689;
  assign n18691 = ~n5308 & ~n18688;
  assign n18692 = ~controllable_hmaster0 & ~n18691;
  assign n18693 = ~n18690 & ~n18692;
  assign n18694 = controllable_hmaster1 & ~n18693;
  assign n18695 = ~controllable_hmaster0 & ~n18689;
  assign n18696 = ~n9210 & ~n18695;
  assign n18697 = ~controllable_hmaster1 & ~n18696;
  assign n18698 = ~n18694 & ~n18697;
  assign n18699 = ~i_hbusreq3 & ~n18698;
  assign n18700 = ~n18683 & ~n18699;
  assign n18701 = ~controllable_hmaster2 & ~n18700;
  assign n18702 = ~n18670 & ~n18701;
  assign n18703 = ~controllable_hgrant3 & ~n18702;
  assign n18704 = ~n18382 & ~n18703;
  assign n18705 = controllable_nhgrant0 & ~n18704;
  assign n18706 = ~n18416 & ~n18705;
  assign n18707 = ~n3281 & ~n18706;
  assign n18708 = ~n3950 & ~n18707;
  assign n18709 = n3378 & ~n18708;
  assign n18710 = ~n9117 & ~n12336;
  assign n18711 = ~controllable_hmaster1 & ~n18710;
  assign n18712 = ~n9116 & ~n18711;
  assign n18713 = i_hbusreq3 & ~n18712;
  assign n18714 = i_hlock0 & ~n17646;
  assign n18715 = ~i_hlock0 & n3417;
  assign n18716 = ~n18714 & ~n18715;
  assign n18717 = ~i_hbusreq0 & ~n18716;
  assign n18718 = ~n17643 & ~n18717;
  assign n18719 = ~i_hbusreq4 & ~n18718;
  assign n18720 = ~n17642 & ~n18719;
  assign n18721 = ~controllable_hgrant4 & ~n18720;
  assign n18722 = ~n3916 & ~n18721;
  assign n18723 = ~i_hbusreq2 & ~n18722;
  assign n18724 = ~n17641 & ~n18723;
  assign n18725 = ~controllable_hgrant2 & ~n18724;
  assign n18726 = ~n3859 & ~n18725;
  assign n18727 = controllable_hmaster1 & ~n18726;
  assign n18728 = controllable_hmaster0 & ~n18726;
  assign n18729 = ~n12347 & ~n18728;
  assign n18730 = ~controllable_hmaster1 & ~n18729;
  assign n18731 = ~n18727 & ~n18730;
  assign n18732 = ~i_hbusreq3 & ~n18731;
  assign n18733 = ~n18713 & ~n18732;
  assign n18734 = controllable_hmaster2 & ~n18733;
  assign n18735 = ~n6269 & ~n9174;
  assign n18736 = ~controllable_hmaster1 & ~n18735;
  assign n18737 = ~n6258 & ~n18736;
  assign n18738 = i_hbusreq3 & ~n18737;
  assign n18739 = ~n6337 & ~n9210;
  assign n18740 = ~controllable_hmaster1 & ~n18739;
  assign n18741 = ~n6297 & ~n18740;
  assign n18742 = ~i_hbusreq3 & ~n18741;
  assign n18743 = ~n18738 & ~n18742;
  assign n18744 = ~controllable_hmaster2 & ~n18743;
  assign n18745 = ~n18734 & ~n18744;
  assign n18746 = ~controllable_hgrant3 & ~n18745;
  assign n18747 = ~n5402 & ~n18746;
  assign n18748 = controllable_nhgrant0 & ~n18747;
  assign n18749 = ~n5534 & ~n18748;
  assign n18750 = ~n3281 & ~n18749;
  assign n18751 = ~n3950 & ~n18750;
  assign n18752 = ~n3378 & ~n18751;
  assign n18753 = ~n18709 & ~n18752;
  assign n18754 = n3492 & ~n18753;
  assign n18755 = ~n3631 & ~n18754;
  assign n18756 = n3485 & ~n18755;
  assign n18757 = ~n3630 & ~n18756;
  assign n18758 = ~n3476 & ~n18757;
  assign n18759 = ~n6401 & ~n18637;
  assign n18760 = ~controllable_hgrant4 & ~n18759;
  assign n18761 = ~n4015 & ~n18760;
  assign n18762 = ~controllable_hgrant2 & ~n18761;
  assign n18763 = ~n5616 & ~n18762;
  assign n18764 = ~controllable_hmaster0 & ~n18763;
  assign n18765 = ~n9253 & ~n18764;
  assign n18766 = ~controllable_hmaster1 & ~n18765;
  assign n18767 = ~n9252 & ~n18766;
  assign n18768 = i_hbusreq3 & ~n18767;
  assign n18769 = ~n12172 & ~n17787;
  assign n18770 = ~i_hbusreq2 & ~n18769;
  assign n18771 = ~n9258 & ~n18770;
  assign n18772 = ~controllable_hgrant2 & ~n18771;
  assign n18773 = ~n5635 & ~n18772;
  assign n18774 = controllable_hmaster1 & ~n18773;
  assign n18775 = controllable_hmaster0 & ~n18773;
  assign n18776 = i_hbusreq2 & ~n18761;
  assign n18777 = i_hbusreq4 & ~n18759;
  assign n18778 = i_hbusreq0 & ~n18759;
  assign n18779 = ~n6421 & ~n18652;
  assign n18780 = i_hlock0 & ~n18779;
  assign n18781 = ~n17779 & ~n18652;
  assign n18782 = ~i_hlock0 & ~n18781;
  assign n18783 = ~n18780 & ~n18782;
  assign n18784 = ~i_hbusreq0 & ~n18783;
  assign n18785 = ~n18778 & ~n18784;
  assign n18786 = ~i_hbusreq4 & ~n18785;
  assign n18787 = ~n18777 & ~n18786;
  assign n18788 = ~controllable_hgrant4 & ~n18787;
  assign n18789 = ~n12181 & ~n18788;
  assign n18790 = ~i_hbusreq2 & ~n18789;
  assign n18791 = ~n18776 & ~n18790;
  assign n18792 = ~controllable_hgrant2 & ~n18791;
  assign n18793 = ~n5635 & ~n18792;
  assign n18794 = ~controllable_hmaster0 & ~n18793;
  assign n18795 = ~n18775 & ~n18794;
  assign n18796 = ~controllable_hmaster1 & ~n18795;
  assign n18797 = ~n18774 & ~n18796;
  assign n18798 = ~i_hbusreq3 & ~n18797;
  assign n18799 = ~n18768 & ~n18798;
  assign n18800 = controllable_hmaster2 & ~n18799;
  assign n18801 = ~n4091 & ~n18760;
  assign n18802 = ~controllable_hgrant2 & ~n18801;
  assign n18803 = ~n5616 & ~n18802;
  assign n18804 = controllable_hmaster0 & ~n18803;
  assign n18805 = ~n5686 & ~n18802;
  assign n18806 = ~controllable_hmaster0 & ~n18805;
  assign n18807 = ~n18804 & ~n18806;
  assign n18808 = controllable_hmaster1 & ~n18807;
  assign n18809 = ~controllable_hmaster0 & ~n18803;
  assign n18810 = ~n9309 & ~n18809;
  assign n18811 = ~controllable_hmaster1 & ~n18810;
  assign n18812 = ~n18808 & ~n18811;
  assign n18813 = i_hbusreq3 & ~n18812;
  assign n18814 = i_hbusreq2 & ~n18801;
  assign n18815 = ~n12172 & ~n18788;
  assign n18816 = ~i_hbusreq2 & ~n18815;
  assign n18817 = ~n18814 & ~n18816;
  assign n18818 = ~controllable_hgrant2 & ~n18817;
  assign n18819 = ~n5635 & ~n18818;
  assign n18820 = controllable_hmaster0 & ~n18819;
  assign n18821 = ~n5722 & ~n18818;
  assign n18822 = ~controllable_hmaster0 & ~n18821;
  assign n18823 = ~n18820 & ~n18822;
  assign n18824 = controllable_hmaster1 & ~n18823;
  assign n18825 = ~n12198 & ~n17843;
  assign n18826 = ~i_hbusreq2 & ~n18825;
  assign n18827 = ~n9325 & ~n18826;
  assign n18828 = ~controllable_hgrant2 & ~n18827;
  assign n18829 = ~n5657 & ~n18828;
  assign n18830 = controllable_hmaster0 & ~n18829;
  assign n18831 = ~controllable_hmaster0 & ~n18819;
  assign n18832 = ~n18830 & ~n18831;
  assign n18833 = ~controllable_hmaster1 & ~n18832;
  assign n18834 = ~n18824 & ~n18833;
  assign n18835 = ~i_hbusreq3 & ~n18834;
  assign n18836 = ~n18813 & ~n18835;
  assign n18837 = ~controllable_hmaster2 & ~n18836;
  assign n18838 = ~n18800 & ~n18837;
  assign n18839 = ~controllable_hgrant3 & ~n18838;
  assign n18840 = ~n18453 & ~n18839;
  assign n18841 = controllable_nhgrant0 & ~n18840;
  assign n18842 = ~n18526 & ~n18841;
  assign n18843 = ~n3281 & ~n18842;
  assign n18844 = ~n4089 & ~n18843;
  assign n18845 = n3378 & ~n18844;
  assign n18846 = ~n9253 & ~n12410;
  assign n18847 = ~controllable_hmaster1 & ~n18846;
  assign n18848 = ~n9252 & ~n18847;
  assign n18849 = i_hbusreq3 & ~n18848;
  assign n18850 = ~n9264 & ~n17777;
  assign n18851 = ~i_hbusreq0 & ~n18850;
  assign n18852 = ~n9260 & ~n18851;
  assign n18853 = ~i_hbusreq4 & ~n18852;
  assign n18854 = ~n9259 & ~n18853;
  assign n18855 = ~controllable_hgrant4 & ~n18854;
  assign n18856 = ~n5863 & ~n18855;
  assign n18857 = ~i_hbusreq2 & ~n18856;
  assign n18858 = ~n9258 & ~n18857;
  assign n18859 = ~controllable_hgrant2 & ~n18858;
  assign n18860 = ~n5862 & ~n18859;
  assign n18861 = controllable_hmaster1 & ~n18860;
  assign n18862 = controllable_hmaster0 & ~n18860;
  assign n18863 = ~n12421 & ~n18862;
  assign n18864 = ~controllable_hmaster1 & ~n18863;
  assign n18865 = ~n18861 & ~n18864;
  assign n18866 = ~i_hbusreq3 & ~n18865;
  assign n18867 = ~n18849 & ~n18866;
  assign n18868 = controllable_hmaster2 & ~n18867;
  assign n18869 = ~n6481 & ~n9309;
  assign n18870 = ~controllable_hmaster1 & ~n18869;
  assign n18871 = ~n6473 & ~n18870;
  assign n18872 = i_hbusreq3 & ~n18871;
  assign n18873 = ~n9334 & ~n17832;
  assign n18874 = ~i_hbusreq0 & ~n18873;
  assign n18875 = ~n9327 & ~n18874;
  assign n18876 = ~i_hbusreq4 & ~n18875;
  assign n18877 = ~n9326 & ~n18876;
  assign n18878 = ~controllable_hgrant4 & n18877;
  assign n18879 = ~n5863 & ~n18878;
  assign n18880 = ~i_hbusreq2 & ~n18879;
  assign n18881 = ~n9325 & ~n18880;
  assign n18882 = ~controllable_hgrant2 & ~n18881;
  assign n18883 = ~n5862 & ~n18882;
  assign n18884 = controllable_hmaster0 & ~n18883;
  assign n18885 = ~n6548 & ~n18884;
  assign n18886 = ~controllable_hmaster1 & ~n18885;
  assign n18887 = ~n6508 & ~n18886;
  assign n18888 = ~i_hbusreq3 & ~n18887;
  assign n18889 = ~n18872 & ~n18888;
  assign n18890 = ~controllable_hmaster2 & ~n18889;
  assign n18891 = ~n18868 & ~n18890;
  assign n18892 = ~controllable_hgrant3 & ~n18891;
  assign n18893 = ~n5861 & ~n18892;
  assign n18894 = controllable_nhgrant0 & ~n18893;
  assign n18895 = ~n6082 & ~n18894;
  assign n18896 = ~n3281 & ~n18895;
  assign n18897 = ~n4089 & ~n18896;
  assign n18898 = ~n3378 & ~n18897;
  assign n18899 = ~n18845 & ~n18898;
  assign n18900 = n3492 & ~n18899;
  assign n18901 = ~n18630 & ~n18900;
  assign n18902 = n3485 & ~n18901;
  assign n18903 = ~n18629 & ~n18902;
  assign n18904 = n3476 & ~n18903;
  assign n18905 = ~n18758 & ~n18904;
  assign n18906 = n3374 & ~n18905;
  assign n18907 = ~n18636 & ~n18906;
  assign n18908 = ~n3655 & ~n18907;
  assign n18909 = ~n18570 & ~n18908;
  assign n18910 = n3652 & ~n18909;
  assign n18911 = ~n6665 & ~n18369;
  assign n18912 = n3492 & ~n18911;
  assign n18913 = ~n3631 & ~n18912;
  assign n18914 = n3485 & ~n18913;
  assign n18915 = ~n3630 & ~n18914;
  assign n18916 = ~n3374 & ~n18915;
  assign n18917 = ~n3821 & ~n9440;
  assign n18918 = ~controllable_hmaster1 & ~n18917;
  assign n18919 = ~n5293 & ~n18918;
  assign n18920 = i_hbusreq3 & ~n18919;
  assign n18921 = ~n5278 & ~n9453;
  assign n18922 = ~controllable_hmaster1 & ~n18921;
  assign n18923 = ~n5313 & ~n18922;
  assign n18924 = ~i_hbusreq3 & ~n18923;
  assign n18925 = ~n18920 & ~n18924;
  assign n18926 = ~controllable_hmaster2 & ~n18925;
  assign n18927 = ~n12065 & ~n18926;
  assign n18928 = ~controllable_hgrant3 & ~n18927;
  assign n18929 = ~n18382 & ~n18928;
  assign n18930 = controllable_nhgrant0 & ~n18929;
  assign n18931 = ~n18416 & ~n18930;
  assign n18932 = ~n3281 & ~n18931;
  assign n18933 = ~n3950 & ~n18932;
  assign n18934 = n3378 & ~n18933;
  assign n18935 = ~n6704 & ~n9440;
  assign n18936 = ~controllable_hmaster1 & ~n18935;
  assign n18937 = ~n6701 & ~n18936;
  assign n18938 = i_hbusreq3 & ~n18937;
  assign n18939 = ~n6717 & ~n9453;
  assign n18940 = ~controllable_hmaster1 & ~n18939;
  assign n18941 = ~n6714 & ~n18940;
  assign n18942 = ~i_hbusreq3 & ~n18941;
  assign n18943 = ~n18938 & ~n18942;
  assign n18944 = ~controllable_hmaster2 & ~n18943;
  assign n18945 = ~n12501 & ~n18944;
  assign n18946 = ~controllable_hgrant3 & ~n18945;
  assign n18947 = ~n5402 & ~n18946;
  assign n18948 = controllable_nhgrant0 & ~n18947;
  assign n18949 = ~n5534 & ~n18948;
  assign n18950 = ~n3281 & ~n18949;
  assign n18951 = ~n3950 & ~n18950;
  assign n18952 = ~n3378 & ~n18951;
  assign n18953 = ~n18934 & ~n18952;
  assign n18954 = n3492 & ~n18953;
  assign n18955 = ~n3631 & ~n18954;
  assign n18956 = n3485 & ~n18955;
  assign n18957 = ~n3630 & ~n18956;
  assign n18958 = ~n3476 & ~n18957;
  assign n18959 = ~n6738 & ~n8989;
  assign n18960 = controllable_hmaster0 & ~n18959;
  assign n18961 = ~n5702 & ~n18960;
  assign n18962 = ~controllable_hmaster1 & ~n18961;
  assign n18963 = ~n5690 & ~n18962;
  assign n18964 = i_hbusreq3 & ~n18963;
  assign n18965 = ~n6745 & ~n18499;
  assign n18966 = controllable_hmaster0 & ~n18965;
  assign n18967 = ~n18502 & ~n18966;
  assign n18968 = ~controllable_hmaster1 & ~n18967;
  assign n18969 = ~n18495 & ~n18968;
  assign n18970 = ~i_hbusreq3 & ~n18969;
  assign n18971 = ~n18964 & ~n18970;
  assign n18972 = ~controllable_hmaster2 & ~n18971;
  assign n18973 = ~n18481 & ~n18972;
  assign n18974 = ~controllable_hgrant3 & ~n18973;
  assign n18975 = ~n18453 & ~n18974;
  assign n18976 = controllable_nhgrant0 & ~n18975;
  assign n18977 = ~n18526 & ~n18976;
  assign n18978 = ~n3281 & ~n18977;
  assign n18979 = ~n4089 & ~n18978;
  assign n18980 = n3378 & ~n18979;
  assign n18981 = ~n6793 & ~n9502;
  assign n18982 = ~controllable_hmaster1 & ~n18981;
  assign n18983 = ~n6790 & ~n18982;
  assign n18984 = i_hbusreq3 & ~n18983;
  assign n18985 = ~n6772 & ~n18544;
  assign n18986 = controllable_hmaster0 & ~n18985;
  assign n18987 = ~n6833 & ~n18986;
  assign n18988 = ~controllable_hmaster1 & ~n18987;
  assign n18989 = ~n6817 & ~n18988;
  assign n18990 = ~i_hbusreq3 & ~n18989;
  assign n18991 = ~n18984 & ~n18990;
  assign n18992 = ~controllable_hmaster2 & ~n18991;
  assign n18993 = ~n12561 & ~n18992;
  assign n18994 = ~controllable_hgrant3 & ~n18993;
  assign n18995 = ~n5861 & ~n18994;
  assign n18996 = controllable_nhgrant0 & ~n18995;
  assign n18997 = ~n6082 & ~n18996;
  assign n18998 = ~n3281 & ~n18997;
  assign n18999 = ~n4089 & ~n18998;
  assign n19000 = ~n3378 & ~n18999;
  assign n19001 = ~n18980 & ~n19000;
  assign n19002 = n3492 & ~n19001;
  assign n19003 = ~n3631 & ~n19002;
  assign n19004 = n3485 & ~n19003;
  assign n19005 = ~n3630 & ~n19004;
  assign n19006 = n3476 & ~n19005;
  assign n19007 = ~n18958 & ~n19006;
  assign n19008 = n3374 & ~n19007;
  assign n19009 = ~n18916 & ~n19008;
  assign n19010 = n3655 & ~n19009;
  assign n19011 = ~n4333 & ~n18580;
  assign n19012 = controllable_hmaster1 & ~n19011;
  assign n19013 = controllable_hmaster0 & ~n19011;
  assign n19014 = ~n3729 & ~n19013;
  assign n19015 = ~controllable_hmaster1 & ~n19014;
  assign n19016 = ~n19012 & ~n19015;
  assign n19017 = i_hbusreq3 & ~n19016;
  assign n19018 = ~n4340 & ~n18605;
  assign n19019 = controllable_hmaster1 & ~n19018;
  assign n19020 = controllable_hmaster0 & ~n19018;
  assign n19021 = ~n3767 & ~n19020;
  assign n19022 = ~controllable_hmaster1 & ~n19021;
  assign n19023 = ~n19019 & ~n19022;
  assign n19024 = ~i_hbusreq3 & ~n19023;
  assign n19025 = ~n19017 & ~n19024;
  assign n19026 = controllable_hmaster2 & ~n19025;
  assign n19027 = ~n6887 & ~n19026;
  assign n19028 = ~controllable_hgrant3 & ~n19027;
  assign n19029 = ~n5037 & ~n19028;
  assign n19030 = controllable_nhgrant0 & ~n19029;
  assign n19031 = ~n5245 & ~n19030;
  assign n19032 = ~n3281 & ~n19031;
  assign n19033 = ~n3783 & ~n19032;
  assign n19034 = ~n3378 & ~n19033;
  assign n19035 = ~n18571 & ~n19034;
  assign n19036 = n3492 & ~n19035;
  assign n19037 = ~n3631 & ~n19036;
  assign n19038 = n3485 & ~n19037;
  assign n19039 = ~n3630 & ~n19038;
  assign n19040 = ~n3476 & ~n19039;
  assign n19041 = ~n18630 & ~n19036;
  assign n19042 = n3485 & ~n19041;
  assign n19043 = ~n18629 & ~n19042;
  assign n19044 = n3476 & ~n19043;
  assign n19045 = ~n19040 & ~n19044;
  assign n19046 = ~n3374 & ~n19045;
  assign n19047 = ~n9594 & ~n18679;
  assign n19048 = ~controllable_hmaster1 & ~n19047;
  assign n19049 = ~n18678 & ~n19048;
  assign n19050 = i_hbusreq3 & ~n19049;
  assign n19051 = ~n9607 & ~n18695;
  assign n19052 = ~controllable_hmaster1 & ~n19051;
  assign n19053 = ~n18694 & ~n19052;
  assign n19054 = ~i_hbusreq3 & ~n19053;
  assign n19055 = ~n19050 & ~n19054;
  assign n19056 = ~controllable_hmaster2 & ~n19055;
  assign n19057 = ~n18670 & ~n19056;
  assign n19058 = ~controllable_hgrant3 & ~n19057;
  assign n19059 = ~n18382 & ~n19058;
  assign n19060 = controllable_nhgrant0 & ~n19059;
  assign n19061 = ~n18416 & ~n19060;
  assign n19062 = ~n3281 & ~n19061;
  assign n19063 = ~n3950 & ~n19062;
  assign n19064 = n3378 & ~n19063;
  assign n19065 = ~n4333 & ~n9114;
  assign n19066 = controllable_hmaster1 & ~n19065;
  assign n19067 = controllable_hmaster0 & ~n19065;
  assign n19068 = ~n12617 & ~n19067;
  assign n19069 = ~controllable_hmaster1 & ~n19068;
  assign n19070 = ~n19066 & ~n19069;
  assign n19071 = i_hbusreq3 & ~n19070;
  assign n19072 = ~n4340 & ~n18725;
  assign n19073 = controllable_hmaster1 & ~n19072;
  assign n19074 = controllable_hmaster0 & ~n19072;
  assign n19075 = ~n12623 & ~n19074;
  assign n19076 = ~controllable_hmaster1 & ~n19075;
  assign n19077 = ~n19073 & ~n19076;
  assign n19078 = ~i_hbusreq3 & ~n19077;
  assign n19079 = ~n19071 & ~n19078;
  assign n19080 = controllable_hmaster2 & ~n19079;
  assign n19081 = ~n6934 & ~n9594;
  assign n19082 = ~controllable_hmaster1 & ~n19081;
  assign n19083 = ~n6931 & ~n19082;
  assign n19084 = i_hbusreq3 & ~n19083;
  assign n19085 = ~n6949 & ~n9607;
  assign n19086 = ~controllable_hmaster1 & ~n19085;
  assign n19087 = ~n6944 & ~n19086;
  assign n19088 = ~i_hbusreq3 & ~n19087;
  assign n19089 = ~n19084 & ~n19088;
  assign n19090 = ~controllable_hmaster2 & ~n19089;
  assign n19091 = ~n19080 & ~n19090;
  assign n19092 = ~controllable_hgrant3 & ~n19091;
  assign n19093 = ~n5402 & ~n19092;
  assign n19094 = controllable_nhgrant0 & ~n19093;
  assign n19095 = ~n5534 & ~n19094;
  assign n19096 = ~n3281 & ~n19095;
  assign n19097 = ~n3950 & ~n19096;
  assign n19098 = ~n3378 & ~n19097;
  assign n19099 = ~n19064 & ~n19098;
  assign n19100 = n3492 & ~n19099;
  assign n19101 = ~n3631 & ~n19100;
  assign n19102 = n3485 & ~n19101;
  assign n19103 = ~n3630 & ~n19102;
  assign n19104 = ~n3476 & ~n19103;
  assign n19105 = ~n6738 & ~n9307;
  assign n19106 = controllable_hmaster0 & ~n19105;
  assign n19107 = ~n18809 & ~n19106;
  assign n19108 = ~controllable_hmaster1 & ~n19107;
  assign n19109 = ~n18808 & ~n19108;
  assign n19110 = i_hbusreq3 & ~n19109;
  assign n19111 = ~n6745 & ~n18828;
  assign n19112 = controllable_hmaster0 & ~n19111;
  assign n19113 = ~n18831 & ~n19112;
  assign n19114 = ~controllable_hmaster1 & ~n19113;
  assign n19115 = ~n18824 & ~n19114;
  assign n19116 = ~i_hbusreq3 & ~n19115;
  assign n19117 = ~n19110 & ~n19116;
  assign n19118 = ~controllable_hmaster2 & ~n19117;
  assign n19119 = ~n18800 & ~n19118;
  assign n19120 = ~controllable_hgrant3 & ~n19119;
  assign n19121 = ~n18453 & ~n19120;
  assign n19122 = controllable_nhgrant0 & ~n19121;
  assign n19123 = ~n18526 & ~n19122;
  assign n19124 = ~n3281 & ~n19123;
  assign n19125 = ~n4089 & ~n19124;
  assign n19126 = n3378 & ~n19125;
  assign n19127 = ~n6762 & ~n9250;
  assign n19128 = controllable_hmaster1 & ~n19127;
  assign n19129 = controllable_hmaster0 & ~n19127;
  assign n19130 = ~n12677 & ~n19129;
  assign n19131 = ~controllable_hmaster1 & ~n19130;
  assign n19132 = ~n19128 & ~n19131;
  assign n19133 = i_hbusreq3 & ~n19132;
  assign n19134 = ~n6772 & ~n18859;
  assign n19135 = controllable_hmaster1 & ~n19134;
  assign n19136 = controllable_hmaster0 & ~n19134;
  assign n19137 = ~n12683 & ~n19136;
  assign n19138 = ~controllable_hmaster1 & ~n19137;
  assign n19139 = ~n19135 & ~n19138;
  assign n19140 = ~i_hbusreq3 & ~n19139;
  assign n19141 = ~n19133 & ~n19140;
  assign n19142 = controllable_hmaster2 & ~n19141;
  assign n19143 = ~n7020 & ~n9654;
  assign n19144 = ~controllable_hmaster1 & ~n19143;
  assign n19145 = ~n7017 & ~n19144;
  assign n19146 = i_hbusreq3 & ~n19145;
  assign n19147 = ~n6772 & ~n18882;
  assign n19148 = controllable_hmaster0 & ~n19147;
  assign n19149 = ~n7034 & ~n19148;
  assign n19150 = ~controllable_hmaster1 & ~n19149;
  assign n19151 = ~n7030 & ~n19150;
  assign n19152 = ~i_hbusreq3 & ~n19151;
  assign n19153 = ~n19146 & ~n19152;
  assign n19154 = ~controllable_hmaster2 & ~n19153;
  assign n19155 = ~n19142 & ~n19154;
  assign n19156 = ~controllable_hgrant3 & ~n19155;
  assign n19157 = ~n5861 & ~n19156;
  assign n19158 = controllable_nhgrant0 & ~n19157;
  assign n19159 = ~n6082 & ~n19158;
  assign n19160 = ~n3281 & ~n19159;
  assign n19161 = ~n4089 & ~n19160;
  assign n19162 = ~n3378 & ~n19161;
  assign n19163 = ~n19126 & ~n19162;
  assign n19164 = n3492 & ~n19163;
  assign n19165 = ~n18630 & ~n19164;
  assign n19166 = n3485 & ~n19165;
  assign n19167 = ~n18629 & ~n19166;
  assign n19168 = n3476 & ~n19167;
  assign n19169 = ~n19104 & ~n19168;
  assign n19170 = n3374 & ~n19169;
  assign n19171 = ~n19046 & ~n19170;
  assign n19172 = ~n3655 & ~n19171;
  assign n19173 = ~n19010 & ~n19172;
  assign n19174 = ~n3652 & ~n19173;
  assign n19175 = ~n18910 & ~n19174;
  assign n19176 = ~n3368 & ~n19175;
  assign n19177 = ~controllable_hmaster1 & ~n12752;
  assign n19178 = ~n5280 & ~n19177;
  assign n19179 = ~i_hbusreq3 & ~n19178;
  assign n19180 = ~n5265 & ~n19179;
  assign n19181 = ~controllable_hmaster2 & ~n19180;
  assign n19182 = ~n12033 & ~n19181;
  assign n19183 = controllable_hgrant3 & ~n19182;
  assign n19184 = ~n5278 & ~n9826;
  assign n19185 = ~controllable_hmaster1 & ~n19184;
  assign n19186 = ~n5313 & ~n19185;
  assign n19187 = ~i_hbusreq3 & ~n19186;
  assign n19188 = ~n18386 & ~n19187;
  assign n19189 = ~controllable_hmaster2 & ~n19188;
  assign n19190 = ~n12741 & ~n19189;
  assign n19191 = ~controllable_hgrant3 & ~n19190;
  assign n19192 = ~n19183 & ~n19191;
  assign n19193 = controllable_nhgrant0 & ~n19192;
  assign n19194 = ~n3400 & ~n19177;
  assign n19195 = ~i_hbusreq3 & ~n19194;
  assign n19196 = ~n3951 & ~n19195;
  assign n19197 = ~controllable_hmaster2 & ~n19196;
  assign n19198 = ~n12033 & ~n19197;
  assign n19199 = controllable_hgrant3 & ~n19198;
  assign n19200 = ~n5348 & ~n9737;
  assign n19201 = ~controllable_hmaster1 & ~n19200;
  assign n19202 = ~n3381 & ~n19201;
  assign n19203 = i_hbusreq3 & ~n19202;
  assign n19204 = ~n5353 & ~n9743;
  assign n19205 = ~controllable_hmaster1 & ~n19204;
  assign n19206 = ~n3400 & ~n19205;
  assign n19207 = ~i_hbusreq3 & ~n19206;
  assign n19208 = ~n19203 & ~n19207;
  assign n19209 = ~controllable_hmaster2 & ~n19208;
  assign n19210 = ~n12033 & ~n19209;
  assign n19211 = ~controllable_hgrant3 & ~n19210;
  assign n19212 = ~n19199 & ~n19211;
  assign n19213 = ~controllable_nhgrant0 & ~n19212;
  assign n19214 = ~n19193 & ~n19213;
  assign n19215 = ~n3281 & ~n19214;
  assign n19216 = ~n3281 & ~n19215;
  assign n19217 = n3378 & ~n19216;
  assign n19218 = ~n5394 & ~n9700;
  assign n19219 = ~controllable_hmaster1 & ~n19218;
  assign n19220 = ~n5379 & ~n19219;
  assign n19221 = ~i_hbusreq3 & ~n19220;
  assign n19222 = ~n5265 & ~n19221;
  assign n19223 = ~controllable_hmaster2 & ~n19222;
  assign n19224 = ~n5370 & ~n19223;
  assign n19225 = controllable_hgrant3 & ~n19224;
  assign n19226 = ~n5478 & ~n9826;
  assign n19227 = ~controllable_hmaster1 & ~n19226;
  assign n19228 = ~n5442 & ~n19227;
  assign n19229 = ~i_hbusreq3 & ~n19228;
  assign n19230 = ~n18424 & ~n19229;
  assign n19231 = ~controllable_hmaster2 & ~n19230;
  assign n19232 = ~n12795 & ~n19231;
  assign n19233 = ~controllable_hgrant3 & ~n19232;
  assign n19234 = ~n19225 & ~n19233;
  assign n19235 = controllable_nhgrant0 & ~n19234;
  assign n19236 = ~n4912 & ~n19219;
  assign n19237 = ~i_hbusreq3 & ~n19236;
  assign n19238 = ~n3951 & ~n19237;
  assign n19239 = ~controllable_hmaster2 & ~n19238;
  assign n19240 = ~n5370 & ~n19239;
  assign n19241 = controllable_hgrant3 & ~n19240;
  assign n19242 = ~n5499 & ~n9737;
  assign n19243 = ~controllable_hmaster1 & ~n19242;
  assign n19244 = ~n5190 & ~n19243;
  assign n19245 = i_hbusreq3 & ~n19244;
  assign n19246 = ~n5524 & ~n9743;
  assign n19247 = ~controllable_hmaster1 & ~n19246;
  assign n19248 = ~n5196 & ~n19247;
  assign n19249 = ~i_hbusreq3 & ~n19248;
  assign n19250 = ~n19245 & ~n19249;
  assign n19251 = ~controllable_hmaster2 & ~n19250;
  assign n19252 = ~n5498 & ~n19251;
  assign n19253 = ~controllable_hgrant3 & ~n19252;
  assign n19254 = ~n19241 & ~n19253;
  assign n19255 = ~controllable_nhgrant0 & ~n19254;
  assign n19256 = ~n19235 & ~n19255;
  assign n19257 = ~n3281 & ~n19256;
  assign n19258 = ~n3281 & ~n19257;
  assign n19259 = ~n3378 & ~n19258;
  assign n19260 = ~n19217 & ~n19259;
  assign n19261 = n3492 & ~n19260;
  assign n19262 = n3492 & ~n19261;
  assign n19263 = n3485 & ~n19262;
  assign n19264 = n3485 & ~n19263;
  assign n19265 = ~n3476 & ~n19264;
  assign n19266 = controllable_hmaster0 & ~n7231;
  assign n19267 = ~n5606 & ~n19266;
  assign n19268 = ~controllable_hmaster1 & ~n19267;
  assign n19269 = ~n5608 & ~n19268;
  assign n19270 = ~i_hbusreq3 & ~n19269;
  assign n19271 = ~n5593 & ~n19270;
  assign n19272 = ~controllable_hmaster2 & ~n19271;
  assign n19273 = ~n12233 & ~n19272;
  assign n19274 = controllable_hgrant3 & ~n19273;
  assign n19275 = ~n7272 & ~n17429;
  assign n19276 = ~controllable_ndecide & ~n19275;
  assign n19277 = ~controllable_ndecide & ~n19276;
  assign n19278 = i_hready & ~n19277;
  assign n19279 = ~n3392 & ~n19278;
  assign n19280 = ~i_hbusreq0 & ~n19279;
  assign n19281 = ~n7271 & ~n19280;
  assign n19282 = ~i_hbusreq4 & ~n19281;
  assign n19283 = ~n7270 & ~n19282;
  assign n19284 = ~controllable_hgrant4 & ~n19283;
  assign n19285 = ~n12172 & ~n19284;
  assign n19286 = ~i_hbusreq2 & ~n19285;
  assign n19287 = ~n7264 & ~n19286;
  assign n19288 = ~controllable_hgrant2 & ~n19287;
  assign n19289 = ~n5635 & ~n19288;
  assign n19290 = controllable_hmaster1 & ~n19289;
  assign n19291 = controllable_hmaster0 & ~n19289;
  assign n19292 = ~n7294 & ~n17429;
  assign n19293 = ~controllable_ndecide & ~n19292;
  assign n19294 = ~controllable_ndecide & ~n19293;
  assign n19295 = i_hready & ~n19294;
  assign n19296 = ~n3392 & ~n19295;
  assign n19297 = ~i_hbusreq0 & ~n19296;
  assign n19298 = ~n7347 & ~n19297;
  assign n19299 = ~i_hbusreq4 & ~n19298;
  assign n19300 = ~n7346 & ~n19299;
  assign n19301 = ~controllable_hgrant4 & ~n19300;
  assign n19302 = ~n12181 & ~n19301;
  assign n19303 = ~i_hbusreq2 & ~n19302;
  assign n19304 = ~n12872 & ~n19303;
  assign n19305 = ~controllable_hgrant2 & ~n19304;
  assign n19306 = ~n5635 & ~n19305;
  assign n19307 = ~controllable_hmaster0 & ~n19306;
  assign n19308 = ~n19291 & ~n19307;
  assign n19309 = ~controllable_hmaster1 & ~n19308;
  assign n19310 = ~n19290 & ~n19309;
  assign n19311 = ~i_hbusreq3 & ~n19310;
  assign n19312 = ~n12864 & ~n19311;
  assign n19313 = controllable_hmaster2 & ~n19312;
  assign n19314 = ~n3495 & ~n7333;
  assign n19315 = ~controllable_hgrant4 & ~n19314;
  assign n19316 = ~n4091 & ~n19315;
  assign n19317 = ~controllable_hgrant2 & ~n19316;
  assign n19318 = ~n5616 & ~n19317;
  assign n19319 = controllable_hmaster0 & ~n19318;
  assign n19320 = ~n7340 & ~n19319;
  assign n19321 = ~controllable_hmaster1 & ~n19320;
  assign n19322 = ~n7330 & ~n19321;
  assign n19323 = i_hbusreq3 & ~n19322;
  assign n19324 = ~n12172 & ~n19301;
  assign n19325 = ~i_hbusreq2 & ~n19324;
  assign n19326 = ~n7345 & ~n19325;
  assign n19327 = ~controllable_hgrant2 & ~n19326;
  assign n19328 = ~n5635 & ~n19327;
  assign n19329 = controllable_hmaster0 & ~n19328;
  assign n19330 = ~n5722 & ~n19327;
  assign n19331 = ~controllable_hmaster0 & ~n19330;
  assign n19332 = ~n19329 & ~n19331;
  assign n19333 = controllable_hmaster1 & ~n19332;
  assign n19334 = i_hbusreq2 & ~n19316;
  assign n19335 = i_hbusreq4 & ~n19314;
  assign n19336 = i_hbusreq0 & ~n19314;
  assign n19337 = ~n7367 & ~n18087;
  assign n19338 = ~controllable_ndecide & n19337;
  assign n19339 = ~controllable_ndecide & ~n19338;
  assign n19340 = i_hready & ~n19339;
  assign n19341 = ~n4577 & ~n19340;
  assign n19342 = i_hlock0 & ~n19341;
  assign n19343 = ~n7367 & ~n17487;
  assign n19344 = ~controllable_ndecide & n19343;
  assign n19345 = ~controllable_ndecide & ~n19344;
  assign n19346 = i_hready & ~n19345;
  assign n19347 = ~n3495 & ~n19346;
  assign n19348 = ~i_hlock0 & ~n19347;
  assign n19349 = ~n19342 & ~n19348;
  assign n19350 = ~i_hbusreq0 & ~n19349;
  assign n19351 = ~n19336 & ~n19350;
  assign n19352 = ~i_hbusreq4 & ~n19351;
  assign n19353 = ~n19335 & ~n19352;
  assign n19354 = ~controllable_hgrant4 & ~n19353;
  assign n19355 = ~n12894 & ~n19354;
  assign n19356 = ~i_hbusreq2 & ~n19355;
  assign n19357 = ~n19334 & ~n19356;
  assign n19358 = ~controllable_hgrant2 & ~n19357;
  assign n19359 = ~n7290 & ~n19358;
  assign n19360 = controllable_hmaster0 & ~n19359;
  assign n19361 = ~controllable_hmaster0 & ~n19328;
  assign n19362 = ~n19360 & ~n19361;
  assign n19363 = ~controllable_hmaster1 & ~n19362;
  assign n19364 = ~n19333 & ~n19363;
  assign n19365 = ~i_hbusreq3 & ~n19364;
  assign n19366 = ~n19323 & ~n19365;
  assign n19367 = ~controllable_hmaster2 & ~n19366;
  assign n19368 = ~n19313 & ~n19367;
  assign n19369 = ~controllable_hgrant3 & ~n19368;
  assign n19370 = ~n19274 & ~n19369;
  assign n19371 = controllable_nhgrant0 & ~n19370;
  assign n19372 = ~n5794 & ~n12927;
  assign n19373 = ~controllable_hmaster1 & ~n19372;
  assign n19374 = ~n5757 & ~n19373;
  assign n19375 = i_hbusreq3 & ~n19374;
  assign n19376 = ~n5799 & ~n12932;
  assign n19377 = ~controllable_hmaster1 & ~n19376;
  assign n19378 = ~n5561 & ~n19377;
  assign n19379 = ~i_hbusreq3 & ~n19378;
  assign n19380 = ~n19375 & ~n19379;
  assign n19381 = ~controllable_hmaster2 & ~n19380;
  assign n19382 = ~n12233 & ~n19381;
  assign n19383 = ~controllable_hgrant3 & ~n19382;
  assign n19384 = ~n19199 & ~n19383;
  assign n19385 = ~controllable_nhgrant0 & ~n19384;
  assign n19386 = ~n19371 & ~n19385;
  assign n19387 = ~n3281 & ~n19386;
  assign n19388 = ~n3281 & ~n19387;
  assign n19389 = n3378 & ~n19388;
  assign n19390 = controllable_hmaster0 & ~n7448;
  assign n19391 = ~n5853 & ~n19390;
  assign n19392 = ~controllable_hmaster1 & ~n19391;
  assign n19393 = ~n5838 & ~n19392;
  assign n19394 = ~i_hbusreq3 & ~n19393;
  assign n19395 = ~n5593 & ~n19394;
  assign n19396 = ~controllable_hmaster2 & ~n19395;
  assign n19397 = ~n5828 & ~n19396;
  assign n19398 = controllable_hgrant3 & ~n19397;
  assign n19399 = ~n5038 & ~n19276;
  assign n19400 = i_hready & ~n19399;
  assign n19401 = ~n5055 & ~n19400;
  assign n19402 = i_hlock0 & ~n19401;
  assign n19403 = ~n7493 & ~n19402;
  assign n19404 = ~i_hbusreq0 & ~n19403;
  assign n19405 = ~n7488 & ~n19404;
  assign n19406 = ~i_hbusreq4 & ~n19405;
  assign n19407 = ~n7487 & ~n19406;
  assign n19408 = ~controllable_hgrant4 & ~n19407;
  assign n19409 = ~n5863 & ~n19408;
  assign n19410 = ~i_hbusreq2 & ~n19409;
  assign n19411 = ~n7479 & ~n19410;
  assign n19412 = ~controllable_hgrant2 & ~n19411;
  assign n19413 = ~n5862 & ~n19412;
  assign n19414 = controllable_hmaster1 & ~n19413;
  assign n19415 = controllable_hmaster0 & ~n19413;
  assign n19416 = ~n3903 & ~n19293;
  assign n19417 = i_hready & ~n19416;
  assign n19418 = ~n3920 & ~n19417;
  assign n19419 = i_hlock0 & ~n19418;
  assign n19420 = ~n7562 & ~n19419;
  assign n19421 = ~i_hbusreq0 & ~n19420;
  assign n19422 = ~n7559 & ~n19421;
  assign n19423 = ~i_hbusreq4 & ~n19422;
  assign n19424 = ~n7558 & ~n19423;
  assign n19425 = ~controllable_hgrant4 & ~n19424;
  assign n19426 = ~n4064 & ~n19425;
  assign n19427 = ~i_hbusreq2 & ~n19426;
  assign n19428 = ~n12990 & ~n19427;
  assign n19429 = ~controllable_hgrant2 & ~n19428;
  assign n19430 = ~n5862 & ~n19429;
  assign n19431 = ~controllable_hmaster0 & ~n19430;
  assign n19432 = ~n19415 & ~n19431;
  assign n19433 = ~controllable_hmaster1 & ~n19432;
  assign n19434 = ~n19414 & ~n19433;
  assign n19435 = ~i_hbusreq3 & ~n19434;
  assign n19436 = ~n12982 & ~n19435;
  assign n19437 = controllable_hmaster2 & ~n19436;
  assign n19438 = ~n3495 & ~n7545;
  assign n19439 = ~controllable_hgrant4 & ~n19438;
  assign n19440 = ~n4091 & ~n19439;
  assign n19441 = ~controllable_hgrant2 & ~n19440;
  assign n19442 = ~n5616 & ~n19441;
  assign n19443 = controllable_hmaster0 & ~n19442;
  assign n19444 = ~n7552 & ~n19443;
  assign n19445 = ~controllable_hmaster1 & ~n19444;
  assign n19446 = ~n7543 & ~n19445;
  assign n19447 = i_hbusreq3 & ~n19446;
  assign n19448 = ~n5863 & ~n19425;
  assign n19449 = ~i_hbusreq2 & ~n19448;
  assign n19450 = ~n7557 & ~n19449;
  assign n19451 = ~controllable_hgrant2 & ~n19450;
  assign n19452 = ~n5862 & ~n19451;
  assign n19453 = controllable_hmaster0 & ~n19452;
  assign n19454 = ~n5950 & ~n19451;
  assign n19455 = ~controllable_hmaster0 & ~n19454;
  assign n19456 = ~n19453 & ~n19455;
  assign n19457 = controllable_hmaster1 & ~n19456;
  assign n19458 = i_hbusreq2 & ~n19440;
  assign n19459 = i_hbusreq4 & ~n19438;
  assign n19460 = i_hbusreq0 & ~n19438;
  assign n19461 = ~n3903 & ~n19338;
  assign n19462 = i_hready & ~n19461;
  assign n19463 = ~n4577 & ~n19462;
  assign n19464 = i_hlock0 & ~n19463;
  assign n19465 = ~i_hlock0 & ~n19438;
  assign n19466 = ~n19464 & ~n19465;
  assign n19467 = ~i_hbusreq0 & ~n19466;
  assign n19468 = ~n19460 & ~n19467;
  assign n19469 = ~i_hbusreq4 & ~n19468;
  assign n19470 = ~n19459 & ~n19469;
  assign n19471 = ~controllable_hgrant4 & ~n19470;
  assign n19472 = ~n13012 & ~n19471;
  assign n19473 = ~i_hbusreq2 & ~n19472;
  assign n19474 = ~n19458 & ~n19473;
  assign n19475 = ~controllable_hgrant2 & ~n19474;
  assign n19476 = ~n7507 & ~n19475;
  assign n19477 = controllable_hmaster0 & ~n19476;
  assign n19478 = ~n5464 & ~n19417;
  assign n19479 = i_hlock0 & ~n19478;
  assign n19480 = ~n7562 & ~n19479;
  assign n19481 = ~i_hbusreq0 & ~n19480;
  assign n19482 = ~n7559 & ~n19481;
  assign n19483 = ~i_hbusreq4 & ~n19482;
  assign n19484 = ~n7558 & ~n19483;
  assign n19485 = ~controllable_hgrant4 & ~n19484;
  assign n19486 = ~n5982 & ~n19485;
  assign n19487 = ~i_hbusreq2 & ~n19486;
  assign n19488 = ~n7557 & ~n19487;
  assign n19489 = ~controllable_hgrant2 & ~n19488;
  assign n19490 = ~n5981 & ~n19489;
  assign n19491 = ~controllable_hmaster0 & ~n19490;
  assign n19492 = ~n19477 & ~n19491;
  assign n19493 = ~controllable_hmaster1 & ~n19492;
  assign n19494 = ~n19457 & ~n19493;
  assign n19495 = ~i_hbusreq3 & ~n19494;
  assign n19496 = ~n19447 & ~n19495;
  assign n19497 = ~controllable_hmaster2 & ~n19496;
  assign n19498 = ~n19437 & ~n19497;
  assign n19499 = ~controllable_hgrant3 & ~n19498;
  assign n19500 = ~n19398 & ~n19499;
  assign n19501 = controllable_nhgrant0 & ~n19500;
  assign n19502 = ~n6044 & ~n13049;
  assign n19503 = ~controllable_hmaster1 & ~n19502;
  assign n19504 = ~n6036 & ~n19503;
  assign n19505 = i_hbusreq3 & ~n19504;
  assign n19506 = ~n6072 & ~n13054;
  assign n19507 = ~controllable_hmaster1 & ~n19506;
  assign n19508 = ~n6049 & ~n19507;
  assign n19509 = ~i_hbusreq3 & ~n19508;
  assign n19510 = ~n19505 & ~n19509;
  assign n19511 = ~controllable_hmaster2 & ~n19510;
  assign n19512 = ~n6035 & ~n19511;
  assign n19513 = ~controllable_hgrant3 & ~n19512;
  assign n19514 = ~n19241 & ~n19513;
  assign n19515 = ~controllable_nhgrant0 & ~n19514;
  assign n19516 = ~n19501 & ~n19515;
  assign n19517 = ~n3281 & ~n19516;
  assign n19518 = ~n3281 & ~n19517;
  assign n19519 = ~n3378 & ~n19518;
  assign n19520 = ~n19389 & ~n19519;
  assign n19521 = n3492 & ~n19520;
  assign n19522 = n3492 & ~n19521;
  assign n19523 = n3485 & ~n19522;
  assign n19524 = n3485 & ~n19523;
  assign n19525 = n3476 & ~n19524;
  assign n19526 = ~n19265 & ~n19525;
  assign n19527 = n3374 & ~n19526;
  assign n19528 = ~n7128 & ~n19527;
  assign n19529 = n3655 & ~n19528;
  assign n19530 = controllable_hgrant1 & ~n4697;
  assign n19531 = controllable_ndecide & ~n19530;
  assign n19532 = ~i_hready & n19531;
  assign n19533 = ~n3846 & ~n19532;
  assign n19534 = ~controllable_hgrant4 & ~n19533;
  assign n19535 = ~n3411 & ~n19534;
  assign n19536 = ~controllable_hgrant2 & ~n19535;
  assign n19537 = ~n3410 & ~n19536;
  assign n19538 = controllable_hmaster1 & ~n19537;
  assign n19539 = controllable_hmaster0 & ~n19537;
  assign n19540 = controllable_hmaster0 & ~n19539;
  assign n19541 = ~controllable_hmaster1 & ~n19540;
  assign n19542 = ~n19538 & ~n19541;
  assign n19543 = i_hbusreq3 & ~n19542;
  assign n19544 = i_hbusreq2 & ~n19535;
  assign n19545 = i_hbusreq4 & ~n19533;
  assign n19546 = i_hbusreq0 & ~n19533;
  assign n19547 = ~n3390 & ~n19531;
  assign n19548 = ~i_hready & ~n19547;
  assign n19549 = ~n3864 & ~n19548;
  assign n19550 = ~i_hbusreq0 & ~n19549;
  assign n19551 = ~n19546 & ~n19550;
  assign n19552 = ~i_hbusreq4 & ~n19551;
  assign n19553 = ~n19545 & ~n19552;
  assign n19554 = ~controllable_hgrant4 & ~n19553;
  assign n19555 = ~n3433 & ~n19554;
  assign n19556 = ~i_hbusreq2 & ~n19555;
  assign n19557 = ~n19544 & ~n19556;
  assign n19558 = ~controllable_hgrant2 & ~n19557;
  assign n19559 = ~n3431 & ~n19558;
  assign n19560 = controllable_hmaster1 & ~n19559;
  assign n19561 = controllable_hmaster0 & ~n19559;
  assign n19562 = controllable_hmaster0 & ~n19561;
  assign n19563 = ~controllable_hmaster1 & ~n19562;
  assign n19564 = ~n19560 & ~n19563;
  assign n19565 = ~i_hbusreq3 & ~n19564;
  assign n19566 = ~n19543 & ~n19565;
  assign n19567 = controllable_hmaster2 & ~n19566;
  assign n19568 = controllable_hmaster2 & ~n19567;
  assign n19569 = ~controllable_hgrant3 & ~n19568;
  assign n19570 = ~n3409 & ~n19569;
  assign n19571 = controllable_nhgrant0 & ~n19570;
  assign n19572 = ~n3466 & ~n19571;
  assign n19573 = ~n3281 & ~n19572;
  assign n19574 = ~n3281 & ~n19573;
  assign n19575 = n3378 & ~n19574;
  assign n19576 = ~n4009 & ~n4697;
  assign n19577 = controllable_ndecide & ~n19576;
  assign n19578 = ~i_hready & n19577;
  assign n19579 = ~n3417 & ~n19578;
  assign n19580 = ~controllable_hgrant4 & ~n19579;
  assign n19581 = ~n3411 & ~n19580;
  assign n19582 = ~controllable_hgrant2 & ~n19581;
  assign n19583 = ~n3410 & ~n19582;
  assign n19584 = controllable_hmaster1 & ~n19583;
  assign n19585 = controllable_hmaster0 & ~n19583;
  assign n19586 = controllable_hmaster0 & ~n19585;
  assign n19587 = ~controllable_hmaster1 & ~n19586;
  assign n19588 = ~n19584 & ~n19587;
  assign n19589 = i_hbusreq3 & ~n19588;
  assign n19590 = i_hbusreq2 & ~n19581;
  assign n19591 = i_hbusreq4 & ~n19579;
  assign n19592 = i_hbusreq0 & ~n19579;
  assign n19593 = ~n3390 & ~n19577;
  assign n19594 = ~i_hready & ~n19593;
  assign n19595 = ~n3440 & ~n19594;
  assign n19596 = i_hlock0 & ~n19595;
  assign n19597 = ~i_hlock0 & ~n19579;
  assign n19598 = ~n19596 & ~n19597;
  assign n19599 = ~i_hbusreq0 & ~n19598;
  assign n19600 = ~n19592 & ~n19599;
  assign n19601 = ~i_hbusreq4 & ~n19600;
  assign n19602 = ~n19591 & ~n19601;
  assign n19603 = ~controllable_hgrant4 & ~n19602;
  assign n19604 = ~n3916 & ~n19603;
  assign n19605 = ~i_hbusreq2 & ~n19604;
  assign n19606 = ~n19590 & ~n19605;
  assign n19607 = ~controllable_hgrant2 & ~n19606;
  assign n19608 = ~n3859 & ~n19607;
  assign n19609 = controllable_hmaster1 & ~n19608;
  assign n19610 = controllable_hmaster0 & ~n19608;
  assign n19611 = controllable_hmaster0 & ~n19610;
  assign n19612 = ~controllable_hmaster1 & ~n19611;
  assign n19613 = ~n19609 & ~n19612;
  assign n19614 = ~i_hbusreq3 & ~n19613;
  assign n19615 = ~n19589 & ~n19614;
  assign n19616 = controllable_hmaster2 & ~n19615;
  assign n19617 = controllable_hmaster2 & ~n19616;
  assign n19618 = ~controllable_hgrant3 & ~n19617;
  assign n19619 = ~n7090 & ~n19618;
  assign n19620 = controllable_nhgrant0 & ~n19619;
  assign n19621 = ~n7118 & ~n19620;
  assign n19622 = ~n3281 & ~n19621;
  assign n19623 = ~n3281 & ~n19622;
  assign n19624 = ~n3378 & ~n19623;
  assign n19625 = ~n19575 & ~n19624;
  assign n19626 = n3492 & ~n19625;
  assign n19627 = n3492 & ~n19626;
  assign n19628 = n3485 & ~n19627;
  assign n19629 = n3485 & ~n19628;
  assign n19630 = ~n3374 & ~n19629;
  assign n19631 = ~i_hready & ~n19532;
  assign n19632 = ~controllable_hgrant4 & ~n19631;
  assign n19633 = ~n3848 & ~n19632;
  assign n19634 = ~controllable_hgrant2 & ~n19633;
  assign n19635 = ~n3410 & ~n19634;
  assign n19636 = ~controllable_hmaster0 & ~n19635;
  assign n19637 = ~n19539 & ~n19636;
  assign n19638 = ~controllable_hmaster1 & ~n19637;
  assign n19639 = ~n19538 & ~n19638;
  assign n19640 = i_hbusreq3 & ~n19639;
  assign n19641 = i_hbusreq2 & ~n19633;
  assign n19642 = i_hbusreq4 & ~n19631;
  assign n19643 = i_hbusreq0 & ~n19631;
  assign n19644 = ~i_hready & ~n19548;
  assign n19645 = ~i_hbusreq0 & ~n19644;
  assign n19646 = ~n19643 & ~n19645;
  assign n19647 = ~i_hbusreq4 & ~n19646;
  assign n19648 = ~n19642 & ~n19647;
  assign n19649 = ~controllable_hgrant4 & ~n19648;
  assign n19650 = ~n12052 & ~n19649;
  assign n19651 = ~i_hbusreq2 & ~n19650;
  assign n19652 = ~n19641 & ~n19651;
  assign n19653 = ~controllable_hgrant2 & ~n19652;
  assign n19654 = ~n3431 & ~n19653;
  assign n19655 = ~controllable_hmaster0 & ~n19654;
  assign n19656 = ~n19561 & ~n19655;
  assign n19657 = ~controllable_hmaster1 & ~n19656;
  assign n19658 = ~n19560 & ~n19657;
  assign n19659 = ~i_hbusreq3 & ~n19658;
  assign n19660 = ~n19640 & ~n19659;
  assign n19661 = controllable_hmaster2 & ~n19660;
  assign n19662 = ~n3411 & ~n19632;
  assign n19663 = ~controllable_hgrant2 & ~n19662;
  assign n19664 = ~n3410 & ~n19663;
  assign n19665 = controllable_hmaster0 & ~n19664;
  assign n19666 = ~n5288 & ~n19663;
  assign n19667 = ~controllable_hmaster0 & ~n19666;
  assign n19668 = ~n19665 & ~n19667;
  assign n19669 = controllable_hmaster1 & ~n19668;
  assign n19670 = ~controllable_hmaster0 & ~n19664;
  assign n19671 = ~n10336 & ~n19670;
  assign n19672 = ~controllable_hmaster1 & ~n19671;
  assign n19673 = ~n19669 & ~n19672;
  assign n19674 = i_hbusreq3 & ~n19673;
  assign n19675 = i_hbusreq2 & ~n19662;
  assign n19676 = ~n3433 & ~n19649;
  assign n19677 = ~i_hbusreq2 & ~n19676;
  assign n19678 = ~n19675 & ~n19677;
  assign n19679 = ~controllable_hgrant2 & ~n19678;
  assign n19680 = ~n3431 & ~n19679;
  assign n19681 = controllable_hmaster0 & ~n19680;
  assign n19682 = ~n5308 & ~n19679;
  assign n19683 = ~controllable_hmaster0 & ~n19682;
  assign n19684 = ~n19681 & ~n19683;
  assign n19685 = controllable_hmaster1 & ~n19684;
  assign n19686 = ~controllable_hmaster0 & ~n19680;
  assign n19687 = ~n10376 & ~n19686;
  assign n19688 = ~controllable_hmaster1 & ~n19687;
  assign n19689 = ~n19685 & ~n19688;
  assign n19690 = ~i_hbusreq3 & ~n19689;
  assign n19691 = ~n19674 & ~n19690;
  assign n19692 = ~controllable_hmaster2 & ~n19691;
  assign n19693 = ~n19661 & ~n19692;
  assign n19694 = ~controllable_hgrant3 & ~n19693;
  assign n19695 = ~n19183 & ~n19694;
  assign n19696 = controllable_nhgrant0 & ~n19695;
  assign n19697 = ~n19213 & ~n19696;
  assign n19698 = ~n3281 & ~n19697;
  assign n19699 = ~n3281 & ~n19698;
  assign n19700 = n3378 & ~n19699;
  assign n19701 = ~n3901 & ~n4697;
  assign n19702 = controllable_ndecide & ~n19701;
  assign n19703 = ~i_hready & n19702;
  assign n19704 = ~i_hready & ~n19703;
  assign n19705 = ~controllable_hgrant4 & ~n19704;
  assign n19706 = ~n3848 & ~n19705;
  assign n19707 = ~controllable_hgrant2 & ~n19706;
  assign n19708 = ~n3410 & ~n19707;
  assign n19709 = ~controllable_hmaster0 & ~n19708;
  assign n19710 = ~n19585 & ~n19709;
  assign n19711 = ~controllable_hmaster1 & ~n19710;
  assign n19712 = ~n19584 & ~n19711;
  assign n19713 = i_hbusreq3 & ~n19712;
  assign n19714 = i_hbusreq2 & ~n19706;
  assign n19715 = i_hbusreq4 & ~n19704;
  assign n19716 = i_hbusreq0 & ~n19704;
  assign n19717 = ~n3390 & ~n19702;
  assign n19718 = ~i_hready & ~n19717;
  assign n19719 = ~i_hready & ~n19718;
  assign n19720 = i_hlock0 & ~n19719;
  assign n19721 = ~i_hlock0 & ~n19704;
  assign n19722 = ~n19720 & ~n19721;
  assign n19723 = ~i_hbusreq0 & ~n19722;
  assign n19724 = ~n19716 & ~n19723;
  assign n19725 = ~i_hbusreq4 & ~n19724;
  assign n19726 = ~n19715 & ~n19725;
  assign n19727 = ~controllable_hgrant4 & ~n19726;
  assign n19728 = ~n3873 & ~n19727;
  assign n19729 = ~i_hbusreq2 & ~n19728;
  assign n19730 = ~n19714 & ~n19729;
  assign n19731 = ~controllable_hgrant2 & ~n19730;
  assign n19732 = ~n3859 & ~n19731;
  assign n19733 = ~controllable_hmaster0 & ~n19732;
  assign n19734 = ~n19610 & ~n19733;
  assign n19735 = ~controllable_hmaster1 & ~n19734;
  assign n19736 = ~n19609 & ~n19735;
  assign n19737 = ~i_hbusreq3 & ~n19736;
  assign n19738 = ~n19713 & ~n19737;
  assign n19739 = controllable_hmaster2 & ~n19738;
  assign n19740 = ~n3411 & ~n19705;
  assign n19741 = ~controllable_hgrant2 & ~n19740;
  assign n19742 = ~n3410 & ~n19741;
  assign n19743 = controllable_hmaster0 & ~n19742;
  assign n19744 = ~n5288 & ~n19741;
  assign n19745 = ~controllable_hmaster0 & ~n19744;
  assign n19746 = ~n19743 & ~n19745;
  assign n19747 = controllable_hmaster1 & ~n19746;
  assign n19748 = ~controllable_hmaster0 & ~n19742;
  assign n19749 = ~n10336 & ~n19748;
  assign n19750 = ~controllable_hmaster1 & ~n19749;
  assign n19751 = ~n19747 & ~n19750;
  assign n19752 = i_hbusreq3 & ~n19751;
  assign n19753 = i_hbusreq2 & ~n19740;
  assign n19754 = ~n3916 & ~n19727;
  assign n19755 = ~i_hbusreq2 & ~n19754;
  assign n19756 = ~n19753 & ~n19755;
  assign n19757 = ~controllable_hgrant2 & ~n19756;
  assign n19758 = ~n3859 & ~n19757;
  assign n19759 = controllable_hmaster0 & ~n19758;
  assign n19760 = ~n5438 & ~n19757;
  assign n19761 = ~controllable_hmaster0 & ~n19760;
  assign n19762 = ~n19759 & ~n19761;
  assign n19763 = controllable_hmaster1 & ~n19762;
  assign n19764 = ~n5382 & ~n19702;
  assign n19765 = ~i_hready & ~n19764;
  assign n19766 = ~i_hready & ~n19765;
  assign n19767 = i_hlock0 & ~n19766;
  assign n19768 = ~n19721 & ~n19767;
  assign n19769 = ~i_hbusreq0 & ~n19768;
  assign n19770 = ~n19716 & ~n19769;
  assign n19771 = ~i_hbusreq4 & ~n19770;
  assign n19772 = ~n19715 & ~n19771;
  assign n19773 = ~controllable_hgrant4 & ~n19772;
  assign n19774 = ~n5462 & ~n19773;
  assign n19775 = ~i_hbusreq2 & ~n19774;
  assign n19776 = ~n19753 & ~n19775;
  assign n19777 = ~controllable_hgrant2 & ~n19776;
  assign n19778 = ~n5461 & ~n19777;
  assign n19779 = ~controllable_hmaster0 & ~n19778;
  assign n19780 = ~n10376 & ~n19779;
  assign n19781 = ~controllable_hmaster1 & ~n19780;
  assign n19782 = ~n19763 & ~n19781;
  assign n19783 = ~i_hbusreq3 & ~n19782;
  assign n19784 = ~n19752 & ~n19783;
  assign n19785 = ~controllable_hmaster2 & ~n19784;
  assign n19786 = ~n19739 & ~n19785;
  assign n19787 = ~controllable_hgrant3 & ~n19786;
  assign n19788 = ~n19225 & ~n19787;
  assign n19789 = controllable_nhgrant0 & ~n19788;
  assign n19790 = ~n19255 & ~n19789;
  assign n19791 = ~n3281 & ~n19790;
  assign n19792 = ~n3281 & ~n19791;
  assign n19793 = ~n3378 & ~n19792;
  assign n19794 = ~n19700 & ~n19793;
  assign n19795 = n3492 & ~n19794;
  assign n19796 = n3492 & ~n19795;
  assign n19797 = n3485 & ~n19796;
  assign n19798 = n3485 & ~n19797;
  assign n19799 = ~n3476 & ~n19798;
  assign n19800 = i_hlock1 & ~n18573;
  assign n19801 = ~i_hlock1 & n5864;
  assign n19802 = ~n19800 & ~n19801;
  assign n19803 = ~controllable_ndecide & ~n19802;
  assign n19804 = ~n3494 & ~n19803;
  assign n19805 = i_hready & ~n19804;
  assign n19806 = ~i_hready & ~n19531;
  assign n19807 = ~n19805 & ~n19806;
  assign n19808 = ~controllable_hgrant4 & n19807;
  assign n19809 = ~n4091 & ~n19808;
  assign n19810 = ~controllable_hgrant2 & ~n19809;
  assign n19811 = ~n5616 & ~n19810;
  assign n19812 = controllable_hmaster1 & ~n19811;
  assign n19813 = controllable_hmaster0 & ~n19811;
  assign n19814 = i_hlock1 & ~n9985;
  assign n19815 = ~i_hlock1 & ~controllable_locked;
  assign n19816 = ~n19814 & ~n19815;
  assign n19817 = ~controllable_ndecide & ~n19816;
  assign n19818 = ~n3494 & ~n19817;
  assign n19819 = i_hready & ~n19818;
  assign n19820 = ~n19806 & ~n19819;
  assign n19821 = ~controllable_hgrant4 & n19820;
  assign n19822 = ~n4015 & ~n19821;
  assign n19823 = ~controllable_hgrant2 & ~n19822;
  assign n19824 = ~n5616 & ~n19823;
  assign n19825 = ~controllable_hmaster0 & ~n19824;
  assign n19826 = ~n19813 & ~n19825;
  assign n19827 = ~controllable_hmaster1 & ~n19826;
  assign n19828 = ~n19812 & ~n19827;
  assign n19829 = i_hbusreq3 & ~n19828;
  assign n19830 = i_hbusreq2 & ~n19809;
  assign n19831 = i_hbusreq4 & ~n19807;
  assign n19832 = i_hbusreq0 & ~n19807;
  assign n19833 = i_hbusreq1 & ~n19802;
  assign n19834 = ~n18087 & ~n19833;
  assign n19835 = ~controllable_ndecide & ~n19834;
  assign n19836 = ~n3494 & ~n19835;
  assign n19837 = i_hready & ~n19836;
  assign n19838 = ~i_hready & n19547;
  assign n19839 = ~n19837 & ~n19838;
  assign n19840 = ~i_hbusreq0 & ~n19839;
  assign n19841 = ~n19832 & ~n19840;
  assign n19842 = ~i_hbusreq4 & ~n19841;
  assign n19843 = ~n19831 & ~n19842;
  assign n19844 = ~controllable_hgrant4 & n19843;
  assign n19845 = ~n12172 & ~n19844;
  assign n19846 = ~i_hbusreq2 & ~n19845;
  assign n19847 = ~n19830 & ~n19846;
  assign n19848 = ~controllable_hgrant2 & ~n19847;
  assign n19849 = ~n5635 & ~n19848;
  assign n19850 = controllable_hmaster1 & ~n19849;
  assign n19851 = controllable_hmaster0 & ~n19849;
  assign n19852 = i_hbusreq2 & ~n19822;
  assign n19853 = i_hbusreq4 & ~n19820;
  assign n19854 = i_hbusreq0 & ~n19820;
  assign n19855 = i_hbusreq1 & ~n19816;
  assign n19856 = ~n18087 & ~n19855;
  assign n19857 = ~controllable_ndecide & ~n19856;
  assign n19858 = ~n3494 & ~n19857;
  assign n19859 = i_hready & ~n19858;
  assign n19860 = ~n19838 & ~n19859;
  assign n19861 = ~i_hbusreq0 & ~n19860;
  assign n19862 = ~n19854 & ~n19861;
  assign n19863 = ~i_hbusreq4 & ~n19862;
  assign n19864 = ~n19853 & ~n19863;
  assign n19865 = ~controllable_hgrant4 & n19864;
  assign n19866 = ~n12181 & ~n19865;
  assign n19867 = ~i_hbusreq2 & ~n19866;
  assign n19868 = ~n19852 & ~n19867;
  assign n19869 = ~controllable_hgrant2 & ~n19868;
  assign n19870 = ~n5635 & ~n19869;
  assign n19871 = ~controllable_hmaster0 & ~n19870;
  assign n19872 = ~n19851 & ~n19871;
  assign n19873 = ~controllable_hmaster1 & ~n19872;
  assign n19874 = ~n19850 & ~n19873;
  assign n19875 = ~i_hbusreq3 & ~n19874;
  assign n19876 = ~n19829 & ~n19875;
  assign n19877 = controllable_hmaster2 & ~n19876;
  assign n19878 = ~n4091 & ~n19821;
  assign n19879 = ~controllable_hgrant2 & ~n19878;
  assign n19880 = ~n5616 & ~n19879;
  assign n19881 = controllable_hmaster0 & ~n19880;
  assign n19882 = ~n5686 & ~n19879;
  assign n19883 = ~controllable_hmaster0 & ~n19882;
  assign n19884 = ~n19881 & ~n19883;
  assign n19885 = controllable_hmaster1 & ~n19884;
  assign n19886 = ~i_hlock1 & ~n5961;
  assign n19887 = ~n19814 & ~n19886;
  assign n19888 = ~controllable_ndecide & ~n19887;
  assign n19889 = ~n3494 & ~n19888;
  assign n19890 = i_hready & ~n19889;
  assign n19891 = i_hready & ~n19890;
  assign n19892 = ~controllable_hgrant4 & n19891;
  assign n19893 = ~n4091 & ~n19892;
  assign n19894 = ~controllable_hgrant2 & ~n19893;
  assign n19895 = ~n5616 & ~n19894;
  assign n19896 = controllable_hmaster0 & ~n19895;
  assign n19897 = ~controllable_hmaster0 & ~n19880;
  assign n19898 = ~n19896 & ~n19897;
  assign n19899 = ~controllable_hmaster1 & ~n19898;
  assign n19900 = ~n19885 & ~n19899;
  assign n19901 = i_hbusreq3 & ~n19900;
  assign n19902 = i_hbusreq2 & ~n19878;
  assign n19903 = ~n12172 & ~n19865;
  assign n19904 = ~i_hbusreq2 & ~n19903;
  assign n19905 = ~n19902 & ~n19904;
  assign n19906 = ~controllable_hgrant2 & ~n19905;
  assign n19907 = ~n5635 & ~n19906;
  assign n19908 = controllable_hmaster0 & ~n19907;
  assign n19909 = ~n5722 & ~n19906;
  assign n19910 = ~controllable_hmaster0 & ~n19909;
  assign n19911 = ~n19908 & ~n19910;
  assign n19912 = controllable_hmaster1 & ~n19911;
  assign n19913 = i_hbusreq2 & ~n19893;
  assign n19914 = i_hbusreq4 & ~n19891;
  assign n19915 = i_hbusreq0 & ~n19891;
  assign n19916 = i_hbusreq1 & ~n19887;
  assign n19917 = ~n18087 & ~n19916;
  assign n19918 = ~controllable_ndecide & ~n19917;
  assign n19919 = ~n3494 & ~n19918;
  assign n19920 = i_hready & ~n19919;
  assign n19921 = ~n10361 & ~n19920;
  assign n19922 = i_hlock0 & ~n19921;
  assign n19923 = ~n17487 & ~n19916;
  assign n19924 = ~controllable_ndecide & ~n19923;
  assign n19925 = ~n3494 & ~n19924;
  assign n19926 = i_hready & ~n19925;
  assign n19927 = i_hready & ~n19926;
  assign n19928 = ~i_hlock0 & ~n19927;
  assign n19929 = ~n19922 & ~n19928;
  assign n19930 = ~i_hbusreq0 & ~n19929;
  assign n19931 = ~n19915 & ~n19930;
  assign n19932 = ~i_hbusreq4 & ~n19931;
  assign n19933 = ~n19914 & ~n19932;
  assign n19934 = ~controllable_hgrant4 & n19933;
  assign n19935 = ~n12894 & ~n19934;
  assign n19936 = ~i_hbusreq2 & ~n19935;
  assign n19937 = ~n19913 & ~n19936;
  assign n19938 = ~controllable_hgrant2 & ~n19937;
  assign n19939 = ~n7290 & ~n19938;
  assign n19940 = controllable_hmaster0 & ~n19939;
  assign n19941 = ~controllable_hmaster0 & ~n19907;
  assign n19942 = ~n19940 & ~n19941;
  assign n19943 = ~controllable_hmaster1 & ~n19942;
  assign n19944 = ~n19912 & ~n19943;
  assign n19945 = ~i_hbusreq3 & ~n19944;
  assign n19946 = ~n19901 & ~n19945;
  assign n19947 = ~controllable_hmaster2 & ~n19946;
  assign n19948 = ~n19877 & ~n19947;
  assign n19949 = ~controllable_hgrant3 & ~n19948;
  assign n19950 = ~n19274 & ~n19949;
  assign n19951 = controllable_nhgrant0 & ~n19950;
  assign n19952 = ~n19385 & ~n19951;
  assign n19953 = ~n3281 & ~n19952;
  assign n19954 = ~n3281 & ~n19953;
  assign n19955 = n3378 & ~n19954;
  assign n19956 = ~n18574 & ~n19803;
  assign n19957 = i_hready & ~n19956;
  assign n19958 = ~i_hready & ~n19577;
  assign n19959 = ~n19957 & ~n19958;
  assign n19960 = ~controllable_hgrant4 & n19959;
  assign n19961 = ~n4091 & ~n19960;
  assign n19962 = ~controllable_hgrant2 & ~n19961;
  assign n19963 = ~n5616 & ~n19962;
  assign n19964 = controllable_hmaster1 & ~n19963;
  assign n19965 = controllable_hmaster0 & ~n19963;
  assign n19966 = controllable_ndecide & ~n9985;
  assign n19967 = ~n19817 & ~n19966;
  assign n19968 = i_hready & ~n19967;
  assign n19969 = ~i_hready & ~n19702;
  assign n19970 = ~n19968 & ~n19969;
  assign n19971 = ~controllable_hgrant4 & n19970;
  assign n19972 = ~n4015 & ~n19971;
  assign n19973 = ~controllable_hgrant2 & ~n19972;
  assign n19974 = ~n5616 & ~n19973;
  assign n19975 = ~controllable_hmaster0 & ~n19974;
  assign n19976 = ~n19965 & ~n19975;
  assign n19977 = ~controllable_hmaster1 & ~n19976;
  assign n19978 = ~n19964 & ~n19977;
  assign n19979 = i_hbusreq3 & ~n19978;
  assign n19980 = i_hbusreq2 & ~n19961;
  assign n19981 = i_hbusreq4 & ~n19959;
  assign n19982 = i_hbusreq0 & ~n19959;
  assign n19983 = ~n18574 & ~n19835;
  assign n19984 = i_hready & ~n19983;
  assign n19985 = ~i_hready & n19593;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = i_hlock0 & ~n19986;
  assign n19988 = ~n10431 & ~n19833;
  assign n19989 = ~controllable_ndecide & ~n19988;
  assign n19990 = ~n18574 & ~n19989;
  assign n19991 = i_hready & ~n19990;
  assign n19992 = ~n19958 & ~n19991;
  assign n19993 = ~i_hlock0 & ~n19992;
  assign n19994 = ~n19987 & ~n19993;
  assign n19995 = ~i_hbusreq0 & ~n19994;
  assign n19996 = ~n19982 & ~n19995;
  assign n19997 = ~i_hbusreq4 & ~n19996;
  assign n19998 = ~n19981 & ~n19997;
  assign n19999 = ~controllable_hgrant4 & n19998;
  assign n20000 = ~n5863 & ~n19999;
  assign n20001 = ~i_hbusreq2 & ~n20000;
  assign n20002 = ~n19980 & ~n20001;
  assign n20003 = ~controllable_hgrant2 & ~n20002;
  assign n20004 = ~n5862 & ~n20003;
  assign n20005 = controllable_hmaster1 & ~n20004;
  assign n20006 = controllable_hmaster0 & ~n20004;
  assign n20007 = i_hbusreq2 & ~n19972;
  assign n20008 = i_hbusreq4 & ~n19970;
  assign n20009 = i_hbusreq0 & ~n19970;
  assign n20010 = ~n19857 & ~n19966;
  assign n20011 = i_hready & ~n20010;
  assign n20012 = ~i_hready & n19717;
  assign n20013 = ~n20011 & ~n20012;
  assign n20014 = i_hlock0 & ~n20013;
  assign n20015 = ~n10157 & ~n19855;
  assign n20016 = ~controllable_ndecide & ~n20015;
  assign n20017 = ~n19966 & ~n20016;
  assign n20018 = i_hready & ~n20017;
  assign n20019 = ~n19969 & ~n20018;
  assign n20020 = ~i_hlock0 & ~n20019;
  assign n20021 = ~n20014 & ~n20020;
  assign n20022 = ~i_hbusreq0 & ~n20021;
  assign n20023 = ~n20009 & ~n20022;
  assign n20024 = ~i_hbusreq4 & ~n20023;
  assign n20025 = ~n20008 & ~n20024;
  assign n20026 = ~controllable_hgrant4 & n20025;
  assign n20027 = ~n4064 & ~n20026;
  assign n20028 = ~i_hbusreq2 & ~n20027;
  assign n20029 = ~n20007 & ~n20028;
  assign n20030 = ~controllable_hgrant2 & ~n20029;
  assign n20031 = ~n5862 & ~n20030;
  assign n20032 = ~controllable_hmaster0 & ~n20031;
  assign n20033 = ~n20006 & ~n20032;
  assign n20034 = ~controllable_hmaster1 & ~n20033;
  assign n20035 = ~n20005 & ~n20034;
  assign n20036 = ~i_hbusreq3 & ~n20035;
  assign n20037 = ~n19979 & ~n20036;
  assign n20038 = controllable_hmaster2 & ~n20037;
  assign n20039 = ~n4091 & ~n19971;
  assign n20040 = ~controllable_hgrant2 & ~n20039;
  assign n20041 = ~n5616 & ~n20040;
  assign n20042 = controllable_hmaster0 & ~n20041;
  assign n20043 = ~n5686 & ~n20040;
  assign n20044 = ~controllable_hmaster0 & ~n20043;
  assign n20045 = ~n20042 & ~n20044;
  assign n20046 = controllable_hmaster1 & ~n20045;
  assign n20047 = ~n19888 & ~n19966;
  assign n20048 = i_hready & ~n20047;
  assign n20049 = i_hready & ~n20048;
  assign n20050 = ~controllable_hgrant4 & n20049;
  assign n20051 = ~n4091 & ~n20050;
  assign n20052 = ~controllable_hgrant2 & ~n20051;
  assign n20053 = ~n5616 & ~n20052;
  assign n20054 = controllable_hmaster0 & ~n20053;
  assign n20055 = ~controllable_hmaster0 & ~n20041;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = ~controllable_hmaster1 & ~n20056;
  assign n20058 = ~n20046 & ~n20057;
  assign n20059 = i_hbusreq3 & ~n20058;
  assign n20060 = i_hbusreq2 & ~n20039;
  assign n20061 = ~n5863 & ~n20026;
  assign n20062 = ~i_hbusreq2 & ~n20061;
  assign n20063 = ~n20060 & ~n20062;
  assign n20064 = ~controllable_hgrant2 & ~n20063;
  assign n20065 = ~n5862 & ~n20064;
  assign n20066 = controllable_hmaster0 & ~n20065;
  assign n20067 = ~n5950 & ~n20064;
  assign n20068 = ~controllable_hmaster0 & ~n20067;
  assign n20069 = ~n20066 & ~n20068;
  assign n20070 = controllable_hmaster1 & ~n20069;
  assign n20071 = i_hbusreq2 & ~n20051;
  assign n20072 = i_hbusreq4 & ~n20049;
  assign n20073 = i_hbusreq0 & ~n20049;
  assign n20074 = ~n19918 & ~n19966;
  assign n20075 = i_hready & ~n20074;
  assign n20076 = ~n10361 & ~n20075;
  assign n20077 = i_hlock0 & ~n20076;
  assign n20078 = ~n5962 & ~n19916;
  assign n20079 = ~controllable_ndecide & ~n20078;
  assign n20080 = ~n19966 & ~n20079;
  assign n20081 = i_hready & ~n20080;
  assign n20082 = i_hready & ~n20081;
  assign n20083 = ~i_hlock0 & ~n20082;
  assign n20084 = ~n20077 & ~n20083;
  assign n20085 = ~i_hbusreq0 & ~n20084;
  assign n20086 = ~n20073 & ~n20085;
  assign n20087 = ~i_hbusreq4 & ~n20086;
  assign n20088 = ~n20072 & ~n20087;
  assign n20089 = ~controllable_hgrant4 & n20088;
  assign n20090 = ~n13012 & ~n20089;
  assign n20091 = ~i_hbusreq2 & ~n20090;
  assign n20092 = ~n20071 & ~n20091;
  assign n20093 = ~controllable_hgrant2 & ~n20092;
  assign n20094 = ~n7507 & ~n20093;
  assign n20095 = controllable_hmaster0 & ~n20094;
  assign n20096 = ~i_hready & n19764;
  assign n20097 = ~n20011 & ~n20096;
  assign n20098 = i_hlock0 & ~n20097;
  assign n20099 = ~n20020 & ~n20098;
  assign n20100 = ~i_hbusreq0 & ~n20099;
  assign n20101 = ~n20009 & ~n20100;
  assign n20102 = ~i_hbusreq4 & ~n20101;
  assign n20103 = ~n20008 & ~n20102;
  assign n20104 = ~controllable_hgrant4 & n20103;
  assign n20105 = ~n5982 & ~n20104;
  assign n20106 = ~i_hbusreq2 & ~n20105;
  assign n20107 = ~n20060 & ~n20106;
  assign n20108 = ~controllable_hgrant2 & ~n20107;
  assign n20109 = ~n5981 & ~n20108;
  assign n20110 = ~controllable_hmaster0 & ~n20109;
  assign n20111 = ~n20095 & ~n20110;
  assign n20112 = ~controllable_hmaster1 & ~n20111;
  assign n20113 = ~n20070 & ~n20112;
  assign n20114 = ~i_hbusreq3 & ~n20113;
  assign n20115 = ~n20059 & ~n20114;
  assign n20116 = ~controllable_hmaster2 & ~n20115;
  assign n20117 = ~n20038 & ~n20116;
  assign n20118 = ~controllable_hgrant3 & ~n20117;
  assign n20119 = ~n19398 & ~n20118;
  assign n20120 = controllable_nhgrant0 & ~n20119;
  assign n20121 = ~n19515 & ~n20120;
  assign n20122 = ~n3281 & ~n20121;
  assign n20123 = ~n3281 & ~n20122;
  assign n20124 = ~n3378 & ~n20123;
  assign n20125 = ~n19955 & ~n20124;
  assign n20126 = n3492 & ~n20125;
  assign n20127 = ~n18151 & ~n20126;
  assign n20128 = n3485 & ~n20127;
  assign n20129 = ~n18150 & ~n20128;
  assign n20130 = n3476 & ~n20129;
  assign n20131 = ~n19799 & ~n20130;
  assign n20132 = n3374 & ~n20131;
  assign n20133 = ~n19630 & ~n20132;
  assign n20134 = ~n3655 & ~n20133;
  assign n20135 = ~n19529 & ~n20134;
  assign n20136 = n3652 & ~n20135;
  assign n20137 = ~n3821 & ~n10774;
  assign n20138 = ~controllable_hmaster1 & ~n20137;
  assign n20139 = ~n5293 & ~n20138;
  assign n20140 = i_hbusreq3 & ~n20139;
  assign n20141 = ~n5278 & ~n10788;
  assign n20142 = ~controllable_hmaster1 & ~n20141;
  assign n20143 = ~n5313 & ~n20142;
  assign n20144 = ~i_hbusreq3 & ~n20143;
  assign n20145 = ~n20140 & ~n20144;
  assign n20146 = ~controllable_hmaster2 & ~n20145;
  assign n20147 = ~n12741 & ~n20146;
  assign n20148 = ~controllable_hgrant3 & ~n20147;
  assign n20149 = ~n19183 & ~n20148;
  assign n20150 = controllable_nhgrant0 & ~n20149;
  assign n20151 = ~n19213 & ~n20150;
  assign n20152 = ~n3281 & ~n20151;
  assign n20153 = ~n3281 & ~n20152;
  assign n20154 = n3378 & ~n20153;
  assign n20155 = ~n6704 & ~n10774;
  assign n20156 = ~controllable_hmaster1 & ~n20155;
  assign n20157 = ~n6701 & ~n20156;
  assign n20158 = i_hbusreq3 & ~n20157;
  assign n20159 = ~n6717 & ~n10788;
  assign n20160 = ~controllable_hmaster1 & ~n20159;
  assign n20161 = ~n6714 & ~n20160;
  assign n20162 = ~i_hbusreq3 & ~n20161;
  assign n20163 = ~n20158 & ~n20162;
  assign n20164 = ~controllable_hmaster2 & ~n20163;
  assign n20165 = ~n13276 & ~n20164;
  assign n20166 = ~controllable_hgrant3 & ~n20165;
  assign n20167 = ~n19225 & ~n20166;
  assign n20168 = controllable_nhgrant0 & ~n20167;
  assign n20169 = ~n19255 & ~n20168;
  assign n20170 = ~n3281 & ~n20169;
  assign n20171 = ~n3281 & ~n20170;
  assign n20172 = ~n3378 & ~n20171;
  assign n20173 = ~n20154 & ~n20172;
  assign n20174 = n3492 & ~n20173;
  assign n20175 = n3492 & ~n20174;
  assign n20176 = n3485 & ~n20175;
  assign n20177 = n3485 & ~n20176;
  assign n20178 = ~n3476 & ~n20177;
  assign n20179 = ~n8029 & ~n19317;
  assign n20180 = controllable_hmaster0 & ~n20179;
  assign n20181 = ~n7340 & ~n20180;
  assign n20182 = ~controllable_hmaster1 & ~n20181;
  assign n20183 = ~n7330 & ~n20182;
  assign n20184 = i_hbusreq3 & ~n20183;
  assign n20185 = ~n8036 & ~n19358;
  assign n20186 = controllable_hmaster0 & ~n20185;
  assign n20187 = ~n19361 & ~n20186;
  assign n20188 = ~controllable_hmaster1 & ~n20187;
  assign n20189 = ~n19333 & ~n20188;
  assign n20190 = ~i_hbusreq3 & ~n20189;
  assign n20191 = ~n20184 & ~n20190;
  assign n20192 = ~controllable_hmaster2 & ~n20191;
  assign n20193 = ~n19313 & ~n20192;
  assign n20194 = ~controllable_hgrant3 & ~n20193;
  assign n20195 = ~n19274 & ~n20194;
  assign n20196 = controllable_nhgrant0 & ~n20195;
  assign n20197 = ~n19385 & ~n20196;
  assign n20198 = ~n3281 & ~n20197;
  assign n20199 = ~n3281 & ~n20198;
  assign n20200 = n3378 & ~n20199;
  assign n20201 = ~n6772 & ~n19412;
  assign n20202 = controllable_hmaster1 & ~n20201;
  assign n20203 = controllable_hmaster0 & ~n20201;
  assign n20204 = ~n6772 & ~n19429;
  assign n20205 = ~controllable_hmaster0 & ~n20204;
  assign n20206 = ~n20203 & ~n20205;
  assign n20207 = ~controllable_hmaster1 & ~n20206;
  assign n20208 = ~n20202 & ~n20207;
  assign n20209 = ~i_hbusreq3 & ~n20208;
  assign n20210 = ~n13328 & ~n20209;
  assign n20211 = controllable_hmaster2 & ~n20210;
  assign n20212 = ~n8056 & ~n19441;
  assign n20213 = controllable_hmaster0 & ~n20212;
  assign n20214 = ~n8083 & ~n20213;
  assign n20215 = ~controllable_hmaster1 & ~n20214;
  assign n20216 = ~n8080 & ~n20215;
  assign n20217 = i_hbusreq3 & ~n20216;
  assign n20218 = ~n6772 & ~n19451;
  assign n20219 = controllable_hmaster0 & ~n20218;
  assign n20220 = ~n6813 & ~n19451;
  assign n20221 = ~controllable_hmaster0 & ~n20220;
  assign n20222 = ~n20219 & ~n20221;
  assign n20223 = controllable_hmaster1 & ~n20222;
  assign n20224 = ~n8066 & ~n19475;
  assign n20225 = controllable_hmaster0 & ~n20224;
  assign n20226 = ~n6831 & ~n19489;
  assign n20227 = ~controllable_hmaster0 & ~n20226;
  assign n20228 = ~n20225 & ~n20227;
  assign n20229 = ~controllable_hmaster1 & ~n20228;
  assign n20230 = ~n20223 & ~n20229;
  assign n20231 = ~i_hbusreq3 & ~n20230;
  assign n20232 = ~n20217 & ~n20231;
  assign n20233 = ~controllable_hmaster2 & ~n20232;
  assign n20234 = ~n20211 & ~n20233;
  assign n20235 = ~controllable_hgrant3 & ~n20234;
  assign n20236 = ~n19398 & ~n20235;
  assign n20237 = controllable_nhgrant0 & ~n20236;
  assign n20238 = ~n19515 & ~n20237;
  assign n20239 = ~n3281 & ~n20238;
  assign n20240 = ~n3281 & ~n20239;
  assign n20241 = ~n3378 & ~n20240;
  assign n20242 = ~n20200 & ~n20241;
  assign n20243 = n3492 & ~n20242;
  assign n20244 = n3492 & ~n20243;
  assign n20245 = n3485 & ~n20244;
  assign n20246 = n3485 & ~n20245;
  assign n20247 = n3476 & ~n20246;
  assign n20248 = ~n20178 & ~n20247;
  assign n20249 = n3374 & ~n20248;
  assign n20250 = ~n7986 & ~n20249;
  assign n20251 = n3655 & ~n20250;
  assign n20252 = ~n4333 & ~n19582;
  assign n20253 = controllable_hmaster1 & ~n20252;
  assign n20254 = controllable_hmaster0 & ~n20252;
  assign n20255 = controllable_hmaster0 & ~n20254;
  assign n20256 = ~controllable_hmaster1 & ~n20255;
  assign n20257 = ~n20253 & ~n20256;
  assign n20258 = i_hbusreq3 & ~n20257;
  assign n20259 = ~n4340 & ~n19607;
  assign n20260 = controllable_hmaster1 & ~n20259;
  assign n20261 = controllable_hmaster0 & ~n20259;
  assign n20262 = controllable_hmaster0 & ~n20261;
  assign n20263 = ~controllable_hmaster1 & ~n20262;
  assign n20264 = ~n20260 & ~n20263;
  assign n20265 = ~i_hbusreq3 & ~n20264;
  assign n20266 = ~n20258 & ~n20265;
  assign n20267 = controllable_hmaster2 & ~n20266;
  assign n20268 = controllable_hmaster2 & ~n20267;
  assign n20269 = ~controllable_hgrant3 & ~n20268;
  assign n20270 = ~n7090 & ~n20269;
  assign n20271 = controllable_nhgrant0 & ~n20270;
  assign n20272 = ~n7118 & ~n20271;
  assign n20273 = ~n3281 & ~n20272;
  assign n20274 = ~n3281 & ~n20273;
  assign n20275 = ~n3378 & ~n20274;
  assign n20276 = ~n19575 & ~n20275;
  assign n20277 = n3492 & ~n20276;
  assign n20278 = n3492 & ~n20277;
  assign n20279 = n3485 & ~n20278;
  assign n20280 = n3485 & ~n20279;
  assign n20281 = ~n3374 & ~n20280;
  assign n20282 = ~n11209 & ~n19670;
  assign n20283 = ~controllable_hmaster1 & ~n20282;
  assign n20284 = ~n19669 & ~n20283;
  assign n20285 = i_hbusreq3 & ~n20284;
  assign n20286 = ~n11222 & ~n19686;
  assign n20287 = ~controllable_hmaster1 & ~n20286;
  assign n20288 = ~n19685 & ~n20287;
  assign n20289 = ~i_hbusreq3 & ~n20288;
  assign n20290 = ~n20285 & ~n20289;
  assign n20291 = ~controllable_hmaster2 & ~n20290;
  assign n20292 = ~n19661 & ~n20291;
  assign n20293 = ~controllable_hgrant3 & ~n20292;
  assign n20294 = ~n19183 & ~n20293;
  assign n20295 = controllable_nhgrant0 & ~n20294;
  assign n20296 = ~n19213 & ~n20295;
  assign n20297 = ~n3281 & ~n20296;
  assign n20298 = ~n3281 & ~n20297;
  assign n20299 = n3378 & ~n20298;
  assign n20300 = ~n4333 & ~n19707;
  assign n20301 = ~controllable_hmaster0 & ~n20300;
  assign n20302 = ~n20254 & ~n20301;
  assign n20303 = ~controllable_hmaster1 & ~n20302;
  assign n20304 = ~n20253 & ~n20303;
  assign n20305 = i_hbusreq3 & ~n20304;
  assign n20306 = ~n4340 & ~n19731;
  assign n20307 = ~controllable_hmaster0 & ~n20306;
  assign n20308 = ~n20261 & ~n20307;
  assign n20309 = ~controllable_hmaster1 & ~n20308;
  assign n20310 = ~n20260 & ~n20309;
  assign n20311 = ~i_hbusreq3 & ~n20310;
  assign n20312 = ~n20305 & ~n20311;
  assign n20313 = controllable_hmaster2 & ~n20312;
  assign n20314 = ~n4333 & ~n19741;
  assign n20315 = controllable_hmaster0 & ~n20314;
  assign n20316 = ~n6697 & ~n19741;
  assign n20317 = ~controllable_hmaster0 & ~n20316;
  assign n20318 = ~n20315 & ~n20317;
  assign n20319 = controllable_hmaster1 & ~n20318;
  assign n20320 = ~controllable_hmaster0 & ~n20314;
  assign n20321 = ~n11209 & ~n20320;
  assign n20322 = ~controllable_hmaster1 & ~n20321;
  assign n20323 = ~n20319 & ~n20322;
  assign n20324 = i_hbusreq3 & ~n20323;
  assign n20325 = ~n4340 & ~n19757;
  assign n20326 = controllable_hmaster0 & ~n20325;
  assign n20327 = ~n6710 & ~n19757;
  assign n20328 = ~controllable_hmaster0 & ~n20327;
  assign n20329 = ~n20326 & ~n20328;
  assign n20330 = controllable_hmaster1 & ~n20329;
  assign n20331 = ~n6947 & ~n19777;
  assign n20332 = ~controllable_hmaster0 & ~n20331;
  assign n20333 = ~n11222 & ~n20332;
  assign n20334 = ~controllable_hmaster1 & ~n20333;
  assign n20335 = ~n20330 & ~n20334;
  assign n20336 = ~i_hbusreq3 & ~n20335;
  assign n20337 = ~n20324 & ~n20336;
  assign n20338 = ~controllable_hmaster2 & ~n20337;
  assign n20339 = ~n20313 & ~n20338;
  assign n20340 = ~controllable_hgrant3 & ~n20339;
  assign n20341 = ~n19225 & ~n20340;
  assign n20342 = controllable_nhgrant0 & ~n20341;
  assign n20343 = ~n19255 & ~n20342;
  assign n20344 = ~n3281 & ~n20343;
  assign n20345 = ~n3281 & ~n20344;
  assign n20346 = ~n3378 & ~n20345;
  assign n20347 = ~n20299 & ~n20346;
  assign n20348 = n3492 & ~n20347;
  assign n20349 = n3492 & ~n20348;
  assign n20350 = n3485 & ~n20349;
  assign n20351 = n3485 & ~n20350;
  assign n20352 = ~n3476 & ~n20351;
  assign n20353 = ~n8029 & ~n19894;
  assign n20354 = controllable_hmaster0 & ~n20353;
  assign n20355 = ~n19897 & ~n20354;
  assign n20356 = ~controllable_hmaster1 & ~n20355;
  assign n20357 = ~n19885 & ~n20356;
  assign n20358 = i_hbusreq3 & ~n20357;
  assign n20359 = ~n8036 & ~n19938;
  assign n20360 = controllable_hmaster0 & ~n20359;
  assign n20361 = ~n19941 & ~n20360;
  assign n20362 = ~controllable_hmaster1 & ~n20361;
  assign n20363 = ~n19912 & ~n20362;
  assign n20364 = ~i_hbusreq3 & ~n20363;
  assign n20365 = ~n20358 & ~n20364;
  assign n20366 = ~controllable_hmaster2 & ~n20365;
  assign n20367 = ~n19877 & ~n20366;
  assign n20368 = ~controllable_hgrant3 & ~n20367;
  assign n20369 = ~n19274 & ~n20368;
  assign n20370 = controllable_nhgrant0 & ~n20369;
  assign n20371 = ~n19385 & ~n20370;
  assign n20372 = ~n3281 & ~n20371;
  assign n20373 = ~n3281 & ~n20372;
  assign n20374 = n3378 & ~n20373;
  assign n20375 = ~n6762 & ~n19962;
  assign n20376 = controllable_hmaster1 & ~n20375;
  assign n20377 = controllable_hmaster0 & ~n20375;
  assign n20378 = ~n6762 & ~n19973;
  assign n20379 = ~controllable_hmaster0 & ~n20378;
  assign n20380 = ~n20377 & ~n20379;
  assign n20381 = ~controllable_hmaster1 & ~n20380;
  assign n20382 = ~n20376 & ~n20381;
  assign n20383 = i_hbusreq3 & ~n20382;
  assign n20384 = ~n6772 & ~n20003;
  assign n20385 = controllable_hmaster1 & ~n20384;
  assign n20386 = controllable_hmaster0 & ~n20384;
  assign n20387 = ~n6772 & ~n20030;
  assign n20388 = ~controllable_hmaster0 & ~n20387;
  assign n20389 = ~n20386 & ~n20388;
  assign n20390 = ~controllable_hmaster1 & ~n20389;
  assign n20391 = ~n20385 & ~n20390;
  assign n20392 = ~i_hbusreq3 & ~n20391;
  assign n20393 = ~n20383 & ~n20392;
  assign n20394 = controllable_hmaster2 & ~n20393;
  assign n20395 = ~n6762 & ~n20040;
  assign n20396 = controllable_hmaster0 & ~n20395;
  assign n20397 = ~n6786 & ~n20040;
  assign n20398 = ~controllable_hmaster0 & ~n20397;
  assign n20399 = ~n20396 & ~n20398;
  assign n20400 = controllable_hmaster1 & ~n20399;
  assign n20401 = ~n8056 & ~n20052;
  assign n20402 = controllable_hmaster0 & ~n20401;
  assign n20403 = ~controllable_hmaster0 & ~n20395;
  assign n20404 = ~n20402 & ~n20403;
  assign n20405 = ~controllable_hmaster1 & ~n20404;
  assign n20406 = ~n20400 & ~n20405;
  assign n20407 = i_hbusreq3 & ~n20406;
  assign n20408 = ~n6772 & ~n20064;
  assign n20409 = controllable_hmaster0 & ~n20408;
  assign n20410 = ~n6813 & ~n20064;
  assign n20411 = ~controllable_hmaster0 & ~n20410;
  assign n20412 = ~n20409 & ~n20411;
  assign n20413 = controllable_hmaster1 & ~n20412;
  assign n20414 = ~n8066 & ~n20093;
  assign n20415 = controllable_hmaster0 & ~n20414;
  assign n20416 = ~n6831 & ~n20108;
  assign n20417 = ~controllable_hmaster0 & ~n20416;
  assign n20418 = ~n20415 & ~n20417;
  assign n20419 = ~controllable_hmaster1 & ~n20418;
  assign n20420 = ~n20413 & ~n20419;
  assign n20421 = ~i_hbusreq3 & ~n20420;
  assign n20422 = ~n20407 & ~n20421;
  assign n20423 = ~controllable_hmaster2 & ~n20422;
  assign n20424 = ~n20394 & ~n20423;
  assign n20425 = ~controllable_hgrant3 & ~n20424;
  assign n20426 = ~n19398 & ~n20425;
  assign n20427 = controllable_nhgrant0 & ~n20426;
  assign n20428 = ~n19515 & ~n20427;
  assign n20429 = ~n3281 & ~n20428;
  assign n20430 = ~n3281 & ~n20429;
  assign n20431 = ~n3378 & ~n20430;
  assign n20432 = ~n20374 & ~n20431;
  assign n20433 = n3492 & ~n20432;
  assign n20434 = ~n18151 & ~n20433;
  assign n20435 = n3485 & ~n20434;
  assign n20436 = ~n18150 & ~n20435;
  assign n20437 = n3476 & ~n20436;
  assign n20438 = ~n20352 & ~n20437;
  assign n20439 = n3374 & ~n20438;
  assign n20440 = ~n20281 & ~n20439;
  assign n20441 = ~n3655 & ~n20440;
  assign n20442 = ~n20251 & ~n20441;
  assign n20443 = ~n3652 & ~n20442;
  assign n20444 = ~n20136 & ~n20443;
  assign n20445 = n3368 & ~n20444;
  assign n20446 = ~n19176 & ~n20445;
  assign n20447 = n3362 & ~n20446;
  assign n20448 = n3492 & ~n18437;
  assign n20449 = ~n3631 & ~n20448;
  assign n20450 = n3485 & ~n20449;
  assign n20451 = ~n3630 & ~n20450;
  assign n20452 = ~n3476 & ~n20451;
  assign n20453 = n3492 & ~n18559;
  assign n20454 = ~n3631 & ~n20453;
  assign n20455 = n3485 & ~n20454;
  assign n20456 = ~n8312 & ~n20455;
  assign n20457 = n3476 & ~n20456;
  assign n20458 = ~n20452 & ~n20457;
  assign n20459 = n3374 & ~n20458;
  assign n20460 = ~n8316 & ~n20459;
  assign n20461 = n3655 & ~n20460;
  assign n20462 = n3492 & ~n18621;
  assign n20463 = ~n3631 & ~n20462;
  assign n20464 = n3485 & ~n20463;
  assign n20465 = ~n3630 & ~n20464;
  assign n20466 = ~n3476 & ~n20465;
  assign n20467 = n3492 & ~n17608;
  assign n20468 = ~n8367 & ~n20467;
  assign n20469 = ~n3485 & ~n20468;
  assign n20470 = ~n18630 & ~n20462;
  assign n20471 = n3485 & ~n20470;
  assign n20472 = ~n20469 & ~n20471;
  assign n20473 = n3476 & ~n20472;
  assign n20474 = ~n20466 & ~n20473;
  assign n20475 = ~n3374 & ~n20474;
  assign n20476 = n3492 & ~n18751;
  assign n20477 = ~n3631 & ~n20476;
  assign n20478 = n3485 & ~n20477;
  assign n20479 = ~n3630 & ~n20478;
  assign n20480 = ~n3476 & ~n20479;
  assign n20481 = n3492 & ~n18897;
  assign n20482 = ~n18630 & ~n20481;
  assign n20483 = n3485 & ~n20482;
  assign n20484 = ~n20469 & ~n20483;
  assign n20485 = n3476 & ~n20484;
  assign n20486 = ~n20480 & ~n20485;
  assign n20487 = n3374 & ~n20486;
  assign n20488 = ~n20475 & ~n20487;
  assign n20489 = ~n3655 & ~n20488;
  assign n20490 = ~n20461 & ~n20489;
  assign n20491 = n3652 & ~n20490;
  assign n20492 = n3492 & ~n18951;
  assign n20493 = ~n3631 & ~n20492;
  assign n20494 = n3485 & ~n20493;
  assign n20495 = ~n3630 & ~n20494;
  assign n20496 = ~n3476 & ~n20495;
  assign n20497 = n3492 & ~n18999;
  assign n20498 = ~n3631 & ~n20497;
  assign n20499 = n3485 & ~n20498;
  assign n20500 = ~n8436 & ~n20499;
  assign n20501 = n3476 & ~n20500;
  assign n20502 = ~n20496 & ~n20501;
  assign n20503 = n3374 & ~n20502;
  assign n20504 = ~n8440 & ~n20503;
  assign n20505 = n3655 & ~n20504;
  assign n20506 = n3492 & ~n19033;
  assign n20507 = ~n3631 & ~n20506;
  assign n20508 = n3485 & ~n20507;
  assign n20509 = ~n3630 & ~n20508;
  assign n20510 = ~n3476 & ~n20509;
  assign n20511 = ~n8491 & ~n20467;
  assign n20512 = ~n3485 & ~n20511;
  assign n20513 = ~n18630 & ~n20506;
  assign n20514 = n3485 & ~n20513;
  assign n20515 = ~n20512 & ~n20514;
  assign n20516 = n3476 & ~n20515;
  assign n20517 = ~n20510 & ~n20516;
  assign n20518 = ~n3374 & ~n20517;
  assign n20519 = n3492 & ~n19097;
  assign n20520 = ~n3631 & ~n20519;
  assign n20521 = n3485 & ~n20520;
  assign n20522 = ~n3630 & ~n20521;
  assign n20523 = ~n3476 & ~n20522;
  assign n20524 = n3492 & ~n19161;
  assign n20525 = ~n18630 & ~n20524;
  assign n20526 = n3485 & ~n20525;
  assign n20527 = ~n20512 & ~n20526;
  assign n20528 = n3476 & ~n20527;
  assign n20529 = ~n20523 & ~n20528;
  assign n20530 = n3374 & ~n20529;
  assign n20531 = ~n20518 & ~n20530;
  assign n20532 = ~n3655 & ~n20531;
  assign n20533 = ~n20505 & ~n20532;
  assign n20534 = ~n3652 & ~n20533;
  assign n20535 = ~n20491 & ~n20534;
  assign n20536 = ~n3368 & ~n20535;
  assign n20537 = n3492 & ~n19258;
  assign n20538 = n3492 & ~n20537;
  assign n20539 = n3485 & ~n20538;
  assign n20540 = n3485 & ~n20539;
  assign n20541 = ~n3476 & ~n20540;
  assign n20542 = n3492 & ~n19518;
  assign n20543 = n3492 & ~n20542;
  assign n20544 = n3485 & ~n20543;
  assign n20545 = ~n8538 & ~n20544;
  assign n20546 = n3476 & ~n20545;
  assign n20547 = ~n20541 & ~n20546;
  assign n20548 = n3374 & ~n20547;
  assign n20549 = ~n8529 & ~n20548;
  assign n20550 = n3655 & ~n20549;
  assign n20551 = n3492 & ~n19623;
  assign n20552 = n3492 & ~n20551;
  assign n20553 = n3485 & ~n20552;
  assign n20554 = n3485 & ~n20553;
  assign n20555 = ~n3476 & ~n20554;
  assign n20556 = ~n8525 & ~n20553;
  assign n20557 = n3476 & ~n20556;
  assign n20558 = ~n20555 & ~n20557;
  assign n20559 = ~n3374 & ~n20558;
  assign n20560 = n3492 & ~n19792;
  assign n20561 = n3492 & ~n20560;
  assign n20562 = n3485 & ~n20561;
  assign n20563 = n3485 & ~n20562;
  assign n20564 = ~n3476 & ~n20563;
  assign n20565 = n3492 & ~n17546;
  assign n20566 = ~n8563 & ~n20565;
  assign n20567 = ~n3485 & ~n20566;
  assign n20568 = n3492 & ~n20123;
  assign n20569 = ~n18151 & ~n20568;
  assign n20570 = n3485 & ~n20569;
  assign n20571 = ~n20567 & ~n20570;
  assign n20572 = n3476 & ~n20571;
  assign n20573 = ~n20564 & ~n20572;
  assign n20574 = n3374 & ~n20573;
  assign n20575 = ~n20559 & ~n20574;
  assign n20576 = ~n3655 & ~n20575;
  assign n20577 = ~n20550 & ~n20576;
  assign n20578 = n3652 & ~n20577;
  assign n20579 = n3492 & ~n20171;
  assign n20580 = n3492 & ~n20579;
  assign n20581 = n3485 & ~n20580;
  assign n20582 = n3485 & ~n20581;
  assign n20583 = ~n3476 & ~n20582;
  assign n20584 = n3492 & ~n20240;
  assign n20585 = n3492 & ~n20584;
  assign n20586 = n3485 & ~n20585;
  assign n20587 = ~n8594 & ~n20586;
  assign n20588 = n3476 & ~n20587;
  assign n20589 = ~n20583 & ~n20588;
  assign n20590 = n3374 & ~n20589;
  assign n20591 = ~n8585 & ~n20590;
  assign n20592 = n3655 & ~n20591;
  assign n20593 = n3492 & ~n20274;
  assign n20594 = n3492 & ~n20593;
  assign n20595 = n3485 & ~n20594;
  assign n20596 = n3485 & ~n20595;
  assign n20597 = ~n3476 & ~n20596;
  assign n20598 = ~n8525 & ~n20595;
  assign n20599 = n3476 & ~n20598;
  assign n20600 = ~n20597 & ~n20599;
  assign n20601 = ~n3374 & ~n20600;
  assign n20602 = n3492 & ~n20345;
  assign n20603 = n3492 & ~n20602;
  assign n20604 = n3485 & ~n20603;
  assign n20605 = n3485 & ~n20604;
  assign n20606 = ~n3476 & ~n20605;
  assign n20607 = ~n8619 & ~n20565;
  assign n20608 = ~n3485 & ~n20607;
  assign n20609 = n3492 & ~n20430;
  assign n20610 = ~n18151 & ~n20609;
  assign n20611 = n3485 & ~n20610;
  assign n20612 = ~n20608 & ~n20611;
  assign n20613 = n3476 & ~n20612;
  assign n20614 = ~n20606 & ~n20613;
  assign n20615 = n3374 & ~n20614;
  assign n20616 = ~n20601 & ~n20615;
  assign n20617 = ~n3655 & ~n20616;
  assign n20618 = ~n20592 & ~n20617;
  assign n20619 = ~n3652 & ~n20618;
  assign n20620 = ~n20578 & ~n20619;
  assign n20621 = n3368 & ~n20620;
  assign n20622 = ~n20536 & ~n20621;
  assign n20623 = ~n3362 & ~n20622;
  assign n20624 = ~n20447 & ~n20623;
  assign n20625 = n3359 & ~n20624;
  assign n20626 = ~n8639 & ~n20455;
  assign n20627 = n3476 & ~n20626;
  assign n20628 = ~n20452 & ~n20627;
  assign n20629 = n3374 & ~n20628;
  assign n20630 = ~n8643 & ~n20629;
  assign n20631 = n3655 & ~n20630;
  assign n20632 = ~n8650 & ~n20471;
  assign n20633 = n3476 & ~n20632;
  assign n20634 = ~n20466 & ~n20633;
  assign n20635 = ~n3374 & ~n20634;
  assign n20636 = ~n8650 & ~n20483;
  assign n20637 = n3476 & ~n20636;
  assign n20638 = ~n20480 & ~n20637;
  assign n20639 = n3374 & ~n20638;
  assign n20640 = ~n20635 & ~n20639;
  assign n20641 = ~n3655 & ~n20640;
  assign n20642 = ~n20631 & ~n20641;
  assign n20643 = n3652 & ~n20642;
  assign n20644 = ~n8663 & ~n20499;
  assign n20645 = n3476 & ~n20644;
  assign n20646 = ~n20496 & ~n20645;
  assign n20647 = n3374 & ~n20646;
  assign n20648 = ~n8667 & ~n20647;
  assign n20649 = n3655 & ~n20648;
  assign n20650 = ~n8674 & ~n20514;
  assign n20651 = n3476 & ~n20650;
  assign n20652 = ~n20510 & ~n20651;
  assign n20653 = ~n3374 & ~n20652;
  assign n20654 = ~n8674 & ~n20526;
  assign n20655 = n3476 & ~n20654;
  assign n20656 = ~n20523 & ~n20655;
  assign n20657 = n3374 & ~n20656;
  assign n20658 = ~n20653 & ~n20657;
  assign n20659 = ~n3655 & ~n20658;
  assign n20660 = ~n20649 & ~n20659;
  assign n20661 = ~n3652 & ~n20660;
  assign n20662 = ~n20643 & ~n20661;
  assign n20663 = ~n3368 & ~n20662;
  assign n20664 = ~n8694 & ~n20544;
  assign n20665 = n3476 & ~n20664;
  assign n20666 = ~n20541 & ~n20665;
  assign n20667 = n3374 & ~n20666;
  assign n20668 = ~n8693 & ~n20667;
  assign n20669 = n3655 & ~n20668;
  assign n20670 = ~n8689 & ~n20553;
  assign n20671 = n3476 & ~n20670;
  assign n20672 = ~n20555 & ~n20671;
  assign n20673 = ~n3374 & ~n20672;
  assign n20674 = ~n8705 & ~n20570;
  assign n20675 = n3476 & ~n20674;
  assign n20676 = ~n20564 & ~n20675;
  assign n20677 = n3374 & ~n20676;
  assign n20678 = ~n20673 & ~n20677;
  assign n20679 = ~n3655 & ~n20678;
  assign n20680 = ~n20669 & ~n20679;
  assign n20681 = n3652 & ~n20680;
  assign n20682 = ~n8718 & ~n20586;
  assign n20683 = n3476 & ~n20682;
  assign n20684 = ~n20583 & ~n20683;
  assign n20685 = n3374 & ~n20684;
  assign n20686 = ~n8717 & ~n20685;
  assign n20687 = n3655 & ~n20686;
  assign n20688 = ~n8689 & ~n20595;
  assign n20689 = n3476 & ~n20688;
  assign n20690 = ~n20597 & ~n20689;
  assign n20691 = ~n3374 & ~n20690;
  assign n20692 = ~n8729 & ~n20611;
  assign n20693 = n3476 & ~n20692;
  assign n20694 = ~n20606 & ~n20693;
  assign n20695 = n3374 & ~n20694;
  assign n20696 = ~n20691 & ~n20695;
  assign n20697 = ~n3655 & ~n20696;
  assign n20698 = ~n20687 & ~n20697;
  assign n20699 = ~n3652 & ~n20698;
  assign n20700 = ~n20681 & ~n20699;
  assign n20701 = n3368 & ~n20700;
  assign n20702 = ~n20663 & ~n20701;
  assign n20703 = n3362 & ~n20702;
  assign n20704 = n3378 & ~n18437;
  assign n20705 = ~n8906 & ~n20704;
  assign n20706 = n3492 & ~n20705;
  assign n20707 = ~n3631 & ~n20706;
  assign n20708 = n3485 & ~n20707;
  assign n20709 = ~n3630 & ~n20708;
  assign n20710 = ~n3476 & ~n20709;
  assign n20711 = n3378 & ~n18559;
  assign n20712 = ~n9100 & ~n20711;
  assign n20713 = n3492 & ~n20712;
  assign n20714 = ~n8309 & ~n20713;
  assign n20715 = n3485 & ~n20714;
  assign n20716 = ~n8639 & ~n20715;
  assign n20717 = n3476 & ~n20716;
  assign n20718 = ~n20710 & ~n20717;
  assign n20719 = n3374 & ~n20718;
  assign n20720 = ~n8801 & ~n20719;
  assign n20721 = n3655 & ~n20720;
  assign n20722 = n3378 & ~n18621;
  assign n20723 = ~n9135 & ~n20722;
  assign n20724 = n3492 & ~n20723;
  assign n20725 = ~n3631 & ~n20724;
  assign n20726 = n3485 & ~n20725;
  assign n20727 = ~n3630 & ~n20726;
  assign n20728 = ~n3476 & ~n20727;
  assign n20729 = ~n8367 & ~n20724;
  assign n20730 = n3485 & ~n20729;
  assign n20731 = ~n8650 & ~n20730;
  assign n20732 = n3476 & ~n20731;
  assign n20733 = ~n20728 & ~n20732;
  assign n20734 = ~n3374 & ~n20733;
  assign n20735 = n3378 & ~n18751;
  assign n20736 = ~n9240 & ~n20735;
  assign n20737 = n3492 & ~n20736;
  assign n20738 = ~n3631 & ~n20737;
  assign n20739 = n3485 & ~n20738;
  assign n20740 = ~n3630 & ~n20739;
  assign n20741 = ~n3476 & ~n20740;
  assign n20742 = n3378 & ~n18897;
  assign n20743 = ~n9374 & ~n20742;
  assign n20744 = n3492 & ~n20743;
  assign n20745 = ~n8367 & ~n20744;
  assign n20746 = n3485 & ~n20745;
  assign n20747 = ~n8650 & ~n20746;
  assign n20748 = n3476 & ~n20747;
  assign n20749 = ~n20741 & ~n20748;
  assign n20750 = n3374 & ~n20749;
  assign n20751 = ~n20734 & ~n20750;
  assign n20752 = ~n3655 & ~n20751;
  assign n20753 = ~n20721 & ~n20752;
  assign n20754 = n3652 & ~n20753;
  assign n20755 = n3378 & ~n18951;
  assign n20756 = ~n9469 & ~n20755;
  assign n20757 = n3492 & ~n20756;
  assign n20758 = ~n3631 & ~n20757;
  assign n20759 = n3485 & ~n20758;
  assign n20760 = ~n3630 & ~n20759;
  assign n20761 = ~n3476 & ~n20760;
  assign n20762 = n3378 & ~n18999;
  assign n20763 = ~n9531 & ~n20762;
  assign n20764 = n3492 & ~n20763;
  assign n20765 = ~n8434 & ~n20764;
  assign n20766 = n3485 & ~n20765;
  assign n20767 = ~n8663 & ~n20766;
  assign n20768 = n3476 & ~n20767;
  assign n20769 = ~n20761 & ~n20768;
  assign n20770 = n3374 & ~n20769;
  assign n20771 = ~n9421 & ~n20770;
  assign n20772 = n3655 & ~n20771;
  assign n20773 = n3378 & ~n19033;
  assign n20774 = ~n9563 & ~n20773;
  assign n20775 = n3492 & ~n20774;
  assign n20776 = ~n3631 & ~n20775;
  assign n20777 = n3485 & ~n20776;
  assign n20778 = ~n3630 & ~n20777;
  assign n20779 = ~n3476 & ~n20778;
  assign n20780 = ~n8491 & ~n20775;
  assign n20781 = n3485 & ~n20780;
  assign n20782 = ~n8674 & ~n20781;
  assign n20783 = n3476 & ~n20782;
  assign n20784 = ~n20779 & ~n20783;
  assign n20785 = ~n3374 & ~n20784;
  assign n20786 = n3378 & ~n19097;
  assign n20787 = ~n9623 & ~n20786;
  assign n20788 = n3492 & ~n20787;
  assign n20789 = ~n3631 & ~n20788;
  assign n20790 = n3485 & ~n20789;
  assign n20791 = ~n3630 & ~n20790;
  assign n20792 = ~n3476 & ~n20791;
  assign n20793 = n3378 & ~n19161;
  assign n20794 = ~n9683 & ~n20793;
  assign n20795 = n3492 & ~n20794;
  assign n20796 = ~n8491 & ~n20795;
  assign n20797 = n3485 & ~n20796;
  assign n20798 = ~n8674 & ~n20797;
  assign n20799 = n3476 & ~n20798;
  assign n20800 = ~n20792 & ~n20799;
  assign n20801 = n3374 & ~n20800;
  assign n20802 = ~n20785 & ~n20801;
  assign n20803 = ~n3655 & ~n20802;
  assign n20804 = ~n20772 & ~n20803;
  assign n20805 = ~n3652 & ~n20804;
  assign n20806 = ~n20754 & ~n20805;
  assign n20807 = ~n3368 & ~n20806;
  assign n20808 = n3378 & ~n19258;
  assign n20809 = ~n9865 & ~n20808;
  assign n20810 = n3492 & ~n20809;
  assign n20811 = n3492 & ~n20810;
  assign n20812 = n3485 & ~n20811;
  assign n20813 = n3485 & ~n20812;
  assign n20814 = ~n3476 & ~n20813;
  assign n20815 = ~n5055 & ~n17433;
  assign n20816 = i_hlock0 & ~n20815;
  assign n20817 = ~n9889 & ~n20816;
  assign n20818 = ~i_hbusreq0 & ~n20817;
  assign n20819 = ~n9885 & ~n20818;
  assign n20820 = ~i_hbusreq4 & ~n20819;
  assign n20821 = ~n9884 & ~n20820;
  assign n20822 = ~controllable_hgrant4 & ~n20821;
  assign n20823 = ~n5863 & ~n20822;
  assign n20824 = ~i_hbusreq2 & ~n20823;
  assign n20825 = ~n9883 & ~n20824;
  assign n20826 = ~controllable_hgrant2 & ~n20825;
  assign n20827 = ~n5862 & ~n20826;
  assign n20828 = controllable_hmaster1 & ~n20827;
  assign n20829 = controllable_hmaster0 & ~n20827;
  assign n20830 = ~n3920 & ~n17433;
  assign n20831 = i_hlock0 & ~n20830;
  assign n20832 = ~n5937 & ~n20831;
  assign n20833 = ~i_hbusreq0 & ~n20832;
  assign n20834 = ~n5933 & ~n20833;
  assign n20835 = ~i_hbusreq4 & ~n20834;
  assign n20836 = ~n5932 & ~n20835;
  assign n20837 = ~controllable_hgrant4 & ~n20836;
  assign n20838 = ~n4064 & ~n20837;
  assign n20839 = ~i_hbusreq2 & ~n20838;
  assign n20840 = ~n12262 & ~n20839;
  assign n20841 = ~controllable_hgrant2 & ~n20840;
  assign n20842 = ~n5862 & ~n20841;
  assign n20843 = ~controllable_hmaster0 & ~n20842;
  assign n20844 = ~n20829 & ~n20843;
  assign n20845 = ~controllable_hmaster1 & ~n20844;
  assign n20846 = ~n20828 & ~n20845;
  assign n20847 = ~i_hbusreq3 & ~n20846;
  assign n20848 = ~n13795 & ~n20847;
  assign n20849 = controllable_hmaster2 & ~n20848;
  assign n20850 = ~n5863 & ~n20837;
  assign n20851 = ~i_hbusreq2 & ~n20850;
  assign n20852 = ~n5931 & ~n20851;
  assign n20853 = ~controllable_hgrant2 & ~n20852;
  assign n20854 = ~n5862 & ~n20853;
  assign n20855 = controllable_hmaster0 & ~n20854;
  assign n20856 = ~n5950 & ~n20853;
  assign n20857 = ~controllable_hmaster0 & ~n20856;
  assign n20858 = ~n20855 & ~n20857;
  assign n20859 = controllable_hmaster1 & ~n20858;
  assign n20860 = ~n5730 & ~n18087;
  assign n20861 = ~controllable_ndecide & n20860;
  assign n20862 = ~n3494 & ~n20861;
  assign n20863 = i_hready & ~n20862;
  assign n20864 = ~n4577 & ~n20863;
  assign n20865 = i_hlock0 & ~n20864;
  assign n20866 = ~n9018 & ~n20865;
  assign n20867 = ~i_hbusreq0 & ~n20866;
  assign n20868 = ~n9009 & ~n20867;
  assign n20869 = ~i_hbusreq4 & ~n20868;
  assign n20870 = ~n9008 & ~n20869;
  assign n20871 = ~controllable_hgrant4 & ~n20870;
  assign n20872 = ~n13012 & ~n20871;
  assign n20873 = ~i_hbusreq2 & ~n20872;
  assign n20874 = ~n9007 & ~n20873;
  assign n20875 = ~controllable_hgrant2 & ~n20874;
  assign n20876 = ~n7507 & ~n20875;
  assign n20877 = controllable_hmaster0 & ~n20876;
  assign n20878 = ~n5464 & ~n17433;
  assign n20879 = i_hlock0 & ~n20878;
  assign n20880 = ~n5937 & ~n20879;
  assign n20881 = ~i_hbusreq0 & ~n20880;
  assign n20882 = ~n5933 & ~n20881;
  assign n20883 = ~i_hbusreq4 & ~n20882;
  assign n20884 = ~n5932 & ~n20883;
  assign n20885 = ~controllable_hgrant4 & ~n20884;
  assign n20886 = ~n5982 & ~n20885;
  assign n20887 = ~i_hbusreq2 & ~n20886;
  assign n20888 = ~n5931 & ~n20887;
  assign n20889 = ~controllable_hgrant2 & ~n20888;
  assign n20890 = ~n5981 & ~n20889;
  assign n20891 = ~controllable_hmaster0 & ~n20890;
  assign n20892 = ~n20877 & ~n20891;
  assign n20893 = ~controllable_hmaster1 & ~n20892;
  assign n20894 = ~n20859 & ~n20893;
  assign n20895 = ~i_hbusreq3 & ~n20894;
  assign n20896 = ~n18534 & ~n20895;
  assign n20897 = ~controllable_hmaster2 & ~n20896;
  assign n20898 = ~n20849 & ~n20897;
  assign n20899 = ~controllable_hgrant3 & ~n20898;
  assign n20900 = ~n19398 & ~n20899;
  assign n20901 = controllable_nhgrant0 & ~n20900;
  assign n20902 = ~n10040 & ~n10215;
  assign n20903 = ~controllable_hmaster1 & ~n20902;
  assign n20904 = ~n9966 & ~n20903;
  assign n20905 = i_hbusreq3 & ~n20904;
  assign n20906 = ~n10061 & ~n13834;
  assign n20907 = ~controllable_hmaster1 & ~n20906;
  assign n20908 = ~n10004 & ~n20907;
  assign n20909 = ~i_hbusreq3 & ~n20908;
  assign n20910 = ~n20905 & ~n20909;
  assign n20911 = ~controllable_hmaster2 & ~n20910;
  assign n20912 = ~n13828 & ~n20911;
  assign n20913 = ~controllable_hgrant3 & ~n20912;
  assign n20914 = ~n19241 & ~n20913;
  assign n20915 = ~controllable_nhgrant0 & ~n20914;
  assign n20916 = ~n20901 & ~n20915;
  assign n20917 = ~n3281 & ~n20916;
  assign n20918 = ~n3281 & ~n20917;
  assign n20919 = n3378 & ~n20918;
  assign n20920 = ~n10244 & ~n20919;
  assign n20921 = n3492 & ~n20920;
  assign n20922 = ~n8536 & ~n20921;
  assign n20923 = n3485 & ~n20922;
  assign n20924 = ~n8694 & ~n20923;
  assign n20925 = n3476 & ~n20924;
  assign n20926 = ~n20814 & ~n20925;
  assign n20927 = n3374 & ~n20926;
  assign n20928 = ~n9769 & ~n20927;
  assign n20929 = n3655 & ~n20928;
  assign n20930 = n3378 & ~n19623;
  assign n20931 = ~n10299 & ~n20930;
  assign n20932 = n3492 & ~n20931;
  assign n20933 = n3492 & ~n20932;
  assign n20934 = n3485 & ~n20933;
  assign n20935 = n3485 & ~n20934;
  assign n20936 = ~n3476 & ~n20935;
  assign n20937 = ~n8523 & ~n20932;
  assign n20938 = n3485 & ~n20937;
  assign n20939 = ~n8689 & ~n20938;
  assign n20940 = n3476 & ~n20939;
  assign n20941 = ~n20936 & ~n20940;
  assign n20942 = ~n3374 & ~n20941;
  assign n20943 = n3378 & ~n19792;
  assign n20944 = ~n10390 & ~n20943;
  assign n20945 = n3492 & ~n20944;
  assign n20946 = n3492 & ~n20945;
  assign n20947 = n3485 & ~n20946;
  assign n20948 = n3485 & ~n20947;
  assign n20949 = ~n3476 & ~n20948;
  assign n20950 = ~n10401 & ~n19958;
  assign n20951 = ~controllable_hgrant4 & n20950;
  assign n20952 = ~n4091 & ~n20951;
  assign n20953 = ~controllable_hgrant2 & ~n20952;
  assign n20954 = ~n5616 & ~n20953;
  assign n20955 = controllable_hmaster1 & ~n20954;
  assign n20956 = controllable_hmaster0 & ~n20954;
  assign n20957 = ~n10401 & ~n19969;
  assign n20958 = ~controllable_hgrant4 & n20957;
  assign n20959 = ~n4015 & ~n20958;
  assign n20960 = ~controllable_hgrant2 & ~n20959;
  assign n20961 = ~n5616 & ~n20960;
  assign n20962 = ~controllable_hmaster0 & ~n20961;
  assign n20963 = ~n20956 & ~n20962;
  assign n20964 = ~controllable_hmaster1 & ~n20963;
  assign n20965 = ~n20955 & ~n20964;
  assign n20966 = i_hbusreq3 & ~n20965;
  assign n20967 = i_hbusreq2 & ~n20952;
  assign n20968 = i_hbusreq4 & ~n20950;
  assign n20969 = i_hbusreq0 & ~n20950;
  assign n20970 = ~n10424 & ~n18087;
  assign n20971 = ~controllable_ndecide & ~n20970;
  assign n20972 = ~controllable_ndecide & ~n20971;
  assign n20973 = i_hready & ~n20972;
  assign n20974 = ~n19985 & ~n20973;
  assign n20975 = i_hlock0 & ~n20974;
  assign n20976 = ~n10435 & ~n19958;
  assign n20977 = ~i_hlock0 & ~n20976;
  assign n20978 = ~n20975 & ~n20977;
  assign n20979 = ~i_hbusreq0 & ~n20978;
  assign n20980 = ~n20969 & ~n20979;
  assign n20981 = ~i_hbusreq4 & ~n20980;
  assign n20982 = ~n20968 & ~n20981;
  assign n20983 = ~controllable_hgrant4 & n20982;
  assign n20984 = ~n5863 & ~n20983;
  assign n20985 = ~i_hbusreq2 & ~n20984;
  assign n20986 = ~n20967 & ~n20985;
  assign n20987 = ~controllable_hgrant2 & ~n20986;
  assign n20988 = ~n5862 & ~n20987;
  assign n20989 = controllable_hmaster1 & ~n20988;
  assign n20990 = controllable_hmaster0 & ~n20988;
  assign n20991 = i_hbusreq2 & ~n20959;
  assign n20992 = i_hbusreq4 & ~n20957;
  assign n20993 = i_hbusreq0 & ~n20957;
  assign n20994 = ~n20012 & ~n20973;
  assign n20995 = i_hlock0 & ~n20994;
  assign n20996 = ~n10460 & ~n19969;
  assign n20997 = ~i_hlock0 & ~n20996;
  assign n20998 = ~n20995 & ~n20997;
  assign n20999 = ~i_hbusreq0 & ~n20998;
  assign n21000 = ~n20993 & ~n20999;
  assign n21001 = ~i_hbusreq4 & ~n21000;
  assign n21002 = ~n20992 & ~n21001;
  assign n21003 = ~controllable_hgrant4 & n21002;
  assign n21004 = ~n4064 & ~n21003;
  assign n21005 = ~i_hbusreq2 & ~n21004;
  assign n21006 = ~n20991 & ~n21005;
  assign n21007 = ~controllable_hgrant2 & ~n21006;
  assign n21008 = ~n5862 & ~n21007;
  assign n21009 = ~controllable_hmaster0 & ~n21008;
  assign n21010 = ~n20990 & ~n21009;
  assign n21011 = ~controllable_hmaster1 & ~n21010;
  assign n21012 = ~n20989 & ~n21011;
  assign n21013 = ~i_hbusreq3 & ~n21012;
  assign n21014 = ~n20966 & ~n21013;
  assign n21015 = controllable_hmaster2 & ~n21014;
  assign n21016 = ~n4091 & ~n20958;
  assign n21017 = ~controllable_hgrant2 & ~n21016;
  assign n21018 = ~n5616 & ~n21017;
  assign n21019 = controllable_hmaster0 & ~n21018;
  assign n21020 = ~n5686 & ~n21017;
  assign n21021 = ~controllable_hmaster0 & ~n21020;
  assign n21022 = ~n21019 & ~n21021;
  assign n21023 = controllable_hmaster1 & ~n21022;
  assign n21024 = ~controllable_hmaster0 & ~n21018;
  assign n21025 = ~n10642 & ~n21024;
  assign n21026 = ~controllable_hmaster1 & ~n21025;
  assign n21027 = ~n21023 & ~n21026;
  assign n21028 = i_hbusreq3 & ~n21027;
  assign n21029 = i_hbusreq2 & ~n21016;
  assign n21030 = ~n5863 & ~n21003;
  assign n21031 = ~i_hbusreq2 & ~n21030;
  assign n21032 = ~n21029 & ~n21031;
  assign n21033 = ~controllable_hgrant2 & ~n21032;
  assign n21034 = ~n5862 & ~n21033;
  assign n21035 = controllable_hmaster0 & ~n21034;
  assign n21036 = ~n5950 & ~n21033;
  assign n21037 = ~controllable_hmaster0 & ~n21036;
  assign n21038 = ~n21035 & ~n21037;
  assign n21039 = controllable_hmaster1 & ~n21038;
  assign n21040 = ~n10535 & ~n18087;
  assign n21041 = ~controllable_ndecide & ~n21040;
  assign n21042 = ~controllable_ndecide & ~n21041;
  assign n21043 = i_hready & ~n21042;
  assign n21044 = ~n10361 & ~n21043;
  assign n21045 = i_hlock0 & ~n21044;
  assign n21046 = ~n10668 & ~n21045;
  assign n21047 = ~i_hbusreq0 & ~n21046;
  assign n21048 = ~n10660 & ~n21047;
  assign n21049 = ~i_hbusreq4 & ~n21048;
  assign n21050 = ~n10659 & ~n21049;
  assign n21051 = ~controllable_hgrant4 & n21050;
  assign n21052 = ~n13012 & ~n21051;
  assign n21053 = ~i_hbusreq2 & ~n21052;
  assign n21054 = ~n10658 & ~n21053;
  assign n21055 = ~controllable_hgrant2 & ~n21054;
  assign n21056 = ~n7507 & ~n21055;
  assign n21057 = controllable_hmaster0 & ~n21056;
  assign n21058 = ~n20096 & ~n20973;
  assign n21059 = i_hlock0 & ~n21058;
  assign n21060 = ~n20997 & ~n21059;
  assign n21061 = ~i_hbusreq0 & ~n21060;
  assign n21062 = ~n20993 & ~n21061;
  assign n21063 = ~i_hbusreq4 & ~n21062;
  assign n21064 = ~n20992 & ~n21063;
  assign n21065 = ~controllable_hgrant4 & n21064;
  assign n21066 = ~n5982 & ~n21065;
  assign n21067 = ~i_hbusreq2 & ~n21066;
  assign n21068 = ~n21029 & ~n21067;
  assign n21069 = ~controllable_hgrant2 & ~n21068;
  assign n21070 = ~n5981 & ~n21069;
  assign n21071 = ~controllable_hmaster0 & ~n21070;
  assign n21072 = ~n21057 & ~n21071;
  assign n21073 = ~controllable_hmaster1 & ~n21072;
  assign n21074 = ~n21039 & ~n21073;
  assign n21075 = ~i_hbusreq3 & ~n21074;
  assign n21076 = ~n21028 & ~n21075;
  assign n21077 = ~controllable_hmaster2 & ~n21076;
  assign n21078 = ~n21015 & ~n21077;
  assign n21079 = ~controllable_hgrant3 & ~n21078;
  assign n21080 = ~n19398 & ~n21079;
  assign n21081 = controllable_nhgrant0 & ~n21080;
  assign n21082 = ~n20915 & ~n21081;
  assign n21083 = ~n3281 & ~n21082;
  assign n21084 = ~n3281 & ~n21083;
  assign n21085 = n3378 & ~n21084;
  assign n21086 = ~n10705 & ~n21085;
  assign n21087 = n3492 & ~n21086;
  assign n21088 = ~n8563 & ~n21087;
  assign n21089 = n3485 & ~n21088;
  assign n21090 = ~n8705 & ~n21089;
  assign n21091 = n3476 & ~n21090;
  assign n21092 = ~n20949 & ~n21091;
  assign n21093 = n3374 & ~n21092;
  assign n21094 = ~n20942 & ~n21093;
  assign n21095 = ~n3655 & ~n21094;
  assign n21096 = ~n20929 & ~n21095;
  assign n21097 = n3652 & ~n21096;
  assign n21098 = n3378 & ~n20171;
  assign n21099 = ~n10802 & ~n21098;
  assign n21100 = n3492 & ~n21099;
  assign n21101 = n3492 & ~n21100;
  assign n21102 = n3485 & ~n21101;
  assign n21103 = n3485 & ~n21102;
  assign n21104 = ~n3476 & ~n21103;
  assign n21105 = ~n10870 & ~n20826;
  assign n21106 = controllable_hmaster1 & ~n21105;
  assign n21107 = controllable_hmaster0 & ~n21105;
  assign n21108 = ~n10870 & ~n20841;
  assign n21109 = ~controllable_hmaster0 & ~n21108;
  assign n21110 = ~n21107 & ~n21109;
  assign n21111 = ~controllable_hmaster1 & ~n21110;
  assign n21112 = ~n21106 & ~n21111;
  assign n21113 = ~i_hbusreq3 & ~n21112;
  assign n21114 = ~n13963 & ~n21113;
  assign n21115 = controllable_hmaster2 & ~n21114;
  assign n21116 = ~n10929 & ~n11072;
  assign n21117 = ~controllable_hmaster1 & ~n21116;
  assign n21118 = ~n10926 & ~n21117;
  assign n21119 = i_hbusreq3 & ~n21118;
  assign n21120 = ~n10870 & ~n20853;
  assign n21121 = controllable_hmaster0 & ~n21120;
  assign n21122 = ~n10972 & ~n20853;
  assign n21123 = ~controllable_hmaster0 & ~n21122;
  assign n21124 = ~n21121 & ~n21123;
  assign n21125 = controllable_hmaster1 & ~n21124;
  assign n21126 = ~n10904 & ~n20875;
  assign n21127 = controllable_hmaster0 & ~n21126;
  assign n21128 = ~n11002 & ~n20889;
  assign n21129 = ~controllable_hmaster0 & ~n21128;
  assign n21130 = ~n21127 & ~n21129;
  assign n21131 = ~controllable_hmaster1 & ~n21130;
  assign n21132 = ~n21125 & ~n21131;
  assign n21133 = ~i_hbusreq3 & ~n21132;
  assign n21134 = ~n21119 & ~n21133;
  assign n21135 = ~controllable_hmaster2 & ~n21134;
  assign n21136 = ~n21115 & ~n21135;
  assign n21137 = ~controllable_hgrant3 & ~n21136;
  assign n21138 = ~n19398 & ~n21137;
  assign n21139 = controllable_nhgrant0 & ~n21138;
  assign n21140 = ~n20915 & ~n21139;
  assign n21141 = ~n3281 & ~n21140;
  assign n21142 = ~n3281 & ~n21141;
  assign n21143 = n3378 & ~n21142;
  assign n21144 = ~n11143 & ~n21143;
  assign n21145 = n3492 & ~n21144;
  assign n21146 = ~n8592 & ~n21145;
  assign n21147 = n3485 & ~n21146;
  assign n21148 = ~n8718 & ~n21147;
  assign n21149 = n3476 & ~n21148;
  assign n21150 = ~n21104 & ~n21149;
  assign n21151 = n3374 & ~n21150;
  assign n21152 = ~n10754 & ~n21151;
  assign n21153 = n3655 & ~n21152;
  assign n21154 = n3378 & ~n20274;
  assign n21155 = ~n11178 & ~n21154;
  assign n21156 = n3492 & ~n21155;
  assign n21157 = n3492 & ~n21156;
  assign n21158 = n3485 & ~n21157;
  assign n21159 = n3485 & ~n21158;
  assign n21160 = ~n3476 & ~n21159;
  assign n21161 = ~n8523 & ~n21156;
  assign n21162 = n3485 & ~n21161;
  assign n21163 = ~n8689 & ~n21162;
  assign n21164 = n3476 & ~n21163;
  assign n21165 = ~n21160 & ~n21164;
  assign n21166 = ~n3374 & ~n21165;
  assign n21167 = n3378 & ~n20345;
  assign n21168 = ~n11236 & ~n21167;
  assign n21169 = n3492 & ~n21168;
  assign n21170 = n3492 & ~n21169;
  assign n21171 = n3485 & ~n21170;
  assign n21172 = n3485 & ~n21171;
  assign n21173 = ~n3476 & ~n21172;
  assign n21174 = ~n10816 & ~n20953;
  assign n21175 = controllable_hmaster1 & ~n21174;
  assign n21176 = controllable_hmaster0 & ~n21174;
  assign n21177 = ~n10816 & ~n20960;
  assign n21178 = ~controllable_hmaster0 & ~n21177;
  assign n21179 = ~n21176 & ~n21178;
  assign n21180 = ~controllable_hmaster1 & ~n21179;
  assign n21181 = ~n21175 & ~n21180;
  assign n21182 = i_hbusreq3 & ~n21181;
  assign n21183 = ~n10870 & ~n20987;
  assign n21184 = controllable_hmaster1 & ~n21183;
  assign n21185 = controllable_hmaster0 & ~n21183;
  assign n21186 = ~n10870 & ~n21007;
  assign n21187 = ~controllable_hmaster0 & ~n21186;
  assign n21188 = ~n21185 & ~n21187;
  assign n21189 = ~controllable_hmaster1 & ~n21188;
  assign n21190 = ~n21184 & ~n21189;
  assign n21191 = ~i_hbusreq3 & ~n21190;
  assign n21192 = ~n21182 & ~n21191;
  assign n21193 = controllable_hmaster2 & ~n21192;
  assign n21194 = ~n10816 & ~n21017;
  assign n21195 = controllable_hmaster0 & ~n21194;
  assign n21196 = ~n10922 & ~n21017;
  assign n21197 = ~controllable_hmaster0 & ~n21196;
  assign n21198 = ~n21195 & ~n21197;
  assign n21199 = controllable_hmaster1 & ~n21198;
  assign n21200 = ~controllable_hmaster0 & ~n21194;
  assign n21201 = ~n11323 & ~n21200;
  assign n21202 = ~controllable_hmaster1 & ~n21201;
  assign n21203 = ~n21199 & ~n21202;
  assign n21204 = i_hbusreq3 & ~n21203;
  assign n21205 = ~n10870 & ~n21033;
  assign n21206 = controllable_hmaster0 & ~n21205;
  assign n21207 = ~n10972 & ~n21033;
  assign n21208 = ~controllable_hmaster0 & ~n21207;
  assign n21209 = ~n21206 & ~n21208;
  assign n21210 = controllable_hmaster1 & ~n21209;
  assign n21211 = ~n10904 & ~n21055;
  assign n21212 = controllable_hmaster0 & ~n21211;
  assign n21213 = ~n11002 & ~n21069;
  assign n21214 = ~controllable_hmaster0 & ~n21213;
  assign n21215 = ~n21212 & ~n21214;
  assign n21216 = ~controllable_hmaster1 & ~n21215;
  assign n21217 = ~n21210 & ~n21216;
  assign n21218 = ~i_hbusreq3 & ~n21217;
  assign n21219 = ~n21204 & ~n21218;
  assign n21220 = ~controllable_hmaster2 & ~n21219;
  assign n21221 = ~n21193 & ~n21220;
  assign n21222 = ~controllable_hgrant3 & ~n21221;
  assign n21223 = ~n19398 & ~n21222;
  assign n21224 = controllable_nhgrant0 & ~n21223;
  assign n21225 = ~n20915 & ~n21224;
  assign n21226 = ~n3281 & ~n21225;
  assign n21227 = ~n3281 & ~n21226;
  assign n21228 = n3378 & ~n21227;
  assign n21229 = ~n11352 & ~n21228;
  assign n21230 = n3492 & ~n21229;
  assign n21231 = ~n8619 & ~n21230;
  assign n21232 = n3485 & ~n21231;
  assign n21233 = ~n8729 & ~n21232;
  assign n21234 = n3476 & ~n21233;
  assign n21235 = ~n21173 & ~n21234;
  assign n21236 = n3374 & ~n21235;
  assign n21237 = ~n21166 & ~n21236;
  assign n21238 = ~n3655 & ~n21237;
  assign n21239 = ~n21153 & ~n21238;
  assign n21240 = ~n3652 & ~n21239;
  assign n21241 = ~n21097 & ~n21240;
  assign n21242 = n3368 & ~n21241;
  assign n21243 = ~n20807 & ~n21242;
  assign n21244 = ~n3362 & ~n21243;
  assign n21245 = ~n20703 & ~n21244;
  assign n21246 = ~n3359 & ~n21245;
  assign n21247 = ~n20625 & ~n21246;
  assign n21248 = ~n3356 & ~n21247;
  assign n21249 = ~n18368 & ~n21248;
  assign n21250 = ~n3345 & ~n21249;
  assign n21251 = ~controllable_hmaster2 & ~n8291;
  assign n21252 = controllable_nhgrant0 & ~n21251;
  assign n21253 = controllable_hgrant3 & ~n21251;
  assign n21254 = ~controllable_hmaster2 & ~n8301;
  assign n21255 = ~controllable_hgrant3 & ~n21254;
  assign n21256 = ~n21253 & ~n21255;
  assign n21257 = ~controllable_nhgrant0 & ~n21256;
  assign n21258 = ~n21252 & ~n21257;
  assign n21259 = ~n3281 & ~n21258;
  assign n21260 = ~n3281 & ~n21259;
  assign n21261 = n3378 & ~n21260;
  assign n21262 = controllable_hmaster2 & ~n3385;
  assign n21263 = ~n8291 & ~n21262;
  assign n21264 = controllable_hgrant3 & ~n21263;
  assign n21265 = controllable_hmaster2 & ~n3429;
  assign n21266 = ~n8291 & ~n21265;
  assign n21267 = ~controllable_hgrant3 & ~n21266;
  assign n21268 = ~n21264 & ~n21267;
  assign n21269 = controllable_nhgrant0 & ~n21268;
  assign n21270 = ~controllable_hmaster1 & ~n11461;
  assign n21271 = ~n8770 & ~n21270;
  assign n21272 = controllable_hmaster2 & ~n21271;
  assign n21273 = ~n8301 & ~n21272;
  assign n21274 = ~controllable_hgrant3 & ~n21273;
  assign n21275 = ~n21264 & ~n21274;
  assign n21276 = ~controllable_nhgrant0 & ~n21275;
  assign n21277 = ~n21269 & ~n21276;
  assign n21278 = ~n3281 & ~n21277;
  assign n21279 = ~n3783 & ~n21278;
  assign n21280 = ~n3378 & ~n21279;
  assign n21281 = ~n21261 & ~n21280;
  assign n21282 = n3492 & ~n21281;
  assign n21283 = ~n3493 & ~n21282;
  assign n21284 = n3485 & ~n21283;
  assign n21285 = ~n3486 & ~n21284;
  assign n21286 = ~n3476 & ~n21285;
  assign n21287 = ~n3378 & ~n8308;
  assign n21288 = ~n21261 & ~n21287;
  assign n21289 = ~n3485 & ~n21288;
  assign n21290 = ~n3492 & ~n21288;
  assign n21291 = ~n21282 & ~n21290;
  assign n21292 = n3485 & ~n21291;
  assign n21293 = ~n21289 & ~n21292;
  assign n21294 = n3476 & ~n21293;
  assign n21295 = ~n21286 & ~n21294;
  assign n21296 = ~n3374 & ~n21295;
  assign n21297 = ~controllable_hmaster0 & ~n5394;
  assign n21298 = ~controllable_hmaster1 & ~n21297;
  assign n21299 = ~controllable_hmaster1 & ~n21298;
  assign n21300 = ~i_hbusreq3 & ~n21299;
  assign n21301 = ~n3825 & ~n21300;
  assign n21302 = ~controllable_hmaster2 & ~n21301;
  assign n21303 = ~controllable_hmaster2 & ~n21302;
  assign n21304 = controllable_hgrant3 & ~n21303;
  assign n21305 = ~controllable_hmaster0 & ~n8827;
  assign n21306 = ~controllable_hmaster1 & ~n21305;
  assign n21307 = ~controllable_hmaster1 & ~n21306;
  assign n21308 = i_hbusreq3 & ~n21307;
  assign n21309 = ~controllable_hmaster0 & ~n8876;
  assign n21310 = ~controllable_hmaster1 & ~n21309;
  assign n21311 = ~controllable_hmaster1 & ~n21310;
  assign n21312 = ~i_hbusreq3 & ~n21311;
  assign n21313 = ~n21308 & ~n21312;
  assign n21314 = ~controllable_hmaster2 & ~n21313;
  assign n21315 = ~controllable_hmaster2 & ~n21314;
  assign n21316 = ~controllable_hgrant3 & ~n21315;
  assign n21317 = ~n21304 & ~n21316;
  assign n21318 = controllable_nhgrant0 & ~n21317;
  assign n21319 = ~controllable_hmaster0 & ~n5499;
  assign n21320 = ~controllable_hmaster1 & ~n21319;
  assign n21321 = ~controllable_hmaster1 & ~n21320;
  assign n21322 = i_hbusreq3 & ~n21321;
  assign n21323 = ~controllable_hmaster0 & ~n5524;
  assign n21324 = ~controllable_hmaster1 & ~n21323;
  assign n21325 = ~controllable_hmaster1 & ~n21324;
  assign n21326 = ~i_hbusreq3 & ~n21325;
  assign n21327 = ~n21322 & ~n21326;
  assign n21328 = ~controllable_hmaster2 & ~n21327;
  assign n21329 = ~controllable_hmaster2 & ~n21328;
  assign n21330 = ~controllable_hgrant3 & ~n21329;
  assign n21331 = ~n21304 & ~n21330;
  assign n21332 = ~controllable_nhgrant0 & ~n21331;
  assign n21333 = ~n21318 & ~n21332;
  assign n21334 = ~n3281 & ~n21333;
  assign n21335 = ~n3281 & ~n21334;
  assign n21336 = n3378 & ~n21335;
  assign n21337 = ~n21262 & ~n21302;
  assign n21338 = controllable_hgrant3 & ~n21337;
  assign n21339 = controllable_hmaster2 & ~n3505;
  assign n21340 = ~n21314 & ~n21339;
  assign n21341 = ~controllable_hgrant3 & ~n21340;
  assign n21342 = ~n21338 & ~n21341;
  assign n21343 = controllable_nhgrant0 & ~n21342;
  assign n21344 = ~n21272 & ~n21328;
  assign n21345 = ~controllable_hgrant3 & ~n21344;
  assign n21346 = ~n21338 & ~n21345;
  assign n21347 = ~controllable_nhgrant0 & ~n21346;
  assign n21348 = ~n21343 & ~n21347;
  assign n21349 = ~n3281 & ~n21348;
  assign n21350 = ~n3950 & ~n21349;
  assign n21351 = ~n3378 & ~n21350;
  assign n21352 = ~n21336 & ~n21351;
  assign n21353 = n3492 & ~n21352;
  assign n21354 = ~n3493 & ~n21353;
  assign n21355 = n3485 & ~n21354;
  assign n21356 = ~n3486 & ~n21355;
  assign n21357 = ~n3476 & ~n21356;
  assign n21358 = ~controllable_hgrant2 & ~n14487;
  assign n21359 = ~controllable_hgrant2 & ~n21358;
  assign n21360 = i_hbusreq3 & ~n21359;
  assign n21361 = ~controllable_hgrant2 & ~n14505;
  assign n21362 = ~controllable_hgrant2 & ~n21361;
  assign n21363 = ~i_hbusreq3 & ~n21362;
  assign n21364 = ~n21360 & ~n21363;
  assign n21365 = controllable_hmaster2 & ~n21364;
  assign n21366 = controllable_hmaster1 & ~n21359;
  assign n21367 = controllable_hmaster0 & ~n21359;
  assign n21368 = ~n6044 & ~n21367;
  assign n21369 = ~controllable_hmaster1 & ~n21368;
  assign n21370 = ~n21366 & ~n21369;
  assign n21371 = i_hbusreq3 & ~n21370;
  assign n21372 = controllable_hmaster1 & ~n21362;
  assign n21373 = controllable_hmaster0 & ~n21362;
  assign n21374 = ~n6072 & ~n21373;
  assign n21375 = ~controllable_hmaster1 & ~n21374;
  assign n21376 = ~n21372 & ~n21375;
  assign n21377 = ~i_hbusreq3 & ~n21376;
  assign n21378 = ~n21371 & ~n21377;
  assign n21379 = ~controllable_hmaster2 & ~n21378;
  assign n21380 = ~n21365 & ~n21379;
  assign n21381 = ~controllable_hgrant3 & ~n21380;
  assign n21382 = ~n21304 & ~n21381;
  assign n21383 = ~controllable_nhgrant0 & ~n21382;
  assign n21384 = ~n21318 & ~n21383;
  assign n21385 = ~n3281 & ~n21384;
  assign n21386 = ~n3281 & ~n21385;
  assign n21387 = n3378 & ~n21386;
  assign n21388 = ~i_hbusreq0 & ~n11083;
  assign n21389 = ~n3563 & ~n21388;
  assign n21390 = ~i_hbusreq4 & ~n21389;
  assign n21391 = ~n3562 & ~n21390;
  assign n21392 = ~controllable_hgrant4 & ~n21391;
  assign n21393 = ~n3411 & ~n21392;
  assign n21394 = ~i_hbusreq2 & ~n21393;
  assign n21395 = ~n3561 & ~n21394;
  assign n21396 = ~controllable_hgrant2 & ~n21395;
  assign n21397 = ~n3410 & ~n21396;
  assign n21398 = controllable_hmaster1 & ~n21397;
  assign n21399 = controllable_hmaster0 & ~n21397;
  assign n21400 = ~i_hbusreq2 & ~n14853;
  assign n21401 = ~n3582 & ~n21400;
  assign n21402 = ~controllable_hgrant2 & ~n21401;
  assign n21403 = ~controllable_hgrant2 & ~n21402;
  assign n21404 = ~controllable_hmaster0 & ~n21403;
  assign n21405 = ~n21399 & ~n21404;
  assign n21406 = ~controllable_hmaster1 & ~n21405;
  assign n21407 = ~n21398 & ~n21406;
  assign n21408 = ~i_hbusreq3 & ~n21407;
  assign n21409 = ~n3560 & ~n21408;
  assign n21410 = controllable_hmaster2 & ~n21409;
  assign n21411 = controllable_hmaster1 & ~n3555;
  assign n21412 = controllable_hmaster0 & ~n3555;
  assign n21413 = ~controllable_hmaster0 & ~n3548;
  assign n21414 = ~n21412 & ~n21413;
  assign n21415 = ~controllable_hmaster1 & ~n21414;
  assign n21416 = ~n21411 & ~n21415;
  assign n21417 = i_hbusreq3 & ~n21416;
  assign n21418 = controllable_hmaster1 & ~n21403;
  assign n21419 = controllable_hmaster0 & ~n21403;
  assign n21420 = ~n8862 & ~n10842;
  assign n21421 = i_hlock0 & ~n21420;
  assign n21422 = ~n3495 & ~n10842;
  assign n21423 = ~i_hlock0 & ~n21422;
  assign n21424 = ~n21421 & ~n21423;
  assign n21425 = ~i_hbusreq0 & ~n21424;
  assign n21426 = ~n3563 & ~n21425;
  assign n21427 = ~i_hbusreq4 & ~n21426;
  assign n21428 = ~n3562 & ~n21427;
  assign n21429 = ~controllable_hgrant4 & ~n21428;
  assign n21430 = ~n5462 & ~n21429;
  assign n21431 = ~i_hbusreq2 & ~n21430;
  assign n21432 = ~n3561 & ~n21431;
  assign n21433 = ~controllable_hgrant2 & ~n21432;
  assign n21434 = ~n5461 & ~n21433;
  assign n21435 = ~controllable_hmaster0 & ~n21434;
  assign n21436 = ~n21419 & ~n21435;
  assign n21437 = ~controllable_hmaster1 & ~n21436;
  assign n21438 = ~n21418 & ~n21437;
  assign n21439 = ~i_hbusreq3 & ~n21438;
  assign n21440 = ~n21417 & ~n21439;
  assign n21441 = ~controllable_hmaster2 & ~n21440;
  assign n21442 = ~n21410 & ~n21441;
  assign n21443 = ~controllable_hgrant3 & ~n21442;
  assign n21444 = ~n21338 & ~n21443;
  assign n21445 = controllable_nhgrant0 & ~n21444;
  assign n21446 = ~controllable_hmaster0 & ~n21359;
  assign n21447 = ~n9061 & ~n21446;
  assign n21448 = ~controllable_hmaster1 & ~n21447;
  assign n21449 = ~n9060 & ~n21448;
  assign n21450 = i_hbusreq3 & ~n21449;
  assign n21451 = ~controllable_hmaster0 & ~n21362;
  assign n21452 = ~n9085 & ~n21451;
  assign n21453 = ~controllable_hmaster1 & ~n21452;
  assign n21454 = ~n9084 & ~n21453;
  assign n21455 = ~i_hbusreq3 & ~n21454;
  assign n21456 = ~n21450 & ~n21455;
  assign n21457 = controllable_hmaster2 & ~n21456;
  assign n21458 = ~n21379 & ~n21457;
  assign n21459 = ~controllable_hgrant3 & ~n21458;
  assign n21460 = ~n21338 & ~n21459;
  assign n21461 = ~controllable_nhgrant0 & ~n21460;
  assign n21462 = ~n21445 & ~n21461;
  assign n21463 = ~n3281 & ~n21462;
  assign n21464 = ~n4089 & ~n21463;
  assign n21465 = ~n3378 & ~n21464;
  assign n21466 = ~n21387 & ~n21465;
  assign n21467 = n3492 & ~n21466;
  assign n21468 = ~n21290 & ~n21467;
  assign n21469 = n3485 & ~n21468;
  assign n21470 = ~n21289 & ~n21469;
  assign n21471 = n3476 & ~n21470;
  assign n21472 = ~n21357 & ~n21471;
  assign n21473 = n3374 & ~n21472;
  assign n21474 = ~n21296 & ~n21473;
  assign n21475 = n3655 & ~n21474;
  assign n21476 = ~controllable_hmaster0 & ~n9175;
  assign n21477 = ~controllable_hmaster1 & ~n21476;
  assign n21478 = ~controllable_hmaster1 & ~n21477;
  assign n21479 = i_hbusreq3 & ~n21478;
  assign n21480 = ~controllable_hmaster0 & ~n9226;
  assign n21481 = ~controllable_hmaster1 & ~n21480;
  assign n21482 = ~controllable_hmaster1 & ~n21481;
  assign n21483 = ~i_hbusreq3 & ~n21482;
  assign n21484 = ~n21479 & ~n21483;
  assign n21485 = ~controllable_hmaster2 & ~n21484;
  assign n21486 = ~controllable_hmaster2 & ~n21485;
  assign n21487 = ~controllable_hgrant3 & ~n21486;
  assign n21488 = ~n21304 & ~n21487;
  assign n21489 = controllable_nhgrant0 & ~n21488;
  assign n21490 = ~n21332 & ~n21489;
  assign n21491 = ~n3281 & ~n21490;
  assign n21492 = ~n3281 & ~n21491;
  assign n21493 = n3378 & ~n21492;
  assign n21494 = ~n21339 & ~n21485;
  assign n21495 = ~controllable_hgrant3 & ~n21494;
  assign n21496 = ~n21338 & ~n21495;
  assign n21497 = controllable_nhgrant0 & ~n21496;
  assign n21498 = ~n21347 & ~n21497;
  assign n21499 = ~n3281 & ~n21498;
  assign n21500 = ~n3950 & ~n21499;
  assign n21501 = ~n3378 & ~n21500;
  assign n21502 = ~n21493 & ~n21501;
  assign n21503 = n3492 & ~n21502;
  assign n21504 = ~n3493 & ~n21503;
  assign n21505 = n3485 & ~n21504;
  assign n21506 = ~n3486 & ~n21505;
  assign n21507 = ~n3476 & ~n21506;
  assign n21508 = ~n21383 & ~n21489;
  assign n21509 = ~n3281 & ~n21508;
  assign n21510 = ~n3281 & ~n21509;
  assign n21511 = n3378 & ~n21510;
  assign n21512 = ~controllable_hmaster0 & ~n11655;
  assign n21513 = ~n21412 & ~n21512;
  assign n21514 = ~controllable_hmaster1 & ~n21513;
  assign n21515 = ~n21411 & ~n21514;
  assign n21516 = i_hbusreq3 & ~n21515;
  assign n21517 = ~n9212 & ~n10842;
  assign n21518 = i_hlock0 & ~n21517;
  assign n21519 = ~n4180 & ~n10842;
  assign n21520 = ~i_hlock0 & ~n21519;
  assign n21521 = ~n21518 & ~n21520;
  assign n21522 = ~i_hbusreq0 & ~n21521;
  assign n21523 = ~n4290 & ~n21522;
  assign n21524 = ~i_hbusreq4 & ~n21523;
  assign n21525 = ~n4289 & ~n21524;
  assign n21526 = ~controllable_hgrant4 & ~n21525;
  assign n21527 = ~n5462 & ~n21526;
  assign n21528 = ~i_hbusreq2 & ~n21527;
  assign n21529 = ~n11661 & ~n21528;
  assign n21530 = ~controllable_hgrant2 & ~n21529;
  assign n21531 = ~n5461 & ~n21530;
  assign n21532 = ~controllable_hmaster0 & ~n21531;
  assign n21533 = ~n21419 & ~n21532;
  assign n21534 = ~controllable_hmaster1 & ~n21533;
  assign n21535 = ~n21418 & ~n21534;
  assign n21536 = ~i_hbusreq3 & ~n21535;
  assign n21537 = ~n21516 & ~n21536;
  assign n21538 = ~controllable_hmaster2 & ~n21537;
  assign n21539 = ~n21410 & ~n21538;
  assign n21540 = ~controllable_hgrant3 & ~n21539;
  assign n21541 = ~n21338 & ~n21540;
  assign n21542 = controllable_nhgrant0 & ~n21541;
  assign n21543 = ~n21461 & ~n21542;
  assign n21544 = ~n3281 & ~n21543;
  assign n21545 = ~n4089 & ~n21544;
  assign n21546 = ~n3378 & ~n21545;
  assign n21547 = ~n21511 & ~n21546;
  assign n21548 = n3492 & ~n21547;
  assign n21549 = ~n21290 & ~n21548;
  assign n21550 = n3485 & ~n21549;
  assign n21551 = ~n21289 & ~n21550;
  assign n21552 = n3476 & ~n21551;
  assign n21553 = ~n21507 & ~n21552;
  assign n21554 = n3374 & ~n21553;
  assign n21555 = ~n21296 & ~n21554;
  assign n21556 = ~n3655 & ~n21555;
  assign n21557 = ~n21475 & ~n21556;
  assign n21558 = n3652 & ~n21557;
  assign n21559 = ~controllable_hmaster0 & ~n9441;
  assign n21560 = ~controllable_hmaster1 & ~n21559;
  assign n21561 = ~controllable_hmaster1 & ~n21560;
  assign n21562 = i_hbusreq3 & ~n21561;
  assign n21563 = ~controllable_hmaster0 & ~n9455;
  assign n21564 = ~controllable_hmaster1 & ~n21563;
  assign n21565 = ~controllable_hmaster1 & ~n21564;
  assign n21566 = ~i_hbusreq3 & ~n21565;
  assign n21567 = ~n21562 & ~n21566;
  assign n21568 = ~controllable_hmaster2 & ~n21567;
  assign n21569 = ~controllable_hmaster2 & ~n21568;
  assign n21570 = ~controllable_hgrant3 & ~n21569;
  assign n21571 = ~n21304 & ~n21570;
  assign n21572 = controllable_nhgrant0 & ~n21571;
  assign n21573 = ~n21332 & ~n21572;
  assign n21574 = ~n3281 & ~n21573;
  assign n21575 = ~n3281 & ~n21574;
  assign n21576 = n3378 & ~n21575;
  assign n21577 = ~n21339 & ~n21568;
  assign n21578 = ~controllable_hgrant3 & ~n21577;
  assign n21579 = ~n21338 & ~n21578;
  assign n21580 = controllable_nhgrant0 & ~n21579;
  assign n21581 = ~n21347 & ~n21580;
  assign n21582 = ~n3281 & ~n21581;
  assign n21583 = ~n3950 & ~n21582;
  assign n21584 = ~n3378 & ~n21583;
  assign n21585 = ~n21576 & ~n21584;
  assign n21586 = n3492 & ~n21585;
  assign n21587 = ~n3493 & ~n21586;
  assign n21588 = n3485 & ~n21587;
  assign n21589 = ~n3486 & ~n21588;
  assign n21590 = ~n3476 & ~n21589;
  assign n21591 = ~n21383 & ~n21572;
  assign n21592 = ~n3281 & ~n21591;
  assign n21593 = ~n3281 & ~n21592;
  assign n21594 = n3378 & ~n21593;
  assign n21595 = ~controllable_hmaster0 & ~n11732;
  assign n21596 = ~n21412 & ~n21595;
  assign n21597 = ~controllable_hmaster1 & ~n21596;
  assign n21598 = ~n21411 & ~n21597;
  assign n21599 = i_hbusreq3 & ~n21598;
  assign n21600 = ~n6947 & ~n21433;
  assign n21601 = ~controllable_hmaster0 & ~n21600;
  assign n21602 = ~n21419 & ~n21601;
  assign n21603 = ~controllable_hmaster1 & ~n21602;
  assign n21604 = ~n21418 & ~n21603;
  assign n21605 = ~i_hbusreq3 & ~n21604;
  assign n21606 = ~n21599 & ~n21605;
  assign n21607 = ~controllable_hmaster2 & ~n21606;
  assign n21608 = ~n21410 & ~n21607;
  assign n21609 = ~controllable_hgrant3 & ~n21608;
  assign n21610 = ~n21338 & ~n21609;
  assign n21611 = controllable_nhgrant0 & ~n21610;
  assign n21612 = ~n21461 & ~n21611;
  assign n21613 = ~n3281 & ~n21612;
  assign n21614 = ~n4089 & ~n21613;
  assign n21615 = ~n3378 & ~n21614;
  assign n21616 = ~n21594 & ~n21615;
  assign n21617 = n3492 & ~n21616;
  assign n21618 = ~n21290 & ~n21617;
  assign n21619 = n3485 & ~n21618;
  assign n21620 = ~n21289 & ~n21619;
  assign n21621 = n3476 & ~n21620;
  assign n21622 = ~n21590 & ~n21621;
  assign n21623 = n3374 & ~n21622;
  assign n21624 = ~n21296 & ~n21623;
  assign n21625 = n3655 & ~n21624;
  assign n21626 = ~controllable_hmaster0 & ~n9595;
  assign n21627 = ~controllable_hmaster1 & ~n21626;
  assign n21628 = ~controllable_hmaster1 & ~n21627;
  assign n21629 = i_hbusreq3 & ~n21628;
  assign n21630 = ~controllable_hmaster0 & ~n9609;
  assign n21631 = ~controllable_hmaster1 & ~n21630;
  assign n21632 = ~controllable_hmaster1 & ~n21631;
  assign n21633 = ~i_hbusreq3 & ~n21632;
  assign n21634 = ~n21629 & ~n21633;
  assign n21635 = ~controllable_hmaster2 & ~n21634;
  assign n21636 = ~controllable_hmaster2 & ~n21635;
  assign n21637 = ~controllable_hgrant3 & ~n21636;
  assign n21638 = ~n21304 & ~n21637;
  assign n21639 = controllable_nhgrant0 & ~n21638;
  assign n21640 = ~n21332 & ~n21639;
  assign n21641 = ~n3281 & ~n21640;
  assign n21642 = ~n3281 & ~n21641;
  assign n21643 = n3378 & ~n21642;
  assign n21644 = ~n21339 & ~n21635;
  assign n21645 = ~controllable_hgrant3 & ~n21644;
  assign n21646 = ~n21338 & ~n21645;
  assign n21647 = controllable_nhgrant0 & ~n21646;
  assign n21648 = ~n21347 & ~n21647;
  assign n21649 = ~n3281 & ~n21648;
  assign n21650 = ~n3950 & ~n21649;
  assign n21651 = ~n3378 & ~n21650;
  assign n21652 = ~n21643 & ~n21651;
  assign n21653 = n3492 & ~n21652;
  assign n21654 = ~n3493 & ~n21653;
  assign n21655 = n3485 & ~n21654;
  assign n21656 = ~n3486 & ~n21655;
  assign n21657 = ~n3476 & ~n21656;
  assign n21658 = ~n21383 & ~n21639;
  assign n21659 = ~n3281 & ~n21658;
  assign n21660 = ~n3281 & ~n21659;
  assign n21661 = n3378 & ~n21660;
  assign n21662 = ~controllable_hmaster0 & ~n11802;
  assign n21663 = ~n21412 & ~n21662;
  assign n21664 = ~controllable_hmaster1 & ~n21663;
  assign n21665 = ~n21411 & ~n21664;
  assign n21666 = i_hbusreq3 & ~n21665;
  assign n21667 = ~n6947 & ~n21530;
  assign n21668 = ~controllable_hmaster0 & ~n21667;
  assign n21669 = ~n21419 & ~n21668;
  assign n21670 = ~controllable_hmaster1 & ~n21669;
  assign n21671 = ~n21418 & ~n21670;
  assign n21672 = ~i_hbusreq3 & ~n21671;
  assign n21673 = ~n21666 & ~n21672;
  assign n21674 = ~controllable_hmaster2 & ~n21673;
  assign n21675 = ~n21410 & ~n21674;
  assign n21676 = ~controllable_hgrant3 & ~n21675;
  assign n21677 = ~n21338 & ~n21676;
  assign n21678 = controllable_nhgrant0 & ~n21677;
  assign n21679 = ~n21461 & ~n21678;
  assign n21680 = ~n3281 & ~n21679;
  assign n21681 = ~n4089 & ~n21680;
  assign n21682 = ~n3378 & ~n21681;
  assign n21683 = ~n21661 & ~n21682;
  assign n21684 = n3492 & ~n21683;
  assign n21685 = ~n21290 & ~n21684;
  assign n21686 = n3485 & ~n21685;
  assign n21687 = ~n21289 & ~n21686;
  assign n21688 = n3476 & ~n21687;
  assign n21689 = ~n21657 & ~n21688;
  assign n21690 = n3374 & ~n21689;
  assign n21691 = ~n21296 & ~n21690;
  assign n21692 = ~n3655 & ~n21691;
  assign n21693 = ~n21625 & ~n21692;
  assign n21694 = ~n3652 & ~n21693;
  assign n21695 = ~n21558 & ~n21694;
  assign n21696 = ~n3368 & ~n21695;
  assign n21697 = ~controllable_hmaster2 & ~n3824;
  assign n21698 = ~controllable_hmaster2 & ~n21697;
  assign n21699 = controllable_hgrant3 & ~n21698;
  assign n21700 = ~controllable_hmaster2 & ~n21307;
  assign n21701 = ~controllable_hmaster2 & ~n21700;
  assign n21702 = ~controllable_hgrant3 & ~n21701;
  assign n21703 = ~n21699 & ~n21702;
  assign n21704 = controllable_nhgrant0 & ~n21703;
  assign n21705 = ~controllable_hmaster0 & ~n9847;
  assign n21706 = ~controllable_hmaster1 & ~n21705;
  assign n21707 = ~controllable_hmaster1 & ~n21706;
  assign n21708 = ~controllable_hmaster2 & ~n21707;
  assign n21709 = ~controllable_hmaster2 & ~n21708;
  assign n21710 = ~controllable_hgrant3 & ~n21709;
  assign n21711 = ~n21699 & ~n21710;
  assign n21712 = ~controllable_nhgrant0 & ~n21711;
  assign n21713 = ~n21704 & ~n21712;
  assign n21714 = ~n3281 & ~n21713;
  assign n21715 = ~n3281 & ~n21714;
  assign n21716 = n3492 & ~n21715;
  assign n21717 = n3492 & ~n21716;
  assign n21718 = n3485 & ~n21717;
  assign n21719 = n3485 & ~n21718;
  assign n21720 = ~n3476 & ~n21719;
  assign n21721 = ~n3485 & ~n21260;
  assign n21722 = ~n3492 & ~n21260;
  assign n21723 = i_hlock0 & ~n3551;
  assign n21724 = ~i_hlock0 & ~n14838;
  assign n21725 = ~n21723 & ~n21724;
  assign n21726 = ~controllable_hgrant4 & ~n21725;
  assign n21727 = ~controllable_hgrant4 & ~n21726;
  assign n21728 = ~controllable_hgrant2 & ~n21727;
  assign n21729 = ~controllable_hgrant2 & ~n21728;
  assign n21730 = controllable_hmaster2 & ~n21729;
  assign n21731 = controllable_hmaster1 & ~n21729;
  assign n21732 = controllable_hmaster0 & ~n21729;
  assign n21733 = ~n10224 & ~n21732;
  assign n21734 = ~controllable_hmaster1 & ~n21733;
  assign n21735 = ~n21731 & ~n21734;
  assign n21736 = ~controllable_hmaster2 & ~n21735;
  assign n21737 = ~n21730 & ~n21736;
  assign n21738 = ~controllable_hgrant3 & ~n21737;
  assign n21739 = ~n21699 & ~n21738;
  assign n21740 = ~controllable_nhgrant0 & ~n21739;
  assign n21741 = ~n21704 & ~n21740;
  assign n21742 = ~n3281 & ~n21741;
  assign n21743 = ~n3281 & ~n21742;
  assign n21744 = n3492 & ~n21743;
  assign n21745 = ~n21722 & ~n21744;
  assign n21746 = n3485 & ~n21745;
  assign n21747 = ~n21721 & ~n21746;
  assign n21748 = n3476 & ~n21747;
  assign n21749 = ~n21720 & ~n21748;
  assign n21750 = n3374 & ~n21749;
  assign n21751 = n3374 & ~n21750;
  assign n21752 = n3655 & ~n21751;
  assign n21753 = ~controllable_hmaster0 & ~n10337;
  assign n21754 = ~controllable_hmaster1 & ~n21753;
  assign n21755 = ~controllable_hmaster1 & ~n21754;
  assign n21756 = ~controllable_hmaster2 & ~n21755;
  assign n21757 = ~controllable_hmaster2 & ~n21756;
  assign n21758 = ~controllable_hgrant3 & ~n21757;
  assign n21759 = ~n21699 & ~n21758;
  assign n21760 = controllable_nhgrant0 & ~n21759;
  assign n21761 = ~n21712 & ~n21760;
  assign n21762 = ~n3281 & ~n21761;
  assign n21763 = ~n3281 & ~n21762;
  assign n21764 = n3492 & ~n21763;
  assign n21765 = n3492 & ~n21764;
  assign n21766 = n3485 & ~n21765;
  assign n21767 = n3485 & ~n21766;
  assign n21768 = ~n3476 & ~n21767;
  assign n21769 = ~n21740 & ~n21760;
  assign n21770 = ~n3281 & ~n21769;
  assign n21771 = ~n3281 & ~n21770;
  assign n21772 = n3492 & ~n21771;
  assign n21773 = ~n21722 & ~n21772;
  assign n21774 = n3485 & ~n21773;
  assign n21775 = ~n21721 & ~n21774;
  assign n21776 = n3476 & ~n21775;
  assign n21777 = ~n21768 & ~n21776;
  assign n21778 = n3374 & ~n21777;
  assign n21779 = n3374 & ~n21778;
  assign n21780 = ~n3655 & ~n21779;
  assign n21781 = ~n21752 & ~n21780;
  assign n21782 = n3652 & ~n21781;
  assign n21783 = ~controllable_hmaster0 & ~n10775;
  assign n21784 = ~controllable_hmaster1 & ~n21783;
  assign n21785 = ~controllable_hmaster1 & ~n21784;
  assign n21786 = ~controllable_hmaster2 & ~n21785;
  assign n21787 = ~controllable_hmaster2 & ~n21786;
  assign n21788 = ~controllable_hgrant3 & ~n21787;
  assign n21789 = ~n21699 & ~n21788;
  assign n21790 = controllable_nhgrant0 & ~n21789;
  assign n21791 = ~n21712 & ~n21790;
  assign n21792 = ~n3281 & ~n21791;
  assign n21793 = ~n3281 & ~n21792;
  assign n21794 = n3492 & ~n21793;
  assign n21795 = n3492 & ~n21794;
  assign n21796 = n3485 & ~n21795;
  assign n21797 = n3485 & ~n21796;
  assign n21798 = ~n3476 & ~n21797;
  assign n21799 = ~n21740 & ~n21790;
  assign n21800 = ~n3281 & ~n21799;
  assign n21801 = ~n3281 & ~n21800;
  assign n21802 = n3492 & ~n21801;
  assign n21803 = ~n21722 & ~n21802;
  assign n21804 = n3485 & ~n21803;
  assign n21805 = ~n21721 & ~n21804;
  assign n21806 = n3476 & ~n21805;
  assign n21807 = ~n21798 & ~n21806;
  assign n21808 = n3374 & ~n21807;
  assign n21809 = n3374 & ~n21808;
  assign n21810 = n3655 & ~n21809;
  assign n21811 = ~controllable_hmaster0 & ~n11210;
  assign n21812 = ~controllable_hmaster1 & ~n21811;
  assign n21813 = ~controllable_hmaster1 & ~n21812;
  assign n21814 = ~controllable_hmaster2 & ~n21813;
  assign n21815 = ~controllable_hmaster2 & ~n21814;
  assign n21816 = ~controllable_hgrant3 & ~n21815;
  assign n21817 = ~n21699 & ~n21816;
  assign n21818 = controllable_nhgrant0 & ~n21817;
  assign n21819 = ~n21712 & ~n21818;
  assign n21820 = ~n3281 & ~n21819;
  assign n21821 = ~n3281 & ~n21820;
  assign n21822 = n3492 & ~n21821;
  assign n21823 = n3492 & ~n21822;
  assign n21824 = n3485 & ~n21823;
  assign n21825 = n3485 & ~n21824;
  assign n21826 = ~n3476 & ~n21825;
  assign n21827 = ~n21740 & ~n21818;
  assign n21828 = ~n3281 & ~n21827;
  assign n21829 = ~n3281 & ~n21828;
  assign n21830 = n3492 & ~n21829;
  assign n21831 = ~n21722 & ~n21830;
  assign n21832 = n3485 & ~n21831;
  assign n21833 = ~n21721 & ~n21832;
  assign n21834 = n3476 & ~n21833;
  assign n21835 = ~n21826 & ~n21834;
  assign n21836 = n3374 & ~n21835;
  assign n21837 = n3374 & ~n21836;
  assign n21838 = ~n3655 & ~n21837;
  assign n21839 = ~n21810 & ~n21838;
  assign n21840 = ~n3652 & ~n21839;
  assign n21841 = ~n21782 & ~n21840;
  assign n21842 = n3368 & ~n21841;
  assign n21843 = ~n21696 & ~n21842;
  assign n21844 = ~n3362 & ~n21843;
  assign n21845 = ~n3362 & ~n21844;
  assign n21846 = ~n3359 & ~n21845;
  assign n21847 = ~n3359 & ~n21846;
  assign n21848 = n3356 & ~n21847;
  assign n21849 = n3378 & ~n21279;
  assign n21850 = ~n3767 & ~n5046;
  assign n21851 = ~controllable_hmaster1 & ~n21850;
  assign n21852 = ~n5045 & ~n21851;
  assign n21853 = ~i_hbusreq3 & ~n21852;
  assign n21854 = ~n5050 & ~n21853;
  assign n21855 = controllable_hmaster2 & ~n21854;
  assign n21856 = ~n5161 & ~n21855;
  assign n21857 = ~controllable_hgrant3 & ~n21856;
  assign n21858 = ~n8750 & ~n21857;
  assign n21859 = controllable_nhgrant0 & ~n21858;
  assign n21860 = ~n8785 & ~n21859;
  assign n21861 = ~n3281 & ~n21860;
  assign n21862 = ~n3783 & ~n21861;
  assign n21863 = ~n3378 & ~n21862;
  assign n21864 = ~n21849 & ~n21863;
  assign n21865 = n3492 & ~n21864;
  assign n21866 = ~n3631 & ~n21865;
  assign n21867 = n3485 & ~n21866;
  assign n21868 = ~n3630 & ~n21867;
  assign n21869 = ~n3476 & ~n21868;
  assign n21870 = ~n8309 & ~n21865;
  assign n21871 = n3485 & ~n21870;
  assign n21872 = ~n8639 & ~n21871;
  assign n21873 = n3476 & ~n21872;
  assign n21874 = ~n21869 & ~n21873;
  assign n21875 = ~n3374 & ~n21874;
  assign n21876 = ~controllable_hgrant4 & ~n3832;
  assign n21877 = ~n3873 & ~n21876;
  assign n21878 = ~i_hbusreq2 & ~n21877;
  assign n21879 = ~n12051 & ~n21878;
  assign n21880 = ~controllable_hgrant2 & ~n21879;
  assign n21881 = ~n3859 & ~n21880;
  assign n21882 = ~controllable_hmaster0 & ~n21881;
  assign n21883 = ~n3502 & ~n21882;
  assign n21884 = ~controllable_hmaster1 & ~n21883;
  assign n21885 = ~n3501 & ~n21884;
  assign n21886 = ~i_hbusreq3 & ~n21885;
  assign n21887 = ~n12050 & ~n21886;
  assign n21888 = controllable_hmaster2 & ~n21887;
  assign n21889 = ~n5303 & ~n8827;
  assign n21890 = ~controllable_hmaster1 & ~n21889;
  assign n21891 = ~n5293 & ~n21890;
  assign n21892 = i_hbusreq3 & ~n21891;
  assign n21893 = ~controllable_hgrant2 & ~n3834;
  assign n21894 = ~n5438 & ~n21893;
  assign n21895 = ~controllable_hmaster0 & ~n21894;
  assign n21896 = ~n4913 & ~n21895;
  assign n21897 = controllable_hmaster1 & ~n21896;
  assign n21898 = i_hlock0 & ~n5321;
  assign n21899 = ~i_hlock0 & ~n5298;
  assign n21900 = ~n21898 & ~n21899;
  assign n21901 = ~i_hbusreq0 & ~n21900;
  assign n21902 = ~n5316 & ~n21901;
  assign n21903 = ~i_hbusreq4 & ~n21902;
  assign n21904 = ~n5315 & ~n21903;
  assign n21905 = ~controllable_hgrant4 & ~n21904;
  assign n21906 = ~n3916 & ~n21905;
  assign n21907 = ~i_hbusreq2 & ~n21906;
  assign n21908 = ~n5314 & ~n21907;
  assign n21909 = ~controllable_hgrant2 & ~n21908;
  assign n21910 = ~n3859 & ~n21909;
  assign n21911 = controllable_hmaster0 & ~n21910;
  assign n21912 = ~n8876 & ~n21911;
  assign n21913 = ~controllable_hmaster1 & ~n21912;
  assign n21914 = ~n21897 & ~n21913;
  assign n21915 = ~i_hbusreq3 & ~n21914;
  assign n21916 = ~n21892 & ~n21915;
  assign n21917 = ~controllable_hmaster2 & ~n21916;
  assign n21918 = ~n21888 & ~n21917;
  assign n21919 = ~controllable_hgrant3 & ~n21918;
  assign n21920 = ~n8810 & ~n21919;
  assign n21921 = controllable_nhgrant0 & ~n21920;
  assign n21922 = ~n8902 & ~n21921;
  assign n21923 = ~n3281 & ~n21922;
  assign n21924 = ~n3950 & ~n21923;
  assign n21925 = n3378 & ~n21924;
  assign n21926 = ~n3502 & ~n12120;
  assign n21927 = ~controllable_hmaster1 & ~n21926;
  assign n21928 = ~n3501 & ~n21927;
  assign n21929 = ~i_hbusreq3 & ~n21928;
  assign n21930 = ~n12113 & ~n21929;
  assign n21931 = controllable_hmaster2 & ~n21930;
  assign n21932 = ~n5433 & ~n8827;
  assign n21933 = ~controllable_hmaster1 & ~n21932;
  assign n21934 = ~n5427 & ~n21933;
  assign n21935 = i_hbusreq3 & ~n21934;
  assign n21936 = ~n5460 & ~n8876;
  assign n21937 = ~controllable_hmaster1 & ~n21936;
  assign n21938 = ~n5442 & ~n21937;
  assign n21939 = ~i_hbusreq3 & ~n21938;
  assign n21940 = ~n21935 & ~n21939;
  assign n21941 = ~controllable_hmaster2 & ~n21940;
  assign n21942 = ~n21931 & ~n21941;
  assign n21943 = ~controllable_hgrant3 & ~n21942;
  assign n21944 = ~n8810 & ~n21943;
  assign n21945 = controllable_nhgrant0 & ~n21944;
  assign n21946 = ~n8902 & ~n21945;
  assign n21947 = ~n3281 & ~n21946;
  assign n21948 = ~n3950 & ~n21947;
  assign n21949 = ~n3378 & ~n21948;
  assign n21950 = ~n21925 & ~n21949;
  assign n21951 = n3492 & ~n21950;
  assign n21952 = ~n3631 & ~n21951;
  assign n21953 = n3485 & ~n21952;
  assign n21954 = ~n3630 & ~n21953;
  assign n21955 = ~n3476 & ~n21954;
  assign n21956 = ~n3392 & ~n8961;
  assign n21957 = i_hlock0 & ~n21956;
  assign n21958 = ~n3379 & ~n5889;
  assign n21959 = ~i_hlock0 & ~n21958;
  assign n21960 = ~n21957 & ~n21959;
  assign n21961 = ~i_hbusreq0 & ~n21960;
  assign n21962 = ~n5709 & ~n21961;
  assign n21963 = ~i_hbusreq4 & ~n21962;
  assign n21964 = ~n5708 & ~n21963;
  assign n21965 = ~controllable_hgrant4 & ~n21964;
  assign n21966 = ~n4064 & ~n21965;
  assign n21967 = ~i_hbusreq2 & ~n21966;
  assign n21968 = ~n12180 & ~n21967;
  assign n21969 = ~controllable_hgrant2 & ~n21968;
  assign n21970 = ~n5862 & ~n21969;
  assign n21971 = ~controllable_hmaster0 & ~n21970;
  assign n21972 = ~n8957 & ~n21971;
  assign n21973 = ~controllable_hmaster1 & ~n21972;
  assign n21974 = ~n8956 & ~n21973;
  assign n21975 = ~i_hbusreq3 & ~n21974;
  assign n21976 = ~n12171 & ~n21975;
  assign n21977 = controllable_hmaster2 & ~n21976;
  assign n21978 = ~n5701 & ~n8992;
  assign n21979 = ~controllable_hmaster1 & ~n21978;
  assign n21980 = ~n5690 & ~n21979;
  assign n21981 = i_hbusreq3 & ~n21980;
  assign n21982 = ~n5863 & ~n21965;
  assign n21983 = ~i_hbusreq2 & ~n21982;
  assign n21984 = ~n5707 & ~n21983;
  assign n21985 = ~controllable_hgrant2 & ~n21984;
  assign n21986 = ~n5862 & ~n21985;
  assign n21987 = controllable_hmaster0 & ~n21986;
  assign n21988 = ~n5950 & ~n21985;
  assign n21989 = ~controllable_hmaster0 & ~n21988;
  assign n21990 = ~n21987 & ~n21989;
  assign n21991 = controllable_hmaster1 & ~n21990;
  assign n21992 = ~n3392 & ~n9014;
  assign n21993 = i_hlock0 & ~n21992;
  assign n21994 = ~n3379 & ~n5966;
  assign n21995 = ~i_hlock0 & ~n21994;
  assign n21996 = ~n21993 & ~n21995;
  assign n21997 = ~i_hbusreq0 & ~n21996;
  assign n21998 = ~n5729 & ~n21997;
  assign n21999 = ~i_hbusreq4 & ~n21998;
  assign n22000 = ~n5728 & ~n21999;
  assign n22001 = ~controllable_hgrant4 & ~n22000;
  assign n22002 = ~n5863 & ~n22001;
  assign n22003 = ~i_hbusreq2 & ~n22002;
  assign n22004 = ~n5727 & ~n22003;
  assign n22005 = ~controllable_hgrant2 & ~n22004;
  assign n22006 = ~n5862 & ~n22005;
  assign n22007 = controllable_hmaster0 & ~n22006;
  assign n22008 = ~n9044 & ~n22007;
  assign n22009 = ~controllable_hmaster1 & ~n22008;
  assign n22010 = ~n21991 & ~n22009;
  assign n22011 = ~i_hbusreq3 & ~n22010;
  assign n22012 = ~n21981 & ~n22011;
  assign n22013 = ~controllable_hmaster2 & ~n22012;
  assign n22014 = ~n21977 & ~n22013;
  assign n22015 = ~controllable_hgrant3 & ~n22014;
  assign n22016 = ~n8935 & ~n22015;
  assign n22017 = controllable_nhgrant0 & ~n22016;
  assign n22018 = ~n9096 & ~n22017;
  assign n22019 = ~n3281 & ~n22018;
  assign n22020 = ~n4089 & ~n22019;
  assign n22021 = n3378 & ~n22020;
  assign n22022 = ~n3920 & ~n8961;
  assign n22023 = i_hlock0 & ~n22022;
  assign n22024 = ~n5937 & ~n22023;
  assign n22025 = ~i_hbusreq0 & ~n22024;
  assign n22026 = ~n5933 & ~n22025;
  assign n22027 = ~i_hbusreq4 & ~n22026;
  assign n22028 = ~n5932 & ~n22027;
  assign n22029 = ~controllable_hgrant4 & ~n22028;
  assign n22030 = ~n4064 & ~n22029;
  assign n22031 = ~i_hbusreq2 & ~n22030;
  assign n22032 = ~n12262 & ~n22031;
  assign n22033 = ~controllable_hgrant2 & ~n22032;
  assign n22034 = ~n5862 & ~n22033;
  assign n22035 = ~controllable_hmaster0 & ~n22034;
  assign n22036 = ~n8957 & ~n22035;
  assign n22037 = ~controllable_hmaster1 & ~n22036;
  assign n22038 = ~n8956 & ~n22037;
  assign n22039 = ~i_hbusreq3 & ~n22038;
  assign n22040 = ~n12261 & ~n22039;
  assign n22041 = controllable_hmaster2 & ~n22040;
  assign n22042 = ~n5925 & ~n8992;
  assign n22043 = ~controllable_hmaster1 & ~n22042;
  assign n22044 = ~n5919 & ~n22043;
  assign n22045 = i_hbusreq3 & ~n22044;
  assign n22046 = ~n5863 & ~n22029;
  assign n22047 = ~i_hbusreq2 & ~n22046;
  assign n22048 = ~n5931 & ~n22047;
  assign n22049 = ~controllable_hgrant2 & ~n22048;
  assign n22050 = ~n5862 & ~n22049;
  assign n22051 = controllable_hmaster0 & ~n22050;
  assign n22052 = ~n5950 & ~n22049;
  assign n22053 = ~controllable_hmaster0 & ~n22052;
  assign n22054 = ~n22051 & ~n22053;
  assign n22055 = controllable_hmaster1 & ~n22054;
  assign n22056 = ~n3920 & ~n9014;
  assign n22057 = i_hlock0 & ~n22056;
  assign n22058 = ~n5968 & ~n22057;
  assign n22059 = ~i_hbusreq0 & ~n22058;
  assign n22060 = ~n5957 & ~n22059;
  assign n22061 = ~i_hbusreq4 & ~n22060;
  assign n22062 = ~n5956 & ~n22061;
  assign n22063 = ~controllable_hgrant4 & ~n22062;
  assign n22064 = ~n5863 & ~n22063;
  assign n22065 = ~i_hbusreq2 & ~n22064;
  assign n22066 = ~n5955 & ~n22065;
  assign n22067 = ~controllable_hgrant2 & ~n22066;
  assign n22068 = ~n5862 & ~n22067;
  assign n22069 = controllable_hmaster0 & ~n22068;
  assign n22070 = ~n9044 & ~n22069;
  assign n22071 = ~controllable_hmaster1 & ~n22070;
  assign n22072 = ~n22055 & ~n22071;
  assign n22073 = ~i_hbusreq3 & ~n22072;
  assign n22074 = ~n22045 & ~n22073;
  assign n22075 = ~controllable_hmaster2 & ~n22074;
  assign n22076 = ~n22041 & ~n22075;
  assign n22077 = ~controllable_hgrant3 & ~n22076;
  assign n22078 = ~n8935 & ~n22077;
  assign n22079 = controllable_nhgrant0 & ~n22078;
  assign n22080 = ~n9096 & ~n22079;
  assign n22081 = ~n3281 & ~n22080;
  assign n22082 = ~n4089 & ~n22081;
  assign n22083 = ~n3378 & ~n22082;
  assign n22084 = ~n22021 & ~n22083;
  assign n22085 = n3492 & ~n22084;
  assign n22086 = ~n8309 & ~n22085;
  assign n22087 = n3485 & ~n22086;
  assign n22088 = ~n8639 & ~n22087;
  assign n22089 = n3476 & ~n22088;
  assign n22090 = ~n21955 & ~n22089;
  assign n22091 = n3374 & ~n22090;
  assign n22092 = ~n21875 & ~n22091;
  assign n22093 = n3655 & ~n22092;
  assign n22094 = ~n3767 & ~n6105;
  assign n22095 = ~controllable_hmaster1 & ~n22094;
  assign n22096 = ~n6104 & ~n22095;
  assign n22097 = ~i_hbusreq3 & ~n22096;
  assign n22098 = ~n6109 & ~n22097;
  assign n22099 = controllable_hmaster2 & ~n22098;
  assign n22100 = ~n6188 & ~n22099;
  assign n22101 = ~controllable_hgrant3 & ~n22100;
  assign n22102 = ~n8750 & ~n22101;
  assign n22103 = controllable_nhgrant0 & ~n22102;
  assign n22104 = ~n8785 & ~n22103;
  assign n22105 = ~n3281 & ~n22104;
  assign n22106 = ~n3783 & ~n22105;
  assign n22107 = ~n3378 & ~n22106;
  assign n22108 = ~n21849 & ~n22107;
  assign n22109 = n3492 & ~n22108;
  assign n22110 = ~n3631 & ~n22109;
  assign n22111 = n3485 & ~n22110;
  assign n22112 = ~n3630 & ~n22111;
  assign n22113 = ~n3476 & ~n22112;
  assign n22114 = ~n8309 & ~n22109;
  assign n22115 = n3485 & ~n22114;
  assign n22116 = ~n8639 & ~n22115;
  assign n22117 = n3476 & ~n22116;
  assign n22118 = ~n22113 & ~n22117;
  assign n22119 = ~n3374 & ~n22118;
  assign n22120 = ~n5303 & ~n9175;
  assign n22121 = ~controllable_hmaster1 & ~n22120;
  assign n22122 = ~n5293 & ~n22121;
  assign n22123 = i_hbusreq3 & ~n22122;
  assign n22124 = ~n9226 & ~n21911;
  assign n22125 = ~controllable_hmaster1 & ~n22124;
  assign n22126 = ~n21897 & ~n22125;
  assign n22127 = ~i_hbusreq3 & ~n22126;
  assign n22128 = ~n22123 & ~n22127;
  assign n22129 = ~controllable_hmaster2 & ~n22128;
  assign n22130 = ~n21888 & ~n22129;
  assign n22131 = ~controllable_hgrant3 & ~n22130;
  assign n22132 = ~n8810 & ~n22131;
  assign n22133 = controllable_nhgrant0 & ~n22132;
  assign n22134 = ~n8902 & ~n22133;
  assign n22135 = ~n3281 & ~n22134;
  assign n22136 = ~n3950 & ~n22135;
  assign n22137 = n3378 & ~n22136;
  assign n22138 = ~n6217 & ~n12347;
  assign n22139 = ~controllable_hmaster1 & ~n22138;
  assign n22140 = ~n6216 & ~n22139;
  assign n22141 = ~i_hbusreq3 & ~n22140;
  assign n22142 = ~n12340 & ~n22141;
  assign n22143 = controllable_hmaster2 & ~n22142;
  assign n22144 = ~n6268 & ~n9175;
  assign n22145 = ~controllable_hmaster1 & ~n22144;
  assign n22146 = ~n6258 & ~n22145;
  assign n22147 = i_hbusreq3 & ~n22146;
  assign n22148 = ~n6321 & ~n9226;
  assign n22149 = ~controllable_hmaster1 & ~n22148;
  assign n22150 = ~n6297 & ~n22149;
  assign n22151 = ~i_hbusreq3 & ~n22150;
  assign n22152 = ~n22147 & ~n22151;
  assign n22153 = ~controllable_hmaster2 & ~n22152;
  assign n22154 = ~n22143 & ~n22153;
  assign n22155 = ~controllable_hgrant3 & ~n22154;
  assign n22156 = ~n8810 & ~n22155;
  assign n22157 = controllable_nhgrant0 & ~n22156;
  assign n22158 = ~n8902 & ~n22157;
  assign n22159 = ~n3281 & ~n22158;
  assign n22160 = ~n3950 & ~n22159;
  assign n22161 = ~n3378 & ~n22160;
  assign n22162 = ~n22137 & ~n22161;
  assign n22163 = n3492 & ~n22162;
  assign n22164 = ~n3631 & ~n22163;
  assign n22165 = n3485 & ~n22164;
  assign n22166 = ~n3630 & ~n22165;
  assign n22167 = ~n3476 & ~n22166;
  assign n22168 = ~controllable_hmaster0 & ~n12380;
  assign n22169 = ~n5701 & ~n22168;
  assign n22170 = ~controllable_hmaster1 & ~n22169;
  assign n22171 = ~n5690 & ~n22170;
  assign n22172 = i_hbusreq3 & ~n22171;
  assign n22173 = ~n8961 & ~n9212;
  assign n22174 = i_hlock0 & ~n22173;
  assign n22175 = ~n4180 & ~n5889;
  assign n22176 = ~i_hlock0 & ~n22175;
  assign n22177 = ~n22174 & ~n22176;
  assign n22178 = ~i_hbusreq0 & ~n22177;
  assign n22179 = ~n6370 & ~n22178;
  assign n22180 = ~i_hbusreq4 & ~n22179;
  assign n22181 = ~n6369 & ~n22180;
  assign n22182 = ~controllable_hgrant4 & ~n22181;
  assign n22183 = ~n5982 & ~n22182;
  assign n22184 = ~i_hbusreq2 & ~n22183;
  assign n22185 = ~n12386 & ~n22184;
  assign n22186 = ~controllable_hgrant2 & ~n22185;
  assign n22187 = ~n5981 & ~n22186;
  assign n22188 = ~controllable_hmaster0 & ~n22187;
  assign n22189 = ~n22007 & ~n22188;
  assign n22190 = ~controllable_hmaster1 & ~n22189;
  assign n22191 = ~n21991 & ~n22190;
  assign n22192 = ~i_hbusreq3 & ~n22191;
  assign n22193 = ~n22172 & ~n22192;
  assign n22194 = ~controllable_hmaster2 & ~n22193;
  assign n22195 = ~n21977 & ~n22194;
  assign n22196 = ~controllable_hgrant3 & ~n22195;
  assign n22197 = ~n8935 & ~n22196;
  assign n22198 = controllable_nhgrant0 & ~n22197;
  assign n22199 = ~n9096 & ~n22198;
  assign n22200 = ~n3281 & ~n22199;
  assign n22201 = ~n4089 & ~n22200;
  assign n22202 = n3378 & ~n22201;
  assign n22203 = ~n4180 & ~n9262;
  assign n22204 = i_hlock0 & ~n22203;
  assign n22205 = ~n6427 & ~n22204;
  assign n22206 = ~i_hbusreq0 & ~n22205;
  assign n22207 = ~n6419 & ~n22206;
  assign n22208 = ~i_hbusreq4 & ~n22207;
  assign n22209 = ~n6418 & ~n22208;
  assign n22210 = ~controllable_hgrant4 & ~n22209;
  assign n22211 = ~n8937 & ~n22210;
  assign n22212 = ~i_hbusreq2 & ~n22211;
  assign n22213 = ~n6417 & ~n22212;
  assign n22214 = ~controllable_hgrant2 & ~n22213;
  assign n22215 = ~n8936 & ~n22214;
  assign n22216 = controllable_hmaster1 & ~n22215;
  assign n22217 = controllable_hmaster0 & ~n22215;
  assign n22218 = ~n6278 & ~n9279;
  assign n22219 = i_hlock0 & ~n22218;
  assign n22220 = ~n6492 & ~n22219;
  assign n22221 = ~i_hbusreq0 & ~n22220;
  assign n22222 = ~n6488 & ~n22221;
  assign n22223 = ~i_hbusreq4 & ~n22222;
  assign n22224 = ~n6487 & ~n22223;
  assign n22225 = ~controllable_hgrant4 & ~n22224;
  assign n22226 = ~n4064 & ~n22225;
  assign n22227 = ~i_hbusreq2 & ~n22226;
  assign n22228 = ~n12415 & ~n22227;
  assign n22229 = ~controllable_hgrant2 & ~n22228;
  assign n22230 = ~n5862 & ~n22229;
  assign n22231 = ~controllable_hmaster0 & ~n22230;
  assign n22232 = ~n22217 & ~n22231;
  assign n22233 = ~controllable_hmaster1 & ~n22232;
  assign n22234 = ~n22216 & ~n22233;
  assign n22235 = ~i_hbusreq3 & ~n22234;
  assign n22236 = ~n12414 & ~n22235;
  assign n22237 = controllable_hmaster2 & ~n22236;
  assign n22238 = ~n6480 & ~n9310;
  assign n22239 = ~controllable_hmaster1 & ~n22238;
  assign n22240 = ~n6473 & ~n22239;
  assign n22241 = i_hbusreq3 & ~n22240;
  assign n22242 = ~n5863 & ~n22225;
  assign n22243 = ~i_hbusreq2 & ~n22242;
  assign n22244 = ~n6486 & ~n22243;
  assign n22245 = ~controllable_hgrant2 & ~n22244;
  assign n22246 = ~n5862 & ~n22245;
  assign n22247 = controllable_hmaster0 & ~n22246;
  assign n22248 = ~n5950 & ~n22245;
  assign n22249 = ~controllable_hmaster0 & ~n22248;
  assign n22250 = ~n22247 & ~n22249;
  assign n22251 = controllable_hmaster1 & ~n22250;
  assign n22252 = ~n6306 & ~n9330;
  assign n22253 = i_hlock0 & ~n22252;
  assign n22254 = ~n6522 & ~n22253;
  assign n22255 = ~i_hbusreq0 & ~n22254;
  assign n22256 = ~n6511 & ~n22255;
  assign n22257 = ~i_hbusreq4 & ~n22256;
  assign n22258 = ~n6510 & ~n22257;
  assign n22259 = ~controllable_hgrant4 & n22258;
  assign n22260 = ~n5863 & ~n22259;
  assign n22261 = ~i_hbusreq2 & ~n22260;
  assign n22262 = ~n6509 & ~n22261;
  assign n22263 = ~controllable_hgrant2 & ~n22262;
  assign n22264 = ~n5862 & ~n22263;
  assign n22265 = controllable_hmaster0 & ~n22264;
  assign n22266 = ~n9360 & ~n22265;
  assign n22267 = ~controllable_hmaster1 & ~n22266;
  assign n22268 = ~n22251 & ~n22267;
  assign n22269 = ~i_hbusreq3 & ~n22268;
  assign n22270 = ~n22241 & ~n22269;
  assign n22271 = ~controllable_hmaster2 & ~n22270;
  assign n22272 = ~n22237 & ~n22271;
  assign n22273 = ~controllable_hgrant3 & ~n22272;
  assign n22274 = ~n8935 & ~n22273;
  assign n22275 = controllable_nhgrant0 & ~n22274;
  assign n22276 = ~n9096 & ~n22275;
  assign n22277 = ~n3281 & ~n22276;
  assign n22278 = ~n4089 & ~n22277;
  assign n22279 = ~n3378 & ~n22278;
  assign n22280 = ~n22202 & ~n22279;
  assign n22281 = n3492 & ~n22280;
  assign n22282 = ~n8309 & ~n22281;
  assign n22283 = n3485 & ~n22282;
  assign n22284 = ~n8639 & ~n22283;
  assign n22285 = n3476 & ~n22284;
  assign n22286 = ~n22167 & ~n22285;
  assign n22287 = n3374 & ~n22286;
  assign n22288 = ~n22119 & ~n22287;
  assign n22289 = ~n3655 & ~n22288;
  assign n22290 = ~n22093 & ~n22289;
  assign n22291 = n3652 & ~n22290;
  assign n22292 = ~n3767 & ~n6577;
  assign n22293 = ~controllable_hmaster1 & ~n22292;
  assign n22294 = ~n6576 & ~n22293;
  assign n22295 = ~i_hbusreq3 & ~n22294;
  assign n22296 = ~n6581 & ~n22295;
  assign n22297 = controllable_hmaster2 & ~n22296;
  assign n22298 = ~n6657 & ~n22297;
  assign n22299 = ~controllable_hgrant3 & ~n22298;
  assign n22300 = ~n8750 & ~n22299;
  assign n22301 = controllable_nhgrant0 & ~n22300;
  assign n22302 = ~n8785 & ~n22301;
  assign n22303 = ~n3281 & ~n22302;
  assign n22304 = ~n3783 & ~n22303;
  assign n22305 = ~n3378 & ~n22304;
  assign n22306 = ~n21849 & ~n22305;
  assign n22307 = n3492 & ~n22306;
  assign n22308 = ~n3631 & ~n22307;
  assign n22309 = n3485 & ~n22308;
  assign n22310 = ~n3630 & ~n22309;
  assign n22311 = ~n3476 & ~n22310;
  assign n22312 = ~n8309 & ~n22307;
  assign n22313 = n3485 & ~n22312;
  assign n22314 = ~n8639 & ~n22313;
  assign n22315 = n3476 & ~n22314;
  assign n22316 = ~n22311 & ~n22315;
  assign n22317 = ~n3374 & ~n22316;
  assign n22318 = ~n5303 & ~n9441;
  assign n22319 = ~controllable_hmaster1 & ~n22318;
  assign n22320 = ~n5293 & ~n22319;
  assign n22321 = i_hbusreq3 & ~n22320;
  assign n22322 = ~n9455 & ~n21911;
  assign n22323 = ~controllable_hmaster1 & ~n22322;
  assign n22324 = ~n21897 & ~n22323;
  assign n22325 = ~i_hbusreq3 & ~n22324;
  assign n22326 = ~n22321 & ~n22325;
  assign n22327 = ~controllable_hmaster2 & ~n22326;
  assign n22328 = ~n21888 & ~n22327;
  assign n22329 = ~controllable_hgrant3 & ~n22328;
  assign n22330 = ~n8810 & ~n22329;
  assign n22331 = controllable_nhgrant0 & ~n22330;
  assign n22332 = ~n8902 & ~n22331;
  assign n22333 = ~n3281 & ~n22332;
  assign n22334 = ~n3950 & ~n22333;
  assign n22335 = n3378 & ~n22334;
  assign n22336 = ~n6682 & ~n12495;
  assign n22337 = ~controllable_hmaster1 & ~n22336;
  assign n22338 = ~n6681 & ~n22337;
  assign n22339 = ~i_hbusreq3 & ~n22338;
  assign n22340 = ~n12493 & ~n22339;
  assign n22341 = controllable_hmaster2 & ~n22340;
  assign n22342 = ~n6703 & ~n9441;
  assign n22343 = ~controllable_hmaster1 & ~n22342;
  assign n22344 = ~n6701 & ~n22343;
  assign n22345 = i_hbusreq3 & ~n22344;
  assign n22346 = ~n6716 & ~n9455;
  assign n22347 = ~controllable_hmaster1 & ~n22346;
  assign n22348 = ~n6714 & ~n22347;
  assign n22349 = ~i_hbusreq3 & ~n22348;
  assign n22350 = ~n22345 & ~n22349;
  assign n22351 = ~controllable_hmaster2 & ~n22350;
  assign n22352 = ~n22341 & ~n22351;
  assign n22353 = ~controllable_hgrant3 & ~n22352;
  assign n22354 = ~n8810 & ~n22353;
  assign n22355 = controllable_nhgrant0 & ~n22354;
  assign n22356 = ~n8902 & ~n22355;
  assign n22357 = ~n3281 & ~n22356;
  assign n22358 = ~n3950 & ~n22357;
  assign n22359 = ~n3378 & ~n22358;
  assign n22360 = ~n22335 & ~n22359;
  assign n22361 = n3492 & ~n22360;
  assign n22362 = ~n3631 & ~n22361;
  assign n22363 = n3485 & ~n22362;
  assign n22364 = ~n3630 & ~n22363;
  assign n22365 = ~n3476 & ~n22364;
  assign n22366 = ~controllable_hmaster0 & ~n12526;
  assign n22367 = ~n5701 & ~n22366;
  assign n22368 = ~controllable_hmaster1 & ~n22367;
  assign n22369 = ~n5690 & ~n22368;
  assign n22370 = i_hbusreq3 & ~n22369;
  assign n22371 = ~n4031 & ~n5464;
  assign n22372 = i_hlock0 & ~n22371;
  assign n22373 = ~i_hlock0 & ~n5759;
  assign n22374 = ~n22372 & ~n22373;
  assign n22375 = ~i_hbusreq0 & ~n22374;
  assign n22376 = ~n5771 & ~n22375;
  assign n22377 = ~i_hbusreq4 & ~n22376;
  assign n22378 = ~n5770 & ~n22377;
  assign n22379 = ~controllable_hgrant4 & ~n22378;
  assign n22380 = ~n5462 & ~n22379;
  assign n22381 = ~i_hbusreq2 & ~n22380;
  assign n22382 = ~n5769 & ~n22381;
  assign n22383 = controllable_hgrant2 & ~n22382;
  assign n22384 = ~n9042 & ~n22383;
  assign n22385 = ~controllable_hmaster0 & ~n22384;
  assign n22386 = ~n22007 & ~n22385;
  assign n22387 = ~controllable_hmaster1 & ~n22386;
  assign n22388 = ~n21991 & ~n22387;
  assign n22389 = ~i_hbusreq3 & ~n22388;
  assign n22390 = ~n22370 & ~n22389;
  assign n22391 = ~controllable_hmaster2 & ~n22390;
  assign n22392 = ~n21977 & ~n22391;
  assign n22393 = ~controllable_hgrant3 & ~n22392;
  assign n22394 = ~n8935 & ~n22393;
  assign n22395 = controllable_nhgrant0 & ~n22394;
  assign n22396 = ~n9096 & ~n22395;
  assign n22397 = ~n3281 & ~n22396;
  assign n22398 = ~n4089 & ~n22397;
  assign n22399 = n3378 & ~n22398;
  assign n22400 = ~n3904 & ~n6018;
  assign n22401 = i_hlock0 & ~n22400;
  assign n22402 = ~n6021 & ~n22401;
  assign n22403 = ~i_hbusreq0 & ~n22402;
  assign n22404 = ~n6016 & ~n22403;
  assign n22405 = ~i_hbusreq4 & ~n22404;
  assign n22406 = ~n6015 & ~n22405;
  assign n22407 = ~controllable_hgrant4 & ~n22406;
  assign n22408 = ~n3411 & ~n22407;
  assign n22409 = ~i_hbusreq2 & ~n22408;
  assign n22410 = ~n6014 & ~n22409;
  assign n22411 = controllable_hgrant2 & ~n22410;
  assign n22412 = ~n8954 & ~n22411;
  assign n22413 = controllable_hmaster1 & ~n22412;
  assign n22414 = controllable_hmaster0 & ~n22412;
  assign n22415 = ~n6772 & ~n22033;
  assign n22416 = ~controllable_hmaster0 & ~n22415;
  assign n22417 = ~n22414 & ~n22416;
  assign n22418 = ~controllable_hmaster1 & ~n22417;
  assign n22419 = ~n22413 & ~n22418;
  assign n22420 = ~i_hbusreq3 & ~n22419;
  assign n22421 = ~n12553 & ~n22420;
  assign n22422 = controllable_hmaster2 & ~n22421;
  assign n22423 = ~n6792 & ~n9503;
  assign n22424 = ~controllable_hmaster1 & ~n22423;
  assign n22425 = ~n6790 & ~n22424;
  assign n22426 = i_hbusreq3 & ~n22425;
  assign n22427 = ~n6772 & ~n22049;
  assign n22428 = controllable_hmaster0 & ~n22427;
  assign n22429 = ~n6813 & ~n22049;
  assign n22430 = ~controllable_hmaster0 & ~n22429;
  assign n22431 = ~n22428 & ~n22430;
  assign n22432 = controllable_hmaster1 & ~n22431;
  assign n22433 = ~n6772 & ~n22067;
  assign n22434 = controllable_hmaster0 & ~n22433;
  assign n22435 = ~n9517 & ~n22434;
  assign n22436 = ~controllable_hmaster1 & ~n22435;
  assign n22437 = ~n22432 & ~n22436;
  assign n22438 = ~i_hbusreq3 & ~n22437;
  assign n22439 = ~n22426 & ~n22438;
  assign n22440 = ~controllable_hmaster2 & ~n22439;
  assign n22441 = ~n22422 & ~n22440;
  assign n22442 = ~controllable_hgrant3 & ~n22441;
  assign n22443 = ~n8935 & ~n22442;
  assign n22444 = controllable_nhgrant0 & ~n22443;
  assign n22445 = ~n9096 & ~n22444;
  assign n22446 = ~n3281 & ~n22445;
  assign n22447 = ~n4089 & ~n22446;
  assign n22448 = ~n3378 & ~n22447;
  assign n22449 = ~n22399 & ~n22448;
  assign n22450 = n3492 & ~n22449;
  assign n22451 = ~n8309 & ~n22450;
  assign n22452 = n3485 & ~n22451;
  assign n22453 = ~n8639 & ~n22452;
  assign n22454 = n3476 & ~n22453;
  assign n22455 = ~n22365 & ~n22454;
  assign n22456 = n3374 & ~n22455;
  assign n22457 = ~n22317 & ~n22456;
  assign n22458 = n3655 & ~n22457;
  assign n22459 = ~n3767 & ~n6860;
  assign n22460 = ~controllable_hmaster1 & ~n22459;
  assign n22461 = ~n6859 & ~n22460;
  assign n22462 = ~i_hbusreq3 & ~n22461;
  assign n22463 = ~n6864 & ~n22462;
  assign n22464 = controllable_hmaster2 & ~n22463;
  assign n22465 = ~n6887 & ~n22464;
  assign n22466 = ~controllable_hgrant3 & ~n22465;
  assign n22467 = ~n8750 & ~n22466;
  assign n22468 = controllable_nhgrant0 & ~n22467;
  assign n22469 = ~n8785 & ~n22468;
  assign n22470 = ~n3281 & ~n22469;
  assign n22471 = ~n3783 & ~n22470;
  assign n22472 = ~n3378 & ~n22471;
  assign n22473 = ~n21849 & ~n22472;
  assign n22474 = n3492 & ~n22473;
  assign n22475 = ~n3631 & ~n22474;
  assign n22476 = n3485 & ~n22475;
  assign n22477 = ~n3630 & ~n22476;
  assign n22478 = ~n3476 & ~n22477;
  assign n22479 = ~n8309 & ~n22474;
  assign n22480 = n3485 & ~n22479;
  assign n22481 = ~n8639 & ~n22480;
  assign n22482 = n3476 & ~n22481;
  assign n22483 = ~n22478 & ~n22482;
  assign n22484 = ~n3374 & ~n22483;
  assign n22485 = ~n5303 & ~n9595;
  assign n22486 = ~controllable_hmaster1 & ~n22485;
  assign n22487 = ~n5293 & ~n22486;
  assign n22488 = i_hbusreq3 & ~n22487;
  assign n22489 = ~n9609 & ~n21911;
  assign n22490 = ~controllable_hmaster1 & ~n22489;
  assign n22491 = ~n21897 & ~n22490;
  assign n22492 = ~i_hbusreq3 & ~n22491;
  assign n22493 = ~n22488 & ~n22492;
  assign n22494 = ~controllable_hmaster2 & ~n22493;
  assign n22495 = ~n21888 & ~n22494;
  assign n22496 = ~controllable_hgrant3 & ~n22495;
  assign n22497 = ~n8810 & ~n22496;
  assign n22498 = controllable_nhgrant0 & ~n22497;
  assign n22499 = ~n8902 & ~n22498;
  assign n22500 = ~n3281 & ~n22499;
  assign n22501 = ~n3950 & ~n22500;
  assign n22502 = n3378 & ~n22501;
  assign n22503 = ~n6912 & ~n12623;
  assign n22504 = ~controllable_hmaster1 & ~n22503;
  assign n22505 = ~n6911 & ~n22504;
  assign n22506 = ~i_hbusreq3 & ~n22505;
  assign n22507 = ~n12621 & ~n22506;
  assign n22508 = controllable_hmaster2 & ~n22507;
  assign n22509 = ~n6933 & ~n9595;
  assign n22510 = ~controllable_hmaster1 & ~n22509;
  assign n22511 = ~n6931 & ~n22510;
  assign n22512 = i_hbusreq3 & ~n22511;
  assign n22513 = ~n6946 & ~n9609;
  assign n22514 = ~controllable_hmaster1 & ~n22513;
  assign n22515 = ~n6944 & ~n22514;
  assign n22516 = ~i_hbusreq3 & ~n22515;
  assign n22517 = ~n22512 & ~n22516;
  assign n22518 = ~controllable_hmaster2 & ~n22517;
  assign n22519 = ~n22508 & ~n22518;
  assign n22520 = ~controllable_hgrant3 & ~n22519;
  assign n22521 = ~n8810 & ~n22520;
  assign n22522 = controllable_nhgrant0 & ~n22521;
  assign n22523 = ~n8902 & ~n22522;
  assign n22524 = ~n3281 & ~n22523;
  assign n22525 = ~n3950 & ~n22524;
  assign n22526 = ~n3378 & ~n22525;
  assign n22527 = ~n22502 & ~n22526;
  assign n22528 = n3492 & ~n22527;
  assign n22529 = ~n3631 & ~n22528;
  assign n22530 = n3485 & ~n22529;
  assign n22531 = ~n3630 & ~n22530;
  assign n22532 = ~n3476 & ~n22531;
  assign n22533 = ~controllable_hmaster0 & ~n12654;
  assign n22534 = ~n5701 & ~n22533;
  assign n22535 = ~controllable_hmaster1 & ~n22534;
  assign n22536 = ~n5690 & ~n22535;
  assign n22537 = i_hbusreq3 & ~n22536;
  assign n22538 = ~n22186 & ~n22383;
  assign n22539 = ~controllable_hmaster0 & ~n22538;
  assign n22540 = ~n22007 & ~n22539;
  assign n22541 = ~controllable_hmaster1 & ~n22540;
  assign n22542 = ~n21991 & ~n22541;
  assign n22543 = ~i_hbusreq3 & ~n22542;
  assign n22544 = ~n22537 & ~n22543;
  assign n22545 = ~controllable_hmaster2 & ~n22544;
  assign n22546 = ~n21977 & ~n22545;
  assign n22547 = ~controllable_hgrant3 & ~n22546;
  assign n22548 = ~n8935 & ~n22547;
  assign n22549 = controllable_nhgrant0 & ~n22548;
  assign n22550 = ~n9096 & ~n22549;
  assign n22551 = ~n3281 & ~n22550;
  assign n22552 = ~n4089 & ~n22551;
  assign n22553 = n3378 & ~n22552;
  assign n22554 = ~n22214 & ~n22411;
  assign n22555 = controllable_hmaster1 & ~n22554;
  assign n22556 = controllable_hmaster0 & ~n22554;
  assign n22557 = ~n6772 & ~n22229;
  assign n22558 = ~controllable_hmaster0 & ~n22557;
  assign n22559 = ~n22556 & ~n22558;
  assign n22560 = ~controllable_hmaster1 & ~n22559;
  assign n22561 = ~n22555 & ~n22560;
  assign n22562 = ~i_hbusreq3 & ~n22561;
  assign n22563 = ~n12681 & ~n22562;
  assign n22564 = controllable_hmaster2 & ~n22563;
  assign n22565 = ~n7019 & ~n9655;
  assign n22566 = ~controllable_hmaster1 & ~n22565;
  assign n22567 = ~n7017 & ~n22566;
  assign n22568 = i_hbusreq3 & ~n22567;
  assign n22569 = ~n6772 & ~n22245;
  assign n22570 = controllable_hmaster0 & ~n22569;
  assign n22571 = ~n6813 & ~n22245;
  assign n22572 = ~controllable_hmaster0 & ~n22571;
  assign n22573 = ~n22570 & ~n22572;
  assign n22574 = controllable_hmaster1 & ~n22573;
  assign n22575 = ~n6772 & ~n22263;
  assign n22576 = controllable_hmaster0 & ~n22575;
  assign n22577 = ~n9669 & ~n22576;
  assign n22578 = ~controllable_hmaster1 & ~n22577;
  assign n22579 = ~n22574 & ~n22578;
  assign n22580 = ~i_hbusreq3 & ~n22579;
  assign n22581 = ~n22568 & ~n22580;
  assign n22582 = ~controllable_hmaster2 & ~n22581;
  assign n22583 = ~n22564 & ~n22582;
  assign n22584 = ~controllable_hgrant3 & ~n22583;
  assign n22585 = ~n8935 & ~n22584;
  assign n22586 = controllable_nhgrant0 & ~n22585;
  assign n22587 = ~n9096 & ~n22586;
  assign n22588 = ~n3281 & ~n22587;
  assign n22589 = ~n4089 & ~n22588;
  assign n22590 = ~n3378 & ~n22589;
  assign n22591 = ~n22553 & ~n22590;
  assign n22592 = n3492 & ~n22591;
  assign n22593 = ~n8309 & ~n22592;
  assign n22594 = n3485 & ~n22593;
  assign n22595 = ~n8639 & ~n22594;
  assign n22596 = n3476 & ~n22595;
  assign n22597 = ~n22532 & ~n22596;
  assign n22598 = n3374 & ~n22597;
  assign n22599 = ~n22484 & ~n22598;
  assign n22600 = ~n3655 & ~n22599;
  assign n22601 = ~n22458 & ~n22600;
  assign n22602 = ~n3652 & ~n22601;
  assign n22603 = ~n22291 & ~n22602;
  assign n22604 = ~n3368 & ~n22603;
  assign n22605 = controllable_hmaster1 & ~n9779;
  assign n22606 = ~controllable_hmaster1 & ~n11838;
  assign n22607 = ~n22605 & ~n22606;
  assign n22608 = ~i_hbusreq3 & ~n22607;
  assign n22609 = ~n7067 & ~n22608;
  assign n22610 = controllable_hmaster2 & ~n22609;
  assign n22611 = controllable_hmaster2 & ~n22610;
  assign n22612 = ~controllable_hgrant3 & ~n22611;
  assign n22613 = ~n9708 & ~n22612;
  assign n22614 = controllable_nhgrant0 & ~n22613;
  assign n22615 = ~n9753 & ~n22614;
  assign n22616 = ~n3281 & ~n22615;
  assign n22617 = ~n3281 & ~n22616;
  assign n22618 = n3378 & ~n22617;
  assign n22619 = ~n4541 & ~n5038;
  assign n22620 = ~i_hready & ~n22619;
  assign n22621 = ~n9710 & ~n22620;
  assign n22622 = i_hlock0 & ~n22621;
  assign n22623 = ~n5058 & ~n22622;
  assign n22624 = ~i_hbusreq0 & ~n22623;
  assign n22625 = ~n5053 & ~n22624;
  assign n22626 = ~i_hbusreq4 & ~n22625;
  assign n22627 = ~n5052 & ~n22626;
  assign n22628 = ~controllable_hgrant4 & ~n22627;
  assign n22629 = ~n4617 & ~n22628;
  assign n22630 = ~i_hbusreq2 & ~n22629;
  assign n22631 = ~n5051 & ~n22630;
  assign n22632 = ~controllable_hgrant2 & ~n22631;
  assign n22633 = ~n4562 & ~n22632;
  assign n22634 = controllable_hmaster1 & ~n22633;
  assign n22635 = controllable_hmaster0 & ~n22633;
  assign n22636 = controllable_hmaster0 & ~n22635;
  assign n22637 = ~controllable_hmaster1 & ~n22636;
  assign n22638 = ~n22634 & ~n22637;
  assign n22639 = ~i_hbusreq3 & ~n22638;
  assign n22640 = ~n7094 & ~n22639;
  assign n22641 = controllable_hmaster2 & ~n22640;
  assign n22642 = controllable_hmaster2 & ~n22641;
  assign n22643 = ~controllable_hgrant3 & ~n22642;
  assign n22644 = ~n9708 & ~n22643;
  assign n22645 = controllable_nhgrant0 & ~n22644;
  assign n22646 = ~n9753 & ~n22645;
  assign n22647 = ~n3281 & ~n22646;
  assign n22648 = ~n3281 & ~n22647;
  assign n22649 = ~n3378 & ~n22648;
  assign n22650 = ~n22618 & ~n22649;
  assign n22651 = n3492 & ~n22650;
  assign n22652 = n3492 & ~n22651;
  assign n22653 = n3485 & ~n22652;
  assign n22654 = n3485 & ~n22653;
  assign n22655 = ~n3374 & ~n22654;
  assign n22656 = ~controllable_hgrant4 & ~n4550;
  assign n22657 = ~n4575 & ~n22656;
  assign n22658 = ~i_hbusreq2 & ~n22657;
  assign n22659 = ~n12051 & ~n22658;
  assign n22660 = ~controllable_hgrant2 & ~n22659;
  assign n22661 = ~n4562 & ~n22660;
  assign n22662 = ~controllable_hmaster0 & ~n22661;
  assign n22663 = ~n9780 & ~n22662;
  assign n22664 = ~controllable_hmaster1 & ~n22663;
  assign n22665 = ~n22605 & ~n22664;
  assign n22666 = ~i_hbusreq3 & ~n22665;
  assign n22667 = ~n12735 & ~n22666;
  assign n22668 = controllable_hmaster2 & ~n22667;
  assign n22669 = ~controllable_hgrant2 & ~n4552;
  assign n22670 = ~n9803 & ~n22669;
  assign n22671 = ~controllable_hmaster0 & ~n22670;
  assign n22672 = ~n9700 & ~n22671;
  assign n22673 = controllable_hmaster1 & ~n22672;
  assign n22674 = ~n4543 & ~n9812;
  assign n22675 = i_hlock0 & ~n22674;
  assign n22676 = ~n21899 & ~n22675;
  assign n22677 = ~i_hbusreq0 & ~n22676;
  assign n22678 = ~n5316 & ~n22677;
  assign n22679 = ~i_hbusreq4 & ~n22678;
  assign n22680 = ~n5315 & ~n22679;
  assign n22681 = ~controllable_hgrant4 & ~n22680;
  assign n22682 = ~n4617 & ~n22681;
  assign n22683 = ~i_hbusreq2 & ~n22682;
  assign n22684 = ~n5314 & ~n22683;
  assign n22685 = ~controllable_hgrant2 & ~n22684;
  assign n22686 = ~n4562 & ~n22685;
  assign n22687 = controllable_hmaster0 & ~n22686;
  assign n22688 = ~n8827 & ~n22687;
  assign n22689 = ~controllable_hmaster1 & ~n22688;
  assign n22690 = ~n22673 & ~n22689;
  assign n22691 = ~i_hbusreq3 & ~n22690;
  assign n22692 = ~n21892 & ~n22691;
  assign n22693 = ~controllable_hmaster2 & ~n22692;
  assign n22694 = ~n22668 & ~n22693;
  assign n22695 = ~controllable_hgrant3 & ~n22694;
  assign n22696 = ~n9790 & ~n22695;
  assign n22697 = controllable_nhgrant0 & ~n22696;
  assign n22698 = ~n9861 & ~n22697;
  assign n22699 = ~n3281 & ~n22698;
  assign n22700 = ~n3281 & ~n22699;
  assign n22701 = n3378 & ~n22700;
  assign n22702 = ~n3903 & ~n4541;
  assign n22703 = ~i_hready & ~n22702;
  assign n22704 = ~i_hready & ~n22703;
  assign n22705 = i_hlock0 & ~n22704;
  assign n22706 = ~n3923 & ~n22705;
  assign n22707 = ~i_hbusreq0 & ~n22706;
  assign n22708 = ~n3918 & ~n22707;
  assign n22709 = ~i_hbusreq4 & ~n22708;
  assign n22710 = ~n3917 & ~n22709;
  assign n22711 = ~controllable_hgrant4 & ~n22710;
  assign n22712 = ~n4575 & ~n22711;
  assign n22713 = ~i_hbusreq2 & ~n22712;
  assign n22714 = ~n12114 & ~n22713;
  assign n22715 = ~controllable_hgrant2 & ~n22714;
  assign n22716 = ~n4562 & ~n22715;
  assign n22717 = ~controllable_hmaster0 & ~n22716;
  assign n22718 = ~n22635 & ~n22717;
  assign n22719 = ~controllable_hmaster1 & ~n22718;
  assign n22720 = ~n22634 & ~n22719;
  assign n22721 = ~i_hbusreq3 & ~n22720;
  assign n22722 = ~n12789 & ~n22721;
  assign n22723 = controllable_hmaster2 & ~n22722;
  assign n22724 = ~n4617 & ~n22711;
  assign n22725 = ~i_hbusreq2 & ~n22724;
  assign n22726 = ~n3915 & ~n22725;
  assign n22727 = ~controllable_hgrant2 & ~n22726;
  assign n22728 = ~n4562 & ~n22727;
  assign n22729 = controllable_hmaster0 & ~n22728;
  assign n22730 = ~n9803 & ~n22727;
  assign n22731 = ~controllable_hmaster0 & ~n22730;
  assign n22732 = ~n22729 & ~n22731;
  assign n22733 = controllable_hmaster1 & ~n22732;
  assign n22734 = ~n9812 & ~n22703;
  assign n22735 = i_hlock0 & ~n22734;
  assign n22736 = ~n5448 & ~n22735;
  assign n22737 = ~i_hbusreq0 & ~n22736;
  assign n22738 = ~n5445 & ~n22737;
  assign n22739 = ~i_hbusreq4 & ~n22738;
  assign n22740 = ~n5444 & ~n22739;
  assign n22741 = ~controllable_hgrant4 & ~n22740;
  assign n22742 = ~n4617 & ~n22741;
  assign n22743 = ~i_hbusreq2 & ~n22742;
  assign n22744 = ~n5443 & ~n22743;
  assign n22745 = ~controllable_hgrant2 & ~n22744;
  assign n22746 = ~n4562 & ~n22745;
  assign n22747 = controllable_hmaster0 & ~n22746;
  assign n22748 = ~n8827 & ~n22747;
  assign n22749 = ~controllable_hmaster1 & ~n22748;
  assign n22750 = ~n22733 & ~n22749;
  assign n22751 = ~i_hbusreq3 & ~n22750;
  assign n22752 = ~n21935 & ~n22751;
  assign n22753 = ~controllable_hmaster2 & ~n22752;
  assign n22754 = ~n22723 & ~n22753;
  assign n22755 = ~controllable_hgrant3 & ~n22754;
  assign n22756 = ~n9790 & ~n22755;
  assign n22757 = controllable_nhgrant0 & ~n22756;
  assign n22758 = ~n9861 & ~n22757;
  assign n22759 = ~n3281 & ~n22758;
  assign n22760 = ~n3281 & ~n22759;
  assign n22761 = ~n3378 & ~n22760;
  assign n22762 = ~n22701 & ~n22761;
  assign n22763 = n3492 & ~n22762;
  assign n22764 = n3492 & ~n22763;
  assign n22765 = n3485 & ~n22764;
  assign n22766 = n3485 & ~n22765;
  assign n22767 = ~n3476 & ~n22766;
  assign n22768 = ~n5885 & ~n7272;
  assign n22769 = ~controllable_ndecide & ~n22768;
  assign n22770 = ~controllable_ndecide & ~n22769;
  assign n22771 = i_hready & ~n22770;
  assign n22772 = ~n4543 & ~n22771;
  assign n22773 = i_hlock0 & ~n22772;
  assign n22774 = ~i_hlock0 & ~n7244;
  assign n22775 = ~n22773 & ~n22774;
  assign n22776 = ~i_hbusreq0 & ~n22775;
  assign n22777 = ~n7271 & ~n22776;
  assign n22778 = ~i_hbusreq4 & ~n22777;
  assign n22779 = ~n7270 & ~n22778;
  assign n22780 = ~controllable_hgrant4 & ~n22779;
  assign n22781 = ~n10112 & ~n22780;
  assign n22782 = ~i_hbusreq2 & ~n22781;
  assign n22783 = ~n7264 & ~n22782;
  assign n22784 = ~controllable_hgrant2 & ~n22783;
  assign n22785 = ~n10111 & ~n22784;
  assign n22786 = controllable_hmaster1 & ~n22785;
  assign n22787 = controllable_hmaster0 & ~n22785;
  assign n22788 = ~n4543 & ~n7253;
  assign n22789 = i_hlock0 & ~n22788;
  assign n22790 = ~i_hlock0 & ~n7321;
  assign n22791 = ~n22789 & ~n22790;
  assign n22792 = ~i_hbusreq0 & ~n22791;
  assign n22793 = ~n7347 & ~n22792;
  assign n22794 = ~i_hbusreq4 & ~n22793;
  assign n22795 = ~n7346 & ~n22794;
  assign n22796 = ~controllable_hgrant4 & ~n22795;
  assign n22797 = ~n4667 & ~n22796;
  assign n22798 = ~i_hbusreq2 & ~n22797;
  assign n22799 = ~n12872 & ~n22798;
  assign n22800 = ~controllable_hgrant2 & ~n22799;
  assign n22801 = ~n10111 & ~n22800;
  assign n22802 = ~controllable_hmaster0 & ~n22801;
  assign n22803 = ~n22787 & ~n22802;
  assign n22804 = ~controllable_hmaster1 & ~n22803;
  assign n22805 = ~n22786 & ~n22804;
  assign n22806 = ~i_hbusreq3 & ~n22805;
  assign n22807 = ~n12864 & ~n22806;
  assign n22808 = controllable_hmaster2 & ~n22807;
  assign n22809 = ~controllable_hmaster0 & ~n12887;
  assign n22810 = ~n7339 & ~n22809;
  assign n22811 = ~controllable_hmaster1 & ~n22810;
  assign n22812 = ~n7330 & ~n22811;
  assign n22813 = i_hbusreq3 & ~n22812;
  assign n22814 = ~n10112 & ~n22796;
  assign n22815 = ~i_hbusreq2 & ~n22814;
  assign n22816 = ~n7345 & ~n22815;
  assign n22817 = ~controllable_hgrant2 & ~n22816;
  assign n22818 = ~n10111 & ~n22817;
  assign n22819 = controllable_hmaster0 & ~n22818;
  assign n22820 = ~n10152 & ~n22817;
  assign n22821 = ~controllable_hmaster0 & ~n22820;
  assign n22822 = ~n22819 & ~n22821;
  assign n22823 = controllable_hmaster1 & ~n22822;
  assign n22824 = ~n7367 & ~n10157;
  assign n22825 = ~controllable_ndecide & n22824;
  assign n22826 = ~controllable_ndecide & ~n22825;
  assign n22827 = i_hready & ~n22826;
  assign n22828 = ~n4543 & ~n22827;
  assign n22829 = i_hlock0 & ~n22828;
  assign n22830 = ~i_hlock0 & ~n7334;
  assign n22831 = ~n22829 & ~n22830;
  assign n22832 = ~i_hbusreq0 & ~n22831;
  assign n22833 = ~n7366 & ~n22832;
  assign n22834 = ~i_hbusreq4 & ~n22833;
  assign n22835 = ~n7365 & ~n22834;
  assign n22836 = ~controllable_hgrant4 & ~n22835;
  assign n22837 = ~n10112 & ~n22836;
  assign n22838 = ~i_hbusreq2 & ~n22837;
  assign n22839 = ~n7364 & ~n22838;
  assign n22840 = ~controllable_hgrant2 & ~n22839;
  assign n22841 = ~n10111 & ~n22840;
  assign n22842 = controllable_hmaster0 & ~n22841;
  assign n22843 = ~n22809 & ~n22842;
  assign n22844 = ~controllable_hmaster1 & ~n22843;
  assign n22845 = ~n22823 & ~n22844;
  assign n22846 = ~i_hbusreq3 & ~n22845;
  assign n22847 = ~n22813 & ~n22846;
  assign n22848 = ~controllable_hmaster2 & ~n22847;
  assign n22849 = ~n22808 & ~n22848;
  assign n22850 = ~controllable_hgrant3 & ~n22849;
  assign n22851 = ~n10110 & ~n22850;
  assign n22852 = controllable_nhgrant0 & ~n22851;
  assign n22853 = ~n10240 & ~n22852;
  assign n22854 = ~n3281 & ~n22853;
  assign n22855 = ~n3281 & ~n22854;
  assign n22856 = n3378 & ~n22855;
  assign n22857 = ~n5038 & ~n22769;
  assign n22858 = i_hready & ~n22857;
  assign n22859 = ~n22620 & ~n22858;
  assign n22860 = i_hlock0 & ~n22859;
  assign n22861 = ~n7493 & ~n22860;
  assign n22862 = ~i_hbusreq0 & ~n22861;
  assign n22863 = ~n7488 & ~n22862;
  assign n22864 = ~i_hbusreq4 & ~n22863;
  assign n22865 = ~n7487 & ~n22864;
  assign n22866 = ~controllable_hgrant4 & ~n22865;
  assign n22867 = ~n10112 & ~n22866;
  assign n22868 = ~i_hbusreq2 & ~n22867;
  assign n22869 = ~n7479 & ~n22868;
  assign n22870 = ~controllable_hgrant2 & ~n22869;
  assign n22871 = ~n10111 & ~n22870;
  assign n22872 = controllable_hmaster1 & ~n22871;
  assign n22873 = controllable_hmaster0 & ~n22871;
  assign n22874 = ~n7468 & ~n22703;
  assign n22875 = i_hlock0 & ~n22874;
  assign n22876 = ~n7562 & ~n22875;
  assign n22877 = ~i_hbusreq0 & ~n22876;
  assign n22878 = ~n7559 & ~n22877;
  assign n22879 = ~i_hbusreq4 & ~n22878;
  assign n22880 = ~n7558 & ~n22879;
  assign n22881 = ~controllable_hgrant4 & ~n22880;
  assign n22882 = ~n4667 & ~n22881;
  assign n22883 = ~i_hbusreq2 & ~n22882;
  assign n22884 = ~n12990 & ~n22883;
  assign n22885 = ~controllable_hgrant2 & ~n22884;
  assign n22886 = ~n10111 & ~n22885;
  assign n22887 = ~controllable_hmaster0 & ~n22886;
  assign n22888 = ~n22873 & ~n22887;
  assign n22889 = ~controllable_hmaster1 & ~n22888;
  assign n22890 = ~n22872 & ~n22889;
  assign n22891 = ~i_hbusreq3 & ~n22890;
  assign n22892 = ~n12982 & ~n22891;
  assign n22893 = controllable_hmaster2 & ~n22892;
  assign n22894 = ~controllable_hmaster0 & ~n13005;
  assign n22895 = ~n7551 & ~n22894;
  assign n22896 = ~controllable_hmaster1 & ~n22895;
  assign n22897 = ~n7543 & ~n22896;
  assign n22898 = i_hbusreq3 & ~n22897;
  assign n22899 = ~n10112 & ~n22881;
  assign n22900 = ~i_hbusreq2 & ~n22899;
  assign n22901 = ~n7557 & ~n22900;
  assign n22902 = ~controllable_hgrant2 & ~n22901;
  assign n22903 = ~n10111 & ~n22902;
  assign n22904 = controllable_hmaster0 & ~n22903;
  assign n22905 = ~n10152 & ~n22902;
  assign n22906 = ~controllable_hmaster0 & ~n22905;
  assign n22907 = ~n22904 & ~n22906;
  assign n22908 = controllable_hmaster1 & ~n22907;
  assign n22909 = ~n3903 & ~n22825;
  assign n22910 = i_hready & ~n22909;
  assign n22911 = ~n22703 & ~n22910;
  assign n22912 = i_hlock0 & ~n22911;
  assign n22913 = ~n7586 & ~n22912;
  assign n22914 = ~i_hbusreq0 & ~n22913;
  assign n22915 = ~n7581 & ~n22914;
  assign n22916 = ~i_hbusreq4 & ~n22915;
  assign n22917 = ~n7580 & ~n22916;
  assign n22918 = ~controllable_hgrant4 & ~n22917;
  assign n22919 = ~n10112 & ~n22918;
  assign n22920 = ~i_hbusreq2 & ~n22919;
  assign n22921 = ~n7579 & ~n22920;
  assign n22922 = ~controllable_hgrant2 & ~n22921;
  assign n22923 = ~n10111 & ~n22922;
  assign n22924 = controllable_hmaster0 & ~n22923;
  assign n22925 = ~n22894 & ~n22924;
  assign n22926 = ~controllable_hmaster1 & ~n22925;
  assign n22927 = ~n22908 & ~n22926;
  assign n22928 = ~i_hbusreq3 & ~n22927;
  assign n22929 = ~n22898 & ~n22928;
  assign n22930 = ~controllable_hmaster2 & ~n22929;
  assign n22931 = ~n22893 & ~n22930;
  assign n22932 = ~controllable_hgrant3 & ~n22931;
  assign n22933 = ~n10110 & ~n22932;
  assign n22934 = controllable_nhgrant0 & ~n22933;
  assign n22935 = ~n10240 & ~n22934;
  assign n22936 = ~n3281 & ~n22935;
  assign n22937 = ~n3281 & ~n22936;
  assign n22938 = ~n3378 & ~n22937;
  assign n22939 = ~n22856 & ~n22938;
  assign n22940 = n3492 & ~n22939;
  assign n22941 = ~n21722 & ~n22940;
  assign n22942 = n3485 & ~n22941;
  assign n22943 = ~n21721 & ~n22942;
  assign n22944 = n3476 & ~n22943;
  assign n22945 = ~n22767 & ~n22944;
  assign n22946 = n3374 & ~n22945;
  assign n22947 = ~n22655 & ~n22946;
  assign n22948 = n3655 & ~n22947;
  assign n22949 = ~n4541 & ~n6097;
  assign n22950 = ~i_hready & ~n22949;
  assign n22951 = ~n9710 & ~n22950;
  assign n22952 = i_hlock0 & ~n22951;
  assign n22953 = ~n6117 & ~n22952;
  assign n22954 = ~i_hbusreq0 & ~n22953;
  assign n22955 = ~n6112 & ~n22954;
  assign n22956 = ~i_hbusreq4 & ~n22955;
  assign n22957 = ~n6111 & ~n22956;
  assign n22958 = ~controllable_hgrant4 & ~n22957;
  assign n22959 = ~n4617 & ~n22958;
  assign n22960 = ~i_hbusreq2 & ~n22959;
  assign n22961 = ~n6110 & ~n22960;
  assign n22962 = ~controllable_hgrant2 & ~n22961;
  assign n22963 = ~n4562 & ~n22962;
  assign n22964 = controllable_hmaster1 & ~n22963;
  assign n22965 = controllable_hmaster0 & ~n22963;
  assign n22966 = controllable_hmaster0 & ~n22965;
  assign n22967 = ~controllable_hmaster1 & ~n22966;
  assign n22968 = ~n22964 & ~n22967;
  assign n22969 = ~i_hbusreq3 & ~n22968;
  assign n22970 = ~n7686 & ~n22969;
  assign n22971 = controllable_hmaster2 & ~n22970;
  assign n22972 = controllable_hmaster2 & ~n22971;
  assign n22973 = ~controllable_hgrant3 & ~n22972;
  assign n22974 = ~n9708 & ~n22973;
  assign n22975 = controllable_nhgrant0 & ~n22974;
  assign n22976 = ~n9753 & ~n22975;
  assign n22977 = ~n3281 & ~n22976;
  assign n22978 = ~n3281 & ~n22977;
  assign n22979 = ~n3378 & ~n22978;
  assign n22980 = ~n22618 & ~n22979;
  assign n22981 = n3492 & ~n22980;
  assign n22982 = n3492 & ~n22981;
  assign n22983 = n3485 & ~n22982;
  assign n22984 = n3485 & ~n22983;
  assign n22985 = ~n3374 & ~n22984;
  assign n22986 = ~n5303 & ~n10337;
  assign n22987 = ~controllable_hmaster1 & ~n22986;
  assign n22988 = ~n5293 & ~n22987;
  assign n22989 = i_hbusreq3 & ~n22988;
  assign n22990 = ~n10337 & ~n22687;
  assign n22991 = ~controllable_hmaster1 & ~n22990;
  assign n22992 = ~n22673 & ~n22991;
  assign n22993 = ~i_hbusreq3 & ~n22992;
  assign n22994 = ~n22989 & ~n22993;
  assign n22995 = ~controllable_hmaster2 & ~n22994;
  assign n22996 = ~n22668 & ~n22995;
  assign n22997 = ~controllable_hgrant3 & ~n22996;
  assign n22998 = ~n9790 & ~n22997;
  assign n22999 = controllable_nhgrant0 & ~n22998;
  assign n23000 = ~n9861 & ~n22999;
  assign n23001 = ~n3281 & ~n23000;
  assign n23002 = ~n3281 & ~n23001;
  assign n23003 = n3378 & ~n23002;
  assign n23004 = ~n4541 & ~n6247;
  assign n23005 = ~i_hready & ~n23004;
  assign n23006 = ~i_hready & ~n23005;
  assign n23007 = i_hlock0 & ~n23006;
  assign n23008 = ~n6281 & ~n23007;
  assign n23009 = ~i_hbusreq0 & ~n23008;
  assign n23010 = ~n6276 & ~n23009;
  assign n23011 = ~i_hbusreq4 & ~n23010;
  assign n23012 = ~n6275 & ~n23011;
  assign n23013 = ~controllable_hgrant4 & ~n23012;
  assign n23014 = ~n4575 & ~n23013;
  assign n23015 = ~i_hbusreq2 & ~n23014;
  assign n23016 = ~n12341 & ~n23015;
  assign n23017 = ~controllable_hgrant2 & ~n23016;
  assign n23018 = ~n4562 & ~n23017;
  assign n23019 = ~controllable_hmaster0 & ~n23018;
  assign n23020 = ~n22965 & ~n23019;
  assign n23021 = ~controllable_hmaster1 & ~n23020;
  assign n23022 = ~n22964 & ~n23021;
  assign n23023 = ~i_hbusreq3 & ~n23022;
  assign n23024 = ~n13100 & ~n23023;
  assign n23025 = controllable_hmaster2 & ~n23024;
  assign n23026 = ~n6268 & ~n10337;
  assign n23027 = ~controllable_hmaster1 & ~n23026;
  assign n23028 = ~n6258 & ~n23027;
  assign n23029 = i_hbusreq3 & ~n23028;
  assign n23030 = ~n4617 & ~n23013;
  assign n23031 = ~i_hbusreq2 & ~n23030;
  assign n23032 = ~n6274 & ~n23031;
  assign n23033 = ~controllable_hgrant2 & ~n23032;
  assign n23034 = ~n4562 & ~n23033;
  assign n23035 = controllable_hmaster0 & ~n23034;
  assign n23036 = ~n9803 & ~n23033;
  assign n23037 = ~controllable_hmaster0 & ~n23036;
  assign n23038 = ~n23035 & ~n23037;
  assign n23039 = controllable_hmaster1 & ~n23038;
  assign n23040 = ~n6260 & ~n10359;
  assign n23041 = ~i_hready & ~n23040;
  assign n23042 = ~n10358 & ~n23041;
  assign n23043 = i_hlock0 & ~n23042;
  assign n23044 = ~n6309 & ~n23043;
  assign n23045 = ~i_hbusreq0 & ~n23044;
  assign n23046 = ~n6300 & ~n23045;
  assign n23047 = ~i_hbusreq4 & ~n23046;
  assign n23048 = ~n6299 & ~n23047;
  assign n23049 = ~controllable_hgrant4 & n23048;
  assign n23050 = ~n4617 & ~n23049;
  assign n23051 = ~i_hbusreq2 & ~n23050;
  assign n23052 = ~n6298 & ~n23051;
  assign n23053 = ~controllable_hgrant2 & ~n23052;
  assign n23054 = ~n4562 & ~n23053;
  assign n23055 = controllable_hmaster0 & ~n23054;
  assign n23056 = ~n10337 & ~n23055;
  assign n23057 = ~controllable_hmaster1 & ~n23056;
  assign n23058 = ~n23039 & ~n23057;
  assign n23059 = ~i_hbusreq3 & ~n23058;
  assign n23060 = ~n23029 & ~n23059;
  assign n23061 = ~controllable_hmaster2 & ~n23060;
  assign n23062 = ~n23025 & ~n23061;
  assign n23063 = ~controllable_hgrant3 & ~n23062;
  assign n23064 = ~n9790 & ~n23063;
  assign n23065 = controllable_nhgrant0 & ~n23064;
  assign n23066 = ~n9861 & ~n23065;
  assign n23067 = ~n3281 & ~n23066;
  assign n23068 = ~n3281 & ~n23067;
  assign n23069 = ~n3378 & ~n23068;
  assign n23070 = ~n23003 & ~n23069;
  assign n23071 = n3492 & ~n23070;
  assign n23072 = n3492 & ~n23071;
  assign n23073 = n3485 & ~n23072;
  assign n23074 = n3485 & ~n23073;
  assign n23075 = ~n3476 & ~n23074;
  assign n23076 = ~controllable_hmaster0 & ~n13133;
  assign n23077 = ~n7339 & ~n23076;
  assign n23078 = ~controllable_hmaster1 & ~n23077;
  assign n23079 = ~n7330 & ~n23078;
  assign n23080 = i_hbusreq3 & ~n23079;
  assign n23081 = ~n22842 & ~n23076;
  assign n23082 = ~controllable_hmaster1 & ~n23081;
  assign n23083 = ~n22823 & ~n23082;
  assign n23084 = ~i_hbusreq3 & ~n23083;
  assign n23085 = ~n23080 & ~n23084;
  assign n23086 = ~controllable_hmaster2 & ~n23085;
  assign n23087 = ~n22808 & ~n23086;
  assign n23088 = ~controllable_hgrant3 & ~n23087;
  assign n23089 = ~n10110 & ~n23088;
  assign n23090 = controllable_nhgrant0 & ~n23089;
  assign n23091 = ~n10240 & ~n23090;
  assign n23092 = ~n3281 & ~n23091;
  assign n23093 = ~n3281 & ~n23092;
  assign n23094 = n3378 & ~n23093;
  assign n23095 = ~n6097 & ~n22769;
  assign n23096 = i_hready & ~n23095;
  assign n23097 = ~n22950 & ~n23096;
  assign n23098 = i_hlock0 & ~n23097;
  assign n23099 = ~n7818 & ~n23098;
  assign n23100 = ~i_hbusreq0 & ~n23099;
  assign n23101 = ~n7813 & ~n23100;
  assign n23102 = ~i_hbusreq4 & ~n23101;
  assign n23103 = ~n7812 & ~n23102;
  assign n23104 = ~controllable_hgrant4 & ~n23103;
  assign n23105 = ~n10112 & ~n23104;
  assign n23106 = ~i_hbusreq2 & ~n23105;
  assign n23107 = ~n7811 & ~n23106;
  assign n23108 = ~controllable_hgrant2 & ~n23107;
  assign n23109 = ~n10111 & ~n23108;
  assign n23110 = controllable_hmaster1 & ~n23109;
  assign n23111 = controllable_hmaster0 & ~n23109;
  assign n23112 = ~n7800 & ~n23005;
  assign n23113 = i_hlock0 & ~n23112;
  assign n23114 = ~n7885 & ~n23113;
  assign n23115 = ~i_hbusreq0 & ~n23114;
  assign n23116 = ~n7882 & ~n23115;
  assign n23117 = ~i_hbusreq4 & ~n23116;
  assign n23118 = ~n7881 & ~n23117;
  assign n23119 = ~controllable_hgrant4 & ~n23118;
  assign n23120 = ~n4667 & ~n23119;
  assign n23121 = ~i_hbusreq2 & ~n23120;
  assign n23122 = ~n13175 & ~n23121;
  assign n23123 = ~controllable_hgrant2 & ~n23122;
  assign n23124 = ~n10111 & ~n23123;
  assign n23125 = ~controllable_hmaster0 & ~n23124;
  assign n23126 = ~n23111 & ~n23125;
  assign n23127 = ~controllable_hmaster1 & ~n23126;
  assign n23128 = ~n23110 & ~n23127;
  assign n23129 = ~i_hbusreq3 & ~n23128;
  assign n23130 = ~n13167 & ~n23129;
  assign n23131 = controllable_hmaster2 & ~n23130;
  assign n23132 = ~controllable_hmaster0 & ~n13190;
  assign n23133 = ~n7874 & ~n23132;
  assign n23134 = ~controllable_hmaster1 & ~n23133;
  assign n23135 = ~n7867 & ~n23134;
  assign n23136 = i_hbusreq3 & ~n23135;
  assign n23137 = ~n10112 & ~n23119;
  assign n23138 = ~i_hbusreq2 & ~n23137;
  assign n23139 = ~n7880 & ~n23138;
  assign n23140 = ~controllable_hgrant2 & ~n23139;
  assign n23141 = ~n10111 & ~n23140;
  assign n23142 = controllable_hmaster0 & ~n23141;
  assign n23143 = ~n10152 & ~n23140;
  assign n23144 = ~controllable_hmaster0 & ~n23143;
  assign n23145 = ~n23142 & ~n23144;
  assign n23146 = controllable_hmaster1 & ~n23145;
  assign n23147 = ~controllable_ndecide & ~n22824;
  assign n23148 = ~n6260 & ~n23147;
  assign n23149 = i_hready & ~n23148;
  assign n23150 = ~n23041 & ~n23149;
  assign n23151 = i_hlock0 & ~n23150;
  assign n23152 = ~n7910 & ~n23151;
  assign n23153 = ~i_hbusreq0 & ~n23152;
  assign n23154 = ~n7904 & ~n23153;
  assign n23155 = ~i_hbusreq4 & ~n23154;
  assign n23156 = ~n7903 & ~n23155;
  assign n23157 = ~controllable_hgrant4 & n23156;
  assign n23158 = ~n10112 & ~n23157;
  assign n23159 = ~i_hbusreq2 & ~n23158;
  assign n23160 = ~n7902 & ~n23159;
  assign n23161 = ~controllable_hgrant2 & ~n23160;
  assign n23162 = ~n10111 & ~n23161;
  assign n23163 = controllable_hmaster0 & ~n23162;
  assign n23164 = ~n23132 & ~n23163;
  assign n23165 = ~controllable_hmaster1 & ~n23164;
  assign n23166 = ~n23146 & ~n23165;
  assign n23167 = ~i_hbusreq3 & ~n23166;
  assign n23168 = ~n23136 & ~n23167;
  assign n23169 = ~controllable_hmaster2 & ~n23168;
  assign n23170 = ~n23131 & ~n23169;
  assign n23171 = ~controllable_hgrant3 & ~n23170;
  assign n23172 = ~n10110 & ~n23171;
  assign n23173 = controllable_nhgrant0 & ~n23172;
  assign n23174 = ~n10240 & ~n23173;
  assign n23175 = ~n3281 & ~n23174;
  assign n23176 = ~n3281 & ~n23175;
  assign n23177 = ~n3378 & ~n23176;
  assign n23178 = ~n23094 & ~n23177;
  assign n23179 = n3492 & ~n23178;
  assign n23180 = ~n21722 & ~n23179;
  assign n23181 = n3485 & ~n23180;
  assign n23182 = ~n21721 & ~n23181;
  assign n23183 = n3476 & ~n23182;
  assign n23184 = ~n23075 & ~n23183;
  assign n23185 = n3374 & ~n23184;
  assign n23186 = ~n22985 & ~n23185;
  assign n23187 = ~n3655 & ~n23186;
  assign n23188 = ~n22948 & ~n23187;
  assign n23189 = n3652 & ~n23188;
  assign n23190 = controllable_hgrant2 & ~n22726;
  assign n23191 = ~n22632 & ~n23190;
  assign n23192 = controllable_hmaster1 & ~n23191;
  assign n23193 = controllable_hmaster0 & ~n23191;
  assign n23194 = controllable_hmaster0 & ~n23193;
  assign n23195 = ~controllable_hmaster1 & ~n23194;
  assign n23196 = ~n23192 & ~n23195;
  assign n23197 = ~i_hbusreq3 & ~n23196;
  assign n23198 = ~n7966 & ~n23197;
  assign n23199 = controllable_hmaster2 & ~n23198;
  assign n23200 = controllable_hmaster2 & ~n23199;
  assign n23201 = ~controllable_hgrant3 & ~n23200;
  assign n23202 = ~n9708 & ~n23201;
  assign n23203 = controllable_nhgrant0 & ~n23202;
  assign n23204 = ~n9753 & ~n23203;
  assign n23205 = ~n3281 & ~n23204;
  assign n23206 = ~n3281 & ~n23205;
  assign n23207 = ~n3378 & ~n23206;
  assign n23208 = ~n22618 & ~n23207;
  assign n23209 = n3492 & ~n23208;
  assign n23210 = n3492 & ~n23209;
  assign n23211 = n3485 & ~n23210;
  assign n23212 = n3485 & ~n23211;
  assign n23213 = ~n3374 & ~n23212;
  assign n23214 = ~n5303 & ~n10775;
  assign n23215 = ~controllable_hmaster1 & ~n23214;
  assign n23216 = ~n5293 & ~n23215;
  assign n23217 = i_hbusreq3 & ~n23216;
  assign n23218 = ~n10775 & ~n22687;
  assign n23219 = ~controllable_hmaster1 & ~n23218;
  assign n23220 = ~n22673 & ~n23219;
  assign n23221 = ~i_hbusreq3 & ~n23220;
  assign n23222 = ~n23217 & ~n23221;
  assign n23223 = ~controllable_hmaster2 & ~n23222;
  assign n23224 = ~n22668 & ~n23223;
  assign n23225 = ~controllable_hgrant3 & ~n23224;
  assign n23226 = ~n9790 & ~n23225;
  assign n23227 = controllable_nhgrant0 & ~n23226;
  assign n23228 = ~n9861 & ~n23227;
  assign n23229 = ~n3281 & ~n23228;
  assign n23230 = ~n3281 & ~n23229;
  assign n23231 = n3378 & ~n23230;
  assign n23232 = ~n22715 & ~n23190;
  assign n23233 = ~controllable_hmaster0 & ~n23232;
  assign n23234 = ~n23193 & ~n23233;
  assign n23235 = ~controllable_hmaster1 & ~n23234;
  assign n23236 = ~n23192 & ~n23235;
  assign n23237 = ~i_hbusreq3 & ~n23236;
  assign n23238 = ~n13270 & ~n23237;
  assign n23239 = controllable_hmaster2 & ~n23238;
  assign n23240 = ~n6703 & ~n10775;
  assign n23241 = ~controllable_hmaster1 & ~n23240;
  assign n23242 = ~n6701 & ~n23241;
  assign n23243 = i_hbusreq3 & ~n23242;
  assign n23244 = controllable_hmaster0 & ~n22726;
  assign n23245 = controllable_hgrant2 & ~n22631;
  assign n23246 = ~n22727 & ~n23245;
  assign n23247 = ~controllable_hmaster0 & ~n23246;
  assign n23248 = ~n23244 & ~n23247;
  assign n23249 = controllable_hmaster1 & ~n23248;
  assign n23250 = ~n22745 & ~n23190;
  assign n23251 = controllable_hmaster0 & ~n23250;
  assign n23252 = ~n10775 & ~n23251;
  assign n23253 = ~controllable_hmaster1 & ~n23252;
  assign n23254 = ~n23249 & ~n23253;
  assign n23255 = ~i_hbusreq3 & ~n23254;
  assign n23256 = ~n23243 & ~n23255;
  assign n23257 = ~controllable_hmaster2 & ~n23256;
  assign n23258 = ~n23239 & ~n23257;
  assign n23259 = ~controllable_hgrant3 & ~n23258;
  assign n23260 = ~n9790 & ~n23259;
  assign n23261 = controllable_nhgrant0 & ~n23260;
  assign n23262 = ~n9861 & ~n23261;
  assign n23263 = ~n3281 & ~n23262;
  assign n23264 = ~n3281 & ~n23263;
  assign n23265 = ~n3378 & ~n23264;
  assign n23266 = ~n23231 & ~n23265;
  assign n23267 = n3492 & ~n23266;
  assign n23268 = n3492 & ~n23267;
  assign n23269 = n3485 & ~n23268;
  assign n23270 = n3485 & ~n23269;
  assign n23271 = ~n3476 & ~n23270;
  assign n23272 = ~controllable_hmaster0 & ~n13301;
  assign n23273 = ~n7339 & ~n23272;
  assign n23274 = ~controllable_hmaster1 & ~n23273;
  assign n23275 = ~n7330 & ~n23274;
  assign n23276 = i_hbusreq3 & ~n23275;
  assign n23277 = ~n22842 & ~n23272;
  assign n23278 = ~controllable_hmaster1 & ~n23277;
  assign n23279 = ~n22823 & ~n23278;
  assign n23280 = ~i_hbusreq3 & ~n23279;
  assign n23281 = ~n23276 & ~n23280;
  assign n23282 = ~controllable_hmaster2 & ~n23281;
  assign n23283 = ~n22808 & ~n23282;
  assign n23284 = ~controllable_hgrant3 & ~n23283;
  assign n23285 = ~n10110 & ~n23284;
  assign n23286 = controllable_nhgrant0 & ~n23285;
  assign n23287 = ~n10240 & ~n23286;
  assign n23288 = ~n3281 & ~n23287;
  assign n23289 = ~n3281 & ~n23288;
  assign n23290 = n3378 & ~n23289;
  assign n23291 = ~n6007 & ~n22703;
  assign n23292 = i_hlock0 & ~n23291;
  assign n23293 = ~n6021 & ~n23292;
  assign n23294 = ~i_hbusreq0 & ~n23293;
  assign n23295 = ~n6016 & ~n23294;
  assign n23296 = ~i_hbusreq4 & ~n23295;
  assign n23297 = ~n6015 & ~n23296;
  assign n23298 = ~controllable_hgrant4 & ~n23297;
  assign n23299 = ~n4617 & ~n23298;
  assign n23300 = ~i_hbusreq2 & ~n23299;
  assign n23301 = ~n6014 & ~n23300;
  assign n23302 = controllable_hgrant2 & ~n23301;
  assign n23303 = ~n22870 & ~n23302;
  assign n23304 = controllable_hmaster1 & ~n23303;
  assign n23305 = controllable_hmaster0 & ~n23303;
  assign n23306 = ~n22885 & ~n23302;
  assign n23307 = ~controllable_hmaster0 & ~n23306;
  assign n23308 = ~n23305 & ~n23307;
  assign n23309 = ~controllable_hmaster1 & ~n23308;
  assign n23310 = ~n23304 & ~n23309;
  assign n23311 = ~i_hbusreq3 & ~n23310;
  assign n23312 = ~n13328 & ~n23311;
  assign n23313 = controllable_hmaster2 & ~n23312;
  assign n23314 = ~controllable_hmaster0 & ~n13340;
  assign n23315 = ~n8082 & ~n23314;
  assign n23316 = ~controllable_hmaster1 & ~n23315;
  assign n23317 = ~n8080 & ~n23316;
  assign n23318 = i_hbusreq3 & ~n23317;
  assign n23319 = ~n22902 & ~n23302;
  assign n23320 = controllable_hmaster0 & ~n23319;
  assign n23321 = ~n4657 & ~n5038;
  assign n23322 = i_hready & ~n23321;
  assign n23323 = ~n22620 & ~n23322;
  assign n23324 = i_hlock0 & ~n23323;
  assign n23325 = ~n6060 & ~n23324;
  assign n23326 = ~i_hbusreq0 & ~n23325;
  assign n23327 = ~n6053 & ~n23326;
  assign n23328 = ~i_hbusreq4 & ~n23327;
  assign n23329 = ~n6052 & ~n23328;
  assign n23330 = ~controllable_hgrant4 & ~n23329;
  assign n23331 = ~n4617 & ~n23330;
  assign n23332 = ~i_hbusreq2 & ~n23331;
  assign n23333 = ~n6051 & ~n23332;
  assign n23334 = controllable_hgrant2 & ~n23333;
  assign n23335 = ~n22902 & ~n23334;
  assign n23336 = ~controllable_hmaster0 & ~n23335;
  assign n23337 = ~n23320 & ~n23336;
  assign n23338 = controllable_hmaster1 & ~n23337;
  assign n23339 = ~n22922 & ~n23302;
  assign n23340 = controllable_hmaster0 & ~n23339;
  assign n23341 = ~n23314 & ~n23340;
  assign n23342 = ~controllable_hmaster1 & ~n23341;
  assign n23343 = ~n23338 & ~n23342;
  assign n23344 = ~i_hbusreq3 & ~n23343;
  assign n23345 = ~n23318 & ~n23344;
  assign n23346 = ~controllable_hmaster2 & ~n23345;
  assign n23347 = ~n23313 & ~n23346;
  assign n23348 = ~controllable_hgrant3 & ~n23347;
  assign n23349 = ~n10110 & ~n23348;
  assign n23350 = controllable_nhgrant0 & ~n23349;
  assign n23351 = ~n10240 & ~n23350;
  assign n23352 = ~n3281 & ~n23351;
  assign n23353 = ~n3281 & ~n23352;
  assign n23354 = ~n3378 & ~n23353;
  assign n23355 = ~n23290 & ~n23354;
  assign n23356 = n3492 & ~n23355;
  assign n23357 = ~n21722 & ~n23356;
  assign n23358 = n3485 & ~n23357;
  assign n23359 = ~n21721 & ~n23358;
  assign n23360 = n3476 & ~n23359;
  assign n23361 = ~n23271 & ~n23360;
  assign n23362 = n3374 & ~n23361;
  assign n23363 = ~n23213 & ~n23362;
  assign n23364 = n3655 & ~n23363;
  assign n23365 = ~n22962 & ~n23190;
  assign n23366 = controllable_hmaster1 & ~n23365;
  assign n23367 = controllable_hmaster0 & ~n23365;
  assign n23368 = controllable_hmaster0 & ~n23367;
  assign n23369 = ~controllable_hmaster1 & ~n23368;
  assign n23370 = ~n23366 & ~n23369;
  assign n23371 = ~i_hbusreq3 & ~n23370;
  assign n23372 = ~n8125 & ~n23371;
  assign n23373 = controllable_hmaster2 & ~n23372;
  assign n23374 = controllable_hmaster2 & ~n23373;
  assign n23375 = ~controllable_hgrant3 & ~n23374;
  assign n23376 = ~n9708 & ~n23375;
  assign n23377 = controllable_nhgrant0 & ~n23376;
  assign n23378 = ~n9753 & ~n23377;
  assign n23379 = ~n3281 & ~n23378;
  assign n23380 = ~n3281 & ~n23379;
  assign n23381 = ~n3378 & ~n23380;
  assign n23382 = ~n22618 & ~n23381;
  assign n23383 = n3492 & ~n23382;
  assign n23384 = n3492 & ~n23383;
  assign n23385 = n3485 & ~n23384;
  assign n23386 = n3485 & ~n23385;
  assign n23387 = ~n3374 & ~n23386;
  assign n23388 = ~n5303 & ~n11210;
  assign n23389 = ~controllable_hmaster1 & ~n23388;
  assign n23390 = ~n5293 & ~n23389;
  assign n23391 = i_hbusreq3 & ~n23390;
  assign n23392 = ~n11210 & ~n22687;
  assign n23393 = ~controllable_hmaster1 & ~n23392;
  assign n23394 = ~n22673 & ~n23393;
  assign n23395 = ~i_hbusreq3 & ~n23394;
  assign n23396 = ~n23391 & ~n23395;
  assign n23397 = ~controllable_hmaster2 & ~n23396;
  assign n23398 = ~n22668 & ~n23397;
  assign n23399 = ~controllable_hgrant3 & ~n23398;
  assign n23400 = ~n9790 & ~n23399;
  assign n23401 = controllable_nhgrant0 & ~n23400;
  assign n23402 = ~n9861 & ~n23401;
  assign n23403 = ~n3281 & ~n23402;
  assign n23404 = ~n3281 & ~n23403;
  assign n23405 = n3378 & ~n23404;
  assign n23406 = ~n23017 & ~n23190;
  assign n23407 = ~controllable_hmaster0 & ~n23406;
  assign n23408 = ~n23367 & ~n23407;
  assign n23409 = ~controllable_hmaster1 & ~n23408;
  assign n23410 = ~n23366 & ~n23409;
  assign n23411 = ~i_hbusreq3 & ~n23410;
  assign n23412 = ~n13401 & ~n23411;
  assign n23413 = controllable_hmaster2 & ~n23412;
  assign n23414 = ~n6933 & ~n11210;
  assign n23415 = ~controllable_hmaster1 & ~n23414;
  assign n23416 = ~n6931 & ~n23415;
  assign n23417 = i_hbusreq3 & ~n23416;
  assign n23418 = ~n23033 & ~n23190;
  assign n23419 = controllable_hmaster0 & ~n23418;
  assign n23420 = ~n23033 & ~n23245;
  assign n23421 = ~controllable_hmaster0 & ~n23420;
  assign n23422 = ~n23419 & ~n23421;
  assign n23423 = controllable_hmaster1 & ~n23422;
  assign n23424 = ~n23053 & ~n23190;
  assign n23425 = controllable_hmaster0 & ~n23424;
  assign n23426 = ~n11210 & ~n23425;
  assign n23427 = ~controllable_hmaster1 & ~n23426;
  assign n23428 = ~n23423 & ~n23427;
  assign n23429 = ~i_hbusreq3 & ~n23428;
  assign n23430 = ~n23417 & ~n23429;
  assign n23431 = ~controllable_hmaster2 & ~n23430;
  assign n23432 = ~n23413 & ~n23431;
  assign n23433 = ~controllable_hgrant3 & ~n23432;
  assign n23434 = ~n9790 & ~n23433;
  assign n23435 = controllable_nhgrant0 & ~n23434;
  assign n23436 = ~n9861 & ~n23435;
  assign n23437 = ~n3281 & ~n23436;
  assign n23438 = ~n3281 & ~n23437;
  assign n23439 = ~n3378 & ~n23438;
  assign n23440 = ~n23405 & ~n23439;
  assign n23441 = n3492 & ~n23440;
  assign n23442 = n3492 & ~n23441;
  assign n23443 = n3485 & ~n23442;
  assign n23444 = n3485 & ~n23443;
  assign n23445 = ~n3476 & ~n23444;
  assign n23446 = ~controllable_hmaster0 & ~n13432;
  assign n23447 = ~n7339 & ~n23446;
  assign n23448 = ~controllable_hmaster1 & ~n23447;
  assign n23449 = ~n7330 & ~n23448;
  assign n23450 = i_hbusreq3 & ~n23449;
  assign n23451 = ~n22842 & ~n23446;
  assign n23452 = ~controllable_hmaster1 & ~n23451;
  assign n23453 = ~n22823 & ~n23452;
  assign n23454 = ~i_hbusreq3 & ~n23453;
  assign n23455 = ~n23450 & ~n23454;
  assign n23456 = ~controllable_hmaster2 & ~n23455;
  assign n23457 = ~n22808 & ~n23456;
  assign n23458 = ~controllable_hgrant3 & ~n23457;
  assign n23459 = ~n10110 & ~n23458;
  assign n23460 = controllable_nhgrant0 & ~n23459;
  assign n23461 = ~n10240 & ~n23460;
  assign n23462 = ~n3281 & ~n23461;
  assign n23463 = ~n3281 & ~n23462;
  assign n23464 = n3378 & ~n23463;
  assign n23465 = ~n23108 & ~n23302;
  assign n23466 = controllable_hmaster1 & ~n23465;
  assign n23467 = controllable_hmaster0 & ~n23465;
  assign n23468 = ~n23123 & ~n23302;
  assign n23469 = ~controllable_hmaster0 & ~n23468;
  assign n23470 = ~n23467 & ~n23469;
  assign n23471 = ~controllable_hmaster1 & ~n23470;
  assign n23472 = ~n23466 & ~n23471;
  assign n23473 = ~i_hbusreq3 & ~n23472;
  assign n23474 = ~n13459 & ~n23473;
  assign n23475 = controllable_hmaster2 & ~n23474;
  assign n23476 = ~controllable_hmaster0 & ~n13471;
  assign n23477 = ~n8237 & ~n23476;
  assign n23478 = ~controllable_hmaster1 & ~n23477;
  assign n23479 = ~n8235 & ~n23478;
  assign n23480 = i_hbusreq3 & ~n23479;
  assign n23481 = ~n23140 & ~n23302;
  assign n23482 = controllable_hmaster0 & ~n23481;
  assign n23483 = ~n23140 & ~n23334;
  assign n23484 = ~controllable_hmaster0 & ~n23483;
  assign n23485 = ~n23482 & ~n23484;
  assign n23486 = controllable_hmaster1 & ~n23485;
  assign n23487 = ~n23161 & ~n23302;
  assign n23488 = controllable_hmaster0 & ~n23487;
  assign n23489 = ~n23476 & ~n23488;
  assign n23490 = ~controllable_hmaster1 & ~n23489;
  assign n23491 = ~n23486 & ~n23490;
  assign n23492 = ~i_hbusreq3 & ~n23491;
  assign n23493 = ~n23480 & ~n23492;
  assign n23494 = ~controllable_hmaster2 & ~n23493;
  assign n23495 = ~n23475 & ~n23494;
  assign n23496 = ~controllable_hgrant3 & ~n23495;
  assign n23497 = ~n10110 & ~n23496;
  assign n23498 = controllable_nhgrant0 & ~n23497;
  assign n23499 = ~n10240 & ~n23498;
  assign n23500 = ~n3281 & ~n23499;
  assign n23501 = ~n3281 & ~n23500;
  assign n23502 = ~n3378 & ~n23501;
  assign n23503 = ~n23464 & ~n23502;
  assign n23504 = n3492 & ~n23503;
  assign n23505 = ~n21722 & ~n23504;
  assign n23506 = n3485 & ~n23505;
  assign n23507 = ~n21721 & ~n23506;
  assign n23508 = n3476 & ~n23507;
  assign n23509 = ~n23445 & ~n23508;
  assign n23510 = n3374 & ~n23509;
  assign n23511 = ~n23387 & ~n23510;
  assign n23512 = ~n3655 & ~n23511;
  assign n23513 = ~n23364 & ~n23512;
  assign n23514 = ~n3652 & ~n23513;
  assign n23515 = ~n23189 & ~n23514;
  assign n23516 = n3368 & ~n23515;
  assign n23517 = ~n22604 & ~n23516;
  assign n23518 = n3362 & ~n23517;
  assign n23519 = n3492 & ~n21862;
  assign n23520 = ~n3631 & ~n23519;
  assign n23521 = n3485 & ~n23520;
  assign n23522 = ~n3630 & ~n23521;
  assign n23523 = ~n3476 & ~n23522;
  assign n23524 = ~n8309 & ~n23519;
  assign n23525 = n3485 & ~n23524;
  assign n23526 = ~n8639 & ~n23525;
  assign n23527 = n3476 & ~n23526;
  assign n23528 = ~n23523 & ~n23527;
  assign n23529 = ~n3374 & ~n23528;
  assign n23530 = n3492 & ~n21948;
  assign n23531 = ~n3631 & ~n23530;
  assign n23532 = n3485 & ~n23531;
  assign n23533 = ~n3630 & ~n23532;
  assign n23534 = ~n3476 & ~n23533;
  assign n23535 = n3492 & ~n22082;
  assign n23536 = ~n8309 & ~n23535;
  assign n23537 = n3485 & ~n23536;
  assign n23538 = ~n8639 & ~n23537;
  assign n23539 = n3476 & ~n23538;
  assign n23540 = ~n23534 & ~n23539;
  assign n23541 = n3374 & ~n23540;
  assign n23542 = ~n23529 & ~n23541;
  assign n23543 = n3655 & ~n23542;
  assign n23544 = n3492 & ~n22106;
  assign n23545 = ~n3631 & ~n23544;
  assign n23546 = n3485 & ~n23545;
  assign n23547 = ~n3630 & ~n23546;
  assign n23548 = ~n3476 & ~n23547;
  assign n23549 = n3492 & ~n8308;
  assign n23550 = ~n8367 & ~n23549;
  assign n23551 = ~n3485 & ~n23550;
  assign n23552 = ~n8309 & ~n23544;
  assign n23553 = n3485 & ~n23552;
  assign n23554 = ~n23551 & ~n23553;
  assign n23555 = n3476 & ~n23554;
  assign n23556 = ~n23548 & ~n23555;
  assign n23557 = ~n3374 & ~n23556;
  assign n23558 = n3492 & ~n22160;
  assign n23559 = ~n3631 & ~n23558;
  assign n23560 = n3485 & ~n23559;
  assign n23561 = ~n3630 & ~n23560;
  assign n23562 = ~n3476 & ~n23561;
  assign n23563 = n3492 & ~n22278;
  assign n23564 = ~n8309 & ~n23563;
  assign n23565 = n3485 & ~n23564;
  assign n23566 = ~n23551 & ~n23565;
  assign n23567 = n3476 & ~n23566;
  assign n23568 = ~n23562 & ~n23567;
  assign n23569 = n3374 & ~n23568;
  assign n23570 = ~n23557 & ~n23569;
  assign n23571 = ~n3655 & ~n23570;
  assign n23572 = ~n23543 & ~n23571;
  assign n23573 = n3652 & ~n23572;
  assign n23574 = n3492 & ~n22304;
  assign n23575 = ~n3631 & ~n23574;
  assign n23576 = n3485 & ~n23575;
  assign n23577 = ~n3630 & ~n23576;
  assign n23578 = ~n3476 & ~n23577;
  assign n23579 = ~n8434 & ~n23549;
  assign n23580 = ~n3485 & ~n23579;
  assign n23581 = ~n8309 & ~n23574;
  assign n23582 = n3485 & ~n23581;
  assign n23583 = ~n23580 & ~n23582;
  assign n23584 = n3476 & ~n23583;
  assign n23585 = ~n23578 & ~n23584;
  assign n23586 = ~n3374 & ~n23585;
  assign n23587 = n3492 & ~n22358;
  assign n23588 = ~n3631 & ~n23587;
  assign n23589 = n3485 & ~n23588;
  assign n23590 = ~n3630 & ~n23589;
  assign n23591 = ~n3476 & ~n23590;
  assign n23592 = n3492 & ~n22447;
  assign n23593 = ~n8309 & ~n23592;
  assign n23594 = n3485 & ~n23593;
  assign n23595 = ~n23580 & ~n23594;
  assign n23596 = n3476 & ~n23595;
  assign n23597 = ~n23591 & ~n23596;
  assign n23598 = n3374 & ~n23597;
  assign n23599 = ~n23586 & ~n23598;
  assign n23600 = n3655 & ~n23599;
  assign n23601 = n3492 & ~n22471;
  assign n23602 = ~n3631 & ~n23601;
  assign n23603 = n3485 & ~n23602;
  assign n23604 = ~n3630 & ~n23603;
  assign n23605 = ~n3476 & ~n23604;
  assign n23606 = ~n8491 & ~n23549;
  assign n23607 = ~n3485 & ~n23606;
  assign n23608 = ~n8309 & ~n23601;
  assign n23609 = n3485 & ~n23608;
  assign n23610 = ~n23607 & ~n23609;
  assign n23611 = n3476 & ~n23610;
  assign n23612 = ~n23605 & ~n23611;
  assign n23613 = ~n3374 & ~n23612;
  assign n23614 = n3492 & ~n22525;
  assign n23615 = ~n3631 & ~n23614;
  assign n23616 = n3485 & ~n23615;
  assign n23617 = ~n3630 & ~n23616;
  assign n23618 = ~n3476 & ~n23617;
  assign n23619 = n3492 & ~n22589;
  assign n23620 = ~n8309 & ~n23619;
  assign n23621 = n3485 & ~n23620;
  assign n23622 = ~n23607 & ~n23621;
  assign n23623 = n3476 & ~n23622;
  assign n23624 = ~n23618 & ~n23623;
  assign n23625 = n3374 & ~n23624;
  assign n23626 = ~n23613 & ~n23625;
  assign n23627 = ~n3655 & ~n23626;
  assign n23628 = ~n23600 & ~n23627;
  assign n23629 = ~n3652 & ~n23628;
  assign n23630 = ~n23573 & ~n23629;
  assign n23631 = ~n3368 & ~n23630;
  assign n23632 = n3492 & ~n22648;
  assign n23633 = n3492 & ~n23632;
  assign n23634 = n3485 & ~n23633;
  assign n23635 = n3485 & ~n23634;
  assign n23636 = ~n3476 & ~n23635;
  assign n23637 = ~n8525 & ~n23634;
  assign n23638 = n3476 & ~n23637;
  assign n23639 = ~n23636 & ~n23638;
  assign n23640 = ~n3374 & ~n23639;
  assign n23641 = n3492 & ~n22760;
  assign n23642 = n3492 & ~n23641;
  assign n23643 = n3485 & ~n23642;
  assign n23644 = n3485 & ~n23643;
  assign n23645 = ~n3476 & ~n23644;
  assign n23646 = n3492 & ~n21260;
  assign n23647 = ~n8536 & ~n23646;
  assign n23648 = ~n3485 & ~n23647;
  assign n23649 = n3492 & ~n22937;
  assign n23650 = ~n21722 & ~n23649;
  assign n23651 = n3485 & ~n23650;
  assign n23652 = ~n23648 & ~n23651;
  assign n23653 = n3476 & ~n23652;
  assign n23654 = ~n23645 & ~n23653;
  assign n23655 = n3374 & ~n23654;
  assign n23656 = ~n23640 & ~n23655;
  assign n23657 = n3655 & ~n23656;
  assign n23658 = n3492 & ~n22978;
  assign n23659 = n3492 & ~n23658;
  assign n23660 = n3485 & ~n23659;
  assign n23661 = n3485 & ~n23660;
  assign n23662 = ~n3476 & ~n23661;
  assign n23663 = ~n8525 & ~n23660;
  assign n23664 = n3476 & ~n23663;
  assign n23665 = ~n23662 & ~n23664;
  assign n23666 = ~n3374 & ~n23665;
  assign n23667 = n3492 & ~n23068;
  assign n23668 = n3492 & ~n23667;
  assign n23669 = n3485 & ~n23668;
  assign n23670 = n3485 & ~n23669;
  assign n23671 = ~n3476 & ~n23670;
  assign n23672 = ~n8563 & ~n23646;
  assign n23673 = ~n3485 & ~n23672;
  assign n23674 = n3492 & ~n23176;
  assign n23675 = ~n21722 & ~n23674;
  assign n23676 = n3485 & ~n23675;
  assign n23677 = ~n23673 & ~n23676;
  assign n23678 = n3476 & ~n23677;
  assign n23679 = ~n23671 & ~n23678;
  assign n23680 = n3374 & ~n23679;
  assign n23681 = ~n23666 & ~n23680;
  assign n23682 = ~n3655 & ~n23681;
  assign n23683 = ~n23657 & ~n23682;
  assign n23684 = n3652 & ~n23683;
  assign n23685 = n3492 & ~n23206;
  assign n23686 = n3492 & ~n23685;
  assign n23687 = n3485 & ~n23686;
  assign n23688 = n3485 & ~n23687;
  assign n23689 = ~n3476 & ~n23688;
  assign n23690 = ~n8525 & ~n23687;
  assign n23691 = n3476 & ~n23690;
  assign n23692 = ~n23689 & ~n23691;
  assign n23693 = ~n3374 & ~n23692;
  assign n23694 = n3492 & ~n23264;
  assign n23695 = n3492 & ~n23694;
  assign n23696 = n3485 & ~n23695;
  assign n23697 = n3485 & ~n23696;
  assign n23698 = ~n3476 & ~n23697;
  assign n23699 = ~n8592 & ~n23646;
  assign n23700 = ~n3485 & ~n23699;
  assign n23701 = n3492 & ~n23353;
  assign n23702 = ~n21722 & ~n23701;
  assign n23703 = n3485 & ~n23702;
  assign n23704 = ~n23700 & ~n23703;
  assign n23705 = n3476 & ~n23704;
  assign n23706 = ~n23698 & ~n23705;
  assign n23707 = n3374 & ~n23706;
  assign n23708 = ~n23693 & ~n23707;
  assign n23709 = n3655 & ~n23708;
  assign n23710 = n3492 & ~n23380;
  assign n23711 = n3492 & ~n23710;
  assign n23712 = n3485 & ~n23711;
  assign n23713 = n3485 & ~n23712;
  assign n23714 = ~n3476 & ~n23713;
  assign n23715 = ~n8525 & ~n23712;
  assign n23716 = n3476 & ~n23715;
  assign n23717 = ~n23714 & ~n23716;
  assign n23718 = ~n3374 & ~n23717;
  assign n23719 = n3492 & ~n23438;
  assign n23720 = n3492 & ~n23719;
  assign n23721 = n3485 & ~n23720;
  assign n23722 = n3485 & ~n23721;
  assign n23723 = ~n3476 & ~n23722;
  assign n23724 = ~n8619 & ~n23646;
  assign n23725 = ~n3485 & ~n23724;
  assign n23726 = n3492 & ~n23501;
  assign n23727 = ~n21722 & ~n23726;
  assign n23728 = n3485 & ~n23727;
  assign n23729 = ~n23725 & ~n23728;
  assign n23730 = n3476 & ~n23729;
  assign n23731 = ~n23723 & ~n23730;
  assign n23732 = n3374 & ~n23731;
  assign n23733 = ~n23718 & ~n23732;
  assign n23734 = ~n3655 & ~n23733;
  assign n23735 = ~n23709 & ~n23734;
  assign n23736 = ~n3652 & ~n23735;
  assign n23737 = ~n23684 & ~n23736;
  assign n23738 = n3368 & ~n23737;
  assign n23739 = ~n23631 & ~n23738;
  assign n23740 = ~n3362 & ~n23739;
  assign n23741 = ~n23518 & ~n23740;
  assign n23742 = n3359 & ~n23741;
  assign n23743 = ~n8650 & ~n23553;
  assign n23744 = n3476 & ~n23743;
  assign n23745 = ~n23548 & ~n23744;
  assign n23746 = ~n3374 & ~n23745;
  assign n23747 = ~n8650 & ~n23565;
  assign n23748 = n3476 & ~n23747;
  assign n23749 = ~n23562 & ~n23748;
  assign n23750 = n3374 & ~n23749;
  assign n23751 = ~n23746 & ~n23750;
  assign n23752 = ~n3655 & ~n23751;
  assign n23753 = ~n23543 & ~n23752;
  assign n23754 = n3652 & ~n23753;
  assign n23755 = ~n8663 & ~n23582;
  assign n23756 = n3476 & ~n23755;
  assign n23757 = ~n23578 & ~n23756;
  assign n23758 = ~n3374 & ~n23757;
  assign n23759 = ~n8663 & ~n23594;
  assign n23760 = n3476 & ~n23759;
  assign n23761 = ~n23591 & ~n23760;
  assign n23762 = n3374 & ~n23761;
  assign n23763 = ~n23758 & ~n23762;
  assign n23764 = n3655 & ~n23763;
  assign n23765 = ~n8674 & ~n23609;
  assign n23766 = n3476 & ~n23765;
  assign n23767 = ~n23605 & ~n23766;
  assign n23768 = ~n3374 & ~n23767;
  assign n23769 = ~n8674 & ~n23621;
  assign n23770 = n3476 & ~n23769;
  assign n23771 = ~n23618 & ~n23770;
  assign n23772 = n3374 & ~n23771;
  assign n23773 = ~n23768 & ~n23772;
  assign n23774 = ~n3655 & ~n23773;
  assign n23775 = ~n23764 & ~n23774;
  assign n23776 = ~n3652 & ~n23775;
  assign n23777 = ~n23754 & ~n23776;
  assign n23778 = ~n3368 & ~n23777;
  assign n23779 = ~n8689 & ~n23634;
  assign n23780 = n3476 & ~n23779;
  assign n23781 = ~n23636 & ~n23780;
  assign n23782 = ~n3374 & ~n23781;
  assign n23783 = ~n8694 & ~n23651;
  assign n23784 = n3476 & ~n23783;
  assign n23785 = ~n23645 & ~n23784;
  assign n23786 = n3374 & ~n23785;
  assign n23787 = ~n23782 & ~n23786;
  assign n23788 = n3655 & ~n23787;
  assign n23789 = ~n8689 & ~n23660;
  assign n23790 = n3476 & ~n23789;
  assign n23791 = ~n23662 & ~n23790;
  assign n23792 = ~n3374 & ~n23791;
  assign n23793 = ~n8705 & ~n23676;
  assign n23794 = n3476 & ~n23793;
  assign n23795 = ~n23671 & ~n23794;
  assign n23796 = n3374 & ~n23795;
  assign n23797 = ~n23792 & ~n23796;
  assign n23798 = ~n3655 & ~n23797;
  assign n23799 = ~n23788 & ~n23798;
  assign n23800 = n3652 & ~n23799;
  assign n23801 = ~n8689 & ~n23687;
  assign n23802 = n3476 & ~n23801;
  assign n23803 = ~n23689 & ~n23802;
  assign n23804 = ~n3374 & ~n23803;
  assign n23805 = ~n8718 & ~n23703;
  assign n23806 = n3476 & ~n23805;
  assign n23807 = ~n23698 & ~n23806;
  assign n23808 = n3374 & ~n23807;
  assign n23809 = ~n23804 & ~n23808;
  assign n23810 = n3655 & ~n23809;
  assign n23811 = ~n8689 & ~n23712;
  assign n23812 = n3476 & ~n23811;
  assign n23813 = ~n23714 & ~n23812;
  assign n23814 = ~n3374 & ~n23813;
  assign n23815 = ~n8729 & ~n23728;
  assign n23816 = n3476 & ~n23815;
  assign n23817 = ~n23723 & ~n23816;
  assign n23818 = n3374 & ~n23817;
  assign n23819 = ~n23814 & ~n23818;
  assign n23820 = ~n3655 & ~n23819;
  assign n23821 = ~n23810 & ~n23820;
  assign n23822 = ~n3652 & ~n23821;
  assign n23823 = ~n23800 & ~n23822;
  assign n23824 = n3368 & ~n23823;
  assign n23825 = ~n23778 & ~n23824;
  assign n23826 = n3362 & ~n23825;
  assign n23827 = n3378 & ~n21862;
  assign n23828 = ~n8789 & ~n23827;
  assign n23829 = n3492 & ~n23828;
  assign n23830 = ~n3631 & ~n23829;
  assign n23831 = n3485 & ~n23830;
  assign n23832 = ~n3630 & ~n23831;
  assign n23833 = ~n3476 & ~n23832;
  assign n23834 = ~n8309 & ~n23829;
  assign n23835 = n3485 & ~n23834;
  assign n23836 = ~n8639 & ~n23835;
  assign n23837 = n3476 & ~n23836;
  assign n23838 = ~n23833 & ~n23837;
  assign n23839 = ~n3374 & ~n23838;
  assign n23840 = n3378 & ~n21948;
  assign n23841 = ~n8906 & ~n23840;
  assign n23842 = n3492 & ~n23841;
  assign n23843 = ~n3631 & ~n23842;
  assign n23844 = n3485 & ~n23843;
  assign n23845 = ~n3630 & ~n23844;
  assign n23846 = ~n3476 & ~n23845;
  assign n23847 = n3378 & ~n22082;
  assign n23848 = ~n9100 & ~n23847;
  assign n23849 = n3492 & ~n23848;
  assign n23850 = ~n8309 & ~n23849;
  assign n23851 = n3485 & ~n23850;
  assign n23852 = ~n8639 & ~n23851;
  assign n23853 = n3476 & ~n23852;
  assign n23854 = ~n23846 & ~n23853;
  assign n23855 = n3374 & ~n23854;
  assign n23856 = ~n23839 & ~n23855;
  assign n23857 = n3655 & ~n23856;
  assign n23858 = n3378 & ~n22106;
  assign n23859 = ~n9135 & ~n23858;
  assign n23860 = n3492 & ~n23859;
  assign n23861 = ~n3631 & ~n23860;
  assign n23862 = n3485 & ~n23861;
  assign n23863 = ~n3630 & ~n23862;
  assign n23864 = ~n3476 & ~n23863;
  assign n23865 = ~n8367 & ~n23860;
  assign n23866 = n3485 & ~n23865;
  assign n23867 = ~n8650 & ~n23866;
  assign n23868 = n3476 & ~n23867;
  assign n23869 = ~n23864 & ~n23868;
  assign n23870 = ~n3374 & ~n23869;
  assign n23871 = n3378 & ~n22160;
  assign n23872 = ~n9240 & ~n23871;
  assign n23873 = n3492 & ~n23872;
  assign n23874 = ~n3631 & ~n23873;
  assign n23875 = n3485 & ~n23874;
  assign n23876 = ~n3630 & ~n23875;
  assign n23877 = ~n3476 & ~n23876;
  assign n23878 = n3378 & ~n22278;
  assign n23879 = ~n9374 & ~n23878;
  assign n23880 = n3492 & ~n23879;
  assign n23881 = ~n8367 & ~n23880;
  assign n23882 = n3485 & ~n23881;
  assign n23883 = ~n8650 & ~n23882;
  assign n23884 = n3476 & ~n23883;
  assign n23885 = ~n23877 & ~n23884;
  assign n23886 = n3374 & ~n23885;
  assign n23887 = ~n23870 & ~n23886;
  assign n23888 = ~n3655 & ~n23887;
  assign n23889 = ~n23857 & ~n23888;
  assign n23890 = n3652 & ~n23889;
  assign n23891 = n3378 & ~n22304;
  assign n23892 = ~n9409 & ~n23891;
  assign n23893 = n3492 & ~n23892;
  assign n23894 = ~n3631 & ~n23893;
  assign n23895 = n3485 & ~n23894;
  assign n23896 = ~n3630 & ~n23895;
  assign n23897 = ~n3476 & ~n23896;
  assign n23898 = ~n8434 & ~n23893;
  assign n23899 = n3485 & ~n23898;
  assign n23900 = ~n8663 & ~n23899;
  assign n23901 = n3476 & ~n23900;
  assign n23902 = ~n23897 & ~n23901;
  assign n23903 = ~n3374 & ~n23902;
  assign n23904 = n3378 & ~n22358;
  assign n23905 = ~n9469 & ~n23904;
  assign n23906 = n3492 & ~n23905;
  assign n23907 = ~n3631 & ~n23906;
  assign n23908 = n3485 & ~n23907;
  assign n23909 = ~n3630 & ~n23908;
  assign n23910 = ~n3476 & ~n23909;
  assign n23911 = n3378 & ~n22447;
  assign n23912 = ~n9531 & ~n23911;
  assign n23913 = n3492 & ~n23912;
  assign n23914 = ~n8434 & ~n23913;
  assign n23915 = n3485 & ~n23914;
  assign n23916 = ~n8663 & ~n23915;
  assign n23917 = n3476 & ~n23916;
  assign n23918 = ~n23910 & ~n23917;
  assign n23919 = n3374 & ~n23918;
  assign n23920 = ~n23903 & ~n23919;
  assign n23921 = n3655 & ~n23920;
  assign n23922 = n3378 & ~n22471;
  assign n23923 = ~n9563 & ~n23922;
  assign n23924 = n3492 & ~n23923;
  assign n23925 = ~n3631 & ~n23924;
  assign n23926 = n3485 & ~n23925;
  assign n23927 = ~n3630 & ~n23926;
  assign n23928 = ~n3476 & ~n23927;
  assign n23929 = ~n8491 & ~n23924;
  assign n23930 = n3485 & ~n23929;
  assign n23931 = ~n8674 & ~n23930;
  assign n23932 = n3476 & ~n23931;
  assign n23933 = ~n23928 & ~n23932;
  assign n23934 = ~n3374 & ~n23933;
  assign n23935 = n3378 & ~n22525;
  assign n23936 = ~n9623 & ~n23935;
  assign n23937 = n3492 & ~n23936;
  assign n23938 = ~n3631 & ~n23937;
  assign n23939 = n3485 & ~n23938;
  assign n23940 = ~n3630 & ~n23939;
  assign n23941 = ~n3476 & ~n23940;
  assign n23942 = n3378 & ~n22589;
  assign n23943 = ~n9683 & ~n23942;
  assign n23944 = n3492 & ~n23943;
  assign n23945 = ~n8491 & ~n23944;
  assign n23946 = n3485 & ~n23945;
  assign n23947 = ~n8674 & ~n23946;
  assign n23948 = n3476 & ~n23947;
  assign n23949 = ~n23941 & ~n23948;
  assign n23950 = n3374 & ~n23949;
  assign n23951 = ~n23934 & ~n23950;
  assign n23952 = ~n3655 & ~n23951;
  assign n23953 = ~n23921 & ~n23952;
  assign n23954 = ~n3652 & ~n23953;
  assign n23955 = ~n23890 & ~n23954;
  assign n23956 = ~n3368 & ~n23955;
  assign n23957 = n3378 & ~n22648;
  assign n23958 = ~n9757 & ~n23957;
  assign n23959 = n3492 & ~n23958;
  assign n23960 = n3492 & ~n23959;
  assign n23961 = n3485 & ~n23960;
  assign n23962 = n3485 & ~n23961;
  assign n23963 = ~n3476 & ~n23962;
  assign n23964 = ~n8523 & ~n23959;
  assign n23965 = n3485 & ~n23964;
  assign n23966 = ~n8689 & ~n23965;
  assign n23967 = n3476 & ~n23966;
  assign n23968 = ~n23963 & ~n23967;
  assign n23969 = ~n3374 & ~n23968;
  assign n23970 = n3378 & ~n22760;
  assign n23971 = ~n9865 & ~n23970;
  assign n23972 = n3492 & ~n23971;
  assign n23973 = n3492 & ~n23972;
  assign n23974 = n3485 & ~n23973;
  assign n23975 = n3485 & ~n23974;
  assign n23976 = ~n3476 & ~n23975;
  assign n23977 = ~n5889 & ~n22620;
  assign n23978 = i_hlock0 & ~n23977;
  assign n23979 = ~n9889 & ~n23978;
  assign n23980 = ~i_hbusreq0 & ~n23979;
  assign n23981 = ~n9885 & ~n23980;
  assign n23982 = ~i_hbusreq4 & ~n23981;
  assign n23983 = ~n9884 & ~n23982;
  assign n23984 = ~controllable_hgrant4 & ~n23983;
  assign n23985 = ~n10112 & ~n23984;
  assign n23986 = ~i_hbusreq2 & ~n23985;
  assign n23987 = ~n9883 & ~n23986;
  assign n23988 = ~controllable_hgrant2 & ~n23987;
  assign n23989 = ~n10111 & ~n23988;
  assign n23990 = controllable_hmaster1 & ~n23989;
  assign n23991 = controllable_hmaster0 & ~n23989;
  assign n23992 = ~n5889 & ~n22703;
  assign n23993 = i_hlock0 & ~n23992;
  assign n23994 = ~n5937 & ~n23993;
  assign n23995 = ~i_hbusreq0 & ~n23994;
  assign n23996 = ~n5933 & ~n23995;
  assign n23997 = ~i_hbusreq4 & ~n23996;
  assign n23998 = ~n5932 & ~n23997;
  assign n23999 = ~controllable_hgrant4 & ~n23998;
  assign n24000 = ~n4667 & ~n23999;
  assign n24001 = ~i_hbusreq2 & ~n24000;
  assign n24002 = ~n12262 & ~n24001;
  assign n24003 = ~controllable_hgrant2 & ~n24002;
  assign n24004 = ~n10111 & ~n24003;
  assign n24005 = ~controllable_hmaster0 & ~n24004;
  assign n24006 = ~n23991 & ~n24005;
  assign n24007 = ~controllable_hmaster1 & ~n24006;
  assign n24008 = ~n23990 & ~n24007;
  assign n24009 = ~i_hbusreq3 & ~n24008;
  assign n24010 = ~n13795 & ~n24009;
  assign n24011 = controllable_hmaster2 & ~n24010;
  assign n24012 = ~n10112 & ~n23999;
  assign n24013 = ~i_hbusreq2 & ~n24012;
  assign n24014 = ~n5931 & ~n24013;
  assign n24015 = ~controllable_hgrant2 & ~n24014;
  assign n24016 = ~n10111 & ~n24015;
  assign n24017 = controllable_hmaster0 & ~n24016;
  assign n24018 = ~n10152 & ~n24015;
  assign n24019 = ~controllable_hmaster0 & ~n24018;
  assign n24020 = ~n24017 & ~n24019;
  assign n24021 = controllable_hmaster1 & ~n24020;
  assign n24022 = ~n10161 & ~n22703;
  assign n24023 = i_hlock0 & ~n24022;
  assign n24024 = ~n5968 & ~n24023;
  assign n24025 = ~i_hbusreq0 & ~n24024;
  assign n24026 = ~n5957 & ~n24025;
  assign n24027 = ~i_hbusreq4 & ~n24026;
  assign n24028 = ~n5956 & ~n24027;
  assign n24029 = ~controllable_hgrant4 & ~n24028;
  assign n24030 = ~n10112 & ~n24029;
  assign n24031 = ~i_hbusreq2 & ~n24030;
  assign n24032 = ~n5955 & ~n24031;
  assign n24033 = ~controllable_hgrant2 & ~n24032;
  assign n24034 = ~n10111 & ~n24033;
  assign n24035 = controllable_hmaster0 & ~n24034;
  assign n24036 = ~n10186 & ~n24035;
  assign n24037 = ~controllable_hmaster1 & ~n24036;
  assign n24038 = ~n24021 & ~n24037;
  assign n24039 = ~i_hbusreq3 & ~n24038;
  assign n24040 = ~n22045 & ~n24039;
  assign n24041 = ~controllable_hmaster2 & ~n24040;
  assign n24042 = ~n24011 & ~n24041;
  assign n24043 = ~controllable_hgrant3 & ~n24042;
  assign n24044 = ~n10110 & ~n24043;
  assign n24045 = controllable_nhgrant0 & ~n24044;
  assign n24046 = ~n10240 & ~n24045;
  assign n24047 = ~n3281 & ~n24046;
  assign n24048 = ~n3281 & ~n24047;
  assign n24049 = n3378 & ~n24048;
  assign n24050 = ~n10244 & ~n24049;
  assign n24051 = n3492 & ~n24050;
  assign n24052 = ~n8536 & ~n24051;
  assign n24053 = n3485 & ~n24052;
  assign n24054 = ~n8694 & ~n24053;
  assign n24055 = n3476 & ~n24054;
  assign n24056 = ~n23976 & ~n24055;
  assign n24057 = n3374 & ~n24056;
  assign n24058 = ~n23969 & ~n24057;
  assign n24059 = n3655 & ~n24058;
  assign n24060 = n3378 & ~n22978;
  assign n24061 = ~n10299 & ~n24060;
  assign n24062 = n3492 & ~n24061;
  assign n24063 = n3492 & ~n24062;
  assign n24064 = n3485 & ~n24063;
  assign n24065 = n3485 & ~n24064;
  assign n24066 = ~n3476 & ~n24065;
  assign n24067 = ~n8523 & ~n24062;
  assign n24068 = n3485 & ~n24067;
  assign n24069 = ~n8689 & ~n24068;
  assign n24070 = n3476 & ~n24069;
  assign n24071 = ~n24066 & ~n24070;
  assign n24072 = ~n3374 & ~n24071;
  assign n24073 = n3378 & ~n23068;
  assign n24074 = ~n10390 & ~n24073;
  assign n24075 = n3492 & ~n24074;
  assign n24076 = n3492 & ~n24075;
  assign n24077 = n3485 & ~n24076;
  assign n24078 = n3485 & ~n24077;
  assign n24079 = ~n3476 & ~n24078;
  assign n24080 = ~i_hready & n22949;
  assign n24081 = ~n10460 & ~n24080;
  assign n24082 = i_hlock0 & ~n24081;
  assign n24083 = ~n10437 & ~n24082;
  assign n24084 = ~i_hbusreq0 & ~n24083;
  assign n24085 = ~n10423 & ~n24084;
  assign n24086 = ~i_hbusreq4 & ~n24085;
  assign n24087 = ~n10422 & ~n24086;
  assign n24088 = ~controllable_hgrant4 & n24087;
  assign n24089 = ~n10112 & ~n24088;
  assign n24090 = ~i_hbusreq2 & ~n24089;
  assign n24091 = ~n10421 & ~n24090;
  assign n24092 = ~controllable_hgrant2 & ~n24091;
  assign n24093 = ~n10111 & ~n24092;
  assign n24094 = controllable_hmaster1 & ~n24093;
  assign n24095 = controllable_hmaster0 & ~n24093;
  assign n24096 = ~i_hready & n23004;
  assign n24097 = ~n10460 & ~n24096;
  assign n24098 = i_hlock0 & ~n24097;
  assign n24099 = ~n10515 & ~n24098;
  assign n24100 = ~i_hbusreq0 & ~n24099;
  assign n24101 = ~n10510 & ~n24100;
  assign n24102 = ~i_hbusreq4 & ~n24101;
  assign n24103 = ~n10509 & ~n24102;
  assign n24104 = ~controllable_hgrant4 & n24103;
  assign n24105 = ~n4667 & ~n24104;
  assign n24106 = ~i_hbusreq2 & ~n24105;
  assign n24107 = ~n13882 & ~n24106;
  assign n24108 = ~controllable_hgrant2 & ~n24107;
  assign n24109 = ~n10111 & ~n24108;
  assign n24110 = ~controllable_hmaster0 & ~n24109;
  assign n24111 = ~n24095 & ~n24110;
  assign n24112 = ~controllable_hmaster1 & ~n24111;
  assign n24113 = ~n24094 & ~n24112;
  assign n24114 = ~i_hbusreq3 & ~n24113;
  assign n24115 = ~n13874 & ~n24114;
  assign n24116 = controllable_hmaster2 & ~n24115;
  assign n24117 = ~n10502 & ~n10643;
  assign n24118 = ~controllable_hmaster1 & ~n24117;
  assign n24119 = ~n10491 & ~n24118;
  assign n24120 = i_hbusreq3 & ~n24119;
  assign n24121 = ~n10112 & ~n24104;
  assign n24122 = ~i_hbusreq2 & ~n24121;
  assign n24123 = ~n10508 & ~n24122;
  assign n24124 = ~controllable_hgrant2 & ~n24123;
  assign n24125 = ~n10111 & ~n24124;
  assign n24126 = controllable_hmaster0 & ~n24125;
  assign n24127 = ~n10152 & ~n24124;
  assign n24128 = ~controllable_hmaster0 & ~n24127;
  assign n24129 = ~n24126 & ~n24128;
  assign n24130 = controllable_hmaster1 & ~n24129;
  assign n24131 = ~n10664 & ~n23041;
  assign n24132 = i_hlock0 & ~n24131;
  assign n24133 = ~n10546 & ~n24132;
  assign n24134 = ~i_hbusreq0 & ~n24133;
  assign n24135 = ~n10534 & ~n24134;
  assign n24136 = ~i_hbusreq4 & ~n24135;
  assign n24137 = ~n10533 & ~n24136;
  assign n24138 = ~controllable_hgrant4 & n24137;
  assign n24139 = ~n10112 & ~n24138;
  assign n24140 = ~i_hbusreq2 & ~n24139;
  assign n24141 = ~n10532 & ~n24140;
  assign n24142 = ~controllable_hgrant2 & ~n24141;
  assign n24143 = ~n10111 & ~n24142;
  assign n24144 = controllable_hmaster0 & ~n24143;
  assign n24145 = ~n10691 & ~n24144;
  assign n24146 = ~controllable_hmaster1 & ~n24145;
  assign n24147 = ~n24130 & ~n24146;
  assign n24148 = ~i_hbusreq3 & ~n24147;
  assign n24149 = ~n24120 & ~n24148;
  assign n24150 = ~controllable_hmaster2 & ~n24149;
  assign n24151 = ~n24116 & ~n24150;
  assign n24152 = ~controllable_hgrant3 & ~n24151;
  assign n24153 = ~n10110 & ~n24152;
  assign n24154 = controllable_nhgrant0 & ~n24153;
  assign n24155 = ~n10240 & ~n24154;
  assign n24156 = ~n3281 & ~n24155;
  assign n24157 = ~n3281 & ~n24156;
  assign n24158 = n3378 & ~n24157;
  assign n24159 = ~n10705 & ~n24158;
  assign n24160 = n3492 & ~n24159;
  assign n24161 = ~n8563 & ~n24160;
  assign n24162 = n3485 & ~n24161;
  assign n24163 = ~n8705 & ~n24162;
  assign n24164 = n3476 & ~n24163;
  assign n24165 = ~n24079 & ~n24164;
  assign n24166 = n3374 & ~n24165;
  assign n24167 = ~n24072 & ~n24166;
  assign n24168 = ~n3655 & ~n24167;
  assign n24169 = ~n24059 & ~n24168;
  assign n24170 = n3652 & ~n24169;
  assign n24171 = n3378 & ~n23206;
  assign n24172 = ~n10742 & ~n24171;
  assign n24173 = n3492 & ~n24172;
  assign n24174 = n3492 & ~n24173;
  assign n24175 = n3485 & ~n24174;
  assign n24176 = n3485 & ~n24175;
  assign n24177 = ~n3476 & ~n24176;
  assign n24178 = ~n8523 & ~n24173;
  assign n24179 = n3485 & ~n24178;
  assign n24180 = ~n8689 & ~n24179;
  assign n24181 = n3476 & ~n24180;
  assign n24182 = ~n24177 & ~n24181;
  assign n24183 = ~n3374 & ~n24182;
  assign n24184 = n3378 & ~n23264;
  assign n24185 = ~n10802 & ~n24184;
  assign n24186 = n3492 & ~n24185;
  assign n24187 = n3492 & ~n24186;
  assign n24188 = n3485 & ~n24187;
  assign n24189 = n3485 & ~n24188;
  assign n24190 = ~n3476 & ~n24189;
  assign n24191 = ~n10842 & ~n22703;
  assign n24192 = i_hlock0 & ~n24191;
  assign n24193 = ~n10844 & ~n24192;
  assign n24194 = ~i_hbusreq0 & ~n24193;
  assign n24195 = ~n10836 & ~n24194;
  assign n24196 = ~i_hbusreq4 & ~n24195;
  assign n24197 = ~n10835 & ~n24196;
  assign n24198 = ~controllable_hgrant4 & ~n24197;
  assign n24199 = ~n4617 & ~n24198;
  assign n24200 = i_hlock2 & ~n24199;
  assign n24201 = ~n9958 & ~n22703;
  assign n24202 = i_hlock0 & ~n24201;
  assign n24203 = ~n9960 & ~n24202;
  assign n24204 = ~i_hbusreq0 & ~n24203;
  assign n24205 = ~n10854 & ~n24204;
  assign n24206 = ~i_hbusreq4 & ~n24205;
  assign n24207 = ~n10853 & ~n24206;
  assign n24208 = ~controllable_hgrant4 & ~n24207;
  assign n24209 = ~n4617 & ~n24208;
  assign n24210 = ~i_hlock2 & ~n24209;
  assign n24211 = ~n24200 & ~n24210;
  assign n24212 = ~i_hbusreq2 & ~n24211;
  assign n24213 = ~n10834 & ~n24212;
  assign n24214 = controllable_hgrant2 & ~n24213;
  assign n24215 = ~n23988 & ~n24214;
  assign n24216 = controllable_hmaster1 & ~n24215;
  assign n24217 = controllable_hmaster0 & ~n24215;
  assign n24218 = ~n24003 & ~n24214;
  assign n24219 = ~controllable_hmaster0 & ~n24218;
  assign n24220 = ~n24217 & ~n24219;
  assign n24221 = ~controllable_hmaster1 & ~n24220;
  assign n24222 = ~n24216 & ~n24221;
  assign n24223 = ~i_hbusreq3 & ~n24222;
  assign n24224 = ~n13963 & ~n24223;
  assign n24225 = controllable_hmaster2 & ~n24224;
  assign n24226 = ~n10928 & ~n11073;
  assign n24227 = ~controllable_hmaster1 & ~n24226;
  assign n24228 = ~n10926 & ~n24227;
  assign n24229 = i_hbusreq3 & ~n24228;
  assign n24230 = ~n24015 & ~n24214;
  assign n24231 = controllable_hmaster0 & ~n24230;
  assign n24232 = ~n10842 & ~n22620;
  assign n24233 = i_hlock0 & ~n24232;
  assign n24234 = ~n10946 & ~n24233;
  assign n24235 = ~i_hbusreq0 & ~n24234;
  assign n24236 = ~n10938 & ~n24235;
  assign n24237 = ~i_hbusreq4 & ~n24236;
  assign n24238 = ~n10937 & ~n24237;
  assign n24239 = ~controllable_hgrant4 & ~n24238;
  assign n24240 = ~n4617 & ~n24239;
  assign n24241 = i_hlock2 & ~n24240;
  assign n24242 = ~n11096 & ~n22620;
  assign n24243 = i_hlock0 & ~n24242;
  assign n24244 = ~n10034 & ~n24243;
  assign n24245 = ~i_hbusreq0 & ~n24244;
  assign n24246 = ~n10956 & ~n24245;
  assign n24247 = ~i_hbusreq4 & ~n24246;
  assign n24248 = ~n10955 & ~n24247;
  assign n24249 = ~controllable_hgrant4 & ~n24248;
  assign n24250 = ~n4617 & ~n24249;
  assign n24251 = ~i_hlock2 & ~n24250;
  assign n24252 = ~n24241 & ~n24251;
  assign n24253 = ~i_hbusreq2 & ~n24252;
  assign n24254 = ~n10936 & ~n24253;
  assign n24255 = controllable_hgrant2 & ~n24254;
  assign n24256 = ~n24015 & ~n24255;
  assign n24257 = ~controllable_hmaster0 & ~n24256;
  assign n24258 = ~n24231 & ~n24257;
  assign n24259 = controllable_hmaster1 & ~n24258;
  assign n24260 = ~n24033 & ~n24214;
  assign n24261 = controllable_hmaster0 & ~n24260;
  assign n24262 = ~n11129 & ~n24261;
  assign n24263 = ~controllable_hmaster1 & ~n24262;
  assign n24264 = ~n24259 & ~n24263;
  assign n24265 = ~i_hbusreq3 & ~n24264;
  assign n24266 = ~n24229 & ~n24265;
  assign n24267 = ~controllable_hmaster2 & ~n24266;
  assign n24268 = ~n24225 & ~n24267;
  assign n24269 = ~controllable_hgrant3 & ~n24268;
  assign n24270 = ~n10110 & ~n24269;
  assign n24271 = controllable_nhgrant0 & ~n24270;
  assign n24272 = ~n10240 & ~n24271;
  assign n24273 = ~n3281 & ~n24272;
  assign n24274 = ~n3281 & ~n24273;
  assign n24275 = n3378 & ~n24274;
  assign n24276 = ~n11143 & ~n24275;
  assign n24277 = n3492 & ~n24276;
  assign n24278 = ~n8592 & ~n24277;
  assign n24279 = n3485 & ~n24278;
  assign n24280 = ~n8718 & ~n24279;
  assign n24281 = n3476 & ~n24280;
  assign n24282 = ~n24190 & ~n24281;
  assign n24283 = n3374 & ~n24282;
  assign n24284 = ~n24183 & ~n24283;
  assign n24285 = n3655 & ~n24284;
  assign n24286 = n3378 & ~n23380;
  assign n24287 = ~n11178 & ~n24286;
  assign n24288 = n3492 & ~n24287;
  assign n24289 = n3492 & ~n24288;
  assign n24290 = n3485 & ~n24289;
  assign n24291 = n3485 & ~n24290;
  assign n24292 = ~n3476 & ~n24291;
  assign n24293 = ~n8523 & ~n24288;
  assign n24294 = n3485 & ~n24293;
  assign n24295 = ~n8689 & ~n24294;
  assign n24296 = n3476 & ~n24295;
  assign n24297 = ~n24292 & ~n24296;
  assign n24298 = ~n3374 & ~n24297;
  assign n24299 = n3378 & ~n23438;
  assign n24300 = ~n11236 & ~n24299;
  assign n24301 = n3492 & ~n24300;
  assign n24302 = n3492 & ~n24301;
  assign n24303 = n3485 & ~n24302;
  assign n24304 = n3485 & ~n24303;
  assign n24305 = ~n3476 & ~n24304;
  assign n24306 = ~n24092 & ~n24214;
  assign n24307 = controllable_hmaster1 & ~n24306;
  assign n24308 = controllable_hmaster0 & ~n24306;
  assign n24309 = ~n24108 & ~n24214;
  assign n24310 = ~controllable_hmaster0 & ~n24309;
  assign n24311 = ~n24308 & ~n24310;
  assign n24312 = ~controllable_hmaster1 & ~n24311;
  assign n24313 = ~n24307 & ~n24312;
  assign n24314 = ~i_hbusreq3 & ~n24313;
  assign n24315 = ~n14025 & ~n24314;
  assign n24316 = controllable_hmaster2 & ~n24315;
  assign n24317 = ~n11270 & ~n11324;
  assign n24318 = ~controllable_hmaster1 & ~n24317;
  assign n24319 = ~n11268 & ~n24318;
  assign n24320 = i_hbusreq3 & ~n24319;
  assign n24321 = ~n24124 & ~n24214;
  assign n24322 = controllable_hmaster0 & ~n24321;
  assign n24323 = ~n24124 & ~n24255;
  assign n24324 = ~controllable_hmaster0 & ~n24323;
  assign n24325 = ~n24322 & ~n24324;
  assign n24326 = controllable_hmaster1 & ~n24325;
  assign n24327 = ~n24142 & ~n24214;
  assign n24328 = controllable_hmaster0 & ~n24327;
  assign n24329 = ~n11338 & ~n24328;
  assign n24330 = ~controllable_hmaster1 & ~n24329;
  assign n24331 = ~n24326 & ~n24330;
  assign n24332 = ~i_hbusreq3 & ~n24331;
  assign n24333 = ~n24320 & ~n24332;
  assign n24334 = ~controllable_hmaster2 & ~n24333;
  assign n24335 = ~n24316 & ~n24334;
  assign n24336 = ~controllable_hgrant3 & ~n24335;
  assign n24337 = ~n10110 & ~n24336;
  assign n24338 = controllable_nhgrant0 & ~n24337;
  assign n24339 = ~n10240 & ~n24338;
  assign n24340 = ~n3281 & ~n24339;
  assign n24341 = ~n3281 & ~n24340;
  assign n24342 = n3378 & ~n24341;
  assign n24343 = ~n11352 & ~n24342;
  assign n24344 = n3492 & ~n24343;
  assign n24345 = ~n8619 & ~n24344;
  assign n24346 = n3485 & ~n24345;
  assign n24347 = ~n8729 & ~n24346;
  assign n24348 = n3476 & ~n24347;
  assign n24349 = ~n24305 & ~n24348;
  assign n24350 = n3374 & ~n24349;
  assign n24351 = ~n24298 & ~n24350;
  assign n24352 = ~n3655 & ~n24351;
  assign n24353 = ~n24285 & ~n24352;
  assign n24354 = ~n3652 & ~n24353;
  assign n24355 = ~n24170 & ~n24354;
  assign n24356 = n3368 & ~n24355;
  assign n24357 = ~n23956 & ~n24356;
  assign n24358 = ~n3362 & ~n24357;
  assign n24359 = ~n23826 & ~n24358;
  assign n24360 = ~n3359 & ~n24359;
  assign n24361 = ~n23742 & ~n24360;
  assign n24362 = ~n3356 & ~n24361;
  assign n24363 = ~n21848 & ~n24362;
  assign n24364 = n3345 & ~n24363;
  assign n24365 = ~n21250 & ~n24364;
  assign n24366 = ~n3341 & ~n24365;
  assign n24367 = controllable_hmaster2 & ~n21262;
  assign n24368 = controllable_hgrant3 & ~n24367;
  assign n24369 = controllable_hmaster2 & ~n21339;
  assign n24370 = ~controllable_hgrant3 & ~n24369;
  assign n24371 = ~n24368 & ~n24370;
  assign n24372 = controllable_nhgrant0 & ~n24371;
  assign n24373 = controllable_hmaster2 & ~n21272;
  assign n24374 = ~controllable_hgrant3 & ~n24373;
  assign n24375 = ~n24368 & ~n24374;
  assign n24376 = ~controllable_nhgrant0 & ~n24375;
  assign n24377 = ~n24372 & ~n24376;
  assign n24378 = ~n3281 & ~n24377;
  assign n24379 = ~n3783 & ~n24378;
  assign n24380 = ~n3378 & ~n24379;
  assign n24381 = ~n3378 & ~n24380;
  assign n24382 = n3492 & ~n24381;
  assign n24383 = ~n3493 & ~n24382;
  assign n24384 = n3485 & ~n24383;
  assign n24385 = ~n3486 & ~n24384;
  assign n24386 = ~n3476 & ~n24385;
  assign n24387 = ~n3281 & ~n8787;
  assign n24388 = n3378 & ~n24387;
  assign n24389 = ~n8789 & ~n24388;
  assign n24390 = n3492 & ~n24389;
  assign n24391 = ~n3493 & ~n24390;
  assign n24392 = n3485 & ~n24391;
  assign n24393 = ~n3486 & ~n24392;
  assign n24394 = n3476 & ~n24393;
  assign n24395 = ~n24386 & ~n24394;
  assign n24396 = ~n3374 & ~n24395;
  assign n24397 = ~n3950 & ~n24378;
  assign n24398 = ~n3378 & ~n24397;
  assign n24399 = ~n3378 & ~n24398;
  assign n24400 = n3492 & ~n24399;
  assign n24401 = ~n3493 & ~n24400;
  assign n24402 = n3485 & ~n24401;
  assign n24403 = ~n3486 & ~n24402;
  assign n24404 = ~n3476 & ~n24403;
  assign n24405 = ~n3281 & ~n9098;
  assign n24406 = n3378 & ~n24405;
  assign n24407 = ~n9100 & ~n24406;
  assign n24408 = n3492 & ~n24407;
  assign n24409 = ~n3493 & ~n24408;
  assign n24410 = n3485 & ~n24409;
  assign n24411 = ~n3486 & ~n24410;
  assign n24412 = n3476 & ~n24411;
  assign n24413 = ~n24404 & ~n24412;
  assign n24414 = n3374 & ~n24413;
  assign n24415 = ~n24396 & ~n24414;
  assign n24416 = n3655 & ~n24415;
  assign n24417 = controllable_hmaster2 & ~n17639;
  assign n24418 = controllable_hmaster2 & ~n24417;
  assign n24419 = ~controllable_hgrant3 & ~n24418;
  assign n24420 = ~n24368 & ~n24419;
  assign n24421 = controllable_nhgrant0 & ~n24420;
  assign n24422 = ~n24376 & ~n24421;
  assign n24423 = ~n3281 & ~n24422;
  assign n24424 = ~n3783 & ~n24423;
  assign n24425 = ~n3378 & ~n24424;
  assign n24426 = ~n3378 & ~n24425;
  assign n24427 = n3492 & ~n24426;
  assign n24428 = ~n3493 & ~n24427;
  assign n24429 = n3485 & ~n24428;
  assign n24430 = ~n3486 & ~n24429;
  assign n24431 = ~n3476 & ~n24430;
  assign n24432 = ~n3281 & ~n9133;
  assign n24433 = n3378 & ~n24432;
  assign n24434 = ~n9135 & ~n24433;
  assign n24435 = n3492 & ~n24434;
  assign n24436 = ~n3493 & ~n24435;
  assign n24437 = n3485 & ~n24436;
  assign n24438 = ~n3486 & ~n24437;
  assign n24439 = n3476 & ~n24438;
  assign n24440 = ~n24431 & ~n24439;
  assign n24441 = ~n3374 & ~n24440;
  assign n24442 = ~n3950 & ~n24423;
  assign n24443 = ~n3378 & ~n24442;
  assign n24444 = ~n3378 & ~n24443;
  assign n24445 = n3492 & ~n24444;
  assign n24446 = ~n3493 & ~n24445;
  assign n24447 = n3485 & ~n24446;
  assign n24448 = ~n3486 & ~n24447;
  assign n24449 = ~n3476 & ~n24448;
  assign n24450 = ~n3281 & ~n9372;
  assign n24451 = n3378 & ~n24450;
  assign n24452 = ~n9374 & ~n24451;
  assign n24453 = n3492 & ~n24452;
  assign n24454 = ~n3493 & ~n24453;
  assign n24455 = n3485 & ~n24454;
  assign n24456 = ~n3486 & ~n24455;
  assign n24457 = n3476 & ~n24456;
  assign n24458 = ~n24449 & ~n24457;
  assign n24459 = n3374 & ~n24458;
  assign n24460 = ~n24441 & ~n24459;
  assign n24461 = ~n3655 & ~n24460;
  assign n24462 = ~n24416 & ~n24461;
  assign n24463 = n3652 & ~n24462;
  assign n24464 = controllable_hmaster2 & ~n14460;
  assign n24465 = controllable_hmaster2 & ~n24464;
  assign n24466 = ~controllable_hgrant3 & ~n24465;
  assign n24467 = ~n24368 & ~n24466;
  assign n24468 = controllable_nhgrant0 & ~n24467;
  assign n24469 = ~n24376 & ~n24468;
  assign n24470 = ~n3281 & ~n24469;
  assign n24471 = ~n3783 & ~n24470;
  assign n24472 = ~n3378 & ~n24471;
  assign n24473 = ~n3378 & ~n24472;
  assign n24474 = n3492 & ~n24473;
  assign n24475 = ~n3493 & ~n24474;
  assign n24476 = n3485 & ~n24475;
  assign n24477 = ~n3486 & ~n24476;
  assign n24478 = ~n3476 & ~n24477;
  assign n24479 = ~n3281 & ~n9407;
  assign n24480 = n3378 & ~n24479;
  assign n24481 = ~n9409 & ~n24480;
  assign n24482 = n3492 & ~n24481;
  assign n24483 = ~n3493 & ~n24482;
  assign n24484 = n3485 & ~n24483;
  assign n24485 = ~n3486 & ~n24484;
  assign n24486 = n3476 & ~n24485;
  assign n24487 = ~n24478 & ~n24486;
  assign n24488 = ~n3374 & ~n24487;
  assign n24489 = ~n3950 & ~n24470;
  assign n24490 = ~n3378 & ~n24489;
  assign n24491 = ~n3378 & ~n24490;
  assign n24492 = n3492 & ~n24491;
  assign n24493 = ~n3493 & ~n24492;
  assign n24494 = n3485 & ~n24493;
  assign n24495 = ~n3486 & ~n24494;
  assign n24496 = ~n3476 & ~n24495;
  assign n24497 = ~n3281 & ~n9529;
  assign n24498 = n3378 & ~n24497;
  assign n24499 = ~n9531 & ~n24498;
  assign n24500 = n3492 & ~n24499;
  assign n24501 = ~n3493 & ~n24500;
  assign n24502 = n3485 & ~n24501;
  assign n24503 = ~n3486 & ~n24502;
  assign n24504 = n3476 & ~n24503;
  assign n24505 = ~n24496 & ~n24504;
  assign n24506 = n3374 & ~n24505;
  assign n24507 = ~n24488 & ~n24506;
  assign n24508 = n3655 & ~n24507;
  assign n24509 = controllable_hmaster0 & ~n9545;
  assign n24510 = ~controllable_hmaster1 & ~n24509;
  assign n24511 = ~n9544 & ~n24510;
  assign n24512 = controllable_hmaster2 & ~n24511;
  assign n24513 = controllable_hmaster2 & ~n24512;
  assign n24514 = ~controllable_hgrant3 & ~n24513;
  assign n24515 = ~n24368 & ~n24514;
  assign n24516 = controllable_nhgrant0 & ~n24515;
  assign n24517 = ~n24376 & ~n24516;
  assign n24518 = ~n3281 & ~n24517;
  assign n24519 = ~n3783 & ~n24518;
  assign n24520 = ~n3378 & ~n24519;
  assign n24521 = ~n3378 & ~n24520;
  assign n24522 = n3492 & ~n24521;
  assign n24523 = ~n3493 & ~n24522;
  assign n24524 = n3485 & ~n24523;
  assign n24525 = ~n3486 & ~n24524;
  assign n24526 = ~n3476 & ~n24525;
  assign n24527 = ~n3281 & ~n9561;
  assign n24528 = n3378 & ~n24527;
  assign n24529 = ~n9563 & ~n24528;
  assign n24530 = n3492 & ~n24529;
  assign n24531 = ~n3493 & ~n24530;
  assign n24532 = n3485 & ~n24531;
  assign n24533 = ~n3486 & ~n24532;
  assign n24534 = n3476 & ~n24533;
  assign n24535 = ~n24526 & ~n24534;
  assign n24536 = ~n3374 & ~n24535;
  assign n24537 = ~n3950 & ~n24518;
  assign n24538 = ~n3378 & ~n24537;
  assign n24539 = ~n3378 & ~n24538;
  assign n24540 = n3492 & ~n24539;
  assign n24541 = ~n3493 & ~n24540;
  assign n24542 = n3485 & ~n24541;
  assign n24543 = ~n3486 & ~n24542;
  assign n24544 = ~n3476 & ~n24543;
  assign n24545 = ~n3281 & ~n9681;
  assign n24546 = n3378 & ~n24545;
  assign n24547 = ~n9683 & ~n24546;
  assign n24548 = n3492 & ~n24547;
  assign n24549 = ~n3493 & ~n24548;
  assign n24550 = n3485 & ~n24549;
  assign n24551 = ~n3486 & ~n24550;
  assign n24552 = n3476 & ~n24551;
  assign n24553 = ~n24544 & ~n24552;
  assign n24554 = n3374 & ~n24553;
  assign n24555 = ~n24536 & ~n24554;
  assign n24556 = ~n3655 & ~n24555;
  assign n24557 = ~n24508 & ~n24556;
  assign n24558 = ~n3652 & ~n24557;
  assign n24559 = ~n24463 & ~n24558;
  assign n24560 = ~n3368 & ~n24559;
  assign n24561 = n3492 & ~n9756;
  assign n24562 = n3492 & ~n24561;
  assign n24563 = n3485 & ~n24562;
  assign n24564 = n3485 & ~n24563;
  assign n24565 = n3476 & ~n24564;
  assign n24566 = n3476 & ~n24565;
  assign n24567 = ~n3374 & ~n24566;
  assign n24568 = n3492 & ~n10243;
  assign n24569 = n3492 & ~n24568;
  assign n24570 = n3485 & ~n24569;
  assign n24571 = n3485 & ~n24570;
  assign n24572 = n3476 & ~n24571;
  assign n24573 = n3476 & ~n24572;
  assign n24574 = n3374 & ~n24573;
  assign n24575 = ~n24567 & ~n24574;
  assign n24576 = n3655 & ~n24575;
  assign n24577 = n3492 & ~n10298;
  assign n24578 = n3492 & ~n24577;
  assign n24579 = n3485 & ~n24578;
  assign n24580 = n3485 & ~n24579;
  assign n24581 = n3476 & ~n24580;
  assign n24582 = n3476 & ~n24581;
  assign n24583 = ~n3374 & ~n24582;
  assign n24584 = n3492 & ~n10704;
  assign n24585 = n3492 & ~n24584;
  assign n24586 = n3485 & ~n24585;
  assign n24587 = n3485 & ~n24586;
  assign n24588 = n3476 & ~n24587;
  assign n24589 = n3476 & ~n24588;
  assign n24590 = n3374 & ~n24589;
  assign n24591 = ~n24583 & ~n24590;
  assign n24592 = ~n3655 & ~n24591;
  assign n24593 = ~n24576 & ~n24592;
  assign n24594 = n3652 & ~n24593;
  assign n24595 = n3492 & ~n10741;
  assign n24596 = n3492 & ~n24595;
  assign n24597 = n3485 & ~n24596;
  assign n24598 = n3485 & ~n24597;
  assign n24599 = n3476 & ~n24598;
  assign n24600 = n3476 & ~n24599;
  assign n24601 = ~n3374 & ~n24600;
  assign n24602 = n3492 & ~n11142;
  assign n24603 = n3492 & ~n24602;
  assign n24604 = n3485 & ~n24603;
  assign n24605 = n3485 & ~n24604;
  assign n24606 = n3476 & ~n24605;
  assign n24607 = n3476 & ~n24606;
  assign n24608 = n3374 & ~n24607;
  assign n24609 = ~n24601 & ~n24608;
  assign n24610 = n3655 & ~n24609;
  assign n24611 = n3492 & ~n11177;
  assign n24612 = n3492 & ~n24611;
  assign n24613 = n3485 & ~n24612;
  assign n24614 = n3485 & ~n24613;
  assign n24615 = n3476 & ~n24614;
  assign n24616 = n3476 & ~n24615;
  assign n24617 = ~n3374 & ~n24616;
  assign n24618 = n3492 & ~n11351;
  assign n24619 = n3492 & ~n24618;
  assign n24620 = n3485 & ~n24619;
  assign n24621 = n3485 & ~n24620;
  assign n24622 = n3476 & ~n24621;
  assign n24623 = n3476 & ~n24622;
  assign n24624 = n3374 & ~n24623;
  assign n24625 = ~n24617 & ~n24624;
  assign n24626 = ~n3655 & ~n24625;
  assign n24627 = ~n24610 & ~n24626;
  assign n24628 = ~n3652 & ~n24627;
  assign n24629 = ~n24594 & ~n24628;
  assign n24630 = n3368 & ~n24629;
  assign n24631 = ~n24560 & ~n24630;
  assign n24632 = ~n3362 & ~n24631;
  assign n24633 = ~n3362 & ~n24632;
  assign n24634 = ~n3359 & ~n24633;
  assign n24635 = ~n3359 & ~n24634;
  assign n24636 = n3356 & ~n24635;
  assign n24637 = n3492 & ~n8788;
  assign n24638 = ~n3631 & ~n24637;
  assign n24639 = n3485 & ~n24638;
  assign n24640 = ~n3630 & ~n24639;
  assign n24641 = ~n3374 & ~n24640;
  assign n24642 = n3492 & ~n8905;
  assign n24643 = ~n3631 & ~n24642;
  assign n24644 = n3485 & ~n24643;
  assign n24645 = ~n3630 & ~n24644;
  assign n24646 = ~n3476 & ~n24645;
  assign n24647 = n3492 & ~n9099;
  assign n24648 = ~n3631 & ~n24647;
  assign n24649 = n3485 & ~n24648;
  assign n24650 = ~n3630 & ~n24649;
  assign n24651 = n3476 & ~n24650;
  assign n24652 = ~n24646 & ~n24651;
  assign n24653 = n3374 & ~n24652;
  assign n24654 = ~n24641 & ~n24653;
  assign n24655 = n3655 & ~n24654;
  assign n24656 = n3492 & ~n9134;
  assign n24657 = ~n3631 & ~n24656;
  assign n24658 = n3485 & ~n24657;
  assign n24659 = ~n3630 & ~n24658;
  assign n24660 = ~n3374 & ~n24659;
  assign n24661 = n3492 & ~n9239;
  assign n24662 = ~n3631 & ~n24661;
  assign n24663 = n3485 & ~n24662;
  assign n24664 = ~n3630 & ~n24663;
  assign n24665 = ~n3476 & ~n24664;
  assign n24666 = n3492 & ~n9373;
  assign n24667 = ~n3631 & ~n24666;
  assign n24668 = n3485 & ~n24667;
  assign n24669 = ~n3630 & ~n24668;
  assign n24670 = n3476 & ~n24669;
  assign n24671 = ~n24665 & ~n24670;
  assign n24672 = n3374 & ~n24671;
  assign n24673 = ~n24660 & ~n24672;
  assign n24674 = ~n3655 & ~n24673;
  assign n24675 = ~n24655 & ~n24674;
  assign n24676 = n3652 & ~n24675;
  assign n24677 = n3492 & ~n9408;
  assign n24678 = ~n3631 & ~n24677;
  assign n24679 = n3485 & ~n24678;
  assign n24680 = ~n3630 & ~n24679;
  assign n24681 = ~n3374 & ~n24680;
  assign n24682 = n3492 & ~n9468;
  assign n24683 = ~n3631 & ~n24682;
  assign n24684 = n3485 & ~n24683;
  assign n24685 = ~n3630 & ~n24684;
  assign n24686 = ~n3476 & ~n24685;
  assign n24687 = n3492 & ~n9530;
  assign n24688 = ~n3631 & ~n24687;
  assign n24689 = n3485 & ~n24688;
  assign n24690 = ~n3630 & ~n24689;
  assign n24691 = n3476 & ~n24690;
  assign n24692 = ~n24686 & ~n24691;
  assign n24693 = n3374 & ~n24692;
  assign n24694 = ~n24681 & ~n24693;
  assign n24695 = n3655 & ~n24694;
  assign n24696 = n3492 & ~n9562;
  assign n24697 = ~n3631 & ~n24696;
  assign n24698 = n3485 & ~n24697;
  assign n24699 = ~n3630 & ~n24698;
  assign n24700 = ~n3374 & ~n24699;
  assign n24701 = n3492 & ~n9622;
  assign n24702 = ~n3631 & ~n24701;
  assign n24703 = n3485 & ~n24702;
  assign n24704 = ~n3630 & ~n24703;
  assign n24705 = ~n3476 & ~n24704;
  assign n24706 = n3492 & ~n9682;
  assign n24707 = ~n3631 & ~n24706;
  assign n24708 = n3485 & ~n24707;
  assign n24709 = ~n3630 & ~n24708;
  assign n24710 = n3476 & ~n24709;
  assign n24711 = ~n24705 & ~n24710;
  assign n24712 = n3374 & ~n24711;
  assign n24713 = ~n24700 & ~n24712;
  assign n24714 = ~n3655 & ~n24713;
  assign n24715 = ~n24695 & ~n24714;
  assign n24716 = ~n3652 & ~n24715;
  assign n24717 = ~n24676 & ~n24716;
  assign n24718 = ~n3368 & ~n24717;
  assign n24719 = ~n3374 & ~n24564;
  assign n24720 = n3492 & ~n9864;
  assign n24721 = n3492 & ~n24720;
  assign n24722 = n3485 & ~n24721;
  assign n24723 = n3485 & ~n24722;
  assign n24724 = ~n3476 & ~n24723;
  assign n24725 = ~n24572 & ~n24724;
  assign n24726 = n3374 & ~n24725;
  assign n24727 = ~n24719 & ~n24726;
  assign n24728 = n3655 & ~n24727;
  assign n24729 = ~n3374 & ~n24580;
  assign n24730 = n3492 & ~n10389;
  assign n24731 = n3492 & ~n24730;
  assign n24732 = n3485 & ~n24731;
  assign n24733 = n3485 & ~n24732;
  assign n24734 = ~n3476 & ~n24733;
  assign n24735 = ~n24588 & ~n24734;
  assign n24736 = n3374 & ~n24735;
  assign n24737 = ~n24729 & ~n24736;
  assign n24738 = ~n3655 & ~n24737;
  assign n24739 = ~n24728 & ~n24738;
  assign n24740 = n3652 & ~n24739;
  assign n24741 = ~n3374 & ~n24598;
  assign n24742 = n3492 & ~n10801;
  assign n24743 = n3492 & ~n24742;
  assign n24744 = n3485 & ~n24743;
  assign n24745 = n3485 & ~n24744;
  assign n24746 = ~n3476 & ~n24745;
  assign n24747 = ~n24606 & ~n24746;
  assign n24748 = n3374 & ~n24747;
  assign n24749 = ~n24741 & ~n24748;
  assign n24750 = n3655 & ~n24749;
  assign n24751 = ~n3374 & ~n24614;
  assign n24752 = n3492 & ~n11235;
  assign n24753 = n3492 & ~n24752;
  assign n24754 = n3485 & ~n24753;
  assign n24755 = n3485 & ~n24754;
  assign n24756 = ~n3476 & ~n24755;
  assign n24757 = ~n24622 & ~n24756;
  assign n24758 = n3374 & ~n24757;
  assign n24759 = ~n24751 & ~n24758;
  assign n24760 = ~n3655 & ~n24759;
  assign n24761 = ~n24750 & ~n24760;
  assign n24762 = ~n3652 & ~n24761;
  assign n24763 = ~n24740 & ~n24762;
  assign n24764 = n3368 & ~n24763;
  assign n24765 = ~n24718 & ~n24764;
  assign n24766 = n3362 & ~n24765;
  assign n24767 = ~n3476 & ~n24640;
  assign n24768 = ~n8312 & ~n24639;
  assign n24769 = n3476 & ~n24768;
  assign n24770 = ~n24767 & ~n24769;
  assign n24771 = ~n3374 & ~n24770;
  assign n24772 = ~n8312 & ~n24649;
  assign n24773 = n3476 & ~n24772;
  assign n24774 = ~n24646 & ~n24773;
  assign n24775 = n3374 & ~n24774;
  assign n24776 = ~n24771 & ~n24775;
  assign n24777 = n3655 & ~n24776;
  assign n24778 = ~n3476 & ~n24659;
  assign n24779 = ~n8369 & ~n24658;
  assign n24780 = n3476 & ~n24779;
  assign n24781 = ~n24778 & ~n24780;
  assign n24782 = ~n3374 & ~n24781;
  assign n24783 = ~n8369 & ~n24668;
  assign n24784 = n3476 & ~n24783;
  assign n24785 = ~n24665 & ~n24784;
  assign n24786 = n3374 & ~n24785;
  assign n24787 = ~n24782 & ~n24786;
  assign n24788 = ~n3655 & ~n24787;
  assign n24789 = ~n24777 & ~n24788;
  assign n24790 = n3652 & ~n24789;
  assign n24791 = ~n3476 & ~n24680;
  assign n24792 = ~n8436 & ~n24679;
  assign n24793 = n3476 & ~n24792;
  assign n24794 = ~n24791 & ~n24793;
  assign n24795 = ~n3374 & ~n24794;
  assign n24796 = ~n8436 & ~n24689;
  assign n24797 = n3476 & ~n24796;
  assign n24798 = ~n24686 & ~n24797;
  assign n24799 = n3374 & ~n24798;
  assign n24800 = ~n24795 & ~n24799;
  assign n24801 = n3655 & ~n24800;
  assign n24802 = ~n3476 & ~n24699;
  assign n24803 = ~n8493 & ~n24698;
  assign n24804 = n3476 & ~n24803;
  assign n24805 = ~n24802 & ~n24804;
  assign n24806 = ~n3374 & ~n24805;
  assign n24807 = ~n8493 & ~n24708;
  assign n24808 = n3476 & ~n24807;
  assign n24809 = ~n24705 & ~n24808;
  assign n24810 = n3374 & ~n24809;
  assign n24811 = ~n24806 & ~n24810;
  assign n24812 = ~n3655 & ~n24811;
  assign n24813 = ~n24801 & ~n24812;
  assign n24814 = ~n3652 & ~n24813;
  assign n24815 = ~n24790 & ~n24814;
  assign n24816 = ~n3368 & ~n24815;
  assign n24817 = ~n3476 & ~n24564;
  assign n24818 = ~n8525 & ~n24563;
  assign n24819 = n3476 & ~n24818;
  assign n24820 = ~n24817 & ~n24819;
  assign n24821 = ~n3374 & ~n24820;
  assign n24822 = ~n8538 & ~n24570;
  assign n24823 = n3476 & ~n24822;
  assign n24824 = ~n24724 & ~n24823;
  assign n24825 = n3374 & ~n24824;
  assign n24826 = ~n24821 & ~n24825;
  assign n24827 = n3655 & ~n24826;
  assign n24828 = ~n3476 & ~n24580;
  assign n24829 = ~n8525 & ~n24579;
  assign n24830 = n3476 & ~n24829;
  assign n24831 = ~n24828 & ~n24830;
  assign n24832 = ~n3374 & ~n24831;
  assign n24833 = ~n8565 & ~n24586;
  assign n24834 = n3476 & ~n24833;
  assign n24835 = ~n24734 & ~n24834;
  assign n24836 = n3374 & ~n24835;
  assign n24837 = ~n24832 & ~n24836;
  assign n24838 = ~n3655 & ~n24837;
  assign n24839 = ~n24827 & ~n24838;
  assign n24840 = n3652 & ~n24839;
  assign n24841 = ~n3476 & ~n24598;
  assign n24842 = ~n8525 & ~n24597;
  assign n24843 = n3476 & ~n24842;
  assign n24844 = ~n24841 & ~n24843;
  assign n24845 = ~n3374 & ~n24844;
  assign n24846 = ~n8594 & ~n24604;
  assign n24847 = n3476 & ~n24846;
  assign n24848 = ~n24746 & ~n24847;
  assign n24849 = n3374 & ~n24848;
  assign n24850 = ~n24845 & ~n24849;
  assign n24851 = n3655 & ~n24850;
  assign n24852 = ~n3476 & ~n24614;
  assign n24853 = ~n8525 & ~n24613;
  assign n24854 = n3476 & ~n24853;
  assign n24855 = ~n24852 & ~n24854;
  assign n24856 = ~n3374 & ~n24855;
  assign n24857 = ~n8621 & ~n24620;
  assign n24858 = n3476 & ~n24857;
  assign n24859 = ~n24756 & ~n24858;
  assign n24860 = n3374 & ~n24859;
  assign n24861 = ~n24856 & ~n24860;
  assign n24862 = ~n3655 & ~n24861;
  assign n24863 = ~n24851 & ~n24862;
  assign n24864 = ~n3652 & ~n24863;
  assign n24865 = ~n24840 & ~n24864;
  assign n24866 = n3368 & ~n24865;
  assign n24867 = ~n24816 & ~n24866;
  assign n24868 = ~n3362 & ~n24867;
  assign n24869 = ~n24766 & ~n24868;
  assign n24870 = n3359 & ~n24869;
  assign n24871 = ~n8639 & ~n24639;
  assign n24872 = n3476 & ~n24871;
  assign n24873 = ~n24767 & ~n24872;
  assign n24874 = ~n3374 & ~n24873;
  assign n24875 = ~n8639 & ~n24649;
  assign n24876 = n3476 & ~n24875;
  assign n24877 = ~n24646 & ~n24876;
  assign n24878 = n3374 & ~n24877;
  assign n24879 = ~n24874 & ~n24878;
  assign n24880 = n3655 & ~n24879;
  assign n24881 = ~n8650 & ~n24658;
  assign n24882 = n3476 & ~n24881;
  assign n24883 = ~n24778 & ~n24882;
  assign n24884 = ~n3374 & ~n24883;
  assign n24885 = ~n8650 & ~n24668;
  assign n24886 = n3476 & ~n24885;
  assign n24887 = ~n24665 & ~n24886;
  assign n24888 = n3374 & ~n24887;
  assign n24889 = ~n24884 & ~n24888;
  assign n24890 = ~n3655 & ~n24889;
  assign n24891 = ~n24880 & ~n24890;
  assign n24892 = n3652 & ~n24891;
  assign n24893 = ~n8663 & ~n24679;
  assign n24894 = n3476 & ~n24893;
  assign n24895 = ~n24791 & ~n24894;
  assign n24896 = ~n3374 & ~n24895;
  assign n24897 = ~n8663 & ~n24689;
  assign n24898 = n3476 & ~n24897;
  assign n24899 = ~n24686 & ~n24898;
  assign n24900 = n3374 & ~n24899;
  assign n24901 = ~n24896 & ~n24900;
  assign n24902 = n3655 & ~n24901;
  assign n24903 = ~n8674 & ~n24698;
  assign n24904 = n3476 & ~n24903;
  assign n24905 = ~n24802 & ~n24904;
  assign n24906 = ~n3374 & ~n24905;
  assign n24907 = ~n8674 & ~n24708;
  assign n24908 = n3476 & ~n24907;
  assign n24909 = ~n24705 & ~n24908;
  assign n24910 = n3374 & ~n24909;
  assign n24911 = ~n24906 & ~n24910;
  assign n24912 = ~n3655 & ~n24911;
  assign n24913 = ~n24902 & ~n24912;
  assign n24914 = ~n3652 & ~n24913;
  assign n24915 = ~n24892 & ~n24914;
  assign n24916 = ~n3368 & ~n24915;
  assign n24917 = ~n8689 & ~n24563;
  assign n24918 = n3476 & ~n24917;
  assign n24919 = ~n24817 & ~n24918;
  assign n24920 = ~n3374 & ~n24919;
  assign n24921 = ~n8694 & ~n24570;
  assign n24922 = n3476 & ~n24921;
  assign n24923 = ~n24724 & ~n24922;
  assign n24924 = n3374 & ~n24923;
  assign n24925 = ~n24920 & ~n24924;
  assign n24926 = n3655 & ~n24925;
  assign n24927 = ~n8689 & ~n24579;
  assign n24928 = n3476 & ~n24927;
  assign n24929 = ~n24828 & ~n24928;
  assign n24930 = ~n3374 & ~n24929;
  assign n24931 = ~n8705 & ~n24586;
  assign n24932 = n3476 & ~n24931;
  assign n24933 = ~n24734 & ~n24932;
  assign n24934 = n3374 & ~n24933;
  assign n24935 = ~n24930 & ~n24934;
  assign n24936 = ~n3655 & ~n24935;
  assign n24937 = ~n24926 & ~n24936;
  assign n24938 = n3652 & ~n24937;
  assign n24939 = ~n8689 & ~n24597;
  assign n24940 = n3476 & ~n24939;
  assign n24941 = ~n24841 & ~n24940;
  assign n24942 = ~n3374 & ~n24941;
  assign n24943 = ~n8718 & ~n24604;
  assign n24944 = n3476 & ~n24943;
  assign n24945 = ~n24746 & ~n24944;
  assign n24946 = n3374 & ~n24945;
  assign n24947 = ~n24942 & ~n24946;
  assign n24948 = n3655 & ~n24947;
  assign n24949 = ~n8689 & ~n24613;
  assign n24950 = n3476 & ~n24949;
  assign n24951 = ~n24852 & ~n24950;
  assign n24952 = ~n3374 & ~n24951;
  assign n24953 = ~n8729 & ~n24620;
  assign n24954 = n3476 & ~n24953;
  assign n24955 = ~n24756 & ~n24954;
  assign n24956 = n3374 & ~n24955;
  assign n24957 = ~n24952 & ~n24956;
  assign n24958 = ~n3655 & ~n24957;
  assign n24959 = ~n24948 & ~n24958;
  assign n24960 = ~n3652 & ~n24959;
  assign n24961 = ~n24938 & ~n24960;
  assign n24962 = n3368 & ~n24961;
  assign n24963 = ~n24916 & ~n24962;
  assign n24964 = n3362 & ~n24963;
  assign n24965 = ~n8309 & ~n24637;
  assign n24966 = n3485 & ~n24965;
  assign n24967 = ~n8639 & ~n24966;
  assign n24968 = n3476 & ~n24967;
  assign n24969 = ~n24767 & ~n24968;
  assign n24970 = ~n3374 & ~n24969;
  assign n24971 = ~n8309 & ~n24647;
  assign n24972 = n3485 & ~n24971;
  assign n24973 = ~n8639 & ~n24972;
  assign n24974 = n3476 & ~n24973;
  assign n24975 = ~n24646 & ~n24974;
  assign n24976 = n3374 & ~n24975;
  assign n24977 = ~n24970 & ~n24976;
  assign n24978 = n3655 & ~n24977;
  assign n24979 = ~n8367 & ~n24656;
  assign n24980 = n3485 & ~n24979;
  assign n24981 = ~n8650 & ~n24980;
  assign n24982 = n3476 & ~n24981;
  assign n24983 = ~n24778 & ~n24982;
  assign n24984 = ~n3374 & ~n24983;
  assign n24985 = ~n8367 & ~n24666;
  assign n24986 = n3485 & ~n24985;
  assign n24987 = ~n8650 & ~n24986;
  assign n24988 = n3476 & ~n24987;
  assign n24989 = ~n24665 & ~n24988;
  assign n24990 = n3374 & ~n24989;
  assign n24991 = ~n24984 & ~n24990;
  assign n24992 = ~n3655 & ~n24991;
  assign n24993 = ~n24978 & ~n24992;
  assign n24994 = n3652 & ~n24993;
  assign n24995 = ~n8434 & ~n24677;
  assign n24996 = n3485 & ~n24995;
  assign n24997 = ~n8663 & ~n24996;
  assign n24998 = n3476 & ~n24997;
  assign n24999 = ~n24791 & ~n24998;
  assign n25000 = ~n3374 & ~n24999;
  assign n25001 = ~n8434 & ~n24687;
  assign n25002 = n3485 & ~n25001;
  assign n25003 = ~n8663 & ~n25002;
  assign n25004 = n3476 & ~n25003;
  assign n25005 = ~n24686 & ~n25004;
  assign n25006 = n3374 & ~n25005;
  assign n25007 = ~n25000 & ~n25006;
  assign n25008 = n3655 & ~n25007;
  assign n25009 = ~n8491 & ~n24696;
  assign n25010 = n3485 & ~n25009;
  assign n25011 = ~n8674 & ~n25010;
  assign n25012 = n3476 & ~n25011;
  assign n25013 = ~n24802 & ~n25012;
  assign n25014 = ~n3374 & ~n25013;
  assign n25015 = ~n8491 & ~n24706;
  assign n25016 = n3485 & ~n25015;
  assign n25017 = ~n8674 & ~n25016;
  assign n25018 = n3476 & ~n25017;
  assign n25019 = ~n24705 & ~n25018;
  assign n25020 = n3374 & ~n25019;
  assign n25021 = ~n25014 & ~n25020;
  assign n25022 = ~n3655 & ~n25021;
  assign n25023 = ~n25008 & ~n25022;
  assign n25024 = ~n3652 & ~n25023;
  assign n25025 = ~n24994 & ~n25024;
  assign n25026 = ~n3368 & ~n25025;
  assign n25027 = ~n8523 & ~n24561;
  assign n25028 = n3485 & ~n25027;
  assign n25029 = ~n8689 & ~n25028;
  assign n25030 = n3476 & ~n25029;
  assign n25031 = ~n24817 & ~n25030;
  assign n25032 = ~n3374 & ~n25031;
  assign n25033 = ~n8536 & ~n24568;
  assign n25034 = n3485 & ~n25033;
  assign n25035 = ~n8694 & ~n25034;
  assign n25036 = n3476 & ~n25035;
  assign n25037 = ~n24724 & ~n25036;
  assign n25038 = n3374 & ~n25037;
  assign n25039 = ~n25032 & ~n25038;
  assign n25040 = n3655 & ~n25039;
  assign n25041 = ~n8523 & ~n24577;
  assign n25042 = n3485 & ~n25041;
  assign n25043 = ~n8689 & ~n25042;
  assign n25044 = n3476 & ~n25043;
  assign n25045 = ~n24828 & ~n25044;
  assign n25046 = ~n3374 & ~n25045;
  assign n25047 = ~n8563 & ~n24584;
  assign n25048 = n3485 & ~n25047;
  assign n25049 = ~n8705 & ~n25048;
  assign n25050 = n3476 & ~n25049;
  assign n25051 = ~n24734 & ~n25050;
  assign n25052 = n3374 & ~n25051;
  assign n25053 = ~n25046 & ~n25052;
  assign n25054 = ~n3655 & ~n25053;
  assign n25055 = ~n25040 & ~n25054;
  assign n25056 = n3652 & ~n25055;
  assign n25057 = ~n8523 & ~n24595;
  assign n25058 = n3485 & ~n25057;
  assign n25059 = ~n8689 & ~n25058;
  assign n25060 = n3476 & ~n25059;
  assign n25061 = ~n24841 & ~n25060;
  assign n25062 = ~n3374 & ~n25061;
  assign n25063 = ~n8592 & ~n24602;
  assign n25064 = n3485 & ~n25063;
  assign n25065 = ~n8718 & ~n25064;
  assign n25066 = n3476 & ~n25065;
  assign n25067 = ~n24746 & ~n25066;
  assign n25068 = n3374 & ~n25067;
  assign n25069 = ~n25062 & ~n25068;
  assign n25070 = n3655 & ~n25069;
  assign n25071 = ~n8523 & ~n24611;
  assign n25072 = n3485 & ~n25071;
  assign n25073 = ~n8689 & ~n25072;
  assign n25074 = n3476 & ~n25073;
  assign n25075 = ~n24852 & ~n25074;
  assign n25076 = ~n3374 & ~n25075;
  assign n25077 = ~n8619 & ~n24618;
  assign n25078 = n3485 & ~n25077;
  assign n25079 = ~n8729 & ~n25078;
  assign n25080 = n3476 & ~n25079;
  assign n25081 = ~n24756 & ~n25080;
  assign n25082 = n3374 & ~n25081;
  assign n25083 = ~n25076 & ~n25082;
  assign n25084 = ~n3655 & ~n25083;
  assign n25085 = ~n25070 & ~n25084;
  assign n25086 = ~n3652 & ~n25085;
  assign n25087 = ~n25056 & ~n25086;
  assign n25088 = n3368 & ~n25087;
  assign n25089 = ~n25026 & ~n25088;
  assign n25090 = ~n3362 & ~n25089;
  assign n25091 = ~n24964 & ~n25090;
  assign n25092 = ~n3359 & ~n25091;
  assign n25093 = ~n24870 & ~n25092;
  assign n25094 = ~n3356 & ~n25093;
  assign n25095 = ~n24636 & ~n25094;
  assign n25096 = ~n3345 & ~n25095;
  assign n25097 = ~n3378 & ~n8789;
  assign n25098 = n3492 & ~n25097;
  assign n25099 = ~n3493 & ~n25098;
  assign n25100 = n3485 & ~n25099;
  assign n25101 = ~n3486 & ~n25100;
  assign n25102 = ~n3476 & ~n25101;
  assign n25103 = ~n3378 & ~n21287;
  assign n25104 = ~n3485 & ~n25103;
  assign n25105 = ~n3492 & ~n25103;
  assign n25106 = ~n25098 & ~n25105;
  assign n25107 = n3485 & ~n25106;
  assign n25108 = ~n25104 & ~n25107;
  assign n25109 = n3476 & ~n25108;
  assign n25110 = ~n25102 & ~n25109;
  assign n25111 = ~n3374 & ~n25110;
  assign n25112 = n3378 & ~n8522;
  assign n25113 = ~n3468 & ~n25112;
  assign n25114 = ~n3485 & ~n25113;
  assign n25115 = ~n3492 & ~n25113;
  assign n25116 = ~n3281 & ~n8904;
  assign n25117 = n3378 & ~n25116;
  assign n25118 = ~n8906 & ~n25117;
  assign n25119 = n3492 & ~n25118;
  assign n25120 = ~n25115 & ~n25119;
  assign n25121 = n3485 & ~n25120;
  assign n25122 = ~n25114 & ~n25121;
  assign n25123 = ~n3476 & ~n25122;
  assign n25124 = n3378 & ~n8535;
  assign n25125 = ~n21287 & ~n25124;
  assign n25126 = ~n3485 & ~n25125;
  assign n25127 = ~n3492 & ~n25125;
  assign n25128 = ~n24408 & ~n25127;
  assign n25129 = n3485 & ~n25128;
  assign n25130 = ~n25126 & ~n25129;
  assign n25131 = n3476 & ~n25130;
  assign n25132 = ~n25123 & ~n25131;
  assign n25133 = n3374 & ~n25132;
  assign n25134 = ~n25111 & ~n25133;
  assign n25135 = n3655 & ~n25134;
  assign n25136 = ~n3378 & ~n9135;
  assign n25137 = n3492 & ~n25136;
  assign n25138 = ~n3493 & ~n25137;
  assign n25139 = n3485 & ~n25138;
  assign n25140 = ~n3486 & ~n25139;
  assign n25141 = ~n3476 & ~n25140;
  assign n25142 = ~n3378 & ~n8366;
  assign n25143 = ~n3378 & ~n25142;
  assign n25144 = ~n3485 & ~n25143;
  assign n25145 = ~n3492 & ~n25143;
  assign n25146 = ~n25137 & ~n25145;
  assign n25147 = n3485 & ~n25146;
  assign n25148 = ~n25144 & ~n25147;
  assign n25149 = n3476 & ~n25148;
  assign n25150 = ~n25141 & ~n25149;
  assign n25151 = ~n3374 & ~n25150;
  assign n25152 = ~n3281 & ~n9238;
  assign n25153 = n3378 & ~n25152;
  assign n25154 = ~n9240 & ~n25153;
  assign n25155 = n3492 & ~n25154;
  assign n25156 = ~n25115 & ~n25155;
  assign n25157 = n3485 & ~n25156;
  assign n25158 = ~n25114 & ~n25157;
  assign n25159 = ~n3476 & ~n25158;
  assign n25160 = n3378 & ~n8562;
  assign n25161 = ~n25142 & ~n25160;
  assign n25162 = ~n3485 & ~n25161;
  assign n25163 = ~n3492 & ~n25161;
  assign n25164 = ~n24453 & ~n25163;
  assign n25165 = n3485 & ~n25164;
  assign n25166 = ~n25162 & ~n25165;
  assign n25167 = n3476 & ~n25166;
  assign n25168 = ~n25159 & ~n25167;
  assign n25169 = n3374 & ~n25168;
  assign n25170 = ~n25151 & ~n25169;
  assign n25171 = ~n3655 & ~n25170;
  assign n25172 = ~n25135 & ~n25171;
  assign n25173 = n3652 & ~n25172;
  assign n25174 = ~n3378 & ~n9409;
  assign n25175 = n3492 & ~n25174;
  assign n25176 = ~n3493 & ~n25175;
  assign n25177 = n3485 & ~n25176;
  assign n25178 = ~n3486 & ~n25177;
  assign n25179 = ~n3476 & ~n25178;
  assign n25180 = ~n3378 & ~n8433;
  assign n25181 = ~n3378 & ~n25180;
  assign n25182 = ~n3485 & ~n25181;
  assign n25183 = ~n3492 & ~n25181;
  assign n25184 = ~n25175 & ~n25183;
  assign n25185 = n3485 & ~n25184;
  assign n25186 = ~n25182 & ~n25185;
  assign n25187 = n3476 & ~n25186;
  assign n25188 = ~n25179 & ~n25187;
  assign n25189 = ~n3374 & ~n25188;
  assign n25190 = ~n3281 & ~n9467;
  assign n25191 = n3378 & ~n25190;
  assign n25192 = ~n9469 & ~n25191;
  assign n25193 = n3492 & ~n25192;
  assign n25194 = ~n25115 & ~n25193;
  assign n25195 = n3485 & ~n25194;
  assign n25196 = ~n25114 & ~n25195;
  assign n25197 = ~n3476 & ~n25196;
  assign n25198 = n3378 & ~n8591;
  assign n25199 = ~n25180 & ~n25198;
  assign n25200 = ~n3485 & ~n25199;
  assign n25201 = ~n3492 & ~n25199;
  assign n25202 = ~n24500 & ~n25201;
  assign n25203 = n3485 & ~n25202;
  assign n25204 = ~n25200 & ~n25203;
  assign n25205 = n3476 & ~n25204;
  assign n25206 = ~n25197 & ~n25205;
  assign n25207 = n3374 & ~n25206;
  assign n25208 = ~n25189 & ~n25207;
  assign n25209 = n3655 & ~n25208;
  assign n25210 = ~n3378 & ~n9563;
  assign n25211 = n3492 & ~n25210;
  assign n25212 = ~n3493 & ~n25211;
  assign n25213 = n3485 & ~n25212;
  assign n25214 = ~n3486 & ~n25213;
  assign n25215 = ~n3476 & ~n25214;
  assign n25216 = ~n3378 & ~n8490;
  assign n25217 = ~n3378 & ~n25216;
  assign n25218 = ~n3485 & ~n25217;
  assign n25219 = ~n3492 & ~n25217;
  assign n25220 = ~n25211 & ~n25219;
  assign n25221 = n3485 & ~n25220;
  assign n25222 = ~n25218 & ~n25221;
  assign n25223 = n3476 & ~n25222;
  assign n25224 = ~n25215 & ~n25223;
  assign n25225 = ~n3374 & ~n25224;
  assign n25226 = ~n3281 & ~n9621;
  assign n25227 = n3378 & ~n25226;
  assign n25228 = ~n9623 & ~n25227;
  assign n25229 = n3492 & ~n25228;
  assign n25230 = ~n25115 & ~n25229;
  assign n25231 = n3485 & ~n25230;
  assign n25232 = ~n25114 & ~n25231;
  assign n25233 = ~n3476 & ~n25232;
  assign n25234 = n3378 & ~n8618;
  assign n25235 = ~n25216 & ~n25234;
  assign n25236 = ~n3485 & ~n25235;
  assign n25237 = ~n3492 & ~n25235;
  assign n25238 = ~n24548 & ~n25237;
  assign n25239 = n3485 & ~n25238;
  assign n25240 = ~n25236 & ~n25239;
  assign n25241 = n3476 & ~n25240;
  assign n25242 = ~n25233 & ~n25241;
  assign n25243 = n3374 & ~n25242;
  assign n25244 = ~n25225 & ~n25243;
  assign n25245 = ~n3655 & ~n25244;
  assign n25246 = ~n25209 & ~n25245;
  assign n25247 = ~n3652 & ~n25246;
  assign n25248 = ~n25173 & ~n25247;
  assign n25249 = ~n3368 & ~n25248;
  assign n25250 = ~n3378 & ~n9757;
  assign n25251 = n3492 & ~n25250;
  assign n25252 = n3492 & ~n25251;
  assign n25253 = n3485 & ~n25252;
  assign n25254 = n3485 & ~n25253;
  assign n25255 = ~n3476 & ~n25254;
  assign n25256 = ~n3378 & ~n8522;
  assign n25257 = ~n3378 & ~n25256;
  assign n25258 = ~n3485 & ~n25257;
  assign n25259 = ~n3492 & ~n25257;
  assign n25260 = ~n25251 & ~n25259;
  assign n25261 = n3485 & ~n25260;
  assign n25262 = ~n25258 & ~n25261;
  assign n25263 = n3476 & ~n25262;
  assign n25264 = ~n25255 & ~n25263;
  assign n25265 = ~n3374 & ~n25264;
  assign n25266 = ~n25038 & ~n25265;
  assign n25267 = n3655 & ~n25266;
  assign n25268 = ~n3378 & ~n10299;
  assign n25269 = n3492 & ~n25268;
  assign n25270 = n3492 & ~n25269;
  assign n25271 = n3485 & ~n25270;
  assign n25272 = n3485 & ~n25271;
  assign n25273 = ~n3476 & ~n25272;
  assign n25274 = ~n25259 & ~n25269;
  assign n25275 = n3485 & ~n25274;
  assign n25276 = ~n25258 & ~n25275;
  assign n25277 = n3476 & ~n25276;
  assign n25278 = ~n25273 & ~n25277;
  assign n25279 = ~n3374 & ~n25278;
  assign n25280 = ~n25052 & ~n25279;
  assign n25281 = ~n3655 & ~n25280;
  assign n25282 = ~n25267 & ~n25281;
  assign n25283 = n3652 & ~n25282;
  assign n25284 = ~n3378 & ~n10742;
  assign n25285 = n3492 & ~n25284;
  assign n25286 = n3492 & ~n25285;
  assign n25287 = n3485 & ~n25286;
  assign n25288 = n3485 & ~n25287;
  assign n25289 = ~n3476 & ~n25288;
  assign n25290 = ~n25259 & ~n25285;
  assign n25291 = n3485 & ~n25290;
  assign n25292 = ~n25258 & ~n25291;
  assign n25293 = n3476 & ~n25292;
  assign n25294 = ~n25289 & ~n25293;
  assign n25295 = ~n3374 & ~n25294;
  assign n25296 = ~n25068 & ~n25295;
  assign n25297 = n3655 & ~n25296;
  assign n25298 = ~n3378 & ~n11178;
  assign n25299 = n3492 & ~n25298;
  assign n25300 = n3492 & ~n25299;
  assign n25301 = n3485 & ~n25300;
  assign n25302 = n3485 & ~n25301;
  assign n25303 = ~n3476 & ~n25302;
  assign n25304 = ~n25259 & ~n25299;
  assign n25305 = n3485 & ~n25304;
  assign n25306 = ~n25258 & ~n25305;
  assign n25307 = n3476 & ~n25306;
  assign n25308 = ~n25303 & ~n25307;
  assign n25309 = ~n3374 & ~n25308;
  assign n25310 = ~n25082 & ~n25309;
  assign n25311 = ~n3655 & ~n25310;
  assign n25312 = ~n25297 & ~n25311;
  assign n25313 = ~n3652 & ~n25312;
  assign n25314 = ~n25283 & ~n25313;
  assign n25315 = n3368 & ~n25314;
  assign n25316 = ~n25249 & ~n25315;
  assign n25317 = ~n3362 & ~n25316;
  assign n25318 = ~n3362 & ~n25317;
  assign n25319 = ~n3359 & ~n25318;
  assign n25320 = ~n3359 & ~n25319;
  assign n25321 = n3356 & ~n25320;
  assign n25322 = ~n3356 & ~n25089;
  assign n25323 = ~n25321 & ~n25322;
  assign n25324 = n3345 & ~n25323;
  assign n25325 = ~n25096 & ~n25324;
  assign n25326 = n3341 & ~n25325;
  assign n25327 = ~n24366 & ~n25326;
  assign n25328 = n3337 & ~n25327;
  assign n25329 = ~n17220 & ~n25328;
  assign n25330 = n3280 & ~n25329;
  assign n25331 = controllable_hgrant3 & ~n3942;
  assign n25332 = ~n3898 & ~n25331;
  assign n25333 = controllable_nhgrant0 & ~n25332;
  assign n25334 = ~n3945 & ~n25333;
  assign n25335 = ~n3281 & ~n25334;
  assign n25336 = ~n3281 & ~n25335;
  assign n25337 = n3378 & ~n25336;
  assign n25338 = controllable_hgrant3 & ~n3984;
  assign n25339 = ~n3971 & ~n25338;
  assign n25340 = controllable_nhgrant0 & ~n25339;
  assign n25341 = ~n3987 & ~n25340;
  assign n25342 = ~n3281 & ~n25341;
  assign n25343 = ~n3950 & ~n25342;
  assign n25344 = ~n3378 & ~n25343;
  assign n25345 = ~n25337 & ~n25344;
  assign n25346 = n3492 & ~n25345;
  assign n25347 = ~n3493 & ~n25346;
  assign n25348 = n3485 & ~n25347;
  assign n25349 = ~n3486 & ~n25348;
  assign n25350 = ~n3476 & ~n25349;
  assign n25351 = ~n4082 & ~n25331;
  assign n25352 = controllable_nhgrant0 & ~n25351;
  assign n25353 = ~n3945 & ~n25352;
  assign n25354 = ~n3281 & ~n25353;
  assign n25355 = ~n3281 & ~n25354;
  assign n25356 = n3378 & ~n25355;
  assign n25357 = ~n4161 & ~n25338;
  assign n25358 = controllable_nhgrant0 & ~n25357;
  assign n25359 = ~n3987 & ~n25358;
  assign n25360 = ~n3281 & ~n25359;
  assign n25361 = ~n4089 & ~n25360;
  assign n25362 = ~n3378 & ~n25361;
  assign n25363 = ~n25356 & ~n25362;
  assign n25364 = n3492 & ~n25363;
  assign n25365 = ~n3493 & ~n25364;
  assign n25366 = n3485 & ~n25365;
  assign n25367 = ~n3486 & ~n25366;
  assign n25368 = n3476 & ~n25367;
  assign n25369 = ~n25350 & ~n25368;
  assign n25370 = n3374 & ~n25369;
  assign n25371 = ~n3820 & ~n25370;
  assign n25372 = n3655 & ~n25371;
  assign n25373 = ~n4218 & ~n25331;
  assign n25374 = controllable_nhgrant0 & ~n25373;
  assign n25375 = ~n3945 & ~n25374;
  assign n25376 = ~n3281 & ~n25375;
  assign n25377 = ~n3281 & ~n25376;
  assign n25378 = n3378 & ~n25377;
  assign n25379 = ~n4236 & ~n25338;
  assign n25380 = controllable_nhgrant0 & ~n25379;
  assign n25381 = ~n3987 & ~n25380;
  assign n25382 = ~n3281 & ~n25381;
  assign n25383 = ~n3950 & ~n25382;
  assign n25384 = ~n3378 & ~n25383;
  assign n25385 = ~n25378 & ~n25384;
  assign n25386 = n3492 & ~n25385;
  assign n25387 = ~n3493 & ~n25386;
  assign n25388 = n3485 & ~n25387;
  assign n25389 = ~n3486 & ~n25388;
  assign n25390 = ~n3476 & ~n25389;
  assign n25391 = ~n4271 & ~n25331;
  assign n25392 = controllable_nhgrant0 & ~n25391;
  assign n25393 = ~n3945 & ~n25392;
  assign n25394 = ~n3281 & ~n25393;
  assign n25395 = ~n3281 & ~n25394;
  assign n25396 = n3378 & ~n25395;
  assign n25397 = ~n4314 & ~n25338;
  assign n25398 = controllable_nhgrant0 & ~n25397;
  assign n25399 = ~n3987 & ~n25398;
  assign n25400 = ~n3281 & ~n25399;
  assign n25401 = ~n4089 & ~n25400;
  assign n25402 = ~n3378 & ~n25401;
  assign n25403 = ~n25396 & ~n25402;
  assign n25404 = n3492 & ~n25403;
  assign n25405 = ~n3493 & ~n25404;
  assign n25406 = n3485 & ~n25405;
  assign n25407 = ~n3486 & ~n25406;
  assign n25408 = n3476 & ~n25407;
  assign n25409 = ~n25390 & ~n25408;
  assign n25410 = n3374 & ~n25409;
  assign n25411 = ~n3820 & ~n25410;
  assign n25412 = ~n3655 & ~n25411;
  assign n25413 = ~n25372 & ~n25412;
  assign n25414 = n3652 & ~n25413;
  assign n25415 = ~n4350 & ~n25331;
  assign n25416 = controllable_nhgrant0 & ~n25415;
  assign n25417 = ~n3945 & ~n25416;
  assign n25418 = ~n3281 & ~n25417;
  assign n25419 = ~n3281 & ~n25418;
  assign n25420 = n3378 & ~n25419;
  assign n25421 = ~n4368 & ~n25338;
  assign n25422 = controllable_nhgrant0 & ~n25421;
  assign n25423 = ~n3987 & ~n25422;
  assign n25424 = ~n3281 & ~n25423;
  assign n25425 = ~n3950 & ~n25424;
  assign n25426 = ~n3378 & ~n25425;
  assign n25427 = ~n25420 & ~n25426;
  assign n25428 = n3492 & ~n25427;
  assign n25429 = ~n3493 & ~n25428;
  assign n25430 = n3485 & ~n25429;
  assign n25431 = ~n3486 & ~n25430;
  assign n25432 = ~n3476 & ~n25431;
  assign n25433 = ~n4396 & ~n25331;
  assign n25434 = controllable_nhgrant0 & ~n25433;
  assign n25435 = ~n3945 & ~n25434;
  assign n25436 = ~n3281 & ~n25435;
  assign n25437 = ~n3281 & ~n25436;
  assign n25438 = n3378 & ~n25437;
  assign n25439 = ~n4418 & ~n25338;
  assign n25440 = controllable_nhgrant0 & ~n25439;
  assign n25441 = ~n3987 & ~n25440;
  assign n25442 = ~n3281 & ~n25441;
  assign n25443 = ~n4089 & ~n25442;
  assign n25444 = ~n3378 & ~n25443;
  assign n25445 = ~n25438 & ~n25444;
  assign n25446 = n3492 & ~n25445;
  assign n25447 = ~n3493 & ~n25446;
  assign n25448 = n3485 & ~n25447;
  assign n25449 = ~n3486 & ~n25448;
  assign n25450 = n3476 & ~n25449;
  assign n25451 = ~n25432 & ~n25450;
  assign n25452 = n3374 & ~n25451;
  assign n25453 = ~n3820 & ~n25452;
  assign n25454 = n3655 & ~n25453;
  assign n25455 = ~n4450 & ~n25331;
  assign n25456 = controllable_nhgrant0 & ~n25455;
  assign n25457 = ~n3945 & ~n25456;
  assign n25458 = ~n3281 & ~n25457;
  assign n25459 = ~n3281 & ~n25458;
  assign n25460 = n3378 & ~n25459;
  assign n25461 = ~n4468 & ~n25338;
  assign n25462 = controllable_nhgrant0 & ~n25461;
  assign n25463 = ~n3987 & ~n25462;
  assign n25464 = ~n3281 & ~n25463;
  assign n25465 = ~n3950 & ~n25464;
  assign n25466 = ~n3378 & ~n25465;
  assign n25467 = ~n25460 & ~n25466;
  assign n25468 = n3492 & ~n25467;
  assign n25469 = ~n3493 & ~n25468;
  assign n25470 = n3485 & ~n25469;
  assign n25471 = ~n3486 & ~n25470;
  assign n25472 = ~n3476 & ~n25471;
  assign n25473 = ~n4496 & ~n25331;
  assign n25474 = controllable_nhgrant0 & ~n25473;
  assign n25475 = ~n3945 & ~n25474;
  assign n25476 = ~n3281 & ~n25475;
  assign n25477 = ~n3281 & ~n25476;
  assign n25478 = n3378 & ~n25477;
  assign n25479 = ~n4518 & ~n25338;
  assign n25480 = controllable_nhgrant0 & ~n25479;
  assign n25481 = ~n3987 & ~n25480;
  assign n25482 = ~n3281 & ~n25481;
  assign n25483 = ~n4089 & ~n25482;
  assign n25484 = ~n3378 & ~n25483;
  assign n25485 = ~n25478 & ~n25484;
  assign n25486 = n3492 & ~n25485;
  assign n25487 = ~n3493 & ~n25486;
  assign n25488 = n3485 & ~n25487;
  assign n25489 = ~n3486 & ~n25488;
  assign n25490 = n3476 & ~n25489;
  assign n25491 = ~n25472 & ~n25490;
  assign n25492 = n3374 & ~n25491;
  assign n25493 = ~n3820 & ~n25492;
  assign n25494 = ~n3655 & ~n25493;
  assign n25495 = ~n25454 & ~n25494;
  assign n25496 = ~n3652 & ~n25495;
  assign n25497 = ~n25414 & ~n25496;
  assign n25498 = ~n3368 & ~n25497;
  assign n25499 = controllable_hgrant3 & ~n4643;
  assign n25500 = ~n4599 & ~n25499;
  assign n25501 = controllable_nhgrant0 & ~n25500;
  assign n25502 = ~n4646 & ~n25501;
  assign n25503 = ~n3281 & ~n25502;
  assign n25504 = ~n3281 & ~n25503;
  assign n25505 = n3492 & ~n25504;
  assign n25506 = n3492 & ~n25505;
  assign n25507 = n3485 & ~n25506;
  assign n25508 = n3485 & ~n25507;
  assign n25509 = ~n3476 & ~n25508;
  assign n25510 = ~n4682 & ~n25499;
  assign n25511 = controllable_nhgrant0 & ~n25510;
  assign n25512 = ~n4646 & ~n25511;
  assign n25513 = ~n3281 & ~n25512;
  assign n25514 = ~n3281 & ~n25513;
  assign n25515 = n3492 & ~n25514;
  assign n25516 = n3492 & ~n25515;
  assign n25517 = n3485 & ~n25516;
  assign n25518 = n3485 & ~n25517;
  assign n25519 = n3476 & ~n25518;
  assign n25520 = ~n25509 & ~n25519;
  assign n25521 = n3374 & ~n25520;
  assign n25522 = n3374 & ~n25521;
  assign n25523 = n3655 & ~n25522;
  assign n25524 = ~n4737 & ~n25499;
  assign n25525 = controllable_nhgrant0 & ~n25524;
  assign n25526 = ~n4646 & ~n25525;
  assign n25527 = ~n3281 & ~n25526;
  assign n25528 = ~n3281 & ~n25527;
  assign n25529 = n3492 & ~n25528;
  assign n25530 = n3492 & ~n25529;
  assign n25531 = n3485 & ~n25530;
  assign n25532 = n3485 & ~n25531;
  assign n25533 = ~n3476 & ~n25532;
  assign n25534 = ~n4770 & ~n25499;
  assign n25535 = controllable_nhgrant0 & ~n25534;
  assign n25536 = ~n4646 & ~n25535;
  assign n25537 = ~n3281 & ~n25536;
  assign n25538 = ~n3281 & ~n25537;
  assign n25539 = n3492 & ~n25538;
  assign n25540 = n3492 & ~n25539;
  assign n25541 = n3485 & ~n25540;
  assign n25542 = n3485 & ~n25541;
  assign n25543 = n3476 & ~n25542;
  assign n25544 = ~n25533 & ~n25543;
  assign n25545 = n3374 & ~n25544;
  assign n25546 = n3374 & ~n25545;
  assign n25547 = ~n3655 & ~n25546;
  assign n25548 = ~n25523 & ~n25547;
  assign n25549 = n3652 & ~n25548;
  assign n25550 = ~n4804 & ~n25499;
  assign n25551 = controllable_nhgrant0 & ~n25550;
  assign n25552 = ~n4646 & ~n25551;
  assign n25553 = ~n3281 & ~n25552;
  assign n25554 = ~n3281 & ~n25553;
  assign n25555 = n3492 & ~n25554;
  assign n25556 = n3492 & ~n25555;
  assign n25557 = n3485 & ~n25556;
  assign n25558 = n3485 & ~n25557;
  assign n25559 = ~n3476 & ~n25558;
  assign n25560 = ~n4830 & ~n25499;
  assign n25561 = controllable_nhgrant0 & ~n25560;
  assign n25562 = ~n4646 & ~n25561;
  assign n25563 = ~n3281 & ~n25562;
  assign n25564 = ~n3281 & ~n25563;
  assign n25565 = n3492 & ~n25564;
  assign n25566 = n3492 & ~n25565;
  assign n25567 = n3485 & ~n25566;
  assign n25568 = n3485 & ~n25567;
  assign n25569 = n3476 & ~n25568;
  assign n25570 = ~n25559 & ~n25569;
  assign n25571 = n3374 & ~n25570;
  assign n25572 = n3374 & ~n25571;
  assign n25573 = n3655 & ~n25572;
  assign n25574 = ~n4860 & ~n25499;
  assign n25575 = controllable_nhgrant0 & ~n25574;
  assign n25576 = ~n4646 & ~n25575;
  assign n25577 = ~n3281 & ~n25576;
  assign n25578 = ~n3281 & ~n25577;
  assign n25579 = n3492 & ~n25578;
  assign n25580 = n3492 & ~n25579;
  assign n25581 = n3485 & ~n25580;
  assign n25582 = n3485 & ~n25581;
  assign n25583 = ~n3476 & ~n25582;
  assign n25584 = ~n4886 & ~n25499;
  assign n25585 = controllable_nhgrant0 & ~n25584;
  assign n25586 = ~n4646 & ~n25585;
  assign n25587 = ~n3281 & ~n25586;
  assign n25588 = ~n3281 & ~n25587;
  assign n25589 = n3492 & ~n25588;
  assign n25590 = n3492 & ~n25589;
  assign n25591 = n3485 & ~n25590;
  assign n25592 = n3485 & ~n25591;
  assign n25593 = n3476 & ~n25592;
  assign n25594 = ~n25583 & ~n25593;
  assign n25595 = n3374 & ~n25594;
  assign n25596 = n3374 & ~n25595;
  assign n25597 = ~n3655 & ~n25596;
  assign n25598 = ~n25573 & ~n25597;
  assign n25599 = ~n3652 & ~n25598;
  assign n25600 = ~n25549 & ~n25599;
  assign n25601 = n3368 & ~n25600;
  assign n25602 = ~n25498 & ~n25601;
  assign n25603 = ~n3362 & ~n25602;
  assign n25604 = ~n3362 & ~n25603;
  assign n25605 = ~n3359 & ~n25604;
  assign n25606 = ~n3359 & ~n25605;
  assign n25607 = n3356 & ~n25606;
  assign n25608 = ~controllable_hgrant2 & ~n6592;
  assign n25609 = ~n4920 & ~n25608;
  assign n25610 = controllable_hmaster0 & ~n25609;
  assign n25611 = ~n4930 & ~n25610;
  assign n25612 = controllable_hmaster1 & ~n25611;
  assign n25613 = ~n4946 & ~n25612;
  assign n25614 = i_hlock3 & ~n25613;
  assign n25615 = ~controllable_hgrant2 & ~n6595;
  assign n25616 = ~n4949 & ~n25615;
  assign n25617 = controllable_hmaster0 & ~n25616;
  assign n25618 = ~n4930 & ~n25617;
  assign n25619 = controllable_hmaster1 & ~n25618;
  assign n25620 = ~n4946 & ~n25619;
  assign n25621 = ~i_hlock3 & ~n25620;
  assign n25622 = ~n25614 & ~n25621;
  assign n25623 = i_hbusreq3 & ~n25622;
  assign n25624 = i_hbusreq2 & ~n6592;
  assign n25625 = ~i_hbusreq2 & ~n6624;
  assign n25626 = ~n25624 & ~n25625;
  assign n25627 = ~controllable_hgrant2 & ~n25626;
  assign n25628 = ~n4968 & ~n25627;
  assign n25629 = controllable_hmaster0 & ~n25628;
  assign n25630 = ~n4990 & ~n25629;
  assign n25631 = controllable_hmaster1 & ~n25630;
  assign n25632 = ~n5009 & ~n25631;
  assign n25633 = i_hlock3 & ~n25632;
  assign n25634 = i_hbusreq2 & ~n6595;
  assign n25635 = ~i_hbusreq2 & ~n6638;
  assign n25636 = ~n25634 & ~n25635;
  assign n25637 = ~controllable_hgrant2 & ~n25636;
  assign n25638 = ~n5015 & ~n25637;
  assign n25639 = controllable_hmaster0 & ~n25638;
  assign n25640 = ~n4990 & ~n25639;
  assign n25641 = controllable_hmaster1 & ~n25640;
  assign n25642 = ~n5009 & ~n25641;
  assign n25643 = ~i_hlock3 & ~n25642;
  assign n25644 = ~n25633 & ~n25643;
  assign n25645 = ~i_hbusreq3 & ~n25644;
  assign n25646 = ~n25623 & ~n25645;
  assign n25647 = ~controllable_hmaster2 & ~n25646;
  assign n25648 = ~n5203 & ~n25647;
  assign n25649 = controllable_hgrant3 & ~n25648;
  assign n25650 = ~n5163 & ~n25649;
  assign n25651 = controllable_nhgrant0 & ~n25650;
  assign n25652 = ~n5245 & ~n25651;
  assign n25653 = ~n3281 & ~n25652;
  assign n25654 = ~n3783 & ~n25653;
  assign n25655 = ~n3378 & ~n25654;
  assign n25656 = ~n4911 & ~n25655;
  assign n25657 = n3492 & ~n25656;
  assign n25658 = ~n3631 & ~n25657;
  assign n25659 = n3485 & ~n25658;
  assign n25660 = ~n3630 & ~n25659;
  assign n25661 = ~n3374 & ~n25660;
  assign n25662 = ~n3983 & ~n5285;
  assign n25663 = controllable_hgrant3 & ~n25662;
  assign n25664 = ~n5340 & ~n25663;
  assign n25665 = controllable_nhgrant0 & ~n25664;
  assign n25666 = ~n5363 & ~n25665;
  assign n25667 = ~n3281 & ~n25666;
  assign n25668 = ~n3950 & ~n25667;
  assign n25669 = n3378 & ~n25668;
  assign n25670 = ~n3910 & ~n5046;
  assign n25671 = controllable_hmaster1 & ~n25670;
  assign n25672 = ~controllable_hmaster1 & ~n3909;
  assign n25673 = ~n25671 & ~n25672;
  assign n25674 = i_hbusreq3 & ~n25673;
  assign n25675 = ~n3935 & ~n5071;
  assign n25676 = controllable_hmaster1 & ~n25675;
  assign n25677 = ~n5197 & ~n5478;
  assign n25678 = ~controllable_hmaster1 & ~n25677;
  assign n25679 = ~n25676 & ~n25678;
  assign n25680 = ~i_hbusreq3 & ~n25679;
  assign n25681 = ~n25674 & ~n25680;
  assign n25682 = ~controllable_hmaster2 & ~n25681;
  assign n25683 = ~n5498 & ~n25682;
  assign n25684 = controllable_hgrant3 & ~n25683;
  assign n25685 = ~n5486 & ~n25684;
  assign n25686 = controllable_nhgrant0 & ~n25685;
  assign n25687 = ~n5534 & ~n25686;
  assign n25688 = ~n3281 & ~n25687;
  assign n25689 = ~n3950 & ~n25688;
  assign n25690 = ~n3378 & ~n25689;
  assign n25691 = ~n25669 & ~n25690;
  assign n25692 = n3492 & ~n25691;
  assign n25693 = ~n3631 & ~n25692;
  assign n25694 = n3485 & ~n25693;
  assign n25695 = ~n3630 & ~n25694;
  assign n25696 = ~n3476 & ~n25695;
  assign n25697 = ~n5613 & ~n5793;
  assign n25698 = controllable_hgrant3 & ~n25697;
  assign n25699 = ~n5754 & ~n25698;
  assign n25700 = controllable_nhgrant0 & ~n25699;
  assign n25701 = ~n5809 & ~n25700;
  assign n25702 = ~n3281 & ~n25701;
  assign n25703 = ~n4089 & ~n25702;
  assign n25704 = n3378 & ~n25703;
  assign n25705 = controllable_hmaster0 & ~n6043;
  assign n25706 = ~n9062 & ~n25705;
  assign n25707 = controllable_hmaster1 & ~n25706;
  assign n25708 = ~controllable_hmaster1 & ~n6012;
  assign n25709 = ~n25707 & ~n25708;
  assign n25710 = i_hbusreq3 & ~n25709;
  assign n25711 = ~controllable_hgrant2 & ~n6812;
  assign n25712 = ~n3859 & ~n25711;
  assign n25713 = controllable_hmaster0 & ~n25712;
  assign n25714 = ~n9086 & ~n25713;
  assign n25715 = controllable_hmaster1 & ~n25714;
  assign n25716 = ~controllable_hgrant2 & ~n6830;
  assign n25717 = ~n5461 & ~n25716;
  assign n25718 = ~controllable_hmaster0 & ~n25717;
  assign n25719 = ~n6050 & ~n25718;
  assign n25720 = ~controllable_hmaster1 & ~n25719;
  assign n25721 = ~n25715 & ~n25720;
  assign n25722 = ~i_hbusreq3 & ~n25721;
  assign n25723 = ~n25710 & ~n25722;
  assign n25724 = ~controllable_hmaster2 & ~n25723;
  assign n25725 = ~n6035 & ~n25724;
  assign n25726 = controllable_hgrant3 & ~n25725;
  assign n25727 = ~n6004 & ~n25726;
  assign n25728 = controllable_nhgrant0 & ~n25727;
  assign n25729 = ~n6082 & ~n25728;
  assign n25730 = ~n3281 & ~n25729;
  assign n25731 = ~n4089 & ~n25730;
  assign n25732 = ~n3378 & ~n25731;
  assign n25733 = ~n25704 & ~n25732;
  assign n25734 = n3492 & ~n25733;
  assign n25735 = ~n3631 & ~n25734;
  assign n25736 = n3485 & ~n25735;
  assign n25737 = ~n3630 & ~n25736;
  assign n25738 = n3476 & ~n25737;
  assign n25739 = ~n25696 & ~n25738;
  assign n25740 = n3374 & ~n25739;
  assign n25741 = ~n25661 & ~n25740;
  assign n25742 = n3655 & ~n25741;
  assign n25743 = ~n6190 & ~n25649;
  assign n25744 = controllable_nhgrant0 & ~n25743;
  assign n25745 = ~n5245 & ~n25744;
  assign n25746 = ~n3281 & ~n25745;
  assign n25747 = ~n3783 & ~n25746;
  assign n25748 = ~n3378 & ~n25747;
  assign n25749 = ~n4911 & ~n25748;
  assign n25750 = n3492 & ~n25749;
  assign n25751 = ~n3631 & ~n25750;
  assign n25752 = n3485 & ~n25751;
  assign n25753 = ~n3630 & ~n25752;
  assign n25754 = ~n3374 & ~n25753;
  assign n25755 = ~n6204 & ~n25663;
  assign n25756 = controllable_nhgrant0 & ~n25755;
  assign n25757 = ~n5363 & ~n25756;
  assign n25758 = ~n3281 & ~n25757;
  assign n25759 = ~n3950 & ~n25758;
  assign n25760 = n3378 & ~n25759;
  assign n25761 = ~n6345 & ~n25684;
  assign n25762 = controllable_nhgrant0 & ~n25761;
  assign n25763 = ~n5534 & ~n25762;
  assign n25764 = ~n3281 & ~n25763;
  assign n25765 = ~n3950 & ~n25764;
  assign n25766 = ~n3378 & ~n25765;
  assign n25767 = ~n25760 & ~n25766;
  assign n25768 = n3492 & ~n25767;
  assign n25769 = ~n3631 & ~n25768;
  assign n25770 = n3485 & ~n25769;
  assign n25771 = ~n3630 & ~n25770;
  assign n25772 = ~n3476 & ~n25771;
  assign n25773 = ~n6394 & ~n25698;
  assign n25774 = controllable_nhgrant0 & ~n25773;
  assign n25775 = ~n5809 & ~n25774;
  assign n25776 = ~n3281 & ~n25775;
  assign n25777 = ~n4089 & ~n25776;
  assign n25778 = n3378 & ~n25777;
  assign n25779 = ~n6556 & ~n25726;
  assign n25780 = controllable_nhgrant0 & ~n25779;
  assign n25781 = ~n6082 & ~n25780;
  assign n25782 = ~n3281 & ~n25781;
  assign n25783 = ~n4089 & ~n25782;
  assign n25784 = ~n3378 & ~n25783;
  assign n25785 = ~n25778 & ~n25784;
  assign n25786 = n3492 & ~n25785;
  assign n25787 = ~n3631 & ~n25786;
  assign n25788 = n3485 & ~n25787;
  assign n25789 = ~n3630 & ~n25788;
  assign n25790 = n3476 & ~n25789;
  assign n25791 = ~n25772 & ~n25790;
  assign n25792 = n3374 & ~n25791;
  assign n25793 = ~n25754 & ~n25792;
  assign n25794 = ~n3655 & ~n25793;
  assign n25795 = ~n25742 & ~n25794;
  assign n25796 = n3652 & ~n25795;
  assign n25797 = ~n6659 & ~n25649;
  assign n25798 = controllable_nhgrant0 & ~n25797;
  assign n25799 = ~n5245 & ~n25798;
  assign n25800 = ~n3281 & ~n25799;
  assign n25801 = ~n3783 & ~n25800;
  assign n25802 = ~n3378 & ~n25801;
  assign n25803 = ~n4911 & ~n25802;
  assign n25804 = n3492 & ~n25803;
  assign n25805 = ~n3631 & ~n25804;
  assign n25806 = n3485 & ~n25805;
  assign n25807 = ~n3630 & ~n25806;
  assign n25808 = ~n3374 & ~n25807;
  assign n25809 = ~n6673 & ~n25663;
  assign n25810 = controllable_nhgrant0 & ~n25809;
  assign n25811 = ~n5363 & ~n25810;
  assign n25812 = ~n3281 & ~n25811;
  assign n25813 = ~n3950 & ~n25812;
  assign n25814 = n3378 & ~n25813;
  assign n25815 = ~n6725 & ~n25684;
  assign n25816 = controllable_nhgrant0 & ~n25815;
  assign n25817 = ~n5534 & ~n25816;
  assign n25818 = ~n3281 & ~n25817;
  assign n25819 = ~n3950 & ~n25818;
  assign n25820 = ~n3378 & ~n25819;
  assign n25821 = ~n25814 & ~n25820;
  assign n25822 = n3492 & ~n25821;
  assign n25823 = ~n3631 & ~n25822;
  assign n25824 = n3485 & ~n25823;
  assign n25825 = ~n3630 & ~n25824;
  assign n25826 = ~n3476 & ~n25825;
  assign n25827 = ~n6755 & ~n25698;
  assign n25828 = controllable_nhgrant0 & ~n25827;
  assign n25829 = ~n5809 & ~n25828;
  assign n25830 = ~n3281 & ~n25829;
  assign n25831 = ~n4089 & ~n25830;
  assign n25832 = n3378 & ~n25831;
  assign n25833 = ~n6841 & ~n25726;
  assign n25834 = controllable_nhgrant0 & ~n25833;
  assign n25835 = ~n6082 & ~n25834;
  assign n25836 = ~n3281 & ~n25835;
  assign n25837 = ~n4089 & ~n25836;
  assign n25838 = ~n3378 & ~n25837;
  assign n25839 = ~n25832 & ~n25838;
  assign n25840 = n3492 & ~n25839;
  assign n25841 = ~n3631 & ~n25840;
  assign n25842 = n3485 & ~n25841;
  assign n25843 = ~n3630 & ~n25842;
  assign n25844 = n3476 & ~n25843;
  assign n25845 = ~n25826 & ~n25844;
  assign n25846 = n3374 & ~n25845;
  assign n25847 = ~n25808 & ~n25846;
  assign n25848 = n3655 & ~n25847;
  assign n25849 = ~n6889 & ~n25649;
  assign n25850 = controllable_nhgrant0 & ~n25849;
  assign n25851 = ~n5245 & ~n25850;
  assign n25852 = ~n3281 & ~n25851;
  assign n25853 = ~n3783 & ~n25852;
  assign n25854 = ~n3378 & ~n25853;
  assign n25855 = ~n4911 & ~n25854;
  assign n25856 = n3492 & ~n25855;
  assign n25857 = ~n3631 & ~n25856;
  assign n25858 = n3485 & ~n25857;
  assign n25859 = ~n3630 & ~n25858;
  assign n25860 = ~n3374 & ~n25859;
  assign n25861 = ~n6903 & ~n25663;
  assign n25862 = controllable_nhgrant0 & ~n25861;
  assign n25863 = ~n5363 & ~n25862;
  assign n25864 = ~n3281 & ~n25863;
  assign n25865 = ~n3950 & ~n25864;
  assign n25866 = n3378 & ~n25865;
  assign n25867 = ~n6957 & ~n25684;
  assign n25868 = controllable_nhgrant0 & ~n25867;
  assign n25869 = ~n5534 & ~n25868;
  assign n25870 = ~n3281 & ~n25869;
  assign n25871 = ~n3950 & ~n25870;
  assign n25872 = ~n3378 & ~n25871;
  assign n25873 = ~n25866 & ~n25872;
  assign n25874 = n3492 & ~n25873;
  assign n25875 = ~n3631 & ~n25874;
  assign n25876 = n3485 & ~n25875;
  assign n25877 = ~n3630 & ~n25876;
  assign n25878 = ~n3476 & ~n25877;
  assign n25879 = ~n6985 & ~n25698;
  assign n25880 = controllable_nhgrant0 & ~n25879;
  assign n25881 = ~n5809 & ~n25880;
  assign n25882 = ~n3281 & ~n25881;
  assign n25883 = ~n4089 & ~n25882;
  assign n25884 = n3378 & ~n25883;
  assign n25885 = ~n7042 & ~n25726;
  assign n25886 = controllable_nhgrant0 & ~n25885;
  assign n25887 = ~n6082 & ~n25886;
  assign n25888 = ~n3281 & ~n25887;
  assign n25889 = ~n4089 & ~n25888;
  assign n25890 = ~n3378 & ~n25889;
  assign n25891 = ~n25884 & ~n25890;
  assign n25892 = n3492 & ~n25891;
  assign n25893 = ~n3631 & ~n25892;
  assign n25894 = n3485 & ~n25893;
  assign n25895 = ~n3630 & ~n25894;
  assign n25896 = n3476 & ~n25895;
  assign n25897 = ~n25878 & ~n25896;
  assign n25898 = n3374 & ~n25897;
  assign n25899 = ~n25860 & ~n25898;
  assign n25900 = ~n3655 & ~n25899;
  assign n25901 = ~n25848 & ~n25900;
  assign n25902 = ~n3652 & ~n25901;
  assign n25903 = ~n25796 & ~n25902;
  assign n25904 = ~n3368 & ~n25903;
  assign n25905 = controllable_hgrant3 & ~n7115;
  assign n25906 = ~n7102 & ~n25905;
  assign n25907 = controllable_nhgrant0 & ~n25906;
  assign n25908 = ~n7118 & ~n25907;
  assign n25909 = ~n3281 & ~n25908;
  assign n25910 = ~n3281 & ~n25909;
  assign n25911 = ~n3378 & ~n25910;
  assign n25912 = ~n7082 & ~n25911;
  assign n25913 = n3492 & ~n25912;
  assign n25914 = n3492 & ~n25913;
  assign n25915 = n3485 & ~n25914;
  assign n25916 = n3485 & ~n25915;
  assign n25917 = ~n3374 & ~n25916;
  assign n25918 = ~n5285 & ~n7162;
  assign n25919 = controllable_hgrant3 & ~n25918;
  assign n25920 = ~n7148 & ~n25919;
  assign n25921 = controllable_nhgrant0 & ~n25920;
  assign n25922 = ~n7166 & ~n25921;
  assign n25923 = ~n3281 & ~n25922;
  assign n25924 = ~n3281 & ~n25923;
  assign n25925 = n3378 & ~n25924;
  assign n25926 = ~n7204 & ~n25682;
  assign n25927 = controllable_hgrant3 & ~n25926;
  assign n25928 = ~n7190 & ~n25927;
  assign n25929 = controllable_nhgrant0 & ~n25928;
  assign n25930 = ~n7208 & ~n25929;
  assign n25931 = ~n3281 & ~n25930;
  assign n25932 = ~n3281 & ~n25931;
  assign n25933 = ~n3378 & ~n25932;
  assign n25934 = ~n25925 & ~n25933;
  assign n25935 = n3492 & ~n25934;
  assign n25936 = n3492 & ~n25935;
  assign n25937 = n3485 & ~n25936;
  assign n25938 = n3485 & ~n25937;
  assign n25939 = ~n3476 & ~n25938;
  assign n25940 = ~n5613 & ~n7428;
  assign n25941 = controllable_hgrant3 & ~n25940;
  assign n25942 = ~n7391 & ~n25941;
  assign n25943 = controllable_nhgrant0 & ~n25942;
  assign n25944 = ~n7432 & ~n25943;
  assign n25945 = ~n3281 & ~n25944;
  assign n25946 = ~n3281 & ~n25945;
  assign n25947 = n3378 & ~n25946;
  assign n25948 = ~n7664 & ~n25724;
  assign n25949 = controllable_hgrant3 & ~n25948;
  assign n25950 = ~n7628 & ~n25949;
  assign n25951 = controllable_nhgrant0 & ~n25950;
  assign n25952 = ~n7668 & ~n25951;
  assign n25953 = ~n3281 & ~n25952;
  assign n25954 = ~n3281 & ~n25953;
  assign n25955 = ~n3378 & ~n25954;
  assign n25956 = ~n25947 & ~n25955;
  assign n25957 = n3492 & ~n25956;
  assign n25958 = n3492 & ~n25957;
  assign n25959 = n3485 & ~n25958;
  assign n25960 = n3485 & ~n25959;
  assign n25961 = n3476 & ~n25960;
  assign n25962 = ~n25939 & ~n25961;
  assign n25963 = n3374 & ~n25962;
  assign n25964 = ~n25917 & ~n25963;
  assign n25965 = n3655 & ~n25964;
  assign n25966 = ~n7694 & ~n25905;
  assign n25967 = controllable_nhgrant0 & ~n25966;
  assign n25968 = ~n7118 & ~n25967;
  assign n25969 = ~n3281 & ~n25968;
  assign n25970 = ~n3281 & ~n25969;
  assign n25971 = ~n3378 & ~n25970;
  assign n25972 = ~n7082 & ~n25971;
  assign n25973 = n3492 & ~n25972;
  assign n25974 = n3492 & ~n25973;
  assign n25975 = n3485 & ~n25974;
  assign n25976 = n3485 & ~n25975;
  assign n25977 = ~n3374 & ~n25976;
  assign n25978 = ~n7718 & ~n25919;
  assign n25979 = controllable_nhgrant0 & ~n25978;
  assign n25980 = ~n7166 & ~n25979;
  assign n25981 = ~n3281 & ~n25980;
  assign n25982 = ~n3281 & ~n25981;
  assign n25983 = n3378 & ~n25982;
  assign n25984 = ~n7736 & ~n25927;
  assign n25985 = controllable_nhgrant0 & ~n25984;
  assign n25986 = ~n7208 & ~n25985;
  assign n25987 = ~n3281 & ~n25986;
  assign n25988 = ~n3281 & ~n25987;
  assign n25989 = ~n3378 & ~n25988;
  assign n25990 = ~n25983 & ~n25989;
  assign n25991 = n3492 & ~n25990;
  assign n25992 = n3492 & ~n25991;
  assign n25993 = n3485 & ~n25992;
  assign n25994 = n3485 & ~n25993;
  assign n25995 = ~n3476 & ~n25994;
  assign n25996 = ~n7785 & ~n25941;
  assign n25997 = controllable_nhgrant0 & ~n25996;
  assign n25998 = ~n7432 & ~n25997;
  assign n25999 = ~n3281 & ~n25998;
  assign n26000 = ~n3281 & ~n25999;
  assign n26001 = n3378 & ~n26000;
  assign n26002 = ~n7944 & ~n25949;
  assign n26003 = controllable_nhgrant0 & ~n26002;
  assign n26004 = ~n7668 & ~n26003;
  assign n26005 = ~n3281 & ~n26004;
  assign n26006 = ~n3281 & ~n26005;
  assign n26007 = ~n3378 & ~n26006;
  assign n26008 = ~n26001 & ~n26007;
  assign n26009 = n3492 & ~n26008;
  assign n26010 = n3492 & ~n26009;
  assign n26011 = n3485 & ~n26010;
  assign n26012 = n3485 & ~n26011;
  assign n26013 = n3476 & ~n26012;
  assign n26014 = ~n25995 & ~n26013;
  assign n26015 = n3374 & ~n26014;
  assign n26016 = ~n25977 & ~n26015;
  assign n26017 = ~n3655 & ~n26016;
  assign n26018 = ~n25965 & ~n26017;
  assign n26019 = n3652 & ~n26018;
  assign n26020 = ~n7974 & ~n25905;
  assign n26021 = controllable_nhgrant0 & ~n26020;
  assign n26022 = ~n7118 & ~n26021;
  assign n26023 = ~n3281 & ~n26022;
  assign n26024 = ~n3281 & ~n26023;
  assign n26025 = ~n3378 & ~n26024;
  assign n26026 = ~n7082 & ~n26025;
  assign n26027 = n3492 & ~n26026;
  assign n26028 = n3492 & ~n26027;
  assign n26029 = n3485 & ~n26028;
  assign n26030 = n3485 & ~n26029;
  assign n26031 = ~n3374 & ~n26030;
  assign n26032 = ~n7998 & ~n25919;
  assign n26033 = controllable_nhgrant0 & ~n26032;
  assign n26034 = ~n7166 & ~n26033;
  assign n26035 = ~n3281 & ~n26034;
  assign n26036 = ~n3281 & ~n26035;
  assign n26037 = n3378 & ~n26036;
  assign n26038 = ~n8016 & ~n25927;
  assign n26039 = controllable_nhgrant0 & ~n26038;
  assign n26040 = ~n7208 & ~n26039;
  assign n26041 = ~n3281 & ~n26040;
  assign n26042 = ~n3281 & ~n26041;
  assign n26043 = ~n3378 & ~n26042;
  assign n26044 = ~n26037 & ~n26043;
  assign n26045 = n3492 & ~n26044;
  assign n26046 = n3492 & ~n26045;
  assign n26047 = n3485 & ~n26046;
  assign n26048 = n3485 & ~n26047;
  assign n26049 = ~n3476 & ~n26048;
  assign n26050 = ~n8046 & ~n25941;
  assign n26051 = controllable_nhgrant0 & ~n26050;
  assign n26052 = ~n7432 & ~n26051;
  assign n26053 = ~n3281 & ~n26052;
  assign n26054 = ~n3281 & ~n26053;
  assign n26055 = n3378 & ~n26054;
  assign n26056 = ~n8105 & ~n25949;
  assign n26057 = controllable_nhgrant0 & ~n26056;
  assign n26058 = ~n7668 & ~n26057;
  assign n26059 = ~n3281 & ~n26058;
  assign n26060 = ~n3281 & ~n26059;
  assign n26061 = ~n3378 & ~n26060;
  assign n26062 = ~n26055 & ~n26061;
  assign n26063 = n3492 & ~n26062;
  assign n26064 = n3492 & ~n26063;
  assign n26065 = n3485 & ~n26064;
  assign n26066 = n3485 & ~n26065;
  assign n26067 = n3476 & ~n26066;
  assign n26068 = ~n26049 & ~n26067;
  assign n26069 = n3374 & ~n26068;
  assign n26070 = ~n26031 & ~n26069;
  assign n26071 = n3655 & ~n26070;
  assign n26072 = ~n8133 & ~n25905;
  assign n26073 = controllable_nhgrant0 & ~n26072;
  assign n26074 = ~n7118 & ~n26073;
  assign n26075 = ~n3281 & ~n26074;
  assign n26076 = ~n3281 & ~n26075;
  assign n26077 = ~n3378 & ~n26076;
  assign n26078 = ~n7082 & ~n26077;
  assign n26079 = n3492 & ~n26078;
  assign n26080 = n3492 & ~n26079;
  assign n26081 = n3485 & ~n26080;
  assign n26082 = n3485 & ~n26081;
  assign n26083 = ~n3374 & ~n26082;
  assign n26084 = ~n8157 & ~n25919;
  assign n26085 = controllable_nhgrant0 & ~n26084;
  assign n26086 = ~n7166 & ~n26085;
  assign n26087 = ~n3281 & ~n26086;
  assign n26088 = ~n3281 & ~n26087;
  assign n26089 = n3378 & ~n26088;
  assign n26090 = ~n8175 & ~n25927;
  assign n26091 = controllable_nhgrant0 & ~n26090;
  assign n26092 = ~n7208 & ~n26091;
  assign n26093 = ~n3281 & ~n26092;
  assign n26094 = ~n3281 & ~n26093;
  assign n26095 = ~n3378 & ~n26094;
  assign n26096 = ~n26089 & ~n26095;
  assign n26097 = n3492 & ~n26096;
  assign n26098 = n3492 & ~n26097;
  assign n26099 = n3485 & ~n26098;
  assign n26100 = n3485 & ~n26099;
  assign n26101 = ~n3476 & ~n26100;
  assign n26102 = ~n8203 & ~n25941;
  assign n26103 = controllable_nhgrant0 & ~n26102;
  assign n26104 = ~n7432 & ~n26103;
  assign n26105 = ~n3281 & ~n26104;
  assign n26106 = ~n3281 & ~n26105;
  assign n26107 = n3378 & ~n26106;
  assign n26108 = ~n8260 & ~n25949;
  assign n26109 = controllable_nhgrant0 & ~n26108;
  assign n26110 = ~n7668 & ~n26109;
  assign n26111 = ~n3281 & ~n26110;
  assign n26112 = ~n3281 & ~n26111;
  assign n26113 = ~n3378 & ~n26112;
  assign n26114 = ~n26107 & ~n26113;
  assign n26115 = n3492 & ~n26114;
  assign n26116 = n3492 & ~n26115;
  assign n26117 = n3485 & ~n26116;
  assign n26118 = n3485 & ~n26117;
  assign n26119 = n3476 & ~n26118;
  assign n26120 = ~n26101 & ~n26119;
  assign n26121 = n3374 & ~n26120;
  assign n26122 = ~n26083 & ~n26121;
  assign n26123 = ~n3655 & ~n26122;
  assign n26124 = ~n26071 & ~n26123;
  assign n26125 = ~n3652 & ~n26124;
  assign n26126 = ~n26019 & ~n26125;
  assign n26127 = n3368 & ~n26126;
  assign n26128 = ~n25904 & ~n26127;
  assign n26129 = n3362 & ~n26128;
  assign n26130 = n3492 & ~n25654;
  assign n26131 = ~n3631 & ~n26130;
  assign n26132 = n3485 & ~n26131;
  assign n26133 = ~n3630 & ~n26132;
  assign n26134 = ~n3476 & ~n26133;
  assign n26135 = controllable_hmaster0 & ~n25610;
  assign n26136 = controllable_hmaster1 & ~n26135;
  assign n26137 = ~n8289 & ~n26136;
  assign n26138 = i_hlock3 & ~n26137;
  assign n26139 = controllable_hmaster0 & ~n25617;
  assign n26140 = controllable_hmaster1 & ~n26139;
  assign n26141 = ~n8289 & ~n26140;
  assign n26142 = ~i_hlock3 & ~n26141;
  assign n26143 = ~n26138 & ~n26142;
  assign n26144 = i_hbusreq3 & ~n26143;
  assign n26145 = controllable_hmaster0 & ~n25629;
  assign n26146 = controllable_hmaster1 & ~n26145;
  assign n26147 = ~n8289 & ~n26146;
  assign n26148 = i_hlock3 & ~n26147;
  assign n26149 = controllable_hmaster0 & ~n25639;
  assign n26150 = controllable_hmaster1 & ~n26149;
  assign n26151 = ~n8289 & ~n26150;
  assign n26152 = ~i_hlock3 & ~n26151;
  assign n26153 = ~n26148 & ~n26152;
  assign n26154 = ~i_hbusreq3 & ~n26153;
  assign n26155 = ~n26144 & ~n26154;
  assign n26156 = ~controllable_hmaster2 & ~n26155;
  assign n26157 = ~n3407 & ~n26156;
  assign n26158 = controllable_hgrant3 & ~n26157;
  assign n26159 = ~n8289 & ~n11402;
  assign n26160 = i_hlock3 & ~n26159;
  assign n26161 = ~n8289 & ~n11406;
  assign n26162 = ~i_hlock3 & ~n26161;
  assign n26163 = ~n26160 & ~n26162;
  assign n26164 = i_hbusreq3 & ~n26163;
  assign n26165 = ~n8289 & ~n11412;
  assign n26166 = i_hlock3 & ~n26165;
  assign n26167 = ~n8289 & ~n11416;
  assign n26168 = ~i_hlock3 & ~n26167;
  assign n26169 = ~n26166 & ~n26168;
  assign n26170 = ~i_hbusreq3 & ~n26169;
  assign n26171 = ~n26164 & ~n26170;
  assign n26172 = ~controllable_hmaster2 & ~n26171;
  assign n26173 = ~n3461 & ~n26172;
  assign n26174 = ~controllable_hgrant3 & ~n26173;
  assign n26175 = ~n26158 & ~n26174;
  assign n26176 = controllable_nhgrant0 & ~n26175;
  assign n26177 = ~n3407 & ~n26172;
  assign n26178 = controllable_hgrant3 & ~n26177;
  assign n26179 = ~n8299 & ~n11402;
  assign n26180 = i_hlock3 & ~n26179;
  assign n26181 = ~n8299 & ~n11406;
  assign n26182 = ~i_hlock3 & ~n26181;
  assign n26183 = ~n26180 & ~n26182;
  assign n26184 = i_hbusreq3 & ~n26183;
  assign n26185 = ~n8299 & ~n11412;
  assign n26186 = i_hlock3 & ~n26185;
  assign n26187 = ~n8299 & ~n11416;
  assign n26188 = ~i_hlock3 & ~n26187;
  assign n26189 = ~n26186 & ~n26188;
  assign n26190 = ~i_hbusreq3 & ~n26189;
  assign n26191 = ~n26184 & ~n26190;
  assign n26192 = ~controllable_hmaster2 & ~n26191;
  assign n26193 = ~n3407 & ~n26192;
  assign n26194 = ~controllable_hgrant3 & ~n26193;
  assign n26195 = ~n26178 & ~n26194;
  assign n26196 = ~controllable_nhgrant0 & ~n26195;
  assign n26197 = ~n26176 & ~n26196;
  assign n26198 = ~n3281 & ~n26197;
  assign n26199 = ~n3783 & ~n26198;
  assign n26200 = ~n3492 & ~n26199;
  assign n26201 = ~n8310 & ~n26200;
  assign n26202 = ~n3485 & ~n26201;
  assign n26203 = ~n26132 & ~n26202;
  assign n26204 = n3476 & ~n26203;
  assign n26205 = ~n26134 & ~n26204;
  assign n26206 = ~n3374 & ~n26205;
  assign n26207 = n3492 & ~n25689;
  assign n26208 = ~n3631 & ~n26207;
  assign n26209 = n3485 & ~n26208;
  assign n26210 = ~n3630 & ~n26209;
  assign n26211 = ~n3476 & ~n26210;
  assign n26212 = n3492 & ~n25731;
  assign n26213 = ~n3631 & ~n26212;
  assign n26214 = n3485 & ~n26213;
  assign n26215 = ~n26202 & ~n26214;
  assign n26216 = n3476 & ~n26215;
  assign n26217 = ~n26211 & ~n26216;
  assign n26218 = n3374 & ~n26217;
  assign n26219 = ~n26206 & ~n26218;
  assign n26220 = n3655 & ~n26219;
  assign n26221 = n3492 & ~n25747;
  assign n26222 = ~n3631 & ~n26221;
  assign n26223 = n3485 & ~n26222;
  assign n26224 = ~n3630 & ~n26223;
  assign n26225 = ~n3476 & ~n26224;
  assign n26226 = ~n4946 & ~n26136;
  assign n26227 = i_hlock3 & ~n26226;
  assign n26228 = ~n4946 & ~n26140;
  assign n26229 = ~i_hlock3 & ~n26228;
  assign n26230 = ~n26227 & ~n26229;
  assign n26231 = i_hbusreq3 & ~n26230;
  assign n26232 = ~n5009 & ~n26146;
  assign n26233 = i_hlock3 & ~n26232;
  assign n26234 = ~n5009 & ~n26150;
  assign n26235 = ~i_hlock3 & ~n26234;
  assign n26236 = ~n26233 & ~n26235;
  assign n26237 = ~i_hbusreq3 & ~n26236;
  assign n26238 = ~n26231 & ~n26237;
  assign n26239 = ~controllable_hmaster2 & ~n26238;
  assign n26240 = ~n3407 & ~n26239;
  assign n26241 = controllable_hgrant3 & ~n26240;
  assign n26242 = ~n6151 & ~n11402;
  assign n26243 = i_hlock3 & ~n26242;
  assign n26244 = ~n6151 & ~n11406;
  assign n26245 = ~i_hlock3 & ~n26244;
  assign n26246 = ~n26243 & ~n26245;
  assign n26247 = i_hbusreq3 & ~n26246;
  assign n26248 = ~n6180 & ~n11412;
  assign n26249 = i_hlock3 & ~n26248;
  assign n26250 = ~n6180 & ~n11416;
  assign n26251 = ~i_hlock3 & ~n26250;
  assign n26252 = ~n26249 & ~n26251;
  assign n26253 = ~i_hbusreq3 & ~n26252;
  assign n26254 = ~n26247 & ~n26253;
  assign n26255 = ~controllable_hmaster2 & ~n26254;
  assign n26256 = ~n3461 & ~n26255;
  assign n26257 = ~controllable_hgrant3 & ~n26256;
  assign n26258 = ~n26241 & ~n26257;
  assign n26259 = controllable_nhgrant0 & ~n26258;
  assign n26260 = ~n4946 & ~n11402;
  assign n26261 = i_hlock3 & ~n26260;
  assign n26262 = ~n4946 & ~n11406;
  assign n26263 = ~i_hlock3 & ~n26262;
  assign n26264 = ~n26261 & ~n26263;
  assign n26265 = i_hbusreq3 & ~n26264;
  assign n26266 = ~n5009 & ~n11412;
  assign n26267 = i_hlock3 & ~n26266;
  assign n26268 = ~n5009 & ~n11416;
  assign n26269 = ~i_hlock3 & ~n26268;
  assign n26270 = ~n26267 & ~n26269;
  assign n26271 = ~i_hbusreq3 & ~n26270;
  assign n26272 = ~n26265 & ~n26271;
  assign n26273 = ~controllable_hmaster2 & ~n26272;
  assign n26274 = ~n3407 & ~n26273;
  assign n26275 = controllable_hgrant3 & ~n26274;
  assign n26276 = ~n5225 & ~n11402;
  assign n26277 = i_hlock3 & ~n26276;
  assign n26278 = ~n5225 & ~n11406;
  assign n26279 = ~i_hlock3 & ~n26278;
  assign n26280 = ~n26277 & ~n26279;
  assign n26281 = i_hbusreq3 & ~n26280;
  assign n26282 = ~n5233 & ~n11412;
  assign n26283 = i_hlock3 & ~n26282;
  assign n26284 = ~n5233 & ~n11416;
  assign n26285 = ~i_hlock3 & ~n26284;
  assign n26286 = ~n26283 & ~n26285;
  assign n26287 = ~i_hbusreq3 & ~n26286;
  assign n26288 = ~n26281 & ~n26287;
  assign n26289 = ~controllable_hmaster2 & ~n26288;
  assign n26290 = ~n3407 & ~n26289;
  assign n26291 = ~controllable_hgrant3 & ~n26290;
  assign n26292 = ~n26275 & ~n26291;
  assign n26293 = ~controllable_nhgrant0 & ~n26292;
  assign n26294 = ~n26259 & ~n26293;
  assign n26295 = ~n3281 & ~n26294;
  assign n26296 = ~n3783 & ~n26295;
  assign n26297 = ~n3492 & ~n26296;
  assign n26298 = ~n8310 & ~n26297;
  assign n26299 = ~n3485 & ~n26298;
  assign n26300 = ~n26223 & ~n26299;
  assign n26301 = n3476 & ~n26300;
  assign n26302 = ~n26225 & ~n26301;
  assign n26303 = ~n3374 & ~n26302;
  assign n26304 = n3492 & ~n25765;
  assign n26305 = ~n3631 & ~n26304;
  assign n26306 = n3485 & ~n26305;
  assign n26307 = ~n3630 & ~n26306;
  assign n26308 = ~n3476 & ~n26307;
  assign n26309 = n3492 & ~n25783;
  assign n26310 = ~n3631 & ~n26309;
  assign n26311 = n3485 & ~n26310;
  assign n26312 = ~n26299 & ~n26311;
  assign n26313 = n3476 & ~n26312;
  assign n26314 = ~n26308 & ~n26313;
  assign n26315 = n3374 & ~n26314;
  assign n26316 = ~n26303 & ~n26315;
  assign n26317 = ~n3655 & ~n26316;
  assign n26318 = ~n26220 & ~n26317;
  assign n26319 = n3652 & ~n26318;
  assign n26320 = n3492 & ~n25801;
  assign n26321 = ~n3631 & ~n26320;
  assign n26322 = n3485 & ~n26321;
  assign n26323 = ~n3630 & ~n26322;
  assign n26324 = ~n3476 & ~n26323;
  assign n26325 = ~n8289 & ~n25612;
  assign n26326 = i_hlock3 & ~n26325;
  assign n26327 = ~n8289 & ~n25619;
  assign n26328 = ~i_hlock3 & ~n26327;
  assign n26329 = ~n26326 & ~n26328;
  assign n26330 = i_hbusreq3 & ~n26329;
  assign n26331 = ~n8289 & ~n25631;
  assign n26332 = i_hlock3 & ~n26331;
  assign n26333 = ~n8289 & ~n25641;
  assign n26334 = ~i_hlock3 & ~n26333;
  assign n26335 = ~n26332 & ~n26334;
  assign n26336 = ~i_hbusreq3 & ~n26335;
  assign n26337 = ~n26330 & ~n26336;
  assign n26338 = ~controllable_hmaster2 & ~n26337;
  assign n26339 = ~n3407 & ~n26338;
  assign n26340 = controllable_hgrant3 & ~n26339;
  assign n26341 = ~n6602 & ~n8289;
  assign n26342 = i_hlock3 & ~n26341;
  assign n26343 = ~n6606 & ~n8289;
  assign n26344 = ~i_hlock3 & ~n26343;
  assign n26345 = ~n26342 & ~n26344;
  assign n26346 = i_hbusreq3 & ~n26345;
  assign n26347 = ~n6647 & ~n8289;
  assign n26348 = i_hlock3 & ~n26347;
  assign n26349 = ~n6651 & ~n8289;
  assign n26350 = ~i_hlock3 & ~n26349;
  assign n26351 = ~n26348 & ~n26350;
  assign n26352 = ~i_hbusreq3 & ~n26351;
  assign n26353 = ~n26346 & ~n26352;
  assign n26354 = ~controllable_hmaster2 & ~n26353;
  assign n26355 = ~n3461 & ~n26354;
  assign n26356 = ~controllable_hgrant3 & ~n26355;
  assign n26357 = ~n26340 & ~n26356;
  assign n26358 = controllable_nhgrant0 & ~n26357;
  assign n26359 = ~n5167 & ~n8289;
  assign n26360 = i_hlock3 & ~n26359;
  assign n26361 = ~n5171 & ~n8289;
  assign n26362 = ~i_hlock3 & ~n26361;
  assign n26363 = ~n26360 & ~n26362;
  assign n26364 = i_hbusreq3 & ~n26363;
  assign n26365 = ~n5177 & ~n8289;
  assign n26366 = i_hlock3 & ~n26365;
  assign n26367 = ~n5181 & ~n8289;
  assign n26368 = ~i_hlock3 & ~n26367;
  assign n26369 = ~n26366 & ~n26368;
  assign n26370 = ~i_hbusreq3 & ~n26369;
  assign n26371 = ~n26364 & ~n26370;
  assign n26372 = ~controllable_hmaster2 & ~n26371;
  assign n26373 = ~n3407 & ~n26372;
  assign n26374 = controllable_hgrant3 & ~n26373;
  assign n26375 = ~n5167 & ~n8299;
  assign n26376 = i_hlock3 & ~n26375;
  assign n26377 = ~n5171 & ~n8299;
  assign n26378 = ~i_hlock3 & ~n26377;
  assign n26379 = ~n26376 & ~n26378;
  assign n26380 = i_hbusreq3 & ~n26379;
  assign n26381 = ~n5177 & ~n8299;
  assign n26382 = i_hlock3 & ~n26381;
  assign n26383 = ~n5181 & ~n8299;
  assign n26384 = ~i_hlock3 & ~n26383;
  assign n26385 = ~n26382 & ~n26384;
  assign n26386 = ~i_hbusreq3 & ~n26385;
  assign n26387 = ~n26380 & ~n26386;
  assign n26388 = ~controllable_hmaster2 & ~n26387;
  assign n26389 = ~n3407 & ~n26388;
  assign n26390 = ~controllable_hgrant3 & ~n26389;
  assign n26391 = ~n26374 & ~n26390;
  assign n26392 = ~controllable_nhgrant0 & ~n26391;
  assign n26393 = ~n26358 & ~n26392;
  assign n26394 = ~n3281 & ~n26393;
  assign n26395 = ~n3783 & ~n26394;
  assign n26396 = ~n3492 & ~n26395;
  assign n26397 = ~n8310 & ~n26396;
  assign n26398 = ~n3485 & ~n26397;
  assign n26399 = ~n26322 & ~n26398;
  assign n26400 = n3476 & ~n26399;
  assign n26401 = ~n26324 & ~n26400;
  assign n26402 = ~n3374 & ~n26401;
  assign n26403 = n3492 & ~n25819;
  assign n26404 = ~n3631 & ~n26403;
  assign n26405 = n3485 & ~n26404;
  assign n26406 = ~n3630 & ~n26405;
  assign n26407 = ~n3476 & ~n26406;
  assign n26408 = n3492 & ~n25837;
  assign n26409 = ~n3631 & ~n26408;
  assign n26410 = n3485 & ~n26409;
  assign n26411 = ~n26398 & ~n26410;
  assign n26412 = n3476 & ~n26411;
  assign n26413 = ~n26407 & ~n26412;
  assign n26414 = n3374 & ~n26413;
  assign n26415 = ~n26402 & ~n26414;
  assign n26416 = n3655 & ~n26415;
  assign n26417 = n3492 & ~n25853;
  assign n26418 = ~n3631 & ~n26417;
  assign n26419 = n3485 & ~n26418;
  assign n26420 = ~n3630 & ~n26419;
  assign n26421 = ~n3476 & ~n26420;
  assign n26422 = ~n3407 & ~n25647;
  assign n26423 = controllable_hgrant3 & ~n26422;
  assign n26424 = ~n3461 & ~n6887;
  assign n26425 = ~controllable_hgrant3 & ~n26424;
  assign n26426 = ~n26423 & ~n26425;
  assign n26427 = controllable_nhgrant0 & ~n26426;
  assign n26428 = ~n3407 & ~n5187;
  assign n26429 = controllable_hgrant3 & ~n26428;
  assign n26430 = ~n3407 & ~n5241;
  assign n26431 = ~controllable_hgrant3 & ~n26430;
  assign n26432 = ~n26429 & ~n26431;
  assign n26433 = ~controllable_nhgrant0 & ~n26432;
  assign n26434 = ~n26427 & ~n26433;
  assign n26435 = ~n3281 & ~n26434;
  assign n26436 = ~n3783 & ~n26435;
  assign n26437 = ~n3492 & ~n26436;
  assign n26438 = ~n8310 & ~n26437;
  assign n26439 = ~n3485 & ~n26438;
  assign n26440 = ~n26419 & ~n26439;
  assign n26441 = n3476 & ~n26440;
  assign n26442 = ~n26421 & ~n26441;
  assign n26443 = ~n3374 & ~n26442;
  assign n26444 = n3492 & ~n25871;
  assign n26445 = ~n3631 & ~n26444;
  assign n26446 = n3485 & ~n26445;
  assign n26447 = ~n3630 & ~n26446;
  assign n26448 = ~n3476 & ~n26447;
  assign n26449 = n3492 & ~n25889;
  assign n26450 = ~n3631 & ~n26449;
  assign n26451 = n3485 & ~n26450;
  assign n26452 = ~n26439 & ~n26451;
  assign n26453 = n3476 & ~n26452;
  assign n26454 = ~n26448 & ~n26453;
  assign n26455 = n3374 & ~n26454;
  assign n26456 = ~n26443 & ~n26455;
  assign n26457 = ~n3655 & ~n26456;
  assign n26458 = ~n26416 & ~n26457;
  assign n26459 = ~n3652 & ~n26458;
  assign n26460 = ~n26319 & ~n26459;
  assign n26461 = ~n3368 & ~n26460;
  assign n26462 = n3492 & ~n25910;
  assign n26463 = n3492 & ~n26462;
  assign n26464 = n3485 & ~n26463;
  assign n26465 = n3485 & ~n26464;
  assign n26466 = ~n3476 & ~n26465;
  assign n26467 = ~n8525 & ~n26464;
  assign n26468 = n3476 & ~n26467;
  assign n26469 = ~n26466 & ~n26468;
  assign n26470 = ~n3374 & ~n26469;
  assign n26471 = n3492 & ~n25932;
  assign n26472 = n3492 & ~n26471;
  assign n26473 = n3485 & ~n26472;
  assign n26474 = n3485 & ~n26473;
  assign n26475 = ~n3476 & ~n26474;
  assign n26476 = ~n3281 & ~n26198;
  assign n26477 = ~n3492 & ~n26476;
  assign n26478 = ~n3492 & ~n26477;
  assign n26479 = ~n3485 & ~n26478;
  assign n26480 = n3492 & ~n25954;
  assign n26481 = n3492 & ~n26480;
  assign n26482 = n3485 & ~n26481;
  assign n26483 = ~n26479 & ~n26482;
  assign n26484 = n3476 & ~n26483;
  assign n26485 = ~n26475 & ~n26484;
  assign n26486 = n3374 & ~n26485;
  assign n26487 = ~n26470 & ~n26486;
  assign n26488 = n3655 & ~n26487;
  assign n26489 = n3492 & ~n25970;
  assign n26490 = n3492 & ~n26489;
  assign n26491 = n3485 & ~n26490;
  assign n26492 = n3485 & ~n26491;
  assign n26493 = ~n3476 & ~n26492;
  assign n26494 = ~n8525 & ~n26491;
  assign n26495 = n3476 & ~n26494;
  assign n26496 = ~n26493 & ~n26495;
  assign n26497 = ~n3374 & ~n26496;
  assign n26498 = n3492 & ~n25988;
  assign n26499 = n3492 & ~n26498;
  assign n26500 = n3485 & ~n26499;
  assign n26501 = n3485 & ~n26500;
  assign n26502 = ~n3476 & ~n26501;
  assign n26503 = ~n3281 & ~n26295;
  assign n26504 = ~n3492 & ~n26503;
  assign n26505 = ~n3492 & ~n26504;
  assign n26506 = ~n3485 & ~n26505;
  assign n26507 = n3492 & ~n26006;
  assign n26508 = n3492 & ~n26507;
  assign n26509 = n3485 & ~n26508;
  assign n26510 = ~n26506 & ~n26509;
  assign n26511 = n3476 & ~n26510;
  assign n26512 = ~n26502 & ~n26511;
  assign n26513 = n3374 & ~n26512;
  assign n26514 = ~n26497 & ~n26513;
  assign n26515 = ~n3655 & ~n26514;
  assign n26516 = ~n26488 & ~n26515;
  assign n26517 = n3652 & ~n26516;
  assign n26518 = n3492 & ~n26024;
  assign n26519 = n3492 & ~n26518;
  assign n26520 = n3485 & ~n26519;
  assign n26521 = n3485 & ~n26520;
  assign n26522 = ~n3476 & ~n26521;
  assign n26523 = ~n8525 & ~n26520;
  assign n26524 = n3476 & ~n26523;
  assign n26525 = ~n26522 & ~n26524;
  assign n26526 = ~n3374 & ~n26525;
  assign n26527 = n3492 & ~n26042;
  assign n26528 = n3492 & ~n26527;
  assign n26529 = n3485 & ~n26528;
  assign n26530 = n3485 & ~n26529;
  assign n26531 = ~n3476 & ~n26530;
  assign n26532 = ~n3281 & ~n26394;
  assign n26533 = ~n3492 & ~n26532;
  assign n26534 = ~n3492 & ~n26533;
  assign n26535 = ~n3485 & ~n26534;
  assign n26536 = n3492 & ~n26060;
  assign n26537 = n3492 & ~n26536;
  assign n26538 = n3485 & ~n26537;
  assign n26539 = ~n26535 & ~n26538;
  assign n26540 = n3476 & ~n26539;
  assign n26541 = ~n26531 & ~n26540;
  assign n26542 = n3374 & ~n26541;
  assign n26543 = ~n26526 & ~n26542;
  assign n26544 = n3655 & ~n26543;
  assign n26545 = n3492 & ~n26076;
  assign n26546 = n3492 & ~n26545;
  assign n26547 = n3485 & ~n26546;
  assign n26548 = n3485 & ~n26547;
  assign n26549 = ~n3476 & ~n26548;
  assign n26550 = ~n8525 & ~n26547;
  assign n26551 = n3476 & ~n26550;
  assign n26552 = ~n26549 & ~n26551;
  assign n26553 = ~n3374 & ~n26552;
  assign n26554 = n3492 & ~n26094;
  assign n26555 = n3492 & ~n26554;
  assign n26556 = n3485 & ~n26555;
  assign n26557 = n3485 & ~n26556;
  assign n26558 = ~n3476 & ~n26557;
  assign n26559 = ~n3281 & ~n26435;
  assign n26560 = ~n3492 & ~n26559;
  assign n26561 = ~n3492 & ~n26560;
  assign n26562 = ~n3485 & ~n26561;
  assign n26563 = n3492 & ~n26112;
  assign n26564 = n3492 & ~n26563;
  assign n26565 = n3485 & ~n26564;
  assign n26566 = ~n26562 & ~n26565;
  assign n26567 = n3476 & ~n26566;
  assign n26568 = ~n26558 & ~n26567;
  assign n26569 = n3374 & ~n26568;
  assign n26570 = ~n26553 & ~n26569;
  assign n26571 = ~n3655 & ~n26570;
  assign n26572 = ~n26544 & ~n26571;
  assign n26573 = ~n3652 & ~n26572;
  assign n26574 = ~n26517 & ~n26573;
  assign n26575 = n3368 & ~n26574;
  assign n26576 = ~n26461 & ~n26575;
  assign n26577 = ~n3362 & ~n26576;
  assign n26578 = ~n26129 & ~n26577;
  assign n26579 = n3359 & ~n26578;
  assign n26580 = ~n3485 & ~n26199;
  assign n26581 = ~n26132 & ~n26580;
  assign n26582 = n3476 & ~n26581;
  assign n26583 = ~n26134 & ~n26582;
  assign n26584 = ~n3374 & ~n26583;
  assign n26585 = ~n26214 & ~n26580;
  assign n26586 = n3476 & ~n26585;
  assign n26587 = ~n26211 & ~n26586;
  assign n26588 = n3374 & ~n26587;
  assign n26589 = ~n26584 & ~n26588;
  assign n26590 = n3655 & ~n26589;
  assign n26591 = ~n3485 & ~n26296;
  assign n26592 = ~n26223 & ~n26591;
  assign n26593 = n3476 & ~n26592;
  assign n26594 = ~n26225 & ~n26593;
  assign n26595 = ~n3374 & ~n26594;
  assign n26596 = ~n26311 & ~n26591;
  assign n26597 = n3476 & ~n26596;
  assign n26598 = ~n26308 & ~n26597;
  assign n26599 = n3374 & ~n26598;
  assign n26600 = ~n26595 & ~n26599;
  assign n26601 = ~n3655 & ~n26600;
  assign n26602 = ~n26590 & ~n26601;
  assign n26603 = n3652 & ~n26602;
  assign n26604 = ~n3485 & ~n26395;
  assign n26605 = ~n26322 & ~n26604;
  assign n26606 = n3476 & ~n26605;
  assign n26607 = ~n26324 & ~n26606;
  assign n26608 = ~n3374 & ~n26607;
  assign n26609 = ~n26410 & ~n26604;
  assign n26610 = n3476 & ~n26609;
  assign n26611 = ~n26407 & ~n26610;
  assign n26612 = n3374 & ~n26611;
  assign n26613 = ~n26608 & ~n26612;
  assign n26614 = n3655 & ~n26613;
  assign n26615 = ~n3485 & ~n26436;
  assign n26616 = ~n26419 & ~n26615;
  assign n26617 = n3476 & ~n26616;
  assign n26618 = ~n26421 & ~n26617;
  assign n26619 = ~n3374 & ~n26618;
  assign n26620 = ~n26451 & ~n26615;
  assign n26621 = n3476 & ~n26620;
  assign n26622 = ~n26448 & ~n26621;
  assign n26623 = n3374 & ~n26622;
  assign n26624 = ~n26619 & ~n26623;
  assign n26625 = ~n3655 & ~n26624;
  assign n26626 = ~n26614 & ~n26625;
  assign n26627 = ~n3652 & ~n26626;
  assign n26628 = ~n26603 & ~n26627;
  assign n26629 = ~n3368 & ~n26628;
  assign n26630 = ~n8689 & ~n26464;
  assign n26631 = n3476 & ~n26630;
  assign n26632 = ~n26466 & ~n26631;
  assign n26633 = ~n3374 & ~n26632;
  assign n26634 = ~n3485 & ~n26476;
  assign n26635 = ~n26482 & ~n26634;
  assign n26636 = n3476 & ~n26635;
  assign n26637 = ~n26475 & ~n26636;
  assign n26638 = n3374 & ~n26637;
  assign n26639 = ~n26633 & ~n26638;
  assign n26640 = n3655 & ~n26639;
  assign n26641 = ~n8689 & ~n26491;
  assign n26642 = n3476 & ~n26641;
  assign n26643 = ~n26493 & ~n26642;
  assign n26644 = ~n3374 & ~n26643;
  assign n26645 = ~n3485 & ~n26503;
  assign n26646 = ~n26509 & ~n26645;
  assign n26647 = n3476 & ~n26646;
  assign n26648 = ~n26502 & ~n26647;
  assign n26649 = n3374 & ~n26648;
  assign n26650 = ~n26644 & ~n26649;
  assign n26651 = ~n3655 & ~n26650;
  assign n26652 = ~n26640 & ~n26651;
  assign n26653 = n3652 & ~n26652;
  assign n26654 = ~n8689 & ~n26520;
  assign n26655 = n3476 & ~n26654;
  assign n26656 = ~n26522 & ~n26655;
  assign n26657 = ~n3374 & ~n26656;
  assign n26658 = ~n3485 & ~n26532;
  assign n26659 = ~n26538 & ~n26658;
  assign n26660 = n3476 & ~n26659;
  assign n26661 = ~n26531 & ~n26660;
  assign n26662 = n3374 & ~n26661;
  assign n26663 = ~n26657 & ~n26662;
  assign n26664 = n3655 & ~n26663;
  assign n26665 = ~n8689 & ~n26547;
  assign n26666 = n3476 & ~n26665;
  assign n26667 = ~n26549 & ~n26666;
  assign n26668 = ~n3374 & ~n26667;
  assign n26669 = ~n3485 & ~n26559;
  assign n26670 = ~n26565 & ~n26669;
  assign n26671 = n3476 & ~n26670;
  assign n26672 = ~n26558 & ~n26671;
  assign n26673 = n3374 & ~n26672;
  assign n26674 = ~n26668 & ~n26673;
  assign n26675 = ~n3655 & ~n26674;
  assign n26676 = ~n26664 & ~n26675;
  assign n26677 = ~n3652 & ~n26676;
  assign n26678 = ~n26653 & ~n26677;
  assign n26679 = n3368 & ~n26678;
  assign n26680 = ~n26629 & ~n26679;
  assign n26681 = n3362 & ~n26680;
  assign n26682 = n3378 & ~n25654;
  assign n26683 = ~n8781 & ~n25647;
  assign n26684 = controllable_hgrant3 & ~n26683;
  assign n26685 = ~n8762 & ~n26684;
  assign n26686 = controllable_nhgrant0 & ~n26685;
  assign n26687 = ~n8785 & ~n26686;
  assign n26688 = ~n3281 & ~n26687;
  assign n26689 = ~n3783 & ~n26688;
  assign n26690 = ~n3378 & ~n26689;
  assign n26691 = ~n26682 & ~n26690;
  assign n26692 = n3492 & ~n26691;
  assign n26693 = ~n3631 & ~n26692;
  assign n26694 = n3485 & ~n26693;
  assign n26695 = ~n3630 & ~n26694;
  assign n26696 = ~n3476 & ~n26695;
  assign n26697 = ~n26200 & ~n26692;
  assign n26698 = n3485 & ~n26697;
  assign n26699 = ~n26580 & ~n26698;
  assign n26700 = n3476 & ~n26699;
  assign n26701 = ~n26696 & ~n26700;
  assign n26702 = ~n3374 & ~n26701;
  assign n26703 = n3378 & ~n25689;
  assign n26704 = ~n8898 & ~n25682;
  assign n26705 = controllable_hgrant3 & ~n26704;
  assign n26706 = ~n8884 & ~n26705;
  assign n26707 = controllable_nhgrant0 & ~n26706;
  assign n26708 = ~n8902 & ~n26707;
  assign n26709 = ~n3281 & ~n26708;
  assign n26710 = ~n3950 & ~n26709;
  assign n26711 = ~n3378 & ~n26710;
  assign n26712 = ~n26703 & ~n26711;
  assign n26713 = n3492 & ~n26712;
  assign n26714 = ~n3631 & ~n26713;
  assign n26715 = n3485 & ~n26714;
  assign n26716 = ~n3630 & ~n26715;
  assign n26717 = ~n3476 & ~n26716;
  assign n26718 = n3378 & ~n25731;
  assign n26719 = ~n9092 & ~n25724;
  assign n26720 = controllable_hgrant3 & ~n26719;
  assign n26721 = ~n9052 & ~n26720;
  assign n26722 = controllable_nhgrant0 & ~n26721;
  assign n26723 = ~n9096 & ~n26722;
  assign n26724 = ~n3281 & ~n26723;
  assign n26725 = ~n4089 & ~n26724;
  assign n26726 = ~n3378 & ~n26725;
  assign n26727 = ~n26718 & ~n26726;
  assign n26728 = n3492 & ~n26727;
  assign n26729 = ~n26200 & ~n26728;
  assign n26730 = n3485 & ~n26729;
  assign n26731 = ~n26580 & ~n26730;
  assign n26732 = n3476 & ~n26731;
  assign n26733 = ~n26717 & ~n26732;
  assign n26734 = n3374 & ~n26733;
  assign n26735 = ~n26702 & ~n26734;
  assign n26736 = n3655 & ~n26735;
  assign n26737 = n3378 & ~n25747;
  assign n26738 = ~n9129 & ~n26684;
  assign n26739 = controllable_nhgrant0 & ~n26738;
  assign n26740 = ~n8785 & ~n26739;
  assign n26741 = ~n3281 & ~n26740;
  assign n26742 = ~n3783 & ~n26741;
  assign n26743 = ~n3378 & ~n26742;
  assign n26744 = ~n26737 & ~n26743;
  assign n26745 = n3492 & ~n26744;
  assign n26746 = ~n3631 & ~n26745;
  assign n26747 = n3485 & ~n26746;
  assign n26748 = ~n3630 & ~n26747;
  assign n26749 = ~n3476 & ~n26748;
  assign n26750 = ~n26297 & ~n26745;
  assign n26751 = n3485 & ~n26750;
  assign n26752 = ~n26591 & ~n26751;
  assign n26753 = n3476 & ~n26752;
  assign n26754 = ~n26749 & ~n26753;
  assign n26755 = ~n3374 & ~n26754;
  assign n26756 = n3378 & ~n25765;
  assign n26757 = ~n9234 & ~n26705;
  assign n26758 = controllable_nhgrant0 & ~n26757;
  assign n26759 = ~n8902 & ~n26758;
  assign n26760 = ~n3281 & ~n26759;
  assign n26761 = ~n3950 & ~n26760;
  assign n26762 = ~n3378 & ~n26761;
  assign n26763 = ~n26756 & ~n26762;
  assign n26764 = n3492 & ~n26763;
  assign n26765 = ~n3631 & ~n26764;
  assign n26766 = n3485 & ~n26765;
  assign n26767 = ~n3630 & ~n26766;
  assign n26768 = ~n3476 & ~n26767;
  assign n26769 = n3378 & ~n25783;
  assign n26770 = ~n9368 & ~n26720;
  assign n26771 = controllable_nhgrant0 & ~n26770;
  assign n26772 = ~n9096 & ~n26771;
  assign n26773 = ~n3281 & ~n26772;
  assign n26774 = ~n4089 & ~n26773;
  assign n26775 = ~n3378 & ~n26774;
  assign n26776 = ~n26769 & ~n26775;
  assign n26777 = n3492 & ~n26776;
  assign n26778 = ~n26297 & ~n26777;
  assign n26779 = n3485 & ~n26778;
  assign n26780 = ~n26591 & ~n26779;
  assign n26781 = n3476 & ~n26780;
  assign n26782 = ~n26768 & ~n26781;
  assign n26783 = n3374 & ~n26782;
  assign n26784 = ~n26755 & ~n26783;
  assign n26785 = ~n3655 & ~n26784;
  assign n26786 = ~n26736 & ~n26785;
  assign n26787 = n3652 & ~n26786;
  assign n26788 = n3378 & ~n25801;
  assign n26789 = ~n9403 & ~n26684;
  assign n26790 = controllable_nhgrant0 & ~n26789;
  assign n26791 = ~n8785 & ~n26790;
  assign n26792 = ~n3281 & ~n26791;
  assign n26793 = ~n3783 & ~n26792;
  assign n26794 = ~n3378 & ~n26793;
  assign n26795 = ~n26788 & ~n26794;
  assign n26796 = n3492 & ~n26795;
  assign n26797 = ~n3631 & ~n26796;
  assign n26798 = n3485 & ~n26797;
  assign n26799 = ~n3630 & ~n26798;
  assign n26800 = ~n3476 & ~n26799;
  assign n26801 = ~n26396 & ~n26796;
  assign n26802 = n3485 & ~n26801;
  assign n26803 = ~n26604 & ~n26802;
  assign n26804 = n3476 & ~n26803;
  assign n26805 = ~n26800 & ~n26804;
  assign n26806 = ~n3374 & ~n26805;
  assign n26807 = n3378 & ~n25819;
  assign n26808 = ~n9463 & ~n26705;
  assign n26809 = controllable_nhgrant0 & ~n26808;
  assign n26810 = ~n8902 & ~n26809;
  assign n26811 = ~n3281 & ~n26810;
  assign n26812 = ~n3950 & ~n26811;
  assign n26813 = ~n3378 & ~n26812;
  assign n26814 = ~n26807 & ~n26813;
  assign n26815 = n3492 & ~n26814;
  assign n26816 = ~n3631 & ~n26815;
  assign n26817 = n3485 & ~n26816;
  assign n26818 = ~n3630 & ~n26817;
  assign n26819 = ~n3476 & ~n26818;
  assign n26820 = n3378 & ~n25837;
  assign n26821 = ~n9525 & ~n26720;
  assign n26822 = controllable_nhgrant0 & ~n26821;
  assign n26823 = ~n9096 & ~n26822;
  assign n26824 = ~n3281 & ~n26823;
  assign n26825 = ~n4089 & ~n26824;
  assign n26826 = ~n3378 & ~n26825;
  assign n26827 = ~n26820 & ~n26826;
  assign n26828 = n3492 & ~n26827;
  assign n26829 = ~n26396 & ~n26828;
  assign n26830 = n3485 & ~n26829;
  assign n26831 = ~n26604 & ~n26830;
  assign n26832 = n3476 & ~n26831;
  assign n26833 = ~n26819 & ~n26832;
  assign n26834 = n3374 & ~n26833;
  assign n26835 = ~n26806 & ~n26834;
  assign n26836 = n3655 & ~n26835;
  assign n26837 = n3378 & ~n25853;
  assign n26838 = ~n9557 & ~n26684;
  assign n26839 = controllable_nhgrant0 & ~n26838;
  assign n26840 = ~n8785 & ~n26839;
  assign n26841 = ~n3281 & ~n26840;
  assign n26842 = ~n3783 & ~n26841;
  assign n26843 = ~n3378 & ~n26842;
  assign n26844 = ~n26837 & ~n26843;
  assign n26845 = n3492 & ~n26844;
  assign n26846 = ~n3631 & ~n26845;
  assign n26847 = n3485 & ~n26846;
  assign n26848 = ~n3630 & ~n26847;
  assign n26849 = ~n3476 & ~n26848;
  assign n26850 = ~n26437 & ~n26845;
  assign n26851 = n3485 & ~n26850;
  assign n26852 = ~n26615 & ~n26851;
  assign n26853 = n3476 & ~n26852;
  assign n26854 = ~n26849 & ~n26853;
  assign n26855 = ~n3374 & ~n26854;
  assign n26856 = n3378 & ~n25871;
  assign n26857 = ~n9617 & ~n26705;
  assign n26858 = controllable_nhgrant0 & ~n26857;
  assign n26859 = ~n8902 & ~n26858;
  assign n26860 = ~n3281 & ~n26859;
  assign n26861 = ~n3950 & ~n26860;
  assign n26862 = ~n3378 & ~n26861;
  assign n26863 = ~n26856 & ~n26862;
  assign n26864 = n3492 & ~n26863;
  assign n26865 = ~n3631 & ~n26864;
  assign n26866 = n3485 & ~n26865;
  assign n26867 = ~n3630 & ~n26866;
  assign n26868 = ~n3476 & ~n26867;
  assign n26869 = n3378 & ~n25889;
  assign n26870 = ~n9677 & ~n26720;
  assign n26871 = controllable_nhgrant0 & ~n26870;
  assign n26872 = ~n9096 & ~n26871;
  assign n26873 = ~n3281 & ~n26872;
  assign n26874 = ~n4089 & ~n26873;
  assign n26875 = ~n3378 & ~n26874;
  assign n26876 = ~n26869 & ~n26875;
  assign n26877 = n3492 & ~n26876;
  assign n26878 = ~n26437 & ~n26877;
  assign n26879 = n3485 & ~n26878;
  assign n26880 = ~n26615 & ~n26879;
  assign n26881 = n3476 & ~n26880;
  assign n26882 = ~n26868 & ~n26881;
  assign n26883 = n3374 & ~n26882;
  assign n26884 = ~n26855 & ~n26883;
  assign n26885 = ~n3655 & ~n26884;
  assign n26886 = ~n26836 & ~n26885;
  assign n26887 = ~n3652 & ~n26886;
  assign n26888 = ~n26787 & ~n26887;
  assign n26889 = ~n3368 & ~n26888;
  assign n26890 = n3378 & ~n25910;
  assign n26891 = controllable_hgrant3 & ~n9750;
  assign n26892 = ~n9733 & ~n26891;
  assign n26893 = controllable_nhgrant0 & ~n26892;
  assign n26894 = ~n9753 & ~n26893;
  assign n26895 = ~n3281 & ~n26894;
  assign n26896 = ~n3281 & ~n26895;
  assign n26897 = ~n3378 & ~n26896;
  assign n26898 = ~n26890 & ~n26897;
  assign n26899 = n3492 & ~n26898;
  assign n26900 = n3492 & ~n26899;
  assign n26901 = n3485 & ~n26900;
  assign n26902 = n3485 & ~n26901;
  assign n26903 = ~n3476 & ~n26902;
  assign n26904 = ~n8523 & ~n26899;
  assign n26905 = n3485 & ~n26904;
  assign n26906 = ~n8689 & ~n26905;
  assign n26907 = n3476 & ~n26906;
  assign n26908 = ~n26903 & ~n26907;
  assign n26909 = ~n3374 & ~n26908;
  assign n26910 = n3378 & ~n25932;
  assign n26911 = ~n3502 & ~n4611;
  assign n26912 = controllable_hmaster1 & ~n26911;
  assign n26913 = ~controllable_hmaster1 & ~n4610;
  assign n26914 = ~n26912 & ~n26913;
  assign n26915 = i_hbusreq3 & ~n26914;
  assign n26916 = ~n4636 & ~n9725;
  assign n26917 = controllable_hmaster1 & ~n26916;
  assign n26918 = ~n4611 & ~n9743;
  assign n26919 = ~controllable_hmaster1 & ~n26918;
  assign n26920 = ~n26917 & ~n26919;
  assign n26921 = ~i_hbusreq3 & ~n26920;
  assign n26922 = ~n26915 & ~n26921;
  assign n26923 = ~controllable_hmaster2 & ~n26922;
  assign n26924 = ~n9846 & ~n26923;
  assign n26925 = controllable_hgrant3 & ~n26924;
  assign n26926 = ~n9834 & ~n26925;
  assign n26927 = controllable_nhgrant0 & ~n26926;
  assign n26928 = ~n9861 & ~n26927;
  assign n26929 = ~n3281 & ~n26928;
  assign n26930 = ~n3281 & ~n26929;
  assign n26931 = ~n3378 & ~n26930;
  assign n26932 = ~n26910 & ~n26931;
  assign n26933 = n3492 & ~n26932;
  assign n26934 = n3492 & ~n26933;
  assign n26935 = n3485 & ~n26934;
  assign n26936 = n3485 & ~n26935;
  assign n26937 = ~n3476 & ~n26936;
  assign n26938 = ~controllable_hgrant2 & ~n10810;
  assign n26939 = ~n3410 & ~n26938;
  assign n26940 = controllable_hmaster1 & ~n26939;
  assign n26941 = controllable_hmaster0 & ~n26939;
  assign n26942 = ~controllable_hgrant2 & ~n10821;
  assign n26943 = ~n3410 & ~n26942;
  assign n26944 = ~controllable_hmaster0 & ~n26943;
  assign n26945 = ~n26941 & ~n26944;
  assign n26946 = ~controllable_hmaster1 & ~n26945;
  assign n26947 = ~n26940 & ~n26946;
  assign n26948 = i_hlock3 & ~n26947;
  assign n26949 = ~controllable_hgrant2 & ~n10813;
  assign n26950 = ~n3410 & ~n26949;
  assign n26951 = controllable_hmaster1 & ~n26950;
  assign n26952 = controllable_hmaster0 & ~n26950;
  assign n26953 = ~controllable_hgrant2 & ~n10824;
  assign n26954 = ~n3410 & ~n26953;
  assign n26955 = ~controllable_hmaster0 & ~n26954;
  assign n26956 = ~n26952 & ~n26955;
  assign n26957 = ~controllable_hmaster1 & ~n26956;
  assign n26958 = ~n26951 & ~n26957;
  assign n26959 = ~i_hlock3 & ~n26958;
  assign n26960 = ~n26948 & ~n26959;
  assign n26961 = i_hbusreq3 & ~n26960;
  assign n26962 = i_hbusreq2 & ~n10810;
  assign n26963 = ~i_hbusreq2 & ~n10851;
  assign n26964 = ~n26962 & ~n26963;
  assign n26965 = ~controllable_hgrant2 & ~n26964;
  assign n26966 = ~n3859 & ~n26965;
  assign n26967 = controllable_hmaster1 & ~n26966;
  assign n26968 = controllable_hmaster0 & ~n26966;
  assign n26969 = i_hbusreq2 & ~n10821;
  assign n26970 = ~i_hbusreq2 & ~n10887;
  assign n26971 = ~n26969 & ~n26970;
  assign n26972 = ~controllable_hgrant2 & ~n26971;
  assign n26973 = ~n4562 & ~n26972;
  assign n26974 = ~controllable_hmaster0 & ~n26973;
  assign n26975 = ~n26968 & ~n26974;
  assign n26976 = ~controllable_hmaster1 & ~n26975;
  assign n26977 = ~n26967 & ~n26976;
  assign n26978 = i_hlock3 & ~n26977;
  assign n26979 = i_hbusreq2 & ~n10813;
  assign n26980 = ~i_hbusreq2 & ~n10865;
  assign n26981 = ~n26979 & ~n26980;
  assign n26982 = ~controllable_hgrant2 & ~n26981;
  assign n26983 = ~n3859 & ~n26982;
  assign n26984 = controllable_hmaster1 & ~n26983;
  assign n26985 = controllable_hmaster0 & ~n26983;
  assign n26986 = i_hbusreq2 & ~n10824;
  assign n26987 = ~i_hbusreq2 & ~n10899;
  assign n26988 = ~n26986 & ~n26987;
  assign n26989 = ~controllable_hgrant2 & ~n26988;
  assign n26990 = ~n4562 & ~n26989;
  assign n26991 = ~controllable_hmaster0 & ~n26990;
  assign n26992 = ~n26985 & ~n26991;
  assign n26993 = ~controllable_hmaster1 & ~n26992;
  assign n26994 = ~n26984 & ~n26993;
  assign n26995 = ~i_hlock3 & ~n26994;
  assign n26996 = ~n26978 & ~n26995;
  assign n26997 = ~i_hbusreq3 & ~n26996;
  assign n26998 = ~n26961 & ~n26997;
  assign n26999 = controllable_hmaster2 & ~n26998;
  assign n27000 = ~controllable_hgrant2 & ~n10916;
  assign n27001 = ~n3410 & ~n27000;
  assign n27002 = controllable_hmaster0 & ~n27001;
  assign n27003 = ~controllable_hmaster0 & ~n26939;
  assign n27004 = ~n27002 & ~n27003;
  assign n27005 = controllable_hmaster1 & ~n27004;
  assign n27006 = ~controllable_hmaster1 & ~n26939;
  assign n27007 = ~n27005 & ~n27006;
  assign n27008 = i_hlock3 & ~n27007;
  assign n27009 = ~controllable_hgrant2 & ~n10919;
  assign n27010 = ~n3410 & ~n27009;
  assign n27011 = controllable_hmaster0 & ~n27010;
  assign n27012 = ~controllable_hmaster0 & ~n26950;
  assign n27013 = ~n27011 & ~n27012;
  assign n27014 = controllable_hmaster1 & ~n27013;
  assign n27015 = ~controllable_hmaster1 & ~n26950;
  assign n27016 = ~n27014 & ~n27015;
  assign n27017 = ~i_hlock3 & ~n27016;
  assign n27018 = ~n27008 & ~n27017;
  assign n27019 = i_hbusreq3 & ~n27018;
  assign n27020 = i_hbusreq2 & ~n10916;
  assign n27021 = ~i_hbusreq2 & ~n10953;
  assign n27022 = ~n27020 & ~n27021;
  assign n27023 = ~controllable_hgrant2 & ~n27022;
  assign n27024 = ~n3859 & ~n27023;
  assign n27025 = controllable_hmaster0 & ~n27024;
  assign n27026 = ~controllable_hmaster0 & ~n26966;
  assign n27027 = ~n27025 & ~n27026;
  assign n27028 = controllable_hmaster1 & ~n27027;
  assign n27029 = ~i_hbusreq2 & ~n10987;
  assign n27030 = ~n26962 & ~n27029;
  assign n27031 = ~controllable_hgrant2 & ~n27030;
  assign n27032 = ~n5461 & ~n27031;
  assign n27033 = ~controllable_hmaster0 & ~n27032;
  assign n27034 = ~n26968 & ~n27033;
  assign n27035 = ~controllable_hmaster1 & ~n27034;
  assign n27036 = ~n27028 & ~n27035;
  assign n27037 = i_hlock3 & ~n27036;
  assign n27038 = i_hbusreq2 & ~n10919;
  assign n27039 = ~i_hbusreq2 & ~n10967;
  assign n27040 = ~n27038 & ~n27039;
  assign n27041 = ~controllable_hgrant2 & ~n27040;
  assign n27042 = ~n3859 & ~n27041;
  assign n27043 = controllable_hmaster0 & ~n27042;
  assign n27044 = ~controllable_hmaster0 & ~n26983;
  assign n27045 = ~n27043 & ~n27044;
  assign n27046 = controllable_hmaster1 & ~n27045;
  assign n27047 = ~i_hbusreq2 & ~n10997;
  assign n27048 = ~n26979 & ~n27047;
  assign n27049 = ~controllable_hgrant2 & ~n27048;
  assign n27050 = ~n5461 & ~n27049;
  assign n27051 = ~controllable_hmaster0 & ~n27050;
  assign n27052 = ~n26985 & ~n27051;
  assign n27053 = ~controllable_hmaster1 & ~n27052;
  assign n27054 = ~n27046 & ~n27053;
  assign n27055 = ~i_hlock3 & ~n27054;
  assign n27056 = ~n27037 & ~n27055;
  assign n27057 = ~i_hbusreq3 & ~n27056;
  assign n27058 = ~n27019 & ~n27057;
  assign n27059 = ~controllable_hmaster2 & ~n27058;
  assign n27060 = ~n26999 & ~n27059;
  assign n27061 = controllable_hgrant3 & ~n27060;
  assign n27062 = ~n9952 & ~n27061;
  assign n27063 = controllable_nhgrant0 & ~n27062;
  assign n27064 = ~n10071 & ~n27063;
  assign n27065 = ~n3281 & ~n27064;
  assign n27066 = ~n3281 & ~n27065;
  assign n27067 = n3378 & ~n27066;
  assign n27068 = i_hlock3 & ~n26943;
  assign n27069 = ~i_hlock3 & ~n26954;
  assign n27070 = ~n27068 & ~n27069;
  assign n27071 = i_hbusreq3 & ~n27070;
  assign n27072 = ~i_hbusreq2 & ~n11034;
  assign n27073 = ~n26969 & ~n27072;
  assign n27074 = ~controllable_hgrant2 & ~n27073;
  assign n27075 = ~n4562 & ~n27074;
  assign n27076 = i_hlock3 & ~n27075;
  assign n27077 = ~i_hbusreq2 & ~n11044;
  assign n27078 = ~n26986 & ~n27077;
  assign n27079 = ~controllable_hgrant2 & ~n27078;
  assign n27080 = ~n4562 & ~n27079;
  assign n27081 = ~i_hlock3 & ~n27080;
  assign n27082 = ~n27076 & ~n27081;
  assign n27083 = ~i_hbusreq3 & ~n27082;
  assign n27084 = ~n27071 & ~n27083;
  assign n27085 = controllable_hmaster2 & ~n27084;
  assign n27086 = ~n3550 & ~n26944;
  assign n27087 = controllable_hmaster1 & ~n27086;
  assign n27088 = ~controllable_hmaster1 & ~n26943;
  assign n27089 = ~n27087 & ~n27088;
  assign n27090 = i_hlock3 & ~n27089;
  assign n27091 = ~controllable_hgrant2 & ~n11063;
  assign n27092 = ~n3410 & ~n27091;
  assign n27093 = controllable_hmaster0 & ~n27092;
  assign n27094 = ~n26955 & ~n27093;
  assign n27095 = controllable_hmaster1 & ~n27094;
  assign n27096 = ~controllable_hmaster1 & ~n26954;
  assign n27097 = ~n27095 & ~n27096;
  assign n27098 = ~i_hlock3 & ~n27097;
  assign n27099 = ~n27090 & ~n27098;
  assign n27100 = i_hbusreq3 & ~n27099;
  assign n27101 = ~i_hbusreq2 & ~n11091;
  assign n27102 = ~n3561 & ~n27101;
  assign n27103 = ~controllable_hgrant2 & ~n27102;
  assign n27104 = ~n4562 & ~n27103;
  assign n27105 = controllable_hmaster0 & ~n27104;
  assign n27106 = ~controllable_hmaster0 & ~n27075;
  assign n27107 = ~n27105 & ~n27106;
  assign n27108 = controllable_hmaster1 & ~n27107;
  assign n27109 = controllable_hmaster0 & ~n27075;
  assign n27110 = ~i_hbusreq2 & ~n11122;
  assign n27111 = ~n26969 & ~n27110;
  assign n27112 = ~controllable_hgrant2 & ~n27111;
  assign n27113 = ~n3410 & ~n27112;
  assign n27114 = ~controllable_hmaster0 & ~n27113;
  assign n27115 = ~n27109 & ~n27114;
  assign n27116 = ~controllable_hmaster1 & ~n27115;
  assign n27117 = ~n27108 & ~n27116;
  assign n27118 = i_hlock3 & ~n27117;
  assign n27119 = i_hbusreq2 & ~n11063;
  assign n27120 = ~i_hbusreq2 & ~n11105;
  assign n27121 = ~n27119 & ~n27120;
  assign n27122 = ~controllable_hgrant2 & ~n27121;
  assign n27123 = ~n4562 & ~n27122;
  assign n27124 = controllable_hmaster0 & ~n27123;
  assign n27125 = ~controllable_hmaster0 & ~n27080;
  assign n27126 = ~n27124 & ~n27125;
  assign n27127 = controllable_hmaster1 & ~n27126;
  assign n27128 = controllable_hmaster0 & ~n27080;
  assign n27129 = ~n26955 & ~n27128;
  assign n27130 = ~controllable_hmaster1 & ~n27129;
  assign n27131 = ~n27127 & ~n27130;
  assign n27132 = ~i_hlock3 & ~n27131;
  assign n27133 = ~n27118 & ~n27132;
  assign n27134 = ~i_hbusreq3 & ~n27133;
  assign n27135 = ~n27100 & ~n27134;
  assign n27136 = ~controllable_hmaster2 & ~n27135;
  assign n27137 = ~n27085 & ~n27136;
  assign n27138 = controllable_hgrant3 & ~n27137;
  assign n27139 = ~n10194 & ~n27138;
  assign n27140 = controllable_nhgrant0 & ~n27139;
  assign n27141 = ~n10240 & ~n27140;
  assign n27142 = ~n3281 & ~n27141;
  assign n27143 = ~n3281 & ~n27142;
  assign n27144 = ~n3378 & ~n27143;
  assign n27145 = ~n27067 & ~n27144;
  assign n27146 = n3492 & ~n27145;
  assign n27147 = ~n26477 & ~n27146;
  assign n27148 = n3485 & ~n27147;
  assign n27149 = ~n26634 & ~n27148;
  assign n27150 = n3476 & ~n27149;
  assign n27151 = ~n26937 & ~n27150;
  assign n27152 = n3374 & ~n27151;
  assign n27153 = ~n26909 & ~n27152;
  assign n27154 = n3655 & ~n27153;
  assign n27155 = n3378 & ~n25970;
  assign n27156 = ~n10293 & ~n26891;
  assign n27157 = controllable_nhgrant0 & ~n27156;
  assign n27158 = ~n9753 & ~n27157;
  assign n27159 = ~n3281 & ~n27158;
  assign n27160 = ~n3281 & ~n27159;
  assign n27161 = ~n3378 & ~n27160;
  assign n27162 = ~n27155 & ~n27161;
  assign n27163 = n3492 & ~n27162;
  assign n27164 = n3492 & ~n27163;
  assign n27165 = n3485 & ~n27164;
  assign n27166 = n3485 & ~n27165;
  assign n27167 = ~n3476 & ~n27166;
  assign n27168 = ~n8523 & ~n27163;
  assign n27169 = n3485 & ~n27168;
  assign n27170 = ~n8689 & ~n27169;
  assign n27171 = n3476 & ~n27170;
  assign n27172 = ~n27167 & ~n27171;
  assign n27173 = ~n3374 & ~n27172;
  assign n27174 = n3378 & ~n25988;
  assign n27175 = ~n10384 & ~n26925;
  assign n27176 = controllable_nhgrant0 & ~n27175;
  assign n27177 = ~n9861 & ~n27176;
  assign n27178 = ~n3281 & ~n27177;
  assign n27179 = ~n3281 & ~n27178;
  assign n27180 = ~n3378 & ~n27179;
  assign n27181 = ~n27174 & ~n27180;
  assign n27182 = n3492 & ~n27181;
  assign n27183 = n3492 & ~n27182;
  assign n27184 = n3485 & ~n27183;
  assign n27185 = n3485 & ~n27184;
  assign n27186 = ~n3476 & ~n27185;
  assign n27187 = ~n10581 & ~n27061;
  assign n27188 = controllable_nhgrant0 & ~n27187;
  assign n27189 = ~n10071 & ~n27188;
  assign n27190 = ~n3281 & ~n27189;
  assign n27191 = ~n3281 & ~n27190;
  assign n27192 = n3378 & ~n27191;
  assign n27193 = ~n10699 & ~n27138;
  assign n27194 = controllable_nhgrant0 & ~n27193;
  assign n27195 = ~n10240 & ~n27194;
  assign n27196 = ~n3281 & ~n27195;
  assign n27197 = ~n3281 & ~n27196;
  assign n27198 = ~n3378 & ~n27197;
  assign n27199 = ~n27192 & ~n27198;
  assign n27200 = n3492 & ~n27199;
  assign n27201 = ~n26504 & ~n27200;
  assign n27202 = n3485 & ~n27201;
  assign n27203 = ~n26645 & ~n27202;
  assign n27204 = n3476 & ~n27203;
  assign n27205 = ~n27186 & ~n27204;
  assign n27206 = n3374 & ~n27205;
  assign n27207 = ~n27173 & ~n27206;
  assign n27208 = ~n3655 & ~n27207;
  assign n27209 = ~n27154 & ~n27208;
  assign n27210 = n3652 & ~n27209;
  assign n27211 = n3378 & ~n26024;
  assign n27212 = ~n10736 & ~n26891;
  assign n27213 = controllable_nhgrant0 & ~n27212;
  assign n27214 = ~n9753 & ~n27213;
  assign n27215 = ~n3281 & ~n27214;
  assign n27216 = ~n3281 & ~n27215;
  assign n27217 = ~n3378 & ~n27216;
  assign n27218 = ~n27211 & ~n27217;
  assign n27219 = n3492 & ~n27218;
  assign n27220 = n3492 & ~n27219;
  assign n27221 = n3485 & ~n27220;
  assign n27222 = n3485 & ~n27221;
  assign n27223 = ~n3476 & ~n27222;
  assign n27224 = ~n8523 & ~n27219;
  assign n27225 = n3485 & ~n27224;
  assign n27226 = ~n8689 & ~n27225;
  assign n27227 = n3476 & ~n27226;
  assign n27228 = ~n27223 & ~n27227;
  assign n27229 = ~n3374 & ~n27228;
  assign n27230 = n3378 & ~n26042;
  assign n27231 = ~n10796 & ~n26925;
  assign n27232 = controllable_nhgrant0 & ~n27231;
  assign n27233 = ~n9861 & ~n27232;
  assign n27234 = ~n3281 & ~n27233;
  assign n27235 = ~n3281 & ~n27234;
  assign n27236 = ~n3378 & ~n27235;
  assign n27237 = ~n27230 & ~n27236;
  assign n27238 = n3492 & ~n27237;
  assign n27239 = n3492 & ~n27238;
  assign n27240 = n3485 & ~n27239;
  assign n27241 = n3485 & ~n27240;
  assign n27242 = ~n3476 & ~n27241;
  assign n27243 = ~n11012 & ~n27061;
  assign n27244 = controllable_nhgrant0 & ~n27243;
  assign n27245 = ~n10071 & ~n27244;
  assign n27246 = ~n3281 & ~n27245;
  assign n27247 = ~n3281 & ~n27246;
  assign n27248 = n3378 & ~n27247;
  assign n27249 = ~n11137 & ~n27138;
  assign n27250 = controllable_nhgrant0 & ~n27249;
  assign n27251 = ~n10240 & ~n27250;
  assign n27252 = ~n3281 & ~n27251;
  assign n27253 = ~n3281 & ~n27252;
  assign n27254 = ~n3378 & ~n27253;
  assign n27255 = ~n27248 & ~n27254;
  assign n27256 = n3492 & ~n27255;
  assign n27257 = ~n26533 & ~n27256;
  assign n27258 = n3485 & ~n27257;
  assign n27259 = ~n26658 & ~n27258;
  assign n27260 = n3476 & ~n27259;
  assign n27261 = ~n27242 & ~n27260;
  assign n27262 = n3374 & ~n27261;
  assign n27263 = ~n27229 & ~n27262;
  assign n27264 = n3655 & ~n27263;
  assign n27265 = n3378 & ~n26076;
  assign n27266 = ~n11172 & ~n26891;
  assign n27267 = controllable_nhgrant0 & ~n27266;
  assign n27268 = ~n9753 & ~n27267;
  assign n27269 = ~n3281 & ~n27268;
  assign n27270 = ~n3281 & ~n27269;
  assign n27271 = ~n3378 & ~n27270;
  assign n27272 = ~n27265 & ~n27271;
  assign n27273 = n3492 & ~n27272;
  assign n27274 = n3492 & ~n27273;
  assign n27275 = n3485 & ~n27274;
  assign n27276 = n3485 & ~n27275;
  assign n27277 = ~n3476 & ~n27276;
  assign n27278 = ~n8523 & ~n27273;
  assign n27279 = n3485 & ~n27278;
  assign n27280 = ~n8689 & ~n27279;
  assign n27281 = n3476 & ~n27280;
  assign n27282 = ~n27277 & ~n27281;
  assign n27283 = ~n3374 & ~n27282;
  assign n27284 = n3378 & ~n26094;
  assign n27285 = ~n11230 & ~n26925;
  assign n27286 = controllable_nhgrant0 & ~n27285;
  assign n27287 = ~n9861 & ~n27286;
  assign n27288 = ~n3281 & ~n27287;
  assign n27289 = ~n3281 & ~n27288;
  assign n27290 = ~n3378 & ~n27289;
  assign n27291 = ~n27284 & ~n27290;
  assign n27292 = n3492 & ~n27291;
  assign n27293 = n3492 & ~n27292;
  assign n27294 = n3485 & ~n27293;
  assign n27295 = n3485 & ~n27294;
  assign n27296 = ~n3476 & ~n27295;
  assign n27297 = ~n11293 & ~n27061;
  assign n27298 = controllable_nhgrant0 & ~n27297;
  assign n27299 = ~n10071 & ~n27298;
  assign n27300 = ~n3281 & ~n27299;
  assign n27301 = ~n3281 & ~n27300;
  assign n27302 = n3378 & ~n27301;
  assign n27303 = ~n11346 & ~n27138;
  assign n27304 = controllable_nhgrant0 & ~n27303;
  assign n27305 = ~n10240 & ~n27304;
  assign n27306 = ~n3281 & ~n27305;
  assign n27307 = ~n3281 & ~n27306;
  assign n27308 = ~n3378 & ~n27307;
  assign n27309 = ~n27302 & ~n27308;
  assign n27310 = n3492 & ~n27309;
  assign n27311 = ~n26560 & ~n27310;
  assign n27312 = n3485 & ~n27311;
  assign n27313 = ~n26669 & ~n27312;
  assign n27314 = n3476 & ~n27313;
  assign n27315 = ~n27296 & ~n27314;
  assign n27316 = n3374 & ~n27315;
  assign n27317 = ~n27283 & ~n27316;
  assign n27318 = ~n3655 & ~n27317;
  assign n27319 = ~n27264 & ~n27318;
  assign n27320 = ~n3652 & ~n27319;
  assign n27321 = ~n27210 & ~n27320;
  assign n27322 = n3368 & ~n27321;
  assign n27323 = ~n26889 & ~n27322;
  assign n27324 = ~n3362 & ~n27323;
  assign n27325 = ~n26681 & ~n27324;
  assign n27326 = ~n3359 & ~n27325;
  assign n27327 = ~n26579 & ~n27326;
  assign n27328 = ~n3356 & ~n27327;
  assign n27329 = ~n25607 & ~n27328;
  assign n27330 = n3345 & ~n27329;
  assign n27331 = ~n3649 & ~n27330;
  assign n27332 = ~n3341 & ~n27331;
  assign n27333 = controllable_hmaster1 & ~n26136;
  assign n27334 = i_hlock3 & ~n27333;
  assign n27335 = controllable_hmaster1 & ~n26140;
  assign n27336 = ~i_hlock3 & ~n27335;
  assign n27337 = ~n27334 & ~n27336;
  assign n27338 = i_hbusreq3 & ~n27337;
  assign n27339 = controllable_hmaster1 & ~n26146;
  assign n27340 = i_hlock3 & ~n27339;
  assign n27341 = controllable_hmaster1 & ~n26150;
  assign n27342 = ~i_hlock3 & ~n27341;
  assign n27343 = ~n27340 & ~n27342;
  assign n27344 = ~i_hbusreq3 & ~n27343;
  assign n27345 = ~n27338 & ~n27344;
  assign n27346 = ~controllable_hmaster2 & ~n27345;
  assign n27347 = ~controllable_hmaster2 & ~n27346;
  assign n27348 = controllable_hgrant3 & ~n27347;
  assign n27349 = ~n11424 & ~n27348;
  assign n27350 = controllable_nhgrant0 & ~n27349;
  assign n27351 = ~n11427 & ~n27350;
  assign n27352 = ~n3281 & ~n27351;
  assign n27353 = ~n3281 & ~n27352;
  assign n27354 = n3378 & ~n27353;
  assign n27355 = i_hbusreq3 & ~n21271;
  assign n27356 = ~controllable_hgrant2 & ~n14398;
  assign n27357 = ~n3431 & ~n27356;
  assign n27358 = controllable_hmaster1 & ~n27357;
  assign n27359 = controllable_hmaster0 & ~n27357;
  assign n27360 = controllable_hmaster0 & ~n27359;
  assign n27361 = ~controllable_hmaster1 & ~n27360;
  assign n27362 = ~n27358 & ~n27361;
  assign n27363 = ~i_hbusreq3 & ~n27362;
  assign n27364 = ~n27355 & ~n27363;
  assign n27365 = controllable_hmaster2 & ~n27364;
  assign n27366 = ~n27346 & ~n27365;
  assign n27367 = controllable_hgrant3 & ~n27366;
  assign n27368 = ~n11435 & ~n27367;
  assign n27369 = controllable_nhgrant0 & ~n27368;
  assign n27370 = ~n11439 & ~n27369;
  assign n27371 = ~n3281 & ~n27370;
  assign n27372 = ~n3783 & ~n27371;
  assign n27373 = ~n3378 & ~n27372;
  assign n27374 = ~n27354 & ~n27373;
  assign n27375 = n3492 & ~n27374;
  assign n27376 = ~n3493 & ~n27375;
  assign n27377 = n3485 & ~n27376;
  assign n27378 = ~n3486 & ~n27377;
  assign n27379 = ~n3476 & ~n27378;
  assign n27380 = ~n3407 & ~n27346;
  assign n27381 = controllable_hgrant3 & ~n27380;
  assign n27382 = ~n11435 & ~n27381;
  assign n27383 = controllable_nhgrant0 & ~n27382;
  assign n27384 = ~n11439 & ~n27383;
  assign n27385 = ~n3281 & ~n27384;
  assign n27386 = ~n3783 & ~n27385;
  assign n27387 = ~n3378 & ~n27386;
  assign n27388 = ~n27354 & ~n27387;
  assign n27389 = ~n3485 & ~n27388;
  assign n27390 = ~n3492 & ~n27388;
  assign n27391 = ~n27375 & ~n27390;
  assign n27392 = n3485 & ~n27391;
  assign n27393 = ~n27389 & ~n27392;
  assign n27394 = n3476 & ~n27393;
  assign n27395 = ~n27379 & ~n27394;
  assign n27396 = ~n3374 & ~n27395;
  assign n27397 = controllable_hmaster1 & ~n7091;
  assign n27398 = controllable_hmaster1 & ~n27397;
  assign n27399 = i_hbusreq3 & ~n27398;
  assign n27400 = controllable_hmaster1 & ~n7095;
  assign n27401 = controllable_hmaster1 & ~n27400;
  assign n27402 = ~i_hbusreq3 & ~n27401;
  assign n27403 = ~n27399 & ~n27402;
  assign n27404 = ~controllable_hmaster2 & ~n27403;
  assign n27405 = ~controllable_hmaster2 & ~n27404;
  assign n27406 = controllable_hgrant3 & ~n27405;
  assign n27407 = ~n11472 & ~n27406;
  assign n27408 = controllable_nhgrant0 & ~n27407;
  assign n27409 = ~n11496 & ~n27408;
  assign n27410 = ~n3281 & ~n27409;
  assign n27411 = ~n3281 & ~n27410;
  assign n27412 = n3378 & ~n27411;
  assign n27413 = ~n27365 & ~n27404;
  assign n27414 = controllable_hgrant3 & ~n27413;
  assign n27415 = ~n11504 & ~n27414;
  assign n27416 = controllable_nhgrant0 & ~n27415;
  assign n27417 = ~n11512 & ~n27416;
  assign n27418 = ~n3281 & ~n27417;
  assign n27419 = ~n3950 & ~n27418;
  assign n27420 = ~n3378 & ~n27419;
  assign n27421 = ~n27412 & ~n27420;
  assign n27422 = n3492 & ~n27421;
  assign n27423 = ~n3493 & ~n27422;
  assign n27424 = n3485 & ~n27423;
  assign n27425 = ~n3486 & ~n27424;
  assign n27426 = ~n3476 & ~n27425;
  assign n27427 = ~n21446 & ~n25705;
  assign n27428 = controllable_hmaster1 & ~n27427;
  assign n27429 = ~controllable_hmaster1 & ~n21359;
  assign n27430 = ~n27428 & ~n27429;
  assign n27431 = i_hbusreq3 & ~n27430;
  assign n27432 = ~n21451 & ~n25713;
  assign n27433 = controllable_hmaster1 & ~n27432;
  assign n27434 = ~controllable_hmaster1 & ~n21362;
  assign n27435 = ~n27433 & ~n27434;
  assign n27436 = ~i_hbusreq3 & ~n27435;
  assign n27437 = ~n27431 & ~n27436;
  assign n27438 = ~controllable_hmaster2 & ~n27437;
  assign n27439 = ~n21365 & ~n27438;
  assign n27440 = controllable_hgrant3 & ~n27439;
  assign n27441 = ~n11472 & ~n27440;
  assign n27442 = controllable_nhgrant0 & ~n27441;
  assign n27443 = ~n11496 & ~n27442;
  assign n27444 = ~n3281 & ~n27443;
  assign n27445 = ~n3281 & ~n27444;
  assign n27446 = n3378 & ~n27445;
  assign n27447 = ~controllable_hgrant2 & ~n14558;
  assign n27448 = ~n3431 & ~n27447;
  assign n27449 = controllable_hmaster1 & ~n27448;
  assign n27450 = controllable_hmaster0 & ~n27448;
  assign n27451 = ~n21451 & ~n27450;
  assign n27452 = ~controllable_hmaster1 & ~n27451;
  assign n27453 = ~n27449 & ~n27452;
  assign n27454 = ~i_hbusreq3 & ~n27453;
  assign n27455 = ~n21450 & ~n27454;
  assign n27456 = controllable_hmaster2 & ~n27455;
  assign n27457 = ~n27438 & ~n27456;
  assign n27458 = controllable_hgrant3 & ~n27457;
  assign n27459 = ~n11598 & ~n27458;
  assign n27460 = controllable_nhgrant0 & ~n27459;
  assign n27461 = ~n11512 & ~n27460;
  assign n27462 = ~n3281 & ~n27461;
  assign n27463 = ~n4089 & ~n27462;
  assign n27464 = ~n3378 & ~n27463;
  assign n27465 = ~n27446 & ~n27464;
  assign n27466 = n3492 & ~n27465;
  assign n27467 = ~n27390 & ~n27466;
  assign n27468 = n3485 & ~n27467;
  assign n27469 = ~n27389 & ~n27468;
  assign n27470 = n3476 & ~n27469;
  assign n27471 = ~n27426 & ~n27470;
  assign n27472 = n3374 & ~n27471;
  assign n27473 = ~n27396 & ~n27472;
  assign n27474 = n3655 & ~n27473;
  assign n27475 = ~n11626 & ~n27406;
  assign n27476 = controllable_nhgrant0 & ~n27475;
  assign n27477 = ~n11496 & ~n27476;
  assign n27478 = ~n3281 & ~n27477;
  assign n27479 = ~n3281 & ~n27478;
  assign n27480 = n3378 & ~n27479;
  assign n27481 = ~n11634 & ~n27414;
  assign n27482 = controllable_nhgrant0 & ~n27481;
  assign n27483 = ~n11512 & ~n27482;
  assign n27484 = ~n3281 & ~n27483;
  assign n27485 = ~n3950 & ~n27484;
  assign n27486 = ~n3378 & ~n27485;
  assign n27487 = ~n27480 & ~n27486;
  assign n27488 = n3492 & ~n27487;
  assign n27489 = ~n3493 & ~n27488;
  assign n27490 = n3485 & ~n27489;
  assign n27491 = ~n3486 & ~n27490;
  assign n27492 = ~n3476 & ~n27491;
  assign n27493 = ~n11626 & ~n27440;
  assign n27494 = controllable_nhgrant0 & ~n27493;
  assign n27495 = ~n11496 & ~n27494;
  assign n27496 = ~n3281 & ~n27495;
  assign n27497 = ~n3281 & ~n27496;
  assign n27498 = n3378 & ~n27497;
  assign n27499 = ~n11675 & ~n27458;
  assign n27500 = controllable_nhgrant0 & ~n27499;
  assign n27501 = ~n11512 & ~n27500;
  assign n27502 = ~n3281 & ~n27501;
  assign n27503 = ~n4089 & ~n27502;
  assign n27504 = ~n3378 & ~n27503;
  assign n27505 = ~n27498 & ~n27504;
  assign n27506 = n3492 & ~n27505;
  assign n27507 = ~n27390 & ~n27506;
  assign n27508 = n3485 & ~n27507;
  assign n27509 = ~n27389 & ~n27508;
  assign n27510 = n3476 & ~n27509;
  assign n27511 = ~n27492 & ~n27510;
  assign n27512 = n3374 & ~n27511;
  assign n27513 = ~n27396 & ~n27512;
  assign n27514 = ~n3655 & ~n27513;
  assign n27515 = ~n27474 & ~n27514;
  assign n27516 = n3652 & ~n27515;
  assign n27517 = ~n11705 & ~n27406;
  assign n27518 = controllable_nhgrant0 & ~n27517;
  assign n27519 = ~n11496 & ~n27518;
  assign n27520 = ~n3281 & ~n27519;
  assign n27521 = ~n3281 & ~n27520;
  assign n27522 = n3378 & ~n27521;
  assign n27523 = ~n11713 & ~n27414;
  assign n27524 = controllable_nhgrant0 & ~n27523;
  assign n27525 = ~n11512 & ~n27524;
  assign n27526 = ~n3281 & ~n27525;
  assign n27527 = ~n3950 & ~n27526;
  assign n27528 = ~n3378 & ~n27527;
  assign n27529 = ~n27522 & ~n27528;
  assign n27530 = n3492 & ~n27529;
  assign n27531 = ~n3493 & ~n27530;
  assign n27532 = n3485 & ~n27531;
  assign n27533 = ~n3486 & ~n27532;
  assign n27534 = ~n3476 & ~n27533;
  assign n27535 = ~n11705 & ~n27440;
  assign n27536 = controllable_nhgrant0 & ~n27535;
  assign n27537 = ~n11496 & ~n27536;
  assign n27538 = ~n3281 & ~n27537;
  assign n27539 = ~n3281 & ~n27538;
  assign n27540 = n3378 & ~n27539;
  assign n27541 = ~n11747 & ~n27458;
  assign n27542 = controllable_nhgrant0 & ~n27541;
  assign n27543 = ~n11512 & ~n27542;
  assign n27544 = ~n3281 & ~n27543;
  assign n27545 = ~n4089 & ~n27544;
  assign n27546 = ~n3378 & ~n27545;
  assign n27547 = ~n27540 & ~n27546;
  assign n27548 = n3492 & ~n27547;
  assign n27549 = ~n27390 & ~n27548;
  assign n27550 = n3485 & ~n27549;
  assign n27551 = ~n27389 & ~n27550;
  assign n27552 = n3476 & ~n27551;
  assign n27553 = ~n27534 & ~n27552;
  assign n27554 = n3374 & ~n27553;
  assign n27555 = ~n27396 & ~n27554;
  assign n27556 = n3655 & ~n27555;
  assign n27557 = ~n11775 & ~n27406;
  assign n27558 = controllable_nhgrant0 & ~n27557;
  assign n27559 = ~n11496 & ~n27558;
  assign n27560 = ~n3281 & ~n27559;
  assign n27561 = ~n3281 & ~n27560;
  assign n27562 = n3378 & ~n27561;
  assign n27563 = ~n11783 & ~n27414;
  assign n27564 = controllable_nhgrant0 & ~n27563;
  assign n27565 = ~n11512 & ~n27564;
  assign n27566 = ~n3281 & ~n27565;
  assign n27567 = ~n3950 & ~n27566;
  assign n27568 = ~n3378 & ~n27567;
  assign n27569 = ~n27562 & ~n27568;
  assign n27570 = n3492 & ~n27569;
  assign n27571 = ~n3493 & ~n27570;
  assign n27572 = n3485 & ~n27571;
  assign n27573 = ~n3486 & ~n27572;
  assign n27574 = ~n3476 & ~n27573;
  assign n27575 = ~n11775 & ~n27440;
  assign n27576 = controllable_nhgrant0 & ~n27575;
  assign n27577 = ~n11496 & ~n27576;
  assign n27578 = ~n3281 & ~n27577;
  assign n27579 = ~n3281 & ~n27578;
  assign n27580 = n3378 & ~n27579;
  assign n27581 = ~n11817 & ~n27458;
  assign n27582 = controllable_nhgrant0 & ~n27581;
  assign n27583 = ~n11512 & ~n27582;
  assign n27584 = ~n3281 & ~n27583;
  assign n27585 = ~n4089 & ~n27584;
  assign n27586 = ~n3378 & ~n27585;
  assign n27587 = ~n27580 & ~n27586;
  assign n27588 = n3492 & ~n27587;
  assign n27589 = ~n27390 & ~n27588;
  assign n27590 = n3485 & ~n27589;
  assign n27591 = ~n27389 & ~n27590;
  assign n27592 = n3476 & ~n27591;
  assign n27593 = ~n27574 & ~n27592;
  assign n27594 = n3374 & ~n27593;
  assign n27595 = ~n27396 & ~n27594;
  assign n27596 = ~n3655 & ~n27595;
  assign n27597 = ~n27556 & ~n27596;
  assign n27598 = ~n3652 & ~n27597;
  assign n27599 = ~n27516 & ~n27598;
  assign n27600 = ~n3368 & ~n27599;
  assign n27601 = controllable_hmaster1 & ~n3503;
  assign n27602 = controllable_hmaster1 & ~n27601;
  assign n27603 = i_hbusreq3 & ~n27602;
  assign n27604 = controllable_hmaster1 & ~n9726;
  assign n27605 = controllable_hmaster1 & ~n27604;
  assign n27606 = ~i_hbusreq3 & ~n27605;
  assign n27607 = ~n27603 & ~n27606;
  assign n27608 = ~controllable_hmaster2 & ~n27607;
  assign n27609 = ~controllable_hmaster2 & ~n27608;
  assign n27610 = controllable_hgrant3 & ~n27609;
  assign n27611 = ~n11853 & ~n27610;
  assign n27612 = controllable_nhgrant0 & ~n27611;
  assign n27613 = ~n11874 & ~n27612;
  assign n27614 = ~n3281 & ~n27613;
  assign n27615 = ~n3281 & ~n27614;
  assign n27616 = n3492 & ~n27615;
  assign n27617 = n3492 & ~n27616;
  assign n27618 = n3485 & ~n27617;
  assign n27619 = n3485 & ~n27618;
  assign n27620 = ~n3476 & ~n27619;
  assign n27621 = ~n3485 & ~n27353;
  assign n27622 = ~n3492 & ~n27353;
  assign n27623 = i_hlock3 & ~n3555;
  assign n27624 = ~controllable_hgrant2 & ~n14840;
  assign n27625 = ~controllable_hgrant2 & ~n27624;
  assign n27626 = ~i_hlock3 & ~n27625;
  assign n27627 = ~n27623 & ~n27626;
  assign n27628 = i_hbusreq3 & ~n27627;
  assign n27629 = i_hlock3 & ~n21403;
  assign n27630 = ~n27626 & ~n27629;
  assign n27631 = ~i_hbusreq3 & ~n27630;
  assign n27632 = ~n27628 & ~n27631;
  assign n27633 = controllable_hmaster2 & ~n27632;
  assign n27634 = i_hlock3 & ~n11582;
  assign n27635 = ~controllable_hmaster0 & ~n27625;
  assign n27636 = ~n27093 & ~n27635;
  assign n27637 = controllable_hmaster1 & ~n27636;
  assign n27638 = ~controllable_hmaster1 & ~n27625;
  assign n27639 = ~n27637 & ~n27638;
  assign n27640 = ~i_hlock3 & ~n27639;
  assign n27641 = ~n27634 & ~n27640;
  assign n27642 = i_hbusreq3 & ~n27641;
  assign n27643 = ~n21404 & ~n27105;
  assign n27644 = controllable_hmaster1 & ~n27643;
  assign n27645 = ~controllable_hmaster1 & ~n21403;
  assign n27646 = ~n27644 & ~n27645;
  assign n27647 = i_hlock3 & ~n27646;
  assign n27648 = ~n27124 & ~n27635;
  assign n27649 = controllable_hmaster1 & ~n27648;
  assign n27650 = ~n27638 & ~n27649;
  assign n27651 = ~i_hlock3 & ~n27650;
  assign n27652 = ~n27647 & ~n27651;
  assign n27653 = ~i_hbusreq3 & ~n27652;
  assign n27654 = ~n27642 & ~n27653;
  assign n27655 = ~controllable_hmaster2 & ~n27654;
  assign n27656 = ~n27633 & ~n27655;
  assign n27657 = controllable_hgrant3 & ~n27656;
  assign n27658 = ~n11853 & ~n27657;
  assign n27659 = controllable_nhgrant0 & ~n27658;
  assign n27660 = ~n11874 & ~n27659;
  assign n27661 = ~n3281 & ~n27660;
  assign n27662 = ~n3281 & ~n27661;
  assign n27663 = n3492 & ~n27662;
  assign n27664 = ~n27622 & ~n27663;
  assign n27665 = n3485 & ~n27664;
  assign n27666 = ~n27621 & ~n27665;
  assign n27667 = n3476 & ~n27666;
  assign n27668 = ~n27620 & ~n27667;
  assign n27669 = n3374 & ~n27668;
  assign n27670 = n3374 & ~n27669;
  assign n27671 = n3655 & ~n27670;
  assign n27672 = ~n11917 & ~n27610;
  assign n27673 = controllable_nhgrant0 & ~n27672;
  assign n27674 = ~n11874 & ~n27673;
  assign n27675 = ~n3281 & ~n27674;
  assign n27676 = ~n3281 & ~n27675;
  assign n27677 = n3492 & ~n27676;
  assign n27678 = n3492 & ~n27677;
  assign n27679 = n3485 & ~n27678;
  assign n27680 = n3485 & ~n27679;
  assign n27681 = ~n3476 & ~n27680;
  assign n27682 = ~n11917 & ~n27657;
  assign n27683 = controllable_nhgrant0 & ~n27682;
  assign n27684 = ~n11874 & ~n27683;
  assign n27685 = ~n3281 & ~n27684;
  assign n27686 = ~n3281 & ~n27685;
  assign n27687 = n3492 & ~n27686;
  assign n27688 = ~n27622 & ~n27687;
  assign n27689 = n3485 & ~n27688;
  assign n27690 = ~n27621 & ~n27689;
  assign n27691 = n3476 & ~n27690;
  assign n27692 = ~n27681 & ~n27691;
  assign n27693 = n3374 & ~n27692;
  assign n27694 = n3374 & ~n27693;
  assign n27695 = ~n3655 & ~n27694;
  assign n27696 = ~n27671 & ~n27695;
  assign n27697 = n3652 & ~n27696;
  assign n27698 = ~n11955 & ~n27610;
  assign n27699 = controllable_nhgrant0 & ~n27698;
  assign n27700 = ~n11874 & ~n27699;
  assign n27701 = ~n3281 & ~n27700;
  assign n27702 = ~n3281 & ~n27701;
  assign n27703 = n3492 & ~n27702;
  assign n27704 = n3492 & ~n27703;
  assign n27705 = n3485 & ~n27704;
  assign n27706 = n3485 & ~n27705;
  assign n27707 = ~n3476 & ~n27706;
  assign n27708 = ~n11955 & ~n27657;
  assign n27709 = controllable_nhgrant0 & ~n27708;
  assign n27710 = ~n11874 & ~n27709;
  assign n27711 = ~n3281 & ~n27710;
  assign n27712 = ~n3281 & ~n27711;
  assign n27713 = n3492 & ~n27712;
  assign n27714 = ~n27622 & ~n27713;
  assign n27715 = n3485 & ~n27714;
  assign n27716 = ~n27621 & ~n27715;
  assign n27717 = n3476 & ~n27716;
  assign n27718 = ~n27707 & ~n27717;
  assign n27719 = n3374 & ~n27718;
  assign n27720 = n3374 & ~n27719;
  assign n27721 = n3655 & ~n27720;
  assign n27722 = ~n11991 & ~n27610;
  assign n27723 = controllable_nhgrant0 & ~n27722;
  assign n27724 = ~n11874 & ~n27723;
  assign n27725 = ~n3281 & ~n27724;
  assign n27726 = ~n3281 & ~n27725;
  assign n27727 = n3492 & ~n27726;
  assign n27728 = n3492 & ~n27727;
  assign n27729 = n3485 & ~n27728;
  assign n27730 = n3485 & ~n27729;
  assign n27731 = ~n3476 & ~n27730;
  assign n27732 = ~n11991 & ~n27657;
  assign n27733 = controllable_nhgrant0 & ~n27732;
  assign n27734 = ~n11874 & ~n27733;
  assign n27735 = ~n3281 & ~n27734;
  assign n27736 = ~n3281 & ~n27735;
  assign n27737 = n3492 & ~n27736;
  assign n27738 = ~n27622 & ~n27737;
  assign n27739 = n3485 & ~n27738;
  assign n27740 = ~n27621 & ~n27739;
  assign n27741 = n3476 & ~n27740;
  assign n27742 = ~n27731 & ~n27741;
  assign n27743 = n3374 & ~n27742;
  assign n27744 = n3374 & ~n27743;
  assign n27745 = ~n3655 & ~n27744;
  assign n27746 = ~n27721 & ~n27745;
  assign n27747 = ~n3652 & ~n27746;
  assign n27748 = ~n27697 & ~n27747;
  assign n27749 = n3368 & ~n27748;
  assign n27750 = ~n27600 & ~n27749;
  assign n27751 = ~n3362 & ~n27750;
  assign n27752 = ~n3362 & ~n27751;
  assign n27753 = ~n3359 & ~n27752;
  assign n27754 = ~n3359 & ~n27753;
  assign n27755 = n3356 & ~n27754;
  assign n27756 = n3378 & ~n27372;
  assign n27757 = controllable_hmaster1 & ~n8837;
  assign n27758 = ~n3697 & ~n8838;
  assign n27759 = ~controllable_hmaster1 & ~n27758;
  assign n27760 = ~n27757 & ~n27759;
  assign n27761 = ~i_hbusreq3 & ~n27760;
  assign n27762 = ~n8775 & ~n27761;
  assign n27763 = controllable_hmaster2 & ~n27762;
  assign n27764 = ~n25647 & ~n27763;
  assign n27765 = controllable_hgrant3 & ~n27764;
  assign n27766 = ~n5163 & ~n27765;
  assign n27767 = controllable_nhgrant0 & ~n27766;
  assign n27768 = ~n5245 & ~n27767;
  assign n27769 = ~n3281 & ~n27768;
  assign n27770 = ~n3783 & ~n27769;
  assign n27771 = ~n3378 & ~n27770;
  assign n27772 = ~n27756 & ~n27771;
  assign n27773 = n3492 & ~n27772;
  assign n27774 = ~n3631 & ~n27773;
  assign n27775 = n3485 & ~n27774;
  assign n27776 = ~n3630 & ~n27775;
  assign n27777 = ~n3476 & ~n27776;
  assign n27778 = ~n3485 & ~n27386;
  assign n27779 = ~n3492 & ~n27386;
  assign n27780 = ~n27773 & ~n27779;
  assign n27781 = n3485 & ~n27780;
  assign n27782 = ~n27778 & ~n27781;
  assign n27783 = n3476 & ~n27782;
  assign n27784 = ~n27777 & ~n27783;
  assign n27785 = ~n3374 & ~n27784;
  assign n27786 = ~controllable_hgrant2 & ~n15278;
  assign n27787 = ~n3431 & ~n27786;
  assign n27788 = ~controllable_hmaster0 & ~n27787;
  assign n27789 = ~n27359 & ~n27788;
  assign n27790 = ~controllable_hmaster1 & ~n27789;
  assign n27791 = ~n27358 & ~n27790;
  assign n27792 = ~i_hbusreq3 & ~n27791;
  assign n27793 = ~n8892 & ~n27792;
  assign n27794 = controllable_hmaster2 & ~n27793;
  assign n27795 = ~n5071 & ~n27788;
  assign n27796 = controllable_hmaster1 & ~n27795;
  assign n27797 = ~controllable_hmaster1 & ~n27787;
  assign n27798 = ~n27796 & ~n27797;
  assign n27799 = ~i_hbusreq3 & ~n27798;
  assign n27800 = ~n25674 & ~n27799;
  assign n27801 = ~controllable_hmaster2 & ~n27800;
  assign n27802 = ~n27794 & ~n27801;
  assign n27803 = controllable_hgrant3 & ~n27802;
  assign n27804 = ~n12077 & ~n27803;
  assign n27805 = controllable_nhgrant0 & ~n27804;
  assign n27806 = ~n12101 & ~n27805;
  assign n27807 = ~n3281 & ~n27806;
  assign n27808 = ~n3950 & ~n27807;
  assign n27809 = n3378 & ~n27808;
  assign n27810 = ~n3935 & ~n8838;
  assign n27811 = ~controllable_hmaster1 & ~n27810;
  assign n27812 = ~n27757 & ~n27811;
  assign n27813 = ~i_hbusreq3 & ~n27812;
  assign n27814 = ~n8892 & ~n27813;
  assign n27815 = controllable_hmaster2 & ~n27814;
  assign n27816 = ~n25682 & ~n27815;
  assign n27817 = controllable_hgrant3 & ~n27816;
  assign n27818 = ~n12138 & ~n27817;
  assign n27819 = controllable_nhgrant0 & ~n27818;
  assign n27820 = ~n5534 & ~n27819;
  assign n27821 = ~n3281 & ~n27820;
  assign n27822 = ~n3950 & ~n27821;
  assign n27823 = ~n3378 & ~n27822;
  assign n27824 = ~n27809 & ~n27823;
  assign n27825 = n3492 & ~n27824;
  assign n27826 = ~n3631 & ~n27825;
  assign n27827 = n3485 & ~n27826;
  assign n27828 = ~n3630 & ~n27827;
  assign n27829 = ~n3476 & ~n27828;
  assign n27830 = ~controllable_hgrant2 & ~n15376;
  assign n27831 = ~n3431 & ~n27830;
  assign n27832 = ~controllable_hmaster0 & ~n27831;
  assign n27833 = ~n27450 & ~n27832;
  assign n27834 = ~controllable_hmaster1 & ~n27833;
  assign n27835 = ~n27449 & ~n27834;
  assign n27836 = ~i_hbusreq3 & ~n27835;
  assign n27837 = ~n9066 & ~n27836;
  assign n27838 = controllable_hmaster2 & ~n27837;
  assign n27839 = ~n25713 & ~n27832;
  assign n27840 = controllable_hmaster1 & ~n27839;
  assign n27841 = ~controllable_hmaster1 & ~n27831;
  assign n27842 = ~n27840 & ~n27841;
  assign n27843 = ~i_hbusreq3 & ~n27842;
  assign n27844 = ~n25710 & ~n27843;
  assign n27845 = ~controllable_hmaster2 & ~n27844;
  assign n27846 = ~n27838 & ~n27845;
  assign n27847 = controllable_hgrant3 & ~n27846;
  assign n27848 = ~n12228 & ~n27847;
  assign n27849 = controllable_nhgrant0 & ~n27848;
  assign n27850 = ~n12249 & ~n27849;
  assign n27851 = ~n3281 & ~n27850;
  assign n27852 = ~n4089 & ~n27851;
  assign n27853 = n3378 & ~n27852;
  assign n27854 = ~controllable_hgrant2 & ~n15432;
  assign n27855 = ~n3859 & ~n27854;
  assign n27856 = controllable_hmaster1 & ~n27855;
  assign n27857 = controllable_hmaster0 & ~n27855;
  assign n27858 = ~n9086 & ~n27857;
  assign n27859 = ~controllable_hmaster1 & ~n27858;
  assign n27860 = ~n27856 & ~n27859;
  assign n27861 = ~i_hbusreq3 & ~n27860;
  assign n27862 = ~n9066 & ~n27861;
  assign n27863 = controllable_hmaster2 & ~n27862;
  assign n27864 = ~n25724 & ~n27863;
  assign n27865 = controllable_hgrant3 & ~n27864;
  assign n27866 = ~n12292 & ~n27865;
  assign n27867 = controllable_nhgrant0 & ~n27866;
  assign n27868 = ~n6082 & ~n27867;
  assign n27869 = ~n3281 & ~n27868;
  assign n27870 = ~n4089 & ~n27869;
  assign n27871 = ~n3378 & ~n27870;
  assign n27872 = ~n27853 & ~n27871;
  assign n27873 = n3492 & ~n27872;
  assign n27874 = ~n27779 & ~n27873;
  assign n27875 = n3485 & ~n27874;
  assign n27876 = ~n27778 & ~n27875;
  assign n27877 = n3476 & ~n27876;
  assign n27878 = ~n27829 & ~n27877;
  assign n27879 = n3374 & ~n27878;
  assign n27880 = ~n27785 & ~n27879;
  assign n27881 = n3655 & ~n27880;
  assign n27882 = ~n6190 & ~n27765;
  assign n27883 = controllable_nhgrant0 & ~n27882;
  assign n27884 = ~n5245 & ~n27883;
  assign n27885 = ~n3281 & ~n27884;
  assign n27886 = ~n3783 & ~n27885;
  assign n27887 = ~n3378 & ~n27886;
  assign n27888 = ~n27756 & ~n27887;
  assign n27889 = n3492 & ~n27888;
  assign n27890 = ~n3631 & ~n27889;
  assign n27891 = n3485 & ~n27890;
  assign n27892 = ~n3630 & ~n27891;
  assign n27893 = ~n3476 & ~n27892;
  assign n27894 = ~n27779 & ~n27889;
  assign n27895 = n3485 & ~n27894;
  assign n27896 = ~n27778 & ~n27895;
  assign n27897 = n3476 & ~n27896;
  assign n27898 = ~n27893 & ~n27897;
  assign n27899 = ~n3374 & ~n27898;
  assign n27900 = ~n12326 & ~n27803;
  assign n27901 = controllable_nhgrant0 & ~n27900;
  assign n27902 = ~n12101 & ~n27901;
  assign n27903 = ~n3281 & ~n27902;
  assign n27904 = ~n3950 & ~n27903;
  assign n27905 = n3378 & ~n27904;
  assign n27906 = ~n12365 & ~n27817;
  assign n27907 = controllable_nhgrant0 & ~n27906;
  assign n27908 = ~n5534 & ~n27907;
  assign n27909 = ~n3281 & ~n27908;
  assign n27910 = ~n3950 & ~n27909;
  assign n27911 = ~n3378 & ~n27910;
  assign n27912 = ~n27905 & ~n27911;
  assign n27913 = n3492 & ~n27912;
  assign n27914 = ~n3631 & ~n27913;
  assign n27915 = n3485 & ~n27914;
  assign n27916 = ~n3630 & ~n27915;
  assign n27917 = ~n3476 & ~n27916;
  assign n27918 = ~n12400 & ~n27847;
  assign n27919 = controllable_nhgrant0 & ~n27918;
  assign n27920 = ~n12249 & ~n27919;
  assign n27921 = ~n3281 & ~n27920;
  assign n27922 = ~n4089 & ~n27921;
  assign n27923 = n3378 & ~n27922;
  assign n27924 = ~n12445 & ~n27865;
  assign n27925 = controllable_nhgrant0 & ~n27924;
  assign n27926 = ~n6082 & ~n27925;
  assign n27927 = ~n3281 & ~n27926;
  assign n27928 = ~n4089 & ~n27927;
  assign n27929 = ~n3378 & ~n27928;
  assign n27930 = ~n27923 & ~n27929;
  assign n27931 = n3492 & ~n27930;
  assign n27932 = ~n27779 & ~n27931;
  assign n27933 = n3485 & ~n27932;
  assign n27934 = ~n27778 & ~n27933;
  assign n27935 = n3476 & ~n27934;
  assign n27936 = ~n27917 & ~n27935;
  assign n27937 = n3374 & ~n27936;
  assign n27938 = ~n27899 & ~n27937;
  assign n27939 = ~n3655 & ~n27938;
  assign n27940 = ~n27881 & ~n27939;
  assign n27941 = n3652 & ~n27940;
  assign n27942 = ~n6659 & ~n27765;
  assign n27943 = controllable_nhgrant0 & ~n27942;
  assign n27944 = ~n5245 & ~n27943;
  assign n27945 = ~n3281 & ~n27944;
  assign n27946 = ~n3783 & ~n27945;
  assign n27947 = ~n3378 & ~n27946;
  assign n27948 = ~n27756 & ~n27947;
  assign n27949 = n3492 & ~n27948;
  assign n27950 = ~n3631 & ~n27949;
  assign n27951 = n3485 & ~n27950;
  assign n27952 = ~n3630 & ~n27951;
  assign n27953 = ~n3476 & ~n27952;
  assign n27954 = ~n27779 & ~n27949;
  assign n27955 = n3485 & ~n27954;
  assign n27956 = ~n27778 & ~n27955;
  assign n27957 = n3476 & ~n27956;
  assign n27958 = ~n27953 & ~n27957;
  assign n27959 = ~n3374 & ~n27958;
  assign n27960 = ~n12481 & ~n27803;
  assign n27961 = controllable_nhgrant0 & ~n27960;
  assign n27962 = ~n12101 & ~n27961;
  assign n27963 = ~n3281 & ~n27962;
  assign n27964 = ~n3950 & ~n27963;
  assign n27965 = n3378 & ~n27964;
  assign n27966 = ~n12513 & ~n27817;
  assign n27967 = controllable_nhgrant0 & ~n27966;
  assign n27968 = ~n5534 & ~n27967;
  assign n27969 = ~n3281 & ~n27968;
  assign n27970 = ~n3950 & ~n27969;
  assign n27971 = ~n3378 & ~n27970;
  assign n27972 = ~n27965 & ~n27971;
  assign n27973 = n3492 & ~n27972;
  assign n27974 = ~n3631 & ~n27973;
  assign n27975 = n3485 & ~n27974;
  assign n27976 = ~n3630 & ~n27975;
  assign n27977 = ~n3476 & ~n27976;
  assign n27978 = ~n12541 & ~n27847;
  assign n27979 = controllable_nhgrant0 & ~n27978;
  assign n27980 = ~n12249 & ~n27979;
  assign n27981 = ~n3281 & ~n27980;
  assign n27982 = ~n4089 & ~n27981;
  assign n27983 = n3378 & ~n27982;
  assign n27984 = ~n12575 & ~n27865;
  assign n27985 = controllable_nhgrant0 & ~n27984;
  assign n27986 = ~n6082 & ~n27985;
  assign n27987 = ~n3281 & ~n27986;
  assign n27988 = ~n4089 & ~n27987;
  assign n27989 = ~n3378 & ~n27988;
  assign n27990 = ~n27983 & ~n27989;
  assign n27991 = n3492 & ~n27990;
  assign n27992 = ~n27779 & ~n27991;
  assign n27993 = n3485 & ~n27992;
  assign n27994 = ~n27778 & ~n27993;
  assign n27995 = n3476 & ~n27994;
  assign n27996 = ~n27977 & ~n27995;
  assign n27997 = n3374 & ~n27996;
  assign n27998 = ~n27959 & ~n27997;
  assign n27999 = n3655 & ~n27998;
  assign n28000 = ~n6889 & ~n27765;
  assign n28001 = controllable_nhgrant0 & ~n28000;
  assign n28002 = ~n5245 & ~n28001;
  assign n28003 = ~n3281 & ~n28002;
  assign n28004 = ~n3783 & ~n28003;
  assign n28005 = ~n3378 & ~n28004;
  assign n28006 = ~n27756 & ~n28005;
  assign n28007 = n3492 & ~n28006;
  assign n28008 = ~n3631 & ~n28007;
  assign n28009 = n3485 & ~n28008;
  assign n28010 = ~n3630 & ~n28009;
  assign n28011 = ~n3476 & ~n28010;
  assign n28012 = ~n27779 & ~n28007;
  assign n28013 = n3485 & ~n28012;
  assign n28014 = ~n27778 & ~n28013;
  assign n28015 = n3476 & ~n28014;
  assign n28016 = ~n28011 & ~n28015;
  assign n28017 = ~n3374 & ~n28016;
  assign n28018 = ~n12609 & ~n27803;
  assign n28019 = controllable_nhgrant0 & ~n28018;
  assign n28020 = ~n12101 & ~n28019;
  assign n28021 = ~n3281 & ~n28020;
  assign n28022 = ~n3950 & ~n28021;
  assign n28023 = n3378 & ~n28022;
  assign n28024 = ~n12641 & ~n27817;
  assign n28025 = controllable_nhgrant0 & ~n28024;
  assign n28026 = ~n5534 & ~n28025;
  assign n28027 = ~n3281 & ~n28026;
  assign n28028 = ~n3950 & ~n28027;
  assign n28029 = ~n3378 & ~n28028;
  assign n28030 = ~n28023 & ~n28029;
  assign n28031 = n3492 & ~n28030;
  assign n28032 = ~n3631 & ~n28031;
  assign n28033 = n3485 & ~n28032;
  assign n28034 = ~n3630 & ~n28033;
  assign n28035 = ~n3476 & ~n28034;
  assign n28036 = ~n12669 & ~n27847;
  assign n28037 = controllable_nhgrant0 & ~n28036;
  assign n28038 = ~n12249 & ~n28037;
  assign n28039 = ~n3281 & ~n28038;
  assign n28040 = ~n4089 & ~n28039;
  assign n28041 = n3378 & ~n28040;
  assign n28042 = ~n12703 & ~n27865;
  assign n28043 = controllable_nhgrant0 & ~n28042;
  assign n28044 = ~n6082 & ~n28043;
  assign n28045 = ~n3281 & ~n28044;
  assign n28046 = ~n4089 & ~n28045;
  assign n28047 = ~n3378 & ~n28046;
  assign n28048 = ~n28041 & ~n28047;
  assign n28049 = n3492 & ~n28048;
  assign n28050 = ~n27779 & ~n28049;
  assign n28051 = n3485 & ~n28050;
  assign n28052 = ~n27778 & ~n28051;
  assign n28053 = n3476 & ~n28052;
  assign n28054 = ~n28035 & ~n28053;
  assign n28055 = n3374 & ~n28054;
  assign n28056 = ~n28017 & ~n28055;
  assign n28057 = ~n3655 & ~n28056;
  assign n28058 = ~n27999 & ~n28057;
  assign n28059 = ~n3652 & ~n28058;
  assign n28060 = ~n27941 & ~n28059;
  assign n28061 = ~n3368 & ~n28060;
  assign n28062 = ~controllable_hgrant2 & ~n15995;
  assign n28063 = ~n3431 & ~n28062;
  assign n28064 = controllable_hmaster1 & ~n28063;
  assign n28065 = controllable_hmaster0 & ~n28063;
  assign n28066 = controllable_hmaster0 & ~n28065;
  assign n28067 = ~controllable_hmaster1 & ~n28066;
  assign n28068 = ~n28064 & ~n28067;
  assign n28069 = ~i_hbusreq3 & ~n28068;
  assign n28070 = ~n9741 & ~n28069;
  assign n28071 = controllable_hmaster2 & ~n28070;
  assign n28072 = controllable_hmaster2 & ~n28071;
  assign n28073 = controllable_hgrant3 & ~n28072;
  assign n28074 = ~n7076 & ~n28073;
  assign n28075 = controllable_nhgrant0 & ~n28074;
  assign n28076 = ~n3466 & ~n28075;
  assign n28077 = ~n3281 & ~n28076;
  assign n28078 = ~n3281 & ~n28077;
  assign n28079 = n3378 & ~n28078;
  assign n28080 = ~controllable_hgrant2 & ~n16030;
  assign n28081 = ~n3859 & ~n28080;
  assign n28082 = controllable_hmaster1 & ~n28081;
  assign n28083 = controllable_hmaster0 & ~n28081;
  assign n28084 = controllable_hmaster0 & ~n28083;
  assign n28085 = ~controllable_hmaster1 & ~n28084;
  assign n28086 = ~n28082 & ~n28085;
  assign n28087 = ~i_hbusreq3 & ~n28086;
  assign n28088 = ~n9741 & ~n28087;
  assign n28089 = controllable_hmaster2 & ~n28088;
  assign n28090 = controllable_hmaster2 & ~n28089;
  assign n28091 = controllable_hgrant3 & ~n28090;
  assign n28092 = ~n7102 & ~n28091;
  assign n28093 = controllable_nhgrant0 & ~n28092;
  assign n28094 = ~n7118 & ~n28093;
  assign n28095 = ~n3281 & ~n28094;
  assign n28096 = ~n3281 & ~n28095;
  assign n28097 = ~n3378 & ~n28096;
  assign n28098 = ~n28079 & ~n28097;
  assign n28099 = n3492 & ~n28098;
  assign n28100 = n3492 & ~n28099;
  assign n28101 = n3485 & ~n28100;
  assign n28102 = n3485 & ~n28101;
  assign n28103 = ~n3374 & ~n28102;
  assign n28104 = ~i_hbusreq3 & ~n28063;
  assign n28105 = ~n9843 & ~n28104;
  assign n28106 = controllable_hmaster2 & ~n28105;
  assign n28107 = ~controllable_hmaster0 & ~n28063;
  assign n28108 = ~n9725 & ~n28107;
  assign n28109 = controllable_hmaster1 & ~n28108;
  assign n28110 = ~controllable_hmaster1 & ~n28063;
  assign n28111 = ~n28109 & ~n28110;
  assign n28112 = ~i_hbusreq3 & ~n28111;
  assign n28113 = ~n26915 & ~n28112;
  assign n28114 = ~controllable_hmaster2 & ~n28113;
  assign n28115 = ~n28106 & ~n28114;
  assign n28116 = controllable_hgrant3 & ~n28115;
  assign n28117 = ~n12749 & ~n28116;
  assign n28118 = controllable_nhgrant0 & ~n28117;
  assign n28119 = ~n12773 & ~n28118;
  assign n28120 = ~n3281 & ~n28119;
  assign n28121 = ~n3281 & ~n28120;
  assign n28122 = n3378 & ~n28121;
  assign n28123 = ~i_hbusreq3 & ~n28081;
  assign n28124 = ~n9843 & ~n28123;
  assign n28125 = controllable_hmaster2 & ~n28124;
  assign n28126 = ~controllable_hmaster0 & ~n28081;
  assign n28127 = ~n9725 & ~n28126;
  assign n28128 = controllable_hmaster1 & ~n28127;
  assign n28129 = ~controllable_hgrant2 & ~n16144;
  assign n28130 = ~n5461 & ~n28129;
  assign n28131 = ~controllable_hmaster0 & ~n28130;
  assign n28132 = ~n28083 & ~n28131;
  assign n28133 = ~controllable_hmaster1 & ~n28132;
  assign n28134 = ~n28128 & ~n28133;
  assign n28135 = ~i_hbusreq3 & ~n28134;
  assign n28136 = ~n26915 & ~n28135;
  assign n28137 = ~controllable_hmaster2 & ~n28136;
  assign n28138 = ~n28125 & ~n28137;
  assign n28139 = controllable_hgrant3 & ~n28138;
  assign n28140 = ~n12803 & ~n28139;
  assign n28141 = controllable_nhgrant0 & ~n28140;
  assign n28142 = ~n12827 & ~n28141;
  assign n28143 = ~n3281 & ~n28142;
  assign n28144 = ~n3281 & ~n28143;
  assign n28145 = ~n3378 & ~n28144;
  assign n28146 = ~n28122 & ~n28145;
  assign n28147 = n3492 & ~n28146;
  assign n28148 = n3492 & ~n28147;
  assign n28149 = n3485 & ~n28148;
  assign n28150 = n3485 & ~n28149;
  assign n28151 = ~n3476 & ~n28150;
  assign n28152 = ~i_hbusreq2 & ~n16183;
  assign n28153 = ~n26969 & ~n28152;
  assign n28154 = ~controllable_hgrant2 & ~n28153;
  assign n28155 = ~n3431 & ~n28154;
  assign n28156 = i_hlock3 & ~n28155;
  assign n28157 = ~i_hbusreq2 & ~n16191;
  assign n28158 = ~n26986 & ~n28157;
  assign n28159 = ~controllable_hgrant2 & ~n28158;
  assign n28160 = ~n3431 & ~n28159;
  assign n28161 = ~i_hlock3 & ~n28160;
  assign n28162 = ~n28156 & ~n28161;
  assign n28163 = ~i_hbusreq3 & ~n28162;
  assign n28164 = ~n27071 & ~n28163;
  assign n28165 = controllable_hmaster2 & ~n28164;
  assign n28166 = ~controllable_hmaster0 & ~n28155;
  assign n28167 = ~n27105 & ~n28166;
  assign n28168 = controllable_hmaster1 & ~n28167;
  assign n28169 = ~controllable_hmaster1 & ~n28155;
  assign n28170 = ~n28168 & ~n28169;
  assign n28171 = i_hlock3 & ~n28170;
  assign n28172 = ~controllable_hmaster0 & ~n28160;
  assign n28173 = ~n27124 & ~n28172;
  assign n28174 = controllable_hmaster1 & ~n28173;
  assign n28175 = ~controllable_hmaster1 & ~n28160;
  assign n28176 = ~n28174 & ~n28175;
  assign n28177 = ~i_hlock3 & ~n28176;
  assign n28178 = ~n28171 & ~n28177;
  assign n28179 = ~i_hbusreq3 & ~n28178;
  assign n28180 = ~n27100 & ~n28179;
  assign n28181 = ~controllable_hmaster2 & ~n28180;
  assign n28182 = ~n28165 & ~n28181;
  assign n28183 = controllable_hgrant3 & ~n28182;
  assign n28184 = ~n12924 & ~n28183;
  assign n28185 = controllable_nhgrant0 & ~n28184;
  assign n28186 = ~n12942 & ~n28185;
  assign n28187 = ~n3281 & ~n28186;
  assign n28188 = ~n3281 & ~n28187;
  assign n28189 = n3378 & ~n28188;
  assign n28190 = ~i_hbusreq2 & ~n16260;
  assign n28191 = ~n26969 & ~n28190;
  assign n28192 = ~controllable_hgrant2 & ~n28191;
  assign n28193 = ~n3859 & ~n28192;
  assign n28194 = i_hlock3 & ~n28193;
  assign n28195 = ~i_hbusreq2 & ~n16269;
  assign n28196 = ~n26986 & ~n28195;
  assign n28197 = ~controllable_hgrant2 & ~n28196;
  assign n28198 = ~n3859 & ~n28197;
  assign n28199 = ~i_hlock3 & ~n28198;
  assign n28200 = ~n28194 & ~n28199;
  assign n28201 = ~i_hbusreq3 & ~n28200;
  assign n28202 = ~n27071 & ~n28201;
  assign n28203 = controllable_hmaster2 & ~n28202;
  assign n28204 = ~controllable_hmaster0 & ~n28193;
  assign n28205 = ~n27105 & ~n28204;
  assign n28206 = controllable_hmaster1 & ~n28205;
  assign n28207 = controllable_hmaster0 & ~n28193;
  assign n28208 = ~i_hbusreq2 & ~n16315;
  assign n28209 = ~n26969 & ~n28208;
  assign n28210 = ~controllable_hgrant2 & ~n28209;
  assign n28211 = ~n5461 & ~n28210;
  assign n28212 = ~controllable_hmaster0 & ~n28211;
  assign n28213 = ~n28207 & ~n28212;
  assign n28214 = ~controllable_hmaster1 & ~n28213;
  assign n28215 = ~n28206 & ~n28214;
  assign n28216 = i_hlock3 & ~n28215;
  assign n28217 = ~controllable_hmaster0 & ~n28198;
  assign n28218 = ~n27124 & ~n28217;
  assign n28219 = controllable_hmaster1 & ~n28218;
  assign n28220 = controllable_hmaster0 & ~n28198;
  assign n28221 = ~i_hbusreq2 & ~n16325;
  assign n28222 = ~n26986 & ~n28221;
  assign n28223 = ~controllable_hgrant2 & ~n28222;
  assign n28224 = ~n5461 & ~n28223;
  assign n28225 = ~controllable_hmaster0 & ~n28224;
  assign n28226 = ~n28220 & ~n28225;
  assign n28227 = ~controllable_hmaster1 & ~n28226;
  assign n28228 = ~n28219 & ~n28227;
  assign n28229 = ~i_hlock3 & ~n28228;
  assign n28230 = ~n28216 & ~n28229;
  assign n28231 = ~i_hbusreq3 & ~n28230;
  assign n28232 = ~n27100 & ~n28231;
  assign n28233 = ~controllable_hmaster2 & ~n28232;
  assign n28234 = ~n28203 & ~n28233;
  assign n28235 = controllable_hgrant3 & ~n28234;
  assign n28236 = ~n13046 & ~n28235;
  assign n28237 = controllable_nhgrant0 & ~n28236;
  assign n28238 = ~n13064 & ~n28237;
  assign n28239 = ~n3281 & ~n28238;
  assign n28240 = ~n3281 & ~n28239;
  assign n28241 = ~n3378 & ~n28240;
  assign n28242 = ~n28189 & ~n28241;
  assign n28243 = n3492 & ~n28242;
  assign n28244 = ~n27622 & ~n28243;
  assign n28245 = n3485 & ~n28244;
  assign n28246 = ~n27621 & ~n28245;
  assign n28247 = n3476 & ~n28246;
  assign n28248 = ~n28151 & ~n28247;
  assign n28249 = n3374 & ~n28248;
  assign n28250 = ~n28103 & ~n28249;
  assign n28251 = n3655 & ~n28250;
  assign n28252 = ~n7694 & ~n28091;
  assign n28253 = controllable_nhgrant0 & ~n28252;
  assign n28254 = ~n7118 & ~n28253;
  assign n28255 = ~n3281 & ~n28254;
  assign n28256 = ~n3281 & ~n28255;
  assign n28257 = ~n3378 & ~n28256;
  assign n28258 = ~n28079 & ~n28257;
  assign n28259 = n3492 & ~n28258;
  assign n28260 = n3492 & ~n28259;
  assign n28261 = n3485 & ~n28260;
  assign n28262 = n3485 & ~n28261;
  assign n28263 = ~n3374 & ~n28262;
  assign n28264 = ~n13090 & ~n28116;
  assign n28265 = controllable_nhgrant0 & ~n28264;
  assign n28266 = ~n12773 & ~n28265;
  assign n28267 = ~n3281 & ~n28266;
  assign n28268 = ~n3281 & ~n28267;
  assign n28269 = n3378 & ~n28268;
  assign n28270 = ~n13118 & ~n28139;
  assign n28271 = controllable_nhgrant0 & ~n28270;
  assign n28272 = ~n12827 & ~n28271;
  assign n28273 = ~n3281 & ~n28272;
  assign n28274 = ~n3281 & ~n28273;
  assign n28275 = ~n3378 & ~n28274;
  assign n28276 = ~n28269 & ~n28275;
  assign n28277 = n3492 & ~n28276;
  assign n28278 = n3492 & ~n28277;
  assign n28279 = n3485 & ~n28278;
  assign n28280 = n3485 & ~n28279;
  assign n28281 = ~n3476 & ~n28280;
  assign n28282 = ~n13153 & ~n28183;
  assign n28283 = controllable_nhgrant0 & ~n28282;
  assign n28284 = ~n12942 & ~n28283;
  assign n28285 = ~n3281 & ~n28284;
  assign n28286 = ~n3281 & ~n28285;
  assign n28287 = n3378 & ~n28286;
  assign n28288 = ~n13230 & ~n28235;
  assign n28289 = controllable_nhgrant0 & ~n28288;
  assign n28290 = ~n13064 & ~n28289;
  assign n28291 = ~n3281 & ~n28290;
  assign n28292 = ~n3281 & ~n28291;
  assign n28293 = ~n3378 & ~n28292;
  assign n28294 = ~n28287 & ~n28293;
  assign n28295 = n3492 & ~n28294;
  assign n28296 = ~n27622 & ~n28295;
  assign n28297 = n3485 & ~n28296;
  assign n28298 = ~n27621 & ~n28297;
  assign n28299 = n3476 & ~n28298;
  assign n28300 = ~n28281 & ~n28299;
  assign n28301 = n3374 & ~n28300;
  assign n28302 = ~n28263 & ~n28301;
  assign n28303 = ~n3655 & ~n28302;
  assign n28304 = ~n28251 & ~n28303;
  assign n28305 = n3652 & ~n28304;
  assign n28306 = ~n7974 & ~n28091;
  assign n28307 = controllable_nhgrant0 & ~n28306;
  assign n28308 = ~n7118 & ~n28307;
  assign n28309 = ~n3281 & ~n28308;
  assign n28310 = ~n3281 & ~n28309;
  assign n28311 = ~n3378 & ~n28310;
  assign n28312 = ~n28079 & ~n28311;
  assign n28313 = n3492 & ~n28312;
  assign n28314 = n3492 & ~n28313;
  assign n28315 = n3485 & ~n28314;
  assign n28316 = n3485 & ~n28315;
  assign n28317 = ~n3374 & ~n28316;
  assign n28318 = ~n13260 & ~n28116;
  assign n28319 = controllable_nhgrant0 & ~n28318;
  assign n28320 = ~n12773 & ~n28319;
  assign n28321 = ~n3281 & ~n28320;
  assign n28322 = ~n3281 & ~n28321;
  assign n28323 = n3378 & ~n28322;
  assign n28324 = ~n13288 & ~n28139;
  assign n28325 = controllable_nhgrant0 & ~n28324;
  assign n28326 = ~n12827 & ~n28325;
  assign n28327 = ~n3281 & ~n28326;
  assign n28328 = ~n3281 & ~n28327;
  assign n28329 = ~n3378 & ~n28328;
  assign n28330 = ~n28323 & ~n28329;
  assign n28331 = n3492 & ~n28330;
  assign n28332 = n3492 & ~n28331;
  assign n28333 = n3485 & ~n28332;
  assign n28334 = n3485 & ~n28333;
  assign n28335 = ~n3476 & ~n28334;
  assign n28336 = ~n13316 & ~n28183;
  assign n28337 = controllable_nhgrant0 & ~n28336;
  assign n28338 = ~n12942 & ~n28337;
  assign n28339 = ~n3281 & ~n28338;
  assign n28340 = ~n3281 & ~n28339;
  assign n28341 = n3378 & ~n28340;
  assign n28342 = ~n13363 & ~n28235;
  assign n28343 = controllable_nhgrant0 & ~n28342;
  assign n28344 = ~n13064 & ~n28343;
  assign n28345 = ~n3281 & ~n28344;
  assign n28346 = ~n3281 & ~n28345;
  assign n28347 = ~n3378 & ~n28346;
  assign n28348 = ~n28341 & ~n28347;
  assign n28349 = n3492 & ~n28348;
  assign n28350 = ~n27622 & ~n28349;
  assign n28351 = n3485 & ~n28350;
  assign n28352 = ~n27621 & ~n28351;
  assign n28353 = n3476 & ~n28352;
  assign n28354 = ~n28335 & ~n28353;
  assign n28355 = n3374 & ~n28354;
  assign n28356 = ~n28317 & ~n28355;
  assign n28357 = n3655 & ~n28356;
  assign n28358 = ~n8133 & ~n28091;
  assign n28359 = controllable_nhgrant0 & ~n28358;
  assign n28360 = ~n7118 & ~n28359;
  assign n28361 = ~n3281 & ~n28360;
  assign n28362 = ~n3281 & ~n28361;
  assign n28363 = ~n3378 & ~n28362;
  assign n28364 = ~n28079 & ~n28363;
  assign n28365 = n3492 & ~n28364;
  assign n28366 = n3492 & ~n28365;
  assign n28367 = n3485 & ~n28366;
  assign n28368 = n3485 & ~n28367;
  assign n28369 = ~n3374 & ~n28368;
  assign n28370 = ~n13391 & ~n28116;
  assign n28371 = controllable_nhgrant0 & ~n28370;
  assign n28372 = ~n12773 & ~n28371;
  assign n28373 = ~n3281 & ~n28372;
  assign n28374 = ~n3281 & ~n28373;
  assign n28375 = n3378 & ~n28374;
  assign n28376 = ~n13419 & ~n28139;
  assign n28377 = controllable_nhgrant0 & ~n28376;
  assign n28378 = ~n12827 & ~n28377;
  assign n28379 = ~n3281 & ~n28378;
  assign n28380 = ~n3281 & ~n28379;
  assign n28381 = ~n3378 & ~n28380;
  assign n28382 = ~n28375 & ~n28381;
  assign n28383 = n3492 & ~n28382;
  assign n28384 = n3492 & ~n28383;
  assign n28385 = n3485 & ~n28384;
  assign n28386 = n3485 & ~n28385;
  assign n28387 = ~n3476 & ~n28386;
  assign n28388 = ~n13447 & ~n28183;
  assign n28389 = controllable_nhgrant0 & ~n28388;
  assign n28390 = ~n12942 & ~n28389;
  assign n28391 = ~n3281 & ~n28390;
  assign n28392 = ~n3281 & ~n28391;
  assign n28393 = n3378 & ~n28392;
  assign n28394 = ~n13494 & ~n28235;
  assign n28395 = controllable_nhgrant0 & ~n28394;
  assign n28396 = ~n13064 & ~n28395;
  assign n28397 = ~n3281 & ~n28396;
  assign n28398 = ~n3281 & ~n28397;
  assign n28399 = ~n3378 & ~n28398;
  assign n28400 = ~n28393 & ~n28399;
  assign n28401 = n3492 & ~n28400;
  assign n28402 = ~n27622 & ~n28401;
  assign n28403 = n3485 & ~n28402;
  assign n28404 = ~n27621 & ~n28403;
  assign n28405 = n3476 & ~n28404;
  assign n28406 = ~n28387 & ~n28405;
  assign n28407 = n3374 & ~n28406;
  assign n28408 = ~n28369 & ~n28407;
  assign n28409 = ~n3655 & ~n28408;
  assign n28410 = ~n28357 & ~n28409;
  assign n28411 = ~n3652 & ~n28410;
  assign n28412 = ~n28305 & ~n28411;
  assign n28413 = n3368 & ~n28412;
  assign n28414 = ~n28061 & ~n28413;
  assign n28415 = n3362 & ~n28414;
  assign n28416 = n3492 & ~n27770;
  assign n28417 = ~n3631 & ~n28416;
  assign n28418 = n3485 & ~n28417;
  assign n28419 = ~n3630 & ~n28418;
  assign n28420 = ~n3476 & ~n28419;
  assign n28421 = n3492 & ~n27386;
  assign n28422 = ~n26200 & ~n28421;
  assign n28423 = ~n3485 & ~n28422;
  assign n28424 = ~n27779 & ~n28416;
  assign n28425 = n3485 & ~n28424;
  assign n28426 = ~n28423 & ~n28425;
  assign n28427 = n3476 & ~n28426;
  assign n28428 = ~n28420 & ~n28427;
  assign n28429 = ~n3374 & ~n28428;
  assign n28430 = n3492 & ~n27822;
  assign n28431 = ~n3631 & ~n28430;
  assign n28432 = n3485 & ~n28431;
  assign n28433 = ~n3630 & ~n28432;
  assign n28434 = ~n3476 & ~n28433;
  assign n28435 = n3492 & ~n27870;
  assign n28436 = ~n27779 & ~n28435;
  assign n28437 = n3485 & ~n28436;
  assign n28438 = ~n28423 & ~n28437;
  assign n28439 = n3476 & ~n28438;
  assign n28440 = ~n28434 & ~n28439;
  assign n28441 = n3374 & ~n28440;
  assign n28442 = ~n28429 & ~n28441;
  assign n28443 = n3655 & ~n28442;
  assign n28444 = n3492 & ~n27886;
  assign n28445 = ~n3631 & ~n28444;
  assign n28446 = n3485 & ~n28445;
  assign n28447 = ~n3630 & ~n28446;
  assign n28448 = ~n3476 & ~n28447;
  assign n28449 = ~n26297 & ~n28421;
  assign n28450 = ~n3485 & ~n28449;
  assign n28451 = ~n27779 & ~n28444;
  assign n28452 = n3485 & ~n28451;
  assign n28453 = ~n28450 & ~n28452;
  assign n28454 = n3476 & ~n28453;
  assign n28455 = ~n28448 & ~n28454;
  assign n28456 = ~n3374 & ~n28455;
  assign n28457 = n3492 & ~n27910;
  assign n28458 = ~n3631 & ~n28457;
  assign n28459 = n3485 & ~n28458;
  assign n28460 = ~n3630 & ~n28459;
  assign n28461 = ~n3476 & ~n28460;
  assign n28462 = n3492 & ~n27928;
  assign n28463 = ~n27779 & ~n28462;
  assign n28464 = n3485 & ~n28463;
  assign n28465 = ~n28450 & ~n28464;
  assign n28466 = n3476 & ~n28465;
  assign n28467 = ~n28461 & ~n28466;
  assign n28468 = n3374 & ~n28467;
  assign n28469 = ~n28456 & ~n28468;
  assign n28470 = ~n3655 & ~n28469;
  assign n28471 = ~n28443 & ~n28470;
  assign n28472 = n3652 & ~n28471;
  assign n28473 = n3492 & ~n27946;
  assign n28474 = ~n3631 & ~n28473;
  assign n28475 = n3485 & ~n28474;
  assign n28476 = ~n3630 & ~n28475;
  assign n28477 = ~n3476 & ~n28476;
  assign n28478 = ~n26396 & ~n28421;
  assign n28479 = ~n3485 & ~n28478;
  assign n28480 = ~n27779 & ~n28473;
  assign n28481 = n3485 & ~n28480;
  assign n28482 = ~n28479 & ~n28481;
  assign n28483 = n3476 & ~n28482;
  assign n28484 = ~n28477 & ~n28483;
  assign n28485 = ~n3374 & ~n28484;
  assign n28486 = n3492 & ~n27970;
  assign n28487 = ~n3631 & ~n28486;
  assign n28488 = n3485 & ~n28487;
  assign n28489 = ~n3630 & ~n28488;
  assign n28490 = ~n3476 & ~n28489;
  assign n28491 = n3492 & ~n27988;
  assign n28492 = ~n27779 & ~n28491;
  assign n28493 = n3485 & ~n28492;
  assign n28494 = ~n28479 & ~n28493;
  assign n28495 = n3476 & ~n28494;
  assign n28496 = ~n28490 & ~n28495;
  assign n28497 = n3374 & ~n28496;
  assign n28498 = ~n28485 & ~n28497;
  assign n28499 = n3655 & ~n28498;
  assign n28500 = n3492 & ~n28004;
  assign n28501 = ~n3631 & ~n28500;
  assign n28502 = n3485 & ~n28501;
  assign n28503 = ~n3630 & ~n28502;
  assign n28504 = ~n3476 & ~n28503;
  assign n28505 = ~n26437 & ~n28421;
  assign n28506 = ~n3485 & ~n28505;
  assign n28507 = ~n27779 & ~n28500;
  assign n28508 = n3485 & ~n28507;
  assign n28509 = ~n28506 & ~n28508;
  assign n28510 = n3476 & ~n28509;
  assign n28511 = ~n28504 & ~n28510;
  assign n28512 = ~n3374 & ~n28511;
  assign n28513 = n3492 & ~n28028;
  assign n28514 = ~n3631 & ~n28513;
  assign n28515 = n3485 & ~n28514;
  assign n28516 = ~n3630 & ~n28515;
  assign n28517 = ~n3476 & ~n28516;
  assign n28518 = n3492 & ~n28046;
  assign n28519 = ~n27779 & ~n28518;
  assign n28520 = n3485 & ~n28519;
  assign n28521 = ~n28506 & ~n28520;
  assign n28522 = n3476 & ~n28521;
  assign n28523 = ~n28517 & ~n28522;
  assign n28524 = n3374 & ~n28523;
  assign n28525 = ~n28512 & ~n28524;
  assign n28526 = ~n3655 & ~n28525;
  assign n28527 = ~n28499 & ~n28526;
  assign n28528 = ~n3652 & ~n28527;
  assign n28529 = ~n28472 & ~n28528;
  assign n28530 = ~n3368 & ~n28529;
  assign n28531 = n3492 & ~n28096;
  assign n28532 = n3492 & ~n28531;
  assign n28533 = n3485 & ~n28532;
  assign n28534 = n3485 & ~n28533;
  assign n28535 = ~n3476 & ~n28534;
  assign n28536 = ~n8525 & ~n28533;
  assign n28537 = n3476 & ~n28536;
  assign n28538 = ~n28535 & ~n28537;
  assign n28539 = ~n3374 & ~n28538;
  assign n28540 = n3492 & ~n28144;
  assign n28541 = n3492 & ~n28540;
  assign n28542 = n3485 & ~n28541;
  assign n28543 = n3485 & ~n28542;
  assign n28544 = ~n3476 & ~n28543;
  assign n28545 = n3492 & ~n27353;
  assign n28546 = ~n26477 & ~n28545;
  assign n28547 = ~n3485 & ~n28546;
  assign n28548 = n3492 & ~n28240;
  assign n28549 = ~n27622 & ~n28548;
  assign n28550 = n3485 & ~n28549;
  assign n28551 = ~n28547 & ~n28550;
  assign n28552 = n3476 & ~n28551;
  assign n28553 = ~n28544 & ~n28552;
  assign n28554 = n3374 & ~n28553;
  assign n28555 = ~n28539 & ~n28554;
  assign n28556 = n3655 & ~n28555;
  assign n28557 = n3492 & ~n28256;
  assign n28558 = n3492 & ~n28557;
  assign n28559 = n3485 & ~n28558;
  assign n28560 = n3485 & ~n28559;
  assign n28561 = ~n3476 & ~n28560;
  assign n28562 = ~n8525 & ~n28559;
  assign n28563 = n3476 & ~n28562;
  assign n28564 = ~n28561 & ~n28563;
  assign n28565 = ~n3374 & ~n28564;
  assign n28566 = n3492 & ~n28274;
  assign n28567 = n3492 & ~n28566;
  assign n28568 = n3485 & ~n28567;
  assign n28569 = n3485 & ~n28568;
  assign n28570 = ~n3476 & ~n28569;
  assign n28571 = ~n26504 & ~n28545;
  assign n28572 = ~n3485 & ~n28571;
  assign n28573 = n3492 & ~n28292;
  assign n28574 = ~n27622 & ~n28573;
  assign n28575 = n3485 & ~n28574;
  assign n28576 = ~n28572 & ~n28575;
  assign n28577 = n3476 & ~n28576;
  assign n28578 = ~n28570 & ~n28577;
  assign n28579 = n3374 & ~n28578;
  assign n28580 = ~n28565 & ~n28579;
  assign n28581 = ~n3655 & ~n28580;
  assign n28582 = ~n28556 & ~n28581;
  assign n28583 = n3652 & ~n28582;
  assign n28584 = n3492 & ~n28310;
  assign n28585 = n3492 & ~n28584;
  assign n28586 = n3485 & ~n28585;
  assign n28587 = n3485 & ~n28586;
  assign n28588 = ~n3476 & ~n28587;
  assign n28589 = ~n8525 & ~n28586;
  assign n28590 = n3476 & ~n28589;
  assign n28591 = ~n28588 & ~n28590;
  assign n28592 = ~n3374 & ~n28591;
  assign n28593 = n3492 & ~n28328;
  assign n28594 = n3492 & ~n28593;
  assign n28595 = n3485 & ~n28594;
  assign n28596 = n3485 & ~n28595;
  assign n28597 = ~n3476 & ~n28596;
  assign n28598 = ~n26533 & ~n28545;
  assign n28599 = ~n3485 & ~n28598;
  assign n28600 = n3492 & ~n28346;
  assign n28601 = ~n27622 & ~n28600;
  assign n28602 = n3485 & ~n28601;
  assign n28603 = ~n28599 & ~n28602;
  assign n28604 = n3476 & ~n28603;
  assign n28605 = ~n28597 & ~n28604;
  assign n28606 = n3374 & ~n28605;
  assign n28607 = ~n28592 & ~n28606;
  assign n28608 = n3655 & ~n28607;
  assign n28609 = n3492 & ~n28362;
  assign n28610 = n3492 & ~n28609;
  assign n28611 = n3485 & ~n28610;
  assign n28612 = n3485 & ~n28611;
  assign n28613 = ~n3476 & ~n28612;
  assign n28614 = ~n8525 & ~n28611;
  assign n28615 = n3476 & ~n28614;
  assign n28616 = ~n28613 & ~n28615;
  assign n28617 = ~n3374 & ~n28616;
  assign n28618 = n3492 & ~n28380;
  assign n28619 = n3492 & ~n28618;
  assign n28620 = n3485 & ~n28619;
  assign n28621 = n3485 & ~n28620;
  assign n28622 = ~n3476 & ~n28621;
  assign n28623 = ~n26560 & ~n28545;
  assign n28624 = ~n3485 & ~n28623;
  assign n28625 = n3492 & ~n28398;
  assign n28626 = ~n27622 & ~n28625;
  assign n28627 = n3485 & ~n28626;
  assign n28628 = ~n28624 & ~n28627;
  assign n28629 = n3476 & ~n28628;
  assign n28630 = ~n28622 & ~n28629;
  assign n28631 = n3374 & ~n28630;
  assign n28632 = ~n28617 & ~n28631;
  assign n28633 = ~n3655 & ~n28632;
  assign n28634 = ~n28608 & ~n28633;
  assign n28635 = ~n3652 & ~n28634;
  assign n28636 = ~n28583 & ~n28635;
  assign n28637 = n3368 & ~n28636;
  assign n28638 = ~n28530 & ~n28637;
  assign n28639 = ~n3362 & ~n28638;
  assign n28640 = ~n28415 & ~n28639;
  assign n28641 = n3359 & ~n28640;
  assign n28642 = ~n26580 & ~n28425;
  assign n28643 = n3476 & ~n28642;
  assign n28644 = ~n28420 & ~n28643;
  assign n28645 = ~n3374 & ~n28644;
  assign n28646 = ~n26580 & ~n28437;
  assign n28647 = n3476 & ~n28646;
  assign n28648 = ~n28434 & ~n28647;
  assign n28649 = n3374 & ~n28648;
  assign n28650 = ~n28645 & ~n28649;
  assign n28651 = n3655 & ~n28650;
  assign n28652 = ~n26591 & ~n28452;
  assign n28653 = n3476 & ~n28652;
  assign n28654 = ~n28448 & ~n28653;
  assign n28655 = ~n3374 & ~n28654;
  assign n28656 = ~n26591 & ~n28464;
  assign n28657 = n3476 & ~n28656;
  assign n28658 = ~n28461 & ~n28657;
  assign n28659 = n3374 & ~n28658;
  assign n28660 = ~n28655 & ~n28659;
  assign n28661 = ~n3655 & ~n28660;
  assign n28662 = ~n28651 & ~n28661;
  assign n28663 = n3652 & ~n28662;
  assign n28664 = ~n26604 & ~n28481;
  assign n28665 = n3476 & ~n28664;
  assign n28666 = ~n28477 & ~n28665;
  assign n28667 = ~n3374 & ~n28666;
  assign n28668 = ~n26604 & ~n28493;
  assign n28669 = n3476 & ~n28668;
  assign n28670 = ~n28490 & ~n28669;
  assign n28671 = n3374 & ~n28670;
  assign n28672 = ~n28667 & ~n28671;
  assign n28673 = n3655 & ~n28672;
  assign n28674 = ~n26615 & ~n28508;
  assign n28675 = n3476 & ~n28674;
  assign n28676 = ~n28504 & ~n28675;
  assign n28677 = ~n3374 & ~n28676;
  assign n28678 = ~n26615 & ~n28520;
  assign n28679 = n3476 & ~n28678;
  assign n28680 = ~n28517 & ~n28679;
  assign n28681 = n3374 & ~n28680;
  assign n28682 = ~n28677 & ~n28681;
  assign n28683 = ~n3655 & ~n28682;
  assign n28684 = ~n28673 & ~n28683;
  assign n28685 = ~n3652 & ~n28684;
  assign n28686 = ~n28663 & ~n28685;
  assign n28687 = ~n3368 & ~n28686;
  assign n28688 = ~n8689 & ~n28533;
  assign n28689 = n3476 & ~n28688;
  assign n28690 = ~n28535 & ~n28689;
  assign n28691 = ~n3374 & ~n28690;
  assign n28692 = ~n26634 & ~n28550;
  assign n28693 = n3476 & ~n28692;
  assign n28694 = ~n28544 & ~n28693;
  assign n28695 = n3374 & ~n28694;
  assign n28696 = ~n28691 & ~n28695;
  assign n28697 = n3655 & ~n28696;
  assign n28698 = ~n8689 & ~n28559;
  assign n28699 = n3476 & ~n28698;
  assign n28700 = ~n28561 & ~n28699;
  assign n28701 = ~n3374 & ~n28700;
  assign n28702 = ~n26645 & ~n28575;
  assign n28703 = n3476 & ~n28702;
  assign n28704 = ~n28570 & ~n28703;
  assign n28705 = n3374 & ~n28704;
  assign n28706 = ~n28701 & ~n28705;
  assign n28707 = ~n3655 & ~n28706;
  assign n28708 = ~n28697 & ~n28707;
  assign n28709 = n3652 & ~n28708;
  assign n28710 = ~n8689 & ~n28586;
  assign n28711 = n3476 & ~n28710;
  assign n28712 = ~n28588 & ~n28711;
  assign n28713 = ~n3374 & ~n28712;
  assign n28714 = ~n26658 & ~n28602;
  assign n28715 = n3476 & ~n28714;
  assign n28716 = ~n28597 & ~n28715;
  assign n28717 = n3374 & ~n28716;
  assign n28718 = ~n28713 & ~n28717;
  assign n28719 = n3655 & ~n28718;
  assign n28720 = ~n8689 & ~n28611;
  assign n28721 = n3476 & ~n28720;
  assign n28722 = ~n28613 & ~n28721;
  assign n28723 = ~n3374 & ~n28722;
  assign n28724 = ~n26669 & ~n28627;
  assign n28725 = n3476 & ~n28724;
  assign n28726 = ~n28622 & ~n28725;
  assign n28727 = n3374 & ~n28726;
  assign n28728 = ~n28723 & ~n28727;
  assign n28729 = ~n3655 & ~n28728;
  assign n28730 = ~n28719 & ~n28729;
  assign n28731 = ~n3652 & ~n28730;
  assign n28732 = ~n28709 & ~n28731;
  assign n28733 = n3368 & ~n28732;
  assign n28734 = ~n28687 & ~n28733;
  assign n28735 = n3362 & ~n28734;
  assign n28736 = n3378 & ~n27770;
  assign n28737 = ~n26690 & ~n28736;
  assign n28738 = n3492 & ~n28737;
  assign n28739 = ~n3631 & ~n28738;
  assign n28740 = n3485 & ~n28739;
  assign n28741 = ~n3630 & ~n28740;
  assign n28742 = ~n3476 & ~n28741;
  assign n28743 = ~n26200 & ~n28738;
  assign n28744 = n3485 & ~n28743;
  assign n28745 = ~n26580 & ~n28744;
  assign n28746 = n3476 & ~n28745;
  assign n28747 = ~n28742 & ~n28746;
  assign n28748 = ~n3374 & ~n28747;
  assign n28749 = n3378 & ~n27822;
  assign n28750 = ~n26711 & ~n28749;
  assign n28751 = n3492 & ~n28750;
  assign n28752 = ~n3631 & ~n28751;
  assign n28753 = n3485 & ~n28752;
  assign n28754 = ~n3630 & ~n28753;
  assign n28755 = ~n3476 & ~n28754;
  assign n28756 = n3378 & ~n27870;
  assign n28757 = ~n26726 & ~n28756;
  assign n28758 = n3492 & ~n28757;
  assign n28759 = ~n26200 & ~n28758;
  assign n28760 = n3485 & ~n28759;
  assign n28761 = ~n26580 & ~n28760;
  assign n28762 = n3476 & ~n28761;
  assign n28763 = ~n28755 & ~n28762;
  assign n28764 = n3374 & ~n28763;
  assign n28765 = ~n28748 & ~n28764;
  assign n28766 = n3655 & ~n28765;
  assign n28767 = n3378 & ~n27886;
  assign n28768 = ~n26743 & ~n28767;
  assign n28769 = n3492 & ~n28768;
  assign n28770 = ~n3631 & ~n28769;
  assign n28771 = n3485 & ~n28770;
  assign n28772 = ~n3630 & ~n28771;
  assign n28773 = ~n3476 & ~n28772;
  assign n28774 = ~n26297 & ~n28769;
  assign n28775 = n3485 & ~n28774;
  assign n28776 = ~n26591 & ~n28775;
  assign n28777 = n3476 & ~n28776;
  assign n28778 = ~n28773 & ~n28777;
  assign n28779 = ~n3374 & ~n28778;
  assign n28780 = n3378 & ~n27910;
  assign n28781 = ~n26762 & ~n28780;
  assign n28782 = n3492 & ~n28781;
  assign n28783 = ~n3631 & ~n28782;
  assign n28784 = n3485 & ~n28783;
  assign n28785 = ~n3630 & ~n28784;
  assign n28786 = ~n3476 & ~n28785;
  assign n28787 = n3378 & ~n27928;
  assign n28788 = ~n26775 & ~n28787;
  assign n28789 = n3492 & ~n28788;
  assign n28790 = ~n26297 & ~n28789;
  assign n28791 = n3485 & ~n28790;
  assign n28792 = ~n26591 & ~n28791;
  assign n28793 = n3476 & ~n28792;
  assign n28794 = ~n28786 & ~n28793;
  assign n28795 = n3374 & ~n28794;
  assign n28796 = ~n28779 & ~n28795;
  assign n28797 = ~n3655 & ~n28796;
  assign n28798 = ~n28766 & ~n28797;
  assign n28799 = n3652 & ~n28798;
  assign n28800 = n3378 & ~n27946;
  assign n28801 = ~n26794 & ~n28800;
  assign n28802 = n3492 & ~n28801;
  assign n28803 = ~n3631 & ~n28802;
  assign n28804 = n3485 & ~n28803;
  assign n28805 = ~n3630 & ~n28804;
  assign n28806 = ~n3476 & ~n28805;
  assign n28807 = ~n26396 & ~n28802;
  assign n28808 = n3485 & ~n28807;
  assign n28809 = ~n26604 & ~n28808;
  assign n28810 = n3476 & ~n28809;
  assign n28811 = ~n28806 & ~n28810;
  assign n28812 = ~n3374 & ~n28811;
  assign n28813 = n3378 & ~n27970;
  assign n28814 = ~n26813 & ~n28813;
  assign n28815 = n3492 & ~n28814;
  assign n28816 = ~n3631 & ~n28815;
  assign n28817 = n3485 & ~n28816;
  assign n28818 = ~n3630 & ~n28817;
  assign n28819 = ~n3476 & ~n28818;
  assign n28820 = n3378 & ~n27988;
  assign n28821 = ~n26826 & ~n28820;
  assign n28822 = n3492 & ~n28821;
  assign n28823 = ~n26396 & ~n28822;
  assign n28824 = n3485 & ~n28823;
  assign n28825 = ~n26604 & ~n28824;
  assign n28826 = n3476 & ~n28825;
  assign n28827 = ~n28819 & ~n28826;
  assign n28828 = n3374 & ~n28827;
  assign n28829 = ~n28812 & ~n28828;
  assign n28830 = n3655 & ~n28829;
  assign n28831 = n3378 & ~n28004;
  assign n28832 = ~n26843 & ~n28831;
  assign n28833 = n3492 & ~n28832;
  assign n28834 = ~n3631 & ~n28833;
  assign n28835 = n3485 & ~n28834;
  assign n28836 = ~n3630 & ~n28835;
  assign n28837 = ~n3476 & ~n28836;
  assign n28838 = ~n26437 & ~n28833;
  assign n28839 = n3485 & ~n28838;
  assign n28840 = ~n26615 & ~n28839;
  assign n28841 = n3476 & ~n28840;
  assign n28842 = ~n28837 & ~n28841;
  assign n28843 = ~n3374 & ~n28842;
  assign n28844 = n3378 & ~n28028;
  assign n28845 = ~n26862 & ~n28844;
  assign n28846 = n3492 & ~n28845;
  assign n28847 = ~n3631 & ~n28846;
  assign n28848 = n3485 & ~n28847;
  assign n28849 = ~n3630 & ~n28848;
  assign n28850 = ~n3476 & ~n28849;
  assign n28851 = n3378 & ~n28046;
  assign n28852 = ~n26875 & ~n28851;
  assign n28853 = n3492 & ~n28852;
  assign n28854 = ~n26437 & ~n28853;
  assign n28855 = n3485 & ~n28854;
  assign n28856 = ~n26615 & ~n28855;
  assign n28857 = n3476 & ~n28856;
  assign n28858 = ~n28850 & ~n28857;
  assign n28859 = n3374 & ~n28858;
  assign n28860 = ~n28843 & ~n28859;
  assign n28861 = ~n3655 & ~n28860;
  assign n28862 = ~n28830 & ~n28861;
  assign n28863 = ~n3652 & ~n28862;
  assign n28864 = ~n28799 & ~n28863;
  assign n28865 = ~n3368 & ~n28864;
  assign n28866 = n3378 & ~n28096;
  assign n28867 = ~n26897 & ~n28866;
  assign n28868 = n3492 & ~n28867;
  assign n28869 = n3492 & ~n28868;
  assign n28870 = n3485 & ~n28869;
  assign n28871 = n3485 & ~n28870;
  assign n28872 = ~n3476 & ~n28871;
  assign n28873 = ~n8523 & ~n28868;
  assign n28874 = n3485 & ~n28873;
  assign n28875 = ~n8689 & ~n28874;
  assign n28876 = n3476 & ~n28875;
  assign n28877 = ~n28872 & ~n28876;
  assign n28878 = ~n3374 & ~n28877;
  assign n28879 = n3378 & ~n28144;
  assign n28880 = ~n26931 & ~n28879;
  assign n28881 = n3492 & ~n28880;
  assign n28882 = n3492 & ~n28881;
  assign n28883 = n3485 & ~n28882;
  assign n28884 = n3485 & ~n28883;
  assign n28885 = ~n3476 & ~n28884;
  assign n28886 = ~n13822 & ~n28235;
  assign n28887 = controllable_nhgrant0 & ~n28886;
  assign n28888 = ~n13845 & ~n28887;
  assign n28889 = ~n3281 & ~n28888;
  assign n28890 = ~n3281 & ~n28889;
  assign n28891 = n3378 & ~n28890;
  assign n28892 = ~n27144 & ~n28891;
  assign n28893 = n3492 & ~n28892;
  assign n28894 = ~n26477 & ~n28893;
  assign n28895 = n3485 & ~n28894;
  assign n28896 = ~n26634 & ~n28895;
  assign n28897 = n3476 & ~n28896;
  assign n28898 = ~n28885 & ~n28897;
  assign n28899 = n3374 & ~n28898;
  assign n28900 = ~n28878 & ~n28899;
  assign n28901 = n3655 & ~n28900;
  assign n28902 = n3378 & ~n28256;
  assign n28903 = ~n27161 & ~n28902;
  assign n28904 = n3492 & ~n28903;
  assign n28905 = n3492 & ~n28904;
  assign n28906 = n3485 & ~n28905;
  assign n28907 = n3485 & ~n28906;
  assign n28908 = ~n3476 & ~n28907;
  assign n28909 = ~n8523 & ~n28904;
  assign n28910 = n3485 & ~n28909;
  assign n28911 = ~n8689 & ~n28910;
  assign n28912 = n3476 & ~n28911;
  assign n28913 = ~n28908 & ~n28912;
  assign n28914 = ~n3374 & ~n28913;
  assign n28915 = n3378 & ~n28274;
  assign n28916 = ~n27180 & ~n28915;
  assign n28917 = n3492 & ~n28916;
  assign n28918 = n3492 & ~n28917;
  assign n28919 = n3485 & ~n28918;
  assign n28920 = n3485 & ~n28919;
  assign n28921 = ~n3476 & ~n28920;
  assign n28922 = ~n13932 & ~n28235;
  assign n28923 = controllable_nhgrant0 & ~n28922;
  assign n28924 = ~n13845 & ~n28923;
  assign n28925 = ~n3281 & ~n28924;
  assign n28926 = ~n3281 & ~n28925;
  assign n28927 = n3378 & ~n28926;
  assign n28928 = ~n27198 & ~n28927;
  assign n28929 = n3492 & ~n28928;
  assign n28930 = ~n26504 & ~n28929;
  assign n28931 = n3485 & ~n28930;
  assign n28932 = ~n26645 & ~n28931;
  assign n28933 = n3476 & ~n28932;
  assign n28934 = ~n28921 & ~n28933;
  assign n28935 = n3374 & ~n28934;
  assign n28936 = ~n28914 & ~n28935;
  assign n28937 = ~n3655 & ~n28936;
  assign n28938 = ~n28901 & ~n28937;
  assign n28939 = n3652 & ~n28938;
  assign n28940 = n3378 & ~n28310;
  assign n28941 = ~n27217 & ~n28940;
  assign n28942 = n3492 & ~n28941;
  assign n28943 = n3492 & ~n28942;
  assign n28944 = n3485 & ~n28943;
  assign n28945 = n3485 & ~n28944;
  assign n28946 = ~n3476 & ~n28945;
  assign n28947 = ~n8523 & ~n28942;
  assign n28948 = n3485 & ~n28947;
  assign n28949 = ~n8689 & ~n28948;
  assign n28950 = n3476 & ~n28949;
  assign n28951 = ~n28946 & ~n28950;
  assign n28952 = ~n3374 & ~n28951;
  assign n28953 = n3378 & ~n28328;
  assign n28954 = ~n27236 & ~n28953;
  assign n28955 = n3492 & ~n28954;
  assign n28956 = n3492 & ~n28955;
  assign n28957 = n3485 & ~n28956;
  assign n28958 = n3485 & ~n28957;
  assign n28959 = ~n3476 & ~n28958;
  assign n28960 = ~n13996 & ~n28235;
  assign n28961 = controllable_nhgrant0 & ~n28960;
  assign n28962 = ~n13845 & ~n28961;
  assign n28963 = ~n3281 & ~n28962;
  assign n28964 = ~n3281 & ~n28963;
  assign n28965 = n3378 & ~n28964;
  assign n28966 = ~n27254 & ~n28965;
  assign n28967 = n3492 & ~n28966;
  assign n28968 = ~n26533 & ~n28967;
  assign n28969 = n3485 & ~n28968;
  assign n28970 = ~n26658 & ~n28969;
  assign n28971 = n3476 & ~n28970;
  assign n28972 = ~n28959 & ~n28971;
  assign n28973 = n3374 & ~n28972;
  assign n28974 = ~n28952 & ~n28973;
  assign n28975 = n3655 & ~n28974;
  assign n28976 = n3378 & ~n28362;
  assign n28977 = ~n27271 & ~n28976;
  assign n28978 = n3492 & ~n28977;
  assign n28979 = n3492 & ~n28978;
  assign n28980 = n3485 & ~n28979;
  assign n28981 = n3485 & ~n28980;
  assign n28982 = ~n3476 & ~n28981;
  assign n28983 = ~n8523 & ~n28978;
  assign n28984 = n3485 & ~n28983;
  assign n28985 = ~n8689 & ~n28984;
  assign n28986 = n3476 & ~n28985;
  assign n28987 = ~n28982 & ~n28986;
  assign n28988 = ~n3374 & ~n28987;
  assign n28989 = n3378 & ~n28380;
  assign n28990 = ~n27290 & ~n28989;
  assign n28991 = n3492 & ~n28990;
  assign n28992 = n3492 & ~n28991;
  assign n28993 = n3485 & ~n28992;
  assign n28994 = n3485 & ~n28993;
  assign n28995 = ~n3476 & ~n28994;
  assign n28996 = ~n14058 & ~n28235;
  assign n28997 = controllable_nhgrant0 & ~n28996;
  assign n28998 = ~n13845 & ~n28997;
  assign n28999 = ~n3281 & ~n28998;
  assign n29000 = ~n3281 & ~n28999;
  assign n29001 = n3378 & ~n29000;
  assign n29002 = ~n27308 & ~n29001;
  assign n29003 = n3492 & ~n29002;
  assign n29004 = ~n26560 & ~n29003;
  assign n29005 = n3485 & ~n29004;
  assign n29006 = ~n26669 & ~n29005;
  assign n29007 = n3476 & ~n29006;
  assign n29008 = ~n28995 & ~n29007;
  assign n29009 = n3374 & ~n29008;
  assign n29010 = ~n28988 & ~n29009;
  assign n29011 = ~n3655 & ~n29010;
  assign n29012 = ~n28975 & ~n29011;
  assign n29013 = ~n3652 & ~n29012;
  assign n29014 = ~n28939 & ~n29013;
  assign n29015 = n3368 & ~n29014;
  assign n29016 = ~n28865 & ~n29015;
  assign n29017 = ~n3362 & ~n29016;
  assign n29018 = ~n28735 & ~n29017;
  assign n29019 = ~n3359 & ~n29018;
  assign n29020 = ~n28641 & ~n29019;
  assign n29021 = ~n3356 & ~n29020;
  assign n29022 = ~n27755 & ~n29021;
  assign n29023 = ~n3345 & ~n29022;
  assign n29024 = controllable_hgrant3 & ~n14163;
  assign n29025 = ~n14152 & ~n29024;
  assign n29026 = controllable_nhgrant0 & ~n29025;
  assign n29027 = ~n14166 & ~n29026;
  assign n29028 = ~n3281 & ~n29027;
  assign n29029 = ~n3281 & ~n29028;
  assign n29030 = n3378 & ~n29029;
  assign n29031 = controllable_hgrant3 & ~n14177;
  assign n29032 = ~n14174 & ~n29031;
  assign n29033 = controllable_nhgrant0 & ~n29032;
  assign n29034 = ~n14180 & ~n29033;
  assign n29035 = ~n3281 & ~n29034;
  assign n29036 = ~n3950 & ~n29035;
  assign n29037 = ~n3378 & ~n29036;
  assign n29038 = ~n29030 & ~n29037;
  assign n29039 = n3492 & ~n29038;
  assign n29040 = ~n3493 & ~n29039;
  assign n29041 = n3485 & ~n29040;
  assign n29042 = ~n3486 & ~n29041;
  assign n29043 = ~n3476 & ~n29042;
  assign n29044 = ~n14218 & ~n29024;
  assign n29045 = controllable_nhgrant0 & ~n29044;
  assign n29046 = ~n14166 & ~n29045;
  assign n29047 = ~n3281 & ~n29046;
  assign n29048 = ~n3281 & ~n29047;
  assign n29049 = n3378 & ~n29048;
  assign n29050 = ~n14265 & ~n29031;
  assign n29051 = controllable_nhgrant0 & ~n29050;
  assign n29052 = ~n14180 & ~n29051;
  assign n29053 = ~n3281 & ~n29052;
  assign n29054 = ~n4089 & ~n29053;
  assign n29055 = ~n3378 & ~n29054;
  assign n29056 = ~n29049 & ~n29055;
  assign n29057 = n3492 & ~n29056;
  assign n29058 = ~n3493 & ~n29057;
  assign n29059 = n3485 & ~n29058;
  assign n29060 = ~n3486 & ~n29059;
  assign n29061 = n3476 & ~n29060;
  assign n29062 = ~n29043 & ~n29061;
  assign n29063 = n3374 & ~n29062;
  assign n29064 = ~n14130 & ~n29063;
  assign n29065 = n3655 & ~n29064;
  assign n29066 = ~n14293 & ~n29024;
  assign n29067 = controllable_nhgrant0 & ~n29066;
  assign n29068 = ~n14166 & ~n29067;
  assign n29069 = ~n3281 & ~n29068;
  assign n29070 = ~n3281 & ~n29069;
  assign n29071 = n3378 & ~n29070;
  assign n29072 = ~n14301 & ~n29031;
  assign n29073 = controllable_nhgrant0 & ~n29072;
  assign n29074 = ~n14180 & ~n29073;
  assign n29075 = ~n3281 & ~n29074;
  assign n29076 = ~n3950 & ~n29075;
  assign n29077 = ~n3378 & ~n29076;
  assign n29078 = ~n29071 & ~n29077;
  assign n29079 = n3492 & ~n29078;
  assign n29080 = ~n3493 & ~n29079;
  assign n29081 = n3485 & ~n29080;
  assign n29082 = ~n3486 & ~n29081;
  assign n29083 = ~n3476 & ~n29082;
  assign n29084 = ~n14329 & ~n29024;
  assign n29085 = controllable_nhgrant0 & ~n29084;
  assign n29086 = ~n14166 & ~n29085;
  assign n29087 = ~n3281 & ~n29086;
  assign n29088 = ~n3281 & ~n29087;
  assign n29089 = n3378 & ~n29088;
  assign n29090 = ~n14351 & ~n29031;
  assign n29091 = controllable_nhgrant0 & ~n29090;
  assign n29092 = ~n14180 & ~n29091;
  assign n29093 = ~n3281 & ~n29092;
  assign n29094 = ~n4089 & ~n29093;
  assign n29095 = ~n3378 & ~n29094;
  assign n29096 = ~n29089 & ~n29095;
  assign n29097 = n3492 & ~n29096;
  assign n29098 = ~n3493 & ~n29097;
  assign n29099 = n3485 & ~n29098;
  assign n29100 = ~n3486 & ~n29099;
  assign n29101 = n3476 & ~n29100;
  assign n29102 = ~n29083 & ~n29101;
  assign n29103 = n3374 & ~n29102;
  assign n29104 = ~n14130 & ~n29103;
  assign n29105 = ~n3655 & ~n29104;
  assign n29106 = ~n29065 & ~n29105;
  assign n29107 = n3652 & ~n29106;
  assign n29108 = ~n14451 & ~n29024;
  assign n29109 = controllable_nhgrant0 & ~n29108;
  assign n29110 = ~n14166 & ~n29109;
  assign n29111 = ~n3281 & ~n29110;
  assign n29112 = ~n3281 & ~n29111;
  assign n29113 = n3378 & ~n29112;
  assign n29114 = ~n14472 & ~n29031;
  assign n29115 = controllable_nhgrant0 & ~n29114;
  assign n29116 = ~n14180 & ~n29115;
  assign n29117 = ~n3281 & ~n29116;
  assign n29118 = ~n3950 & ~n29117;
  assign n29119 = ~n3378 & ~n29118;
  assign n29120 = ~n29113 & ~n29119;
  assign n29121 = n3492 & ~n29120;
  assign n29122 = ~n3493 & ~n29121;
  assign n29123 = n3485 & ~n29122;
  assign n29124 = ~n3486 & ~n29123;
  assign n29125 = ~n3476 & ~n29124;
  assign n29126 = ~n14530 & ~n29024;
  assign n29127 = controllable_nhgrant0 & ~n29126;
  assign n29128 = ~n14166 & ~n29127;
  assign n29129 = ~n3281 & ~n29128;
  assign n29130 = ~n3281 & ~n29129;
  assign n29131 = n3378 & ~n29130;
  assign n29132 = ~n14590 & ~n29031;
  assign n29133 = controllable_nhgrant0 & ~n29132;
  assign n29134 = ~n14180 & ~n29133;
  assign n29135 = ~n3281 & ~n29134;
  assign n29136 = ~n4089 & ~n29135;
  assign n29137 = ~n3378 & ~n29136;
  assign n29138 = ~n29131 & ~n29137;
  assign n29139 = n3492 & ~n29138;
  assign n29140 = ~n14433 & ~n29139;
  assign n29141 = n3485 & ~n29140;
  assign n29142 = ~n14432 & ~n29141;
  assign n29143 = n3476 & ~n29142;
  assign n29144 = ~n29125 & ~n29143;
  assign n29145 = n3374 & ~n29144;
  assign n29146 = ~n14439 & ~n29145;
  assign n29147 = n3655 & ~n29146;
  assign n29148 = ~n14618 & ~n29024;
  assign n29149 = controllable_nhgrant0 & ~n29148;
  assign n29150 = ~n14166 & ~n29149;
  assign n29151 = ~n3281 & ~n29150;
  assign n29152 = ~n3281 & ~n29151;
  assign n29153 = n3378 & ~n29152;
  assign n29154 = ~n14626 & ~n29031;
  assign n29155 = controllable_nhgrant0 & ~n29154;
  assign n29156 = ~n14180 & ~n29155;
  assign n29157 = ~n3281 & ~n29156;
  assign n29158 = ~n3950 & ~n29157;
  assign n29159 = ~n3378 & ~n29158;
  assign n29160 = ~n29153 & ~n29159;
  assign n29161 = n3492 & ~n29160;
  assign n29162 = ~n3493 & ~n29161;
  assign n29163 = n3485 & ~n29162;
  assign n29164 = ~n3486 & ~n29163;
  assign n29165 = ~n3476 & ~n29164;
  assign n29166 = ~n14654 & ~n29024;
  assign n29167 = controllable_nhgrant0 & ~n29166;
  assign n29168 = ~n14166 & ~n29167;
  assign n29169 = ~n3281 & ~n29168;
  assign n29170 = ~n3281 & ~n29169;
  assign n29171 = n3378 & ~n29170;
  assign n29172 = ~n14676 & ~n29031;
  assign n29173 = controllable_nhgrant0 & ~n29172;
  assign n29174 = ~n14180 & ~n29173;
  assign n29175 = ~n3281 & ~n29174;
  assign n29176 = ~n4089 & ~n29175;
  assign n29177 = ~n3378 & ~n29176;
  assign n29178 = ~n29171 & ~n29177;
  assign n29179 = n3492 & ~n29178;
  assign n29180 = ~n14433 & ~n29179;
  assign n29181 = n3485 & ~n29180;
  assign n29182 = ~n14432 & ~n29181;
  assign n29183 = n3476 & ~n29182;
  assign n29184 = ~n29165 & ~n29183;
  assign n29185 = n3374 & ~n29184;
  assign n29186 = ~n14439 & ~n29185;
  assign n29187 = ~n3655 & ~n29186;
  assign n29188 = ~n29147 & ~n29187;
  assign n29189 = ~n3652 & ~n29188;
  assign n29190 = ~n29107 & ~n29189;
  assign n29191 = ~n3368 & ~n29190;
  assign n29192 = controllable_hgrant3 & ~n14722;
  assign n29193 = ~n14711 & ~n29192;
  assign n29194 = controllable_nhgrant0 & ~n29193;
  assign n29195 = ~n14725 & ~n29194;
  assign n29196 = ~n3281 & ~n29195;
  assign n29197 = ~n3281 & ~n29196;
  assign n29198 = n3492 & ~n29197;
  assign n29199 = n3492 & ~n29198;
  assign n29200 = n3485 & ~n29199;
  assign n29201 = n3485 & ~n29200;
  assign n29202 = ~n3476 & ~n29201;
  assign n29203 = ~n14744 & ~n29192;
  assign n29204 = controllable_nhgrant0 & ~n29203;
  assign n29205 = ~n14725 & ~n29204;
  assign n29206 = ~n3281 & ~n29205;
  assign n29207 = ~n3281 & ~n29206;
  assign n29208 = n3492 & ~n29207;
  assign n29209 = n3492 & ~n29208;
  assign n29210 = n3485 & ~n29209;
  assign n29211 = n3485 & ~n29210;
  assign n29212 = n3476 & ~n29211;
  assign n29213 = ~n29202 & ~n29212;
  assign n29214 = n3374 & ~n29213;
  assign n29215 = n3374 & ~n29214;
  assign n29216 = n3655 & ~n29215;
  assign n29217 = ~n14770 & ~n29192;
  assign n29218 = controllable_nhgrant0 & ~n29217;
  assign n29219 = ~n14725 & ~n29218;
  assign n29220 = ~n3281 & ~n29219;
  assign n29221 = ~n3281 & ~n29220;
  assign n29222 = n3492 & ~n29221;
  assign n29223 = n3492 & ~n29222;
  assign n29224 = n3485 & ~n29223;
  assign n29225 = n3485 & ~n29224;
  assign n29226 = ~n3476 & ~n29225;
  assign n29227 = ~n14796 & ~n29192;
  assign n29228 = controllable_nhgrant0 & ~n29227;
  assign n29229 = ~n14725 & ~n29228;
  assign n29230 = ~n3281 & ~n29229;
  assign n29231 = ~n3281 & ~n29230;
  assign n29232 = n3492 & ~n29231;
  assign n29233 = n3492 & ~n29232;
  assign n29234 = n3485 & ~n29233;
  assign n29235 = n3485 & ~n29234;
  assign n29236 = n3476 & ~n29235;
  assign n29237 = ~n29226 & ~n29236;
  assign n29238 = n3374 & ~n29237;
  assign n29239 = n3374 & ~n29238;
  assign n29240 = ~n3655 & ~n29239;
  assign n29241 = ~n29216 & ~n29240;
  assign n29242 = n3652 & ~n29241;
  assign n29243 = ~n14824 & ~n29192;
  assign n29244 = controllable_nhgrant0 & ~n29243;
  assign n29245 = ~n14725 & ~n29244;
  assign n29246 = ~n3281 & ~n29245;
  assign n29247 = ~n3281 & ~n29246;
  assign n29248 = n3492 & ~n29247;
  assign n29249 = n3492 & ~n29248;
  assign n29250 = n3485 & ~n29249;
  assign n29251 = n3485 & ~n29250;
  assign n29252 = ~n3476 & ~n29251;
  assign n29253 = ~n14882 & ~n29192;
  assign n29254 = controllable_nhgrant0 & ~n29253;
  assign n29255 = ~n14725 & ~n29254;
  assign n29256 = ~n3281 & ~n29255;
  assign n29257 = ~n3281 & ~n29256;
  assign n29258 = n3492 & ~n29257;
  assign n29259 = ~n14836 & ~n29258;
  assign n29260 = n3485 & ~n29259;
  assign n29261 = ~n14835 & ~n29260;
  assign n29262 = n3476 & ~n29261;
  assign n29263 = ~n29252 & ~n29262;
  assign n29264 = n3374 & ~n29263;
  assign n29265 = n3374 & ~n29264;
  assign n29266 = n3655 & ~n29265;
  assign n29267 = ~n14908 & ~n29192;
  assign n29268 = controllable_nhgrant0 & ~n29267;
  assign n29269 = ~n14725 & ~n29268;
  assign n29270 = ~n3281 & ~n29269;
  assign n29271 = ~n3281 & ~n29270;
  assign n29272 = n3492 & ~n29271;
  assign n29273 = n3492 & ~n29272;
  assign n29274 = n3485 & ~n29273;
  assign n29275 = n3485 & ~n29274;
  assign n29276 = ~n3476 & ~n29275;
  assign n29277 = ~n14934 & ~n29192;
  assign n29278 = controllable_nhgrant0 & ~n29277;
  assign n29279 = ~n14725 & ~n29278;
  assign n29280 = ~n3281 & ~n29279;
  assign n29281 = ~n3281 & ~n29280;
  assign n29282 = n3492 & ~n29281;
  assign n29283 = ~n14836 & ~n29282;
  assign n29284 = n3485 & ~n29283;
  assign n29285 = ~n14835 & ~n29284;
  assign n29286 = n3476 & ~n29285;
  assign n29287 = ~n29276 & ~n29286;
  assign n29288 = n3374 & ~n29287;
  assign n29289 = n3374 & ~n29288;
  assign n29290 = ~n3655 & ~n29289;
  assign n29291 = ~n29266 & ~n29290;
  assign n29292 = ~n3652 & ~n29291;
  assign n29293 = ~n29242 & ~n29292;
  assign n29294 = n3368 & ~n29293;
  assign n29295 = ~n29191 & ~n29294;
  assign n29296 = ~n3362 & ~n29295;
  assign n29297 = ~n3362 & ~n29296;
  assign n29298 = ~n3359 & ~n29297;
  assign n29299 = ~n3359 & ~n29298;
  assign n29300 = n3356 & ~n29299;
  assign n29301 = ~n14959 & ~n25655;
  assign n29302 = n3492 & ~n29301;
  assign n29303 = ~n3631 & ~n29302;
  assign n29304 = n3485 & ~n29303;
  assign n29305 = ~n3630 & ~n29304;
  assign n29306 = ~n3374 & ~n29305;
  assign n29307 = ~n3910 & ~n5260;
  assign n29308 = controllable_hmaster1 & ~n29307;
  assign n29309 = ~n5263 & ~n29308;
  assign n29310 = i_hbusreq3 & ~n29309;
  assign n29311 = ~n3935 & ~n5277;
  assign n29312 = controllable_hmaster1 & ~n29311;
  assign n29313 = ~n5281 & ~n29312;
  assign n29314 = ~i_hbusreq3 & ~n29313;
  assign n29315 = ~n29310 & ~n29314;
  assign n29316 = ~controllable_hmaster2 & ~n29315;
  assign n29317 = ~n12033 & ~n29316;
  assign n29318 = controllable_hgrant3 & ~n29317;
  assign n29319 = ~n14985 & ~n29318;
  assign n29320 = controllable_nhgrant0 & ~n29319;
  assign n29321 = ~n15006 & ~n29320;
  assign n29322 = ~n3281 & ~n29321;
  assign n29323 = ~n3950 & ~n29322;
  assign n29324 = n3378 & ~n29323;
  assign n29325 = ~n15022 & ~n25684;
  assign n29326 = controllable_nhgrant0 & ~n29325;
  assign n29327 = ~n5534 & ~n29326;
  assign n29328 = ~n3281 & ~n29327;
  assign n29329 = ~n3950 & ~n29328;
  assign n29330 = ~n3378 & ~n29329;
  assign n29331 = ~n29324 & ~n29330;
  assign n29332 = n3492 & ~n29331;
  assign n29333 = ~n3631 & ~n29332;
  assign n29334 = n3485 & ~n29333;
  assign n29335 = ~n3630 & ~n29334;
  assign n29336 = ~n3476 & ~n29335;
  assign n29337 = ~n5587 & ~n5764;
  assign n29338 = controllable_hmaster1 & ~n29337;
  assign n29339 = ~n5591 & ~n29338;
  assign n29340 = i_hbusreq3 & ~n29339;
  assign n29341 = ~n5605 & ~n5787;
  assign n29342 = controllable_hmaster1 & ~n29341;
  assign n29343 = ~n5609 & ~n29342;
  assign n29344 = ~i_hbusreq3 & ~n29343;
  assign n29345 = ~n29340 & ~n29344;
  assign n29346 = ~controllable_hmaster2 & ~n29345;
  assign n29347 = ~n12233 & ~n29346;
  assign n29348 = controllable_hgrant3 & ~n29347;
  assign n29349 = ~n15074 & ~n29348;
  assign n29350 = controllable_nhgrant0 & ~n29349;
  assign n29351 = ~n15088 & ~n29350;
  assign n29352 = ~n3281 & ~n29351;
  assign n29353 = ~n4089 & ~n29352;
  assign n29354 = n3378 & ~n29353;
  assign n29355 = ~n15106 & ~n25726;
  assign n29356 = controllable_nhgrant0 & ~n29355;
  assign n29357 = ~n6082 & ~n29356;
  assign n29358 = ~n3281 & ~n29357;
  assign n29359 = ~n4089 & ~n29358;
  assign n29360 = ~n3378 & ~n29359;
  assign n29361 = ~n29354 & ~n29360;
  assign n29362 = n3492 & ~n29361;
  assign n29363 = ~n3631 & ~n29362;
  assign n29364 = n3485 & ~n29363;
  assign n29365 = ~n3630 & ~n29364;
  assign n29366 = n3476 & ~n29365;
  assign n29367 = ~n29336 & ~n29366;
  assign n29368 = n3374 & ~n29367;
  assign n29369 = ~n29306 & ~n29368;
  assign n29370 = n3655 & ~n29369;
  assign n29371 = ~n14959 & ~n25748;
  assign n29372 = n3492 & ~n29371;
  assign n29373 = ~n3631 & ~n29372;
  assign n29374 = n3485 & ~n29373;
  assign n29375 = ~n3630 & ~n29374;
  assign n29376 = ~n3374 & ~n29375;
  assign n29377 = ~n15140 & ~n29318;
  assign n29378 = controllable_nhgrant0 & ~n29377;
  assign n29379 = ~n15006 & ~n29378;
  assign n29380 = ~n3281 & ~n29379;
  assign n29381 = ~n3950 & ~n29380;
  assign n29382 = n3378 & ~n29381;
  assign n29383 = ~n15158 & ~n25684;
  assign n29384 = controllable_nhgrant0 & ~n29383;
  assign n29385 = ~n5534 & ~n29384;
  assign n29386 = ~n3281 & ~n29385;
  assign n29387 = ~n3950 & ~n29386;
  assign n29388 = ~n3378 & ~n29387;
  assign n29389 = ~n29382 & ~n29388;
  assign n29390 = n3492 & ~n29389;
  assign n29391 = ~n3631 & ~n29390;
  assign n29392 = n3485 & ~n29391;
  assign n29393 = ~n3630 & ~n29392;
  assign n29394 = ~n3476 & ~n29393;
  assign n29395 = ~n15186 & ~n29348;
  assign n29396 = controllable_nhgrant0 & ~n29395;
  assign n29397 = ~n15088 & ~n29396;
  assign n29398 = ~n3281 & ~n29397;
  assign n29399 = ~n4089 & ~n29398;
  assign n29400 = n3378 & ~n29399;
  assign n29401 = ~n15206 & ~n25726;
  assign n29402 = controllable_nhgrant0 & ~n29401;
  assign n29403 = ~n6082 & ~n29402;
  assign n29404 = ~n3281 & ~n29403;
  assign n29405 = ~n4089 & ~n29404;
  assign n29406 = ~n3378 & ~n29405;
  assign n29407 = ~n29400 & ~n29406;
  assign n29408 = n3492 & ~n29407;
  assign n29409 = ~n3631 & ~n29408;
  assign n29410 = n3485 & ~n29409;
  assign n29411 = ~n3630 & ~n29410;
  assign n29412 = n3476 & ~n29411;
  assign n29413 = ~n29394 & ~n29412;
  assign n29414 = n3374 & ~n29413;
  assign n29415 = ~n29376 & ~n29414;
  assign n29416 = ~n3655 & ~n29415;
  assign n29417 = ~n29370 & ~n29416;
  assign n29418 = n3652 & ~n29417;
  assign n29419 = ~n15244 & ~n25649;
  assign n29420 = controllable_nhgrant0 & ~n29419;
  assign n29421 = ~n5245 & ~n29420;
  assign n29422 = ~n3281 & ~n29421;
  assign n29423 = ~n3783 & ~n29422;
  assign n29424 = ~n3378 & ~n29423;
  assign n29425 = ~n15225 & ~n29424;
  assign n29426 = n3492 & ~n29425;
  assign n29427 = ~n3631 & ~n29426;
  assign n29428 = n3485 & ~n29427;
  assign n29429 = ~n3630 & ~n29428;
  assign n29430 = ~n3476 & ~n29429;
  assign n29431 = ~n15258 & ~n29426;
  assign n29432 = n3485 & ~n29431;
  assign n29433 = ~n15257 & ~n29432;
  assign n29434 = n3476 & ~n29433;
  assign n29435 = ~n29430 & ~n29434;
  assign n29436 = ~n3374 & ~n29435;
  assign n29437 = ~n15313 & ~n29318;
  assign n29438 = controllable_nhgrant0 & ~n29437;
  assign n29439 = ~n15006 & ~n29438;
  assign n29440 = ~n3281 & ~n29439;
  assign n29441 = ~n3950 & ~n29440;
  assign n29442 = n3378 & ~n29441;
  assign n29443 = ~n15344 & ~n25684;
  assign n29444 = controllable_nhgrant0 & ~n29443;
  assign n29445 = ~n5534 & ~n29444;
  assign n29446 = ~n3281 & ~n29445;
  assign n29447 = ~n3950 & ~n29446;
  assign n29448 = ~n3378 & ~n29447;
  assign n29449 = ~n29442 & ~n29448;
  assign n29450 = n3492 & ~n29449;
  assign n29451 = ~n3631 & ~n29450;
  assign n29452 = n3485 & ~n29451;
  assign n29453 = ~n3630 & ~n29452;
  assign n29454 = ~n3476 & ~n29453;
  assign n29455 = ~n15413 & ~n29348;
  assign n29456 = controllable_nhgrant0 & ~n29455;
  assign n29457 = ~n15088 & ~n29456;
  assign n29458 = ~n3281 & ~n29457;
  assign n29459 = ~n4089 & ~n29458;
  assign n29460 = n3378 & ~n29459;
  assign n29461 = ~n15456 & ~n25726;
  assign n29462 = controllable_nhgrant0 & ~n29461;
  assign n29463 = ~n6082 & ~n29462;
  assign n29464 = ~n3281 & ~n29463;
  assign n29465 = ~n4089 & ~n29464;
  assign n29466 = ~n3378 & ~n29465;
  assign n29467 = ~n29460 & ~n29466;
  assign n29468 = n3492 & ~n29467;
  assign n29469 = ~n15258 & ~n29468;
  assign n29470 = n3485 & ~n29469;
  assign n29471 = ~n15257 & ~n29470;
  assign n29472 = n3476 & ~n29471;
  assign n29473 = ~n29454 & ~n29472;
  assign n29474 = n3374 & ~n29473;
  assign n29475 = ~n29436 & ~n29474;
  assign n29476 = n3655 & ~n29475;
  assign n29477 = ~n15490 & ~n25649;
  assign n29478 = controllable_nhgrant0 & ~n29477;
  assign n29479 = ~n5245 & ~n29478;
  assign n29480 = ~n3281 & ~n29479;
  assign n29481 = ~n3783 & ~n29480;
  assign n29482 = ~n3378 & ~n29481;
  assign n29483 = ~n15225 & ~n29482;
  assign n29484 = n3492 & ~n29483;
  assign n29485 = ~n3631 & ~n29484;
  assign n29486 = n3485 & ~n29485;
  assign n29487 = ~n3630 & ~n29486;
  assign n29488 = ~n3476 & ~n29487;
  assign n29489 = ~n15258 & ~n29484;
  assign n29490 = n3485 & ~n29489;
  assign n29491 = ~n15257 & ~n29490;
  assign n29492 = n3476 & ~n29491;
  assign n29493 = ~n29488 & ~n29492;
  assign n29494 = ~n3374 & ~n29493;
  assign n29495 = ~n15520 & ~n29318;
  assign n29496 = controllable_nhgrant0 & ~n29495;
  assign n29497 = ~n15006 & ~n29496;
  assign n29498 = ~n3281 & ~n29497;
  assign n29499 = ~n3950 & ~n29498;
  assign n29500 = n3378 & ~n29499;
  assign n29501 = ~n15554 & ~n25684;
  assign n29502 = controllable_nhgrant0 & ~n29501;
  assign n29503 = ~n5534 & ~n29502;
  assign n29504 = ~n3281 & ~n29503;
  assign n29505 = ~n3950 & ~n29504;
  assign n29506 = ~n3378 & ~n29505;
  assign n29507 = ~n29500 & ~n29506;
  assign n29508 = n3492 & ~n29507;
  assign n29509 = ~n3631 & ~n29508;
  assign n29510 = n3485 & ~n29509;
  assign n29511 = ~n3630 & ~n29510;
  assign n29512 = ~n3476 & ~n29511;
  assign n29513 = ~n15582 & ~n29348;
  assign n29514 = controllable_nhgrant0 & ~n29513;
  assign n29515 = ~n15088 & ~n29514;
  assign n29516 = ~n3281 & ~n29515;
  assign n29517 = ~n4089 & ~n29516;
  assign n29518 = n3378 & ~n29517;
  assign n29519 = ~n15618 & ~n25726;
  assign n29520 = controllable_nhgrant0 & ~n29519;
  assign n29521 = ~n6082 & ~n29520;
  assign n29522 = ~n3281 & ~n29521;
  assign n29523 = ~n4089 & ~n29522;
  assign n29524 = ~n3378 & ~n29523;
  assign n29525 = ~n29518 & ~n29524;
  assign n29526 = n3492 & ~n29525;
  assign n29527 = ~n15258 & ~n29526;
  assign n29528 = n3485 & ~n29527;
  assign n29529 = ~n15257 & ~n29528;
  assign n29530 = n3476 & ~n29529;
  assign n29531 = ~n29512 & ~n29530;
  assign n29532 = n3374 & ~n29531;
  assign n29533 = ~n29494 & ~n29532;
  assign n29534 = ~n3655 & ~n29533;
  assign n29535 = ~n29476 & ~n29534;
  assign n29536 = ~n3652 & ~n29535;
  assign n29537 = ~n29418 & ~n29536;
  assign n29538 = ~n3368 & ~n29537;
  assign n29539 = ~n4611 & ~n5260;
  assign n29540 = controllable_hmaster1 & ~n29539;
  assign n29541 = ~n5263 & ~n29540;
  assign n29542 = i_hbusreq3 & ~n29541;
  assign n29543 = ~n4636 & ~n5277;
  assign n29544 = controllable_hmaster1 & ~n29543;
  assign n29545 = ~n5281 & ~n29544;
  assign n29546 = ~i_hbusreq3 & ~n29545;
  assign n29547 = ~n29542 & ~n29546;
  assign n29548 = ~controllable_hmaster2 & ~n29547;
  assign n29549 = ~n12033 & ~n29548;
  assign n29550 = controllable_hgrant3 & ~n29549;
  assign n29551 = ~n15654 & ~n29550;
  assign n29552 = controllable_nhgrant0 & ~n29551;
  assign n29553 = ~n15675 & ~n29552;
  assign n29554 = ~n3281 & ~n29553;
  assign n29555 = ~n3281 & ~n29554;
  assign n29556 = n3378 & ~n29555;
  assign n29557 = ~n4611 & ~n5046;
  assign n29558 = controllable_hmaster1 & ~n29557;
  assign n29559 = ~n25672 & ~n29558;
  assign n29560 = i_hbusreq3 & ~n29559;
  assign n29561 = ~n4636 & ~n5071;
  assign n29562 = controllable_hmaster1 & ~n29561;
  assign n29563 = ~n25678 & ~n29562;
  assign n29564 = ~i_hbusreq3 & ~n29563;
  assign n29565 = ~n29560 & ~n29564;
  assign n29566 = ~controllable_hmaster2 & ~n29565;
  assign n29567 = ~n5498 & ~n29566;
  assign n29568 = controllable_hgrant3 & ~n29567;
  assign n29569 = ~n15695 & ~n29568;
  assign n29570 = controllable_nhgrant0 & ~n29569;
  assign n29571 = ~n15716 & ~n29570;
  assign n29572 = ~n3281 & ~n29571;
  assign n29573 = ~n3281 & ~n29572;
  assign n29574 = ~n3378 & ~n29573;
  assign n29575 = ~n29556 & ~n29574;
  assign n29576 = n3492 & ~n29575;
  assign n29577 = n3492 & ~n29576;
  assign n29578 = n3485 & ~n29577;
  assign n29579 = n3485 & ~n29578;
  assign n29580 = ~n3476 & ~n29579;
  assign n29581 = ~n5587 & ~n7399;
  assign n29582 = controllable_hmaster1 & ~n29581;
  assign n29583 = ~n5591 & ~n29582;
  assign n29584 = i_hbusreq3 & ~n29583;
  assign n29585 = ~n5605 & ~n7422;
  assign n29586 = controllable_hmaster1 & ~n29585;
  assign n29587 = ~n5609 & ~n29586;
  assign n29588 = ~i_hbusreq3 & ~n29587;
  assign n29589 = ~n29584 & ~n29588;
  assign n29590 = ~controllable_hmaster2 & ~n29589;
  assign n29591 = ~n12233 & ~n29590;
  assign n29592 = controllable_hgrant3 & ~n29591;
  assign n29593 = ~n15769 & ~n29592;
  assign n29594 = controllable_nhgrant0 & ~n29593;
  assign n29595 = ~n15783 & ~n29594;
  assign n29596 = ~n3281 & ~n29595;
  assign n29597 = ~n3281 & ~n29596;
  assign n29598 = n3378 & ~n29597;
  assign n29599 = ~n7636 & ~n25705;
  assign n29600 = controllable_hmaster1 & ~n29599;
  assign n29601 = ~n25708 & ~n29600;
  assign n29602 = i_hbusreq3 & ~n29601;
  assign n29603 = ~n7658 & ~n25713;
  assign n29604 = controllable_hmaster1 & ~n29603;
  assign n29605 = ~n25720 & ~n29604;
  assign n29606 = ~i_hbusreq3 & ~n29605;
  assign n29607 = ~n29602 & ~n29606;
  assign n29608 = ~controllable_hmaster2 & ~n29607;
  assign n29609 = ~n6035 & ~n29608;
  assign n29610 = controllable_hgrant3 & ~n29609;
  assign n29611 = ~n15832 & ~n29610;
  assign n29612 = controllable_nhgrant0 & ~n29611;
  assign n29613 = ~n15846 & ~n29612;
  assign n29614 = ~n3281 & ~n29613;
  assign n29615 = ~n3281 & ~n29614;
  assign n29616 = ~n3378 & ~n29615;
  assign n29617 = ~n29598 & ~n29616;
  assign n29618 = n3492 & ~n29617;
  assign n29619 = n3492 & ~n29618;
  assign n29620 = n3485 & ~n29619;
  assign n29621 = n3485 & ~n29620;
  assign n29622 = n3476 & ~n29621;
  assign n29623 = ~n29580 & ~n29622;
  assign n29624 = n3374 & ~n29623;
  assign n29625 = ~n25917 & ~n29624;
  assign n29626 = n3655 & ~n29625;
  assign n29627 = ~n15872 & ~n29550;
  assign n29628 = controllable_nhgrant0 & ~n29627;
  assign n29629 = ~n15675 & ~n29628;
  assign n29630 = ~n3281 & ~n29629;
  assign n29631 = ~n3281 & ~n29630;
  assign n29632 = n3378 & ~n29631;
  assign n29633 = ~n15890 & ~n29568;
  assign n29634 = controllable_nhgrant0 & ~n29633;
  assign n29635 = ~n15716 & ~n29634;
  assign n29636 = ~n3281 & ~n29635;
  assign n29637 = ~n3281 & ~n29636;
  assign n29638 = ~n3378 & ~n29637;
  assign n29639 = ~n29632 & ~n29638;
  assign n29640 = n3492 & ~n29639;
  assign n29641 = n3492 & ~n29640;
  assign n29642 = n3485 & ~n29641;
  assign n29643 = n3485 & ~n29642;
  assign n29644 = ~n3476 & ~n29643;
  assign n29645 = ~n15918 & ~n29592;
  assign n29646 = controllable_nhgrant0 & ~n29645;
  assign n29647 = ~n15783 & ~n29646;
  assign n29648 = ~n3281 & ~n29647;
  assign n29649 = ~n3281 & ~n29648;
  assign n29650 = n3378 & ~n29649;
  assign n29651 = ~n15959 & ~n29610;
  assign n29652 = controllable_nhgrant0 & ~n29651;
  assign n29653 = ~n15846 & ~n29652;
  assign n29654 = ~n3281 & ~n29653;
  assign n29655 = ~n3281 & ~n29654;
  assign n29656 = ~n3378 & ~n29655;
  assign n29657 = ~n29650 & ~n29656;
  assign n29658 = n3492 & ~n29657;
  assign n29659 = n3492 & ~n29658;
  assign n29660 = n3485 & ~n29659;
  assign n29661 = n3485 & ~n29660;
  assign n29662 = n3476 & ~n29661;
  assign n29663 = ~n29644 & ~n29662;
  assign n29664 = n3374 & ~n29663;
  assign n29665 = ~n25977 & ~n29664;
  assign n29666 = ~n3655 & ~n29665;
  assign n29667 = ~n29626 & ~n29666;
  assign n29668 = n3652 & ~n29667;
  assign n29669 = ~n16042 & ~n25905;
  assign n29670 = controllable_nhgrant0 & ~n29669;
  assign n29671 = ~n7118 & ~n29670;
  assign n29672 = ~n3281 & ~n29671;
  assign n29673 = ~n3281 & ~n29672;
  assign n29674 = ~n3378 & ~n29673;
  assign n29675 = ~n16013 & ~n29674;
  assign n29676 = n3492 & ~n29675;
  assign n29677 = n3492 & ~n29676;
  assign n29678 = n3485 & ~n29677;
  assign n29679 = n3485 & ~n29678;
  assign n29680 = ~n3374 & ~n29679;
  assign n29681 = ~n16094 & ~n29550;
  assign n29682 = controllable_nhgrant0 & ~n29681;
  assign n29683 = ~n15675 & ~n29682;
  assign n29684 = ~n3281 & ~n29683;
  assign n29685 = ~n3281 & ~n29684;
  assign n29686 = n3378 & ~n29685;
  assign n29687 = ~n16155 & ~n29568;
  assign n29688 = controllable_nhgrant0 & ~n29687;
  assign n29689 = ~n15716 & ~n29688;
  assign n29690 = ~n3281 & ~n29689;
  assign n29691 = ~n3281 & ~n29690;
  assign n29692 = ~n3378 & ~n29691;
  assign n29693 = ~n29686 & ~n29692;
  assign n29694 = n3492 & ~n29693;
  assign n29695 = n3492 & ~n29694;
  assign n29696 = n3485 & ~n29695;
  assign n29697 = n3485 & ~n29696;
  assign n29698 = ~n3476 & ~n29697;
  assign n29699 = ~n16237 & ~n29592;
  assign n29700 = controllable_nhgrant0 & ~n29699;
  assign n29701 = ~n15783 & ~n29700;
  assign n29702 = ~n3281 & ~n29701;
  assign n29703 = ~n3281 & ~n29702;
  assign n29704 = n3378 & ~n29703;
  assign n29705 = ~n16340 & ~n29610;
  assign n29706 = controllable_nhgrant0 & ~n29705;
  assign n29707 = ~n15846 & ~n29706;
  assign n29708 = ~n3281 & ~n29707;
  assign n29709 = ~n3281 & ~n29708;
  assign n29710 = ~n3378 & ~n29709;
  assign n29711 = ~n29704 & ~n29710;
  assign n29712 = n3492 & ~n29711;
  assign n29713 = ~n14836 & ~n29712;
  assign n29714 = n3485 & ~n29713;
  assign n29715 = ~n14835 & ~n29714;
  assign n29716 = n3476 & ~n29715;
  assign n29717 = ~n29698 & ~n29716;
  assign n29718 = n3374 & ~n29717;
  assign n29719 = ~n29680 & ~n29718;
  assign n29720 = n3655 & ~n29719;
  assign n29721 = ~n16374 & ~n25905;
  assign n29722 = controllable_nhgrant0 & ~n29721;
  assign n29723 = ~n7118 & ~n29722;
  assign n29724 = ~n3281 & ~n29723;
  assign n29725 = ~n3281 & ~n29724;
  assign n29726 = ~n3378 & ~n29725;
  assign n29727 = ~n16013 & ~n29726;
  assign n29728 = n3492 & ~n29727;
  assign n29729 = n3492 & ~n29728;
  assign n29730 = n3485 & ~n29729;
  assign n29731 = n3485 & ~n29730;
  assign n29732 = ~n3374 & ~n29731;
  assign n29733 = ~n16398 & ~n29550;
  assign n29734 = controllable_nhgrant0 & ~n29733;
  assign n29735 = ~n15675 & ~n29734;
  assign n29736 = ~n3281 & ~n29735;
  assign n29737 = ~n3281 & ~n29736;
  assign n29738 = n3378 & ~n29737;
  assign n29739 = ~n16445 & ~n29568;
  assign n29740 = controllable_nhgrant0 & ~n29739;
  assign n29741 = ~n15716 & ~n29740;
  assign n29742 = ~n3281 & ~n29741;
  assign n29743 = ~n3281 & ~n29742;
  assign n29744 = ~n3378 & ~n29743;
  assign n29745 = ~n29738 & ~n29744;
  assign n29746 = n3492 & ~n29745;
  assign n29747 = n3492 & ~n29746;
  assign n29748 = n3485 & ~n29747;
  assign n29749 = n3485 & ~n29748;
  assign n29750 = ~n3476 & ~n29749;
  assign n29751 = ~n16473 & ~n29592;
  assign n29752 = controllable_nhgrant0 & ~n29751;
  assign n29753 = ~n15783 & ~n29752;
  assign n29754 = ~n3281 & ~n29753;
  assign n29755 = ~n3281 & ~n29754;
  assign n29756 = n3378 & ~n29755;
  assign n29757 = ~n16530 & ~n29610;
  assign n29758 = controllable_nhgrant0 & ~n29757;
  assign n29759 = ~n15846 & ~n29758;
  assign n29760 = ~n3281 & ~n29759;
  assign n29761 = ~n3281 & ~n29760;
  assign n29762 = ~n3378 & ~n29761;
  assign n29763 = ~n29756 & ~n29762;
  assign n29764 = n3492 & ~n29763;
  assign n29765 = ~n14836 & ~n29764;
  assign n29766 = n3485 & ~n29765;
  assign n29767 = ~n14835 & ~n29766;
  assign n29768 = n3476 & ~n29767;
  assign n29769 = ~n29750 & ~n29768;
  assign n29770 = n3374 & ~n29769;
  assign n29771 = ~n29732 & ~n29770;
  assign n29772 = ~n3655 & ~n29771;
  assign n29773 = ~n29720 & ~n29772;
  assign n29774 = ~n3652 & ~n29773;
  assign n29775 = ~n29668 & ~n29774;
  assign n29776 = n3368 & ~n29775;
  assign n29777 = ~n29538 & ~n29776;
  assign n29778 = n3362 & ~n29777;
  assign n29779 = n3492 & ~n29329;
  assign n29780 = ~n3631 & ~n29779;
  assign n29781 = n3485 & ~n29780;
  assign n29782 = ~n3630 & ~n29781;
  assign n29783 = ~n3476 & ~n29782;
  assign n29784 = n3492 & ~n29359;
  assign n29785 = ~n3631 & ~n29784;
  assign n29786 = n3485 & ~n29785;
  assign n29787 = ~n26202 & ~n29786;
  assign n29788 = n3476 & ~n29787;
  assign n29789 = ~n29783 & ~n29788;
  assign n29790 = n3374 & ~n29789;
  assign n29791 = ~n26206 & ~n29790;
  assign n29792 = n3655 & ~n29791;
  assign n29793 = n3492 & ~n29387;
  assign n29794 = ~n3631 & ~n29793;
  assign n29795 = n3485 & ~n29794;
  assign n29796 = ~n3630 & ~n29795;
  assign n29797 = ~n3476 & ~n29796;
  assign n29798 = n3492 & ~n29405;
  assign n29799 = ~n3631 & ~n29798;
  assign n29800 = n3485 & ~n29799;
  assign n29801 = ~n26299 & ~n29800;
  assign n29802 = n3476 & ~n29801;
  assign n29803 = ~n29797 & ~n29802;
  assign n29804 = n3374 & ~n29803;
  assign n29805 = ~n26303 & ~n29804;
  assign n29806 = ~n3655 & ~n29805;
  assign n29807 = ~n29792 & ~n29806;
  assign n29808 = n3652 & ~n29807;
  assign n29809 = n3492 & ~n29423;
  assign n29810 = ~n3631 & ~n29809;
  assign n29811 = n3485 & ~n29810;
  assign n29812 = ~n3630 & ~n29811;
  assign n29813 = ~n3476 & ~n29812;
  assign n29814 = ~n16588 & ~n26396;
  assign n29815 = ~n3485 & ~n29814;
  assign n29816 = ~n15258 & ~n29809;
  assign n29817 = n3485 & ~n29816;
  assign n29818 = ~n29815 & ~n29817;
  assign n29819 = n3476 & ~n29818;
  assign n29820 = ~n29813 & ~n29819;
  assign n29821 = ~n3374 & ~n29820;
  assign n29822 = n3492 & ~n29447;
  assign n29823 = ~n3631 & ~n29822;
  assign n29824 = n3485 & ~n29823;
  assign n29825 = ~n3630 & ~n29824;
  assign n29826 = ~n3476 & ~n29825;
  assign n29827 = n3492 & ~n29465;
  assign n29828 = ~n15258 & ~n29827;
  assign n29829 = n3485 & ~n29828;
  assign n29830 = ~n29815 & ~n29829;
  assign n29831 = n3476 & ~n29830;
  assign n29832 = ~n29826 & ~n29831;
  assign n29833 = n3374 & ~n29832;
  assign n29834 = ~n29821 & ~n29833;
  assign n29835 = n3655 & ~n29834;
  assign n29836 = n3492 & ~n29481;
  assign n29837 = ~n3631 & ~n29836;
  assign n29838 = n3485 & ~n29837;
  assign n29839 = ~n3630 & ~n29838;
  assign n29840 = ~n3476 & ~n29839;
  assign n29841 = ~n16588 & ~n26437;
  assign n29842 = ~n3485 & ~n29841;
  assign n29843 = ~n15258 & ~n29836;
  assign n29844 = n3485 & ~n29843;
  assign n29845 = ~n29842 & ~n29844;
  assign n29846 = n3476 & ~n29845;
  assign n29847 = ~n29840 & ~n29846;
  assign n29848 = ~n3374 & ~n29847;
  assign n29849 = n3492 & ~n29505;
  assign n29850 = ~n3631 & ~n29849;
  assign n29851 = n3485 & ~n29850;
  assign n29852 = ~n3630 & ~n29851;
  assign n29853 = ~n3476 & ~n29852;
  assign n29854 = n3492 & ~n29523;
  assign n29855 = ~n15258 & ~n29854;
  assign n29856 = n3485 & ~n29855;
  assign n29857 = ~n29842 & ~n29856;
  assign n29858 = n3476 & ~n29857;
  assign n29859 = ~n29853 & ~n29858;
  assign n29860 = n3374 & ~n29859;
  assign n29861 = ~n29848 & ~n29860;
  assign n29862 = ~n3655 & ~n29861;
  assign n29863 = ~n29835 & ~n29862;
  assign n29864 = ~n3652 & ~n29863;
  assign n29865 = ~n29808 & ~n29864;
  assign n29866 = ~n3368 & ~n29865;
  assign n29867 = n3492 & ~n29573;
  assign n29868 = n3492 & ~n29867;
  assign n29869 = n3485 & ~n29868;
  assign n29870 = n3485 & ~n29869;
  assign n29871 = ~n3476 & ~n29870;
  assign n29872 = n3492 & ~n29615;
  assign n29873 = n3492 & ~n29872;
  assign n29874 = n3485 & ~n29873;
  assign n29875 = ~n26479 & ~n29874;
  assign n29876 = n3476 & ~n29875;
  assign n29877 = ~n29871 & ~n29876;
  assign n29878 = n3374 & ~n29877;
  assign n29879 = ~n26470 & ~n29878;
  assign n29880 = n3655 & ~n29879;
  assign n29881 = n3492 & ~n29637;
  assign n29882 = n3492 & ~n29881;
  assign n29883 = n3485 & ~n29882;
  assign n29884 = n3485 & ~n29883;
  assign n29885 = ~n3476 & ~n29884;
  assign n29886 = n3492 & ~n29655;
  assign n29887 = n3492 & ~n29886;
  assign n29888 = n3485 & ~n29887;
  assign n29889 = ~n26506 & ~n29888;
  assign n29890 = n3476 & ~n29889;
  assign n29891 = ~n29885 & ~n29890;
  assign n29892 = n3374 & ~n29891;
  assign n29893 = ~n26497 & ~n29892;
  assign n29894 = ~n3655 & ~n29893;
  assign n29895 = ~n29880 & ~n29894;
  assign n29896 = n3652 & ~n29895;
  assign n29897 = n3492 & ~n29673;
  assign n29898 = n3492 & ~n29897;
  assign n29899 = n3485 & ~n29898;
  assign n29900 = n3485 & ~n29899;
  assign n29901 = ~n3476 & ~n29900;
  assign n29902 = ~n8525 & ~n29899;
  assign n29903 = n3476 & ~n29902;
  assign n29904 = ~n29901 & ~n29903;
  assign n29905 = ~n3374 & ~n29904;
  assign n29906 = n3492 & ~n29691;
  assign n29907 = n3492 & ~n29906;
  assign n29908 = n3485 & ~n29907;
  assign n29909 = n3485 & ~n29908;
  assign n29910 = ~n3476 & ~n29909;
  assign n29911 = ~n16686 & ~n26533;
  assign n29912 = ~n3485 & ~n29911;
  assign n29913 = n3492 & ~n29709;
  assign n29914 = ~n14836 & ~n29913;
  assign n29915 = n3485 & ~n29914;
  assign n29916 = ~n29912 & ~n29915;
  assign n29917 = n3476 & ~n29916;
  assign n29918 = ~n29910 & ~n29917;
  assign n29919 = n3374 & ~n29918;
  assign n29920 = ~n29905 & ~n29919;
  assign n29921 = n3655 & ~n29920;
  assign n29922 = n3492 & ~n29725;
  assign n29923 = n3492 & ~n29922;
  assign n29924 = n3485 & ~n29923;
  assign n29925 = n3485 & ~n29924;
  assign n29926 = ~n3476 & ~n29925;
  assign n29927 = ~n8525 & ~n29924;
  assign n29928 = n3476 & ~n29927;
  assign n29929 = ~n29926 & ~n29928;
  assign n29930 = ~n3374 & ~n29929;
  assign n29931 = n3492 & ~n29743;
  assign n29932 = n3492 & ~n29931;
  assign n29933 = n3485 & ~n29932;
  assign n29934 = n3485 & ~n29933;
  assign n29935 = ~n3476 & ~n29934;
  assign n29936 = ~n16686 & ~n26560;
  assign n29937 = ~n3485 & ~n29936;
  assign n29938 = n3492 & ~n29761;
  assign n29939 = ~n14836 & ~n29938;
  assign n29940 = n3485 & ~n29939;
  assign n29941 = ~n29937 & ~n29940;
  assign n29942 = n3476 & ~n29941;
  assign n29943 = ~n29935 & ~n29942;
  assign n29944 = n3374 & ~n29943;
  assign n29945 = ~n29930 & ~n29944;
  assign n29946 = ~n3655 & ~n29945;
  assign n29947 = ~n29921 & ~n29946;
  assign n29948 = ~n3652 & ~n29947;
  assign n29949 = ~n29896 & ~n29948;
  assign n29950 = n3368 & ~n29949;
  assign n29951 = ~n29866 & ~n29950;
  assign n29952 = ~n3362 & ~n29951;
  assign n29953 = ~n29778 & ~n29952;
  assign n29954 = n3359 & ~n29953;
  assign n29955 = ~n26580 & ~n29786;
  assign n29956 = n3476 & ~n29955;
  assign n29957 = ~n29783 & ~n29956;
  assign n29958 = n3374 & ~n29957;
  assign n29959 = ~n26584 & ~n29958;
  assign n29960 = n3655 & ~n29959;
  assign n29961 = ~n26591 & ~n29800;
  assign n29962 = n3476 & ~n29961;
  assign n29963 = ~n29797 & ~n29962;
  assign n29964 = n3374 & ~n29963;
  assign n29965 = ~n26595 & ~n29964;
  assign n29966 = ~n3655 & ~n29965;
  assign n29967 = ~n29960 & ~n29966;
  assign n29968 = n3652 & ~n29967;
  assign n29969 = ~n26604 & ~n29817;
  assign n29970 = n3476 & ~n29969;
  assign n29971 = ~n29813 & ~n29970;
  assign n29972 = ~n3374 & ~n29971;
  assign n29973 = ~n26604 & ~n29829;
  assign n29974 = n3476 & ~n29973;
  assign n29975 = ~n29826 & ~n29974;
  assign n29976 = n3374 & ~n29975;
  assign n29977 = ~n29972 & ~n29976;
  assign n29978 = n3655 & ~n29977;
  assign n29979 = ~n26615 & ~n29844;
  assign n29980 = n3476 & ~n29979;
  assign n29981 = ~n29840 & ~n29980;
  assign n29982 = ~n3374 & ~n29981;
  assign n29983 = ~n26615 & ~n29856;
  assign n29984 = n3476 & ~n29983;
  assign n29985 = ~n29853 & ~n29984;
  assign n29986 = n3374 & ~n29985;
  assign n29987 = ~n29982 & ~n29986;
  assign n29988 = ~n3655 & ~n29987;
  assign n29989 = ~n29978 & ~n29988;
  assign n29990 = ~n3652 & ~n29989;
  assign n29991 = ~n29968 & ~n29990;
  assign n29992 = ~n3368 & ~n29991;
  assign n29993 = ~n26634 & ~n29874;
  assign n29994 = n3476 & ~n29993;
  assign n29995 = ~n29871 & ~n29994;
  assign n29996 = n3374 & ~n29995;
  assign n29997 = ~n26633 & ~n29996;
  assign n29998 = n3655 & ~n29997;
  assign n29999 = ~n26645 & ~n29888;
  assign n30000 = n3476 & ~n29999;
  assign n30001 = ~n29885 & ~n30000;
  assign n30002 = n3374 & ~n30001;
  assign n30003 = ~n26644 & ~n30002;
  assign n30004 = ~n3655 & ~n30003;
  assign n30005 = ~n29998 & ~n30004;
  assign n30006 = n3652 & ~n30005;
  assign n30007 = ~n8689 & ~n29899;
  assign n30008 = n3476 & ~n30007;
  assign n30009 = ~n29901 & ~n30008;
  assign n30010 = ~n3374 & ~n30009;
  assign n30011 = ~n26658 & ~n29915;
  assign n30012 = n3476 & ~n30011;
  assign n30013 = ~n29910 & ~n30012;
  assign n30014 = n3374 & ~n30013;
  assign n30015 = ~n30010 & ~n30014;
  assign n30016 = n3655 & ~n30015;
  assign n30017 = ~n8689 & ~n29924;
  assign n30018 = n3476 & ~n30017;
  assign n30019 = ~n29926 & ~n30018;
  assign n30020 = ~n3374 & ~n30019;
  assign n30021 = ~n26669 & ~n29940;
  assign n30022 = n3476 & ~n30021;
  assign n30023 = ~n29935 & ~n30022;
  assign n30024 = n3374 & ~n30023;
  assign n30025 = ~n30020 & ~n30024;
  assign n30026 = ~n3655 & ~n30025;
  assign n30027 = ~n30016 & ~n30026;
  assign n30028 = ~n3652 & ~n30027;
  assign n30029 = ~n30006 & ~n30028;
  assign n30030 = n3368 & ~n30029;
  assign n30031 = ~n29992 & ~n30030;
  assign n30032 = n3362 & ~n30031;
  assign n30033 = n3378 & ~n29329;
  assign n30034 = ~n26711 & ~n30033;
  assign n30035 = n3492 & ~n30034;
  assign n30036 = ~n3631 & ~n30035;
  assign n30037 = n3485 & ~n30036;
  assign n30038 = ~n3630 & ~n30037;
  assign n30039 = ~n3476 & ~n30038;
  assign n30040 = n3378 & ~n29359;
  assign n30041 = ~n26726 & ~n30040;
  assign n30042 = n3492 & ~n30041;
  assign n30043 = ~n26200 & ~n30042;
  assign n30044 = n3485 & ~n30043;
  assign n30045 = ~n26580 & ~n30044;
  assign n30046 = n3476 & ~n30045;
  assign n30047 = ~n30039 & ~n30046;
  assign n30048 = n3374 & ~n30047;
  assign n30049 = ~n26702 & ~n30048;
  assign n30050 = n3655 & ~n30049;
  assign n30051 = n3378 & ~n29387;
  assign n30052 = ~n26762 & ~n30051;
  assign n30053 = n3492 & ~n30052;
  assign n30054 = ~n3631 & ~n30053;
  assign n30055 = n3485 & ~n30054;
  assign n30056 = ~n3630 & ~n30055;
  assign n30057 = ~n3476 & ~n30056;
  assign n30058 = n3378 & ~n29405;
  assign n30059 = ~n26775 & ~n30058;
  assign n30060 = n3492 & ~n30059;
  assign n30061 = ~n26297 & ~n30060;
  assign n30062 = n3485 & ~n30061;
  assign n30063 = ~n26591 & ~n30062;
  assign n30064 = n3476 & ~n30063;
  assign n30065 = ~n30057 & ~n30064;
  assign n30066 = n3374 & ~n30065;
  assign n30067 = ~n26755 & ~n30066;
  assign n30068 = ~n3655 & ~n30067;
  assign n30069 = ~n30050 & ~n30068;
  assign n30070 = n3652 & ~n30069;
  assign n30071 = n3378 & ~n29423;
  assign n30072 = ~n26794 & ~n30071;
  assign n30073 = n3492 & ~n30072;
  assign n30074 = ~n3631 & ~n30073;
  assign n30075 = n3485 & ~n30074;
  assign n30076 = ~n3630 & ~n30075;
  assign n30077 = ~n3476 & ~n30076;
  assign n30078 = ~n26396 & ~n30073;
  assign n30079 = n3485 & ~n30078;
  assign n30080 = ~n26604 & ~n30079;
  assign n30081 = n3476 & ~n30080;
  assign n30082 = ~n30077 & ~n30081;
  assign n30083 = ~n3374 & ~n30082;
  assign n30084 = n3378 & ~n29447;
  assign n30085 = ~n26813 & ~n30084;
  assign n30086 = n3492 & ~n30085;
  assign n30087 = ~n3631 & ~n30086;
  assign n30088 = n3485 & ~n30087;
  assign n30089 = ~n3630 & ~n30088;
  assign n30090 = ~n3476 & ~n30089;
  assign n30091 = n3378 & ~n29465;
  assign n30092 = ~n26826 & ~n30091;
  assign n30093 = n3492 & ~n30092;
  assign n30094 = ~n26396 & ~n30093;
  assign n30095 = n3485 & ~n30094;
  assign n30096 = ~n26604 & ~n30095;
  assign n30097 = n3476 & ~n30096;
  assign n30098 = ~n30090 & ~n30097;
  assign n30099 = n3374 & ~n30098;
  assign n30100 = ~n30083 & ~n30099;
  assign n30101 = n3655 & ~n30100;
  assign n30102 = n3378 & ~n29481;
  assign n30103 = ~n26843 & ~n30102;
  assign n30104 = n3492 & ~n30103;
  assign n30105 = ~n3631 & ~n30104;
  assign n30106 = n3485 & ~n30105;
  assign n30107 = ~n3630 & ~n30106;
  assign n30108 = ~n3476 & ~n30107;
  assign n30109 = ~n26437 & ~n30104;
  assign n30110 = n3485 & ~n30109;
  assign n30111 = ~n26615 & ~n30110;
  assign n30112 = n3476 & ~n30111;
  assign n30113 = ~n30108 & ~n30112;
  assign n30114 = ~n3374 & ~n30113;
  assign n30115 = n3378 & ~n29505;
  assign n30116 = ~n26862 & ~n30115;
  assign n30117 = n3492 & ~n30116;
  assign n30118 = ~n3631 & ~n30117;
  assign n30119 = n3485 & ~n30118;
  assign n30120 = ~n3630 & ~n30119;
  assign n30121 = ~n3476 & ~n30120;
  assign n30122 = n3378 & ~n29523;
  assign n30123 = ~n26875 & ~n30122;
  assign n30124 = n3492 & ~n30123;
  assign n30125 = ~n26437 & ~n30124;
  assign n30126 = n3485 & ~n30125;
  assign n30127 = ~n26615 & ~n30126;
  assign n30128 = n3476 & ~n30127;
  assign n30129 = ~n30121 & ~n30128;
  assign n30130 = n3374 & ~n30129;
  assign n30131 = ~n30114 & ~n30130;
  assign n30132 = ~n3655 & ~n30131;
  assign n30133 = ~n30101 & ~n30132;
  assign n30134 = ~n3652 & ~n30133;
  assign n30135 = ~n30070 & ~n30134;
  assign n30136 = ~n3368 & ~n30135;
  assign n30137 = n3378 & ~n29573;
  assign n30138 = ~n26931 & ~n30137;
  assign n30139 = n3492 & ~n30138;
  assign n30140 = n3492 & ~n30139;
  assign n30141 = n3485 & ~n30140;
  assign n30142 = n3485 & ~n30141;
  assign n30143 = ~n3476 & ~n30142;
  assign n30144 = i_hlock3 & ~n26939;
  assign n30145 = ~i_hlock3 & ~n26950;
  assign n30146 = ~n30144 & ~n30145;
  assign n30147 = i_hbusreq3 & ~n30146;
  assign n30148 = i_hlock3 & ~n26966;
  assign n30149 = ~i_hlock3 & ~n26983;
  assign n30150 = ~n30148 & ~n30149;
  assign n30151 = ~i_hbusreq3 & ~n30150;
  assign n30152 = ~n30147 & ~n30151;
  assign n30153 = controllable_hmaster2 & ~n30152;
  assign n30154 = ~n26944 & ~n27002;
  assign n30155 = controllable_hmaster1 & ~n30154;
  assign n30156 = ~n27006 & ~n30155;
  assign n30157 = i_hlock3 & ~n30156;
  assign n30158 = ~n26955 & ~n27011;
  assign n30159 = controllable_hmaster1 & ~n30158;
  assign n30160 = ~n27015 & ~n30159;
  assign n30161 = ~i_hlock3 & ~n30160;
  assign n30162 = ~n30157 & ~n30161;
  assign n30163 = i_hbusreq3 & ~n30162;
  assign n30164 = ~n26974 & ~n27025;
  assign n30165 = controllable_hmaster1 & ~n30164;
  assign n30166 = ~n27035 & ~n30165;
  assign n30167 = i_hlock3 & ~n30166;
  assign n30168 = ~n26991 & ~n27043;
  assign n30169 = controllable_hmaster1 & ~n30168;
  assign n30170 = ~n27053 & ~n30169;
  assign n30171 = ~i_hlock3 & ~n30170;
  assign n30172 = ~n30167 & ~n30171;
  assign n30173 = ~i_hbusreq3 & ~n30172;
  assign n30174 = ~n30163 & ~n30173;
  assign n30175 = ~controllable_hmaster2 & ~n30174;
  assign n30176 = ~n30153 & ~n30175;
  assign n30177 = controllable_hgrant3 & ~n30176;
  assign n30178 = ~n16948 & ~n30177;
  assign n30179 = controllable_nhgrant0 & ~n30178;
  assign n30180 = ~n16962 & ~n30179;
  assign n30181 = ~n3281 & ~n30180;
  assign n30182 = ~n3281 & ~n30181;
  assign n30183 = n3378 & ~n30182;
  assign n30184 = ~n27144 & ~n30183;
  assign n30185 = n3492 & ~n30184;
  assign n30186 = ~n26477 & ~n30185;
  assign n30187 = n3485 & ~n30186;
  assign n30188 = ~n26634 & ~n30187;
  assign n30189 = n3476 & ~n30188;
  assign n30190 = ~n30143 & ~n30189;
  assign n30191 = n3374 & ~n30190;
  assign n30192 = ~n26909 & ~n30191;
  assign n30193 = n3655 & ~n30192;
  assign n30194 = n3378 & ~n29637;
  assign n30195 = ~n27180 & ~n30194;
  assign n30196 = n3492 & ~n30195;
  assign n30197 = n3492 & ~n30196;
  assign n30198 = n3485 & ~n30197;
  assign n30199 = n3485 & ~n30198;
  assign n30200 = ~n3476 & ~n30199;
  assign n30201 = ~n17016 & ~n30177;
  assign n30202 = controllable_nhgrant0 & ~n30201;
  assign n30203 = ~n16962 & ~n30202;
  assign n30204 = ~n3281 & ~n30203;
  assign n30205 = ~n3281 & ~n30204;
  assign n30206 = n3378 & ~n30205;
  assign n30207 = ~n27198 & ~n30206;
  assign n30208 = n3492 & ~n30207;
  assign n30209 = ~n26504 & ~n30208;
  assign n30210 = n3485 & ~n30209;
  assign n30211 = ~n26645 & ~n30210;
  assign n30212 = n3476 & ~n30211;
  assign n30213 = ~n30200 & ~n30212;
  assign n30214 = n3374 & ~n30213;
  assign n30215 = ~n27173 & ~n30214;
  assign n30216 = ~n3655 & ~n30215;
  assign n30217 = ~n30193 & ~n30216;
  assign n30218 = n3652 & ~n30217;
  assign n30219 = n3378 & ~n29673;
  assign n30220 = ~n27217 & ~n30219;
  assign n30221 = n3492 & ~n30220;
  assign n30222 = n3492 & ~n30221;
  assign n30223 = n3485 & ~n30222;
  assign n30224 = n3485 & ~n30223;
  assign n30225 = ~n3476 & ~n30224;
  assign n30226 = ~n8523 & ~n30221;
  assign n30227 = n3485 & ~n30226;
  assign n30228 = ~n8689 & ~n30227;
  assign n30229 = n3476 & ~n30228;
  assign n30230 = ~n30225 & ~n30229;
  assign n30231 = ~n3374 & ~n30230;
  assign n30232 = n3378 & ~n29691;
  assign n30233 = ~n27236 & ~n30232;
  assign n30234 = n3492 & ~n30233;
  assign n30235 = n3492 & ~n30234;
  assign n30236 = n3485 & ~n30235;
  assign n30237 = n3485 & ~n30236;
  assign n30238 = ~n3476 & ~n30237;
  assign n30239 = ~n17103 & ~n30177;
  assign n30240 = controllable_nhgrant0 & ~n30239;
  assign n30241 = ~n16962 & ~n30240;
  assign n30242 = ~n3281 & ~n30241;
  assign n30243 = ~n3281 & ~n30242;
  assign n30244 = n3378 & ~n30243;
  assign n30245 = ~n27254 & ~n30244;
  assign n30246 = n3492 & ~n30245;
  assign n30247 = ~n26533 & ~n30246;
  assign n30248 = n3485 & ~n30247;
  assign n30249 = ~n26658 & ~n30248;
  assign n30250 = n3476 & ~n30249;
  assign n30251 = ~n30238 & ~n30250;
  assign n30252 = n3374 & ~n30251;
  assign n30253 = ~n30231 & ~n30252;
  assign n30254 = n3655 & ~n30253;
  assign n30255 = n3378 & ~n29725;
  assign n30256 = ~n27271 & ~n30255;
  assign n30257 = n3492 & ~n30256;
  assign n30258 = n3492 & ~n30257;
  assign n30259 = n3485 & ~n30258;
  assign n30260 = n3485 & ~n30259;
  assign n30261 = ~n3476 & ~n30260;
  assign n30262 = ~n8523 & ~n30257;
  assign n30263 = n3485 & ~n30262;
  assign n30264 = ~n8689 & ~n30263;
  assign n30265 = n3476 & ~n30264;
  assign n30266 = ~n30261 & ~n30265;
  assign n30267 = ~n3374 & ~n30266;
  assign n30268 = n3378 & ~n29743;
  assign n30269 = ~n27290 & ~n30268;
  assign n30270 = n3492 & ~n30269;
  assign n30271 = n3492 & ~n30270;
  assign n30272 = n3485 & ~n30271;
  assign n30273 = n3485 & ~n30272;
  assign n30274 = ~n3476 & ~n30273;
  assign n30275 = ~n17188 & ~n30177;
  assign n30276 = controllable_nhgrant0 & ~n30275;
  assign n30277 = ~n16962 & ~n30276;
  assign n30278 = ~n3281 & ~n30277;
  assign n30279 = ~n3281 & ~n30278;
  assign n30280 = n3378 & ~n30279;
  assign n30281 = ~n27308 & ~n30280;
  assign n30282 = n3492 & ~n30281;
  assign n30283 = ~n26560 & ~n30282;
  assign n30284 = n3485 & ~n30283;
  assign n30285 = ~n26669 & ~n30284;
  assign n30286 = n3476 & ~n30285;
  assign n30287 = ~n30274 & ~n30286;
  assign n30288 = n3374 & ~n30287;
  assign n30289 = ~n30267 & ~n30288;
  assign n30290 = ~n3655 & ~n30289;
  assign n30291 = ~n30254 & ~n30290;
  assign n30292 = ~n3652 & ~n30291;
  assign n30293 = ~n30218 & ~n30292;
  assign n30294 = n3368 & ~n30293;
  assign n30295 = ~n30136 & ~n30294;
  assign n30296 = ~n3362 & ~n30295;
  assign n30297 = ~n30032 & ~n30296;
  assign n30298 = ~n3359 & ~n30297;
  assign n30299 = ~n29954 & ~n30298;
  assign n30300 = ~n3356 & ~n30299;
  assign n30301 = ~n29300 & ~n30300;
  assign n30302 = n3345 & ~n30301;
  assign n30303 = ~n29023 & ~n30302;
  assign n30304 = n3341 & ~n30303;
  assign n30305 = ~n27332 & ~n30304;
  assign n30306 = ~n3337 & ~n30305;
  assign n30307 = controllable_hgrant3 & ~n17297;
  assign n30308 = ~n17288 & ~n30307;
  assign n30309 = controllable_nhgrant0 & ~n30308;
  assign n30310 = ~n17300 & ~n30309;
  assign n30311 = ~n3281 & ~n30310;
  assign n30312 = ~n3281 & ~n30311;
  assign n30313 = n3378 & ~n30312;
  assign n30314 = controllable_hgrant3 & ~n17311;
  assign n30315 = ~n17308 & ~n30314;
  assign n30316 = controllable_nhgrant0 & ~n30315;
  assign n30317 = ~n17314 & ~n30316;
  assign n30318 = ~n3281 & ~n30317;
  assign n30319 = ~n3950 & ~n30318;
  assign n30320 = ~n3378 & ~n30319;
  assign n30321 = ~n30313 & ~n30320;
  assign n30322 = n3492 & ~n30321;
  assign n30323 = ~n3493 & ~n30322;
  assign n30324 = n3485 & ~n30323;
  assign n30325 = ~n3486 & ~n30324;
  assign n30326 = ~n3476 & ~n30325;
  assign n30327 = ~n17406 & ~n30307;
  assign n30328 = controllable_nhgrant0 & ~n30327;
  assign n30329 = ~n17300 & ~n30328;
  assign n30330 = ~n3281 & ~n30329;
  assign n30331 = ~n3281 & ~n30330;
  assign n30332 = n3378 & ~n30331;
  assign n30333 = ~n17513 & ~n30314;
  assign n30334 = controllable_nhgrant0 & ~n30333;
  assign n30335 = ~n17314 & ~n30334;
  assign n30336 = ~n3281 & ~n30335;
  assign n30337 = ~n4089 & ~n30336;
  assign n30338 = ~n3378 & ~n30337;
  assign n30339 = ~n30332 & ~n30338;
  assign n30340 = n3492 & ~n30339;
  assign n30341 = ~n3493 & ~n30340;
  assign n30342 = n3485 & ~n30341;
  assign n30343 = ~n3486 & ~n30342;
  assign n30344 = n3476 & ~n30343;
  assign n30345 = ~n30326 & ~n30344;
  assign n30346 = n3374 & ~n30345;
  assign n30347 = ~n17268 & ~n30346;
  assign n30348 = n3655 & ~n30347;
  assign n30349 = ~n17630 & ~n30307;
  assign n30350 = controllable_nhgrant0 & ~n30349;
  assign n30351 = ~n17300 & ~n30350;
  assign n30352 = ~n3281 & ~n30351;
  assign n30353 = ~n3281 & ~n30352;
  assign n30354 = n3378 & ~n30353;
  assign n30355 = ~n17666 & ~n30314;
  assign n30356 = controllable_nhgrant0 & ~n30355;
  assign n30357 = ~n17314 & ~n30356;
  assign n30358 = ~n3281 & ~n30357;
  assign n30359 = ~n3950 & ~n30358;
  assign n30360 = ~n3378 & ~n30359;
  assign n30361 = ~n30354 & ~n30360;
  assign n30362 = n3492 & ~n30361;
  assign n30363 = ~n3493 & ~n30362;
  assign n30364 = n3485 & ~n30363;
  assign n30365 = ~n3486 & ~n30364;
  assign n30366 = ~n3476 & ~n30365;
  assign n30367 = ~n17753 & ~n30307;
  assign n30368 = controllable_nhgrant0 & ~n30367;
  assign n30369 = ~n17300 & ~n30368;
  assign n30370 = ~n3281 & ~n30369;
  assign n30371 = ~n3281 & ~n30370;
  assign n30372 = n3378 & ~n30371;
  assign n30373 = ~n17857 & ~n30314;
  assign n30374 = controllable_nhgrant0 & ~n30373;
  assign n30375 = ~n17314 & ~n30374;
  assign n30376 = ~n3281 & ~n30375;
  assign n30377 = ~n4089 & ~n30376;
  assign n30378 = ~n3378 & ~n30377;
  assign n30379 = ~n30372 & ~n30378;
  assign n30380 = n3492 & ~n30379;
  assign n30381 = ~n17612 & ~n30380;
  assign n30382 = n3485 & ~n30381;
  assign n30383 = ~n17611 & ~n30382;
  assign n30384 = n3476 & ~n30383;
  assign n30385 = ~n30366 & ~n30384;
  assign n30386 = n3374 & ~n30385;
  assign n30387 = ~n17618 & ~n30386;
  assign n30388 = ~n3655 & ~n30387;
  assign n30389 = ~n30348 & ~n30388;
  assign n30390 = n3652 & ~n30389;
  assign n30391 = ~n17887 & ~n30307;
  assign n30392 = controllable_nhgrant0 & ~n30391;
  assign n30393 = ~n17300 & ~n30392;
  assign n30394 = ~n3281 & ~n30393;
  assign n30395 = ~n3281 & ~n30394;
  assign n30396 = n3378 & ~n30395;
  assign n30397 = ~n17895 & ~n30314;
  assign n30398 = controllable_nhgrant0 & ~n30397;
  assign n30399 = ~n17314 & ~n30398;
  assign n30400 = ~n3281 & ~n30399;
  assign n30401 = ~n3950 & ~n30400;
  assign n30402 = ~n3378 & ~n30401;
  assign n30403 = ~n30396 & ~n30402;
  assign n30404 = n3492 & ~n30403;
  assign n30405 = ~n3493 & ~n30404;
  assign n30406 = n3485 & ~n30405;
  assign n30407 = ~n3486 & ~n30406;
  assign n30408 = ~n3476 & ~n30407;
  assign n30409 = ~n17923 & ~n30307;
  assign n30410 = controllable_nhgrant0 & ~n30409;
  assign n30411 = ~n17300 & ~n30410;
  assign n30412 = ~n3281 & ~n30411;
  assign n30413 = ~n3281 & ~n30412;
  assign n30414 = n3378 & ~n30413;
  assign n30415 = ~n17945 & ~n30314;
  assign n30416 = controllable_nhgrant0 & ~n30415;
  assign n30417 = ~n17314 & ~n30416;
  assign n30418 = ~n3281 & ~n30417;
  assign n30419 = ~n4089 & ~n30418;
  assign n30420 = ~n3378 & ~n30419;
  assign n30421 = ~n30414 & ~n30420;
  assign n30422 = n3492 & ~n30421;
  assign n30423 = ~n3493 & ~n30422;
  assign n30424 = n3485 & ~n30423;
  assign n30425 = ~n3486 & ~n30424;
  assign n30426 = n3476 & ~n30425;
  assign n30427 = ~n30408 & ~n30426;
  assign n30428 = n3374 & ~n30427;
  assign n30429 = ~n17268 & ~n30428;
  assign n30430 = n3655 & ~n30429;
  assign n30431 = ~n17973 & ~n30307;
  assign n30432 = controllable_nhgrant0 & ~n30431;
  assign n30433 = ~n17300 & ~n30432;
  assign n30434 = ~n3281 & ~n30433;
  assign n30435 = ~n3281 & ~n30434;
  assign n30436 = n3378 & ~n30435;
  assign n30437 = ~n17981 & ~n30314;
  assign n30438 = controllable_nhgrant0 & ~n30437;
  assign n30439 = ~n17314 & ~n30438;
  assign n30440 = ~n3281 & ~n30439;
  assign n30441 = ~n3950 & ~n30440;
  assign n30442 = ~n3378 & ~n30441;
  assign n30443 = ~n30436 & ~n30442;
  assign n30444 = n3492 & ~n30443;
  assign n30445 = ~n3493 & ~n30444;
  assign n30446 = n3485 & ~n30445;
  assign n30447 = ~n3486 & ~n30446;
  assign n30448 = ~n3476 & ~n30447;
  assign n30449 = ~n18009 & ~n30307;
  assign n30450 = controllable_nhgrant0 & ~n30449;
  assign n30451 = ~n17300 & ~n30450;
  assign n30452 = ~n3281 & ~n30451;
  assign n30453 = ~n3281 & ~n30452;
  assign n30454 = n3378 & ~n30453;
  assign n30455 = ~n18031 & ~n30314;
  assign n30456 = controllable_nhgrant0 & ~n30455;
  assign n30457 = ~n17314 & ~n30456;
  assign n30458 = ~n3281 & ~n30457;
  assign n30459 = ~n4089 & ~n30458;
  assign n30460 = ~n3378 & ~n30459;
  assign n30461 = ~n30454 & ~n30460;
  assign n30462 = n3492 & ~n30461;
  assign n30463 = ~n17612 & ~n30462;
  assign n30464 = n3485 & ~n30463;
  assign n30465 = ~n17611 & ~n30464;
  assign n30466 = n3476 & ~n30465;
  assign n30467 = ~n30448 & ~n30466;
  assign n30468 = n3374 & ~n30467;
  assign n30469 = ~n17618 & ~n30468;
  assign n30470 = ~n3655 & ~n30469;
  assign n30471 = ~n30430 & ~n30470;
  assign n30472 = ~n3652 & ~n30471;
  assign n30473 = ~n30390 & ~n30472;
  assign n30474 = ~n3368 & ~n30473;
  assign n30475 = controllable_hgrant3 & ~n18074;
  assign n30476 = ~n18065 & ~n30475;
  assign n30477 = controllable_nhgrant0 & ~n30476;
  assign n30478 = ~n18077 & ~n30477;
  assign n30479 = ~n3281 & ~n30478;
  assign n30480 = ~n3281 & ~n30479;
  assign n30481 = n3492 & ~n30480;
  assign n30482 = n3492 & ~n30481;
  assign n30483 = n3485 & ~n30482;
  assign n30484 = n3485 & ~n30483;
  assign n30485 = ~n3476 & ~n30484;
  assign n30486 = ~n18113 & ~n30475;
  assign n30487 = controllable_nhgrant0 & ~n30486;
  assign n30488 = ~n18077 & ~n30487;
  assign n30489 = ~n3281 & ~n30488;
  assign n30490 = ~n3281 & ~n30489;
  assign n30491 = n3492 & ~n30490;
  assign n30492 = n3492 & ~n30491;
  assign n30493 = n3485 & ~n30492;
  assign n30494 = n3485 & ~n30493;
  assign n30495 = n3476 & ~n30494;
  assign n30496 = ~n30485 & ~n30495;
  assign n30497 = n3374 & ~n30496;
  assign n30498 = n3374 & ~n30497;
  assign n30499 = n3655 & ~n30498;
  assign n30500 = ~n18139 & ~n30475;
  assign n30501 = controllable_nhgrant0 & ~n30500;
  assign n30502 = ~n18077 & ~n30501;
  assign n30503 = ~n3281 & ~n30502;
  assign n30504 = ~n3281 & ~n30503;
  assign n30505 = n3492 & ~n30504;
  assign n30506 = n3492 & ~n30505;
  assign n30507 = n3485 & ~n30506;
  assign n30508 = n3485 & ~n30507;
  assign n30509 = ~n3476 & ~n30508;
  assign n30510 = ~n18238 & ~n30475;
  assign n30511 = controllable_nhgrant0 & ~n30510;
  assign n30512 = ~n18077 & ~n30511;
  assign n30513 = ~n3281 & ~n30512;
  assign n30514 = ~n3281 & ~n30513;
  assign n30515 = n3492 & ~n30514;
  assign n30516 = ~n18151 & ~n30515;
  assign n30517 = n3485 & ~n30516;
  assign n30518 = ~n18150 & ~n30517;
  assign n30519 = n3476 & ~n30518;
  assign n30520 = ~n30509 & ~n30519;
  assign n30521 = n3374 & ~n30520;
  assign n30522 = n3374 & ~n30521;
  assign n30523 = ~n3655 & ~n30522;
  assign n30524 = ~n30499 & ~n30523;
  assign n30525 = n3652 & ~n30524;
  assign n30526 = ~n18266 & ~n30475;
  assign n30527 = controllable_nhgrant0 & ~n30526;
  assign n30528 = ~n18077 & ~n30527;
  assign n30529 = ~n3281 & ~n30528;
  assign n30530 = ~n3281 & ~n30529;
  assign n30531 = n3492 & ~n30530;
  assign n30532 = n3492 & ~n30531;
  assign n30533 = n3485 & ~n30532;
  assign n30534 = n3485 & ~n30533;
  assign n30535 = ~n3476 & ~n30534;
  assign n30536 = ~n18292 & ~n30475;
  assign n30537 = controllable_nhgrant0 & ~n30536;
  assign n30538 = ~n18077 & ~n30537;
  assign n30539 = ~n3281 & ~n30538;
  assign n30540 = ~n3281 & ~n30539;
  assign n30541 = n3492 & ~n30540;
  assign n30542 = n3492 & ~n30541;
  assign n30543 = n3485 & ~n30542;
  assign n30544 = n3485 & ~n30543;
  assign n30545 = n3476 & ~n30544;
  assign n30546 = ~n30535 & ~n30545;
  assign n30547 = n3374 & ~n30546;
  assign n30548 = n3374 & ~n30547;
  assign n30549 = n3655 & ~n30548;
  assign n30550 = ~n18318 & ~n30475;
  assign n30551 = controllable_nhgrant0 & ~n30550;
  assign n30552 = ~n18077 & ~n30551;
  assign n30553 = ~n3281 & ~n30552;
  assign n30554 = ~n3281 & ~n30553;
  assign n30555 = n3492 & ~n30554;
  assign n30556 = n3492 & ~n30555;
  assign n30557 = n3485 & ~n30556;
  assign n30558 = n3485 & ~n30557;
  assign n30559 = ~n3476 & ~n30558;
  assign n30560 = ~n18344 & ~n30475;
  assign n30561 = controllable_nhgrant0 & ~n30560;
  assign n30562 = ~n18077 & ~n30561;
  assign n30563 = ~n3281 & ~n30562;
  assign n30564 = ~n3281 & ~n30563;
  assign n30565 = n3492 & ~n30564;
  assign n30566 = ~n18151 & ~n30565;
  assign n30567 = n3485 & ~n30566;
  assign n30568 = ~n18150 & ~n30567;
  assign n30569 = n3476 & ~n30568;
  assign n30570 = ~n30559 & ~n30569;
  assign n30571 = n3374 & ~n30570;
  assign n30572 = n3374 & ~n30571;
  assign n30573 = ~n3655 & ~n30572;
  assign n30574 = ~n30549 & ~n30573;
  assign n30575 = ~n3652 & ~n30574;
  assign n30576 = ~n30525 & ~n30575;
  assign n30577 = n3368 & ~n30576;
  assign n30578 = ~n30474 & ~n30577;
  assign n30579 = ~n3362 & ~n30578;
  assign n30580 = ~n3362 & ~n30579;
  assign n30581 = ~n3359 & ~n30580;
  assign n30582 = ~n3359 & ~n30581;
  assign n30583 = n3356 & ~n30582;
  assign n30584 = ~n18369 & ~n25655;
  assign n30585 = n3492 & ~n30584;
  assign n30586 = ~n3631 & ~n30585;
  assign n30587 = n3485 & ~n30586;
  assign n30588 = ~n3630 & ~n30587;
  assign n30589 = ~n3374 & ~n30588;
  assign n30590 = ~controllable_hmaster1 & ~n12088;
  assign n30591 = ~n5262 & ~n30590;
  assign n30592 = i_hbusreq3 & ~n30591;
  assign n30593 = ~controllable_hmaster1 & ~n12092;
  assign n30594 = ~n5280 & ~n30593;
  assign n30595 = ~i_hbusreq3 & ~n30594;
  assign n30596 = ~n30592 & ~n30595;
  assign n30597 = ~controllable_hmaster2 & ~n30596;
  assign n30598 = ~n12033 & ~n30597;
  assign n30599 = controllable_hgrant3 & ~n30598;
  assign n30600 = ~n18394 & ~n30599;
  assign n30601 = controllable_nhgrant0 & ~n30600;
  assign n30602 = ~n18416 & ~n30601;
  assign n30603 = ~n3281 & ~n30602;
  assign n30604 = ~n3950 & ~n30603;
  assign n30605 = n3378 & ~n30604;
  assign n30606 = ~n18432 & ~n25684;
  assign n30607 = controllable_nhgrant0 & ~n30606;
  assign n30608 = ~n5534 & ~n30607;
  assign n30609 = ~n3281 & ~n30608;
  assign n30610 = ~n3950 & ~n30609;
  assign n30611 = ~n3378 & ~n30610;
  assign n30612 = ~n30605 & ~n30611;
  assign n30613 = n3492 & ~n30612;
  assign n30614 = ~n3631 & ~n30613;
  assign n30615 = n3485 & ~n30614;
  assign n30616 = ~n3630 & ~n30615;
  assign n30617 = ~n3476 & ~n30616;
  assign n30618 = ~controllable_hmaster1 & ~n12235;
  assign n30619 = ~n5590 & ~n30618;
  assign n30620 = i_hbusreq3 & ~n30619;
  assign n30621 = ~controllable_hmaster1 & ~n12240;
  assign n30622 = ~n5608 & ~n30621;
  assign n30623 = ~i_hbusreq3 & ~n30622;
  assign n30624 = ~n30620 & ~n30623;
  assign n30625 = ~controllable_hmaster2 & ~n30624;
  assign n30626 = ~n12233 & ~n30625;
  assign n30627 = controllable_hgrant3 & ~n30626;
  assign n30628 = ~n18510 & ~n30627;
  assign n30629 = controllable_nhgrant0 & ~n30628;
  assign n30630 = ~n18526 & ~n30629;
  assign n30631 = ~n3281 & ~n30630;
  assign n30632 = ~n4089 & ~n30631;
  assign n30633 = n3378 & ~n30632;
  assign n30634 = ~n18554 & ~n25726;
  assign n30635 = controllable_nhgrant0 & ~n30634;
  assign n30636 = ~n6082 & ~n30635;
  assign n30637 = ~n3281 & ~n30636;
  assign n30638 = ~n4089 & ~n30637;
  assign n30639 = ~n3378 & ~n30638;
  assign n30640 = ~n30633 & ~n30639;
  assign n30641 = n3492 & ~n30640;
  assign n30642 = ~n3631 & ~n30641;
  assign n30643 = n3485 & ~n30642;
  assign n30644 = ~n3630 & ~n30643;
  assign n30645 = n3476 & ~n30644;
  assign n30646 = ~n30617 & ~n30645;
  assign n30647 = n3374 & ~n30646;
  assign n30648 = ~n30589 & ~n30647;
  assign n30649 = n3655 & ~n30648;
  assign n30650 = ~n18616 & ~n25649;
  assign n30651 = controllable_nhgrant0 & ~n30650;
  assign n30652 = ~n5245 & ~n30651;
  assign n30653 = ~n3281 & ~n30652;
  assign n30654 = ~n3783 & ~n30653;
  assign n30655 = ~n3378 & ~n30654;
  assign n30656 = ~n18571 & ~n30655;
  assign n30657 = n3492 & ~n30656;
  assign n30658 = ~n3631 & ~n30657;
  assign n30659 = n3485 & ~n30658;
  assign n30660 = ~n3630 & ~n30659;
  assign n30661 = ~n3476 & ~n30660;
  assign n30662 = ~n18630 & ~n30657;
  assign n30663 = n3485 & ~n30662;
  assign n30664 = ~n18629 & ~n30663;
  assign n30665 = n3476 & ~n30664;
  assign n30666 = ~n30661 & ~n30665;
  assign n30667 = ~n3374 & ~n30666;
  assign n30668 = ~n18703 & ~n30599;
  assign n30669 = controllable_nhgrant0 & ~n30668;
  assign n30670 = ~n18416 & ~n30669;
  assign n30671 = ~n3281 & ~n30670;
  assign n30672 = ~n3950 & ~n30671;
  assign n30673 = n3378 & ~n30672;
  assign n30674 = ~n18746 & ~n25684;
  assign n30675 = controllable_nhgrant0 & ~n30674;
  assign n30676 = ~n5534 & ~n30675;
  assign n30677 = ~n3281 & ~n30676;
  assign n30678 = ~n3950 & ~n30677;
  assign n30679 = ~n3378 & ~n30678;
  assign n30680 = ~n30673 & ~n30679;
  assign n30681 = n3492 & ~n30680;
  assign n30682 = ~n3631 & ~n30681;
  assign n30683 = n3485 & ~n30682;
  assign n30684 = ~n3630 & ~n30683;
  assign n30685 = ~n3476 & ~n30684;
  assign n30686 = ~n18839 & ~n30627;
  assign n30687 = controllable_nhgrant0 & ~n30686;
  assign n30688 = ~n18526 & ~n30687;
  assign n30689 = ~n3281 & ~n30688;
  assign n30690 = ~n4089 & ~n30689;
  assign n30691 = n3378 & ~n30690;
  assign n30692 = ~n18892 & ~n25726;
  assign n30693 = controllable_nhgrant0 & ~n30692;
  assign n30694 = ~n6082 & ~n30693;
  assign n30695 = ~n3281 & ~n30694;
  assign n30696 = ~n4089 & ~n30695;
  assign n30697 = ~n3378 & ~n30696;
  assign n30698 = ~n30691 & ~n30697;
  assign n30699 = n3492 & ~n30698;
  assign n30700 = ~n18630 & ~n30699;
  assign n30701 = n3485 & ~n30700;
  assign n30702 = ~n18629 & ~n30701;
  assign n30703 = n3476 & ~n30702;
  assign n30704 = ~n30685 & ~n30703;
  assign n30705 = n3374 & ~n30704;
  assign n30706 = ~n30667 & ~n30705;
  assign n30707 = ~n3655 & ~n30706;
  assign n30708 = ~n30649 & ~n30707;
  assign n30709 = n3652 & ~n30708;
  assign n30710 = ~n18369 & ~n25802;
  assign n30711 = n3492 & ~n30710;
  assign n30712 = ~n3631 & ~n30711;
  assign n30713 = n3485 & ~n30712;
  assign n30714 = ~n3630 & ~n30713;
  assign n30715 = ~n3374 & ~n30714;
  assign n30716 = ~n18928 & ~n30599;
  assign n30717 = controllable_nhgrant0 & ~n30716;
  assign n30718 = ~n18416 & ~n30717;
  assign n30719 = ~n3281 & ~n30718;
  assign n30720 = ~n3950 & ~n30719;
  assign n30721 = n3378 & ~n30720;
  assign n30722 = ~n18946 & ~n25684;
  assign n30723 = controllable_nhgrant0 & ~n30722;
  assign n30724 = ~n5534 & ~n30723;
  assign n30725 = ~n3281 & ~n30724;
  assign n30726 = ~n3950 & ~n30725;
  assign n30727 = ~n3378 & ~n30726;
  assign n30728 = ~n30721 & ~n30727;
  assign n30729 = n3492 & ~n30728;
  assign n30730 = ~n3631 & ~n30729;
  assign n30731 = n3485 & ~n30730;
  assign n30732 = ~n3630 & ~n30731;
  assign n30733 = ~n3476 & ~n30732;
  assign n30734 = ~n18974 & ~n30627;
  assign n30735 = controllable_nhgrant0 & ~n30734;
  assign n30736 = ~n18526 & ~n30735;
  assign n30737 = ~n3281 & ~n30736;
  assign n30738 = ~n4089 & ~n30737;
  assign n30739 = n3378 & ~n30738;
  assign n30740 = ~n18994 & ~n25726;
  assign n30741 = controllable_nhgrant0 & ~n30740;
  assign n30742 = ~n6082 & ~n30741;
  assign n30743 = ~n3281 & ~n30742;
  assign n30744 = ~n4089 & ~n30743;
  assign n30745 = ~n3378 & ~n30744;
  assign n30746 = ~n30739 & ~n30745;
  assign n30747 = n3492 & ~n30746;
  assign n30748 = ~n3631 & ~n30747;
  assign n30749 = n3485 & ~n30748;
  assign n30750 = ~n3630 & ~n30749;
  assign n30751 = n3476 & ~n30750;
  assign n30752 = ~n30733 & ~n30751;
  assign n30753 = n3374 & ~n30752;
  assign n30754 = ~n30715 & ~n30753;
  assign n30755 = n3655 & ~n30754;
  assign n30756 = ~n19028 & ~n25649;
  assign n30757 = controllable_nhgrant0 & ~n30756;
  assign n30758 = ~n5245 & ~n30757;
  assign n30759 = ~n3281 & ~n30758;
  assign n30760 = ~n3783 & ~n30759;
  assign n30761 = ~n3378 & ~n30760;
  assign n30762 = ~n18571 & ~n30761;
  assign n30763 = n3492 & ~n30762;
  assign n30764 = ~n3631 & ~n30763;
  assign n30765 = n3485 & ~n30764;
  assign n30766 = ~n3630 & ~n30765;
  assign n30767 = ~n3476 & ~n30766;
  assign n30768 = ~n18630 & ~n30763;
  assign n30769 = n3485 & ~n30768;
  assign n30770 = ~n18629 & ~n30769;
  assign n30771 = n3476 & ~n30770;
  assign n30772 = ~n30767 & ~n30771;
  assign n30773 = ~n3374 & ~n30772;
  assign n30774 = ~n19058 & ~n30599;
  assign n30775 = controllable_nhgrant0 & ~n30774;
  assign n30776 = ~n18416 & ~n30775;
  assign n30777 = ~n3281 & ~n30776;
  assign n30778 = ~n3950 & ~n30777;
  assign n30779 = n3378 & ~n30778;
  assign n30780 = ~n19092 & ~n25684;
  assign n30781 = controllable_nhgrant0 & ~n30780;
  assign n30782 = ~n5534 & ~n30781;
  assign n30783 = ~n3281 & ~n30782;
  assign n30784 = ~n3950 & ~n30783;
  assign n30785 = ~n3378 & ~n30784;
  assign n30786 = ~n30779 & ~n30785;
  assign n30787 = n3492 & ~n30786;
  assign n30788 = ~n3631 & ~n30787;
  assign n30789 = n3485 & ~n30788;
  assign n30790 = ~n3630 & ~n30789;
  assign n30791 = ~n3476 & ~n30790;
  assign n30792 = ~n19120 & ~n30627;
  assign n30793 = controllable_nhgrant0 & ~n30792;
  assign n30794 = ~n18526 & ~n30793;
  assign n30795 = ~n3281 & ~n30794;
  assign n30796 = ~n4089 & ~n30795;
  assign n30797 = n3378 & ~n30796;
  assign n30798 = ~n19156 & ~n25726;
  assign n30799 = controllable_nhgrant0 & ~n30798;
  assign n30800 = ~n6082 & ~n30799;
  assign n30801 = ~n3281 & ~n30800;
  assign n30802 = ~n4089 & ~n30801;
  assign n30803 = ~n3378 & ~n30802;
  assign n30804 = ~n30797 & ~n30803;
  assign n30805 = n3492 & ~n30804;
  assign n30806 = ~n18630 & ~n30805;
  assign n30807 = n3485 & ~n30806;
  assign n30808 = ~n18629 & ~n30807;
  assign n30809 = n3476 & ~n30808;
  assign n30810 = ~n30791 & ~n30809;
  assign n30811 = n3374 & ~n30810;
  assign n30812 = ~n30773 & ~n30811;
  assign n30813 = ~n3655 & ~n30812;
  assign n30814 = ~n30755 & ~n30813;
  assign n30815 = ~n3652 & ~n30814;
  assign n30816 = ~n30709 & ~n30815;
  assign n30817 = ~n3368 & ~n30816;
  assign n30818 = ~controllable_hmaster1 & ~n12760;
  assign n30819 = ~n5262 & ~n30818;
  assign n30820 = i_hbusreq3 & ~n30819;
  assign n30821 = ~controllable_hmaster1 & ~n12764;
  assign n30822 = ~n5280 & ~n30821;
  assign n30823 = ~i_hbusreq3 & ~n30822;
  assign n30824 = ~n30820 & ~n30823;
  assign n30825 = ~controllable_hmaster2 & ~n30824;
  assign n30826 = ~n12033 & ~n30825;
  assign n30827 = controllable_hgrant3 & ~n30826;
  assign n30828 = ~n19191 & ~n30827;
  assign n30829 = controllable_nhgrant0 & ~n30828;
  assign n30830 = ~n19213 & ~n30829;
  assign n30831 = ~n3281 & ~n30830;
  assign n30832 = ~n3281 & ~n30831;
  assign n30833 = n3378 & ~n30832;
  assign n30834 = ~controllable_hmaster1 & ~n12814;
  assign n30835 = ~n25671 & ~n30834;
  assign n30836 = i_hbusreq3 & ~n30835;
  assign n30837 = ~n5478 & ~n9743;
  assign n30838 = ~controllable_hmaster1 & ~n30837;
  assign n30839 = ~n25676 & ~n30838;
  assign n30840 = ~i_hbusreq3 & ~n30839;
  assign n30841 = ~n30836 & ~n30840;
  assign n30842 = ~controllable_hmaster2 & ~n30841;
  assign n30843 = ~n5498 & ~n30842;
  assign n30844 = controllable_hgrant3 & ~n30843;
  assign n30845 = ~n19233 & ~n30844;
  assign n30846 = controllable_nhgrant0 & ~n30845;
  assign n30847 = ~n19255 & ~n30846;
  assign n30848 = ~n3281 & ~n30847;
  assign n30849 = ~n3281 & ~n30848;
  assign n30850 = ~n3378 & ~n30849;
  assign n30851 = ~n30833 & ~n30850;
  assign n30852 = n3492 & ~n30851;
  assign n30853 = n3492 & ~n30852;
  assign n30854 = n3485 & ~n30853;
  assign n30855 = n3485 & ~n30854;
  assign n30856 = ~n3476 & ~n30855;
  assign n30857 = ~controllable_hmaster1 & ~n12928;
  assign n30858 = ~n5590 & ~n30857;
  assign n30859 = i_hbusreq3 & ~n30858;
  assign n30860 = ~controllable_hmaster1 & ~n12933;
  assign n30861 = ~n5608 & ~n30860;
  assign n30862 = ~i_hbusreq3 & ~n30861;
  assign n30863 = ~n30859 & ~n30862;
  assign n30864 = ~controllable_hmaster2 & ~n30863;
  assign n30865 = ~n12233 & ~n30864;
  assign n30866 = controllable_hgrant3 & ~n30865;
  assign n30867 = ~n19369 & ~n30866;
  assign n30868 = controllable_nhgrant0 & ~n30867;
  assign n30869 = ~n19385 & ~n30868;
  assign n30870 = ~n3281 & ~n30869;
  assign n30871 = ~n3281 & ~n30870;
  assign n30872 = n3378 & ~n30871;
  assign n30873 = ~controllable_hmaster1 & ~n13050;
  assign n30874 = ~n25707 & ~n30873;
  assign n30875 = i_hbusreq3 & ~n30874;
  assign n30876 = ~n13054 & ~n25718;
  assign n30877 = ~controllable_hmaster1 & ~n30876;
  assign n30878 = ~n25715 & ~n30877;
  assign n30879 = ~i_hbusreq3 & ~n30878;
  assign n30880 = ~n30875 & ~n30879;
  assign n30881 = ~controllable_hmaster2 & ~n30880;
  assign n30882 = ~n6035 & ~n30881;
  assign n30883 = controllable_hgrant3 & ~n30882;
  assign n30884 = ~n19499 & ~n30883;
  assign n30885 = controllable_nhgrant0 & ~n30884;
  assign n30886 = ~n19515 & ~n30885;
  assign n30887 = ~n3281 & ~n30886;
  assign n30888 = ~n3281 & ~n30887;
  assign n30889 = ~n3378 & ~n30888;
  assign n30890 = ~n30872 & ~n30889;
  assign n30891 = n3492 & ~n30890;
  assign n30892 = n3492 & ~n30891;
  assign n30893 = n3485 & ~n30892;
  assign n30894 = n3485 & ~n30893;
  assign n30895 = n3476 & ~n30894;
  assign n30896 = ~n30856 & ~n30895;
  assign n30897 = n3374 & ~n30896;
  assign n30898 = ~n25917 & ~n30897;
  assign n30899 = n3655 & ~n30898;
  assign n30900 = ~n19618 & ~n25905;
  assign n30901 = controllable_nhgrant0 & ~n30900;
  assign n30902 = ~n7118 & ~n30901;
  assign n30903 = ~n3281 & ~n30902;
  assign n30904 = ~n3281 & ~n30903;
  assign n30905 = ~n3378 & ~n30904;
  assign n30906 = ~n19575 & ~n30905;
  assign n30907 = n3492 & ~n30906;
  assign n30908 = n3492 & ~n30907;
  assign n30909 = n3485 & ~n30908;
  assign n30910 = n3485 & ~n30909;
  assign n30911 = ~n3374 & ~n30910;
  assign n30912 = ~n19694 & ~n30827;
  assign n30913 = controllable_nhgrant0 & ~n30912;
  assign n30914 = ~n19213 & ~n30913;
  assign n30915 = ~n3281 & ~n30914;
  assign n30916 = ~n3281 & ~n30915;
  assign n30917 = n3378 & ~n30916;
  assign n30918 = ~n19787 & ~n30844;
  assign n30919 = controllable_nhgrant0 & ~n30918;
  assign n30920 = ~n19255 & ~n30919;
  assign n30921 = ~n3281 & ~n30920;
  assign n30922 = ~n3281 & ~n30921;
  assign n30923 = ~n3378 & ~n30922;
  assign n30924 = ~n30917 & ~n30923;
  assign n30925 = n3492 & ~n30924;
  assign n30926 = n3492 & ~n30925;
  assign n30927 = n3485 & ~n30926;
  assign n30928 = n3485 & ~n30927;
  assign n30929 = ~n3476 & ~n30928;
  assign n30930 = ~n19949 & ~n30866;
  assign n30931 = controllable_nhgrant0 & ~n30930;
  assign n30932 = ~n19385 & ~n30931;
  assign n30933 = ~n3281 & ~n30932;
  assign n30934 = ~n3281 & ~n30933;
  assign n30935 = n3378 & ~n30934;
  assign n30936 = ~n20118 & ~n30883;
  assign n30937 = controllable_nhgrant0 & ~n30936;
  assign n30938 = ~n19515 & ~n30937;
  assign n30939 = ~n3281 & ~n30938;
  assign n30940 = ~n3281 & ~n30939;
  assign n30941 = ~n3378 & ~n30940;
  assign n30942 = ~n30935 & ~n30941;
  assign n30943 = n3492 & ~n30942;
  assign n30944 = ~n18151 & ~n30943;
  assign n30945 = n3485 & ~n30944;
  assign n30946 = ~n18150 & ~n30945;
  assign n30947 = n3476 & ~n30946;
  assign n30948 = ~n30929 & ~n30947;
  assign n30949 = n3374 & ~n30948;
  assign n30950 = ~n30911 & ~n30949;
  assign n30951 = ~n3655 & ~n30950;
  assign n30952 = ~n30899 & ~n30951;
  assign n30953 = n3652 & ~n30952;
  assign n30954 = ~n20148 & ~n30827;
  assign n30955 = controllable_nhgrant0 & ~n30954;
  assign n30956 = ~n19213 & ~n30955;
  assign n30957 = ~n3281 & ~n30956;
  assign n30958 = ~n3281 & ~n30957;
  assign n30959 = n3378 & ~n30958;
  assign n30960 = ~n20166 & ~n30844;
  assign n30961 = controllable_nhgrant0 & ~n30960;
  assign n30962 = ~n19255 & ~n30961;
  assign n30963 = ~n3281 & ~n30962;
  assign n30964 = ~n3281 & ~n30963;
  assign n30965 = ~n3378 & ~n30964;
  assign n30966 = ~n30959 & ~n30965;
  assign n30967 = n3492 & ~n30966;
  assign n30968 = n3492 & ~n30967;
  assign n30969 = n3485 & ~n30968;
  assign n30970 = n3485 & ~n30969;
  assign n30971 = ~n3476 & ~n30970;
  assign n30972 = ~n20194 & ~n30866;
  assign n30973 = controllable_nhgrant0 & ~n30972;
  assign n30974 = ~n19385 & ~n30973;
  assign n30975 = ~n3281 & ~n30974;
  assign n30976 = ~n3281 & ~n30975;
  assign n30977 = n3378 & ~n30976;
  assign n30978 = ~n20235 & ~n30883;
  assign n30979 = controllable_nhgrant0 & ~n30978;
  assign n30980 = ~n19515 & ~n30979;
  assign n30981 = ~n3281 & ~n30980;
  assign n30982 = ~n3281 & ~n30981;
  assign n30983 = ~n3378 & ~n30982;
  assign n30984 = ~n30977 & ~n30983;
  assign n30985 = n3492 & ~n30984;
  assign n30986 = n3492 & ~n30985;
  assign n30987 = n3485 & ~n30986;
  assign n30988 = n3485 & ~n30987;
  assign n30989 = n3476 & ~n30988;
  assign n30990 = ~n30971 & ~n30989;
  assign n30991 = n3374 & ~n30990;
  assign n30992 = ~n26031 & ~n30991;
  assign n30993 = n3655 & ~n30992;
  assign n30994 = ~n20269 & ~n25905;
  assign n30995 = controllable_nhgrant0 & ~n30994;
  assign n30996 = ~n7118 & ~n30995;
  assign n30997 = ~n3281 & ~n30996;
  assign n30998 = ~n3281 & ~n30997;
  assign n30999 = ~n3378 & ~n30998;
  assign n31000 = ~n19575 & ~n30999;
  assign n31001 = n3492 & ~n31000;
  assign n31002 = n3492 & ~n31001;
  assign n31003 = n3485 & ~n31002;
  assign n31004 = n3485 & ~n31003;
  assign n31005 = ~n3374 & ~n31004;
  assign n31006 = ~n20293 & ~n30827;
  assign n31007 = controllable_nhgrant0 & ~n31006;
  assign n31008 = ~n19213 & ~n31007;
  assign n31009 = ~n3281 & ~n31008;
  assign n31010 = ~n3281 & ~n31009;
  assign n31011 = n3378 & ~n31010;
  assign n31012 = ~n20340 & ~n30844;
  assign n31013 = controllable_nhgrant0 & ~n31012;
  assign n31014 = ~n19255 & ~n31013;
  assign n31015 = ~n3281 & ~n31014;
  assign n31016 = ~n3281 & ~n31015;
  assign n31017 = ~n3378 & ~n31016;
  assign n31018 = ~n31011 & ~n31017;
  assign n31019 = n3492 & ~n31018;
  assign n31020 = n3492 & ~n31019;
  assign n31021 = n3485 & ~n31020;
  assign n31022 = n3485 & ~n31021;
  assign n31023 = ~n3476 & ~n31022;
  assign n31024 = ~n20368 & ~n30866;
  assign n31025 = controllable_nhgrant0 & ~n31024;
  assign n31026 = ~n19385 & ~n31025;
  assign n31027 = ~n3281 & ~n31026;
  assign n31028 = ~n3281 & ~n31027;
  assign n31029 = n3378 & ~n31028;
  assign n31030 = ~n20425 & ~n30883;
  assign n31031 = controllable_nhgrant0 & ~n31030;
  assign n31032 = ~n19515 & ~n31031;
  assign n31033 = ~n3281 & ~n31032;
  assign n31034 = ~n3281 & ~n31033;
  assign n31035 = ~n3378 & ~n31034;
  assign n31036 = ~n31029 & ~n31035;
  assign n31037 = n3492 & ~n31036;
  assign n31038 = ~n18151 & ~n31037;
  assign n31039 = n3485 & ~n31038;
  assign n31040 = ~n18150 & ~n31039;
  assign n31041 = n3476 & ~n31040;
  assign n31042 = ~n31023 & ~n31041;
  assign n31043 = n3374 & ~n31042;
  assign n31044 = ~n31005 & ~n31043;
  assign n31045 = ~n3655 & ~n31044;
  assign n31046 = ~n30993 & ~n31045;
  assign n31047 = ~n3652 & ~n31046;
  assign n31048 = ~n30953 & ~n31047;
  assign n31049 = n3368 & ~n31048;
  assign n31050 = ~n30817 & ~n31049;
  assign n31051 = n3362 & ~n31050;
  assign n31052 = n3492 & ~n30610;
  assign n31053 = ~n3631 & ~n31052;
  assign n31054 = n3485 & ~n31053;
  assign n31055 = ~n3630 & ~n31054;
  assign n31056 = ~n3476 & ~n31055;
  assign n31057 = n3492 & ~n30638;
  assign n31058 = ~n3631 & ~n31057;
  assign n31059 = n3485 & ~n31058;
  assign n31060 = ~n26202 & ~n31059;
  assign n31061 = n3476 & ~n31060;
  assign n31062 = ~n31056 & ~n31061;
  assign n31063 = n3374 & ~n31062;
  assign n31064 = ~n26206 & ~n31063;
  assign n31065 = n3655 & ~n31064;
  assign n31066 = n3492 & ~n30654;
  assign n31067 = ~n3631 & ~n31066;
  assign n31068 = n3485 & ~n31067;
  assign n31069 = ~n3630 & ~n31068;
  assign n31070 = ~n3476 & ~n31069;
  assign n31071 = ~n20467 & ~n26297;
  assign n31072 = ~n3485 & ~n31071;
  assign n31073 = ~n18630 & ~n31066;
  assign n31074 = n3485 & ~n31073;
  assign n31075 = ~n31072 & ~n31074;
  assign n31076 = n3476 & ~n31075;
  assign n31077 = ~n31070 & ~n31076;
  assign n31078 = ~n3374 & ~n31077;
  assign n31079 = n3492 & ~n30678;
  assign n31080 = ~n3631 & ~n31079;
  assign n31081 = n3485 & ~n31080;
  assign n31082 = ~n3630 & ~n31081;
  assign n31083 = ~n3476 & ~n31082;
  assign n31084 = n3492 & ~n30696;
  assign n31085 = ~n18630 & ~n31084;
  assign n31086 = n3485 & ~n31085;
  assign n31087 = ~n31072 & ~n31086;
  assign n31088 = n3476 & ~n31087;
  assign n31089 = ~n31083 & ~n31088;
  assign n31090 = n3374 & ~n31089;
  assign n31091 = ~n31078 & ~n31090;
  assign n31092 = ~n3655 & ~n31091;
  assign n31093 = ~n31065 & ~n31092;
  assign n31094 = n3652 & ~n31093;
  assign n31095 = n3492 & ~n30726;
  assign n31096 = ~n3631 & ~n31095;
  assign n31097 = n3485 & ~n31096;
  assign n31098 = ~n3630 & ~n31097;
  assign n31099 = ~n3476 & ~n31098;
  assign n31100 = n3492 & ~n30744;
  assign n31101 = ~n3631 & ~n31100;
  assign n31102 = n3485 & ~n31101;
  assign n31103 = ~n26398 & ~n31102;
  assign n31104 = n3476 & ~n31103;
  assign n31105 = ~n31099 & ~n31104;
  assign n31106 = n3374 & ~n31105;
  assign n31107 = ~n26402 & ~n31106;
  assign n31108 = n3655 & ~n31107;
  assign n31109 = n3492 & ~n30760;
  assign n31110 = ~n3631 & ~n31109;
  assign n31111 = n3485 & ~n31110;
  assign n31112 = ~n3630 & ~n31111;
  assign n31113 = ~n3476 & ~n31112;
  assign n31114 = ~n20467 & ~n26437;
  assign n31115 = ~n3485 & ~n31114;
  assign n31116 = ~n18630 & ~n31109;
  assign n31117 = n3485 & ~n31116;
  assign n31118 = ~n31115 & ~n31117;
  assign n31119 = n3476 & ~n31118;
  assign n31120 = ~n31113 & ~n31119;
  assign n31121 = ~n3374 & ~n31120;
  assign n31122 = n3492 & ~n30784;
  assign n31123 = ~n3631 & ~n31122;
  assign n31124 = n3485 & ~n31123;
  assign n31125 = ~n3630 & ~n31124;
  assign n31126 = ~n3476 & ~n31125;
  assign n31127 = n3492 & ~n30802;
  assign n31128 = ~n18630 & ~n31127;
  assign n31129 = n3485 & ~n31128;
  assign n31130 = ~n31115 & ~n31129;
  assign n31131 = n3476 & ~n31130;
  assign n31132 = ~n31126 & ~n31131;
  assign n31133 = n3374 & ~n31132;
  assign n31134 = ~n31121 & ~n31133;
  assign n31135 = ~n3655 & ~n31134;
  assign n31136 = ~n31108 & ~n31135;
  assign n31137 = ~n3652 & ~n31136;
  assign n31138 = ~n31094 & ~n31137;
  assign n31139 = ~n3368 & ~n31138;
  assign n31140 = n3492 & ~n30849;
  assign n31141 = n3492 & ~n31140;
  assign n31142 = n3485 & ~n31141;
  assign n31143 = n3485 & ~n31142;
  assign n31144 = ~n3476 & ~n31143;
  assign n31145 = n3492 & ~n30888;
  assign n31146 = n3492 & ~n31145;
  assign n31147 = n3485 & ~n31146;
  assign n31148 = ~n26479 & ~n31147;
  assign n31149 = n3476 & ~n31148;
  assign n31150 = ~n31144 & ~n31149;
  assign n31151 = n3374 & ~n31150;
  assign n31152 = ~n26470 & ~n31151;
  assign n31153 = n3655 & ~n31152;
  assign n31154 = n3492 & ~n30904;
  assign n31155 = n3492 & ~n31154;
  assign n31156 = n3485 & ~n31155;
  assign n31157 = n3485 & ~n31156;
  assign n31158 = ~n3476 & ~n31157;
  assign n31159 = ~n8525 & ~n31156;
  assign n31160 = n3476 & ~n31159;
  assign n31161 = ~n31158 & ~n31160;
  assign n31162 = ~n3374 & ~n31161;
  assign n31163 = n3492 & ~n30922;
  assign n31164 = n3492 & ~n31163;
  assign n31165 = n3485 & ~n31164;
  assign n31166 = n3485 & ~n31165;
  assign n31167 = ~n3476 & ~n31166;
  assign n31168 = ~n20565 & ~n26504;
  assign n31169 = ~n3485 & ~n31168;
  assign n31170 = n3492 & ~n30940;
  assign n31171 = ~n18151 & ~n31170;
  assign n31172 = n3485 & ~n31171;
  assign n31173 = ~n31169 & ~n31172;
  assign n31174 = n3476 & ~n31173;
  assign n31175 = ~n31167 & ~n31174;
  assign n31176 = n3374 & ~n31175;
  assign n31177 = ~n31162 & ~n31176;
  assign n31178 = ~n3655 & ~n31177;
  assign n31179 = ~n31153 & ~n31178;
  assign n31180 = n3652 & ~n31179;
  assign n31181 = n3492 & ~n30964;
  assign n31182 = n3492 & ~n31181;
  assign n31183 = n3485 & ~n31182;
  assign n31184 = n3485 & ~n31183;
  assign n31185 = ~n3476 & ~n31184;
  assign n31186 = n3492 & ~n30982;
  assign n31187 = n3492 & ~n31186;
  assign n31188 = n3485 & ~n31187;
  assign n31189 = ~n26535 & ~n31188;
  assign n31190 = n3476 & ~n31189;
  assign n31191 = ~n31185 & ~n31190;
  assign n31192 = n3374 & ~n31191;
  assign n31193 = ~n26526 & ~n31192;
  assign n31194 = n3655 & ~n31193;
  assign n31195 = n3492 & ~n30998;
  assign n31196 = n3492 & ~n31195;
  assign n31197 = n3485 & ~n31196;
  assign n31198 = n3485 & ~n31197;
  assign n31199 = ~n3476 & ~n31198;
  assign n31200 = ~n8525 & ~n31197;
  assign n31201 = n3476 & ~n31200;
  assign n31202 = ~n31199 & ~n31201;
  assign n31203 = ~n3374 & ~n31202;
  assign n31204 = n3492 & ~n31016;
  assign n31205 = n3492 & ~n31204;
  assign n31206 = n3485 & ~n31205;
  assign n31207 = n3485 & ~n31206;
  assign n31208 = ~n3476 & ~n31207;
  assign n31209 = ~n20565 & ~n26560;
  assign n31210 = ~n3485 & ~n31209;
  assign n31211 = n3492 & ~n31034;
  assign n31212 = ~n18151 & ~n31211;
  assign n31213 = n3485 & ~n31212;
  assign n31214 = ~n31210 & ~n31213;
  assign n31215 = n3476 & ~n31214;
  assign n31216 = ~n31208 & ~n31215;
  assign n31217 = n3374 & ~n31216;
  assign n31218 = ~n31203 & ~n31217;
  assign n31219 = ~n3655 & ~n31218;
  assign n31220 = ~n31194 & ~n31219;
  assign n31221 = ~n3652 & ~n31220;
  assign n31222 = ~n31180 & ~n31221;
  assign n31223 = n3368 & ~n31222;
  assign n31224 = ~n31139 & ~n31223;
  assign n31225 = ~n3362 & ~n31224;
  assign n31226 = ~n31051 & ~n31225;
  assign n31227 = n3359 & ~n31226;
  assign n31228 = ~n26580 & ~n31059;
  assign n31229 = n3476 & ~n31228;
  assign n31230 = ~n31056 & ~n31229;
  assign n31231 = n3374 & ~n31230;
  assign n31232 = ~n26584 & ~n31231;
  assign n31233 = n3655 & ~n31232;
  assign n31234 = ~n26591 & ~n31074;
  assign n31235 = n3476 & ~n31234;
  assign n31236 = ~n31070 & ~n31235;
  assign n31237 = ~n3374 & ~n31236;
  assign n31238 = ~n26591 & ~n31086;
  assign n31239 = n3476 & ~n31238;
  assign n31240 = ~n31083 & ~n31239;
  assign n31241 = n3374 & ~n31240;
  assign n31242 = ~n31237 & ~n31241;
  assign n31243 = ~n3655 & ~n31242;
  assign n31244 = ~n31233 & ~n31243;
  assign n31245 = n3652 & ~n31244;
  assign n31246 = ~n26604 & ~n31102;
  assign n31247 = n3476 & ~n31246;
  assign n31248 = ~n31099 & ~n31247;
  assign n31249 = n3374 & ~n31248;
  assign n31250 = ~n26608 & ~n31249;
  assign n31251 = n3655 & ~n31250;
  assign n31252 = ~n26615 & ~n31117;
  assign n31253 = n3476 & ~n31252;
  assign n31254 = ~n31113 & ~n31253;
  assign n31255 = ~n3374 & ~n31254;
  assign n31256 = ~n26615 & ~n31129;
  assign n31257 = n3476 & ~n31256;
  assign n31258 = ~n31126 & ~n31257;
  assign n31259 = n3374 & ~n31258;
  assign n31260 = ~n31255 & ~n31259;
  assign n31261 = ~n3655 & ~n31260;
  assign n31262 = ~n31251 & ~n31261;
  assign n31263 = ~n3652 & ~n31262;
  assign n31264 = ~n31245 & ~n31263;
  assign n31265 = ~n3368 & ~n31264;
  assign n31266 = ~n26634 & ~n31147;
  assign n31267 = n3476 & ~n31266;
  assign n31268 = ~n31144 & ~n31267;
  assign n31269 = n3374 & ~n31268;
  assign n31270 = ~n26633 & ~n31269;
  assign n31271 = n3655 & ~n31270;
  assign n31272 = ~n8689 & ~n31156;
  assign n31273 = n3476 & ~n31272;
  assign n31274 = ~n31158 & ~n31273;
  assign n31275 = ~n3374 & ~n31274;
  assign n31276 = ~n26645 & ~n31172;
  assign n31277 = n3476 & ~n31276;
  assign n31278 = ~n31167 & ~n31277;
  assign n31279 = n3374 & ~n31278;
  assign n31280 = ~n31275 & ~n31279;
  assign n31281 = ~n3655 & ~n31280;
  assign n31282 = ~n31271 & ~n31281;
  assign n31283 = n3652 & ~n31282;
  assign n31284 = ~n26658 & ~n31188;
  assign n31285 = n3476 & ~n31284;
  assign n31286 = ~n31185 & ~n31285;
  assign n31287 = n3374 & ~n31286;
  assign n31288 = ~n26657 & ~n31287;
  assign n31289 = n3655 & ~n31288;
  assign n31290 = ~n8689 & ~n31197;
  assign n31291 = n3476 & ~n31290;
  assign n31292 = ~n31199 & ~n31291;
  assign n31293 = ~n3374 & ~n31292;
  assign n31294 = ~n26669 & ~n31213;
  assign n31295 = n3476 & ~n31294;
  assign n31296 = ~n31208 & ~n31295;
  assign n31297 = n3374 & ~n31296;
  assign n31298 = ~n31293 & ~n31297;
  assign n31299 = ~n3655 & ~n31298;
  assign n31300 = ~n31289 & ~n31299;
  assign n31301 = ~n3652 & ~n31300;
  assign n31302 = ~n31283 & ~n31301;
  assign n31303 = n3368 & ~n31302;
  assign n31304 = ~n31265 & ~n31303;
  assign n31305 = n3362 & ~n31304;
  assign n31306 = n3378 & ~n30610;
  assign n31307 = ~n26711 & ~n31306;
  assign n31308 = n3492 & ~n31307;
  assign n31309 = ~n3631 & ~n31308;
  assign n31310 = n3485 & ~n31309;
  assign n31311 = ~n3630 & ~n31310;
  assign n31312 = ~n3476 & ~n31311;
  assign n31313 = n3378 & ~n30638;
  assign n31314 = ~n26726 & ~n31313;
  assign n31315 = n3492 & ~n31314;
  assign n31316 = ~n26200 & ~n31315;
  assign n31317 = n3485 & ~n31316;
  assign n31318 = ~n26580 & ~n31317;
  assign n31319 = n3476 & ~n31318;
  assign n31320 = ~n31312 & ~n31319;
  assign n31321 = n3374 & ~n31320;
  assign n31322 = ~n26702 & ~n31321;
  assign n31323 = n3655 & ~n31322;
  assign n31324 = n3378 & ~n30654;
  assign n31325 = ~n26743 & ~n31324;
  assign n31326 = n3492 & ~n31325;
  assign n31327 = ~n3631 & ~n31326;
  assign n31328 = n3485 & ~n31327;
  assign n31329 = ~n3630 & ~n31328;
  assign n31330 = ~n3476 & ~n31329;
  assign n31331 = ~n26297 & ~n31326;
  assign n31332 = n3485 & ~n31331;
  assign n31333 = ~n26591 & ~n31332;
  assign n31334 = n3476 & ~n31333;
  assign n31335 = ~n31330 & ~n31334;
  assign n31336 = ~n3374 & ~n31335;
  assign n31337 = n3378 & ~n30678;
  assign n31338 = ~n26762 & ~n31337;
  assign n31339 = n3492 & ~n31338;
  assign n31340 = ~n3631 & ~n31339;
  assign n31341 = n3485 & ~n31340;
  assign n31342 = ~n3630 & ~n31341;
  assign n31343 = ~n3476 & ~n31342;
  assign n31344 = n3378 & ~n30696;
  assign n31345 = ~n26775 & ~n31344;
  assign n31346 = n3492 & ~n31345;
  assign n31347 = ~n26297 & ~n31346;
  assign n31348 = n3485 & ~n31347;
  assign n31349 = ~n26591 & ~n31348;
  assign n31350 = n3476 & ~n31349;
  assign n31351 = ~n31343 & ~n31350;
  assign n31352 = n3374 & ~n31351;
  assign n31353 = ~n31336 & ~n31352;
  assign n31354 = ~n3655 & ~n31353;
  assign n31355 = ~n31323 & ~n31354;
  assign n31356 = n3652 & ~n31355;
  assign n31357 = n3378 & ~n30726;
  assign n31358 = ~n26813 & ~n31357;
  assign n31359 = n3492 & ~n31358;
  assign n31360 = ~n3631 & ~n31359;
  assign n31361 = n3485 & ~n31360;
  assign n31362 = ~n3630 & ~n31361;
  assign n31363 = ~n3476 & ~n31362;
  assign n31364 = n3378 & ~n30744;
  assign n31365 = ~n26826 & ~n31364;
  assign n31366 = n3492 & ~n31365;
  assign n31367 = ~n26396 & ~n31366;
  assign n31368 = n3485 & ~n31367;
  assign n31369 = ~n26604 & ~n31368;
  assign n31370 = n3476 & ~n31369;
  assign n31371 = ~n31363 & ~n31370;
  assign n31372 = n3374 & ~n31371;
  assign n31373 = ~n26806 & ~n31372;
  assign n31374 = n3655 & ~n31373;
  assign n31375 = n3378 & ~n30760;
  assign n31376 = ~n26843 & ~n31375;
  assign n31377 = n3492 & ~n31376;
  assign n31378 = ~n3631 & ~n31377;
  assign n31379 = n3485 & ~n31378;
  assign n31380 = ~n3630 & ~n31379;
  assign n31381 = ~n3476 & ~n31380;
  assign n31382 = ~n26437 & ~n31377;
  assign n31383 = n3485 & ~n31382;
  assign n31384 = ~n26615 & ~n31383;
  assign n31385 = n3476 & ~n31384;
  assign n31386 = ~n31381 & ~n31385;
  assign n31387 = ~n3374 & ~n31386;
  assign n31388 = n3378 & ~n30784;
  assign n31389 = ~n26862 & ~n31388;
  assign n31390 = n3492 & ~n31389;
  assign n31391 = ~n3631 & ~n31390;
  assign n31392 = n3485 & ~n31391;
  assign n31393 = ~n3630 & ~n31392;
  assign n31394 = ~n3476 & ~n31393;
  assign n31395 = n3378 & ~n30802;
  assign n31396 = ~n26875 & ~n31395;
  assign n31397 = n3492 & ~n31396;
  assign n31398 = ~n26437 & ~n31397;
  assign n31399 = n3485 & ~n31398;
  assign n31400 = ~n26615 & ~n31399;
  assign n31401 = n3476 & ~n31400;
  assign n31402 = ~n31394 & ~n31401;
  assign n31403 = n3374 & ~n31402;
  assign n31404 = ~n31387 & ~n31403;
  assign n31405 = ~n3655 & ~n31404;
  assign n31406 = ~n31374 & ~n31405;
  assign n31407 = ~n3652 & ~n31406;
  assign n31408 = ~n31356 & ~n31407;
  assign n31409 = ~n3368 & ~n31408;
  assign n31410 = n3378 & ~n30849;
  assign n31411 = ~n26931 & ~n31410;
  assign n31412 = n3492 & ~n31411;
  assign n31413 = n3492 & ~n31412;
  assign n31414 = n3485 & ~n31413;
  assign n31415 = n3485 & ~n31414;
  assign n31416 = ~n3476 & ~n31415;
  assign n31417 = controllable_hmaster0 & ~n26943;
  assign n31418 = ~n27003 & ~n31417;
  assign n31419 = ~controllable_hmaster1 & ~n31418;
  assign n31420 = ~n27005 & ~n31419;
  assign n31421 = i_hlock3 & ~n31420;
  assign n31422 = controllable_hmaster0 & ~n26954;
  assign n31423 = ~n27012 & ~n31422;
  assign n31424 = ~controllable_hmaster1 & ~n31423;
  assign n31425 = ~n27014 & ~n31424;
  assign n31426 = ~i_hlock3 & ~n31425;
  assign n31427 = ~n31421 & ~n31426;
  assign n31428 = i_hbusreq3 & ~n31427;
  assign n31429 = controllable_hmaster0 & ~n26973;
  assign n31430 = ~n27033 & ~n31429;
  assign n31431 = ~controllable_hmaster1 & ~n31430;
  assign n31432 = ~n27028 & ~n31431;
  assign n31433 = i_hlock3 & ~n31432;
  assign n31434 = controllable_hmaster0 & ~n26990;
  assign n31435 = ~n27051 & ~n31434;
  assign n31436 = ~controllable_hmaster1 & ~n31435;
  assign n31437 = ~n27046 & ~n31436;
  assign n31438 = ~i_hlock3 & ~n31437;
  assign n31439 = ~n31433 & ~n31438;
  assign n31440 = ~i_hbusreq3 & ~n31439;
  assign n31441 = ~n31428 & ~n31440;
  assign n31442 = ~controllable_hmaster2 & ~n31441;
  assign n31443 = ~n30153 & ~n31442;
  assign n31444 = controllable_hgrant3 & ~n31443;
  assign n31445 = ~n20899 & ~n31444;
  assign n31446 = controllable_nhgrant0 & ~n31445;
  assign n31447 = ~n20915 & ~n31446;
  assign n31448 = ~n3281 & ~n31447;
  assign n31449 = ~n3281 & ~n31448;
  assign n31450 = n3378 & ~n31449;
  assign n31451 = ~n27144 & ~n31450;
  assign n31452 = n3492 & ~n31451;
  assign n31453 = ~n26477 & ~n31452;
  assign n31454 = n3485 & ~n31453;
  assign n31455 = ~n26634 & ~n31454;
  assign n31456 = n3476 & ~n31455;
  assign n31457 = ~n31416 & ~n31456;
  assign n31458 = n3374 & ~n31457;
  assign n31459 = ~n26909 & ~n31458;
  assign n31460 = n3655 & ~n31459;
  assign n31461 = n3378 & ~n30904;
  assign n31462 = ~n27161 & ~n31461;
  assign n31463 = n3492 & ~n31462;
  assign n31464 = n3492 & ~n31463;
  assign n31465 = n3485 & ~n31464;
  assign n31466 = n3485 & ~n31465;
  assign n31467 = ~n3476 & ~n31466;
  assign n31468 = ~n8523 & ~n31463;
  assign n31469 = n3485 & ~n31468;
  assign n31470 = ~n8689 & ~n31469;
  assign n31471 = n3476 & ~n31470;
  assign n31472 = ~n31467 & ~n31471;
  assign n31473 = ~n3374 & ~n31472;
  assign n31474 = n3378 & ~n30922;
  assign n31475 = ~n27180 & ~n31474;
  assign n31476 = n3492 & ~n31475;
  assign n31477 = n3492 & ~n31476;
  assign n31478 = n3485 & ~n31477;
  assign n31479 = n3485 & ~n31478;
  assign n31480 = ~n3476 & ~n31479;
  assign n31481 = ~n21079 & ~n31444;
  assign n31482 = controllable_nhgrant0 & ~n31481;
  assign n31483 = ~n20915 & ~n31482;
  assign n31484 = ~n3281 & ~n31483;
  assign n31485 = ~n3281 & ~n31484;
  assign n31486 = n3378 & ~n31485;
  assign n31487 = ~n27198 & ~n31486;
  assign n31488 = n3492 & ~n31487;
  assign n31489 = ~n26504 & ~n31488;
  assign n31490 = n3485 & ~n31489;
  assign n31491 = ~n26645 & ~n31490;
  assign n31492 = n3476 & ~n31491;
  assign n31493 = ~n31480 & ~n31492;
  assign n31494 = n3374 & ~n31493;
  assign n31495 = ~n31473 & ~n31494;
  assign n31496 = ~n3655 & ~n31495;
  assign n31497 = ~n31460 & ~n31496;
  assign n31498 = n3652 & ~n31497;
  assign n31499 = n3378 & ~n30964;
  assign n31500 = ~n27236 & ~n31499;
  assign n31501 = n3492 & ~n31500;
  assign n31502 = n3492 & ~n31501;
  assign n31503 = n3485 & ~n31502;
  assign n31504 = n3485 & ~n31503;
  assign n31505 = ~n3476 & ~n31504;
  assign n31506 = ~n21137 & ~n31444;
  assign n31507 = controllable_nhgrant0 & ~n31506;
  assign n31508 = ~n20915 & ~n31507;
  assign n31509 = ~n3281 & ~n31508;
  assign n31510 = ~n3281 & ~n31509;
  assign n31511 = n3378 & ~n31510;
  assign n31512 = ~n27254 & ~n31511;
  assign n31513 = n3492 & ~n31512;
  assign n31514 = ~n26533 & ~n31513;
  assign n31515 = n3485 & ~n31514;
  assign n31516 = ~n26658 & ~n31515;
  assign n31517 = n3476 & ~n31516;
  assign n31518 = ~n31505 & ~n31517;
  assign n31519 = n3374 & ~n31518;
  assign n31520 = ~n27229 & ~n31519;
  assign n31521 = n3655 & ~n31520;
  assign n31522 = n3378 & ~n30998;
  assign n31523 = ~n27271 & ~n31522;
  assign n31524 = n3492 & ~n31523;
  assign n31525 = n3492 & ~n31524;
  assign n31526 = n3485 & ~n31525;
  assign n31527 = n3485 & ~n31526;
  assign n31528 = ~n3476 & ~n31527;
  assign n31529 = ~n8523 & ~n31524;
  assign n31530 = n3485 & ~n31529;
  assign n31531 = ~n8689 & ~n31530;
  assign n31532 = n3476 & ~n31531;
  assign n31533 = ~n31528 & ~n31532;
  assign n31534 = ~n3374 & ~n31533;
  assign n31535 = n3378 & ~n31016;
  assign n31536 = ~n27290 & ~n31535;
  assign n31537 = n3492 & ~n31536;
  assign n31538 = n3492 & ~n31537;
  assign n31539 = n3485 & ~n31538;
  assign n31540 = n3485 & ~n31539;
  assign n31541 = ~n3476 & ~n31540;
  assign n31542 = ~n21222 & ~n31444;
  assign n31543 = controllable_nhgrant0 & ~n31542;
  assign n31544 = ~n20915 & ~n31543;
  assign n31545 = ~n3281 & ~n31544;
  assign n31546 = ~n3281 & ~n31545;
  assign n31547 = n3378 & ~n31546;
  assign n31548 = ~n27308 & ~n31547;
  assign n31549 = n3492 & ~n31548;
  assign n31550 = ~n26560 & ~n31549;
  assign n31551 = n3485 & ~n31550;
  assign n31552 = ~n26669 & ~n31551;
  assign n31553 = n3476 & ~n31552;
  assign n31554 = ~n31541 & ~n31553;
  assign n31555 = n3374 & ~n31554;
  assign n31556 = ~n31534 & ~n31555;
  assign n31557 = ~n3655 & ~n31556;
  assign n31558 = ~n31521 & ~n31557;
  assign n31559 = ~n3652 & ~n31558;
  assign n31560 = ~n31498 & ~n31559;
  assign n31561 = n3368 & ~n31560;
  assign n31562 = ~n31409 & ~n31561;
  assign n31563 = ~n3362 & ~n31562;
  assign n31564 = ~n31305 & ~n31563;
  assign n31565 = ~n3359 & ~n31564;
  assign n31566 = ~n31227 & ~n31565;
  assign n31567 = ~n3356 & ~n31566;
  assign n31568 = ~n30583 & ~n31567;
  assign n31569 = ~n3345 & ~n31568;
  assign n31570 = ~controllable_hmaster0 & ~n5478;
  assign n31571 = ~controllable_hmaster1 & ~n31570;
  assign n31572 = ~controllable_hmaster1 & ~n31571;
  assign n31573 = ~i_hbusreq3 & ~n31572;
  assign n31574 = ~n3914 & ~n31573;
  assign n31575 = ~controllable_hmaster2 & ~n31574;
  assign n31576 = ~controllable_hmaster2 & ~n31575;
  assign n31577 = controllable_hgrant3 & ~n31576;
  assign n31578 = ~n21316 & ~n31577;
  assign n31579 = controllable_nhgrant0 & ~n31578;
  assign n31580 = ~n21332 & ~n31579;
  assign n31581 = ~n3281 & ~n31580;
  assign n31582 = ~n3281 & ~n31581;
  assign n31583 = n3378 & ~n31582;
  assign n31584 = ~n21262 & ~n31575;
  assign n31585 = controllable_hgrant3 & ~n31584;
  assign n31586 = ~n21341 & ~n31585;
  assign n31587 = controllable_nhgrant0 & ~n31586;
  assign n31588 = ~n21347 & ~n31587;
  assign n31589 = ~n3281 & ~n31588;
  assign n31590 = ~n3950 & ~n31589;
  assign n31591 = ~n3378 & ~n31590;
  assign n31592 = ~n31583 & ~n31591;
  assign n31593 = n3492 & ~n31592;
  assign n31594 = ~n3493 & ~n31593;
  assign n31595 = n3485 & ~n31594;
  assign n31596 = ~n3486 & ~n31595;
  assign n31597 = ~n3476 & ~n31596;
  assign n31598 = ~n21383 & ~n31579;
  assign n31599 = ~n3281 & ~n31598;
  assign n31600 = ~n3281 & ~n31599;
  assign n31601 = n3378 & ~n31600;
  assign n31602 = ~n21443 & ~n31585;
  assign n31603 = controllable_nhgrant0 & ~n31602;
  assign n31604 = ~n21461 & ~n31603;
  assign n31605 = ~n3281 & ~n31604;
  assign n31606 = ~n4089 & ~n31605;
  assign n31607 = ~n3378 & ~n31606;
  assign n31608 = ~n31601 & ~n31607;
  assign n31609 = n3492 & ~n31608;
  assign n31610 = ~n21290 & ~n31609;
  assign n31611 = n3485 & ~n31610;
  assign n31612 = ~n21289 & ~n31611;
  assign n31613 = n3476 & ~n31612;
  assign n31614 = ~n31597 & ~n31613;
  assign n31615 = n3374 & ~n31614;
  assign n31616 = ~n21296 & ~n31615;
  assign n31617 = n3655 & ~n31616;
  assign n31618 = ~n21487 & ~n31577;
  assign n31619 = controllable_nhgrant0 & ~n31618;
  assign n31620 = ~n21332 & ~n31619;
  assign n31621 = ~n3281 & ~n31620;
  assign n31622 = ~n3281 & ~n31621;
  assign n31623 = n3378 & ~n31622;
  assign n31624 = ~n21495 & ~n31585;
  assign n31625 = controllable_nhgrant0 & ~n31624;
  assign n31626 = ~n21347 & ~n31625;
  assign n31627 = ~n3281 & ~n31626;
  assign n31628 = ~n3950 & ~n31627;
  assign n31629 = ~n3378 & ~n31628;
  assign n31630 = ~n31623 & ~n31629;
  assign n31631 = n3492 & ~n31630;
  assign n31632 = ~n3493 & ~n31631;
  assign n31633 = n3485 & ~n31632;
  assign n31634 = ~n3486 & ~n31633;
  assign n31635 = ~n3476 & ~n31634;
  assign n31636 = ~n21383 & ~n31619;
  assign n31637 = ~n3281 & ~n31636;
  assign n31638 = ~n3281 & ~n31637;
  assign n31639 = n3378 & ~n31638;
  assign n31640 = ~n21540 & ~n31585;
  assign n31641 = controllable_nhgrant0 & ~n31640;
  assign n31642 = ~n21461 & ~n31641;
  assign n31643 = ~n3281 & ~n31642;
  assign n31644 = ~n4089 & ~n31643;
  assign n31645 = ~n3378 & ~n31644;
  assign n31646 = ~n31639 & ~n31645;
  assign n31647 = n3492 & ~n31646;
  assign n31648 = ~n21290 & ~n31647;
  assign n31649 = n3485 & ~n31648;
  assign n31650 = ~n21289 & ~n31649;
  assign n31651 = n3476 & ~n31650;
  assign n31652 = ~n31635 & ~n31651;
  assign n31653 = n3374 & ~n31652;
  assign n31654 = ~n21296 & ~n31653;
  assign n31655 = ~n3655 & ~n31654;
  assign n31656 = ~n31617 & ~n31655;
  assign n31657 = n3652 & ~n31656;
  assign n31658 = ~n21570 & ~n31577;
  assign n31659 = controllable_nhgrant0 & ~n31658;
  assign n31660 = ~n21332 & ~n31659;
  assign n31661 = ~n3281 & ~n31660;
  assign n31662 = ~n3281 & ~n31661;
  assign n31663 = n3378 & ~n31662;
  assign n31664 = ~n21578 & ~n31585;
  assign n31665 = controllable_nhgrant0 & ~n31664;
  assign n31666 = ~n21347 & ~n31665;
  assign n31667 = ~n3281 & ~n31666;
  assign n31668 = ~n3950 & ~n31667;
  assign n31669 = ~n3378 & ~n31668;
  assign n31670 = ~n31663 & ~n31669;
  assign n31671 = n3492 & ~n31670;
  assign n31672 = ~n3493 & ~n31671;
  assign n31673 = n3485 & ~n31672;
  assign n31674 = ~n3486 & ~n31673;
  assign n31675 = ~n3476 & ~n31674;
  assign n31676 = ~n21383 & ~n31659;
  assign n31677 = ~n3281 & ~n31676;
  assign n31678 = ~n3281 & ~n31677;
  assign n31679 = n3378 & ~n31678;
  assign n31680 = ~n21609 & ~n31585;
  assign n31681 = controllable_nhgrant0 & ~n31680;
  assign n31682 = ~n21461 & ~n31681;
  assign n31683 = ~n3281 & ~n31682;
  assign n31684 = ~n4089 & ~n31683;
  assign n31685 = ~n3378 & ~n31684;
  assign n31686 = ~n31679 & ~n31685;
  assign n31687 = n3492 & ~n31686;
  assign n31688 = ~n21290 & ~n31687;
  assign n31689 = n3485 & ~n31688;
  assign n31690 = ~n21289 & ~n31689;
  assign n31691 = n3476 & ~n31690;
  assign n31692 = ~n31675 & ~n31691;
  assign n31693 = n3374 & ~n31692;
  assign n31694 = ~n21296 & ~n31693;
  assign n31695 = n3655 & ~n31694;
  assign n31696 = ~n21637 & ~n31577;
  assign n31697 = controllable_nhgrant0 & ~n31696;
  assign n31698 = ~n21332 & ~n31697;
  assign n31699 = ~n3281 & ~n31698;
  assign n31700 = ~n3281 & ~n31699;
  assign n31701 = n3378 & ~n31700;
  assign n31702 = ~n21645 & ~n31585;
  assign n31703 = controllable_nhgrant0 & ~n31702;
  assign n31704 = ~n21347 & ~n31703;
  assign n31705 = ~n3281 & ~n31704;
  assign n31706 = ~n3950 & ~n31705;
  assign n31707 = ~n3378 & ~n31706;
  assign n31708 = ~n31701 & ~n31707;
  assign n31709 = n3492 & ~n31708;
  assign n31710 = ~n3493 & ~n31709;
  assign n31711 = n3485 & ~n31710;
  assign n31712 = ~n3486 & ~n31711;
  assign n31713 = ~n3476 & ~n31712;
  assign n31714 = ~n21383 & ~n31697;
  assign n31715 = ~n3281 & ~n31714;
  assign n31716 = ~n3281 & ~n31715;
  assign n31717 = n3378 & ~n31716;
  assign n31718 = ~n21676 & ~n31585;
  assign n31719 = controllable_nhgrant0 & ~n31718;
  assign n31720 = ~n21461 & ~n31719;
  assign n31721 = ~n3281 & ~n31720;
  assign n31722 = ~n4089 & ~n31721;
  assign n31723 = ~n3378 & ~n31722;
  assign n31724 = ~n31717 & ~n31723;
  assign n31725 = n3492 & ~n31724;
  assign n31726 = ~n21290 & ~n31725;
  assign n31727 = n3485 & ~n31726;
  assign n31728 = ~n21289 & ~n31727;
  assign n31729 = n3476 & ~n31728;
  assign n31730 = ~n31713 & ~n31729;
  assign n31731 = n3374 & ~n31730;
  assign n31732 = ~n21296 & ~n31731;
  assign n31733 = ~n3655 & ~n31732;
  assign n31734 = ~n31695 & ~n31733;
  assign n31735 = ~n3652 & ~n31734;
  assign n31736 = ~n31657 & ~n31735;
  assign n31737 = ~n3368 & ~n31736;
  assign n31738 = ~controllable_hmaster2 & ~n4614;
  assign n31739 = ~controllable_hmaster2 & ~n31738;
  assign n31740 = controllable_hgrant3 & ~n31739;
  assign n31741 = ~n21702 & ~n31740;
  assign n31742 = controllable_nhgrant0 & ~n31741;
  assign n31743 = ~n21712 & ~n31742;
  assign n31744 = ~n3281 & ~n31743;
  assign n31745 = ~n3281 & ~n31744;
  assign n31746 = n3492 & ~n31745;
  assign n31747 = n3492 & ~n31746;
  assign n31748 = n3485 & ~n31747;
  assign n31749 = n3485 & ~n31748;
  assign n31750 = ~n3476 & ~n31749;
  assign n31751 = ~n21740 & ~n31742;
  assign n31752 = ~n3281 & ~n31751;
  assign n31753 = ~n3281 & ~n31752;
  assign n31754 = n3492 & ~n31753;
  assign n31755 = ~n21722 & ~n31754;
  assign n31756 = n3485 & ~n31755;
  assign n31757 = ~n21721 & ~n31756;
  assign n31758 = n3476 & ~n31757;
  assign n31759 = ~n31750 & ~n31758;
  assign n31760 = n3374 & ~n31759;
  assign n31761 = n3374 & ~n31760;
  assign n31762 = n3655 & ~n31761;
  assign n31763 = ~n21758 & ~n31740;
  assign n31764 = controllable_nhgrant0 & ~n31763;
  assign n31765 = ~n21712 & ~n31764;
  assign n31766 = ~n3281 & ~n31765;
  assign n31767 = ~n3281 & ~n31766;
  assign n31768 = n3492 & ~n31767;
  assign n31769 = n3492 & ~n31768;
  assign n31770 = n3485 & ~n31769;
  assign n31771 = n3485 & ~n31770;
  assign n31772 = ~n3476 & ~n31771;
  assign n31773 = ~n21740 & ~n31764;
  assign n31774 = ~n3281 & ~n31773;
  assign n31775 = ~n3281 & ~n31774;
  assign n31776 = n3492 & ~n31775;
  assign n31777 = ~n21722 & ~n31776;
  assign n31778 = n3485 & ~n31777;
  assign n31779 = ~n21721 & ~n31778;
  assign n31780 = n3476 & ~n31779;
  assign n31781 = ~n31772 & ~n31780;
  assign n31782 = n3374 & ~n31781;
  assign n31783 = n3374 & ~n31782;
  assign n31784 = ~n3655 & ~n31783;
  assign n31785 = ~n31762 & ~n31784;
  assign n31786 = n3652 & ~n31785;
  assign n31787 = ~n21788 & ~n31740;
  assign n31788 = controllable_nhgrant0 & ~n31787;
  assign n31789 = ~n21712 & ~n31788;
  assign n31790 = ~n3281 & ~n31789;
  assign n31791 = ~n3281 & ~n31790;
  assign n31792 = n3492 & ~n31791;
  assign n31793 = n3492 & ~n31792;
  assign n31794 = n3485 & ~n31793;
  assign n31795 = n3485 & ~n31794;
  assign n31796 = ~n3476 & ~n31795;
  assign n31797 = ~n21740 & ~n31788;
  assign n31798 = ~n3281 & ~n31797;
  assign n31799 = ~n3281 & ~n31798;
  assign n31800 = n3492 & ~n31799;
  assign n31801 = ~n21722 & ~n31800;
  assign n31802 = n3485 & ~n31801;
  assign n31803 = ~n21721 & ~n31802;
  assign n31804 = n3476 & ~n31803;
  assign n31805 = ~n31796 & ~n31804;
  assign n31806 = n3374 & ~n31805;
  assign n31807 = n3374 & ~n31806;
  assign n31808 = n3655 & ~n31807;
  assign n31809 = ~n21816 & ~n31740;
  assign n31810 = controllable_nhgrant0 & ~n31809;
  assign n31811 = ~n21712 & ~n31810;
  assign n31812 = ~n3281 & ~n31811;
  assign n31813 = ~n3281 & ~n31812;
  assign n31814 = n3492 & ~n31813;
  assign n31815 = n3492 & ~n31814;
  assign n31816 = n3485 & ~n31815;
  assign n31817 = n3485 & ~n31816;
  assign n31818 = ~n3476 & ~n31817;
  assign n31819 = ~n21740 & ~n31810;
  assign n31820 = ~n3281 & ~n31819;
  assign n31821 = ~n3281 & ~n31820;
  assign n31822 = n3492 & ~n31821;
  assign n31823 = ~n21722 & ~n31822;
  assign n31824 = n3485 & ~n31823;
  assign n31825 = ~n21721 & ~n31824;
  assign n31826 = n3476 & ~n31825;
  assign n31827 = ~n31818 & ~n31826;
  assign n31828 = n3374 & ~n31827;
  assign n31829 = n3374 & ~n31828;
  assign n31830 = ~n3655 & ~n31829;
  assign n31831 = ~n31808 & ~n31830;
  assign n31832 = ~n3652 & ~n31831;
  assign n31833 = ~n31786 & ~n31832;
  assign n31834 = n3368 & ~n31833;
  assign n31835 = ~n31737 & ~n31834;
  assign n31836 = ~n3362 & ~n31835;
  assign n31837 = ~n3362 & ~n31836;
  assign n31838 = ~n3359 & ~n31837;
  assign n31839 = ~n3359 & ~n31838;
  assign n31840 = n3356 & ~n31839;
  assign n31841 = ~n3697 & ~n5191;
  assign n31842 = ~controllable_hmaster1 & ~n31841;
  assign n31843 = ~n5190 & ~n31842;
  assign n31844 = ~i_hbusreq3 & ~n31843;
  assign n31845 = ~n5195 & ~n31844;
  assign n31846 = controllable_hmaster2 & ~n31845;
  assign n31847 = ~n25647 & ~n31846;
  assign n31848 = controllable_hgrant3 & ~n31847;
  assign n31849 = ~n21857 & ~n31848;
  assign n31850 = controllable_nhgrant0 & ~n31849;
  assign n31851 = ~n8785 & ~n31850;
  assign n31852 = ~n3281 & ~n31851;
  assign n31853 = ~n3783 & ~n31852;
  assign n31854 = ~n3378 & ~n31853;
  assign n31855 = ~n21849 & ~n31854;
  assign n31856 = n3492 & ~n31855;
  assign n31857 = ~n3631 & ~n31856;
  assign n31858 = n3485 & ~n31857;
  assign n31859 = ~n3630 & ~n31858;
  assign n31860 = ~n3476 & ~n31859;
  assign n31861 = ~n8309 & ~n31856;
  assign n31862 = n3485 & ~n31861;
  assign n31863 = ~n8639 & ~n31862;
  assign n31864 = n3476 & ~n31863;
  assign n31865 = ~n31860 & ~n31864;
  assign n31866 = ~n3374 & ~n31865;
  assign n31867 = ~n3975 & ~n5262;
  assign n31868 = i_hbusreq3 & ~n31867;
  assign n31869 = ~n4913 & ~n5478;
  assign n31870 = ~controllable_hmaster1 & ~n31869;
  assign n31871 = ~n5379 & ~n31870;
  assign n31872 = ~i_hbusreq3 & ~n31871;
  assign n31873 = ~n31868 & ~n31872;
  assign n31874 = ~controllable_hmaster2 & ~n31873;
  assign n31875 = ~n8808 & ~n31874;
  assign n31876 = controllable_hgrant3 & ~n31875;
  assign n31877 = ~n21919 & ~n31876;
  assign n31878 = controllable_nhgrant0 & ~n31877;
  assign n31879 = ~n8902 & ~n31878;
  assign n31880 = ~n3281 & ~n31879;
  assign n31881 = ~n3950 & ~n31880;
  assign n31882 = n3378 & ~n31881;
  assign n31883 = ~n3935 & ~n5191;
  assign n31884 = ~controllable_hmaster1 & ~n31883;
  assign n31885 = ~n5190 & ~n31884;
  assign n31886 = ~i_hbusreq3 & ~n31885;
  assign n31887 = ~n5495 & ~n31886;
  assign n31888 = controllable_hmaster2 & ~n31887;
  assign n31889 = ~n25682 & ~n31888;
  assign n31890 = controllable_hgrant3 & ~n31889;
  assign n31891 = ~n21943 & ~n31890;
  assign n31892 = controllable_nhgrant0 & ~n31891;
  assign n31893 = ~n8902 & ~n31892;
  assign n31894 = ~n3281 & ~n31893;
  assign n31895 = ~n3950 & ~n31894;
  assign n31896 = ~n3378 & ~n31895;
  assign n31897 = ~n31882 & ~n31896;
  assign n31898 = n3492 & ~n31897;
  assign n31899 = ~n3631 & ~n31898;
  assign n31900 = n3485 & ~n31899;
  assign n31901 = ~n3630 & ~n31900;
  assign n31902 = ~n3476 & ~n31901;
  assign n31903 = ~n5590 & ~n5766;
  assign n31904 = i_hbusreq3 & ~n31903;
  assign n31905 = ~controllable_hgrant2 & ~n22382;
  assign n31906 = ~n5461 & ~n31905;
  assign n31907 = ~controllable_hmaster0 & ~n31906;
  assign n31908 = ~n5839 & ~n31907;
  assign n31909 = ~controllable_hmaster1 & ~n31908;
  assign n31910 = ~n5838 & ~n31909;
  assign n31911 = ~i_hbusreq3 & ~n31910;
  assign n31912 = ~n31904 & ~n31911;
  assign n31913 = ~controllable_hmaster2 & ~n31912;
  assign n31914 = ~n8933 & ~n31913;
  assign n31915 = controllable_hgrant3 & ~n31914;
  assign n31916 = ~n22015 & ~n31915;
  assign n31917 = controllable_nhgrant0 & ~n31916;
  assign n31918 = ~n9096 & ~n31917;
  assign n31919 = ~n3281 & ~n31918;
  assign n31920 = ~n4089 & ~n31919;
  assign n31921 = n3378 & ~n31920;
  assign n31922 = ~controllable_hgrant2 & ~n22410;
  assign n31923 = ~n3410 & ~n31922;
  assign n31924 = controllable_hmaster1 & ~n31923;
  assign n31925 = controllable_hmaster0 & ~n31923;
  assign n31926 = ~n9086 & ~n31925;
  assign n31927 = ~controllable_hmaster1 & ~n31926;
  assign n31928 = ~n31924 & ~n31927;
  assign n31929 = ~i_hbusreq3 & ~n31928;
  assign n31930 = ~n6013 & ~n31929;
  assign n31931 = controllable_hmaster2 & ~n31930;
  assign n31932 = ~n25724 & ~n31931;
  assign n31933 = controllable_hgrant3 & ~n31932;
  assign n31934 = ~n22077 & ~n31933;
  assign n31935 = controllable_nhgrant0 & ~n31934;
  assign n31936 = ~n9096 & ~n31935;
  assign n31937 = ~n3281 & ~n31936;
  assign n31938 = ~n4089 & ~n31937;
  assign n31939 = ~n3378 & ~n31938;
  assign n31940 = ~n31921 & ~n31939;
  assign n31941 = n3492 & ~n31940;
  assign n31942 = ~n8309 & ~n31941;
  assign n31943 = n3485 & ~n31942;
  assign n31944 = ~n8639 & ~n31943;
  assign n31945 = n3476 & ~n31944;
  assign n31946 = ~n31902 & ~n31945;
  assign n31947 = n3374 & ~n31946;
  assign n31948 = ~n31866 & ~n31947;
  assign n31949 = n3655 & ~n31948;
  assign n31950 = ~n22101 & ~n31848;
  assign n31951 = controllable_nhgrant0 & ~n31950;
  assign n31952 = ~n8785 & ~n31951;
  assign n31953 = ~n3281 & ~n31952;
  assign n31954 = ~n3783 & ~n31953;
  assign n31955 = ~n3378 & ~n31954;
  assign n31956 = ~n21849 & ~n31955;
  assign n31957 = n3492 & ~n31956;
  assign n31958 = ~n3631 & ~n31957;
  assign n31959 = n3485 & ~n31958;
  assign n31960 = ~n3630 & ~n31959;
  assign n31961 = ~n3476 & ~n31960;
  assign n31962 = ~n8309 & ~n31957;
  assign n31963 = n3485 & ~n31962;
  assign n31964 = ~n8639 & ~n31963;
  assign n31965 = n3476 & ~n31964;
  assign n31966 = ~n31961 & ~n31965;
  assign n31967 = ~n3374 & ~n31966;
  assign n31968 = ~n22131 & ~n31876;
  assign n31969 = controllable_nhgrant0 & ~n31968;
  assign n31970 = ~n8902 & ~n31969;
  assign n31971 = ~n3281 & ~n31970;
  assign n31972 = ~n3950 & ~n31971;
  assign n31973 = n3378 & ~n31972;
  assign n31974 = ~n22155 & ~n31890;
  assign n31975 = controllable_nhgrant0 & ~n31974;
  assign n31976 = ~n8902 & ~n31975;
  assign n31977 = ~n3281 & ~n31976;
  assign n31978 = ~n3950 & ~n31977;
  assign n31979 = ~n3378 & ~n31978;
  assign n31980 = ~n31973 & ~n31979;
  assign n31981 = n3492 & ~n31980;
  assign n31982 = ~n3631 & ~n31981;
  assign n31983 = n3485 & ~n31982;
  assign n31984 = ~n3630 & ~n31983;
  assign n31985 = ~n3476 & ~n31984;
  assign n31986 = ~n22196 & ~n31915;
  assign n31987 = controllable_nhgrant0 & ~n31986;
  assign n31988 = ~n9096 & ~n31987;
  assign n31989 = ~n3281 & ~n31988;
  assign n31990 = ~n4089 & ~n31989;
  assign n31991 = n3378 & ~n31990;
  assign n31992 = ~n22273 & ~n31933;
  assign n31993 = controllable_nhgrant0 & ~n31992;
  assign n31994 = ~n9096 & ~n31993;
  assign n31995 = ~n3281 & ~n31994;
  assign n31996 = ~n4089 & ~n31995;
  assign n31997 = ~n3378 & ~n31996;
  assign n31998 = ~n31991 & ~n31997;
  assign n31999 = n3492 & ~n31998;
  assign n32000 = ~n8309 & ~n31999;
  assign n32001 = n3485 & ~n32000;
  assign n32002 = ~n8639 & ~n32001;
  assign n32003 = n3476 & ~n32002;
  assign n32004 = ~n31985 & ~n32003;
  assign n32005 = n3374 & ~n32004;
  assign n32006 = ~n31967 & ~n32005;
  assign n32007 = ~n3655 & ~n32006;
  assign n32008 = ~n31949 & ~n32007;
  assign n32009 = n3652 & ~n32008;
  assign n32010 = ~n22299 & ~n31848;
  assign n32011 = controllable_nhgrant0 & ~n32010;
  assign n32012 = ~n8785 & ~n32011;
  assign n32013 = ~n3281 & ~n32012;
  assign n32014 = ~n3783 & ~n32013;
  assign n32015 = ~n3378 & ~n32014;
  assign n32016 = ~n21849 & ~n32015;
  assign n32017 = n3492 & ~n32016;
  assign n32018 = ~n3631 & ~n32017;
  assign n32019 = n3485 & ~n32018;
  assign n32020 = ~n3630 & ~n32019;
  assign n32021 = ~n3476 & ~n32020;
  assign n32022 = ~n8309 & ~n32017;
  assign n32023 = n3485 & ~n32022;
  assign n32024 = ~n8639 & ~n32023;
  assign n32025 = n3476 & ~n32024;
  assign n32026 = ~n32021 & ~n32025;
  assign n32027 = ~n3374 & ~n32026;
  assign n32028 = ~n22329 & ~n31876;
  assign n32029 = controllable_nhgrant0 & ~n32028;
  assign n32030 = ~n8902 & ~n32029;
  assign n32031 = ~n3281 & ~n32030;
  assign n32032 = ~n3950 & ~n32031;
  assign n32033 = n3378 & ~n32032;
  assign n32034 = ~n22353 & ~n31890;
  assign n32035 = controllable_nhgrant0 & ~n32034;
  assign n32036 = ~n8902 & ~n32035;
  assign n32037 = ~n3281 & ~n32036;
  assign n32038 = ~n3950 & ~n32037;
  assign n32039 = ~n3378 & ~n32038;
  assign n32040 = ~n32033 & ~n32039;
  assign n32041 = n3492 & ~n32040;
  assign n32042 = ~n3631 & ~n32041;
  assign n32043 = n3485 & ~n32042;
  assign n32044 = ~n3630 & ~n32043;
  assign n32045 = ~n3476 & ~n32044;
  assign n32046 = ~n22393 & ~n31915;
  assign n32047 = controllable_nhgrant0 & ~n32046;
  assign n32048 = ~n9096 & ~n32047;
  assign n32049 = ~n3281 & ~n32048;
  assign n32050 = ~n4089 & ~n32049;
  assign n32051 = n3378 & ~n32050;
  assign n32052 = ~n22442 & ~n31933;
  assign n32053 = controllable_nhgrant0 & ~n32052;
  assign n32054 = ~n9096 & ~n32053;
  assign n32055 = ~n3281 & ~n32054;
  assign n32056 = ~n4089 & ~n32055;
  assign n32057 = ~n3378 & ~n32056;
  assign n32058 = ~n32051 & ~n32057;
  assign n32059 = n3492 & ~n32058;
  assign n32060 = ~n8309 & ~n32059;
  assign n32061 = n3485 & ~n32060;
  assign n32062 = ~n8639 & ~n32061;
  assign n32063 = n3476 & ~n32062;
  assign n32064 = ~n32045 & ~n32063;
  assign n32065 = n3374 & ~n32064;
  assign n32066 = ~n32027 & ~n32065;
  assign n32067 = n3655 & ~n32066;
  assign n32068 = ~n22466 & ~n31848;
  assign n32069 = controllable_nhgrant0 & ~n32068;
  assign n32070 = ~n8785 & ~n32069;
  assign n32071 = ~n3281 & ~n32070;
  assign n32072 = ~n3783 & ~n32071;
  assign n32073 = ~n3378 & ~n32072;
  assign n32074 = ~n21849 & ~n32073;
  assign n32075 = n3492 & ~n32074;
  assign n32076 = ~n3631 & ~n32075;
  assign n32077 = n3485 & ~n32076;
  assign n32078 = ~n3630 & ~n32077;
  assign n32079 = ~n3476 & ~n32078;
  assign n32080 = ~n8309 & ~n32075;
  assign n32081 = n3485 & ~n32080;
  assign n32082 = ~n8639 & ~n32081;
  assign n32083 = n3476 & ~n32082;
  assign n32084 = ~n32079 & ~n32083;
  assign n32085 = ~n3374 & ~n32084;
  assign n32086 = ~n22496 & ~n31876;
  assign n32087 = controllable_nhgrant0 & ~n32086;
  assign n32088 = ~n8902 & ~n32087;
  assign n32089 = ~n3281 & ~n32088;
  assign n32090 = ~n3950 & ~n32089;
  assign n32091 = n3378 & ~n32090;
  assign n32092 = ~n22520 & ~n31890;
  assign n32093 = controllable_nhgrant0 & ~n32092;
  assign n32094 = ~n8902 & ~n32093;
  assign n32095 = ~n3281 & ~n32094;
  assign n32096 = ~n3950 & ~n32095;
  assign n32097 = ~n3378 & ~n32096;
  assign n32098 = ~n32091 & ~n32097;
  assign n32099 = n3492 & ~n32098;
  assign n32100 = ~n3631 & ~n32099;
  assign n32101 = n3485 & ~n32100;
  assign n32102 = ~n3630 & ~n32101;
  assign n32103 = ~n3476 & ~n32102;
  assign n32104 = ~n22547 & ~n31915;
  assign n32105 = controllable_nhgrant0 & ~n32104;
  assign n32106 = ~n9096 & ~n32105;
  assign n32107 = ~n3281 & ~n32106;
  assign n32108 = ~n4089 & ~n32107;
  assign n32109 = n3378 & ~n32108;
  assign n32110 = ~n22584 & ~n31933;
  assign n32111 = controllable_nhgrant0 & ~n32110;
  assign n32112 = ~n9096 & ~n32111;
  assign n32113 = ~n3281 & ~n32112;
  assign n32114 = ~n4089 & ~n32113;
  assign n32115 = ~n3378 & ~n32114;
  assign n32116 = ~n32109 & ~n32115;
  assign n32117 = n3492 & ~n32116;
  assign n32118 = ~n8309 & ~n32117;
  assign n32119 = n3485 & ~n32118;
  assign n32120 = ~n8639 & ~n32119;
  assign n32121 = n3476 & ~n32120;
  assign n32122 = ~n32103 & ~n32121;
  assign n32123 = n3374 & ~n32122;
  assign n32124 = ~n32085 & ~n32123;
  assign n32125 = ~n3655 & ~n32124;
  assign n32126 = ~n32067 & ~n32125;
  assign n32127 = ~n3652 & ~n32126;
  assign n32128 = ~n32009 & ~n32127;
  assign n32129 = ~n3368 & ~n32128;
  assign n32130 = controllable_hmaster1 & ~n22728;
  assign n32131 = controllable_hmaster0 & ~n22729;
  assign n32132 = ~controllable_hmaster1 & ~n32131;
  assign n32133 = ~n32130 & ~n32132;
  assign n32134 = ~i_hbusreq3 & ~n32133;
  assign n32135 = ~n7108 & ~n32134;
  assign n32136 = controllable_hmaster2 & ~n32135;
  assign n32137 = controllable_hmaster2 & ~n32136;
  assign n32138 = controllable_hgrant3 & ~n32137;
  assign n32139 = ~n22643 & ~n32138;
  assign n32140 = controllable_nhgrant0 & ~n32139;
  assign n32141 = ~n9753 & ~n32140;
  assign n32142 = ~n3281 & ~n32141;
  assign n32143 = ~n3281 & ~n32142;
  assign n32144 = ~n3378 & ~n32143;
  assign n32145 = ~n22618 & ~n32144;
  assign n32146 = n3492 & ~n32145;
  assign n32147 = n3492 & ~n32146;
  assign n32148 = n3485 & ~n32147;
  assign n32149 = n3485 & ~n32148;
  assign n32150 = ~n3374 & ~n32149;
  assign n32151 = ~n5262 & ~n7154;
  assign n32152 = i_hbusreq3 & ~n32151;
  assign n32153 = ~n4611 & ~n9700;
  assign n32154 = ~controllable_hmaster1 & ~n32153;
  assign n32155 = ~n9782 & ~n32154;
  assign n32156 = ~i_hbusreq3 & ~n32155;
  assign n32157 = ~n32152 & ~n32156;
  assign n32158 = ~controllable_hmaster2 & ~n32157;
  assign n32159 = ~n9773 & ~n32158;
  assign n32160 = controllable_hgrant3 & ~n32159;
  assign n32161 = ~n22695 & ~n32160;
  assign n32162 = controllable_nhgrant0 & ~n32161;
  assign n32163 = ~n9861 & ~n32162;
  assign n32164 = ~n3281 & ~n32163;
  assign n32165 = ~n3281 & ~n32164;
  assign n32166 = n3378 & ~n32165;
  assign n32167 = ~i_hbusreq3 & ~n22728;
  assign n32168 = ~n5495 & ~n32167;
  assign n32169 = controllable_hmaster2 & ~n32168;
  assign n32170 = ~n7196 & ~n25671;
  assign n32171 = i_hbusreq3 & ~n32170;
  assign n32172 = ~controllable_hmaster0 & ~n22728;
  assign n32173 = ~n22635 & ~n32172;
  assign n32174 = controllable_hmaster1 & ~n32173;
  assign n32175 = ~n4611 & ~n22729;
  assign n32176 = ~controllable_hmaster1 & ~n32175;
  assign n32177 = ~n32174 & ~n32176;
  assign n32178 = ~i_hbusreq3 & ~n32177;
  assign n32179 = ~n32171 & ~n32178;
  assign n32180 = ~controllable_hmaster2 & ~n32179;
  assign n32181 = ~n32169 & ~n32180;
  assign n32182 = controllable_hgrant3 & ~n32181;
  assign n32183 = ~n22755 & ~n32182;
  assign n32184 = controllable_nhgrant0 & ~n32183;
  assign n32185 = ~n9861 & ~n32184;
  assign n32186 = ~n3281 & ~n32185;
  assign n32187 = ~n3281 & ~n32186;
  assign n32188 = ~n3378 & ~n32187;
  assign n32189 = ~n32166 & ~n32188;
  assign n32190 = n3492 & ~n32189;
  assign n32191 = n3492 & ~n32190;
  assign n32192 = n3485 & ~n32191;
  assign n32193 = n3485 & ~n32192;
  assign n32194 = ~n3476 & ~n32193;
  assign n32195 = ~n5590 & ~n7401;
  assign n32196 = i_hbusreq3 & ~n32195;
  assign n32197 = ~n7399 & ~n10102;
  assign n32198 = ~controllable_hmaster1 & ~n32197;
  assign n32199 = ~n10101 & ~n32198;
  assign n32200 = ~i_hbusreq3 & ~n32199;
  assign n32201 = ~n32196 & ~n32200;
  assign n32202 = ~controllable_hmaster2 & ~n32201;
  assign n32203 = ~n10091 & ~n32202;
  assign n32204 = controllable_hgrant3 & ~n32203;
  assign n32205 = ~n22850 & ~n32204;
  assign n32206 = controllable_nhgrant0 & ~n32205;
  assign n32207 = ~n10240 & ~n32206;
  assign n32208 = ~n3281 & ~n32207;
  assign n32209 = ~n3281 & ~n32208;
  assign n32210 = n3378 & ~n32209;
  assign n32211 = ~controllable_hgrant2 & ~n23301;
  assign n32212 = ~n4562 & ~n32211;
  assign n32213 = ~i_hbusreq3 & ~n32212;
  assign n32214 = ~n6013 & ~n32213;
  assign n32215 = controllable_hmaster2 & ~n32214;
  assign n32216 = ~n7638 & ~n25707;
  assign n32217 = i_hbusreq3 & ~n32216;
  assign n32218 = ~controllable_hgrant2 & ~n23333;
  assign n32219 = ~n4562 & ~n32218;
  assign n32220 = controllable_hmaster0 & ~n32219;
  assign n32221 = ~controllable_hmaster0 & ~n32212;
  assign n32222 = ~n32220 & ~n32221;
  assign n32223 = controllable_hmaster1 & ~n32222;
  assign n32224 = controllable_hmaster0 & ~n32212;
  assign n32225 = ~n7636 & ~n32224;
  assign n32226 = ~controllable_hmaster1 & ~n32225;
  assign n32227 = ~n32223 & ~n32226;
  assign n32228 = ~i_hbusreq3 & ~n32227;
  assign n32229 = ~n32217 & ~n32228;
  assign n32230 = ~controllable_hmaster2 & ~n32229;
  assign n32231 = ~n32215 & ~n32230;
  assign n32232 = controllable_hgrant3 & ~n32231;
  assign n32233 = ~n22932 & ~n32232;
  assign n32234 = controllable_nhgrant0 & ~n32233;
  assign n32235 = ~n10240 & ~n32234;
  assign n32236 = ~n3281 & ~n32235;
  assign n32237 = ~n3281 & ~n32236;
  assign n32238 = ~n3378 & ~n32237;
  assign n32239 = ~n32210 & ~n32238;
  assign n32240 = n3492 & ~n32239;
  assign n32241 = ~n21722 & ~n32240;
  assign n32242 = n3485 & ~n32241;
  assign n32243 = ~n21721 & ~n32242;
  assign n32244 = n3476 & ~n32243;
  assign n32245 = ~n32194 & ~n32244;
  assign n32246 = n3374 & ~n32245;
  assign n32247 = ~n32150 & ~n32246;
  assign n32248 = n3655 & ~n32247;
  assign n32249 = ~n22973 & ~n32138;
  assign n32250 = controllable_nhgrant0 & ~n32249;
  assign n32251 = ~n9753 & ~n32250;
  assign n32252 = ~n3281 & ~n32251;
  assign n32253 = ~n3281 & ~n32252;
  assign n32254 = ~n3378 & ~n32253;
  assign n32255 = ~n22618 & ~n32254;
  assign n32256 = n3492 & ~n32255;
  assign n32257 = n3492 & ~n32256;
  assign n32258 = n3485 & ~n32257;
  assign n32259 = n3485 & ~n32258;
  assign n32260 = ~n3374 & ~n32259;
  assign n32261 = ~n22997 & ~n32160;
  assign n32262 = controllable_nhgrant0 & ~n32261;
  assign n32263 = ~n9861 & ~n32262;
  assign n32264 = ~n3281 & ~n32263;
  assign n32265 = ~n3281 & ~n32264;
  assign n32266 = n3378 & ~n32265;
  assign n32267 = ~n23063 & ~n32182;
  assign n32268 = controllable_nhgrant0 & ~n32267;
  assign n32269 = ~n9861 & ~n32268;
  assign n32270 = ~n3281 & ~n32269;
  assign n32271 = ~n3281 & ~n32270;
  assign n32272 = ~n3378 & ~n32271;
  assign n32273 = ~n32266 & ~n32272;
  assign n32274 = n3492 & ~n32273;
  assign n32275 = n3492 & ~n32274;
  assign n32276 = n3485 & ~n32275;
  assign n32277 = n3485 & ~n32276;
  assign n32278 = ~n3476 & ~n32277;
  assign n32279 = ~n23088 & ~n32204;
  assign n32280 = controllable_nhgrant0 & ~n32279;
  assign n32281 = ~n10240 & ~n32280;
  assign n32282 = ~n3281 & ~n32281;
  assign n32283 = ~n3281 & ~n32282;
  assign n32284 = n3378 & ~n32283;
  assign n32285 = ~n23171 & ~n32232;
  assign n32286 = controllable_nhgrant0 & ~n32285;
  assign n32287 = ~n10240 & ~n32286;
  assign n32288 = ~n3281 & ~n32287;
  assign n32289 = ~n3281 & ~n32288;
  assign n32290 = ~n3378 & ~n32289;
  assign n32291 = ~n32284 & ~n32290;
  assign n32292 = n3492 & ~n32291;
  assign n32293 = ~n21722 & ~n32292;
  assign n32294 = n3485 & ~n32293;
  assign n32295 = ~n21721 & ~n32294;
  assign n32296 = n3476 & ~n32295;
  assign n32297 = ~n32278 & ~n32296;
  assign n32298 = n3374 & ~n32297;
  assign n32299 = ~n32260 & ~n32298;
  assign n32300 = ~n3655 & ~n32299;
  assign n32301 = ~n32248 & ~n32300;
  assign n32302 = n3652 & ~n32301;
  assign n32303 = ~n23201 & ~n32138;
  assign n32304 = controllable_nhgrant0 & ~n32303;
  assign n32305 = ~n9753 & ~n32304;
  assign n32306 = ~n3281 & ~n32305;
  assign n32307 = ~n3281 & ~n32306;
  assign n32308 = ~n3378 & ~n32307;
  assign n32309 = ~n22618 & ~n32308;
  assign n32310 = n3492 & ~n32309;
  assign n32311 = n3492 & ~n32310;
  assign n32312 = n3485 & ~n32311;
  assign n32313 = n3485 & ~n32312;
  assign n32314 = ~n3374 & ~n32313;
  assign n32315 = ~n23225 & ~n32160;
  assign n32316 = controllable_nhgrant0 & ~n32315;
  assign n32317 = ~n9861 & ~n32316;
  assign n32318 = ~n3281 & ~n32317;
  assign n32319 = ~n3281 & ~n32318;
  assign n32320 = n3378 & ~n32319;
  assign n32321 = ~n23259 & ~n32182;
  assign n32322 = controllable_nhgrant0 & ~n32321;
  assign n32323 = ~n9861 & ~n32322;
  assign n32324 = ~n3281 & ~n32323;
  assign n32325 = ~n3281 & ~n32324;
  assign n32326 = ~n3378 & ~n32325;
  assign n32327 = ~n32320 & ~n32326;
  assign n32328 = n3492 & ~n32327;
  assign n32329 = n3492 & ~n32328;
  assign n32330 = n3485 & ~n32329;
  assign n32331 = n3485 & ~n32330;
  assign n32332 = ~n3476 & ~n32331;
  assign n32333 = ~n23284 & ~n32204;
  assign n32334 = controllable_nhgrant0 & ~n32333;
  assign n32335 = ~n10240 & ~n32334;
  assign n32336 = ~n3281 & ~n32335;
  assign n32337 = ~n3281 & ~n32336;
  assign n32338 = n3378 & ~n32337;
  assign n32339 = ~n23348 & ~n32232;
  assign n32340 = controllable_nhgrant0 & ~n32339;
  assign n32341 = ~n10240 & ~n32340;
  assign n32342 = ~n3281 & ~n32341;
  assign n32343 = ~n3281 & ~n32342;
  assign n32344 = ~n3378 & ~n32343;
  assign n32345 = ~n32338 & ~n32344;
  assign n32346 = n3492 & ~n32345;
  assign n32347 = ~n21722 & ~n32346;
  assign n32348 = n3485 & ~n32347;
  assign n32349 = ~n21721 & ~n32348;
  assign n32350 = n3476 & ~n32349;
  assign n32351 = ~n32332 & ~n32350;
  assign n32352 = n3374 & ~n32351;
  assign n32353 = ~n32314 & ~n32352;
  assign n32354 = n3655 & ~n32353;
  assign n32355 = ~n23375 & ~n32138;
  assign n32356 = controllable_nhgrant0 & ~n32355;
  assign n32357 = ~n9753 & ~n32356;
  assign n32358 = ~n3281 & ~n32357;
  assign n32359 = ~n3281 & ~n32358;
  assign n32360 = ~n3378 & ~n32359;
  assign n32361 = ~n22618 & ~n32360;
  assign n32362 = n3492 & ~n32361;
  assign n32363 = n3492 & ~n32362;
  assign n32364 = n3485 & ~n32363;
  assign n32365 = n3485 & ~n32364;
  assign n32366 = ~n3374 & ~n32365;
  assign n32367 = ~n23399 & ~n32160;
  assign n32368 = controllable_nhgrant0 & ~n32367;
  assign n32369 = ~n9861 & ~n32368;
  assign n32370 = ~n3281 & ~n32369;
  assign n32371 = ~n3281 & ~n32370;
  assign n32372 = n3378 & ~n32371;
  assign n32373 = ~n23433 & ~n32182;
  assign n32374 = controllable_nhgrant0 & ~n32373;
  assign n32375 = ~n9861 & ~n32374;
  assign n32376 = ~n3281 & ~n32375;
  assign n32377 = ~n3281 & ~n32376;
  assign n32378 = ~n3378 & ~n32377;
  assign n32379 = ~n32372 & ~n32378;
  assign n32380 = n3492 & ~n32379;
  assign n32381 = n3492 & ~n32380;
  assign n32382 = n3485 & ~n32381;
  assign n32383 = n3485 & ~n32382;
  assign n32384 = ~n3476 & ~n32383;
  assign n32385 = ~n23458 & ~n32204;
  assign n32386 = controllable_nhgrant0 & ~n32385;
  assign n32387 = ~n10240 & ~n32386;
  assign n32388 = ~n3281 & ~n32387;
  assign n32389 = ~n3281 & ~n32388;
  assign n32390 = n3378 & ~n32389;
  assign n32391 = ~n23496 & ~n32232;
  assign n32392 = controllable_nhgrant0 & ~n32391;
  assign n32393 = ~n10240 & ~n32392;
  assign n32394 = ~n3281 & ~n32393;
  assign n32395 = ~n3281 & ~n32394;
  assign n32396 = ~n3378 & ~n32395;
  assign n32397 = ~n32390 & ~n32396;
  assign n32398 = n3492 & ~n32397;
  assign n32399 = ~n21722 & ~n32398;
  assign n32400 = n3485 & ~n32399;
  assign n32401 = ~n21721 & ~n32400;
  assign n32402 = n3476 & ~n32401;
  assign n32403 = ~n32384 & ~n32402;
  assign n32404 = n3374 & ~n32403;
  assign n32405 = ~n32366 & ~n32404;
  assign n32406 = ~n3655 & ~n32405;
  assign n32407 = ~n32354 & ~n32406;
  assign n32408 = ~n3652 & ~n32407;
  assign n32409 = ~n32302 & ~n32408;
  assign n32410 = n3368 & ~n32409;
  assign n32411 = ~n32129 & ~n32410;
  assign n32412 = n3362 & ~n32411;
  assign n32413 = n3492 & ~n31853;
  assign n32414 = ~n3631 & ~n32413;
  assign n32415 = n3485 & ~n32414;
  assign n32416 = ~n3630 & ~n32415;
  assign n32417 = ~n3476 & ~n32416;
  assign n32418 = ~n23549 & ~n26200;
  assign n32419 = ~n3485 & ~n32418;
  assign n32420 = ~n8309 & ~n32413;
  assign n32421 = n3485 & ~n32420;
  assign n32422 = ~n32419 & ~n32421;
  assign n32423 = n3476 & ~n32422;
  assign n32424 = ~n32417 & ~n32423;
  assign n32425 = ~n3374 & ~n32424;
  assign n32426 = n3492 & ~n31895;
  assign n32427 = ~n3631 & ~n32426;
  assign n32428 = n3485 & ~n32427;
  assign n32429 = ~n3630 & ~n32428;
  assign n32430 = ~n3476 & ~n32429;
  assign n32431 = n3492 & ~n31938;
  assign n32432 = ~n8309 & ~n32431;
  assign n32433 = n3485 & ~n32432;
  assign n32434 = ~n32419 & ~n32433;
  assign n32435 = n3476 & ~n32434;
  assign n32436 = ~n32430 & ~n32435;
  assign n32437 = n3374 & ~n32436;
  assign n32438 = ~n32425 & ~n32437;
  assign n32439 = n3655 & ~n32438;
  assign n32440 = n3492 & ~n31954;
  assign n32441 = ~n3631 & ~n32440;
  assign n32442 = n3485 & ~n32441;
  assign n32443 = ~n3630 & ~n32442;
  assign n32444 = ~n3476 & ~n32443;
  assign n32445 = ~n23549 & ~n26297;
  assign n32446 = ~n3485 & ~n32445;
  assign n32447 = ~n8309 & ~n32440;
  assign n32448 = n3485 & ~n32447;
  assign n32449 = ~n32446 & ~n32448;
  assign n32450 = n3476 & ~n32449;
  assign n32451 = ~n32444 & ~n32450;
  assign n32452 = ~n3374 & ~n32451;
  assign n32453 = n3492 & ~n31978;
  assign n32454 = ~n3631 & ~n32453;
  assign n32455 = n3485 & ~n32454;
  assign n32456 = ~n3630 & ~n32455;
  assign n32457 = ~n3476 & ~n32456;
  assign n32458 = n3492 & ~n31996;
  assign n32459 = ~n8309 & ~n32458;
  assign n32460 = n3485 & ~n32459;
  assign n32461 = ~n32446 & ~n32460;
  assign n32462 = n3476 & ~n32461;
  assign n32463 = ~n32457 & ~n32462;
  assign n32464 = n3374 & ~n32463;
  assign n32465 = ~n32452 & ~n32464;
  assign n32466 = ~n3655 & ~n32465;
  assign n32467 = ~n32439 & ~n32466;
  assign n32468 = n3652 & ~n32467;
  assign n32469 = n3492 & ~n32014;
  assign n32470 = ~n3631 & ~n32469;
  assign n32471 = n3485 & ~n32470;
  assign n32472 = ~n3630 & ~n32471;
  assign n32473 = ~n3476 & ~n32472;
  assign n32474 = ~n23549 & ~n26396;
  assign n32475 = ~n3485 & ~n32474;
  assign n32476 = ~n8309 & ~n32469;
  assign n32477 = n3485 & ~n32476;
  assign n32478 = ~n32475 & ~n32477;
  assign n32479 = n3476 & ~n32478;
  assign n32480 = ~n32473 & ~n32479;
  assign n32481 = ~n3374 & ~n32480;
  assign n32482 = n3492 & ~n32038;
  assign n32483 = ~n3631 & ~n32482;
  assign n32484 = n3485 & ~n32483;
  assign n32485 = ~n3630 & ~n32484;
  assign n32486 = ~n3476 & ~n32485;
  assign n32487 = n3492 & ~n32056;
  assign n32488 = ~n8309 & ~n32487;
  assign n32489 = n3485 & ~n32488;
  assign n32490 = ~n32475 & ~n32489;
  assign n32491 = n3476 & ~n32490;
  assign n32492 = ~n32486 & ~n32491;
  assign n32493 = n3374 & ~n32492;
  assign n32494 = ~n32481 & ~n32493;
  assign n32495 = n3655 & ~n32494;
  assign n32496 = n3492 & ~n32072;
  assign n32497 = ~n3631 & ~n32496;
  assign n32498 = n3485 & ~n32497;
  assign n32499 = ~n3630 & ~n32498;
  assign n32500 = ~n3476 & ~n32499;
  assign n32501 = ~n23549 & ~n26437;
  assign n32502 = ~n3485 & ~n32501;
  assign n32503 = ~n8309 & ~n32496;
  assign n32504 = n3485 & ~n32503;
  assign n32505 = ~n32502 & ~n32504;
  assign n32506 = n3476 & ~n32505;
  assign n32507 = ~n32500 & ~n32506;
  assign n32508 = ~n3374 & ~n32507;
  assign n32509 = n3492 & ~n32096;
  assign n32510 = ~n3631 & ~n32509;
  assign n32511 = n3485 & ~n32510;
  assign n32512 = ~n3630 & ~n32511;
  assign n32513 = ~n3476 & ~n32512;
  assign n32514 = n3492 & ~n32114;
  assign n32515 = ~n8309 & ~n32514;
  assign n32516 = n3485 & ~n32515;
  assign n32517 = ~n32502 & ~n32516;
  assign n32518 = n3476 & ~n32517;
  assign n32519 = ~n32513 & ~n32518;
  assign n32520 = n3374 & ~n32519;
  assign n32521 = ~n32508 & ~n32520;
  assign n32522 = ~n3655 & ~n32521;
  assign n32523 = ~n32495 & ~n32522;
  assign n32524 = ~n3652 & ~n32523;
  assign n32525 = ~n32468 & ~n32524;
  assign n32526 = ~n3368 & ~n32525;
  assign n32527 = n3492 & ~n32143;
  assign n32528 = n3492 & ~n32527;
  assign n32529 = n3485 & ~n32528;
  assign n32530 = n3485 & ~n32529;
  assign n32531 = ~n3476 & ~n32530;
  assign n32532 = ~n8525 & ~n32529;
  assign n32533 = n3476 & ~n32532;
  assign n32534 = ~n32531 & ~n32533;
  assign n32535 = ~n3374 & ~n32534;
  assign n32536 = n3492 & ~n32187;
  assign n32537 = n3492 & ~n32536;
  assign n32538 = n3485 & ~n32537;
  assign n32539 = n3485 & ~n32538;
  assign n32540 = ~n3476 & ~n32539;
  assign n32541 = ~n23646 & ~n26477;
  assign n32542 = ~n3485 & ~n32541;
  assign n32543 = n3492 & ~n32237;
  assign n32544 = ~n21722 & ~n32543;
  assign n32545 = n3485 & ~n32544;
  assign n32546 = ~n32542 & ~n32545;
  assign n32547 = n3476 & ~n32546;
  assign n32548 = ~n32540 & ~n32547;
  assign n32549 = n3374 & ~n32548;
  assign n32550 = ~n32535 & ~n32549;
  assign n32551 = n3655 & ~n32550;
  assign n32552 = n3492 & ~n32253;
  assign n32553 = n3492 & ~n32552;
  assign n32554 = n3485 & ~n32553;
  assign n32555 = n3485 & ~n32554;
  assign n32556 = ~n3476 & ~n32555;
  assign n32557 = ~n8525 & ~n32554;
  assign n32558 = n3476 & ~n32557;
  assign n32559 = ~n32556 & ~n32558;
  assign n32560 = ~n3374 & ~n32559;
  assign n32561 = n3492 & ~n32271;
  assign n32562 = n3492 & ~n32561;
  assign n32563 = n3485 & ~n32562;
  assign n32564 = n3485 & ~n32563;
  assign n32565 = ~n3476 & ~n32564;
  assign n32566 = ~n23646 & ~n26504;
  assign n32567 = ~n3485 & ~n32566;
  assign n32568 = n3492 & ~n32289;
  assign n32569 = ~n21722 & ~n32568;
  assign n32570 = n3485 & ~n32569;
  assign n32571 = ~n32567 & ~n32570;
  assign n32572 = n3476 & ~n32571;
  assign n32573 = ~n32565 & ~n32572;
  assign n32574 = n3374 & ~n32573;
  assign n32575 = ~n32560 & ~n32574;
  assign n32576 = ~n3655 & ~n32575;
  assign n32577 = ~n32551 & ~n32576;
  assign n32578 = n3652 & ~n32577;
  assign n32579 = n3492 & ~n32307;
  assign n32580 = n3492 & ~n32579;
  assign n32581 = n3485 & ~n32580;
  assign n32582 = n3485 & ~n32581;
  assign n32583 = ~n3476 & ~n32582;
  assign n32584 = ~n8525 & ~n32581;
  assign n32585 = n3476 & ~n32584;
  assign n32586 = ~n32583 & ~n32585;
  assign n32587 = ~n3374 & ~n32586;
  assign n32588 = n3492 & ~n32325;
  assign n32589 = n3492 & ~n32588;
  assign n32590 = n3485 & ~n32589;
  assign n32591 = n3485 & ~n32590;
  assign n32592 = ~n3476 & ~n32591;
  assign n32593 = ~n23646 & ~n26533;
  assign n32594 = ~n3485 & ~n32593;
  assign n32595 = n3492 & ~n32343;
  assign n32596 = ~n21722 & ~n32595;
  assign n32597 = n3485 & ~n32596;
  assign n32598 = ~n32594 & ~n32597;
  assign n32599 = n3476 & ~n32598;
  assign n32600 = ~n32592 & ~n32599;
  assign n32601 = n3374 & ~n32600;
  assign n32602 = ~n32587 & ~n32601;
  assign n32603 = n3655 & ~n32602;
  assign n32604 = n3492 & ~n32359;
  assign n32605 = n3492 & ~n32604;
  assign n32606 = n3485 & ~n32605;
  assign n32607 = n3485 & ~n32606;
  assign n32608 = ~n3476 & ~n32607;
  assign n32609 = ~n8525 & ~n32606;
  assign n32610 = n3476 & ~n32609;
  assign n32611 = ~n32608 & ~n32610;
  assign n32612 = ~n3374 & ~n32611;
  assign n32613 = n3492 & ~n32377;
  assign n32614 = n3492 & ~n32613;
  assign n32615 = n3485 & ~n32614;
  assign n32616 = n3485 & ~n32615;
  assign n32617 = ~n3476 & ~n32616;
  assign n32618 = ~n23646 & ~n26560;
  assign n32619 = ~n3485 & ~n32618;
  assign n32620 = n3492 & ~n32395;
  assign n32621 = ~n21722 & ~n32620;
  assign n32622 = n3485 & ~n32621;
  assign n32623 = ~n32619 & ~n32622;
  assign n32624 = n3476 & ~n32623;
  assign n32625 = ~n32617 & ~n32624;
  assign n32626 = n3374 & ~n32625;
  assign n32627 = ~n32612 & ~n32626;
  assign n32628 = ~n3655 & ~n32627;
  assign n32629 = ~n32603 & ~n32628;
  assign n32630 = ~n3652 & ~n32629;
  assign n32631 = ~n32578 & ~n32630;
  assign n32632 = n3368 & ~n32631;
  assign n32633 = ~n32526 & ~n32632;
  assign n32634 = ~n3362 & ~n32633;
  assign n32635 = ~n32412 & ~n32634;
  assign n32636 = n3359 & ~n32635;
  assign n32637 = ~n26580 & ~n32421;
  assign n32638 = n3476 & ~n32637;
  assign n32639 = ~n32417 & ~n32638;
  assign n32640 = ~n3374 & ~n32639;
  assign n32641 = ~n26580 & ~n32433;
  assign n32642 = n3476 & ~n32641;
  assign n32643 = ~n32430 & ~n32642;
  assign n32644 = n3374 & ~n32643;
  assign n32645 = ~n32640 & ~n32644;
  assign n32646 = n3655 & ~n32645;
  assign n32647 = ~n26591 & ~n32448;
  assign n32648 = n3476 & ~n32647;
  assign n32649 = ~n32444 & ~n32648;
  assign n32650 = ~n3374 & ~n32649;
  assign n32651 = ~n26591 & ~n32460;
  assign n32652 = n3476 & ~n32651;
  assign n32653 = ~n32457 & ~n32652;
  assign n32654 = n3374 & ~n32653;
  assign n32655 = ~n32650 & ~n32654;
  assign n32656 = ~n3655 & ~n32655;
  assign n32657 = ~n32646 & ~n32656;
  assign n32658 = n3652 & ~n32657;
  assign n32659 = ~n26604 & ~n32477;
  assign n32660 = n3476 & ~n32659;
  assign n32661 = ~n32473 & ~n32660;
  assign n32662 = ~n3374 & ~n32661;
  assign n32663 = ~n26604 & ~n32489;
  assign n32664 = n3476 & ~n32663;
  assign n32665 = ~n32486 & ~n32664;
  assign n32666 = n3374 & ~n32665;
  assign n32667 = ~n32662 & ~n32666;
  assign n32668 = n3655 & ~n32667;
  assign n32669 = ~n26615 & ~n32504;
  assign n32670 = n3476 & ~n32669;
  assign n32671 = ~n32500 & ~n32670;
  assign n32672 = ~n3374 & ~n32671;
  assign n32673 = ~n26615 & ~n32516;
  assign n32674 = n3476 & ~n32673;
  assign n32675 = ~n32513 & ~n32674;
  assign n32676 = n3374 & ~n32675;
  assign n32677 = ~n32672 & ~n32676;
  assign n32678 = ~n3655 & ~n32677;
  assign n32679 = ~n32668 & ~n32678;
  assign n32680 = ~n3652 & ~n32679;
  assign n32681 = ~n32658 & ~n32680;
  assign n32682 = ~n3368 & ~n32681;
  assign n32683 = ~n8689 & ~n32529;
  assign n32684 = n3476 & ~n32683;
  assign n32685 = ~n32531 & ~n32684;
  assign n32686 = ~n3374 & ~n32685;
  assign n32687 = ~n26634 & ~n32545;
  assign n32688 = n3476 & ~n32687;
  assign n32689 = ~n32540 & ~n32688;
  assign n32690 = n3374 & ~n32689;
  assign n32691 = ~n32686 & ~n32690;
  assign n32692 = n3655 & ~n32691;
  assign n32693 = ~n8689 & ~n32554;
  assign n32694 = n3476 & ~n32693;
  assign n32695 = ~n32556 & ~n32694;
  assign n32696 = ~n3374 & ~n32695;
  assign n32697 = ~n26645 & ~n32570;
  assign n32698 = n3476 & ~n32697;
  assign n32699 = ~n32565 & ~n32698;
  assign n32700 = n3374 & ~n32699;
  assign n32701 = ~n32696 & ~n32700;
  assign n32702 = ~n3655 & ~n32701;
  assign n32703 = ~n32692 & ~n32702;
  assign n32704 = n3652 & ~n32703;
  assign n32705 = ~n8689 & ~n32581;
  assign n32706 = n3476 & ~n32705;
  assign n32707 = ~n32583 & ~n32706;
  assign n32708 = ~n3374 & ~n32707;
  assign n32709 = ~n26658 & ~n32597;
  assign n32710 = n3476 & ~n32709;
  assign n32711 = ~n32592 & ~n32710;
  assign n32712 = n3374 & ~n32711;
  assign n32713 = ~n32708 & ~n32712;
  assign n32714 = n3655 & ~n32713;
  assign n32715 = ~n8689 & ~n32606;
  assign n32716 = n3476 & ~n32715;
  assign n32717 = ~n32608 & ~n32716;
  assign n32718 = ~n3374 & ~n32717;
  assign n32719 = ~n26669 & ~n32622;
  assign n32720 = n3476 & ~n32719;
  assign n32721 = ~n32617 & ~n32720;
  assign n32722 = n3374 & ~n32721;
  assign n32723 = ~n32718 & ~n32722;
  assign n32724 = ~n3655 & ~n32723;
  assign n32725 = ~n32714 & ~n32724;
  assign n32726 = ~n3652 & ~n32725;
  assign n32727 = ~n32704 & ~n32726;
  assign n32728 = n3368 & ~n32727;
  assign n32729 = ~n32682 & ~n32728;
  assign n32730 = n3362 & ~n32729;
  assign n32731 = n3378 & ~n31853;
  assign n32732 = ~n26690 & ~n32731;
  assign n32733 = n3492 & ~n32732;
  assign n32734 = ~n3631 & ~n32733;
  assign n32735 = n3485 & ~n32734;
  assign n32736 = ~n3630 & ~n32735;
  assign n32737 = ~n3476 & ~n32736;
  assign n32738 = ~n26200 & ~n32733;
  assign n32739 = n3485 & ~n32738;
  assign n32740 = ~n26580 & ~n32739;
  assign n32741 = n3476 & ~n32740;
  assign n32742 = ~n32737 & ~n32741;
  assign n32743 = ~n3374 & ~n32742;
  assign n32744 = n3378 & ~n31895;
  assign n32745 = ~n26711 & ~n32744;
  assign n32746 = n3492 & ~n32745;
  assign n32747 = ~n3631 & ~n32746;
  assign n32748 = n3485 & ~n32747;
  assign n32749 = ~n3630 & ~n32748;
  assign n32750 = ~n3476 & ~n32749;
  assign n32751 = n3378 & ~n31938;
  assign n32752 = ~n26726 & ~n32751;
  assign n32753 = n3492 & ~n32752;
  assign n32754 = ~n26200 & ~n32753;
  assign n32755 = n3485 & ~n32754;
  assign n32756 = ~n26580 & ~n32755;
  assign n32757 = n3476 & ~n32756;
  assign n32758 = ~n32750 & ~n32757;
  assign n32759 = n3374 & ~n32758;
  assign n32760 = ~n32743 & ~n32759;
  assign n32761 = n3655 & ~n32760;
  assign n32762 = n3378 & ~n31954;
  assign n32763 = ~n26743 & ~n32762;
  assign n32764 = n3492 & ~n32763;
  assign n32765 = ~n3631 & ~n32764;
  assign n32766 = n3485 & ~n32765;
  assign n32767 = ~n3630 & ~n32766;
  assign n32768 = ~n3476 & ~n32767;
  assign n32769 = ~n26297 & ~n32764;
  assign n32770 = n3485 & ~n32769;
  assign n32771 = ~n26591 & ~n32770;
  assign n32772 = n3476 & ~n32771;
  assign n32773 = ~n32768 & ~n32772;
  assign n32774 = ~n3374 & ~n32773;
  assign n32775 = n3378 & ~n31978;
  assign n32776 = ~n26762 & ~n32775;
  assign n32777 = n3492 & ~n32776;
  assign n32778 = ~n3631 & ~n32777;
  assign n32779 = n3485 & ~n32778;
  assign n32780 = ~n3630 & ~n32779;
  assign n32781 = ~n3476 & ~n32780;
  assign n32782 = n3378 & ~n31996;
  assign n32783 = ~n26775 & ~n32782;
  assign n32784 = n3492 & ~n32783;
  assign n32785 = ~n26297 & ~n32784;
  assign n32786 = n3485 & ~n32785;
  assign n32787 = ~n26591 & ~n32786;
  assign n32788 = n3476 & ~n32787;
  assign n32789 = ~n32781 & ~n32788;
  assign n32790 = n3374 & ~n32789;
  assign n32791 = ~n32774 & ~n32790;
  assign n32792 = ~n3655 & ~n32791;
  assign n32793 = ~n32761 & ~n32792;
  assign n32794 = n3652 & ~n32793;
  assign n32795 = n3378 & ~n32014;
  assign n32796 = ~n26794 & ~n32795;
  assign n32797 = n3492 & ~n32796;
  assign n32798 = ~n3631 & ~n32797;
  assign n32799 = n3485 & ~n32798;
  assign n32800 = ~n3630 & ~n32799;
  assign n32801 = ~n3476 & ~n32800;
  assign n32802 = ~n26396 & ~n32797;
  assign n32803 = n3485 & ~n32802;
  assign n32804 = ~n26604 & ~n32803;
  assign n32805 = n3476 & ~n32804;
  assign n32806 = ~n32801 & ~n32805;
  assign n32807 = ~n3374 & ~n32806;
  assign n32808 = n3378 & ~n32038;
  assign n32809 = ~n26813 & ~n32808;
  assign n32810 = n3492 & ~n32809;
  assign n32811 = ~n3631 & ~n32810;
  assign n32812 = n3485 & ~n32811;
  assign n32813 = ~n3630 & ~n32812;
  assign n32814 = ~n3476 & ~n32813;
  assign n32815 = n3378 & ~n32056;
  assign n32816 = ~n26826 & ~n32815;
  assign n32817 = n3492 & ~n32816;
  assign n32818 = ~n26396 & ~n32817;
  assign n32819 = n3485 & ~n32818;
  assign n32820 = ~n26604 & ~n32819;
  assign n32821 = n3476 & ~n32820;
  assign n32822 = ~n32814 & ~n32821;
  assign n32823 = n3374 & ~n32822;
  assign n32824 = ~n32807 & ~n32823;
  assign n32825 = n3655 & ~n32824;
  assign n32826 = n3378 & ~n32072;
  assign n32827 = ~n26843 & ~n32826;
  assign n32828 = n3492 & ~n32827;
  assign n32829 = ~n3631 & ~n32828;
  assign n32830 = n3485 & ~n32829;
  assign n32831 = ~n3630 & ~n32830;
  assign n32832 = ~n3476 & ~n32831;
  assign n32833 = ~n26437 & ~n32828;
  assign n32834 = n3485 & ~n32833;
  assign n32835 = ~n26615 & ~n32834;
  assign n32836 = n3476 & ~n32835;
  assign n32837 = ~n32832 & ~n32836;
  assign n32838 = ~n3374 & ~n32837;
  assign n32839 = n3378 & ~n32096;
  assign n32840 = ~n26862 & ~n32839;
  assign n32841 = n3492 & ~n32840;
  assign n32842 = ~n3631 & ~n32841;
  assign n32843 = n3485 & ~n32842;
  assign n32844 = ~n3630 & ~n32843;
  assign n32845 = ~n3476 & ~n32844;
  assign n32846 = n3378 & ~n32114;
  assign n32847 = ~n26875 & ~n32846;
  assign n32848 = n3492 & ~n32847;
  assign n32849 = ~n26437 & ~n32848;
  assign n32850 = n3485 & ~n32849;
  assign n32851 = ~n26615 & ~n32850;
  assign n32852 = n3476 & ~n32851;
  assign n32853 = ~n32845 & ~n32852;
  assign n32854 = n3374 & ~n32853;
  assign n32855 = ~n32838 & ~n32854;
  assign n32856 = ~n3655 & ~n32855;
  assign n32857 = ~n32825 & ~n32856;
  assign n32858 = ~n3652 & ~n32857;
  assign n32859 = ~n32794 & ~n32858;
  assign n32860 = ~n3368 & ~n32859;
  assign n32861 = n3378 & ~n32143;
  assign n32862 = ~n26897 & ~n32861;
  assign n32863 = n3492 & ~n32862;
  assign n32864 = n3492 & ~n32863;
  assign n32865 = n3485 & ~n32864;
  assign n32866 = n3485 & ~n32865;
  assign n32867 = ~n3476 & ~n32866;
  assign n32868 = ~n8523 & ~n32863;
  assign n32869 = n3485 & ~n32868;
  assign n32870 = ~n8689 & ~n32869;
  assign n32871 = n3476 & ~n32870;
  assign n32872 = ~n32867 & ~n32871;
  assign n32873 = ~n3374 & ~n32872;
  assign n32874 = n3378 & ~n32187;
  assign n32875 = ~n26931 & ~n32874;
  assign n32876 = n3492 & ~n32875;
  assign n32877 = n3492 & ~n32876;
  assign n32878 = n3485 & ~n32877;
  assign n32879 = n3485 & ~n32878;
  assign n32880 = ~n3476 & ~n32879;
  assign n32881 = ~i_hbusreq2 & ~n24199;
  assign n32882 = ~n26962 & ~n32881;
  assign n32883 = ~controllable_hgrant2 & ~n32882;
  assign n32884 = ~n4562 & ~n32883;
  assign n32885 = i_hlock3 & ~n32884;
  assign n32886 = ~i_hbusreq2 & ~n24209;
  assign n32887 = ~n26979 & ~n32886;
  assign n32888 = ~controllable_hgrant2 & ~n32887;
  assign n32889 = ~n4562 & ~n32888;
  assign n32890 = ~i_hlock3 & ~n32889;
  assign n32891 = ~n32885 & ~n32890;
  assign n32892 = ~i_hbusreq3 & ~n32891;
  assign n32893 = ~n30147 & ~n32892;
  assign n32894 = controllable_hmaster2 & ~n32893;
  assign n32895 = ~n26946 & ~n27005;
  assign n32896 = i_hlock3 & ~n32895;
  assign n32897 = ~n26957 & ~n27014;
  assign n32898 = ~i_hlock3 & ~n32897;
  assign n32899 = ~n32896 & ~n32898;
  assign n32900 = i_hbusreq3 & ~n32899;
  assign n32901 = ~i_hbusreq2 & ~n24240;
  assign n32902 = ~n27020 & ~n32901;
  assign n32903 = ~controllable_hgrant2 & ~n32902;
  assign n32904 = ~n4562 & ~n32903;
  assign n32905 = controllable_hmaster0 & ~n32904;
  assign n32906 = ~controllable_hmaster0 & ~n32884;
  assign n32907 = ~n32905 & ~n32906;
  assign n32908 = controllable_hmaster1 & ~n32907;
  assign n32909 = controllable_hmaster0 & ~n32884;
  assign n32910 = ~n27114 & ~n32909;
  assign n32911 = ~controllable_hmaster1 & ~n32910;
  assign n32912 = ~n32908 & ~n32911;
  assign n32913 = i_hlock3 & ~n32912;
  assign n32914 = ~i_hbusreq2 & ~n24250;
  assign n32915 = ~n27038 & ~n32914;
  assign n32916 = ~controllable_hgrant2 & ~n32915;
  assign n32917 = ~n4562 & ~n32916;
  assign n32918 = controllable_hmaster0 & ~n32917;
  assign n32919 = ~controllable_hmaster0 & ~n32889;
  assign n32920 = ~n32918 & ~n32919;
  assign n32921 = controllable_hmaster1 & ~n32920;
  assign n32922 = controllable_hmaster0 & ~n32889;
  assign n32923 = ~n26955 & ~n32922;
  assign n32924 = ~controllable_hmaster1 & ~n32923;
  assign n32925 = ~n32921 & ~n32924;
  assign n32926 = ~i_hlock3 & ~n32925;
  assign n32927 = ~n32913 & ~n32926;
  assign n32928 = ~i_hbusreq3 & ~n32927;
  assign n32929 = ~n32900 & ~n32928;
  assign n32930 = ~controllable_hmaster2 & ~n32929;
  assign n32931 = ~n32894 & ~n32930;
  assign n32932 = controllable_hgrant3 & ~n32931;
  assign n32933 = ~n24043 & ~n32932;
  assign n32934 = controllable_nhgrant0 & ~n32933;
  assign n32935 = ~n10240 & ~n32934;
  assign n32936 = ~n3281 & ~n32935;
  assign n32937 = ~n3281 & ~n32936;
  assign n32938 = n3378 & ~n32937;
  assign n32939 = ~n27144 & ~n32938;
  assign n32940 = n3492 & ~n32939;
  assign n32941 = ~n26477 & ~n32940;
  assign n32942 = n3485 & ~n32941;
  assign n32943 = ~n26634 & ~n32942;
  assign n32944 = n3476 & ~n32943;
  assign n32945 = ~n32880 & ~n32944;
  assign n32946 = n3374 & ~n32945;
  assign n32947 = ~n32873 & ~n32946;
  assign n32948 = n3655 & ~n32947;
  assign n32949 = n3378 & ~n32253;
  assign n32950 = ~n27161 & ~n32949;
  assign n32951 = n3492 & ~n32950;
  assign n32952 = n3492 & ~n32951;
  assign n32953 = n3485 & ~n32952;
  assign n32954 = n3485 & ~n32953;
  assign n32955 = ~n3476 & ~n32954;
  assign n32956 = ~n8523 & ~n32951;
  assign n32957 = n3485 & ~n32956;
  assign n32958 = ~n8689 & ~n32957;
  assign n32959 = n3476 & ~n32958;
  assign n32960 = ~n32955 & ~n32959;
  assign n32961 = ~n3374 & ~n32960;
  assign n32962 = n3378 & ~n32271;
  assign n32963 = ~n27180 & ~n32962;
  assign n32964 = n3492 & ~n32963;
  assign n32965 = n3492 & ~n32964;
  assign n32966 = n3485 & ~n32965;
  assign n32967 = n3485 & ~n32966;
  assign n32968 = ~n3476 & ~n32967;
  assign n32969 = ~n24152 & ~n32932;
  assign n32970 = controllable_nhgrant0 & ~n32969;
  assign n32971 = ~n10240 & ~n32970;
  assign n32972 = ~n3281 & ~n32971;
  assign n32973 = ~n3281 & ~n32972;
  assign n32974 = n3378 & ~n32973;
  assign n32975 = ~n27198 & ~n32974;
  assign n32976 = n3492 & ~n32975;
  assign n32977 = ~n26504 & ~n32976;
  assign n32978 = n3485 & ~n32977;
  assign n32979 = ~n26645 & ~n32978;
  assign n32980 = n3476 & ~n32979;
  assign n32981 = ~n32968 & ~n32980;
  assign n32982 = n3374 & ~n32981;
  assign n32983 = ~n32961 & ~n32982;
  assign n32984 = ~n3655 & ~n32983;
  assign n32985 = ~n32948 & ~n32984;
  assign n32986 = n3652 & ~n32985;
  assign n32987 = n3378 & ~n32307;
  assign n32988 = ~n27217 & ~n32987;
  assign n32989 = n3492 & ~n32988;
  assign n32990 = n3492 & ~n32989;
  assign n32991 = n3485 & ~n32990;
  assign n32992 = n3485 & ~n32991;
  assign n32993 = ~n3476 & ~n32992;
  assign n32994 = ~n8523 & ~n32989;
  assign n32995 = n3485 & ~n32994;
  assign n32996 = ~n8689 & ~n32995;
  assign n32997 = n3476 & ~n32996;
  assign n32998 = ~n32993 & ~n32997;
  assign n32999 = ~n3374 & ~n32998;
  assign n33000 = n3378 & ~n32325;
  assign n33001 = ~n27236 & ~n33000;
  assign n33002 = n3492 & ~n33001;
  assign n33003 = n3492 & ~n33002;
  assign n33004 = n3485 & ~n33003;
  assign n33005 = n3485 & ~n33004;
  assign n33006 = ~n3476 & ~n33005;
  assign n33007 = ~n24269 & ~n32932;
  assign n33008 = controllable_nhgrant0 & ~n33007;
  assign n33009 = ~n10240 & ~n33008;
  assign n33010 = ~n3281 & ~n33009;
  assign n33011 = ~n3281 & ~n33010;
  assign n33012 = n3378 & ~n33011;
  assign n33013 = ~n27254 & ~n33012;
  assign n33014 = n3492 & ~n33013;
  assign n33015 = ~n26533 & ~n33014;
  assign n33016 = n3485 & ~n33015;
  assign n33017 = ~n26658 & ~n33016;
  assign n33018 = n3476 & ~n33017;
  assign n33019 = ~n33006 & ~n33018;
  assign n33020 = n3374 & ~n33019;
  assign n33021 = ~n32999 & ~n33020;
  assign n33022 = n3655 & ~n33021;
  assign n33023 = n3378 & ~n32359;
  assign n33024 = ~n27271 & ~n33023;
  assign n33025 = n3492 & ~n33024;
  assign n33026 = n3492 & ~n33025;
  assign n33027 = n3485 & ~n33026;
  assign n33028 = n3485 & ~n33027;
  assign n33029 = ~n3476 & ~n33028;
  assign n33030 = ~n8523 & ~n33025;
  assign n33031 = n3485 & ~n33030;
  assign n33032 = ~n8689 & ~n33031;
  assign n33033 = n3476 & ~n33032;
  assign n33034 = ~n33029 & ~n33033;
  assign n33035 = ~n3374 & ~n33034;
  assign n33036 = n3378 & ~n32377;
  assign n33037 = ~n27290 & ~n33036;
  assign n33038 = n3492 & ~n33037;
  assign n33039 = n3492 & ~n33038;
  assign n33040 = n3485 & ~n33039;
  assign n33041 = n3485 & ~n33040;
  assign n33042 = ~n3476 & ~n33041;
  assign n33043 = ~n24336 & ~n32932;
  assign n33044 = controllable_nhgrant0 & ~n33043;
  assign n33045 = ~n10240 & ~n33044;
  assign n33046 = ~n3281 & ~n33045;
  assign n33047 = ~n3281 & ~n33046;
  assign n33048 = n3378 & ~n33047;
  assign n33049 = ~n27308 & ~n33048;
  assign n33050 = n3492 & ~n33049;
  assign n33051 = ~n26560 & ~n33050;
  assign n33052 = n3485 & ~n33051;
  assign n33053 = ~n26669 & ~n33052;
  assign n33054 = n3476 & ~n33053;
  assign n33055 = ~n33042 & ~n33054;
  assign n33056 = n3374 & ~n33055;
  assign n33057 = ~n33035 & ~n33056;
  assign n33058 = ~n3655 & ~n33057;
  assign n33059 = ~n33022 & ~n33058;
  assign n33060 = ~n3652 & ~n33059;
  assign n33061 = ~n32986 & ~n33060;
  assign n33062 = n3368 & ~n33061;
  assign n33063 = ~n32860 & ~n33062;
  assign n33064 = ~n3362 & ~n33063;
  assign n33065 = ~n32730 & ~n33064;
  assign n33066 = ~n3359 & ~n33065;
  assign n33067 = ~n32636 & ~n33066;
  assign n33068 = ~n3356 & ~n33067;
  assign n33069 = ~n31840 & ~n33068;
  assign n33070 = n3345 & ~n33069;
  assign n33071 = ~n31569 & ~n33070;
  assign n33072 = ~n3341 & ~n33071;
  assign n33073 = controllable_hgrant3 & ~n24373;
  assign n33074 = ~n24370 & ~n33073;
  assign n33075 = controllable_nhgrant0 & ~n33074;
  assign n33076 = ~n24376 & ~n33075;
  assign n33077 = ~n3281 & ~n33076;
  assign n33078 = ~n3783 & ~n33077;
  assign n33079 = ~n3378 & ~n33078;
  assign n33080 = ~n3378 & ~n33079;
  assign n33081 = n3492 & ~n33080;
  assign n33082 = ~n3493 & ~n33081;
  assign n33083 = n3485 & ~n33082;
  assign n33084 = ~n3486 & ~n33083;
  assign n33085 = ~n3476 & ~n33084;
  assign n33086 = ~n3281 & ~n26688;
  assign n33087 = n3378 & ~n33086;
  assign n33088 = ~n26690 & ~n33087;
  assign n33089 = n3492 & ~n33088;
  assign n33090 = ~n3493 & ~n33089;
  assign n33091 = n3485 & ~n33090;
  assign n33092 = ~n3486 & ~n33091;
  assign n33093 = n3476 & ~n33092;
  assign n33094 = ~n33085 & ~n33093;
  assign n33095 = ~n3374 & ~n33094;
  assign n33096 = ~n3950 & ~n33077;
  assign n33097 = ~n3378 & ~n33096;
  assign n33098 = ~n3378 & ~n33097;
  assign n33099 = n3492 & ~n33098;
  assign n33100 = ~n3493 & ~n33099;
  assign n33101 = n3485 & ~n33100;
  assign n33102 = ~n3486 & ~n33101;
  assign n33103 = ~n3476 & ~n33102;
  assign n33104 = ~n3281 & ~n26724;
  assign n33105 = n3378 & ~n33104;
  assign n33106 = ~n26726 & ~n33105;
  assign n33107 = n3492 & ~n33106;
  assign n33108 = ~n3493 & ~n33107;
  assign n33109 = n3485 & ~n33108;
  assign n33110 = ~n3486 & ~n33109;
  assign n33111 = n3476 & ~n33110;
  assign n33112 = ~n33103 & ~n33111;
  assign n33113 = n3374 & ~n33112;
  assign n33114 = ~n33095 & ~n33113;
  assign n33115 = n3655 & ~n33114;
  assign n33116 = ~n24419 & ~n33073;
  assign n33117 = controllable_nhgrant0 & ~n33116;
  assign n33118 = ~n24376 & ~n33117;
  assign n33119 = ~n3281 & ~n33118;
  assign n33120 = ~n3783 & ~n33119;
  assign n33121 = ~n3378 & ~n33120;
  assign n33122 = ~n3378 & ~n33121;
  assign n33123 = n3492 & ~n33122;
  assign n33124 = ~n3493 & ~n33123;
  assign n33125 = n3485 & ~n33124;
  assign n33126 = ~n3486 & ~n33125;
  assign n33127 = ~n3476 & ~n33126;
  assign n33128 = ~n3281 & ~n26741;
  assign n33129 = n3378 & ~n33128;
  assign n33130 = ~n26743 & ~n33129;
  assign n33131 = n3492 & ~n33130;
  assign n33132 = ~n3493 & ~n33131;
  assign n33133 = n3485 & ~n33132;
  assign n33134 = ~n3486 & ~n33133;
  assign n33135 = n3476 & ~n33134;
  assign n33136 = ~n33127 & ~n33135;
  assign n33137 = ~n3374 & ~n33136;
  assign n33138 = ~n3950 & ~n33119;
  assign n33139 = ~n3378 & ~n33138;
  assign n33140 = ~n3378 & ~n33139;
  assign n33141 = n3492 & ~n33140;
  assign n33142 = ~n3493 & ~n33141;
  assign n33143 = n3485 & ~n33142;
  assign n33144 = ~n3486 & ~n33143;
  assign n33145 = ~n3476 & ~n33144;
  assign n33146 = ~n3281 & ~n26773;
  assign n33147 = n3378 & ~n33146;
  assign n33148 = ~n26775 & ~n33147;
  assign n33149 = n3492 & ~n33148;
  assign n33150 = ~n3493 & ~n33149;
  assign n33151 = n3485 & ~n33150;
  assign n33152 = ~n3486 & ~n33151;
  assign n33153 = n3476 & ~n33152;
  assign n33154 = ~n33145 & ~n33153;
  assign n33155 = n3374 & ~n33154;
  assign n33156 = ~n33137 & ~n33155;
  assign n33157 = ~n3655 & ~n33156;
  assign n33158 = ~n33115 & ~n33157;
  assign n33159 = n3652 & ~n33158;
  assign n33160 = ~n24466 & ~n33073;
  assign n33161 = controllable_nhgrant0 & ~n33160;
  assign n33162 = ~n24376 & ~n33161;
  assign n33163 = ~n3281 & ~n33162;
  assign n33164 = ~n3783 & ~n33163;
  assign n33165 = ~n3378 & ~n33164;
  assign n33166 = ~n3378 & ~n33165;
  assign n33167 = n3492 & ~n33166;
  assign n33168 = ~n3493 & ~n33167;
  assign n33169 = n3485 & ~n33168;
  assign n33170 = ~n3486 & ~n33169;
  assign n33171 = ~n3476 & ~n33170;
  assign n33172 = ~n3281 & ~n26792;
  assign n33173 = n3378 & ~n33172;
  assign n33174 = ~n26794 & ~n33173;
  assign n33175 = n3492 & ~n33174;
  assign n33176 = ~n3493 & ~n33175;
  assign n33177 = n3485 & ~n33176;
  assign n33178 = ~n3486 & ~n33177;
  assign n33179 = n3476 & ~n33178;
  assign n33180 = ~n33171 & ~n33179;
  assign n33181 = ~n3374 & ~n33180;
  assign n33182 = ~n3950 & ~n33163;
  assign n33183 = ~n3378 & ~n33182;
  assign n33184 = ~n3378 & ~n33183;
  assign n33185 = n3492 & ~n33184;
  assign n33186 = ~n3493 & ~n33185;
  assign n33187 = n3485 & ~n33186;
  assign n33188 = ~n3486 & ~n33187;
  assign n33189 = ~n3476 & ~n33188;
  assign n33190 = ~n3281 & ~n26824;
  assign n33191 = n3378 & ~n33190;
  assign n33192 = ~n26826 & ~n33191;
  assign n33193 = n3492 & ~n33192;
  assign n33194 = ~n3493 & ~n33193;
  assign n33195 = n3485 & ~n33194;
  assign n33196 = ~n3486 & ~n33195;
  assign n33197 = n3476 & ~n33196;
  assign n33198 = ~n33189 & ~n33197;
  assign n33199 = n3374 & ~n33198;
  assign n33200 = ~n33181 & ~n33199;
  assign n33201 = n3655 & ~n33200;
  assign n33202 = ~n24514 & ~n33073;
  assign n33203 = controllable_nhgrant0 & ~n33202;
  assign n33204 = ~n24376 & ~n33203;
  assign n33205 = ~n3281 & ~n33204;
  assign n33206 = ~n3783 & ~n33205;
  assign n33207 = ~n3378 & ~n33206;
  assign n33208 = ~n3378 & ~n33207;
  assign n33209 = n3492 & ~n33208;
  assign n33210 = ~n3493 & ~n33209;
  assign n33211 = n3485 & ~n33210;
  assign n33212 = ~n3486 & ~n33211;
  assign n33213 = ~n3476 & ~n33212;
  assign n33214 = ~n3281 & ~n26841;
  assign n33215 = n3378 & ~n33214;
  assign n33216 = ~n26843 & ~n33215;
  assign n33217 = n3492 & ~n33216;
  assign n33218 = ~n3493 & ~n33217;
  assign n33219 = n3485 & ~n33218;
  assign n33220 = ~n3486 & ~n33219;
  assign n33221 = n3476 & ~n33220;
  assign n33222 = ~n33213 & ~n33221;
  assign n33223 = ~n3374 & ~n33222;
  assign n33224 = ~n3950 & ~n33205;
  assign n33225 = ~n3378 & ~n33224;
  assign n33226 = ~n3378 & ~n33225;
  assign n33227 = n3492 & ~n33226;
  assign n33228 = ~n3493 & ~n33227;
  assign n33229 = n3485 & ~n33228;
  assign n33230 = ~n3486 & ~n33229;
  assign n33231 = ~n3476 & ~n33230;
  assign n33232 = ~n3281 & ~n26873;
  assign n33233 = n3378 & ~n33232;
  assign n33234 = ~n26875 & ~n33233;
  assign n33235 = n3492 & ~n33234;
  assign n33236 = ~n3493 & ~n33235;
  assign n33237 = n3485 & ~n33236;
  assign n33238 = ~n3486 & ~n33237;
  assign n33239 = n3476 & ~n33238;
  assign n33240 = ~n33231 & ~n33239;
  assign n33241 = n3374 & ~n33240;
  assign n33242 = ~n33223 & ~n33241;
  assign n33243 = ~n3655 & ~n33242;
  assign n33244 = ~n33201 & ~n33243;
  assign n33245 = ~n3652 & ~n33244;
  assign n33246 = ~n33159 & ~n33245;
  assign n33247 = ~n3368 & ~n33246;
  assign n33248 = n3492 & ~n26896;
  assign n33249 = n3492 & ~n33248;
  assign n33250 = n3485 & ~n33249;
  assign n33251 = n3485 & ~n33250;
  assign n33252 = n3476 & ~n33251;
  assign n33253 = n3476 & ~n33252;
  assign n33254 = ~n3374 & ~n33253;
  assign n33255 = n3492 & ~n27143;
  assign n33256 = n3492 & ~n33255;
  assign n33257 = n3485 & ~n33256;
  assign n33258 = n3485 & ~n33257;
  assign n33259 = n3476 & ~n33258;
  assign n33260 = n3476 & ~n33259;
  assign n33261 = n3374 & ~n33260;
  assign n33262 = ~n33254 & ~n33261;
  assign n33263 = n3655 & ~n33262;
  assign n33264 = n3492 & ~n27160;
  assign n33265 = n3492 & ~n33264;
  assign n33266 = n3485 & ~n33265;
  assign n33267 = n3485 & ~n33266;
  assign n33268 = n3476 & ~n33267;
  assign n33269 = n3476 & ~n33268;
  assign n33270 = ~n3374 & ~n33269;
  assign n33271 = n3492 & ~n27197;
  assign n33272 = n3492 & ~n33271;
  assign n33273 = n3485 & ~n33272;
  assign n33274 = n3485 & ~n33273;
  assign n33275 = n3476 & ~n33274;
  assign n33276 = n3476 & ~n33275;
  assign n33277 = n3374 & ~n33276;
  assign n33278 = ~n33270 & ~n33277;
  assign n33279 = ~n3655 & ~n33278;
  assign n33280 = ~n33263 & ~n33279;
  assign n33281 = n3652 & ~n33280;
  assign n33282 = n3492 & ~n27216;
  assign n33283 = n3492 & ~n33282;
  assign n33284 = n3485 & ~n33283;
  assign n33285 = n3485 & ~n33284;
  assign n33286 = n3476 & ~n33285;
  assign n33287 = n3476 & ~n33286;
  assign n33288 = ~n3374 & ~n33287;
  assign n33289 = n3492 & ~n27253;
  assign n33290 = n3492 & ~n33289;
  assign n33291 = n3485 & ~n33290;
  assign n33292 = n3485 & ~n33291;
  assign n33293 = n3476 & ~n33292;
  assign n33294 = n3476 & ~n33293;
  assign n33295 = n3374 & ~n33294;
  assign n33296 = ~n33288 & ~n33295;
  assign n33297 = n3655 & ~n33296;
  assign n33298 = n3492 & ~n27270;
  assign n33299 = n3492 & ~n33298;
  assign n33300 = n3485 & ~n33299;
  assign n33301 = n3485 & ~n33300;
  assign n33302 = n3476 & ~n33301;
  assign n33303 = n3476 & ~n33302;
  assign n33304 = ~n3374 & ~n33303;
  assign n33305 = n3492 & ~n27307;
  assign n33306 = n3492 & ~n33305;
  assign n33307 = n3485 & ~n33306;
  assign n33308 = n3485 & ~n33307;
  assign n33309 = n3476 & ~n33308;
  assign n33310 = n3476 & ~n33309;
  assign n33311 = n3374 & ~n33310;
  assign n33312 = ~n33304 & ~n33311;
  assign n33313 = ~n3655 & ~n33312;
  assign n33314 = ~n33297 & ~n33313;
  assign n33315 = ~n3652 & ~n33314;
  assign n33316 = ~n33281 & ~n33315;
  assign n33317 = n3368 & ~n33316;
  assign n33318 = ~n33247 & ~n33317;
  assign n33319 = ~n3362 & ~n33318;
  assign n33320 = ~n3362 & ~n33319;
  assign n33321 = ~n3359 & ~n33320;
  assign n33322 = ~n3359 & ~n33321;
  assign n33323 = n3356 & ~n33322;
  assign n33324 = n3492 & ~n26689;
  assign n33325 = ~n3631 & ~n33324;
  assign n33326 = n3485 & ~n33325;
  assign n33327 = ~n3630 & ~n33326;
  assign n33328 = ~n3374 & ~n33327;
  assign n33329 = n3492 & ~n26710;
  assign n33330 = ~n3631 & ~n33329;
  assign n33331 = n3485 & ~n33330;
  assign n33332 = ~n3630 & ~n33331;
  assign n33333 = ~n3476 & ~n33332;
  assign n33334 = n3492 & ~n26725;
  assign n33335 = ~n3631 & ~n33334;
  assign n33336 = n3485 & ~n33335;
  assign n33337 = ~n3630 & ~n33336;
  assign n33338 = n3476 & ~n33337;
  assign n33339 = ~n33333 & ~n33338;
  assign n33340 = n3374 & ~n33339;
  assign n33341 = ~n33328 & ~n33340;
  assign n33342 = n3655 & ~n33341;
  assign n33343 = n3492 & ~n26742;
  assign n33344 = ~n3631 & ~n33343;
  assign n33345 = n3485 & ~n33344;
  assign n33346 = ~n3630 & ~n33345;
  assign n33347 = ~n3374 & ~n33346;
  assign n33348 = n3492 & ~n26761;
  assign n33349 = ~n3631 & ~n33348;
  assign n33350 = n3485 & ~n33349;
  assign n33351 = ~n3630 & ~n33350;
  assign n33352 = ~n3476 & ~n33351;
  assign n33353 = n3492 & ~n26774;
  assign n33354 = ~n3631 & ~n33353;
  assign n33355 = n3485 & ~n33354;
  assign n33356 = ~n3630 & ~n33355;
  assign n33357 = n3476 & ~n33356;
  assign n33358 = ~n33352 & ~n33357;
  assign n33359 = n3374 & ~n33358;
  assign n33360 = ~n33347 & ~n33359;
  assign n33361 = ~n3655 & ~n33360;
  assign n33362 = ~n33342 & ~n33361;
  assign n33363 = n3652 & ~n33362;
  assign n33364 = n3492 & ~n26793;
  assign n33365 = ~n3631 & ~n33364;
  assign n33366 = n3485 & ~n33365;
  assign n33367 = ~n3630 & ~n33366;
  assign n33368 = ~n3374 & ~n33367;
  assign n33369 = n3492 & ~n26812;
  assign n33370 = ~n3631 & ~n33369;
  assign n33371 = n3485 & ~n33370;
  assign n33372 = ~n3630 & ~n33371;
  assign n33373 = ~n3476 & ~n33372;
  assign n33374 = n3492 & ~n26825;
  assign n33375 = ~n3631 & ~n33374;
  assign n33376 = n3485 & ~n33375;
  assign n33377 = ~n3630 & ~n33376;
  assign n33378 = n3476 & ~n33377;
  assign n33379 = ~n33373 & ~n33378;
  assign n33380 = n3374 & ~n33379;
  assign n33381 = ~n33368 & ~n33380;
  assign n33382 = n3655 & ~n33381;
  assign n33383 = n3492 & ~n26842;
  assign n33384 = ~n3631 & ~n33383;
  assign n33385 = n3485 & ~n33384;
  assign n33386 = ~n3630 & ~n33385;
  assign n33387 = ~n3374 & ~n33386;
  assign n33388 = n3492 & ~n26861;
  assign n33389 = ~n3631 & ~n33388;
  assign n33390 = n3485 & ~n33389;
  assign n33391 = ~n3630 & ~n33390;
  assign n33392 = ~n3476 & ~n33391;
  assign n33393 = n3492 & ~n26874;
  assign n33394 = ~n3631 & ~n33393;
  assign n33395 = n3485 & ~n33394;
  assign n33396 = ~n3630 & ~n33395;
  assign n33397 = n3476 & ~n33396;
  assign n33398 = ~n33392 & ~n33397;
  assign n33399 = n3374 & ~n33398;
  assign n33400 = ~n33387 & ~n33399;
  assign n33401 = ~n3655 & ~n33400;
  assign n33402 = ~n33382 & ~n33401;
  assign n33403 = ~n3652 & ~n33402;
  assign n33404 = ~n33363 & ~n33403;
  assign n33405 = ~n3368 & ~n33404;
  assign n33406 = ~n3374 & ~n33251;
  assign n33407 = n3492 & ~n26930;
  assign n33408 = n3492 & ~n33407;
  assign n33409 = n3485 & ~n33408;
  assign n33410 = n3485 & ~n33409;
  assign n33411 = ~n3476 & ~n33410;
  assign n33412 = ~n33259 & ~n33411;
  assign n33413 = n3374 & ~n33412;
  assign n33414 = ~n33406 & ~n33413;
  assign n33415 = n3655 & ~n33414;
  assign n33416 = ~n3374 & ~n33267;
  assign n33417 = n3492 & ~n27179;
  assign n33418 = n3492 & ~n33417;
  assign n33419 = n3485 & ~n33418;
  assign n33420 = n3485 & ~n33419;
  assign n33421 = ~n3476 & ~n33420;
  assign n33422 = ~n33275 & ~n33421;
  assign n33423 = n3374 & ~n33422;
  assign n33424 = ~n33416 & ~n33423;
  assign n33425 = ~n3655 & ~n33424;
  assign n33426 = ~n33415 & ~n33425;
  assign n33427 = n3652 & ~n33426;
  assign n33428 = ~n3374 & ~n33285;
  assign n33429 = n3492 & ~n27235;
  assign n33430 = n3492 & ~n33429;
  assign n33431 = n3485 & ~n33430;
  assign n33432 = n3485 & ~n33431;
  assign n33433 = ~n3476 & ~n33432;
  assign n33434 = ~n33293 & ~n33433;
  assign n33435 = n3374 & ~n33434;
  assign n33436 = ~n33428 & ~n33435;
  assign n33437 = n3655 & ~n33436;
  assign n33438 = ~n3374 & ~n33301;
  assign n33439 = n3492 & ~n27289;
  assign n33440 = n3492 & ~n33439;
  assign n33441 = n3485 & ~n33440;
  assign n33442 = n3485 & ~n33441;
  assign n33443 = ~n3476 & ~n33442;
  assign n33444 = ~n33309 & ~n33443;
  assign n33445 = n3374 & ~n33444;
  assign n33446 = ~n33438 & ~n33445;
  assign n33447 = ~n3655 & ~n33446;
  assign n33448 = ~n33437 & ~n33447;
  assign n33449 = ~n3652 & ~n33448;
  assign n33450 = ~n33427 & ~n33449;
  assign n33451 = n3368 & ~n33450;
  assign n33452 = ~n33405 & ~n33451;
  assign n33453 = n3362 & ~n33452;
  assign n33454 = ~n3476 & ~n33327;
  assign n33455 = ~n26202 & ~n33326;
  assign n33456 = n3476 & ~n33455;
  assign n33457 = ~n33454 & ~n33456;
  assign n33458 = ~n3374 & ~n33457;
  assign n33459 = ~n26202 & ~n33336;
  assign n33460 = n3476 & ~n33459;
  assign n33461 = ~n33333 & ~n33460;
  assign n33462 = n3374 & ~n33461;
  assign n33463 = ~n33458 & ~n33462;
  assign n33464 = n3655 & ~n33463;
  assign n33465 = ~n3476 & ~n33346;
  assign n33466 = ~n26299 & ~n33345;
  assign n33467 = n3476 & ~n33466;
  assign n33468 = ~n33465 & ~n33467;
  assign n33469 = ~n3374 & ~n33468;
  assign n33470 = ~n26299 & ~n33355;
  assign n33471 = n3476 & ~n33470;
  assign n33472 = ~n33352 & ~n33471;
  assign n33473 = n3374 & ~n33472;
  assign n33474 = ~n33469 & ~n33473;
  assign n33475 = ~n3655 & ~n33474;
  assign n33476 = ~n33464 & ~n33475;
  assign n33477 = n3652 & ~n33476;
  assign n33478 = ~n3476 & ~n33367;
  assign n33479 = ~n26398 & ~n33366;
  assign n33480 = n3476 & ~n33479;
  assign n33481 = ~n33478 & ~n33480;
  assign n33482 = ~n3374 & ~n33481;
  assign n33483 = ~n26398 & ~n33376;
  assign n33484 = n3476 & ~n33483;
  assign n33485 = ~n33373 & ~n33484;
  assign n33486 = n3374 & ~n33485;
  assign n33487 = ~n33482 & ~n33486;
  assign n33488 = n3655 & ~n33487;
  assign n33489 = ~n3476 & ~n33386;
  assign n33490 = ~n26439 & ~n33385;
  assign n33491 = n3476 & ~n33490;
  assign n33492 = ~n33489 & ~n33491;
  assign n33493 = ~n3374 & ~n33492;
  assign n33494 = ~n26439 & ~n33395;
  assign n33495 = n3476 & ~n33494;
  assign n33496 = ~n33392 & ~n33495;
  assign n33497 = n3374 & ~n33496;
  assign n33498 = ~n33493 & ~n33497;
  assign n33499 = ~n3655 & ~n33498;
  assign n33500 = ~n33488 & ~n33499;
  assign n33501 = ~n3652 & ~n33500;
  assign n33502 = ~n33477 & ~n33501;
  assign n33503 = ~n3368 & ~n33502;
  assign n33504 = ~n3476 & ~n33251;
  assign n33505 = ~n8525 & ~n33250;
  assign n33506 = n3476 & ~n33505;
  assign n33507 = ~n33504 & ~n33506;
  assign n33508 = ~n3374 & ~n33507;
  assign n33509 = ~n26479 & ~n33257;
  assign n33510 = n3476 & ~n33509;
  assign n33511 = ~n33411 & ~n33510;
  assign n33512 = n3374 & ~n33511;
  assign n33513 = ~n33508 & ~n33512;
  assign n33514 = n3655 & ~n33513;
  assign n33515 = ~n3476 & ~n33267;
  assign n33516 = ~n8525 & ~n33266;
  assign n33517 = n3476 & ~n33516;
  assign n33518 = ~n33515 & ~n33517;
  assign n33519 = ~n3374 & ~n33518;
  assign n33520 = ~n26506 & ~n33273;
  assign n33521 = n3476 & ~n33520;
  assign n33522 = ~n33421 & ~n33521;
  assign n33523 = n3374 & ~n33522;
  assign n33524 = ~n33519 & ~n33523;
  assign n33525 = ~n3655 & ~n33524;
  assign n33526 = ~n33514 & ~n33525;
  assign n33527 = n3652 & ~n33526;
  assign n33528 = ~n3476 & ~n33285;
  assign n33529 = ~n8525 & ~n33284;
  assign n33530 = n3476 & ~n33529;
  assign n33531 = ~n33528 & ~n33530;
  assign n33532 = ~n3374 & ~n33531;
  assign n33533 = ~n26535 & ~n33291;
  assign n33534 = n3476 & ~n33533;
  assign n33535 = ~n33433 & ~n33534;
  assign n33536 = n3374 & ~n33535;
  assign n33537 = ~n33532 & ~n33536;
  assign n33538 = n3655 & ~n33537;
  assign n33539 = ~n3476 & ~n33301;
  assign n33540 = ~n8525 & ~n33300;
  assign n33541 = n3476 & ~n33540;
  assign n33542 = ~n33539 & ~n33541;
  assign n33543 = ~n3374 & ~n33542;
  assign n33544 = ~n26562 & ~n33307;
  assign n33545 = n3476 & ~n33544;
  assign n33546 = ~n33443 & ~n33545;
  assign n33547 = n3374 & ~n33546;
  assign n33548 = ~n33543 & ~n33547;
  assign n33549 = ~n3655 & ~n33548;
  assign n33550 = ~n33538 & ~n33549;
  assign n33551 = ~n3652 & ~n33550;
  assign n33552 = ~n33527 & ~n33551;
  assign n33553 = n3368 & ~n33552;
  assign n33554 = ~n33503 & ~n33553;
  assign n33555 = ~n3362 & ~n33554;
  assign n33556 = ~n33453 & ~n33555;
  assign n33557 = n3359 & ~n33556;
  assign n33558 = ~n26580 & ~n33326;
  assign n33559 = n3476 & ~n33558;
  assign n33560 = ~n33454 & ~n33559;
  assign n33561 = ~n3374 & ~n33560;
  assign n33562 = ~n26580 & ~n33336;
  assign n33563 = n3476 & ~n33562;
  assign n33564 = ~n33333 & ~n33563;
  assign n33565 = n3374 & ~n33564;
  assign n33566 = ~n33561 & ~n33565;
  assign n33567 = n3655 & ~n33566;
  assign n33568 = ~n26591 & ~n33345;
  assign n33569 = n3476 & ~n33568;
  assign n33570 = ~n33465 & ~n33569;
  assign n33571 = ~n3374 & ~n33570;
  assign n33572 = ~n26591 & ~n33355;
  assign n33573 = n3476 & ~n33572;
  assign n33574 = ~n33352 & ~n33573;
  assign n33575 = n3374 & ~n33574;
  assign n33576 = ~n33571 & ~n33575;
  assign n33577 = ~n3655 & ~n33576;
  assign n33578 = ~n33567 & ~n33577;
  assign n33579 = n3652 & ~n33578;
  assign n33580 = ~n26604 & ~n33366;
  assign n33581 = n3476 & ~n33580;
  assign n33582 = ~n33478 & ~n33581;
  assign n33583 = ~n3374 & ~n33582;
  assign n33584 = ~n26604 & ~n33376;
  assign n33585 = n3476 & ~n33584;
  assign n33586 = ~n33373 & ~n33585;
  assign n33587 = n3374 & ~n33586;
  assign n33588 = ~n33583 & ~n33587;
  assign n33589 = n3655 & ~n33588;
  assign n33590 = ~n26615 & ~n33385;
  assign n33591 = n3476 & ~n33590;
  assign n33592 = ~n33489 & ~n33591;
  assign n33593 = ~n3374 & ~n33592;
  assign n33594 = ~n26615 & ~n33395;
  assign n33595 = n3476 & ~n33594;
  assign n33596 = ~n33392 & ~n33595;
  assign n33597 = n3374 & ~n33596;
  assign n33598 = ~n33593 & ~n33597;
  assign n33599 = ~n3655 & ~n33598;
  assign n33600 = ~n33589 & ~n33599;
  assign n33601 = ~n3652 & ~n33600;
  assign n33602 = ~n33579 & ~n33601;
  assign n33603 = ~n3368 & ~n33602;
  assign n33604 = ~n8689 & ~n33250;
  assign n33605 = n3476 & ~n33604;
  assign n33606 = ~n33504 & ~n33605;
  assign n33607 = ~n3374 & ~n33606;
  assign n33608 = ~n26634 & ~n33257;
  assign n33609 = n3476 & ~n33608;
  assign n33610 = ~n33411 & ~n33609;
  assign n33611 = n3374 & ~n33610;
  assign n33612 = ~n33607 & ~n33611;
  assign n33613 = n3655 & ~n33612;
  assign n33614 = ~n8689 & ~n33266;
  assign n33615 = n3476 & ~n33614;
  assign n33616 = ~n33515 & ~n33615;
  assign n33617 = ~n3374 & ~n33616;
  assign n33618 = ~n26645 & ~n33273;
  assign n33619 = n3476 & ~n33618;
  assign n33620 = ~n33421 & ~n33619;
  assign n33621 = n3374 & ~n33620;
  assign n33622 = ~n33617 & ~n33621;
  assign n33623 = ~n3655 & ~n33622;
  assign n33624 = ~n33613 & ~n33623;
  assign n33625 = n3652 & ~n33624;
  assign n33626 = ~n8689 & ~n33284;
  assign n33627 = n3476 & ~n33626;
  assign n33628 = ~n33528 & ~n33627;
  assign n33629 = ~n3374 & ~n33628;
  assign n33630 = ~n26658 & ~n33291;
  assign n33631 = n3476 & ~n33630;
  assign n33632 = ~n33433 & ~n33631;
  assign n33633 = n3374 & ~n33632;
  assign n33634 = ~n33629 & ~n33633;
  assign n33635 = n3655 & ~n33634;
  assign n33636 = ~n8689 & ~n33300;
  assign n33637 = n3476 & ~n33636;
  assign n33638 = ~n33539 & ~n33637;
  assign n33639 = ~n3374 & ~n33638;
  assign n33640 = ~n26669 & ~n33307;
  assign n33641 = n3476 & ~n33640;
  assign n33642 = ~n33443 & ~n33641;
  assign n33643 = n3374 & ~n33642;
  assign n33644 = ~n33639 & ~n33643;
  assign n33645 = ~n3655 & ~n33644;
  assign n33646 = ~n33635 & ~n33645;
  assign n33647 = ~n3652 & ~n33646;
  assign n33648 = ~n33625 & ~n33647;
  assign n33649 = n3368 & ~n33648;
  assign n33650 = ~n33603 & ~n33649;
  assign n33651 = n3362 & ~n33650;
  assign n33652 = ~n26200 & ~n33324;
  assign n33653 = n3485 & ~n33652;
  assign n33654 = ~n26580 & ~n33653;
  assign n33655 = n3476 & ~n33654;
  assign n33656 = ~n33454 & ~n33655;
  assign n33657 = ~n3374 & ~n33656;
  assign n33658 = ~n26200 & ~n33334;
  assign n33659 = n3485 & ~n33658;
  assign n33660 = ~n26580 & ~n33659;
  assign n33661 = n3476 & ~n33660;
  assign n33662 = ~n33333 & ~n33661;
  assign n33663 = n3374 & ~n33662;
  assign n33664 = ~n33657 & ~n33663;
  assign n33665 = n3655 & ~n33664;
  assign n33666 = ~n26297 & ~n33343;
  assign n33667 = n3485 & ~n33666;
  assign n33668 = ~n26591 & ~n33667;
  assign n33669 = n3476 & ~n33668;
  assign n33670 = ~n33465 & ~n33669;
  assign n33671 = ~n3374 & ~n33670;
  assign n33672 = ~n26297 & ~n33353;
  assign n33673 = n3485 & ~n33672;
  assign n33674 = ~n26591 & ~n33673;
  assign n33675 = n3476 & ~n33674;
  assign n33676 = ~n33352 & ~n33675;
  assign n33677 = n3374 & ~n33676;
  assign n33678 = ~n33671 & ~n33677;
  assign n33679 = ~n3655 & ~n33678;
  assign n33680 = ~n33665 & ~n33679;
  assign n33681 = n3652 & ~n33680;
  assign n33682 = ~n26396 & ~n33364;
  assign n33683 = n3485 & ~n33682;
  assign n33684 = ~n26604 & ~n33683;
  assign n33685 = n3476 & ~n33684;
  assign n33686 = ~n33478 & ~n33685;
  assign n33687 = ~n3374 & ~n33686;
  assign n33688 = ~n26396 & ~n33374;
  assign n33689 = n3485 & ~n33688;
  assign n33690 = ~n26604 & ~n33689;
  assign n33691 = n3476 & ~n33690;
  assign n33692 = ~n33373 & ~n33691;
  assign n33693 = n3374 & ~n33692;
  assign n33694 = ~n33687 & ~n33693;
  assign n33695 = n3655 & ~n33694;
  assign n33696 = ~n26437 & ~n33383;
  assign n33697 = n3485 & ~n33696;
  assign n33698 = ~n26615 & ~n33697;
  assign n33699 = n3476 & ~n33698;
  assign n33700 = ~n33489 & ~n33699;
  assign n33701 = ~n3374 & ~n33700;
  assign n33702 = ~n26437 & ~n33393;
  assign n33703 = n3485 & ~n33702;
  assign n33704 = ~n26615 & ~n33703;
  assign n33705 = n3476 & ~n33704;
  assign n33706 = ~n33392 & ~n33705;
  assign n33707 = n3374 & ~n33706;
  assign n33708 = ~n33701 & ~n33707;
  assign n33709 = ~n3655 & ~n33708;
  assign n33710 = ~n33695 & ~n33709;
  assign n33711 = ~n3652 & ~n33710;
  assign n33712 = ~n33681 & ~n33711;
  assign n33713 = ~n3368 & ~n33712;
  assign n33714 = ~n8523 & ~n33248;
  assign n33715 = n3485 & ~n33714;
  assign n33716 = ~n8689 & ~n33715;
  assign n33717 = n3476 & ~n33716;
  assign n33718 = ~n33504 & ~n33717;
  assign n33719 = ~n3374 & ~n33718;
  assign n33720 = ~n26477 & ~n33255;
  assign n33721 = n3485 & ~n33720;
  assign n33722 = ~n26634 & ~n33721;
  assign n33723 = n3476 & ~n33722;
  assign n33724 = ~n33411 & ~n33723;
  assign n33725 = n3374 & ~n33724;
  assign n33726 = ~n33719 & ~n33725;
  assign n33727 = n3655 & ~n33726;
  assign n33728 = ~n8523 & ~n33264;
  assign n33729 = n3485 & ~n33728;
  assign n33730 = ~n8689 & ~n33729;
  assign n33731 = n3476 & ~n33730;
  assign n33732 = ~n33515 & ~n33731;
  assign n33733 = ~n3374 & ~n33732;
  assign n33734 = ~n26504 & ~n33271;
  assign n33735 = n3485 & ~n33734;
  assign n33736 = ~n26645 & ~n33735;
  assign n33737 = n3476 & ~n33736;
  assign n33738 = ~n33421 & ~n33737;
  assign n33739 = n3374 & ~n33738;
  assign n33740 = ~n33733 & ~n33739;
  assign n33741 = ~n3655 & ~n33740;
  assign n33742 = ~n33727 & ~n33741;
  assign n33743 = n3652 & ~n33742;
  assign n33744 = ~n8523 & ~n33282;
  assign n33745 = n3485 & ~n33744;
  assign n33746 = ~n8689 & ~n33745;
  assign n33747 = n3476 & ~n33746;
  assign n33748 = ~n33528 & ~n33747;
  assign n33749 = ~n3374 & ~n33748;
  assign n33750 = ~n26533 & ~n33289;
  assign n33751 = n3485 & ~n33750;
  assign n33752 = ~n26658 & ~n33751;
  assign n33753 = n3476 & ~n33752;
  assign n33754 = ~n33433 & ~n33753;
  assign n33755 = n3374 & ~n33754;
  assign n33756 = ~n33749 & ~n33755;
  assign n33757 = n3655 & ~n33756;
  assign n33758 = ~n8523 & ~n33298;
  assign n33759 = n3485 & ~n33758;
  assign n33760 = ~n8689 & ~n33759;
  assign n33761 = n3476 & ~n33760;
  assign n33762 = ~n33539 & ~n33761;
  assign n33763 = ~n3374 & ~n33762;
  assign n33764 = ~n26560 & ~n33305;
  assign n33765 = n3485 & ~n33764;
  assign n33766 = ~n26669 & ~n33765;
  assign n33767 = n3476 & ~n33766;
  assign n33768 = ~n33443 & ~n33767;
  assign n33769 = n3374 & ~n33768;
  assign n33770 = ~n33763 & ~n33769;
  assign n33771 = ~n3655 & ~n33770;
  assign n33772 = ~n33757 & ~n33771;
  assign n33773 = ~n3652 & ~n33772;
  assign n33774 = ~n33743 & ~n33773;
  assign n33775 = n3368 & ~n33774;
  assign n33776 = ~n33713 & ~n33775;
  assign n33777 = ~n3362 & ~n33776;
  assign n33778 = ~n33651 & ~n33777;
  assign n33779 = ~n3359 & ~n33778;
  assign n33780 = ~n33557 & ~n33779;
  assign n33781 = ~n3356 & ~n33780;
  assign n33782 = ~n33323 & ~n33781;
  assign n33783 = ~n3345 & ~n33782;
  assign n33784 = ~n3378 & ~n26690;
  assign n33785 = n3492 & ~n33784;
  assign n33786 = ~n3493 & ~n33785;
  assign n33787 = n3485 & ~n33786;
  assign n33788 = ~n3486 & ~n33787;
  assign n33789 = ~n3476 & ~n33788;
  assign n33790 = ~n3378 & ~n26199;
  assign n33791 = ~n3378 & ~n33790;
  assign n33792 = ~n3485 & ~n33791;
  assign n33793 = ~n3492 & ~n33791;
  assign n33794 = ~n33785 & ~n33793;
  assign n33795 = n3485 & ~n33794;
  assign n33796 = ~n33792 & ~n33795;
  assign n33797 = n3476 & ~n33796;
  assign n33798 = ~n33789 & ~n33797;
  assign n33799 = ~n3374 & ~n33798;
  assign n33800 = ~n3281 & ~n26709;
  assign n33801 = n3378 & ~n33800;
  assign n33802 = ~n26711 & ~n33801;
  assign n33803 = n3492 & ~n33802;
  assign n33804 = ~n25115 & ~n33803;
  assign n33805 = n3485 & ~n33804;
  assign n33806 = ~n25114 & ~n33805;
  assign n33807 = ~n3476 & ~n33806;
  assign n33808 = n3378 & ~n26476;
  assign n33809 = ~n33790 & ~n33808;
  assign n33810 = ~n3485 & ~n33809;
  assign n33811 = ~n3492 & ~n33809;
  assign n33812 = ~n33107 & ~n33811;
  assign n33813 = n3485 & ~n33812;
  assign n33814 = ~n33810 & ~n33813;
  assign n33815 = n3476 & ~n33814;
  assign n33816 = ~n33807 & ~n33815;
  assign n33817 = n3374 & ~n33816;
  assign n33818 = ~n33799 & ~n33817;
  assign n33819 = n3655 & ~n33818;
  assign n33820 = ~n3378 & ~n26743;
  assign n33821 = n3492 & ~n33820;
  assign n33822 = ~n3493 & ~n33821;
  assign n33823 = n3485 & ~n33822;
  assign n33824 = ~n3486 & ~n33823;
  assign n33825 = ~n3476 & ~n33824;
  assign n33826 = ~n3378 & ~n26296;
  assign n33827 = ~n3378 & ~n33826;
  assign n33828 = ~n3485 & ~n33827;
  assign n33829 = ~n3492 & ~n33827;
  assign n33830 = ~n33821 & ~n33829;
  assign n33831 = n3485 & ~n33830;
  assign n33832 = ~n33828 & ~n33831;
  assign n33833 = n3476 & ~n33832;
  assign n33834 = ~n33825 & ~n33833;
  assign n33835 = ~n3374 & ~n33834;
  assign n33836 = ~n3281 & ~n26760;
  assign n33837 = n3378 & ~n33836;
  assign n33838 = ~n26762 & ~n33837;
  assign n33839 = n3492 & ~n33838;
  assign n33840 = ~n25115 & ~n33839;
  assign n33841 = n3485 & ~n33840;
  assign n33842 = ~n25114 & ~n33841;
  assign n33843 = ~n3476 & ~n33842;
  assign n33844 = n3378 & ~n26503;
  assign n33845 = ~n33826 & ~n33844;
  assign n33846 = ~n3485 & ~n33845;
  assign n33847 = ~n3492 & ~n33845;
  assign n33848 = ~n33149 & ~n33847;
  assign n33849 = n3485 & ~n33848;
  assign n33850 = ~n33846 & ~n33849;
  assign n33851 = n3476 & ~n33850;
  assign n33852 = ~n33843 & ~n33851;
  assign n33853 = n3374 & ~n33852;
  assign n33854 = ~n33835 & ~n33853;
  assign n33855 = ~n3655 & ~n33854;
  assign n33856 = ~n33819 & ~n33855;
  assign n33857 = n3652 & ~n33856;
  assign n33858 = ~n3378 & ~n26794;
  assign n33859 = n3492 & ~n33858;
  assign n33860 = ~n3493 & ~n33859;
  assign n33861 = n3485 & ~n33860;
  assign n33862 = ~n3486 & ~n33861;
  assign n33863 = ~n3476 & ~n33862;
  assign n33864 = ~n3378 & ~n26395;
  assign n33865 = ~n3378 & ~n33864;
  assign n33866 = ~n3485 & ~n33865;
  assign n33867 = ~n3492 & ~n33865;
  assign n33868 = ~n33859 & ~n33867;
  assign n33869 = n3485 & ~n33868;
  assign n33870 = ~n33866 & ~n33869;
  assign n33871 = n3476 & ~n33870;
  assign n33872 = ~n33863 & ~n33871;
  assign n33873 = ~n3374 & ~n33872;
  assign n33874 = ~n3281 & ~n26811;
  assign n33875 = n3378 & ~n33874;
  assign n33876 = ~n26813 & ~n33875;
  assign n33877 = n3492 & ~n33876;
  assign n33878 = ~n25115 & ~n33877;
  assign n33879 = n3485 & ~n33878;
  assign n33880 = ~n25114 & ~n33879;
  assign n33881 = ~n3476 & ~n33880;
  assign n33882 = n3378 & ~n26532;
  assign n33883 = ~n33864 & ~n33882;
  assign n33884 = ~n3485 & ~n33883;
  assign n33885 = ~n3492 & ~n33883;
  assign n33886 = ~n33193 & ~n33885;
  assign n33887 = n3485 & ~n33886;
  assign n33888 = ~n33884 & ~n33887;
  assign n33889 = n3476 & ~n33888;
  assign n33890 = ~n33881 & ~n33889;
  assign n33891 = n3374 & ~n33890;
  assign n33892 = ~n33873 & ~n33891;
  assign n33893 = n3655 & ~n33892;
  assign n33894 = ~n3378 & ~n26843;
  assign n33895 = n3492 & ~n33894;
  assign n33896 = ~n3493 & ~n33895;
  assign n33897 = n3485 & ~n33896;
  assign n33898 = ~n3486 & ~n33897;
  assign n33899 = ~n3476 & ~n33898;
  assign n33900 = ~n3378 & ~n26436;
  assign n33901 = ~n3378 & ~n33900;
  assign n33902 = ~n3485 & ~n33901;
  assign n33903 = ~n3492 & ~n33901;
  assign n33904 = ~n33895 & ~n33903;
  assign n33905 = n3485 & ~n33904;
  assign n33906 = ~n33902 & ~n33905;
  assign n33907 = n3476 & ~n33906;
  assign n33908 = ~n33899 & ~n33907;
  assign n33909 = ~n3374 & ~n33908;
  assign n33910 = ~n3281 & ~n26860;
  assign n33911 = n3378 & ~n33910;
  assign n33912 = ~n26862 & ~n33911;
  assign n33913 = n3492 & ~n33912;
  assign n33914 = ~n25115 & ~n33913;
  assign n33915 = n3485 & ~n33914;
  assign n33916 = ~n25114 & ~n33915;
  assign n33917 = ~n3476 & ~n33916;
  assign n33918 = n3378 & ~n26559;
  assign n33919 = ~n33900 & ~n33918;
  assign n33920 = ~n3485 & ~n33919;
  assign n33921 = ~n3492 & ~n33919;
  assign n33922 = ~n33235 & ~n33921;
  assign n33923 = n3485 & ~n33922;
  assign n33924 = ~n33920 & ~n33923;
  assign n33925 = n3476 & ~n33924;
  assign n33926 = ~n33917 & ~n33925;
  assign n33927 = n3374 & ~n33926;
  assign n33928 = ~n33909 & ~n33927;
  assign n33929 = ~n3655 & ~n33928;
  assign n33930 = ~n33893 & ~n33929;
  assign n33931 = ~n3652 & ~n33930;
  assign n33932 = ~n33857 & ~n33931;
  assign n33933 = ~n3368 & ~n33932;
  assign n33934 = ~n3378 & ~n26897;
  assign n33935 = n3492 & ~n33934;
  assign n33936 = n3492 & ~n33935;
  assign n33937 = n3485 & ~n33936;
  assign n33938 = n3485 & ~n33937;
  assign n33939 = ~n3476 & ~n33938;
  assign n33940 = ~n25259 & ~n33935;
  assign n33941 = n3485 & ~n33940;
  assign n33942 = ~n25258 & ~n33941;
  assign n33943 = n3476 & ~n33942;
  assign n33944 = ~n33939 & ~n33943;
  assign n33945 = ~n3374 & ~n33944;
  assign n33946 = ~n33725 & ~n33945;
  assign n33947 = n3655 & ~n33946;
  assign n33948 = ~n3378 & ~n27161;
  assign n33949 = n3492 & ~n33948;
  assign n33950 = n3492 & ~n33949;
  assign n33951 = n3485 & ~n33950;
  assign n33952 = n3485 & ~n33951;
  assign n33953 = ~n3476 & ~n33952;
  assign n33954 = ~n25259 & ~n33949;
  assign n33955 = n3485 & ~n33954;
  assign n33956 = ~n25258 & ~n33955;
  assign n33957 = n3476 & ~n33956;
  assign n33958 = ~n33953 & ~n33957;
  assign n33959 = ~n3374 & ~n33958;
  assign n33960 = ~n33739 & ~n33959;
  assign n33961 = ~n3655 & ~n33960;
  assign n33962 = ~n33947 & ~n33961;
  assign n33963 = n3652 & ~n33962;
  assign n33964 = ~n3378 & ~n27217;
  assign n33965 = n3492 & ~n33964;
  assign n33966 = n3492 & ~n33965;
  assign n33967 = n3485 & ~n33966;
  assign n33968 = n3485 & ~n33967;
  assign n33969 = ~n3476 & ~n33968;
  assign n33970 = ~n25259 & ~n33965;
  assign n33971 = n3485 & ~n33970;
  assign n33972 = ~n25258 & ~n33971;
  assign n33973 = n3476 & ~n33972;
  assign n33974 = ~n33969 & ~n33973;
  assign n33975 = ~n3374 & ~n33974;
  assign n33976 = ~n33755 & ~n33975;
  assign n33977 = n3655 & ~n33976;
  assign n33978 = ~n3378 & ~n27271;
  assign n33979 = n3492 & ~n33978;
  assign n33980 = n3492 & ~n33979;
  assign n33981 = n3485 & ~n33980;
  assign n33982 = n3485 & ~n33981;
  assign n33983 = ~n3476 & ~n33982;
  assign n33984 = ~n25259 & ~n33979;
  assign n33985 = n3485 & ~n33984;
  assign n33986 = ~n25258 & ~n33985;
  assign n33987 = n3476 & ~n33986;
  assign n33988 = ~n33983 & ~n33987;
  assign n33989 = ~n3374 & ~n33988;
  assign n33990 = ~n33769 & ~n33989;
  assign n33991 = ~n3655 & ~n33990;
  assign n33992 = ~n33977 & ~n33991;
  assign n33993 = ~n3652 & ~n33992;
  assign n33994 = ~n33963 & ~n33993;
  assign n33995 = n3368 & ~n33994;
  assign n33996 = ~n33933 & ~n33995;
  assign n33997 = ~n3362 & ~n33996;
  assign n33998 = ~n3362 & ~n33997;
  assign n33999 = ~n3359 & ~n33998;
  assign n34000 = ~n3359 & ~n33999;
  assign n34001 = n3356 & ~n34000;
  assign n34002 = ~n3356 & ~n33776;
  assign n34003 = ~n34001 & ~n34002;
  assign n34004 = n3345 & ~n34003;
  assign n34005 = ~n33783 & ~n34004;
  assign n34006 = n3341 & ~n34005;
  assign n34007 = ~n33072 & ~n34006;
  assign n34008 = n3337 & ~n34007;
  assign n34009 = ~n30306 & ~n34008;
  assign n34010 = ~n3280 & ~n34009;
  assign n34011 = ~n25330 & ~n34010;
  assign n34012 = n3277 & n34011;
  assign n34013 = n3277 & ~n34012;
  assign n34014 = n3266 & ~n34013;
  assign n34015 = i_hlock4 & ~n5210;
  assign n34016 = ~i_hlock4 & ~n5216;
  assign n34017 = ~n34015 & ~n34016;
  assign n34018 = controllable_hgrant4 & ~n34017;
  assign n34019 = ~n3725 & ~n34018;
  assign n34020 = ~controllable_hgrant2 & ~n34019;
  assign n34021 = ~n3706 & ~n34020;
  assign n34022 = ~controllable_hmaster0 & ~n34021;
  assign n34023 = ~controllable_hmaster0 & ~n34022;
  assign n34024 = ~controllable_hmaster1 & ~n34023;
  assign n34025 = ~controllable_hmaster1 & ~n34024;
  assign n34026 = i_hbusreq3 & ~n34025;
  assign n34027 = i_hbusreq2 & ~n34019;
  assign n34028 = i_hbusreq4 & ~n34017;
  assign n34029 = i_hlock4 & ~n6620;
  assign n34030 = ~i_hlock4 & ~n6634;
  assign n34031 = ~n34029 & ~n34030;
  assign n34032 = ~i_hbusreq4 & ~n34031;
  assign n34033 = ~n34028 & ~n34032;
  assign n34034 = controllable_hgrant4 & ~n34033;
  assign n34035 = ~n3761 & ~n34034;
  assign n34036 = ~i_hbusreq2 & ~n34035;
  assign n34037 = ~n34027 & ~n34036;
  assign n34038 = ~controllable_hgrant2 & ~n34037;
  assign n34039 = ~n3734 & ~n34038;
  assign n34040 = ~controllable_hmaster0 & ~n34039;
  assign n34041 = ~controllable_hmaster0 & ~n34040;
  assign n34042 = ~controllable_hmaster1 & ~n34041;
  assign n34043 = ~controllable_hmaster1 & ~n34042;
  assign n34044 = ~i_hbusreq3 & ~n34043;
  assign n34045 = ~n34026 & ~n34044;
  assign n34046 = controllable_hmaster2 & ~n34045;
  assign n34047 = controllable_hmaster2 & ~n34046;
  assign n34048 = ~controllable_hgrant3 & ~n34047;
  assign n34049 = ~n3705 & ~n34048;
  assign n34050 = controllable_nhgrant0 & ~n34049;
  assign n34051 = ~n3778 & ~n34050;
  assign n34052 = ~n3281 & ~n34051;
  assign n34053 = ~n3281 & ~n34052;
  assign n34054 = n3378 & ~n34053;
  assign n34055 = controllable_hgrant4 & ~n3849;
  assign n34056 = ~n3421 & ~n34055;
  assign n34057 = ~controllable_hgrant2 & ~n34056;
  assign n34058 = ~n3410 & ~n34057;
  assign n34059 = controllable_hmaster1 & ~n34058;
  assign n34060 = controllable_hmaster0 & ~n34058;
  assign n34061 = ~n34022 & ~n34060;
  assign n34062 = ~controllable_hmaster1 & ~n34061;
  assign n34063 = ~n34059 & ~n34062;
  assign n34064 = i_hbusreq3 & ~n34063;
  assign n34065 = i_hbusreq2 & ~n34056;
  assign n34066 = controllable_hgrant4 & ~n14394;
  assign n34067 = ~n3448 & ~n34066;
  assign n34068 = ~i_hbusreq2 & ~n34067;
  assign n34069 = ~n34065 & ~n34068;
  assign n34070 = ~controllable_hgrant2 & ~n34069;
  assign n34071 = ~n3431 & ~n34070;
  assign n34072 = controllable_hmaster1 & ~n34071;
  assign n34073 = controllable_hmaster0 & ~n34071;
  assign n34074 = ~n34040 & ~n34073;
  assign n34075 = ~controllable_hmaster1 & ~n34074;
  assign n34076 = ~n34072 & ~n34075;
  assign n34077 = ~i_hbusreq3 & ~n34076;
  assign n34078 = ~n34064 & ~n34077;
  assign n34079 = controllable_hmaster2 & ~n34078;
  assign n34080 = controllable_hmaster2 & ~n34079;
  assign n34081 = ~controllable_hgrant3 & ~n34080;
  assign n34082 = ~n3795 & ~n34081;
  assign n34083 = controllable_nhgrant0 & ~n34082;
  assign n34084 = ~n3810 & ~n34083;
  assign n34085 = ~n3281 & ~n34084;
  assign n34086 = ~n3783 & ~n34085;
  assign n34087 = ~n3378 & ~n34086;
  assign n34088 = ~n34054 & ~n34087;
  assign n34089 = n3492 & ~n34088;
  assign n34090 = ~n3493 & ~n34089;
  assign n34091 = n3485 & ~n34090;
  assign n34092 = ~n3486 & ~n34091;
  assign n34093 = ~n3476 & ~n34092;
  assign n34094 = ~n3426 & ~n34022;
  assign n34095 = ~controllable_hmaster1 & ~n34094;
  assign n34096 = ~n3425 & ~n34095;
  assign n34097 = i_hbusreq3 & ~n34096;
  assign n34098 = ~n3455 & ~n34040;
  assign n34099 = ~controllable_hmaster1 & ~n34098;
  assign n34100 = ~n3454 & ~n34099;
  assign n34101 = ~i_hbusreq3 & ~n34100;
  assign n34102 = ~n34097 & ~n34101;
  assign n34103 = controllable_hmaster2 & ~n34102;
  assign n34104 = controllable_hmaster2 & ~n34103;
  assign n34105 = ~controllable_hgrant3 & ~n34104;
  assign n34106 = ~n3795 & ~n34105;
  assign n34107 = controllable_nhgrant0 & ~n34106;
  assign n34108 = ~n3810 & ~n34107;
  assign n34109 = ~n3281 & ~n34108;
  assign n34110 = ~n3783 & ~n34109;
  assign n34111 = ~n3378 & ~n34110;
  assign n34112 = ~n34054 & ~n34111;
  assign n34113 = ~n3485 & ~n34112;
  assign n34114 = ~n3492 & ~n34112;
  assign n34115 = ~n34089 & ~n34114;
  assign n34116 = n3485 & ~n34115;
  assign n34117 = ~n34113 & ~n34116;
  assign n34118 = n3476 & ~n34117;
  assign n34119 = ~n34093 & ~n34118;
  assign n34120 = ~n3374 & ~n34119;
  assign n34121 = controllable_hgrant4 & ~n5040;
  assign n34122 = ~n3850 & ~n34121;
  assign n34123 = ~controllable_hgrant2 & ~n34122;
  assign n34124 = ~n3410 & ~n34123;
  assign n34125 = ~controllable_hmaster0 & ~n34124;
  assign n34126 = ~controllable_hmaster0 & ~n34125;
  assign n34127 = ~controllable_hmaster1 & ~n34126;
  assign n34128 = ~controllable_hmaster1 & ~n34127;
  assign n34129 = i_hbusreq3 & ~n34128;
  assign n34130 = i_hbusreq2 & ~n34122;
  assign n34131 = controllable_hgrant4 & ~n5063;
  assign n34132 = ~n3884 & ~n34131;
  assign n34133 = ~i_hbusreq2 & ~n34132;
  assign n34134 = ~n34130 & ~n34133;
  assign n34135 = ~controllable_hgrant2 & ~n34134;
  assign n34136 = ~n3859 & ~n34135;
  assign n34137 = ~controllable_hmaster0 & ~n34136;
  assign n34138 = ~controllable_hmaster0 & ~n34137;
  assign n34139 = ~controllable_hmaster1 & ~n34138;
  assign n34140 = ~controllable_hmaster1 & ~n34139;
  assign n34141 = ~i_hbusreq3 & ~n34140;
  assign n34142 = ~n34129 & ~n34141;
  assign n34143 = controllable_hmaster2 & ~n34142;
  assign n34144 = controllable_hmaster2 & ~n34143;
  assign n34145 = ~controllable_hgrant3 & ~n34144;
  assign n34146 = ~n3843 & ~n34145;
  assign n34147 = controllable_nhgrant0 & ~n34146;
  assign n34148 = ~n3945 & ~n34147;
  assign n34149 = ~n3281 & ~n34148;
  assign n34150 = ~n3281 & ~n34149;
  assign n34151 = n3378 & ~n34150;
  assign n34152 = ~n3497 & ~n34055;
  assign n34153 = ~controllable_hgrant2 & ~n34152;
  assign n34154 = ~n3410 & ~n34153;
  assign n34155 = controllable_hmaster1 & ~n34154;
  assign n34156 = controllable_hmaster0 & ~n34154;
  assign n34157 = ~n34125 & ~n34156;
  assign n34158 = ~controllable_hmaster1 & ~n34157;
  assign n34159 = ~n34155 & ~n34158;
  assign n34160 = i_hbusreq3 & ~n34159;
  assign n34161 = i_hbusreq2 & ~n34152;
  assign n34162 = ~n3517 & ~n34066;
  assign n34163 = ~i_hbusreq2 & ~n34162;
  assign n34164 = ~n34161 & ~n34163;
  assign n34165 = ~controllable_hgrant2 & ~n34164;
  assign n34166 = ~n3431 & ~n34165;
  assign n34167 = controllable_hmaster1 & ~n34166;
  assign n34168 = controllable_hmaster0 & ~n34166;
  assign n34169 = ~n34137 & ~n34168;
  assign n34170 = ~controllable_hmaster1 & ~n34169;
  assign n34171 = ~n34167 & ~n34170;
  assign n34172 = ~i_hbusreq3 & ~n34171;
  assign n34173 = ~n34160 & ~n34172;
  assign n34174 = controllable_hmaster2 & ~n34173;
  assign n34175 = controllable_hmaster2 & ~n34174;
  assign n34176 = ~controllable_hgrant3 & ~n34175;
  assign n34177 = ~n3959 & ~n34176;
  assign n34178 = controllable_nhgrant0 & ~n34177;
  assign n34179 = ~n3987 & ~n34178;
  assign n34180 = ~n3281 & ~n34179;
  assign n34181 = ~n3950 & ~n34180;
  assign n34182 = ~n3378 & ~n34181;
  assign n34183 = ~n34151 & ~n34182;
  assign n34184 = n3492 & ~n34183;
  assign n34185 = ~n3493 & ~n34184;
  assign n34186 = n3485 & ~n34185;
  assign n34187 = ~n3486 & ~n34186;
  assign n34188 = ~n3476 & ~n34187;
  assign n34189 = controllable_hgrant4 & ~n14485;
  assign n34190 = controllable_hgrant4 & ~n34189;
  assign n34191 = ~controllable_hgrant2 & ~n34190;
  assign n34192 = ~controllable_hgrant2 & ~n34191;
  assign n34193 = controllable_hmaster1 & ~n34192;
  assign n34194 = controllable_hmaster0 & ~n34192;
  assign n34195 = controllable_hgrant4 & ~n6039;
  assign n34196 = ~n3850 & ~n34195;
  assign n34197 = ~controllable_hgrant2 & ~n34196;
  assign n34198 = ~n3410 & ~n34197;
  assign n34199 = ~controllable_hmaster0 & ~n34198;
  assign n34200 = ~n34194 & ~n34199;
  assign n34201 = ~controllable_hmaster1 & ~n34200;
  assign n34202 = ~n34193 & ~n34201;
  assign n34203 = i_hbusreq3 & ~n34202;
  assign n34204 = i_hbusreq2 & ~n34190;
  assign n34205 = controllable_hgrant4 & ~n14501;
  assign n34206 = controllable_hgrant4 & ~n34205;
  assign n34207 = ~i_hbusreq2 & ~n34206;
  assign n34208 = ~n34204 & ~n34207;
  assign n34209 = ~controllable_hgrant2 & ~n34208;
  assign n34210 = ~controllable_hgrant2 & ~n34209;
  assign n34211 = controllable_hmaster1 & ~n34210;
  assign n34212 = controllable_hmaster0 & ~n34210;
  assign n34213 = i_hbusreq2 & ~n34196;
  assign n34214 = controllable_hgrant4 & ~n6808;
  assign n34215 = ~n3884 & ~n34214;
  assign n34216 = ~i_hbusreq2 & ~n34215;
  assign n34217 = ~n34213 & ~n34216;
  assign n34218 = ~controllable_hgrant2 & ~n34217;
  assign n34219 = ~n3859 & ~n34218;
  assign n34220 = ~controllable_hmaster0 & ~n34219;
  assign n34221 = ~n34212 & ~n34220;
  assign n34222 = ~controllable_hmaster1 & ~n34221;
  assign n34223 = ~n34211 & ~n34222;
  assign n34224 = ~i_hbusreq3 & ~n34223;
  assign n34225 = ~n34203 & ~n34224;
  assign n34226 = controllable_hmaster2 & ~n34225;
  assign n34227 = i_hbusreq3 & ~n34192;
  assign n34228 = ~i_hbusreq3 & ~n34210;
  assign n34229 = ~n34227 & ~n34228;
  assign n34230 = ~controllable_hmaster2 & ~n34229;
  assign n34231 = ~n34226 & ~n34230;
  assign n34232 = ~controllable_hgrant3 & ~n34231;
  assign n34233 = ~n3843 & ~n34232;
  assign n34234 = controllable_nhgrant0 & ~n34233;
  assign n34235 = ~n3945 & ~n34234;
  assign n34236 = ~n3281 & ~n34235;
  assign n34237 = ~n3281 & ~n34236;
  assign n34238 = n3378 & ~n34237;
  assign n34239 = controllable_hgrant4 & ~n9055;
  assign n34240 = ~n3545 & ~n34239;
  assign n34241 = ~controllable_hgrant2 & ~n34240;
  assign n34242 = ~n3410 & ~n34241;
  assign n34243 = controllable_hmaster1 & ~n34242;
  assign n34244 = controllable_hmaster0 & ~n34242;
  assign n34245 = ~n3545 & ~n34195;
  assign n34246 = ~controllable_hgrant2 & ~n34245;
  assign n34247 = ~n3410 & ~n34246;
  assign n34248 = ~controllable_hmaster0 & ~n34247;
  assign n34249 = ~n34244 & ~n34248;
  assign n34250 = ~controllable_hmaster1 & ~n34249;
  assign n34251 = ~n34243 & ~n34250;
  assign n34252 = i_hbusreq3 & ~n34251;
  assign n34253 = i_hbusreq2 & ~n34240;
  assign n34254 = controllable_hgrant4 & ~n14554;
  assign n34255 = ~n3574 & ~n34254;
  assign n34256 = ~i_hbusreq2 & ~n34255;
  assign n34257 = ~n34253 & ~n34256;
  assign n34258 = ~controllable_hgrant2 & ~n34257;
  assign n34259 = ~n3431 & ~n34258;
  assign n34260 = controllable_hmaster1 & ~n34259;
  assign n34261 = controllable_hmaster0 & ~n34259;
  assign n34262 = i_hbusreq2 & ~n34245;
  assign n34263 = ~n4134 & ~n34214;
  assign n34264 = ~i_hbusreq2 & ~n34263;
  assign n34265 = ~n34262 & ~n34264;
  assign n34266 = ~controllable_hgrant2 & ~n34265;
  assign n34267 = ~n3859 & ~n34266;
  assign n34268 = ~controllable_hmaster0 & ~n34267;
  assign n34269 = ~n34261 & ~n34268;
  assign n34270 = ~controllable_hmaster1 & ~n34269;
  assign n34271 = ~n34260 & ~n34270;
  assign n34272 = ~i_hbusreq3 & ~n34271;
  assign n34273 = ~n34252 & ~n34272;
  assign n34274 = controllable_hmaster2 & ~n34273;
  assign n34275 = ~n3552 & ~n34189;
  assign n34276 = ~controllable_hgrant2 & ~n34275;
  assign n34277 = ~controllable_hgrant2 & ~n34276;
  assign n34278 = i_hbusreq3 & ~n34277;
  assign n34279 = i_hbusreq2 & ~n34275;
  assign n34280 = ~n3590 & ~n34205;
  assign n34281 = ~i_hbusreq2 & ~n34280;
  assign n34282 = ~n34279 & ~n34281;
  assign n34283 = ~controllable_hgrant2 & ~n34282;
  assign n34284 = ~controllable_hgrant2 & ~n34283;
  assign n34285 = ~i_hbusreq3 & ~n34284;
  assign n34286 = ~n34278 & ~n34285;
  assign n34287 = ~controllable_hmaster2 & ~n34286;
  assign n34288 = ~n34274 & ~n34287;
  assign n34289 = ~controllable_hgrant3 & ~n34288;
  assign n34290 = ~n3959 & ~n34289;
  assign n34291 = controllable_nhgrant0 & ~n34290;
  assign n34292 = ~n3987 & ~n34291;
  assign n34293 = ~n3281 & ~n34292;
  assign n34294 = ~n4089 & ~n34293;
  assign n34295 = ~n3378 & ~n34294;
  assign n34296 = ~n34238 & ~n34295;
  assign n34297 = n3492 & ~n34296;
  assign n34298 = ~n34114 & ~n34297;
  assign n34299 = n3485 & ~n34298;
  assign n34300 = ~n34113 & ~n34299;
  assign n34301 = n3476 & ~n34300;
  assign n34302 = ~n34188 & ~n34301;
  assign n34303 = n3374 & ~n34302;
  assign n34304 = ~n34120 & ~n34303;
  assign n34305 = n3655 & ~n34304;
  assign n34306 = ~n4182 & ~n34121;
  assign n34307 = ~controllable_hgrant2 & ~n34306;
  assign n34308 = ~n3410 & ~n34307;
  assign n34309 = ~controllable_hmaster0 & ~n34308;
  assign n34310 = ~controllable_hmaster0 & ~n34309;
  assign n34311 = ~controllable_hmaster1 & ~n34310;
  assign n34312 = ~controllable_hmaster1 & ~n34311;
  assign n34313 = i_hbusreq3 & ~n34312;
  assign n34314 = i_hbusreq2 & ~n34306;
  assign n34315 = ~n4204 & ~n34131;
  assign n34316 = ~i_hbusreq2 & ~n34315;
  assign n34317 = ~n34314 & ~n34316;
  assign n34318 = ~controllable_hgrant2 & ~n34317;
  assign n34319 = ~n3859 & ~n34318;
  assign n34320 = ~controllable_hmaster0 & ~n34319;
  assign n34321 = ~controllable_hmaster0 & ~n34320;
  assign n34322 = ~controllable_hmaster1 & ~n34321;
  assign n34323 = ~controllable_hmaster1 & ~n34322;
  assign n34324 = ~i_hbusreq3 & ~n34323;
  assign n34325 = ~n34313 & ~n34324;
  assign n34326 = controllable_hmaster2 & ~n34325;
  assign n34327 = controllable_hmaster2 & ~n34326;
  assign n34328 = ~controllable_hgrant3 & ~n34327;
  assign n34329 = ~n3843 & ~n34328;
  assign n34330 = controllable_nhgrant0 & ~n34329;
  assign n34331 = ~n3945 & ~n34330;
  assign n34332 = ~n3281 & ~n34331;
  assign n34333 = ~n3281 & ~n34332;
  assign n34334 = n3378 & ~n34333;
  assign n34335 = ~n34156 & ~n34309;
  assign n34336 = ~controllable_hmaster1 & ~n34335;
  assign n34337 = ~n34155 & ~n34336;
  assign n34338 = i_hbusreq3 & ~n34337;
  assign n34339 = ~n34168 & ~n34320;
  assign n34340 = ~controllable_hmaster1 & ~n34339;
  assign n34341 = ~n34167 & ~n34340;
  assign n34342 = ~i_hbusreq3 & ~n34341;
  assign n34343 = ~n34338 & ~n34342;
  assign n34344 = controllable_hmaster2 & ~n34343;
  assign n34345 = controllable_hmaster2 & ~n34344;
  assign n34346 = ~controllable_hgrant3 & ~n34345;
  assign n34347 = ~n3959 & ~n34346;
  assign n34348 = controllable_nhgrant0 & ~n34347;
  assign n34349 = ~n3987 & ~n34348;
  assign n34350 = ~n3281 & ~n34349;
  assign n34351 = ~n3950 & ~n34350;
  assign n34352 = ~n3378 & ~n34351;
  assign n34353 = ~n34334 & ~n34352;
  assign n34354 = n3492 & ~n34353;
  assign n34355 = ~n3493 & ~n34354;
  assign n34356 = n3485 & ~n34355;
  assign n34357 = ~n3486 & ~n34356;
  assign n34358 = ~n3476 & ~n34357;
  assign n34359 = ~n4182 & ~n34195;
  assign n34360 = ~controllable_hgrant2 & ~n34359;
  assign n34361 = ~n3410 & ~n34360;
  assign n34362 = ~controllable_hmaster0 & ~n34361;
  assign n34363 = ~n34194 & ~n34362;
  assign n34364 = ~controllable_hmaster1 & ~n34363;
  assign n34365 = ~n34193 & ~n34364;
  assign n34366 = i_hbusreq3 & ~n34365;
  assign n34367 = i_hbusreq2 & ~n34359;
  assign n34368 = ~n4204 & ~n34214;
  assign n34369 = ~i_hbusreq2 & ~n34368;
  assign n34370 = ~n34367 & ~n34369;
  assign n34371 = ~controllable_hgrant2 & ~n34370;
  assign n34372 = ~n3859 & ~n34371;
  assign n34373 = ~controllable_hmaster0 & ~n34372;
  assign n34374 = ~n34212 & ~n34373;
  assign n34375 = ~controllable_hmaster1 & ~n34374;
  assign n34376 = ~n34211 & ~n34375;
  assign n34377 = ~i_hbusreq3 & ~n34376;
  assign n34378 = ~n34366 & ~n34377;
  assign n34379 = controllable_hmaster2 & ~n34378;
  assign n34380 = ~n34230 & ~n34379;
  assign n34381 = ~controllable_hgrant3 & ~n34380;
  assign n34382 = ~n3843 & ~n34381;
  assign n34383 = controllable_nhgrant0 & ~n34382;
  assign n34384 = ~n3945 & ~n34383;
  assign n34385 = ~n3281 & ~n34384;
  assign n34386 = ~n3281 & ~n34385;
  assign n34387 = n3378 & ~n34386;
  assign n34388 = ~n4279 & ~n34195;
  assign n34389 = ~controllable_hgrant2 & ~n34388;
  assign n34390 = ~n3410 & ~n34389;
  assign n34391 = ~controllable_hmaster0 & ~n34390;
  assign n34392 = ~n34244 & ~n34391;
  assign n34393 = ~controllable_hmaster1 & ~n34392;
  assign n34394 = ~n34243 & ~n34393;
  assign n34395 = i_hbusreq3 & ~n34394;
  assign n34396 = i_hbusreq2 & ~n34388;
  assign n34397 = ~n4300 & ~n34214;
  assign n34398 = ~i_hbusreq2 & ~n34397;
  assign n34399 = ~n34396 & ~n34398;
  assign n34400 = ~controllable_hgrant2 & ~n34399;
  assign n34401 = ~n3859 & ~n34400;
  assign n34402 = ~controllable_hmaster0 & ~n34401;
  assign n34403 = ~n34261 & ~n34402;
  assign n34404 = ~controllable_hmaster1 & ~n34403;
  assign n34405 = ~n34260 & ~n34404;
  assign n34406 = ~i_hbusreq3 & ~n34405;
  assign n34407 = ~n34395 & ~n34406;
  assign n34408 = controllable_hmaster2 & ~n34407;
  assign n34409 = ~n34287 & ~n34408;
  assign n34410 = ~controllable_hgrant3 & ~n34409;
  assign n34411 = ~n3959 & ~n34410;
  assign n34412 = controllable_nhgrant0 & ~n34411;
  assign n34413 = ~n3987 & ~n34412;
  assign n34414 = ~n3281 & ~n34413;
  assign n34415 = ~n4089 & ~n34414;
  assign n34416 = ~n3378 & ~n34415;
  assign n34417 = ~n34387 & ~n34416;
  assign n34418 = n3492 & ~n34417;
  assign n34419 = ~n34114 & ~n34418;
  assign n34420 = n3485 & ~n34419;
  assign n34421 = ~n34113 & ~n34420;
  assign n34422 = n3476 & ~n34421;
  assign n34423 = ~n34358 & ~n34422;
  assign n34424 = n3374 & ~n34423;
  assign n34425 = ~n34120 & ~n34424;
  assign n34426 = ~n3655 & ~n34425;
  assign n34427 = ~n34305 & ~n34426;
  assign n34428 = n3652 & ~n34427;
  assign n34429 = ~n4333 & ~n34123;
  assign n34430 = ~controllable_hmaster0 & ~n34429;
  assign n34431 = ~controllable_hmaster0 & ~n34430;
  assign n34432 = ~controllable_hmaster1 & ~n34431;
  assign n34433 = ~controllable_hmaster1 & ~n34432;
  assign n34434 = i_hbusreq3 & ~n34433;
  assign n34435 = ~n4340 & ~n34135;
  assign n34436 = ~controllable_hmaster0 & ~n34435;
  assign n34437 = ~controllable_hmaster0 & ~n34436;
  assign n34438 = ~controllable_hmaster1 & ~n34437;
  assign n34439 = ~controllable_hmaster1 & ~n34438;
  assign n34440 = ~i_hbusreq3 & ~n34439;
  assign n34441 = ~n34434 & ~n34440;
  assign n34442 = controllable_hmaster2 & ~n34441;
  assign n34443 = controllable_hmaster2 & ~n34442;
  assign n34444 = ~controllable_hgrant3 & ~n34443;
  assign n34445 = ~n3843 & ~n34444;
  assign n34446 = controllable_nhgrant0 & ~n34445;
  assign n34447 = ~n3945 & ~n34446;
  assign n34448 = ~n3281 & ~n34447;
  assign n34449 = ~n3281 & ~n34448;
  assign n34450 = n3378 & ~n34449;
  assign n34451 = ~n34156 & ~n34430;
  assign n34452 = ~controllable_hmaster1 & ~n34451;
  assign n34453 = ~n34155 & ~n34452;
  assign n34454 = i_hbusreq3 & ~n34453;
  assign n34455 = ~n34168 & ~n34436;
  assign n34456 = ~controllable_hmaster1 & ~n34455;
  assign n34457 = ~n34167 & ~n34456;
  assign n34458 = ~i_hbusreq3 & ~n34457;
  assign n34459 = ~n34454 & ~n34458;
  assign n34460 = controllable_hmaster2 & ~n34459;
  assign n34461 = controllable_hmaster2 & ~n34460;
  assign n34462 = ~controllable_hgrant3 & ~n34461;
  assign n34463 = ~n3959 & ~n34462;
  assign n34464 = controllable_nhgrant0 & ~n34463;
  assign n34465 = ~n3987 & ~n34464;
  assign n34466 = ~n3281 & ~n34465;
  assign n34467 = ~n3950 & ~n34466;
  assign n34468 = ~n3378 & ~n34467;
  assign n34469 = ~n34450 & ~n34468;
  assign n34470 = n3492 & ~n34469;
  assign n34471 = ~n3493 & ~n34470;
  assign n34472 = n3485 & ~n34471;
  assign n34473 = ~n3486 & ~n34472;
  assign n34474 = ~n3476 & ~n34473;
  assign n34475 = ~n4333 & ~n34197;
  assign n34476 = ~controllable_hmaster0 & ~n34475;
  assign n34477 = ~n34194 & ~n34476;
  assign n34478 = ~controllable_hmaster1 & ~n34477;
  assign n34479 = ~n34193 & ~n34478;
  assign n34480 = i_hbusreq3 & ~n34479;
  assign n34481 = ~n4340 & ~n34218;
  assign n34482 = ~controllable_hmaster0 & ~n34481;
  assign n34483 = ~n34212 & ~n34482;
  assign n34484 = ~controllable_hmaster1 & ~n34483;
  assign n34485 = ~n34211 & ~n34484;
  assign n34486 = ~i_hbusreq3 & ~n34485;
  assign n34487 = ~n34480 & ~n34486;
  assign n34488 = controllable_hmaster2 & ~n34487;
  assign n34489 = ~n34230 & ~n34488;
  assign n34490 = ~controllable_hgrant3 & ~n34489;
  assign n34491 = ~n3843 & ~n34490;
  assign n34492 = controllable_nhgrant0 & ~n34491;
  assign n34493 = ~n3945 & ~n34492;
  assign n34494 = ~n3281 & ~n34493;
  assign n34495 = ~n3281 & ~n34494;
  assign n34496 = n3378 & ~n34495;
  assign n34497 = ~n4333 & ~n34246;
  assign n34498 = ~controllable_hmaster0 & ~n34497;
  assign n34499 = ~n34244 & ~n34498;
  assign n34500 = ~controllable_hmaster1 & ~n34499;
  assign n34501 = ~n34243 & ~n34500;
  assign n34502 = i_hbusreq3 & ~n34501;
  assign n34503 = ~n4340 & ~n34266;
  assign n34504 = ~controllable_hmaster0 & ~n34503;
  assign n34505 = ~n34261 & ~n34504;
  assign n34506 = ~controllable_hmaster1 & ~n34505;
  assign n34507 = ~n34260 & ~n34506;
  assign n34508 = ~i_hbusreq3 & ~n34507;
  assign n34509 = ~n34502 & ~n34508;
  assign n34510 = controllable_hmaster2 & ~n34509;
  assign n34511 = ~n34287 & ~n34510;
  assign n34512 = ~controllable_hgrant3 & ~n34511;
  assign n34513 = ~n3959 & ~n34512;
  assign n34514 = controllable_nhgrant0 & ~n34513;
  assign n34515 = ~n3987 & ~n34514;
  assign n34516 = ~n3281 & ~n34515;
  assign n34517 = ~n4089 & ~n34516;
  assign n34518 = ~n3378 & ~n34517;
  assign n34519 = ~n34496 & ~n34518;
  assign n34520 = n3492 & ~n34519;
  assign n34521 = ~n34114 & ~n34520;
  assign n34522 = n3485 & ~n34521;
  assign n34523 = ~n34113 & ~n34522;
  assign n34524 = n3476 & ~n34523;
  assign n34525 = ~n34474 & ~n34524;
  assign n34526 = n3374 & ~n34525;
  assign n34527 = ~n34120 & ~n34526;
  assign n34528 = n3655 & ~n34527;
  assign n34529 = ~n4333 & ~n34307;
  assign n34530 = ~controllable_hmaster0 & ~n34529;
  assign n34531 = ~controllable_hmaster0 & ~n34530;
  assign n34532 = ~controllable_hmaster1 & ~n34531;
  assign n34533 = ~controllable_hmaster1 & ~n34532;
  assign n34534 = i_hbusreq3 & ~n34533;
  assign n34535 = ~n4340 & ~n34318;
  assign n34536 = ~controllable_hmaster0 & ~n34535;
  assign n34537 = ~controllable_hmaster0 & ~n34536;
  assign n34538 = ~controllable_hmaster1 & ~n34537;
  assign n34539 = ~controllable_hmaster1 & ~n34538;
  assign n34540 = ~i_hbusreq3 & ~n34539;
  assign n34541 = ~n34534 & ~n34540;
  assign n34542 = controllable_hmaster2 & ~n34541;
  assign n34543 = controllable_hmaster2 & ~n34542;
  assign n34544 = ~controllable_hgrant3 & ~n34543;
  assign n34545 = ~n3843 & ~n34544;
  assign n34546 = controllable_nhgrant0 & ~n34545;
  assign n34547 = ~n3945 & ~n34546;
  assign n34548 = ~n3281 & ~n34547;
  assign n34549 = ~n3281 & ~n34548;
  assign n34550 = n3378 & ~n34549;
  assign n34551 = ~n34156 & ~n34530;
  assign n34552 = ~controllable_hmaster1 & ~n34551;
  assign n34553 = ~n34155 & ~n34552;
  assign n34554 = i_hbusreq3 & ~n34553;
  assign n34555 = ~n34168 & ~n34536;
  assign n34556 = ~controllable_hmaster1 & ~n34555;
  assign n34557 = ~n34167 & ~n34556;
  assign n34558 = ~i_hbusreq3 & ~n34557;
  assign n34559 = ~n34554 & ~n34558;
  assign n34560 = controllable_hmaster2 & ~n34559;
  assign n34561 = controllable_hmaster2 & ~n34560;
  assign n34562 = ~controllable_hgrant3 & ~n34561;
  assign n34563 = ~n3959 & ~n34562;
  assign n34564 = controllable_nhgrant0 & ~n34563;
  assign n34565 = ~n3987 & ~n34564;
  assign n34566 = ~n3281 & ~n34565;
  assign n34567 = ~n3950 & ~n34566;
  assign n34568 = ~n3378 & ~n34567;
  assign n34569 = ~n34550 & ~n34568;
  assign n34570 = n3492 & ~n34569;
  assign n34571 = ~n3493 & ~n34570;
  assign n34572 = n3485 & ~n34571;
  assign n34573 = ~n3486 & ~n34572;
  assign n34574 = ~n3476 & ~n34573;
  assign n34575 = ~n4333 & ~n34360;
  assign n34576 = ~controllable_hmaster0 & ~n34575;
  assign n34577 = ~n34194 & ~n34576;
  assign n34578 = ~controllable_hmaster1 & ~n34577;
  assign n34579 = ~n34193 & ~n34578;
  assign n34580 = i_hbusreq3 & ~n34579;
  assign n34581 = ~n4340 & ~n34371;
  assign n34582 = ~controllable_hmaster0 & ~n34581;
  assign n34583 = ~n34212 & ~n34582;
  assign n34584 = ~controllable_hmaster1 & ~n34583;
  assign n34585 = ~n34211 & ~n34584;
  assign n34586 = ~i_hbusreq3 & ~n34585;
  assign n34587 = ~n34580 & ~n34586;
  assign n34588 = controllable_hmaster2 & ~n34587;
  assign n34589 = ~n34230 & ~n34588;
  assign n34590 = ~controllable_hgrant3 & ~n34589;
  assign n34591 = ~n3843 & ~n34590;
  assign n34592 = controllable_nhgrant0 & ~n34591;
  assign n34593 = ~n3945 & ~n34592;
  assign n34594 = ~n3281 & ~n34593;
  assign n34595 = ~n3281 & ~n34594;
  assign n34596 = n3378 & ~n34595;
  assign n34597 = ~n4333 & ~n34389;
  assign n34598 = ~controllable_hmaster0 & ~n34597;
  assign n34599 = ~n34244 & ~n34598;
  assign n34600 = ~controllable_hmaster1 & ~n34599;
  assign n34601 = ~n34243 & ~n34600;
  assign n34602 = i_hbusreq3 & ~n34601;
  assign n34603 = ~n4340 & ~n34400;
  assign n34604 = ~controllable_hmaster0 & ~n34603;
  assign n34605 = ~n34261 & ~n34604;
  assign n34606 = ~controllable_hmaster1 & ~n34605;
  assign n34607 = ~n34260 & ~n34606;
  assign n34608 = ~i_hbusreq3 & ~n34607;
  assign n34609 = ~n34602 & ~n34608;
  assign n34610 = controllable_hmaster2 & ~n34609;
  assign n34611 = ~n34287 & ~n34610;
  assign n34612 = ~controllable_hgrant3 & ~n34611;
  assign n34613 = ~n3959 & ~n34612;
  assign n34614 = controllable_nhgrant0 & ~n34613;
  assign n34615 = ~n3987 & ~n34614;
  assign n34616 = ~n3281 & ~n34615;
  assign n34617 = ~n4089 & ~n34616;
  assign n34618 = ~n3378 & ~n34617;
  assign n34619 = ~n34596 & ~n34618;
  assign n34620 = n3492 & ~n34619;
  assign n34621 = ~n34114 & ~n34620;
  assign n34622 = n3485 & ~n34621;
  assign n34623 = ~n34113 & ~n34622;
  assign n34624 = n3476 & ~n34623;
  assign n34625 = ~n34574 & ~n34624;
  assign n34626 = n3374 & ~n34625;
  assign n34627 = ~n34120 & ~n34626;
  assign n34628 = ~n3655 & ~n34627;
  assign n34629 = ~n34528 & ~n34628;
  assign n34630 = ~n3652 & ~n34629;
  assign n34631 = ~n34428 & ~n34630;
  assign n34632 = ~n3368 & ~n34631;
  assign n34633 = controllable_hgrant4 & ~n3496;
  assign n34634 = ~n3850 & ~n34633;
  assign n34635 = ~controllable_hgrant2 & ~n34634;
  assign n34636 = ~n3410 & ~n34635;
  assign n34637 = ~controllable_hmaster0 & ~n34636;
  assign n34638 = ~controllable_hmaster0 & ~n34637;
  assign n34639 = ~controllable_hmaster1 & ~n34638;
  assign n34640 = ~controllable_hmaster1 & ~n34639;
  assign n34641 = i_hbusreq3 & ~n34640;
  assign n34642 = i_hbusreq2 & ~n34634;
  assign n34643 = controllable_hgrant4 & ~n9717;
  assign n34644 = ~n4585 & ~n34643;
  assign n34645 = ~i_hbusreq2 & ~n34644;
  assign n34646 = ~n34642 & ~n34645;
  assign n34647 = ~controllable_hgrant2 & ~n34646;
  assign n34648 = ~n4562 & ~n34647;
  assign n34649 = ~controllable_hmaster0 & ~n34648;
  assign n34650 = ~controllable_hmaster0 & ~n34649;
  assign n34651 = ~controllable_hmaster1 & ~n34650;
  assign n34652 = ~controllable_hmaster1 & ~n34651;
  assign n34653 = ~i_hbusreq3 & ~n34652;
  assign n34654 = ~n34641 & ~n34653;
  assign n34655 = controllable_hmaster2 & ~n34654;
  assign n34656 = controllable_hmaster2 & ~n34655;
  assign n34657 = ~controllable_hgrant3 & ~n34656;
  assign n34658 = ~n4561 & ~n34657;
  assign n34659 = controllable_nhgrant0 & ~n34658;
  assign n34660 = ~n4646 & ~n34659;
  assign n34661 = ~n3281 & ~n34660;
  assign n34662 = ~n3281 & ~n34661;
  assign n34663 = n3492 & ~n34662;
  assign n34664 = n3492 & ~n34663;
  assign n34665 = n3485 & ~n34664;
  assign n34666 = n3485 & ~n34665;
  assign n34667 = ~n3476 & ~n34666;
  assign n34668 = ~n3485 & ~n34053;
  assign n34669 = ~n3492 & ~n34053;
  assign n34670 = i_hlock4 & ~n3551;
  assign n34671 = ~i_hlock4 & ~n14838;
  assign n34672 = ~n34670 & ~n34671;
  assign n34673 = controllable_hgrant4 & ~n34672;
  assign n34674 = controllable_hgrant4 & ~n34673;
  assign n34675 = ~controllable_hgrant2 & ~n34674;
  assign n34676 = ~controllable_hgrant2 & ~n34675;
  assign n34677 = controllable_hmaster1 & ~n34676;
  assign n34678 = controllable_hmaster0 & ~n34676;
  assign n34679 = i_hlock4 & ~n3544;
  assign n34680 = ~i_hlock4 & ~n10217;
  assign n34681 = ~n34679 & ~n34680;
  assign n34682 = controllable_hgrant4 & ~n34681;
  assign n34683 = ~n3850 & ~n34682;
  assign n34684 = ~controllable_hgrant2 & ~n34683;
  assign n34685 = ~n3410 & ~n34684;
  assign n34686 = ~controllable_hmaster0 & ~n34685;
  assign n34687 = ~n34678 & ~n34686;
  assign n34688 = ~controllable_hmaster1 & ~n34687;
  assign n34689 = ~n34677 & ~n34688;
  assign n34690 = i_hbusreq3 & ~n34689;
  assign n34691 = i_hbusreq2 & ~n34674;
  assign n34692 = i_hbusreq4 & ~n34672;
  assign n34693 = i_hlock4 & ~n14849;
  assign n34694 = ~n34671 & ~n34693;
  assign n34695 = ~i_hbusreq4 & ~n34694;
  assign n34696 = ~n34692 & ~n34695;
  assign n34697 = controllable_hgrant4 & ~n34696;
  assign n34698 = controllable_hgrant4 & ~n34697;
  assign n34699 = ~i_hbusreq2 & ~n34698;
  assign n34700 = ~n34691 & ~n34699;
  assign n34701 = ~controllable_hgrant2 & ~n34700;
  assign n34702 = ~controllable_hgrant2 & ~n34701;
  assign n34703 = controllable_hmaster1 & ~n34702;
  assign n34704 = controllable_hmaster0 & ~n34702;
  assign n34705 = i_hbusreq2 & ~n34683;
  assign n34706 = i_hbusreq4 & ~n34681;
  assign n34707 = i_hlock4 & ~n11087;
  assign n34708 = ~i_hlock4 & ~n11101;
  assign n34709 = ~n34707 & ~n34708;
  assign n34710 = ~i_hbusreq4 & ~n34709;
  assign n34711 = ~n34706 & ~n34710;
  assign n34712 = controllable_hgrant4 & ~n34711;
  assign n34713 = ~n4585 & ~n34712;
  assign n34714 = ~i_hbusreq2 & ~n34713;
  assign n34715 = ~n34705 & ~n34714;
  assign n34716 = ~controllable_hgrant2 & ~n34715;
  assign n34717 = ~n4562 & ~n34716;
  assign n34718 = ~controllable_hmaster0 & ~n34717;
  assign n34719 = ~n34704 & ~n34718;
  assign n34720 = ~controllable_hmaster1 & ~n34719;
  assign n34721 = ~n34703 & ~n34720;
  assign n34722 = ~i_hbusreq3 & ~n34721;
  assign n34723 = ~n34690 & ~n34722;
  assign n34724 = controllable_hmaster2 & ~n34723;
  assign n34725 = i_hbusreq3 & ~n34676;
  assign n34726 = ~i_hbusreq3 & ~n34702;
  assign n34727 = ~n34725 & ~n34726;
  assign n34728 = ~controllable_hmaster2 & ~n34727;
  assign n34729 = ~n34724 & ~n34728;
  assign n34730 = ~controllable_hgrant3 & ~n34729;
  assign n34731 = ~n4561 & ~n34730;
  assign n34732 = controllable_nhgrant0 & ~n34731;
  assign n34733 = ~n4646 & ~n34732;
  assign n34734 = ~n3281 & ~n34733;
  assign n34735 = ~n3281 & ~n34734;
  assign n34736 = n3492 & ~n34735;
  assign n34737 = ~n34669 & ~n34736;
  assign n34738 = n3485 & ~n34737;
  assign n34739 = ~n34668 & ~n34738;
  assign n34740 = n3476 & ~n34739;
  assign n34741 = ~n34667 & ~n34740;
  assign n34742 = n3374 & ~n34741;
  assign n34743 = n3374 & ~n34742;
  assign n34744 = n3655 & ~n34743;
  assign n34745 = ~n4701 & ~n34633;
  assign n34746 = ~controllable_hgrant2 & ~n34745;
  assign n34747 = ~n3410 & ~n34746;
  assign n34748 = ~controllable_hmaster0 & ~n34747;
  assign n34749 = ~controllable_hmaster0 & ~n34748;
  assign n34750 = ~controllable_hmaster1 & ~n34749;
  assign n34751 = ~controllable_hmaster1 & ~n34750;
  assign n34752 = i_hbusreq3 & ~n34751;
  assign n34753 = i_hbusreq2 & ~n34745;
  assign n34754 = ~n4723 & ~n34643;
  assign n34755 = ~i_hbusreq2 & ~n34754;
  assign n34756 = ~n34753 & ~n34755;
  assign n34757 = ~controllable_hgrant2 & ~n34756;
  assign n34758 = ~n4562 & ~n34757;
  assign n34759 = ~controllable_hmaster0 & ~n34758;
  assign n34760 = ~controllable_hmaster0 & ~n34759;
  assign n34761 = ~controllable_hmaster1 & ~n34760;
  assign n34762 = ~controllable_hmaster1 & ~n34761;
  assign n34763 = ~i_hbusreq3 & ~n34762;
  assign n34764 = ~n34752 & ~n34763;
  assign n34765 = controllable_hmaster2 & ~n34764;
  assign n34766 = controllable_hmaster2 & ~n34765;
  assign n34767 = ~controllable_hgrant3 & ~n34766;
  assign n34768 = ~n4561 & ~n34767;
  assign n34769 = controllable_nhgrant0 & ~n34768;
  assign n34770 = ~n4646 & ~n34769;
  assign n34771 = ~n3281 & ~n34770;
  assign n34772 = ~n3281 & ~n34771;
  assign n34773 = n3492 & ~n34772;
  assign n34774 = n3492 & ~n34773;
  assign n34775 = n3485 & ~n34774;
  assign n34776 = n3485 & ~n34775;
  assign n34777 = ~n3476 & ~n34776;
  assign n34778 = ~n4701 & ~n34682;
  assign n34779 = ~controllable_hgrant2 & ~n34778;
  assign n34780 = ~n3410 & ~n34779;
  assign n34781 = ~controllable_hmaster0 & ~n34780;
  assign n34782 = ~n34678 & ~n34781;
  assign n34783 = ~controllable_hmaster1 & ~n34782;
  assign n34784 = ~n34677 & ~n34783;
  assign n34785 = i_hbusreq3 & ~n34784;
  assign n34786 = i_hbusreq2 & ~n34778;
  assign n34787 = ~n4723 & ~n34712;
  assign n34788 = ~i_hbusreq2 & ~n34787;
  assign n34789 = ~n34786 & ~n34788;
  assign n34790 = ~controllable_hgrant2 & ~n34789;
  assign n34791 = ~n4562 & ~n34790;
  assign n34792 = ~controllable_hmaster0 & ~n34791;
  assign n34793 = ~n34704 & ~n34792;
  assign n34794 = ~controllable_hmaster1 & ~n34793;
  assign n34795 = ~n34703 & ~n34794;
  assign n34796 = ~i_hbusreq3 & ~n34795;
  assign n34797 = ~n34785 & ~n34796;
  assign n34798 = controllable_hmaster2 & ~n34797;
  assign n34799 = ~n34728 & ~n34798;
  assign n34800 = ~controllable_hgrant3 & ~n34799;
  assign n34801 = ~n4561 & ~n34800;
  assign n34802 = controllable_nhgrant0 & ~n34801;
  assign n34803 = ~n4646 & ~n34802;
  assign n34804 = ~n3281 & ~n34803;
  assign n34805 = ~n3281 & ~n34804;
  assign n34806 = n3492 & ~n34805;
  assign n34807 = ~n34669 & ~n34806;
  assign n34808 = n3485 & ~n34807;
  assign n34809 = ~n34668 & ~n34808;
  assign n34810 = n3476 & ~n34809;
  assign n34811 = ~n34777 & ~n34810;
  assign n34812 = n3374 & ~n34811;
  assign n34813 = n3374 & ~n34812;
  assign n34814 = ~n3655 & ~n34813;
  assign n34815 = ~n34744 & ~n34814;
  assign n34816 = n3652 & ~n34815;
  assign n34817 = ~n4787 & ~n34635;
  assign n34818 = ~controllable_hmaster0 & ~n34817;
  assign n34819 = ~controllable_hmaster0 & ~n34818;
  assign n34820 = ~controllable_hmaster1 & ~n34819;
  assign n34821 = ~controllable_hmaster1 & ~n34820;
  assign n34822 = i_hbusreq3 & ~n34821;
  assign n34823 = ~n4794 & ~n34647;
  assign n34824 = ~controllable_hmaster0 & ~n34823;
  assign n34825 = ~controllable_hmaster0 & ~n34824;
  assign n34826 = ~controllable_hmaster1 & ~n34825;
  assign n34827 = ~controllable_hmaster1 & ~n34826;
  assign n34828 = ~i_hbusreq3 & ~n34827;
  assign n34829 = ~n34822 & ~n34828;
  assign n34830 = controllable_hmaster2 & ~n34829;
  assign n34831 = controllable_hmaster2 & ~n34830;
  assign n34832 = ~controllable_hgrant3 & ~n34831;
  assign n34833 = ~n4561 & ~n34832;
  assign n34834 = controllable_nhgrant0 & ~n34833;
  assign n34835 = ~n4646 & ~n34834;
  assign n34836 = ~n3281 & ~n34835;
  assign n34837 = ~n3281 & ~n34836;
  assign n34838 = n3492 & ~n34837;
  assign n34839 = n3492 & ~n34838;
  assign n34840 = n3485 & ~n34839;
  assign n34841 = n3485 & ~n34840;
  assign n34842 = ~n3476 & ~n34841;
  assign n34843 = ~n4787 & ~n34684;
  assign n34844 = ~controllable_hmaster0 & ~n34843;
  assign n34845 = ~n34678 & ~n34844;
  assign n34846 = ~controllable_hmaster1 & ~n34845;
  assign n34847 = ~n34677 & ~n34846;
  assign n34848 = i_hbusreq3 & ~n34847;
  assign n34849 = ~n4794 & ~n34716;
  assign n34850 = ~controllable_hmaster0 & ~n34849;
  assign n34851 = ~n34704 & ~n34850;
  assign n34852 = ~controllable_hmaster1 & ~n34851;
  assign n34853 = ~n34703 & ~n34852;
  assign n34854 = ~i_hbusreq3 & ~n34853;
  assign n34855 = ~n34848 & ~n34854;
  assign n34856 = controllable_hmaster2 & ~n34855;
  assign n34857 = ~n34728 & ~n34856;
  assign n34858 = ~controllable_hgrant3 & ~n34857;
  assign n34859 = ~n4561 & ~n34858;
  assign n34860 = controllable_nhgrant0 & ~n34859;
  assign n34861 = ~n4646 & ~n34860;
  assign n34862 = ~n3281 & ~n34861;
  assign n34863 = ~n3281 & ~n34862;
  assign n34864 = n3492 & ~n34863;
  assign n34865 = ~n34669 & ~n34864;
  assign n34866 = n3485 & ~n34865;
  assign n34867 = ~n34668 & ~n34866;
  assign n34868 = n3476 & ~n34867;
  assign n34869 = ~n34842 & ~n34868;
  assign n34870 = n3374 & ~n34869;
  assign n34871 = n3374 & ~n34870;
  assign n34872 = n3655 & ~n34871;
  assign n34873 = ~n4787 & ~n34746;
  assign n34874 = ~controllable_hmaster0 & ~n34873;
  assign n34875 = ~controllable_hmaster0 & ~n34874;
  assign n34876 = ~controllable_hmaster1 & ~n34875;
  assign n34877 = ~controllable_hmaster1 & ~n34876;
  assign n34878 = i_hbusreq3 & ~n34877;
  assign n34879 = ~n4794 & ~n34757;
  assign n34880 = ~controllable_hmaster0 & ~n34879;
  assign n34881 = ~controllable_hmaster0 & ~n34880;
  assign n34882 = ~controllable_hmaster1 & ~n34881;
  assign n34883 = ~controllable_hmaster1 & ~n34882;
  assign n34884 = ~i_hbusreq3 & ~n34883;
  assign n34885 = ~n34878 & ~n34884;
  assign n34886 = controllable_hmaster2 & ~n34885;
  assign n34887 = controllable_hmaster2 & ~n34886;
  assign n34888 = ~controllable_hgrant3 & ~n34887;
  assign n34889 = ~n4561 & ~n34888;
  assign n34890 = controllable_nhgrant0 & ~n34889;
  assign n34891 = ~n4646 & ~n34890;
  assign n34892 = ~n3281 & ~n34891;
  assign n34893 = ~n3281 & ~n34892;
  assign n34894 = n3492 & ~n34893;
  assign n34895 = n3492 & ~n34894;
  assign n34896 = n3485 & ~n34895;
  assign n34897 = n3485 & ~n34896;
  assign n34898 = ~n3476 & ~n34897;
  assign n34899 = ~n4787 & ~n34779;
  assign n34900 = ~controllable_hmaster0 & ~n34899;
  assign n34901 = ~n34678 & ~n34900;
  assign n34902 = ~controllable_hmaster1 & ~n34901;
  assign n34903 = ~n34677 & ~n34902;
  assign n34904 = i_hbusreq3 & ~n34903;
  assign n34905 = ~n4794 & ~n34790;
  assign n34906 = ~controllable_hmaster0 & ~n34905;
  assign n34907 = ~n34704 & ~n34906;
  assign n34908 = ~controllable_hmaster1 & ~n34907;
  assign n34909 = ~n34703 & ~n34908;
  assign n34910 = ~i_hbusreq3 & ~n34909;
  assign n34911 = ~n34904 & ~n34910;
  assign n34912 = controllable_hmaster2 & ~n34911;
  assign n34913 = ~n34728 & ~n34912;
  assign n34914 = ~controllable_hgrant3 & ~n34913;
  assign n34915 = ~n4561 & ~n34914;
  assign n34916 = controllable_nhgrant0 & ~n34915;
  assign n34917 = ~n4646 & ~n34916;
  assign n34918 = ~n3281 & ~n34917;
  assign n34919 = ~n3281 & ~n34918;
  assign n34920 = n3492 & ~n34919;
  assign n34921 = ~n34669 & ~n34920;
  assign n34922 = n3485 & ~n34921;
  assign n34923 = ~n34668 & ~n34922;
  assign n34924 = n3476 & ~n34923;
  assign n34925 = ~n34898 & ~n34924;
  assign n34926 = n3374 & ~n34925;
  assign n34927 = n3374 & ~n34926;
  assign n34928 = ~n3655 & ~n34927;
  assign n34929 = ~n34872 & ~n34928;
  assign n34930 = ~n3652 & ~n34929;
  assign n34931 = ~n34816 & ~n34930;
  assign n34932 = n3368 & ~n34931;
  assign n34933 = ~n34632 & ~n34932;
  assign n34934 = ~n3362 & ~n34933;
  assign n34935 = ~n3362 & ~n34934;
  assign n34936 = ~n3359 & ~n34935;
  assign n34937 = ~n3359 & ~n34936;
  assign n34938 = n3356 & ~n34937;
  assign n34939 = n3378 & ~n34086;
  assign n34940 = ~n5041 & ~n34055;
  assign n34941 = ~controllable_hgrant2 & ~n34940;
  assign n34942 = ~n3410 & ~n34941;
  assign n34943 = controllable_hmaster1 & ~n34942;
  assign n34944 = controllable_hmaster0 & ~n34942;
  assign n34945 = ~n34022 & ~n34944;
  assign n34946 = ~controllable_hmaster1 & ~n34945;
  assign n34947 = ~n34943 & ~n34946;
  assign n34948 = i_hbusreq3 & ~n34947;
  assign n34949 = i_hbusreq2 & ~n34940;
  assign n34950 = controllable_hgrant4 & ~n3883;
  assign n34951 = ~n5064 & ~n34950;
  assign n34952 = ~i_hbusreq2 & ~n34951;
  assign n34953 = ~n34949 & ~n34952;
  assign n34954 = ~controllable_hgrant2 & ~n34953;
  assign n34955 = ~n3859 & ~n34954;
  assign n34956 = controllable_hmaster1 & ~n34955;
  assign n34957 = controllable_hmaster0 & ~n34955;
  assign n34958 = ~n34040 & ~n34957;
  assign n34959 = ~controllable_hmaster1 & ~n34958;
  assign n34960 = ~n34956 & ~n34959;
  assign n34961 = ~i_hbusreq3 & ~n34960;
  assign n34962 = ~n34948 & ~n34961;
  assign n34963 = controllable_hmaster2 & ~n34962;
  assign n34964 = ~n5161 & ~n34963;
  assign n34965 = ~controllable_hgrant3 & ~n34964;
  assign n34966 = ~n5037 & ~n34965;
  assign n34967 = controllable_nhgrant0 & ~n34966;
  assign n34968 = ~n5245 & ~n34967;
  assign n34969 = ~n3281 & ~n34968;
  assign n34970 = ~n3783 & ~n34969;
  assign n34971 = ~n3378 & ~n34970;
  assign n34972 = ~n34939 & ~n34971;
  assign n34973 = n3492 & ~n34972;
  assign n34974 = ~n3631 & ~n34973;
  assign n34975 = n3485 & ~n34974;
  assign n34976 = ~n3630 & ~n34975;
  assign n34977 = ~n3476 & ~n34976;
  assign n34978 = ~n3485 & ~n34110;
  assign n34979 = ~n3492 & ~n34110;
  assign n34980 = ~n34973 & ~n34979;
  assign n34981 = n3485 & ~n34980;
  assign n34982 = ~n34978 & ~n34981;
  assign n34983 = n3476 & ~n34982;
  assign n34984 = ~n34977 & ~n34983;
  assign n34985 = ~n3374 & ~n34984;
  assign n34986 = controllable_hgrant4 & ~n3905;
  assign n34987 = ~n12042 & ~n34986;
  assign n34988 = ~controllable_hgrant2 & ~n34987;
  assign n34989 = ~n3410 & ~n34988;
  assign n34990 = controllable_hmaster0 & ~n34989;
  assign n34991 = ~n5288 & ~n34988;
  assign n34992 = ~controllable_hmaster0 & ~n34991;
  assign n34993 = ~n34990 & ~n34992;
  assign n34994 = controllable_hmaster1 & ~n34993;
  assign n34995 = ~n5299 & ~n34986;
  assign n34996 = ~controllable_hgrant2 & ~n34995;
  assign n34997 = ~n3410 & ~n34996;
  assign n34998 = controllable_hmaster0 & ~n34997;
  assign n34999 = ~controllable_hmaster0 & ~n34989;
  assign n35000 = ~n34998 & ~n34999;
  assign n35001 = ~controllable_hmaster1 & ~n35000;
  assign n35002 = ~n34994 & ~n35001;
  assign n35003 = i_hbusreq3 & ~n35002;
  assign n35004 = i_hbusreq2 & ~n34987;
  assign n35005 = controllable_hgrant4 & ~n15274;
  assign n35006 = ~n12053 & ~n35005;
  assign n35007 = ~i_hbusreq2 & ~n35006;
  assign n35008 = ~n35004 & ~n35007;
  assign n35009 = ~controllable_hgrant2 & ~n35008;
  assign n35010 = ~n3431 & ~n35009;
  assign n35011 = controllable_hmaster0 & ~n35010;
  assign n35012 = ~n5308 & ~n35009;
  assign n35013 = ~controllable_hmaster0 & ~n35012;
  assign n35014 = ~n35011 & ~n35013;
  assign n35015 = controllable_hmaster1 & ~n35014;
  assign n35016 = i_hbusreq2 & ~n34995;
  assign n35017 = ~n5326 & ~n35005;
  assign n35018 = ~i_hbusreq2 & ~n35017;
  assign n35019 = ~n35016 & ~n35018;
  assign n35020 = ~controllable_hgrant2 & ~n35019;
  assign n35021 = ~n3431 & ~n35020;
  assign n35022 = controllable_hmaster0 & ~n35021;
  assign n35023 = ~controllable_hmaster0 & ~n35010;
  assign n35024 = ~n35022 & ~n35023;
  assign n35025 = ~controllable_hmaster1 & ~n35024;
  assign n35026 = ~n35015 & ~n35025;
  assign n35027 = ~i_hbusreq3 & ~n35026;
  assign n35028 = ~n35003 & ~n35027;
  assign n35029 = ~controllable_hmaster2 & ~n35028;
  assign n35030 = ~n34174 & ~n35029;
  assign n35031 = ~controllable_hgrant3 & ~n35030;
  assign n35032 = ~n5287 & ~n35031;
  assign n35033 = controllable_nhgrant0 & ~n35032;
  assign n35034 = ~n5363 & ~n35033;
  assign n35035 = ~n3281 & ~n35034;
  assign n35036 = ~n3950 & ~n35035;
  assign n35037 = n3378 & ~n35036;
  assign n35038 = ~n5410 & ~n34950;
  assign n35039 = ~i_hbusreq2 & ~n35038;
  assign n35040 = ~n34161 & ~n35039;
  assign n35041 = ~controllable_hgrant2 & ~n35040;
  assign n35042 = ~n3859 & ~n35041;
  assign n35043 = controllable_hmaster1 & ~n35042;
  assign n35044 = controllable_hmaster0 & ~n35042;
  assign n35045 = ~n34137 & ~n35044;
  assign n35046 = ~controllable_hmaster1 & ~n35045;
  assign n35047 = ~n35043 & ~n35046;
  assign n35048 = ~i_hbusreq3 & ~n35047;
  assign n35049 = ~n34160 & ~n35048;
  assign n35050 = controllable_hmaster2 & ~n35049;
  assign n35051 = ~controllable_hgrant2 & ~n3905;
  assign n35052 = ~n3410 & ~n35051;
  assign n35053 = controllable_hmaster0 & ~n35052;
  assign n35054 = ~n5288 & ~n35051;
  assign n35055 = ~controllable_hmaster0 & ~n35054;
  assign n35056 = ~n35053 & ~n35055;
  assign n35057 = controllable_hmaster1 & ~n35056;
  assign n35058 = ~n5429 & ~n34986;
  assign n35059 = ~controllable_hgrant2 & ~n35058;
  assign n35060 = ~n3410 & ~n35059;
  assign n35061 = controllable_hmaster0 & ~n35060;
  assign n35062 = ~controllable_hmaster0 & ~n35052;
  assign n35063 = ~n35061 & ~n35062;
  assign n35064 = ~controllable_hmaster1 & ~n35063;
  assign n35065 = ~n35057 & ~n35064;
  assign n35066 = i_hbusreq3 & ~n35065;
  assign n35067 = i_hbusreq2 & ~n3905;
  assign n35068 = ~i_hbusreq2 & ~n3928;
  assign n35069 = ~n35067 & ~n35068;
  assign n35070 = ~controllable_hgrant2 & ~n35069;
  assign n35071 = ~n3859 & ~n35070;
  assign n35072 = controllable_hmaster0 & ~n35071;
  assign n35073 = ~n5438 & ~n35070;
  assign n35074 = ~controllable_hmaster0 & ~n35073;
  assign n35075 = ~n35072 & ~n35074;
  assign n35076 = controllable_hmaster1 & ~n35075;
  assign n35077 = i_hbusreq2 & ~n35058;
  assign n35078 = controllable_hgrant4 & ~n3928;
  assign n35079 = ~n5454 & ~n35078;
  assign n35080 = ~i_hbusreq2 & ~n35079;
  assign n35081 = ~n35077 & ~n35080;
  assign n35082 = ~controllable_hgrant2 & ~n35081;
  assign n35083 = ~n3859 & ~n35082;
  assign n35084 = controllable_hmaster0 & ~n35083;
  assign n35085 = ~i_hbusreq2 & ~n5471;
  assign n35086 = ~n35067 & ~n35085;
  assign n35087 = ~controllable_hgrant2 & ~n35086;
  assign n35088 = ~n5461 & ~n35087;
  assign n35089 = ~controllable_hmaster0 & ~n35088;
  assign n35090 = ~n35084 & ~n35089;
  assign n35091 = ~controllable_hmaster1 & ~n35090;
  assign n35092 = ~n35076 & ~n35091;
  assign n35093 = ~i_hbusreq3 & ~n35092;
  assign n35094 = ~n35066 & ~n35093;
  assign n35095 = ~controllable_hmaster2 & ~n35094;
  assign n35096 = ~n35050 & ~n35095;
  assign n35097 = ~controllable_hgrant3 & ~n35096;
  assign n35098 = ~n5402 & ~n35097;
  assign n35099 = controllable_nhgrant0 & ~n35098;
  assign n35100 = ~n5534 & ~n35099;
  assign n35101 = ~n3281 & ~n35100;
  assign n35102 = ~n3950 & ~n35101;
  assign n35103 = ~n3378 & ~n35102;
  assign n35104 = ~n35037 & ~n35103;
  assign n35105 = n3492 & ~n35104;
  assign n35106 = ~n3631 & ~n35105;
  assign n35107 = n3485 & ~n35106;
  assign n35108 = ~n3630 & ~n35107;
  assign n35109 = ~n3476 & ~n35108;
  assign n35110 = ~n5621 & ~n34239;
  assign n35111 = ~controllable_hgrant2 & ~n35110;
  assign n35112 = ~n5616 & ~n35111;
  assign n35113 = controllable_hmaster1 & ~n35112;
  assign n35114 = controllable_hmaster0 & ~n35112;
  assign n35115 = ~n5621 & ~n34195;
  assign n35116 = ~controllable_hgrant2 & ~n35115;
  assign n35117 = ~n5616 & ~n35116;
  assign n35118 = ~controllable_hmaster0 & ~n35117;
  assign n35119 = ~n35114 & ~n35118;
  assign n35120 = ~controllable_hmaster1 & ~n35119;
  assign n35121 = ~n35113 & ~n35120;
  assign n35122 = i_hbusreq3 & ~n35121;
  assign n35123 = i_hbusreq2 & ~n35110;
  assign n35124 = ~n5649 & ~n34254;
  assign n35125 = ~i_hbusreq2 & ~n35124;
  assign n35126 = ~n35123 & ~n35125;
  assign n35127 = ~controllable_hgrant2 & ~n35126;
  assign n35128 = ~n5635 & ~n35127;
  assign n35129 = controllable_hmaster1 & ~n35128;
  assign n35130 = controllable_hmaster0 & ~n35128;
  assign n35131 = i_hbusreq2 & ~n35115;
  assign n35132 = ~n5667 & ~n34214;
  assign n35133 = ~i_hbusreq2 & ~n35132;
  assign n35134 = ~n35131 & ~n35133;
  assign n35135 = ~controllable_hgrant2 & ~n35134;
  assign n35136 = ~n5657 & ~n35135;
  assign n35137 = ~controllable_hmaster0 & ~n35136;
  assign n35138 = ~n35130 & ~n35137;
  assign n35139 = ~controllable_hmaster1 & ~n35138;
  assign n35140 = ~n35129 & ~n35139;
  assign n35141 = ~i_hbusreq3 & ~n35140;
  assign n35142 = ~n35122 & ~n35141;
  assign n35143 = controllable_hmaster2 & ~n35142;
  assign n35144 = controllable_hgrant4 & ~n6008;
  assign n35145 = ~n5681 & ~n35144;
  assign n35146 = ~controllable_hgrant2 & ~n35145;
  assign n35147 = ~n5616 & ~n35146;
  assign n35148 = controllable_hmaster0 & ~n35147;
  assign n35149 = ~n5686 & ~n35146;
  assign n35150 = ~controllable_hmaster0 & ~n35149;
  assign n35151 = ~n35148 & ~n35150;
  assign n35152 = controllable_hmaster1 & ~n35151;
  assign n35153 = ~n5697 & ~n35144;
  assign n35154 = ~controllable_hgrant2 & ~n35153;
  assign n35155 = ~n5616 & ~n35154;
  assign n35156 = controllable_hmaster0 & ~n35155;
  assign n35157 = ~controllable_hmaster0 & ~n35147;
  assign n35158 = ~n35156 & ~n35157;
  assign n35159 = ~controllable_hmaster1 & ~n35158;
  assign n35160 = ~n35152 & ~n35159;
  assign n35161 = i_hbusreq3 & ~n35160;
  assign n35162 = i_hbusreq2 & ~n35145;
  assign n35163 = controllable_hgrant4 & ~n15372;
  assign n35164 = ~n5715 & ~n35163;
  assign n35165 = ~i_hbusreq2 & ~n35164;
  assign n35166 = ~n35162 & ~n35165;
  assign n35167 = ~controllable_hgrant2 & ~n35166;
  assign n35168 = ~n5635 & ~n35167;
  assign n35169 = controllable_hmaster0 & ~n35168;
  assign n35170 = ~n5722 & ~n35167;
  assign n35171 = ~controllable_hmaster0 & ~n35170;
  assign n35172 = ~n35169 & ~n35171;
  assign n35173 = controllable_hmaster1 & ~n35172;
  assign n35174 = i_hbusreq2 & ~n35153;
  assign n35175 = ~n5739 & ~n35163;
  assign n35176 = ~i_hbusreq2 & ~n35175;
  assign n35177 = ~n35174 & ~n35176;
  assign n35178 = ~controllable_hgrant2 & ~n35177;
  assign n35179 = ~n5635 & ~n35178;
  assign n35180 = controllable_hmaster0 & ~n35179;
  assign n35181 = ~controllable_hmaster0 & ~n35168;
  assign n35182 = ~n35180 & ~n35181;
  assign n35183 = ~controllable_hmaster1 & ~n35182;
  assign n35184 = ~n35173 & ~n35183;
  assign n35185 = ~i_hbusreq3 & ~n35184;
  assign n35186 = ~n35161 & ~n35185;
  assign n35187 = ~controllable_hmaster2 & ~n35186;
  assign n35188 = ~n35143 & ~n35187;
  assign n35189 = ~controllable_hgrant3 & ~n35188;
  assign n35190 = ~n5615 & ~n35189;
  assign n35191 = controllable_nhgrant0 & ~n35190;
  assign n35192 = ~n5809 & ~n35191;
  assign n35193 = ~n3281 & ~n35192;
  assign n35194 = ~n4089 & ~n35193;
  assign n35195 = n3378 & ~n35194;
  assign n35196 = controllable_hgrant4 & ~n15428;
  assign n35197 = ~n5877 & ~n35196;
  assign n35198 = ~i_hbusreq2 & ~n35197;
  assign n35199 = ~n35123 & ~n35198;
  assign n35200 = ~controllable_hgrant2 & ~n35199;
  assign n35201 = ~n5862 & ~n35200;
  assign n35202 = controllable_hmaster1 & ~n35201;
  assign n35203 = controllable_hmaster0 & ~n35201;
  assign n35204 = ~n5897 & ~n34214;
  assign n35205 = ~i_hbusreq2 & ~n35204;
  assign n35206 = ~n35131 & ~n35205;
  assign n35207 = ~controllable_hgrant2 & ~n35206;
  assign n35208 = ~n5862 & ~n35207;
  assign n35209 = ~controllable_hmaster0 & ~n35208;
  assign n35210 = ~n35203 & ~n35209;
  assign n35211 = ~controllable_hmaster1 & ~n35210;
  assign n35212 = ~n35202 & ~n35211;
  assign n35213 = ~i_hbusreq3 & ~n35212;
  assign n35214 = ~n35122 & ~n35213;
  assign n35215 = controllable_hmaster2 & ~n35214;
  assign n35216 = ~n5911 & ~n35144;
  assign n35217 = ~controllable_hgrant2 & ~n35216;
  assign n35218 = ~n5616 & ~n35217;
  assign n35219 = controllable_hmaster0 & ~n35218;
  assign n35220 = ~n5686 & ~n35217;
  assign n35221 = ~controllable_hmaster0 & ~n35220;
  assign n35222 = ~n35219 & ~n35221;
  assign n35223 = controllable_hmaster1 & ~n35222;
  assign n35224 = ~n5921 & ~n35144;
  assign n35225 = ~controllable_hgrant2 & ~n35224;
  assign n35226 = ~n5616 & ~n35225;
  assign n35227 = controllable_hmaster0 & ~n35226;
  assign n35228 = ~controllable_hmaster0 & ~n35218;
  assign n35229 = ~n35227 & ~n35228;
  assign n35230 = ~controllable_hmaster1 & ~n35229;
  assign n35231 = ~n35223 & ~n35230;
  assign n35232 = i_hbusreq3 & ~n35231;
  assign n35233 = i_hbusreq2 & ~n35216;
  assign n35234 = controllable_hgrant4 & ~n6026;
  assign n35235 = ~n5943 & ~n35234;
  assign n35236 = ~i_hbusreq2 & ~n35235;
  assign n35237 = ~n35233 & ~n35236;
  assign n35238 = ~controllable_hgrant2 & ~n35237;
  assign n35239 = ~n5862 & ~n35238;
  assign n35240 = controllable_hmaster0 & ~n35239;
  assign n35241 = ~n5950 & ~n35238;
  assign n35242 = ~controllable_hmaster0 & ~n35241;
  assign n35243 = ~n35240 & ~n35242;
  assign n35244 = controllable_hmaster1 & ~n35243;
  assign n35245 = i_hbusreq2 & ~n35224;
  assign n35246 = ~n5974 & ~n35234;
  assign n35247 = ~i_hbusreq2 & ~n35246;
  assign n35248 = ~n35245 & ~n35247;
  assign n35249 = ~controllable_hgrant2 & ~n35248;
  assign n35250 = ~n5862 & ~n35249;
  assign n35251 = controllable_hmaster0 & ~n35250;
  assign n35252 = controllable_hgrant4 & ~n6826;
  assign n35253 = ~n5990 & ~n35252;
  assign n35254 = ~i_hbusreq2 & ~n35253;
  assign n35255 = ~n35233 & ~n35254;
  assign n35256 = ~controllable_hgrant2 & ~n35255;
  assign n35257 = ~n5981 & ~n35256;
  assign n35258 = ~controllable_hmaster0 & ~n35257;
  assign n35259 = ~n35251 & ~n35258;
  assign n35260 = ~controllable_hmaster1 & ~n35259;
  assign n35261 = ~n35244 & ~n35260;
  assign n35262 = ~i_hbusreq3 & ~n35261;
  assign n35263 = ~n35232 & ~n35262;
  assign n35264 = ~controllable_hmaster2 & ~n35263;
  assign n35265 = ~n35215 & ~n35264;
  assign n35266 = ~controllable_hgrant3 & ~n35265;
  assign n35267 = ~n5861 & ~n35266;
  assign n35268 = controllable_nhgrant0 & ~n35267;
  assign n35269 = ~n6082 & ~n35268;
  assign n35270 = ~n3281 & ~n35269;
  assign n35271 = ~n4089 & ~n35270;
  assign n35272 = ~n3378 & ~n35271;
  assign n35273 = ~n35195 & ~n35272;
  assign n35274 = n3492 & ~n35273;
  assign n35275 = ~n34979 & ~n35274;
  assign n35276 = n3485 & ~n35275;
  assign n35277 = ~n34978 & ~n35276;
  assign n35278 = n3476 & ~n35277;
  assign n35279 = ~n35109 & ~n35278;
  assign n35280 = n3374 & ~n35279;
  assign n35281 = ~n34985 & ~n35280;
  assign n35282 = n3655 & ~n35281;
  assign n35283 = ~n6100 & ~n34055;
  assign n35284 = ~controllable_hgrant2 & ~n35283;
  assign n35285 = ~n3410 & ~n35284;
  assign n35286 = controllable_hmaster1 & ~n35285;
  assign n35287 = controllable_hmaster0 & ~n35285;
  assign n35288 = ~n34022 & ~n35287;
  assign n35289 = ~controllable_hmaster1 & ~n35288;
  assign n35290 = ~n35286 & ~n35289;
  assign n35291 = i_hbusreq3 & ~n35290;
  assign n35292 = i_hbusreq2 & ~n35283;
  assign n35293 = ~n6123 & ~n34950;
  assign n35294 = ~i_hbusreq2 & ~n35293;
  assign n35295 = ~n35292 & ~n35294;
  assign n35296 = ~controllable_hgrant2 & ~n35295;
  assign n35297 = ~n3859 & ~n35296;
  assign n35298 = controllable_hmaster1 & ~n35297;
  assign n35299 = controllable_hmaster0 & ~n35297;
  assign n35300 = ~n34040 & ~n35299;
  assign n35301 = ~controllable_hmaster1 & ~n35300;
  assign n35302 = ~n35298 & ~n35301;
  assign n35303 = ~i_hbusreq3 & ~n35302;
  assign n35304 = ~n35291 & ~n35303;
  assign n35305 = controllable_hmaster2 & ~n35304;
  assign n35306 = ~n6188 & ~n35305;
  assign n35307 = ~controllable_hgrant3 & ~n35306;
  assign n35308 = ~n5037 & ~n35307;
  assign n35309 = controllable_nhgrant0 & ~n35308;
  assign n35310 = ~n5245 & ~n35309;
  assign n35311 = ~n3281 & ~n35310;
  assign n35312 = ~n3783 & ~n35311;
  assign n35313 = ~n3378 & ~n35312;
  assign n35314 = ~n34939 & ~n35313;
  assign n35315 = n3492 & ~n35314;
  assign n35316 = ~n3631 & ~n35315;
  assign n35317 = n3485 & ~n35316;
  assign n35318 = ~n3630 & ~n35317;
  assign n35319 = ~n3476 & ~n35318;
  assign n35320 = ~n34979 & ~n35315;
  assign n35321 = n3485 & ~n35320;
  assign n35322 = ~n34978 & ~n35321;
  assign n35323 = n3476 & ~n35322;
  assign n35324 = ~n35319 & ~n35323;
  assign n35325 = ~n3374 & ~n35324;
  assign n35326 = ~n34344 & ~n35029;
  assign n35327 = ~controllable_hgrant3 & ~n35326;
  assign n35328 = ~n5287 & ~n35327;
  assign n35329 = controllable_nhgrant0 & ~n35328;
  assign n35330 = ~n5363 & ~n35329;
  assign n35331 = ~n3281 & ~n35330;
  assign n35332 = ~n3950 & ~n35331;
  assign n35333 = n3378 & ~n35332;
  assign n35334 = ~n6212 & ~n34055;
  assign n35335 = ~controllable_hgrant2 & ~n35334;
  assign n35336 = ~n3410 & ~n35335;
  assign n35337 = controllable_hmaster1 & ~n35336;
  assign n35338 = controllable_hmaster0 & ~n35336;
  assign n35339 = ~n34309 & ~n35338;
  assign n35340 = ~controllable_hmaster1 & ~n35339;
  assign n35341 = ~n35337 & ~n35340;
  assign n35342 = i_hbusreq3 & ~n35341;
  assign n35343 = i_hbusreq2 & ~n35334;
  assign n35344 = ~n6233 & ~n34950;
  assign n35345 = ~i_hbusreq2 & ~n35344;
  assign n35346 = ~n35343 & ~n35345;
  assign n35347 = ~controllable_hgrant2 & ~n35346;
  assign n35348 = ~n3859 & ~n35347;
  assign n35349 = controllable_hmaster1 & ~n35348;
  assign n35350 = controllable_hmaster0 & ~n35348;
  assign n35351 = ~n34320 & ~n35350;
  assign n35352 = ~controllable_hmaster1 & ~n35351;
  assign n35353 = ~n35349 & ~n35352;
  assign n35354 = ~i_hbusreq3 & ~n35353;
  assign n35355 = ~n35342 & ~n35354;
  assign n35356 = controllable_hmaster2 & ~n35355;
  assign n35357 = ~n6250 & ~n34986;
  assign n35358 = ~controllable_hgrant2 & ~n35357;
  assign n35359 = ~n3410 & ~n35358;
  assign n35360 = controllable_hmaster0 & ~n35359;
  assign n35361 = ~n5288 & ~n35358;
  assign n35362 = ~controllable_hmaster0 & ~n35361;
  assign n35363 = ~n35360 & ~n35362;
  assign n35364 = controllable_hmaster1 & ~n35363;
  assign n35365 = ~n6264 & ~n34986;
  assign n35366 = ~controllable_hgrant2 & ~n35365;
  assign n35367 = ~n3410 & ~n35366;
  assign n35368 = controllable_hmaster0 & ~n35367;
  assign n35369 = ~controllable_hmaster0 & ~n35359;
  assign n35370 = ~n35368 & ~n35369;
  assign n35371 = ~controllable_hmaster1 & ~n35370;
  assign n35372 = ~n35364 & ~n35371;
  assign n35373 = i_hbusreq3 & ~n35372;
  assign n35374 = i_hbusreq2 & ~n35357;
  assign n35375 = ~n6287 & ~n35078;
  assign n35376 = ~i_hbusreq2 & ~n35375;
  assign n35377 = ~n35374 & ~n35376;
  assign n35378 = ~controllable_hgrant2 & ~n35377;
  assign n35379 = ~n3859 & ~n35378;
  assign n35380 = controllable_hmaster0 & ~n35379;
  assign n35381 = ~n5438 & ~n35378;
  assign n35382 = ~controllable_hmaster0 & ~n35381;
  assign n35383 = ~n35380 & ~n35382;
  assign n35384 = controllable_hmaster1 & ~n35383;
  assign n35385 = i_hbusreq2 & ~n35365;
  assign n35386 = ~n6315 & ~n35078;
  assign n35387 = ~i_hbusreq2 & ~n35386;
  assign n35388 = ~n35385 & ~n35387;
  assign n35389 = ~controllable_hgrant2 & ~n35388;
  assign n35390 = ~n3859 & ~n35389;
  assign n35391 = controllable_hmaster0 & ~n35390;
  assign n35392 = controllable_hgrant4 & ~n5471;
  assign n35393 = ~n6331 & ~n35392;
  assign n35394 = ~i_hbusreq2 & ~n35393;
  assign n35395 = ~n35374 & ~n35394;
  assign n35396 = ~controllable_hgrant2 & ~n35395;
  assign n35397 = ~n5461 & ~n35396;
  assign n35398 = ~controllable_hmaster0 & ~n35397;
  assign n35399 = ~n35391 & ~n35398;
  assign n35400 = ~controllable_hmaster1 & ~n35399;
  assign n35401 = ~n35384 & ~n35400;
  assign n35402 = ~i_hbusreq3 & ~n35401;
  assign n35403 = ~n35373 & ~n35402;
  assign n35404 = ~controllable_hmaster2 & ~n35403;
  assign n35405 = ~n35356 & ~n35404;
  assign n35406 = ~controllable_hgrant3 & ~n35405;
  assign n35407 = ~n5402 & ~n35406;
  assign n35408 = controllable_nhgrant0 & ~n35407;
  assign n35409 = ~n5534 & ~n35408;
  assign n35410 = ~n3281 & ~n35409;
  assign n35411 = ~n3950 & ~n35410;
  assign n35412 = ~n3378 & ~n35411;
  assign n35413 = ~n35333 & ~n35412;
  assign n35414 = n3492 & ~n35413;
  assign n35415 = ~n3631 & ~n35414;
  assign n35416 = n3485 & ~n35415;
  assign n35417 = ~n3630 & ~n35416;
  assign n35418 = ~n3476 & ~n35417;
  assign n35419 = ~n6359 & ~n34195;
  assign n35420 = ~controllable_hgrant2 & ~n35419;
  assign n35421 = ~n5616 & ~n35420;
  assign n35422 = ~controllable_hmaster0 & ~n35421;
  assign n35423 = ~n35114 & ~n35422;
  assign n35424 = ~controllable_hmaster1 & ~n35423;
  assign n35425 = ~n35113 & ~n35424;
  assign n35426 = i_hbusreq3 & ~n35425;
  assign n35427 = i_hbusreq2 & ~n35419;
  assign n35428 = ~n6380 & ~n34214;
  assign n35429 = ~i_hbusreq2 & ~n35428;
  assign n35430 = ~n35427 & ~n35429;
  assign n35431 = ~controllable_hgrant2 & ~n35430;
  assign n35432 = ~n5657 & ~n35431;
  assign n35433 = ~controllable_hmaster0 & ~n35432;
  assign n35434 = ~n35130 & ~n35433;
  assign n35435 = ~controllable_hmaster1 & ~n35434;
  assign n35436 = ~n35129 & ~n35435;
  assign n35437 = ~i_hbusreq3 & ~n35436;
  assign n35438 = ~n35426 & ~n35437;
  assign n35439 = controllable_hmaster2 & ~n35438;
  assign n35440 = ~n35187 & ~n35439;
  assign n35441 = ~controllable_hgrant3 & ~n35440;
  assign n35442 = ~n5615 & ~n35441;
  assign n35443 = controllable_nhgrant0 & ~n35442;
  assign n35444 = ~n5809 & ~n35443;
  assign n35445 = ~n3281 & ~n35444;
  assign n35446 = ~n4089 & ~n35445;
  assign n35447 = n3378 & ~n35446;
  assign n35448 = ~n6403 & ~n34239;
  assign n35449 = ~controllable_hgrant2 & ~n35448;
  assign n35450 = ~n5616 & ~n35449;
  assign n35451 = controllable_hmaster1 & ~n35450;
  assign n35452 = controllable_hmaster0 & ~n35450;
  assign n35453 = ~n6403 & ~n34195;
  assign n35454 = ~controllable_hgrant2 & ~n35453;
  assign n35455 = ~n5616 & ~n35454;
  assign n35456 = ~controllable_hmaster0 & ~n35455;
  assign n35457 = ~n35452 & ~n35456;
  assign n35458 = ~controllable_hmaster1 & ~n35457;
  assign n35459 = ~n35451 & ~n35458;
  assign n35460 = i_hbusreq3 & ~n35459;
  assign n35461 = i_hbusreq2 & ~n35448;
  assign n35462 = ~n6433 & ~n35196;
  assign n35463 = ~i_hbusreq2 & ~n35462;
  assign n35464 = ~n35461 & ~n35463;
  assign n35465 = ~controllable_hgrant2 & ~n35464;
  assign n35466 = ~n5862 & ~n35465;
  assign n35467 = controllable_hmaster1 & ~n35466;
  assign n35468 = controllable_hmaster0 & ~n35466;
  assign n35469 = i_hbusreq2 & ~n35453;
  assign n35470 = ~n6451 & ~n34214;
  assign n35471 = ~i_hbusreq2 & ~n35470;
  assign n35472 = ~n35469 & ~n35471;
  assign n35473 = ~controllable_hgrant2 & ~n35472;
  assign n35474 = ~n5862 & ~n35473;
  assign n35475 = ~controllable_hmaster0 & ~n35474;
  assign n35476 = ~n35468 & ~n35475;
  assign n35477 = ~controllable_hmaster1 & ~n35476;
  assign n35478 = ~n35467 & ~n35477;
  assign n35479 = ~i_hbusreq3 & ~n35478;
  assign n35480 = ~n35460 & ~n35479;
  assign n35481 = controllable_hmaster2 & ~n35480;
  assign n35482 = ~n6465 & ~n35144;
  assign n35483 = ~controllable_hgrant2 & ~n35482;
  assign n35484 = ~n5616 & ~n35483;
  assign n35485 = controllable_hmaster0 & ~n35484;
  assign n35486 = ~n5686 & ~n35483;
  assign n35487 = ~controllable_hmaster0 & ~n35486;
  assign n35488 = ~n35485 & ~n35487;
  assign n35489 = controllable_hmaster1 & ~n35488;
  assign n35490 = ~n6476 & ~n35144;
  assign n35491 = ~controllable_hgrant2 & ~n35490;
  assign n35492 = ~n5616 & ~n35491;
  assign n35493 = controllable_hmaster0 & ~n35492;
  assign n35494 = ~controllable_hmaster0 & ~n35484;
  assign n35495 = ~n35493 & ~n35494;
  assign n35496 = ~controllable_hmaster1 & ~n35495;
  assign n35497 = ~n35489 & ~n35496;
  assign n35498 = i_hbusreq3 & ~n35497;
  assign n35499 = i_hbusreq2 & ~n35482;
  assign n35500 = ~n6498 & ~n35234;
  assign n35501 = ~i_hbusreq2 & ~n35500;
  assign n35502 = ~n35499 & ~n35501;
  assign n35503 = ~controllable_hgrant2 & ~n35502;
  assign n35504 = ~n5862 & ~n35503;
  assign n35505 = controllable_hmaster0 & ~n35504;
  assign n35506 = ~n5950 & ~n35503;
  assign n35507 = ~controllable_hmaster0 & ~n35506;
  assign n35508 = ~n35505 & ~n35507;
  assign n35509 = controllable_hmaster1 & ~n35508;
  assign n35510 = i_hbusreq2 & ~n35490;
  assign n35511 = ~n6528 & ~n35234;
  assign n35512 = ~i_hbusreq2 & ~n35511;
  assign n35513 = ~n35510 & ~n35512;
  assign n35514 = ~controllable_hgrant2 & ~n35513;
  assign n35515 = ~n5862 & ~n35514;
  assign n35516 = controllable_hmaster0 & ~n35515;
  assign n35517 = ~n6542 & ~n35252;
  assign n35518 = ~i_hbusreq2 & ~n35517;
  assign n35519 = ~n35499 & ~n35518;
  assign n35520 = ~controllable_hgrant2 & ~n35519;
  assign n35521 = ~n5981 & ~n35520;
  assign n35522 = ~controllable_hmaster0 & ~n35521;
  assign n35523 = ~n35516 & ~n35522;
  assign n35524 = ~controllable_hmaster1 & ~n35523;
  assign n35525 = ~n35509 & ~n35524;
  assign n35526 = ~i_hbusreq3 & ~n35525;
  assign n35527 = ~n35498 & ~n35526;
  assign n35528 = ~controllable_hmaster2 & ~n35527;
  assign n35529 = ~n35481 & ~n35528;
  assign n35530 = ~controllable_hgrant3 & ~n35529;
  assign n35531 = ~n5861 & ~n35530;
  assign n35532 = controllable_nhgrant0 & ~n35531;
  assign n35533 = ~n6082 & ~n35532;
  assign n35534 = ~n3281 & ~n35533;
  assign n35535 = ~n4089 & ~n35534;
  assign n35536 = ~n3378 & ~n35535;
  assign n35537 = ~n35447 & ~n35536;
  assign n35538 = n3492 & ~n35537;
  assign n35539 = ~n34979 & ~n35538;
  assign n35540 = n3485 & ~n35539;
  assign n35541 = ~n34978 & ~n35540;
  assign n35542 = n3476 & ~n35541;
  assign n35543 = ~n35418 & ~n35542;
  assign n35544 = n3374 & ~n35543;
  assign n35545 = ~n35325 & ~n35544;
  assign n35546 = ~n3655 & ~n35545;
  assign n35547 = ~n35282 & ~n35546;
  assign n35548 = n3652 & ~n35547;
  assign n35549 = ~n4333 & ~n34941;
  assign n35550 = controllable_hmaster1 & ~n35549;
  assign n35551 = controllable_hmaster0 & ~n35549;
  assign n35552 = ~n34022 & ~n35551;
  assign n35553 = ~controllable_hmaster1 & ~n35552;
  assign n35554 = ~n35550 & ~n35553;
  assign n35555 = i_hbusreq3 & ~n35554;
  assign n35556 = ~n4340 & ~n34954;
  assign n35557 = controllable_hmaster1 & ~n35556;
  assign n35558 = controllable_hmaster0 & ~n35556;
  assign n35559 = ~n34040 & ~n35558;
  assign n35560 = ~controllable_hmaster1 & ~n35559;
  assign n35561 = ~n35557 & ~n35560;
  assign n35562 = ~i_hbusreq3 & ~n35561;
  assign n35563 = ~n35555 & ~n35562;
  assign n35564 = controllable_hmaster2 & ~n35563;
  assign n35565 = ~n6657 & ~n35564;
  assign n35566 = ~controllable_hgrant3 & ~n35565;
  assign n35567 = ~n5037 & ~n35566;
  assign n35568 = controllable_nhgrant0 & ~n35567;
  assign n35569 = ~n5245 & ~n35568;
  assign n35570 = ~n3281 & ~n35569;
  assign n35571 = ~n3783 & ~n35570;
  assign n35572 = ~n3378 & ~n35571;
  assign n35573 = ~n34939 & ~n35572;
  assign n35574 = n3492 & ~n35573;
  assign n35575 = ~n3631 & ~n35574;
  assign n35576 = n3485 & ~n35575;
  assign n35577 = ~n3630 & ~n35576;
  assign n35578 = ~n3476 & ~n35577;
  assign n35579 = ~n34979 & ~n35574;
  assign n35580 = n3485 & ~n35579;
  assign n35581 = ~n34978 & ~n35580;
  assign n35582 = n3476 & ~n35581;
  assign n35583 = ~n35578 & ~n35582;
  assign n35584 = ~n3374 & ~n35583;
  assign n35585 = ~n34460 & ~n35029;
  assign n35586 = ~controllable_hgrant3 & ~n35585;
  assign n35587 = ~n5287 & ~n35586;
  assign n35588 = controllable_nhgrant0 & ~n35587;
  assign n35589 = ~n5363 & ~n35588;
  assign n35590 = ~n3281 & ~n35589;
  assign n35591 = ~n3950 & ~n35590;
  assign n35592 = n3378 & ~n35591;
  assign n35593 = ~n4333 & ~n34153;
  assign n35594 = controllable_hmaster1 & ~n35593;
  assign n35595 = controllable_hmaster0 & ~n35593;
  assign n35596 = ~n34430 & ~n35595;
  assign n35597 = ~controllable_hmaster1 & ~n35596;
  assign n35598 = ~n35594 & ~n35597;
  assign n35599 = i_hbusreq3 & ~n35598;
  assign n35600 = ~n4340 & ~n35041;
  assign n35601 = controllable_hmaster1 & ~n35600;
  assign n35602 = controllable_hmaster0 & ~n35600;
  assign n35603 = ~n34436 & ~n35602;
  assign n35604 = ~controllable_hmaster1 & ~n35603;
  assign n35605 = ~n35601 & ~n35604;
  assign n35606 = ~i_hbusreq3 & ~n35605;
  assign n35607 = ~n35599 & ~n35606;
  assign n35608 = controllable_hmaster2 & ~n35607;
  assign n35609 = ~n4333 & ~n35051;
  assign n35610 = controllable_hmaster0 & ~n35609;
  assign n35611 = ~n6697 & ~n35051;
  assign n35612 = ~controllable_hmaster0 & ~n35611;
  assign n35613 = ~n35610 & ~n35612;
  assign n35614 = controllable_hmaster1 & ~n35613;
  assign n35615 = ~n4333 & ~n35059;
  assign n35616 = controllable_hmaster0 & ~n35615;
  assign n35617 = ~controllable_hmaster0 & ~n35609;
  assign n35618 = ~n35616 & ~n35617;
  assign n35619 = ~controllable_hmaster1 & ~n35618;
  assign n35620 = ~n35614 & ~n35619;
  assign n35621 = i_hbusreq3 & ~n35620;
  assign n35622 = ~n4340 & ~n35070;
  assign n35623 = controllable_hmaster0 & ~n35622;
  assign n35624 = ~n6710 & ~n35070;
  assign n35625 = ~controllable_hmaster0 & ~n35624;
  assign n35626 = ~n35623 & ~n35625;
  assign n35627 = controllable_hmaster1 & ~n35626;
  assign n35628 = ~n4340 & ~n35082;
  assign n35629 = controllable_hmaster0 & ~n35628;
  assign n35630 = ~n6947 & ~n35087;
  assign n35631 = ~controllable_hmaster0 & ~n35630;
  assign n35632 = ~n35629 & ~n35631;
  assign n35633 = ~controllable_hmaster1 & ~n35632;
  assign n35634 = ~n35627 & ~n35633;
  assign n35635 = ~i_hbusreq3 & ~n35634;
  assign n35636 = ~n35621 & ~n35635;
  assign n35637 = ~controllable_hmaster2 & ~n35636;
  assign n35638 = ~n35608 & ~n35637;
  assign n35639 = ~controllable_hgrant3 & ~n35638;
  assign n35640 = ~n5402 & ~n35639;
  assign n35641 = controllable_nhgrant0 & ~n35640;
  assign n35642 = ~n5534 & ~n35641;
  assign n35643 = ~n3281 & ~n35642;
  assign n35644 = ~n3950 & ~n35643;
  assign n35645 = ~n3378 & ~n35644;
  assign n35646 = ~n35592 & ~n35645;
  assign n35647 = n3492 & ~n35646;
  assign n35648 = ~n3631 & ~n35647;
  assign n35649 = n3485 & ~n35648;
  assign n35650 = ~n3630 & ~n35649;
  assign n35651 = ~n3476 & ~n35650;
  assign n35652 = ~n6738 & ~n35116;
  assign n35653 = ~controllable_hmaster0 & ~n35652;
  assign n35654 = ~n35114 & ~n35653;
  assign n35655 = ~controllable_hmaster1 & ~n35654;
  assign n35656 = ~n35113 & ~n35655;
  assign n35657 = i_hbusreq3 & ~n35656;
  assign n35658 = ~n6745 & ~n35135;
  assign n35659 = ~controllable_hmaster0 & ~n35658;
  assign n35660 = ~n35130 & ~n35659;
  assign n35661 = ~controllable_hmaster1 & ~n35660;
  assign n35662 = ~n35129 & ~n35661;
  assign n35663 = ~i_hbusreq3 & ~n35662;
  assign n35664 = ~n35657 & ~n35663;
  assign n35665 = controllable_hmaster2 & ~n35664;
  assign n35666 = ~n35187 & ~n35665;
  assign n35667 = ~controllable_hgrant3 & ~n35666;
  assign n35668 = ~n5615 & ~n35667;
  assign n35669 = controllable_nhgrant0 & ~n35668;
  assign n35670 = ~n5809 & ~n35669;
  assign n35671 = ~n3281 & ~n35670;
  assign n35672 = ~n4089 & ~n35671;
  assign n35673 = n3378 & ~n35672;
  assign n35674 = ~n6762 & ~n35111;
  assign n35675 = controllable_hmaster1 & ~n35674;
  assign n35676 = controllable_hmaster0 & ~n35674;
  assign n35677 = ~n6762 & ~n35116;
  assign n35678 = ~controllable_hmaster0 & ~n35677;
  assign n35679 = ~n35676 & ~n35678;
  assign n35680 = ~controllable_hmaster1 & ~n35679;
  assign n35681 = ~n35675 & ~n35680;
  assign n35682 = i_hbusreq3 & ~n35681;
  assign n35683 = ~n6772 & ~n35200;
  assign n35684 = controllable_hmaster1 & ~n35683;
  assign n35685 = controllable_hmaster0 & ~n35683;
  assign n35686 = ~n6772 & ~n35207;
  assign n35687 = ~controllable_hmaster0 & ~n35686;
  assign n35688 = ~n35685 & ~n35687;
  assign n35689 = ~controllable_hmaster1 & ~n35688;
  assign n35690 = ~n35684 & ~n35689;
  assign n35691 = ~i_hbusreq3 & ~n35690;
  assign n35692 = ~n35682 & ~n35691;
  assign n35693 = controllable_hmaster2 & ~n35692;
  assign n35694 = ~n6762 & ~n35217;
  assign n35695 = controllable_hmaster0 & ~n35694;
  assign n35696 = ~n6786 & ~n35217;
  assign n35697 = ~controllable_hmaster0 & ~n35696;
  assign n35698 = ~n35695 & ~n35697;
  assign n35699 = controllable_hmaster1 & ~n35698;
  assign n35700 = ~n6762 & ~n35225;
  assign n35701 = controllable_hmaster0 & ~n35700;
  assign n35702 = ~controllable_hmaster0 & ~n35694;
  assign n35703 = ~n35701 & ~n35702;
  assign n35704 = ~controllable_hmaster1 & ~n35703;
  assign n35705 = ~n35699 & ~n35704;
  assign n35706 = i_hbusreq3 & ~n35705;
  assign n35707 = ~n6772 & ~n35238;
  assign n35708 = controllable_hmaster0 & ~n35707;
  assign n35709 = ~n6813 & ~n35238;
  assign n35710 = ~controllable_hmaster0 & ~n35709;
  assign n35711 = ~n35708 & ~n35710;
  assign n35712 = controllable_hmaster1 & ~n35711;
  assign n35713 = ~n6772 & ~n35249;
  assign n35714 = controllable_hmaster0 & ~n35713;
  assign n35715 = ~n6831 & ~n35256;
  assign n35716 = ~controllable_hmaster0 & ~n35715;
  assign n35717 = ~n35714 & ~n35716;
  assign n35718 = ~controllable_hmaster1 & ~n35717;
  assign n35719 = ~n35712 & ~n35718;
  assign n35720 = ~i_hbusreq3 & ~n35719;
  assign n35721 = ~n35706 & ~n35720;
  assign n35722 = ~controllable_hmaster2 & ~n35721;
  assign n35723 = ~n35693 & ~n35722;
  assign n35724 = ~controllable_hgrant3 & ~n35723;
  assign n35725 = ~n5861 & ~n35724;
  assign n35726 = controllable_nhgrant0 & ~n35725;
  assign n35727 = ~n6082 & ~n35726;
  assign n35728 = ~n3281 & ~n35727;
  assign n35729 = ~n4089 & ~n35728;
  assign n35730 = ~n3378 & ~n35729;
  assign n35731 = ~n35673 & ~n35730;
  assign n35732 = n3492 & ~n35731;
  assign n35733 = ~n34979 & ~n35732;
  assign n35734 = n3485 & ~n35733;
  assign n35735 = ~n34978 & ~n35734;
  assign n35736 = n3476 & ~n35735;
  assign n35737 = ~n35651 & ~n35736;
  assign n35738 = n3374 & ~n35737;
  assign n35739 = ~n35584 & ~n35738;
  assign n35740 = n3655 & ~n35739;
  assign n35741 = ~n4333 & ~n35284;
  assign n35742 = controllable_hmaster1 & ~n35741;
  assign n35743 = controllable_hmaster0 & ~n35741;
  assign n35744 = ~n34022 & ~n35743;
  assign n35745 = ~controllable_hmaster1 & ~n35744;
  assign n35746 = ~n35742 & ~n35745;
  assign n35747 = i_hbusreq3 & ~n35746;
  assign n35748 = ~n4340 & ~n35296;
  assign n35749 = controllable_hmaster1 & ~n35748;
  assign n35750 = controllable_hmaster0 & ~n35748;
  assign n35751 = ~n34040 & ~n35750;
  assign n35752 = ~controllable_hmaster1 & ~n35751;
  assign n35753 = ~n35749 & ~n35752;
  assign n35754 = ~i_hbusreq3 & ~n35753;
  assign n35755 = ~n35747 & ~n35754;
  assign n35756 = controllable_hmaster2 & ~n35755;
  assign n35757 = ~n6887 & ~n35756;
  assign n35758 = ~controllable_hgrant3 & ~n35757;
  assign n35759 = ~n5037 & ~n35758;
  assign n35760 = controllable_nhgrant0 & ~n35759;
  assign n35761 = ~n5245 & ~n35760;
  assign n35762 = ~n3281 & ~n35761;
  assign n35763 = ~n3783 & ~n35762;
  assign n35764 = ~n3378 & ~n35763;
  assign n35765 = ~n34939 & ~n35764;
  assign n35766 = n3492 & ~n35765;
  assign n35767 = ~n3631 & ~n35766;
  assign n35768 = n3485 & ~n35767;
  assign n35769 = ~n3630 & ~n35768;
  assign n35770 = ~n3476 & ~n35769;
  assign n35771 = ~n34979 & ~n35766;
  assign n35772 = n3485 & ~n35771;
  assign n35773 = ~n34978 & ~n35772;
  assign n35774 = n3476 & ~n35773;
  assign n35775 = ~n35770 & ~n35774;
  assign n35776 = ~n3374 & ~n35775;
  assign n35777 = ~n34560 & ~n35029;
  assign n35778 = ~controllable_hgrant3 & ~n35777;
  assign n35779 = ~n5287 & ~n35778;
  assign n35780 = controllable_nhgrant0 & ~n35779;
  assign n35781 = ~n5363 & ~n35780;
  assign n35782 = ~n3281 & ~n35781;
  assign n35783 = ~n3950 & ~n35782;
  assign n35784 = n3378 & ~n35783;
  assign n35785 = ~n4333 & ~n35335;
  assign n35786 = controllable_hmaster1 & ~n35785;
  assign n35787 = controllable_hmaster0 & ~n35785;
  assign n35788 = ~n34530 & ~n35787;
  assign n35789 = ~controllable_hmaster1 & ~n35788;
  assign n35790 = ~n35786 & ~n35789;
  assign n35791 = i_hbusreq3 & ~n35790;
  assign n35792 = ~n4340 & ~n35347;
  assign n35793 = controllable_hmaster1 & ~n35792;
  assign n35794 = controllable_hmaster0 & ~n35792;
  assign n35795 = ~n34536 & ~n35794;
  assign n35796 = ~controllable_hmaster1 & ~n35795;
  assign n35797 = ~n35793 & ~n35796;
  assign n35798 = ~i_hbusreq3 & ~n35797;
  assign n35799 = ~n35791 & ~n35798;
  assign n35800 = controllable_hmaster2 & ~n35799;
  assign n35801 = ~n4333 & ~n35358;
  assign n35802 = controllable_hmaster0 & ~n35801;
  assign n35803 = ~n6697 & ~n35358;
  assign n35804 = ~controllable_hmaster0 & ~n35803;
  assign n35805 = ~n35802 & ~n35804;
  assign n35806 = controllable_hmaster1 & ~n35805;
  assign n35807 = ~n4333 & ~n35366;
  assign n35808 = controllable_hmaster0 & ~n35807;
  assign n35809 = ~controllable_hmaster0 & ~n35801;
  assign n35810 = ~n35808 & ~n35809;
  assign n35811 = ~controllable_hmaster1 & ~n35810;
  assign n35812 = ~n35806 & ~n35811;
  assign n35813 = i_hbusreq3 & ~n35812;
  assign n35814 = ~n4340 & ~n35378;
  assign n35815 = controllable_hmaster0 & ~n35814;
  assign n35816 = ~n6710 & ~n35378;
  assign n35817 = ~controllable_hmaster0 & ~n35816;
  assign n35818 = ~n35815 & ~n35817;
  assign n35819 = controllable_hmaster1 & ~n35818;
  assign n35820 = ~n4340 & ~n35389;
  assign n35821 = controllable_hmaster0 & ~n35820;
  assign n35822 = ~n6947 & ~n35396;
  assign n35823 = ~controllable_hmaster0 & ~n35822;
  assign n35824 = ~n35821 & ~n35823;
  assign n35825 = ~controllable_hmaster1 & ~n35824;
  assign n35826 = ~n35819 & ~n35825;
  assign n35827 = ~i_hbusreq3 & ~n35826;
  assign n35828 = ~n35813 & ~n35827;
  assign n35829 = ~controllable_hmaster2 & ~n35828;
  assign n35830 = ~n35800 & ~n35829;
  assign n35831 = ~controllable_hgrant3 & ~n35830;
  assign n35832 = ~n5402 & ~n35831;
  assign n35833 = controllable_nhgrant0 & ~n35832;
  assign n35834 = ~n5534 & ~n35833;
  assign n35835 = ~n3281 & ~n35834;
  assign n35836 = ~n3950 & ~n35835;
  assign n35837 = ~n3378 & ~n35836;
  assign n35838 = ~n35784 & ~n35837;
  assign n35839 = n3492 & ~n35838;
  assign n35840 = ~n3631 & ~n35839;
  assign n35841 = n3485 & ~n35840;
  assign n35842 = ~n3630 & ~n35841;
  assign n35843 = ~n3476 & ~n35842;
  assign n35844 = ~n6738 & ~n35420;
  assign n35845 = ~controllable_hmaster0 & ~n35844;
  assign n35846 = ~n35114 & ~n35845;
  assign n35847 = ~controllable_hmaster1 & ~n35846;
  assign n35848 = ~n35113 & ~n35847;
  assign n35849 = i_hbusreq3 & ~n35848;
  assign n35850 = ~n6745 & ~n35431;
  assign n35851 = ~controllable_hmaster0 & ~n35850;
  assign n35852 = ~n35130 & ~n35851;
  assign n35853 = ~controllable_hmaster1 & ~n35852;
  assign n35854 = ~n35129 & ~n35853;
  assign n35855 = ~i_hbusreq3 & ~n35854;
  assign n35856 = ~n35849 & ~n35855;
  assign n35857 = controllable_hmaster2 & ~n35856;
  assign n35858 = ~n35187 & ~n35857;
  assign n35859 = ~controllable_hgrant3 & ~n35858;
  assign n35860 = ~n5615 & ~n35859;
  assign n35861 = controllable_nhgrant0 & ~n35860;
  assign n35862 = ~n5809 & ~n35861;
  assign n35863 = ~n3281 & ~n35862;
  assign n35864 = ~n4089 & ~n35863;
  assign n35865 = n3378 & ~n35864;
  assign n35866 = ~n6762 & ~n35449;
  assign n35867 = controllable_hmaster1 & ~n35866;
  assign n35868 = controllable_hmaster0 & ~n35866;
  assign n35869 = ~n6762 & ~n35454;
  assign n35870 = ~controllable_hmaster0 & ~n35869;
  assign n35871 = ~n35868 & ~n35870;
  assign n35872 = ~controllable_hmaster1 & ~n35871;
  assign n35873 = ~n35867 & ~n35872;
  assign n35874 = i_hbusreq3 & ~n35873;
  assign n35875 = ~n6772 & ~n35465;
  assign n35876 = controllable_hmaster1 & ~n35875;
  assign n35877 = controllable_hmaster0 & ~n35875;
  assign n35878 = ~n6772 & ~n35473;
  assign n35879 = ~controllable_hmaster0 & ~n35878;
  assign n35880 = ~n35877 & ~n35879;
  assign n35881 = ~controllable_hmaster1 & ~n35880;
  assign n35882 = ~n35876 & ~n35881;
  assign n35883 = ~i_hbusreq3 & ~n35882;
  assign n35884 = ~n35874 & ~n35883;
  assign n35885 = controllable_hmaster2 & ~n35884;
  assign n35886 = ~n6762 & ~n35483;
  assign n35887 = controllable_hmaster0 & ~n35886;
  assign n35888 = ~n6786 & ~n35483;
  assign n35889 = ~controllable_hmaster0 & ~n35888;
  assign n35890 = ~n35887 & ~n35889;
  assign n35891 = controllable_hmaster1 & ~n35890;
  assign n35892 = ~n6762 & ~n35491;
  assign n35893 = controllable_hmaster0 & ~n35892;
  assign n35894 = ~controllable_hmaster0 & ~n35886;
  assign n35895 = ~n35893 & ~n35894;
  assign n35896 = ~controllable_hmaster1 & ~n35895;
  assign n35897 = ~n35891 & ~n35896;
  assign n35898 = i_hbusreq3 & ~n35897;
  assign n35899 = ~n6772 & ~n35503;
  assign n35900 = controllable_hmaster0 & ~n35899;
  assign n35901 = ~n6813 & ~n35503;
  assign n35902 = ~controllable_hmaster0 & ~n35901;
  assign n35903 = ~n35900 & ~n35902;
  assign n35904 = controllable_hmaster1 & ~n35903;
  assign n35905 = ~n6772 & ~n35514;
  assign n35906 = controllable_hmaster0 & ~n35905;
  assign n35907 = ~n6831 & ~n35520;
  assign n35908 = ~controllable_hmaster0 & ~n35907;
  assign n35909 = ~n35906 & ~n35908;
  assign n35910 = ~controllable_hmaster1 & ~n35909;
  assign n35911 = ~n35904 & ~n35910;
  assign n35912 = ~i_hbusreq3 & ~n35911;
  assign n35913 = ~n35898 & ~n35912;
  assign n35914 = ~controllable_hmaster2 & ~n35913;
  assign n35915 = ~n35885 & ~n35914;
  assign n35916 = ~controllable_hgrant3 & ~n35915;
  assign n35917 = ~n5861 & ~n35916;
  assign n35918 = controllable_nhgrant0 & ~n35917;
  assign n35919 = ~n6082 & ~n35918;
  assign n35920 = ~n3281 & ~n35919;
  assign n35921 = ~n4089 & ~n35920;
  assign n35922 = ~n3378 & ~n35921;
  assign n35923 = ~n35865 & ~n35922;
  assign n35924 = n3492 & ~n35923;
  assign n35925 = ~n34979 & ~n35924;
  assign n35926 = n3485 & ~n35925;
  assign n35927 = ~n34978 & ~n35926;
  assign n35928 = n3476 & ~n35927;
  assign n35929 = ~n35843 & ~n35928;
  assign n35930 = n3374 & ~n35929;
  assign n35931 = ~n35776 & ~n35930;
  assign n35932 = ~n3655 & ~n35931;
  assign n35933 = ~n35740 & ~n35932;
  assign n35934 = ~n3652 & ~n35933;
  assign n35935 = ~n35548 & ~n35934;
  assign n35936 = ~n3368 & ~n35935;
  assign n35937 = controllable_hgrant4 & ~n4606;
  assign n35938 = ~n5256 & ~n35937;
  assign n35939 = ~controllable_hgrant2 & ~n35938;
  assign n35940 = ~n3410 & ~n35939;
  assign n35941 = controllable_hmaster1 & ~n35940;
  assign n35942 = controllable_hmaster0 & ~n35940;
  assign n35943 = controllable_hmaster0 & ~n35942;
  assign n35944 = ~controllable_hmaster1 & ~n35943;
  assign n35945 = ~n35941 & ~n35944;
  assign n35946 = i_hbusreq3 & ~n35945;
  assign n35947 = i_hbusreq2 & ~n35938;
  assign n35948 = controllable_hgrant4 & ~n15991;
  assign n35949 = ~n5271 & ~n35948;
  assign n35950 = ~i_hbusreq2 & ~n35949;
  assign n35951 = ~n35947 & ~n35950;
  assign n35952 = ~controllable_hgrant2 & ~n35951;
  assign n35953 = ~n3431 & ~n35952;
  assign n35954 = controllable_hmaster1 & ~n35953;
  assign n35955 = controllable_hmaster0 & ~n35953;
  assign n35956 = controllable_hmaster0 & ~n35955;
  assign n35957 = ~controllable_hmaster1 & ~n35956;
  assign n35958 = ~n35954 & ~n35957;
  assign n35959 = ~i_hbusreq3 & ~n35958;
  assign n35960 = ~n35946 & ~n35959;
  assign n35961 = controllable_hmaster2 & ~n35960;
  assign n35962 = controllable_hmaster2 & ~n35961;
  assign n35963 = ~controllable_hgrant3 & ~n35962;
  assign n35964 = ~n3409 & ~n35963;
  assign n35965 = controllable_nhgrant0 & ~n35964;
  assign n35966 = ~n3466 & ~n35965;
  assign n35967 = ~n3281 & ~n35966;
  assign n35968 = ~n3281 & ~n35967;
  assign n35969 = n3378 & ~n35968;
  assign n35970 = ~n5041 & ~n35937;
  assign n35971 = ~controllable_hgrant2 & ~n35970;
  assign n35972 = ~n3410 & ~n35971;
  assign n35973 = controllable_hmaster1 & ~n35972;
  assign n35974 = controllable_hmaster0 & ~n35972;
  assign n35975 = controllable_hmaster0 & ~n35974;
  assign n35976 = ~controllable_hmaster1 & ~n35975;
  assign n35977 = ~n35973 & ~n35976;
  assign n35978 = i_hbusreq3 & ~n35977;
  assign n35979 = i_hbusreq2 & ~n35970;
  assign n35980 = controllable_hgrant4 & ~n16026;
  assign n35981 = ~n5064 & ~n35980;
  assign n35982 = ~i_hbusreq2 & ~n35981;
  assign n35983 = ~n35979 & ~n35982;
  assign n35984 = ~controllable_hgrant2 & ~n35983;
  assign n35985 = ~n3859 & ~n35984;
  assign n35986 = controllable_hmaster1 & ~n35985;
  assign n35987 = controllable_hmaster0 & ~n35985;
  assign n35988 = controllable_hmaster0 & ~n35987;
  assign n35989 = ~controllable_hmaster1 & ~n35988;
  assign n35990 = ~n35986 & ~n35989;
  assign n35991 = ~i_hbusreq3 & ~n35990;
  assign n35992 = ~n35978 & ~n35991;
  assign n35993 = controllable_hmaster2 & ~n35992;
  assign n35994 = controllable_hmaster2 & ~n35993;
  assign n35995 = ~controllable_hgrant3 & ~n35994;
  assign n35996 = ~n7090 & ~n35995;
  assign n35997 = controllable_nhgrant0 & ~n35996;
  assign n35998 = ~n7118 & ~n35997;
  assign n35999 = ~n3281 & ~n35998;
  assign n36000 = ~n3281 & ~n35999;
  assign n36001 = ~n3378 & ~n36000;
  assign n36002 = ~n35969 & ~n36001;
  assign n36003 = n3492 & ~n36002;
  assign n36004 = n3492 & ~n36003;
  assign n36005 = n3485 & ~n36004;
  assign n36006 = n3485 & ~n36005;
  assign n36007 = ~n3374 & ~n36006;
  assign n36008 = ~n34637 & ~n35942;
  assign n36009 = ~controllable_hmaster1 & ~n36008;
  assign n36010 = ~n35941 & ~n36009;
  assign n36011 = i_hbusreq3 & ~n36010;
  assign n36012 = ~n34649 & ~n35955;
  assign n36013 = ~controllable_hmaster1 & ~n36012;
  assign n36014 = ~n35954 & ~n36013;
  assign n36015 = ~i_hbusreq3 & ~n36014;
  assign n36016 = ~n36011 & ~n36015;
  assign n36017 = controllable_hmaster2 & ~n36016;
  assign n36018 = ~n12042 & ~n35937;
  assign n36019 = ~controllable_hgrant2 & ~n36018;
  assign n36020 = ~n3410 & ~n36019;
  assign n36021 = controllable_hmaster0 & ~n36020;
  assign n36022 = ~n5288 & ~n36019;
  assign n36023 = ~controllable_hmaster0 & ~n36022;
  assign n36024 = ~n36021 & ~n36023;
  assign n36025 = controllable_hmaster1 & ~n36024;
  assign n36026 = ~n5299 & ~n35937;
  assign n36027 = ~controllable_hgrant2 & ~n36026;
  assign n36028 = ~n3410 & ~n36027;
  assign n36029 = controllable_hmaster0 & ~n36028;
  assign n36030 = ~controllable_hmaster0 & ~n36020;
  assign n36031 = ~n36029 & ~n36030;
  assign n36032 = ~controllable_hmaster1 & ~n36031;
  assign n36033 = ~n36025 & ~n36032;
  assign n36034 = i_hbusreq3 & ~n36033;
  assign n36035 = i_hbusreq2 & ~n36018;
  assign n36036 = ~n12053 & ~n35948;
  assign n36037 = ~i_hbusreq2 & ~n36036;
  assign n36038 = ~n36035 & ~n36037;
  assign n36039 = ~controllable_hgrant2 & ~n36038;
  assign n36040 = ~n3431 & ~n36039;
  assign n36041 = controllable_hmaster0 & ~n36040;
  assign n36042 = ~n5308 & ~n36039;
  assign n36043 = ~controllable_hmaster0 & ~n36042;
  assign n36044 = ~n36041 & ~n36043;
  assign n36045 = controllable_hmaster1 & ~n36044;
  assign n36046 = i_hbusreq2 & ~n36026;
  assign n36047 = ~n5326 & ~n35948;
  assign n36048 = ~i_hbusreq2 & ~n36047;
  assign n36049 = ~n36046 & ~n36048;
  assign n36050 = ~controllable_hgrant2 & ~n36049;
  assign n36051 = ~n3431 & ~n36050;
  assign n36052 = controllable_hmaster0 & ~n36051;
  assign n36053 = ~controllable_hmaster0 & ~n36040;
  assign n36054 = ~n36052 & ~n36053;
  assign n36055 = ~controllable_hmaster1 & ~n36054;
  assign n36056 = ~n36045 & ~n36055;
  assign n36057 = ~i_hbusreq3 & ~n36056;
  assign n36058 = ~n36034 & ~n36057;
  assign n36059 = ~controllable_hmaster2 & ~n36058;
  assign n36060 = ~n36017 & ~n36059;
  assign n36061 = ~controllable_hgrant3 & ~n36060;
  assign n36062 = ~n7136 & ~n36061;
  assign n36063 = controllable_nhgrant0 & ~n36062;
  assign n36064 = ~n7166 & ~n36063;
  assign n36065 = ~n3281 & ~n36064;
  assign n36066 = ~n3281 & ~n36065;
  assign n36067 = n3378 & ~n36066;
  assign n36068 = ~n34637 & ~n35974;
  assign n36069 = ~controllable_hmaster1 & ~n36068;
  assign n36070 = ~n35973 & ~n36069;
  assign n36071 = i_hbusreq3 & ~n36070;
  assign n36072 = ~n34649 & ~n35987;
  assign n36073 = ~controllable_hmaster1 & ~n36072;
  assign n36074 = ~n35986 & ~n36073;
  assign n36075 = ~i_hbusreq3 & ~n36074;
  assign n36076 = ~n36071 & ~n36075;
  assign n36077 = controllable_hmaster2 & ~n36076;
  assign n36078 = ~n3906 & ~n35937;
  assign n36079 = ~controllable_hgrant2 & ~n36078;
  assign n36080 = ~n3410 & ~n36079;
  assign n36081 = controllable_hmaster0 & ~n36080;
  assign n36082 = ~n5288 & ~n36079;
  assign n36083 = ~controllable_hmaster0 & ~n36082;
  assign n36084 = ~n36081 & ~n36083;
  assign n36085 = controllable_hmaster1 & ~n36084;
  assign n36086 = ~n5429 & ~n35937;
  assign n36087 = ~controllable_hgrant2 & ~n36086;
  assign n36088 = ~n3410 & ~n36087;
  assign n36089 = controllable_hmaster0 & ~n36088;
  assign n36090 = ~controllable_hmaster0 & ~n36080;
  assign n36091 = ~n36089 & ~n36090;
  assign n36092 = ~controllable_hmaster1 & ~n36091;
  assign n36093 = ~n36085 & ~n36092;
  assign n36094 = i_hbusreq3 & ~n36093;
  assign n36095 = i_hbusreq2 & ~n36078;
  assign n36096 = ~n3929 & ~n35980;
  assign n36097 = ~i_hbusreq2 & ~n36096;
  assign n36098 = ~n36095 & ~n36097;
  assign n36099 = ~controllable_hgrant2 & ~n36098;
  assign n36100 = ~n3859 & ~n36099;
  assign n36101 = controllable_hmaster0 & ~n36100;
  assign n36102 = ~n5438 & ~n36099;
  assign n36103 = ~controllable_hmaster0 & ~n36102;
  assign n36104 = ~n36101 & ~n36103;
  assign n36105 = controllable_hmaster1 & ~n36104;
  assign n36106 = i_hbusreq2 & ~n36086;
  assign n36107 = ~n5454 & ~n35980;
  assign n36108 = ~i_hbusreq2 & ~n36107;
  assign n36109 = ~n36106 & ~n36108;
  assign n36110 = ~controllable_hgrant2 & ~n36109;
  assign n36111 = ~n3859 & ~n36110;
  assign n36112 = controllable_hmaster0 & ~n36111;
  assign n36113 = controllable_hgrant4 & ~n16140;
  assign n36114 = ~n5472 & ~n36113;
  assign n36115 = ~i_hbusreq2 & ~n36114;
  assign n36116 = ~n36095 & ~n36115;
  assign n36117 = ~controllable_hgrant2 & ~n36116;
  assign n36118 = ~n5461 & ~n36117;
  assign n36119 = ~controllable_hmaster0 & ~n36118;
  assign n36120 = ~n36112 & ~n36119;
  assign n36121 = ~controllable_hmaster1 & ~n36120;
  assign n36122 = ~n36105 & ~n36121;
  assign n36123 = ~i_hbusreq3 & ~n36122;
  assign n36124 = ~n36094 & ~n36123;
  assign n36125 = ~controllable_hmaster2 & ~n36124;
  assign n36126 = ~n36077 & ~n36125;
  assign n36127 = ~controllable_hgrant3 & ~n36126;
  assign n36128 = ~n7178 & ~n36127;
  assign n36129 = controllable_nhgrant0 & ~n36128;
  assign n36130 = ~n7208 & ~n36129;
  assign n36131 = ~n3281 & ~n36130;
  assign n36132 = ~n3281 & ~n36131;
  assign n36133 = ~n3378 & ~n36132;
  assign n36134 = ~n36067 & ~n36133;
  assign n36135 = n3492 & ~n36134;
  assign n36136 = n3492 & ~n36135;
  assign n36137 = n3485 & ~n36136;
  assign n36138 = n3485 & ~n36137;
  assign n36139 = ~n3476 & ~n36138;
  assign n36140 = i_hlock4 & ~n9968;
  assign n36141 = ~i_hlock4 & ~n9970;
  assign n36142 = ~n36140 & ~n36141;
  assign n36143 = controllable_hgrant4 & ~n36142;
  assign n36144 = ~n7245 & ~n36143;
  assign n36145 = ~controllable_hgrant2 & ~n36144;
  assign n36146 = ~n5616 & ~n36145;
  assign n36147 = controllable_hmaster1 & ~n36146;
  assign n36148 = controllable_hmaster0 & ~n36146;
  assign n36149 = ~n7255 & ~n34682;
  assign n36150 = ~controllable_hgrant2 & ~n36149;
  assign n36151 = ~n5616 & ~n36150;
  assign n36152 = ~controllable_hmaster0 & ~n36151;
  assign n36153 = ~n36148 & ~n36152;
  assign n36154 = ~controllable_hmaster1 & ~n36153;
  assign n36155 = ~n36147 & ~n36154;
  assign n36156 = i_hbusreq3 & ~n36155;
  assign n36157 = i_hbusreq2 & ~n36144;
  assign n36158 = i_hbusreq4 & ~n36142;
  assign n36159 = i_hlock4 & ~n16179;
  assign n36160 = ~i_hlock4 & ~n16187;
  assign n36161 = ~n36159 & ~n36160;
  assign n36162 = ~i_hbusreq4 & ~n36161;
  assign n36163 = ~n36158 & ~n36162;
  assign n36164 = controllable_hgrant4 & ~n36163;
  assign n36165 = ~n7282 & ~n36164;
  assign n36166 = ~i_hbusreq2 & ~n36165;
  assign n36167 = ~n36157 & ~n36166;
  assign n36168 = ~controllable_hgrant2 & ~n36167;
  assign n36169 = ~n5635 & ~n36168;
  assign n36170 = controllable_hmaster1 & ~n36169;
  assign n36171 = controllable_hmaster0 & ~n36169;
  assign n36172 = i_hbusreq2 & ~n36149;
  assign n36173 = ~n7308 & ~n34712;
  assign n36174 = ~i_hbusreq2 & ~n36173;
  assign n36175 = ~n36172 & ~n36174;
  assign n36176 = ~controllable_hgrant2 & ~n36175;
  assign n36177 = ~n7290 & ~n36176;
  assign n36178 = ~controllable_hmaster0 & ~n36177;
  assign n36179 = ~n36171 & ~n36178;
  assign n36180 = ~controllable_hmaster1 & ~n36179;
  assign n36181 = ~n36170 & ~n36180;
  assign n36182 = ~i_hbusreq3 & ~n36181;
  assign n36183 = ~n36156 & ~n36182;
  assign n36184 = controllable_hmaster2 & ~n36183;
  assign n36185 = ~n7322 & ~n36143;
  assign n36186 = ~controllable_hgrant2 & ~n36185;
  assign n36187 = ~n5616 & ~n36186;
  assign n36188 = controllable_hmaster0 & ~n36187;
  assign n36189 = ~n5686 & ~n36186;
  assign n36190 = ~controllable_hmaster0 & ~n36189;
  assign n36191 = ~n36188 & ~n36190;
  assign n36192 = controllable_hmaster1 & ~n36191;
  assign n36193 = ~n7335 & ~n36143;
  assign n36194 = ~controllable_hgrant2 & ~n36193;
  assign n36195 = ~n5616 & ~n36194;
  assign n36196 = controllable_hmaster0 & ~n36195;
  assign n36197 = ~controllable_hmaster0 & ~n36187;
  assign n36198 = ~n36196 & ~n36197;
  assign n36199 = ~controllable_hmaster1 & ~n36198;
  assign n36200 = ~n36192 & ~n36199;
  assign n36201 = i_hbusreq3 & ~n36200;
  assign n36202 = i_hbusreq2 & ~n36185;
  assign n36203 = ~n7353 & ~n36164;
  assign n36204 = ~i_hbusreq2 & ~n36203;
  assign n36205 = ~n36202 & ~n36204;
  assign n36206 = ~controllable_hgrant2 & ~n36205;
  assign n36207 = ~n5635 & ~n36206;
  assign n36208 = controllable_hmaster0 & ~n36207;
  assign n36209 = ~n5722 & ~n36206;
  assign n36210 = ~controllable_hmaster0 & ~n36209;
  assign n36211 = ~n36208 & ~n36210;
  assign n36212 = controllable_hmaster1 & ~n36211;
  assign n36213 = i_hbusreq2 & ~n36193;
  assign n36214 = ~n7376 & ~n36164;
  assign n36215 = ~i_hbusreq2 & ~n36214;
  assign n36216 = ~n36213 & ~n36215;
  assign n36217 = ~controllable_hgrant2 & ~n36216;
  assign n36218 = ~n5635 & ~n36217;
  assign n36219 = controllable_hmaster0 & ~n36218;
  assign n36220 = ~controllable_hmaster0 & ~n36207;
  assign n36221 = ~n36219 & ~n36220;
  assign n36222 = ~controllable_hmaster1 & ~n36221;
  assign n36223 = ~n36212 & ~n36222;
  assign n36224 = ~i_hbusreq3 & ~n36223;
  assign n36225 = ~n36201 & ~n36224;
  assign n36226 = ~controllable_hmaster2 & ~n36225;
  assign n36227 = ~n36184 & ~n36226;
  assign n36228 = ~controllable_hgrant3 & ~n36227;
  assign n36229 = ~n7240 & ~n36228;
  assign n36230 = controllable_nhgrant0 & ~n36229;
  assign n36231 = ~n7432 & ~n36230;
  assign n36232 = ~n3281 & ~n36231;
  assign n36233 = ~n3281 & ~n36232;
  assign n36234 = n3378 & ~n36233;
  assign n36235 = ~n7461 & ~n36143;
  assign n36236 = ~controllable_hgrant2 & ~n36235;
  assign n36237 = ~n5616 & ~n36236;
  assign n36238 = controllable_hmaster1 & ~n36237;
  assign n36239 = controllable_hmaster0 & ~n36237;
  assign n36240 = ~n7470 & ~n34682;
  assign n36241 = ~controllable_hgrant2 & ~n36240;
  assign n36242 = ~n5616 & ~n36241;
  assign n36243 = ~controllable_hmaster0 & ~n36242;
  assign n36244 = ~n36239 & ~n36243;
  assign n36245 = ~controllable_hmaster1 & ~n36244;
  assign n36246 = ~n36238 & ~n36245;
  assign n36247 = i_hbusreq3 & ~n36246;
  assign n36248 = i_hbusreq2 & ~n36235;
  assign n36249 = i_hlock4 & ~n16256;
  assign n36250 = ~i_hlock4 & ~n16265;
  assign n36251 = ~n36249 & ~n36250;
  assign n36252 = ~i_hbusreq4 & ~n36251;
  assign n36253 = ~n36158 & ~n36252;
  assign n36254 = controllable_hgrant4 & ~n36253;
  assign n36255 = ~n7499 & ~n36254;
  assign n36256 = ~i_hbusreq2 & ~n36255;
  assign n36257 = ~n36248 & ~n36256;
  assign n36258 = ~controllable_hgrant2 & ~n36257;
  assign n36259 = ~n5862 & ~n36258;
  assign n36260 = controllable_hmaster1 & ~n36259;
  assign n36261 = controllable_hmaster0 & ~n36259;
  assign n36262 = i_hbusreq2 & ~n36240;
  assign n36263 = ~n7521 & ~n34712;
  assign n36264 = ~i_hbusreq2 & ~n36263;
  assign n36265 = ~n36262 & ~n36264;
  assign n36266 = ~controllable_hgrant2 & ~n36265;
  assign n36267 = ~n7507 & ~n36266;
  assign n36268 = ~controllable_hmaster0 & ~n36267;
  assign n36269 = ~n36261 & ~n36268;
  assign n36270 = ~controllable_hmaster1 & ~n36269;
  assign n36271 = ~n36260 & ~n36270;
  assign n36272 = ~i_hbusreq3 & ~n36271;
  assign n36273 = ~n36247 & ~n36272;
  assign n36274 = controllable_hmaster2 & ~n36273;
  assign n36275 = ~n7535 & ~n36143;
  assign n36276 = ~controllable_hgrant2 & ~n36275;
  assign n36277 = ~n5616 & ~n36276;
  assign n36278 = controllable_hmaster0 & ~n36277;
  assign n36279 = ~n5686 & ~n36276;
  assign n36280 = ~controllable_hmaster0 & ~n36279;
  assign n36281 = ~n36278 & ~n36280;
  assign n36282 = controllable_hmaster1 & ~n36281;
  assign n36283 = ~n7547 & ~n36143;
  assign n36284 = ~controllable_hgrant2 & ~n36283;
  assign n36285 = ~n5616 & ~n36284;
  assign n36286 = controllable_hmaster0 & ~n36285;
  assign n36287 = ~controllable_hmaster0 & ~n36277;
  assign n36288 = ~n36286 & ~n36287;
  assign n36289 = ~controllable_hmaster1 & ~n36288;
  assign n36290 = ~n36282 & ~n36289;
  assign n36291 = i_hbusreq3 & ~n36290;
  assign n36292 = i_hbusreq2 & ~n36275;
  assign n36293 = ~n7568 & ~n36254;
  assign n36294 = ~i_hbusreq2 & ~n36293;
  assign n36295 = ~n36292 & ~n36294;
  assign n36296 = ~controllable_hgrant2 & ~n36295;
  assign n36297 = ~n5862 & ~n36296;
  assign n36298 = controllable_hmaster0 & ~n36297;
  assign n36299 = ~n5950 & ~n36296;
  assign n36300 = ~controllable_hmaster0 & ~n36299;
  assign n36301 = ~n36298 & ~n36300;
  assign n36302 = controllable_hmaster1 & ~n36301;
  assign n36303 = i_hbusreq2 & ~n36283;
  assign n36304 = ~n7592 & ~n36254;
  assign n36305 = ~i_hbusreq2 & ~n36304;
  assign n36306 = ~n36303 & ~n36305;
  assign n36307 = ~controllable_hgrant2 & ~n36306;
  assign n36308 = ~n5862 & ~n36307;
  assign n36309 = controllable_hmaster0 & ~n36308;
  assign n36310 = i_hlock4 & ~n16311;
  assign n36311 = ~i_hlock4 & ~n16321;
  assign n36312 = ~n36310 & ~n36311;
  assign n36313 = ~i_hbusreq4 & ~n36312;
  assign n36314 = ~n36158 & ~n36313;
  assign n36315 = controllable_hgrant4 & ~n36314;
  assign n36316 = ~n7614 & ~n36315;
  assign n36317 = ~i_hbusreq2 & ~n36316;
  assign n36318 = ~n36292 & ~n36317;
  assign n36319 = ~controllable_hgrant2 & ~n36318;
  assign n36320 = ~n5981 & ~n36319;
  assign n36321 = ~controllable_hmaster0 & ~n36320;
  assign n36322 = ~n36309 & ~n36321;
  assign n36323 = ~controllable_hmaster1 & ~n36322;
  assign n36324 = ~n36302 & ~n36323;
  assign n36325 = ~i_hbusreq3 & ~n36324;
  assign n36326 = ~n36291 & ~n36325;
  assign n36327 = ~controllable_hmaster2 & ~n36326;
  assign n36328 = ~n36274 & ~n36327;
  assign n36329 = ~controllable_hgrant3 & ~n36328;
  assign n36330 = ~n7457 & ~n36329;
  assign n36331 = controllable_nhgrant0 & ~n36330;
  assign n36332 = ~n7668 & ~n36331;
  assign n36333 = ~n3281 & ~n36332;
  assign n36334 = ~n3281 & ~n36333;
  assign n36335 = ~n3378 & ~n36334;
  assign n36336 = ~n36234 & ~n36335;
  assign n36337 = n3492 & ~n36336;
  assign n36338 = ~n34669 & ~n36337;
  assign n36339 = n3485 & ~n36338;
  assign n36340 = ~n34668 & ~n36339;
  assign n36341 = n3476 & ~n36340;
  assign n36342 = ~n36139 & ~n36341;
  assign n36343 = n3374 & ~n36342;
  assign n36344 = ~n36007 & ~n36343;
  assign n36345 = n3655 & ~n36344;
  assign n36346 = ~n6100 & ~n35937;
  assign n36347 = ~controllable_hgrant2 & ~n36346;
  assign n36348 = ~n3410 & ~n36347;
  assign n36349 = controllable_hmaster1 & ~n36348;
  assign n36350 = controllable_hmaster0 & ~n36348;
  assign n36351 = controllable_hmaster0 & ~n36350;
  assign n36352 = ~controllable_hmaster1 & ~n36351;
  assign n36353 = ~n36349 & ~n36352;
  assign n36354 = i_hbusreq3 & ~n36353;
  assign n36355 = i_hbusreq2 & ~n36346;
  assign n36356 = ~n6123 & ~n35980;
  assign n36357 = ~i_hbusreq2 & ~n36356;
  assign n36358 = ~n36355 & ~n36357;
  assign n36359 = ~controllable_hgrant2 & ~n36358;
  assign n36360 = ~n3859 & ~n36359;
  assign n36361 = controllable_hmaster1 & ~n36360;
  assign n36362 = controllable_hmaster0 & ~n36360;
  assign n36363 = controllable_hmaster0 & ~n36362;
  assign n36364 = ~controllable_hmaster1 & ~n36363;
  assign n36365 = ~n36361 & ~n36364;
  assign n36366 = ~i_hbusreq3 & ~n36365;
  assign n36367 = ~n36354 & ~n36366;
  assign n36368 = controllable_hmaster2 & ~n36367;
  assign n36369 = controllable_hmaster2 & ~n36368;
  assign n36370 = ~controllable_hgrant3 & ~n36369;
  assign n36371 = ~n7090 & ~n36370;
  assign n36372 = controllable_nhgrant0 & ~n36371;
  assign n36373 = ~n7118 & ~n36372;
  assign n36374 = ~n3281 & ~n36373;
  assign n36375 = ~n3281 & ~n36374;
  assign n36376 = ~n3378 & ~n36375;
  assign n36377 = ~n35969 & ~n36376;
  assign n36378 = n3492 & ~n36377;
  assign n36379 = n3492 & ~n36378;
  assign n36380 = n3485 & ~n36379;
  assign n36381 = n3485 & ~n36380;
  assign n36382 = ~n3374 & ~n36381;
  assign n36383 = ~n34748 & ~n35942;
  assign n36384 = ~controllable_hmaster1 & ~n36383;
  assign n36385 = ~n35941 & ~n36384;
  assign n36386 = i_hbusreq3 & ~n36385;
  assign n36387 = ~n34759 & ~n35955;
  assign n36388 = ~controllable_hmaster1 & ~n36387;
  assign n36389 = ~n35954 & ~n36388;
  assign n36390 = ~i_hbusreq3 & ~n36389;
  assign n36391 = ~n36386 & ~n36390;
  assign n36392 = controllable_hmaster2 & ~n36391;
  assign n36393 = ~n36059 & ~n36392;
  assign n36394 = ~controllable_hgrant3 & ~n36393;
  assign n36395 = ~n7136 & ~n36394;
  assign n36396 = controllable_nhgrant0 & ~n36395;
  assign n36397 = ~n7166 & ~n36396;
  assign n36398 = ~n3281 & ~n36397;
  assign n36399 = ~n3281 & ~n36398;
  assign n36400 = n3378 & ~n36399;
  assign n36401 = ~n34748 & ~n36350;
  assign n36402 = ~controllable_hmaster1 & ~n36401;
  assign n36403 = ~n36349 & ~n36402;
  assign n36404 = i_hbusreq3 & ~n36403;
  assign n36405 = ~n34759 & ~n36362;
  assign n36406 = ~controllable_hmaster1 & ~n36405;
  assign n36407 = ~n36361 & ~n36406;
  assign n36408 = ~i_hbusreq3 & ~n36407;
  assign n36409 = ~n36404 & ~n36408;
  assign n36410 = controllable_hmaster2 & ~n36409;
  assign n36411 = ~n6250 & ~n35937;
  assign n36412 = ~controllable_hgrant2 & ~n36411;
  assign n36413 = ~n3410 & ~n36412;
  assign n36414 = controllable_hmaster0 & ~n36413;
  assign n36415 = ~n5288 & ~n36412;
  assign n36416 = ~controllable_hmaster0 & ~n36415;
  assign n36417 = ~n36414 & ~n36416;
  assign n36418 = controllable_hmaster1 & ~n36417;
  assign n36419 = ~n6264 & ~n35937;
  assign n36420 = ~controllable_hgrant2 & ~n36419;
  assign n36421 = ~n3410 & ~n36420;
  assign n36422 = controllable_hmaster0 & ~n36421;
  assign n36423 = ~controllable_hmaster0 & ~n36413;
  assign n36424 = ~n36422 & ~n36423;
  assign n36425 = ~controllable_hmaster1 & ~n36424;
  assign n36426 = ~n36418 & ~n36425;
  assign n36427 = i_hbusreq3 & ~n36426;
  assign n36428 = i_hbusreq2 & ~n36411;
  assign n36429 = ~n6287 & ~n35980;
  assign n36430 = ~i_hbusreq2 & ~n36429;
  assign n36431 = ~n36428 & ~n36430;
  assign n36432 = ~controllable_hgrant2 & ~n36431;
  assign n36433 = ~n3859 & ~n36432;
  assign n36434 = controllable_hmaster0 & ~n36433;
  assign n36435 = ~n5438 & ~n36432;
  assign n36436 = ~controllable_hmaster0 & ~n36435;
  assign n36437 = ~n36434 & ~n36436;
  assign n36438 = controllable_hmaster1 & ~n36437;
  assign n36439 = i_hbusreq2 & ~n36419;
  assign n36440 = ~n6315 & ~n35980;
  assign n36441 = ~i_hbusreq2 & ~n36440;
  assign n36442 = ~n36439 & ~n36441;
  assign n36443 = ~controllable_hgrant2 & ~n36442;
  assign n36444 = ~n3859 & ~n36443;
  assign n36445 = controllable_hmaster0 & ~n36444;
  assign n36446 = ~n6331 & ~n36113;
  assign n36447 = ~i_hbusreq2 & ~n36446;
  assign n36448 = ~n36428 & ~n36447;
  assign n36449 = ~controllable_hgrant2 & ~n36448;
  assign n36450 = ~n5461 & ~n36449;
  assign n36451 = ~controllable_hmaster0 & ~n36450;
  assign n36452 = ~n36445 & ~n36451;
  assign n36453 = ~controllable_hmaster1 & ~n36452;
  assign n36454 = ~n36438 & ~n36453;
  assign n36455 = ~i_hbusreq3 & ~n36454;
  assign n36456 = ~n36427 & ~n36455;
  assign n36457 = ~controllable_hmaster2 & ~n36456;
  assign n36458 = ~n36410 & ~n36457;
  assign n36459 = ~controllable_hgrant3 & ~n36458;
  assign n36460 = ~n7178 & ~n36459;
  assign n36461 = controllable_nhgrant0 & ~n36460;
  assign n36462 = ~n7208 & ~n36461;
  assign n36463 = ~n3281 & ~n36462;
  assign n36464 = ~n3281 & ~n36463;
  assign n36465 = ~n3378 & ~n36464;
  assign n36466 = ~n36400 & ~n36465;
  assign n36467 = n3492 & ~n36466;
  assign n36468 = n3492 & ~n36467;
  assign n36469 = n3485 & ~n36468;
  assign n36470 = n3485 & ~n36469;
  assign n36471 = ~n3476 & ~n36470;
  assign n36472 = ~n7750 & ~n34682;
  assign n36473 = ~controllable_hgrant2 & ~n36472;
  assign n36474 = ~n5616 & ~n36473;
  assign n36475 = ~controllable_hmaster0 & ~n36474;
  assign n36476 = ~n36148 & ~n36475;
  assign n36477 = ~controllable_hmaster1 & ~n36476;
  assign n36478 = ~n36147 & ~n36477;
  assign n36479 = i_hbusreq3 & ~n36478;
  assign n36480 = i_hbusreq2 & ~n36472;
  assign n36481 = ~n7771 & ~n34712;
  assign n36482 = ~i_hbusreq2 & ~n36481;
  assign n36483 = ~n36480 & ~n36482;
  assign n36484 = ~controllable_hgrant2 & ~n36483;
  assign n36485 = ~n7290 & ~n36484;
  assign n36486 = ~controllable_hmaster0 & ~n36485;
  assign n36487 = ~n36171 & ~n36486;
  assign n36488 = ~controllable_hmaster1 & ~n36487;
  assign n36489 = ~n36170 & ~n36488;
  assign n36490 = ~i_hbusreq3 & ~n36489;
  assign n36491 = ~n36479 & ~n36490;
  assign n36492 = controllable_hmaster2 & ~n36491;
  assign n36493 = ~n36226 & ~n36492;
  assign n36494 = ~controllable_hgrant3 & ~n36493;
  assign n36495 = ~n7240 & ~n36494;
  assign n36496 = controllable_nhgrant0 & ~n36495;
  assign n36497 = ~n7432 & ~n36496;
  assign n36498 = ~n3281 & ~n36497;
  assign n36499 = ~n3281 & ~n36498;
  assign n36500 = n3378 & ~n36499;
  assign n36501 = ~n7794 & ~n36143;
  assign n36502 = ~controllable_hgrant2 & ~n36501;
  assign n36503 = ~n5616 & ~n36502;
  assign n36504 = controllable_hmaster1 & ~n36503;
  assign n36505 = controllable_hmaster0 & ~n36503;
  assign n36506 = ~n7802 & ~n34682;
  assign n36507 = ~controllable_hgrant2 & ~n36506;
  assign n36508 = ~n5616 & ~n36507;
  assign n36509 = ~controllable_hmaster0 & ~n36508;
  assign n36510 = ~n36505 & ~n36509;
  assign n36511 = ~controllable_hmaster1 & ~n36510;
  assign n36512 = ~n36504 & ~n36511;
  assign n36513 = i_hbusreq3 & ~n36512;
  assign n36514 = i_hbusreq2 & ~n36501;
  assign n36515 = ~n7824 & ~n36254;
  assign n36516 = ~i_hbusreq2 & ~n36515;
  assign n36517 = ~n36514 & ~n36516;
  assign n36518 = ~controllable_hgrant2 & ~n36517;
  assign n36519 = ~n5862 & ~n36518;
  assign n36520 = controllable_hmaster1 & ~n36519;
  assign n36521 = controllable_hmaster0 & ~n36519;
  assign n36522 = i_hbusreq2 & ~n36506;
  assign n36523 = ~n7845 & ~n34712;
  assign n36524 = ~i_hbusreq2 & ~n36523;
  assign n36525 = ~n36522 & ~n36524;
  assign n36526 = ~controllable_hgrant2 & ~n36525;
  assign n36527 = ~n7507 & ~n36526;
  assign n36528 = ~controllable_hmaster0 & ~n36527;
  assign n36529 = ~n36521 & ~n36528;
  assign n36530 = ~controllable_hmaster1 & ~n36529;
  assign n36531 = ~n36520 & ~n36530;
  assign n36532 = ~i_hbusreq3 & ~n36531;
  assign n36533 = ~n36513 & ~n36532;
  assign n36534 = controllable_hmaster2 & ~n36533;
  assign n36535 = ~n7859 & ~n36143;
  assign n36536 = ~controllable_hgrant2 & ~n36535;
  assign n36537 = ~n5616 & ~n36536;
  assign n36538 = controllable_hmaster0 & ~n36537;
  assign n36539 = ~n5686 & ~n36536;
  assign n36540 = ~controllable_hmaster0 & ~n36539;
  assign n36541 = ~n36538 & ~n36540;
  assign n36542 = controllable_hmaster1 & ~n36541;
  assign n36543 = ~n7870 & ~n36143;
  assign n36544 = ~controllable_hgrant2 & ~n36543;
  assign n36545 = ~n5616 & ~n36544;
  assign n36546 = controllable_hmaster0 & ~n36545;
  assign n36547 = ~controllable_hmaster0 & ~n36537;
  assign n36548 = ~n36546 & ~n36547;
  assign n36549 = ~controllable_hmaster1 & ~n36548;
  assign n36550 = ~n36542 & ~n36549;
  assign n36551 = i_hbusreq3 & ~n36550;
  assign n36552 = i_hbusreq2 & ~n36535;
  assign n36553 = ~n7891 & ~n36254;
  assign n36554 = ~i_hbusreq2 & ~n36553;
  assign n36555 = ~n36552 & ~n36554;
  assign n36556 = ~controllable_hgrant2 & ~n36555;
  assign n36557 = ~n5862 & ~n36556;
  assign n36558 = controllable_hmaster0 & ~n36557;
  assign n36559 = ~n5950 & ~n36556;
  assign n36560 = ~controllable_hmaster0 & ~n36559;
  assign n36561 = ~n36558 & ~n36560;
  assign n36562 = controllable_hmaster1 & ~n36561;
  assign n36563 = i_hbusreq2 & ~n36543;
  assign n36564 = ~n7916 & ~n36254;
  assign n36565 = ~i_hbusreq2 & ~n36564;
  assign n36566 = ~n36563 & ~n36565;
  assign n36567 = ~controllable_hgrant2 & ~n36566;
  assign n36568 = ~n5862 & ~n36567;
  assign n36569 = controllable_hmaster0 & ~n36568;
  assign n36570 = ~n7930 & ~n36315;
  assign n36571 = ~i_hbusreq2 & ~n36570;
  assign n36572 = ~n36552 & ~n36571;
  assign n36573 = ~controllable_hgrant2 & ~n36572;
  assign n36574 = ~n5981 & ~n36573;
  assign n36575 = ~controllable_hmaster0 & ~n36574;
  assign n36576 = ~n36569 & ~n36575;
  assign n36577 = ~controllable_hmaster1 & ~n36576;
  assign n36578 = ~n36562 & ~n36577;
  assign n36579 = ~i_hbusreq3 & ~n36578;
  assign n36580 = ~n36551 & ~n36579;
  assign n36581 = ~controllable_hmaster2 & ~n36580;
  assign n36582 = ~n36534 & ~n36581;
  assign n36583 = ~controllable_hgrant3 & ~n36582;
  assign n36584 = ~n7457 & ~n36583;
  assign n36585 = controllable_nhgrant0 & ~n36584;
  assign n36586 = ~n7668 & ~n36585;
  assign n36587 = ~n3281 & ~n36586;
  assign n36588 = ~n3281 & ~n36587;
  assign n36589 = ~n3378 & ~n36588;
  assign n36590 = ~n36500 & ~n36589;
  assign n36591 = n3492 & ~n36590;
  assign n36592 = ~n34669 & ~n36591;
  assign n36593 = n3485 & ~n36592;
  assign n36594 = ~n34668 & ~n36593;
  assign n36595 = n3476 & ~n36594;
  assign n36596 = ~n36471 & ~n36595;
  assign n36597 = n3374 & ~n36596;
  assign n36598 = ~n36382 & ~n36597;
  assign n36599 = ~n3655 & ~n36598;
  assign n36600 = ~n36345 & ~n36599;
  assign n36601 = n3652 & ~n36600;
  assign n36602 = ~n4333 & ~n35971;
  assign n36603 = controllable_hmaster1 & ~n36602;
  assign n36604 = controllable_hmaster0 & ~n36602;
  assign n36605 = controllable_hmaster0 & ~n36604;
  assign n36606 = ~controllable_hmaster1 & ~n36605;
  assign n36607 = ~n36603 & ~n36606;
  assign n36608 = i_hbusreq3 & ~n36607;
  assign n36609 = ~n4340 & ~n35984;
  assign n36610 = controllable_hmaster1 & ~n36609;
  assign n36611 = controllable_hmaster0 & ~n36609;
  assign n36612 = controllable_hmaster0 & ~n36611;
  assign n36613 = ~controllable_hmaster1 & ~n36612;
  assign n36614 = ~n36610 & ~n36613;
  assign n36615 = ~i_hbusreq3 & ~n36614;
  assign n36616 = ~n36608 & ~n36615;
  assign n36617 = controllable_hmaster2 & ~n36616;
  assign n36618 = controllable_hmaster2 & ~n36617;
  assign n36619 = ~controllable_hgrant3 & ~n36618;
  assign n36620 = ~n7090 & ~n36619;
  assign n36621 = controllable_nhgrant0 & ~n36620;
  assign n36622 = ~n7118 & ~n36621;
  assign n36623 = ~n3281 & ~n36622;
  assign n36624 = ~n3281 & ~n36623;
  assign n36625 = ~n3378 & ~n36624;
  assign n36626 = ~n35969 & ~n36625;
  assign n36627 = n3492 & ~n36626;
  assign n36628 = n3492 & ~n36627;
  assign n36629 = n3485 & ~n36628;
  assign n36630 = n3485 & ~n36629;
  assign n36631 = ~n3374 & ~n36630;
  assign n36632 = ~n34818 & ~n35942;
  assign n36633 = ~controllable_hmaster1 & ~n36632;
  assign n36634 = ~n35941 & ~n36633;
  assign n36635 = i_hbusreq3 & ~n36634;
  assign n36636 = ~n34824 & ~n35955;
  assign n36637 = ~controllable_hmaster1 & ~n36636;
  assign n36638 = ~n35954 & ~n36637;
  assign n36639 = ~i_hbusreq3 & ~n36638;
  assign n36640 = ~n36635 & ~n36639;
  assign n36641 = controllable_hmaster2 & ~n36640;
  assign n36642 = ~n36059 & ~n36641;
  assign n36643 = ~controllable_hgrant3 & ~n36642;
  assign n36644 = ~n7136 & ~n36643;
  assign n36645 = controllable_nhgrant0 & ~n36644;
  assign n36646 = ~n7166 & ~n36645;
  assign n36647 = ~n3281 & ~n36646;
  assign n36648 = ~n3281 & ~n36647;
  assign n36649 = n3378 & ~n36648;
  assign n36650 = ~n34818 & ~n36604;
  assign n36651 = ~controllable_hmaster1 & ~n36650;
  assign n36652 = ~n36603 & ~n36651;
  assign n36653 = i_hbusreq3 & ~n36652;
  assign n36654 = ~n34824 & ~n36611;
  assign n36655 = ~controllable_hmaster1 & ~n36654;
  assign n36656 = ~n36610 & ~n36655;
  assign n36657 = ~i_hbusreq3 & ~n36656;
  assign n36658 = ~n36653 & ~n36657;
  assign n36659 = controllable_hmaster2 & ~n36658;
  assign n36660 = ~n4333 & ~n36079;
  assign n36661 = controllable_hmaster0 & ~n36660;
  assign n36662 = ~n6697 & ~n36079;
  assign n36663 = ~controllable_hmaster0 & ~n36662;
  assign n36664 = ~n36661 & ~n36663;
  assign n36665 = controllable_hmaster1 & ~n36664;
  assign n36666 = ~n4333 & ~n36087;
  assign n36667 = controllable_hmaster0 & ~n36666;
  assign n36668 = ~controllable_hmaster0 & ~n36660;
  assign n36669 = ~n36667 & ~n36668;
  assign n36670 = ~controllable_hmaster1 & ~n36669;
  assign n36671 = ~n36665 & ~n36670;
  assign n36672 = i_hbusreq3 & ~n36671;
  assign n36673 = ~n4340 & ~n36099;
  assign n36674 = controllable_hmaster0 & ~n36673;
  assign n36675 = ~n6710 & ~n36099;
  assign n36676 = ~controllable_hmaster0 & ~n36675;
  assign n36677 = ~n36674 & ~n36676;
  assign n36678 = controllable_hmaster1 & ~n36677;
  assign n36679 = ~n4340 & ~n36110;
  assign n36680 = controllable_hmaster0 & ~n36679;
  assign n36681 = ~n6947 & ~n36117;
  assign n36682 = ~controllable_hmaster0 & ~n36681;
  assign n36683 = ~n36680 & ~n36682;
  assign n36684 = ~controllable_hmaster1 & ~n36683;
  assign n36685 = ~n36678 & ~n36684;
  assign n36686 = ~i_hbusreq3 & ~n36685;
  assign n36687 = ~n36672 & ~n36686;
  assign n36688 = ~controllable_hmaster2 & ~n36687;
  assign n36689 = ~n36659 & ~n36688;
  assign n36690 = ~controllable_hgrant3 & ~n36689;
  assign n36691 = ~n7178 & ~n36690;
  assign n36692 = controllable_nhgrant0 & ~n36691;
  assign n36693 = ~n7208 & ~n36692;
  assign n36694 = ~n3281 & ~n36693;
  assign n36695 = ~n3281 & ~n36694;
  assign n36696 = ~n3378 & ~n36695;
  assign n36697 = ~n36649 & ~n36696;
  assign n36698 = n3492 & ~n36697;
  assign n36699 = n3492 & ~n36698;
  assign n36700 = n3485 & ~n36699;
  assign n36701 = n3485 & ~n36700;
  assign n36702 = ~n3476 & ~n36701;
  assign n36703 = ~n8029 & ~n36150;
  assign n36704 = ~controllable_hmaster0 & ~n36703;
  assign n36705 = ~n36148 & ~n36704;
  assign n36706 = ~controllable_hmaster1 & ~n36705;
  assign n36707 = ~n36147 & ~n36706;
  assign n36708 = i_hbusreq3 & ~n36707;
  assign n36709 = ~n8036 & ~n36176;
  assign n36710 = ~controllable_hmaster0 & ~n36709;
  assign n36711 = ~n36171 & ~n36710;
  assign n36712 = ~controllable_hmaster1 & ~n36711;
  assign n36713 = ~n36170 & ~n36712;
  assign n36714 = ~i_hbusreq3 & ~n36713;
  assign n36715 = ~n36708 & ~n36714;
  assign n36716 = controllable_hmaster2 & ~n36715;
  assign n36717 = ~n36226 & ~n36716;
  assign n36718 = ~controllable_hgrant3 & ~n36717;
  assign n36719 = ~n7240 & ~n36718;
  assign n36720 = controllable_nhgrant0 & ~n36719;
  assign n36721 = ~n7432 & ~n36720;
  assign n36722 = ~n3281 & ~n36721;
  assign n36723 = ~n3281 & ~n36722;
  assign n36724 = n3378 & ~n36723;
  assign n36725 = ~n6762 & ~n36236;
  assign n36726 = controllable_hmaster1 & ~n36725;
  assign n36727 = controllable_hmaster0 & ~n36725;
  assign n36728 = ~n8056 & ~n36241;
  assign n36729 = ~controllable_hmaster0 & ~n36728;
  assign n36730 = ~n36727 & ~n36729;
  assign n36731 = ~controllable_hmaster1 & ~n36730;
  assign n36732 = ~n36726 & ~n36731;
  assign n36733 = i_hbusreq3 & ~n36732;
  assign n36734 = ~n6772 & ~n36258;
  assign n36735 = controllable_hmaster1 & ~n36734;
  assign n36736 = controllable_hmaster0 & ~n36734;
  assign n36737 = ~n8066 & ~n36266;
  assign n36738 = ~controllable_hmaster0 & ~n36737;
  assign n36739 = ~n36736 & ~n36738;
  assign n36740 = ~controllable_hmaster1 & ~n36739;
  assign n36741 = ~n36735 & ~n36740;
  assign n36742 = ~i_hbusreq3 & ~n36741;
  assign n36743 = ~n36733 & ~n36742;
  assign n36744 = controllable_hmaster2 & ~n36743;
  assign n36745 = ~n6762 & ~n36276;
  assign n36746 = controllable_hmaster0 & ~n36745;
  assign n36747 = ~n6786 & ~n36276;
  assign n36748 = ~controllable_hmaster0 & ~n36747;
  assign n36749 = ~n36746 & ~n36748;
  assign n36750 = controllable_hmaster1 & ~n36749;
  assign n36751 = ~n6762 & ~n36284;
  assign n36752 = controllable_hmaster0 & ~n36751;
  assign n36753 = ~controllable_hmaster0 & ~n36745;
  assign n36754 = ~n36752 & ~n36753;
  assign n36755 = ~controllable_hmaster1 & ~n36754;
  assign n36756 = ~n36750 & ~n36755;
  assign n36757 = i_hbusreq3 & ~n36756;
  assign n36758 = ~n6772 & ~n36296;
  assign n36759 = controllable_hmaster0 & ~n36758;
  assign n36760 = ~n6813 & ~n36296;
  assign n36761 = ~controllable_hmaster0 & ~n36760;
  assign n36762 = ~n36759 & ~n36761;
  assign n36763 = controllable_hmaster1 & ~n36762;
  assign n36764 = ~n6772 & ~n36307;
  assign n36765 = controllable_hmaster0 & ~n36764;
  assign n36766 = ~n6831 & ~n36319;
  assign n36767 = ~controllable_hmaster0 & ~n36766;
  assign n36768 = ~n36765 & ~n36767;
  assign n36769 = ~controllable_hmaster1 & ~n36768;
  assign n36770 = ~n36763 & ~n36769;
  assign n36771 = ~i_hbusreq3 & ~n36770;
  assign n36772 = ~n36757 & ~n36771;
  assign n36773 = ~controllable_hmaster2 & ~n36772;
  assign n36774 = ~n36744 & ~n36773;
  assign n36775 = ~controllable_hgrant3 & ~n36774;
  assign n36776 = ~n7457 & ~n36775;
  assign n36777 = controllable_nhgrant0 & ~n36776;
  assign n36778 = ~n7668 & ~n36777;
  assign n36779 = ~n3281 & ~n36778;
  assign n36780 = ~n3281 & ~n36779;
  assign n36781 = ~n3378 & ~n36780;
  assign n36782 = ~n36724 & ~n36781;
  assign n36783 = n3492 & ~n36782;
  assign n36784 = ~n34669 & ~n36783;
  assign n36785 = n3485 & ~n36784;
  assign n36786 = ~n34668 & ~n36785;
  assign n36787 = n3476 & ~n36786;
  assign n36788 = ~n36702 & ~n36787;
  assign n36789 = n3374 & ~n36788;
  assign n36790 = ~n36631 & ~n36789;
  assign n36791 = n3655 & ~n36790;
  assign n36792 = ~n4333 & ~n36347;
  assign n36793 = controllable_hmaster1 & ~n36792;
  assign n36794 = controllable_hmaster0 & ~n36792;
  assign n36795 = controllable_hmaster0 & ~n36794;
  assign n36796 = ~controllable_hmaster1 & ~n36795;
  assign n36797 = ~n36793 & ~n36796;
  assign n36798 = i_hbusreq3 & ~n36797;
  assign n36799 = ~n4340 & ~n36359;
  assign n36800 = controllable_hmaster1 & ~n36799;
  assign n36801 = controllable_hmaster0 & ~n36799;
  assign n36802 = controllable_hmaster0 & ~n36801;
  assign n36803 = ~controllable_hmaster1 & ~n36802;
  assign n36804 = ~n36800 & ~n36803;
  assign n36805 = ~i_hbusreq3 & ~n36804;
  assign n36806 = ~n36798 & ~n36805;
  assign n36807 = controllable_hmaster2 & ~n36806;
  assign n36808 = controllable_hmaster2 & ~n36807;
  assign n36809 = ~controllable_hgrant3 & ~n36808;
  assign n36810 = ~n7090 & ~n36809;
  assign n36811 = controllable_nhgrant0 & ~n36810;
  assign n36812 = ~n7118 & ~n36811;
  assign n36813 = ~n3281 & ~n36812;
  assign n36814 = ~n3281 & ~n36813;
  assign n36815 = ~n3378 & ~n36814;
  assign n36816 = ~n35969 & ~n36815;
  assign n36817 = n3492 & ~n36816;
  assign n36818 = n3492 & ~n36817;
  assign n36819 = n3485 & ~n36818;
  assign n36820 = n3485 & ~n36819;
  assign n36821 = ~n3374 & ~n36820;
  assign n36822 = ~n34874 & ~n35942;
  assign n36823 = ~controllable_hmaster1 & ~n36822;
  assign n36824 = ~n35941 & ~n36823;
  assign n36825 = i_hbusreq3 & ~n36824;
  assign n36826 = ~n34880 & ~n35955;
  assign n36827 = ~controllable_hmaster1 & ~n36826;
  assign n36828 = ~n35954 & ~n36827;
  assign n36829 = ~i_hbusreq3 & ~n36828;
  assign n36830 = ~n36825 & ~n36829;
  assign n36831 = controllable_hmaster2 & ~n36830;
  assign n36832 = ~n36059 & ~n36831;
  assign n36833 = ~controllable_hgrant3 & ~n36832;
  assign n36834 = ~n7136 & ~n36833;
  assign n36835 = controllable_nhgrant0 & ~n36834;
  assign n36836 = ~n7166 & ~n36835;
  assign n36837 = ~n3281 & ~n36836;
  assign n36838 = ~n3281 & ~n36837;
  assign n36839 = n3378 & ~n36838;
  assign n36840 = ~n34874 & ~n36794;
  assign n36841 = ~controllable_hmaster1 & ~n36840;
  assign n36842 = ~n36793 & ~n36841;
  assign n36843 = i_hbusreq3 & ~n36842;
  assign n36844 = ~n34880 & ~n36801;
  assign n36845 = ~controllable_hmaster1 & ~n36844;
  assign n36846 = ~n36800 & ~n36845;
  assign n36847 = ~i_hbusreq3 & ~n36846;
  assign n36848 = ~n36843 & ~n36847;
  assign n36849 = controllable_hmaster2 & ~n36848;
  assign n36850 = ~n4333 & ~n36412;
  assign n36851 = controllable_hmaster0 & ~n36850;
  assign n36852 = ~n6697 & ~n36412;
  assign n36853 = ~controllable_hmaster0 & ~n36852;
  assign n36854 = ~n36851 & ~n36853;
  assign n36855 = controllable_hmaster1 & ~n36854;
  assign n36856 = ~n4333 & ~n36420;
  assign n36857 = controllable_hmaster0 & ~n36856;
  assign n36858 = ~controllable_hmaster0 & ~n36850;
  assign n36859 = ~n36857 & ~n36858;
  assign n36860 = ~controllable_hmaster1 & ~n36859;
  assign n36861 = ~n36855 & ~n36860;
  assign n36862 = i_hbusreq3 & ~n36861;
  assign n36863 = ~n4340 & ~n36432;
  assign n36864 = controllable_hmaster0 & ~n36863;
  assign n36865 = ~n6710 & ~n36432;
  assign n36866 = ~controllable_hmaster0 & ~n36865;
  assign n36867 = ~n36864 & ~n36866;
  assign n36868 = controllable_hmaster1 & ~n36867;
  assign n36869 = ~n4340 & ~n36443;
  assign n36870 = controllable_hmaster0 & ~n36869;
  assign n36871 = ~n6947 & ~n36449;
  assign n36872 = ~controllable_hmaster0 & ~n36871;
  assign n36873 = ~n36870 & ~n36872;
  assign n36874 = ~controllable_hmaster1 & ~n36873;
  assign n36875 = ~n36868 & ~n36874;
  assign n36876 = ~i_hbusreq3 & ~n36875;
  assign n36877 = ~n36862 & ~n36876;
  assign n36878 = ~controllable_hmaster2 & ~n36877;
  assign n36879 = ~n36849 & ~n36878;
  assign n36880 = ~controllable_hgrant3 & ~n36879;
  assign n36881 = ~n7178 & ~n36880;
  assign n36882 = controllable_nhgrant0 & ~n36881;
  assign n36883 = ~n7208 & ~n36882;
  assign n36884 = ~n3281 & ~n36883;
  assign n36885 = ~n3281 & ~n36884;
  assign n36886 = ~n3378 & ~n36885;
  assign n36887 = ~n36839 & ~n36886;
  assign n36888 = n3492 & ~n36887;
  assign n36889 = n3492 & ~n36888;
  assign n36890 = n3485 & ~n36889;
  assign n36891 = n3485 & ~n36890;
  assign n36892 = ~n3476 & ~n36891;
  assign n36893 = ~n8029 & ~n36473;
  assign n36894 = ~controllable_hmaster0 & ~n36893;
  assign n36895 = ~n36148 & ~n36894;
  assign n36896 = ~controllable_hmaster1 & ~n36895;
  assign n36897 = ~n36147 & ~n36896;
  assign n36898 = i_hbusreq3 & ~n36897;
  assign n36899 = ~n8036 & ~n36484;
  assign n36900 = ~controllable_hmaster0 & ~n36899;
  assign n36901 = ~n36171 & ~n36900;
  assign n36902 = ~controllable_hmaster1 & ~n36901;
  assign n36903 = ~n36170 & ~n36902;
  assign n36904 = ~i_hbusreq3 & ~n36903;
  assign n36905 = ~n36898 & ~n36904;
  assign n36906 = controllable_hmaster2 & ~n36905;
  assign n36907 = ~n36226 & ~n36906;
  assign n36908 = ~controllable_hgrant3 & ~n36907;
  assign n36909 = ~n7240 & ~n36908;
  assign n36910 = controllable_nhgrant0 & ~n36909;
  assign n36911 = ~n7432 & ~n36910;
  assign n36912 = ~n3281 & ~n36911;
  assign n36913 = ~n3281 & ~n36912;
  assign n36914 = n3378 & ~n36913;
  assign n36915 = ~n6762 & ~n36502;
  assign n36916 = controllable_hmaster1 & ~n36915;
  assign n36917 = controllable_hmaster0 & ~n36915;
  assign n36918 = ~n8056 & ~n36507;
  assign n36919 = ~controllable_hmaster0 & ~n36918;
  assign n36920 = ~n36917 & ~n36919;
  assign n36921 = ~controllable_hmaster1 & ~n36920;
  assign n36922 = ~n36916 & ~n36921;
  assign n36923 = i_hbusreq3 & ~n36922;
  assign n36924 = ~n6772 & ~n36518;
  assign n36925 = controllable_hmaster1 & ~n36924;
  assign n36926 = controllable_hmaster0 & ~n36924;
  assign n36927 = ~n8066 & ~n36526;
  assign n36928 = ~controllable_hmaster0 & ~n36927;
  assign n36929 = ~n36926 & ~n36928;
  assign n36930 = ~controllable_hmaster1 & ~n36929;
  assign n36931 = ~n36925 & ~n36930;
  assign n36932 = ~i_hbusreq3 & ~n36931;
  assign n36933 = ~n36923 & ~n36932;
  assign n36934 = controllable_hmaster2 & ~n36933;
  assign n36935 = ~n6762 & ~n36536;
  assign n36936 = controllable_hmaster0 & ~n36935;
  assign n36937 = ~n6786 & ~n36536;
  assign n36938 = ~controllable_hmaster0 & ~n36937;
  assign n36939 = ~n36936 & ~n36938;
  assign n36940 = controllable_hmaster1 & ~n36939;
  assign n36941 = ~n6762 & ~n36544;
  assign n36942 = controllable_hmaster0 & ~n36941;
  assign n36943 = ~controllable_hmaster0 & ~n36935;
  assign n36944 = ~n36942 & ~n36943;
  assign n36945 = ~controllable_hmaster1 & ~n36944;
  assign n36946 = ~n36940 & ~n36945;
  assign n36947 = i_hbusreq3 & ~n36946;
  assign n36948 = ~n6772 & ~n36556;
  assign n36949 = controllable_hmaster0 & ~n36948;
  assign n36950 = ~n6813 & ~n36556;
  assign n36951 = ~controllable_hmaster0 & ~n36950;
  assign n36952 = ~n36949 & ~n36951;
  assign n36953 = controllable_hmaster1 & ~n36952;
  assign n36954 = ~n6772 & ~n36567;
  assign n36955 = controllable_hmaster0 & ~n36954;
  assign n36956 = ~n6831 & ~n36573;
  assign n36957 = ~controllable_hmaster0 & ~n36956;
  assign n36958 = ~n36955 & ~n36957;
  assign n36959 = ~controllable_hmaster1 & ~n36958;
  assign n36960 = ~n36953 & ~n36959;
  assign n36961 = ~i_hbusreq3 & ~n36960;
  assign n36962 = ~n36947 & ~n36961;
  assign n36963 = ~controllable_hmaster2 & ~n36962;
  assign n36964 = ~n36934 & ~n36963;
  assign n36965 = ~controllable_hgrant3 & ~n36964;
  assign n36966 = ~n7457 & ~n36965;
  assign n36967 = controllable_nhgrant0 & ~n36966;
  assign n36968 = ~n7668 & ~n36967;
  assign n36969 = ~n3281 & ~n36968;
  assign n36970 = ~n3281 & ~n36969;
  assign n36971 = ~n3378 & ~n36970;
  assign n36972 = ~n36914 & ~n36971;
  assign n36973 = n3492 & ~n36972;
  assign n36974 = ~n34669 & ~n36973;
  assign n36975 = n3485 & ~n36974;
  assign n36976 = ~n34668 & ~n36975;
  assign n36977 = n3476 & ~n36976;
  assign n36978 = ~n36892 & ~n36977;
  assign n36979 = n3374 & ~n36978;
  assign n36980 = ~n36821 & ~n36979;
  assign n36981 = ~n3655 & ~n36980;
  assign n36982 = ~n36791 & ~n36981;
  assign n36983 = ~n3652 & ~n36982;
  assign n36984 = ~n36601 & ~n36983;
  assign n36985 = n3368 & ~n36984;
  assign n36986 = ~n35936 & ~n36985;
  assign n36987 = n3362 & ~n36986;
  assign n36988 = n3492 & ~n34970;
  assign n36989 = ~n3631 & ~n36988;
  assign n36990 = n3485 & ~n36989;
  assign n36991 = ~n3630 & ~n36990;
  assign n36992 = ~n3476 & ~n36991;
  assign n36993 = ~n3793 & ~n8291;
  assign n36994 = controllable_hgrant3 & ~n36993;
  assign n36995 = ~n8291 & ~n34103;
  assign n36996 = ~controllable_hgrant3 & ~n36995;
  assign n36997 = ~n36994 & ~n36996;
  assign n36998 = controllable_nhgrant0 & ~n36997;
  assign n36999 = ~n3793 & ~n8301;
  assign n37000 = ~controllable_hgrant3 & ~n36999;
  assign n37001 = ~n36994 & ~n37000;
  assign n37002 = ~controllable_nhgrant0 & ~n37001;
  assign n37003 = ~n36998 & ~n37002;
  assign n37004 = ~n3281 & ~n37003;
  assign n37005 = ~n3783 & ~n37004;
  assign n37006 = ~n3492 & ~n37005;
  assign n37007 = n3492 & ~n34110;
  assign n37008 = ~n37006 & ~n37007;
  assign n37009 = ~n3485 & ~n37008;
  assign n37010 = ~n34979 & ~n36988;
  assign n37011 = n3485 & ~n37010;
  assign n37012 = ~n37009 & ~n37011;
  assign n37013 = n3476 & ~n37012;
  assign n37014 = ~n36992 & ~n37013;
  assign n37015 = ~n3374 & ~n37014;
  assign n37016 = n3492 & ~n35102;
  assign n37017 = ~n3631 & ~n37016;
  assign n37018 = n3485 & ~n37017;
  assign n37019 = ~n3630 & ~n37018;
  assign n37020 = ~n3476 & ~n37019;
  assign n37021 = n3492 & ~n35271;
  assign n37022 = ~n34979 & ~n37021;
  assign n37023 = n3485 & ~n37022;
  assign n37024 = ~n37009 & ~n37023;
  assign n37025 = n3476 & ~n37024;
  assign n37026 = ~n37020 & ~n37025;
  assign n37027 = n3374 & ~n37026;
  assign n37028 = ~n37015 & ~n37027;
  assign n37029 = n3655 & ~n37028;
  assign n37030 = n3492 & ~n35312;
  assign n37031 = ~n3631 & ~n37030;
  assign n37032 = n3485 & ~n37031;
  assign n37033 = ~n3630 & ~n37032;
  assign n37034 = ~n3476 & ~n37033;
  assign n37035 = ~n3793 & ~n8341;
  assign n37036 = controllable_hgrant3 & ~n37035;
  assign n37037 = ~n8349 & ~n34103;
  assign n37038 = ~controllable_hgrant3 & ~n37037;
  assign n37039 = ~n37036 & ~n37038;
  assign n37040 = controllable_nhgrant0 & ~n37039;
  assign n37041 = ~n3793 & ~n8359;
  assign n37042 = ~controllable_hgrant3 & ~n37041;
  assign n37043 = ~n37036 & ~n37042;
  assign n37044 = ~controllable_nhgrant0 & ~n37043;
  assign n37045 = ~n37040 & ~n37044;
  assign n37046 = ~n3281 & ~n37045;
  assign n37047 = ~n3783 & ~n37046;
  assign n37048 = ~n3492 & ~n37047;
  assign n37049 = ~n37007 & ~n37048;
  assign n37050 = ~n3485 & ~n37049;
  assign n37051 = ~n34979 & ~n37030;
  assign n37052 = n3485 & ~n37051;
  assign n37053 = ~n37050 & ~n37052;
  assign n37054 = n3476 & ~n37053;
  assign n37055 = ~n37034 & ~n37054;
  assign n37056 = ~n3374 & ~n37055;
  assign n37057 = n3492 & ~n35411;
  assign n37058 = ~n3631 & ~n37057;
  assign n37059 = n3485 & ~n37058;
  assign n37060 = ~n3630 & ~n37059;
  assign n37061 = ~n3476 & ~n37060;
  assign n37062 = n3492 & ~n35535;
  assign n37063 = ~n34979 & ~n37062;
  assign n37064 = n3485 & ~n37063;
  assign n37065 = ~n37050 & ~n37064;
  assign n37066 = n3476 & ~n37065;
  assign n37067 = ~n37061 & ~n37066;
  assign n37068 = n3374 & ~n37067;
  assign n37069 = ~n37056 & ~n37068;
  assign n37070 = ~n3655 & ~n37069;
  assign n37071 = ~n37029 & ~n37070;
  assign n37072 = n3652 & ~n37071;
  assign n37073 = n3492 & ~n35571;
  assign n37074 = ~n3631 & ~n37073;
  assign n37075 = n3485 & ~n37074;
  assign n37076 = ~n3630 & ~n37075;
  assign n37077 = ~n3476 & ~n37076;
  assign n37078 = ~n3793 & ~n8404;
  assign n37079 = controllable_hgrant3 & ~n37078;
  assign n37080 = ~n8416 & ~n34103;
  assign n37081 = ~controllable_hgrant3 & ~n37080;
  assign n37082 = ~n37079 & ~n37081;
  assign n37083 = controllable_nhgrant0 & ~n37082;
  assign n37084 = ~n3793 & ~n8426;
  assign n37085 = ~controllable_hgrant3 & ~n37084;
  assign n37086 = ~n37079 & ~n37085;
  assign n37087 = ~controllable_nhgrant0 & ~n37086;
  assign n37088 = ~n37083 & ~n37087;
  assign n37089 = ~n3281 & ~n37088;
  assign n37090 = ~n3783 & ~n37089;
  assign n37091 = ~n3492 & ~n37090;
  assign n37092 = ~n37007 & ~n37091;
  assign n37093 = ~n3485 & ~n37092;
  assign n37094 = ~n34979 & ~n37073;
  assign n37095 = n3485 & ~n37094;
  assign n37096 = ~n37093 & ~n37095;
  assign n37097 = n3476 & ~n37096;
  assign n37098 = ~n37077 & ~n37097;
  assign n37099 = ~n3374 & ~n37098;
  assign n37100 = n3492 & ~n35644;
  assign n37101 = ~n3631 & ~n37100;
  assign n37102 = n3485 & ~n37101;
  assign n37103 = ~n3630 & ~n37102;
  assign n37104 = ~n3476 & ~n37103;
  assign n37105 = n3492 & ~n35729;
  assign n37106 = ~n34979 & ~n37105;
  assign n37107 = n3485 & ~n37106;
  assign n37108 = ~n37093 & ~n37107;
  assign n37109 = n3476 & ~n37108;
  assign n37110 = ~n37104 & ~n37109;
  assign n37111 = n3374 & ~n37110;
  assign n37112 = ~n37099 & ~n37111;
  assign n37113 = n3655 & ~n37112;
  assign n37114 = n3492 & ~n35763;
  assign n37115 = ~n3631 & ~n37114;
  assign n37116 = n3485 & ~n37115;
  assign n37117 = ~n3630 & ~n37116;
  assign n37118 = ~n3476 & ~n37117;
  assign n37119 = ~n3793 & ~n8465;
  assign n37120 = controllable_hgrant3 & ~n37119;
  assign n37121 = ~n8473 & ~n34103;
  assign n37122 = ~controllable_hgrant3 & ~n37121;
  assign n37123 = ~n37120 & ~n37122;
  assign n37124 = controllable_nhgrant0 & ~n37123;
  assign n37125 = ~n3793 & ~n8483;
  assign n37126 = ~controllable_hgrant3 & ~n37125;
  assign n37127 = ~n37120 & ~n37126;
  assign n37128 = ~controllable_nhgrant0 & ~n37127;
  assign n37129 = ~n37124 & ~n37128;
  assign n37130 = ~n3281 & ~n37129;
  assign n37131 = ~n3783 & ~n37130;
  assign n37132 = ~n3492 & ~n37131;
  assign n37133 = ~n37007 & ~n37132;
  assign n37134 = ~n3485 & ~n37133;
  assign n37135 = ~n34979 & ~n37114;
  assign n37136 = n3485 & ~n37135;
  assign n37137 = ~n37134 & ~n37136;
  assign n37138 = n3476 & ~n37137;
  assign n37139 = ~n37118 & ~n37138;
  assign n37140 = ~n3374 & ~n37139;
  assign n37141 = n3492 & ~n35836;
  assign n37142 = ~n3631 & ~n37141;
  assign n37143 = n3485 & ~n37142;
  assign n37144 = ~n3630 & ~n37143;
  assign n37145 = ~n3476 & ~n37144;
  assign n37146 = n3492 & ~n35921;
  assign n37147 = ~n34979 & ~n37146;
  assign n37148 = n3485 & ~n37147;
  assign n37149 = ~n37134 & ~n37148;
  assign n37150 = n3476 & ~n37149;
  assign n37151 = ~n37145 & ~n37150;
  assign n37152 = n3374 & ~n37151;
  assign n37153 = ~n37140 & ~n37152;
  assign n37154 = ~n3655 & ~n37153;
  assign n37155 = ~n37113 & ~n37154;
  assign n37156 = ~n3652 & ~n37155;
  assign n37157 = ~n37072 & ~n37156;
  assign n37158 = ~n3368 & ~n37157;
  assign n37159 = n3492 & ~n36000;
  assign n37160 = n3492 & ~n37159;
  assign n37161 = n3485 & ~n37160;
  assign n37162 = n3485 & ~n37161;
  assign n37163 = ~n3476 & ~n37162;
  assign n37164 = ~n8525 & ~n37161;
  assign n37165 = n3476 & ~n37164;
  assign n37166 = ~n37163 & ~n37165;
  assign n37167 = ~n3374 & ~n37166;
  assign n37168 = n3492 & ~n36132;
  assign n37169 = n3492 & ~n37168;
  assign n37170 = n3485 & ~n37169;
  assign n37171 = n3485 & ~n37170;
  assign n37172 = ~n3476 & ~n37171;
  assign n37173 = ~n3281 & ~n37004;
  assign n37174 = ~n3492 & ~n37173;
  assign n37175 = n3492 & ~n34053;
  assign n37176 = ~n37174 & ~n37175;
  assign n37177 = ~n3485 & ~n37176;
  assign n37178 = n3492 & ~n36334;
  assign n37179 = ~n34669 & ~n37178;
  assign n37180 = n3485 & ~n37179;
  assign n37181 = ~n37177 & ~n37180;
  assign n37182 = n3476 & ~n37181;
  assign n37183 = ~n37172 & ~n37182;
  assign n37184 = n3374 & ~n37183;
  assign n37185 = ~n37167 & ~n37184;
  assign n37186 = n3655 & ~n37185;
  assign n37187 = n3492 & ~n36375;
  assign n37188 = n3492 & ~n37187;
  assign n37189 = n3485 & ~n37188;
  assign n37190 = n3485 & ~n37189;
  assign n37191 = ~n3476 & ~n37190;
  assign n37192 = ~n8525 & ~n37189;
  assign n37193 = n3476 & ~n37192;
  assign n37194 = ~n37191 & ~n37193;
  assign n37195 = ~n3374 & ~n37194;
  assign n37196 = n3492 & ~n36464;
  assign n37197 = n3492 & ~n37196;
  assign n37198 = n3485 & ~n37197;
  assign n37199 = n3485 & ~n37198;
  assign n37200 = ~n3476 & ~n37199;
  assign n37201 = ~n3281 & ~n37046;
  assign n37202 = ~n3492 & ~n37201;
  assign n37203 = ~n37175 & ~n37202;
  assign n37204 = ~n3485 & ~n37203;
  assign n37205 = n3492 & ~n36588;
  assign n37206 = ~n34669 & ~n37205;
  assign n37207 = n3485 & ~n37206;
  assign n37208 = ~n37204 & ~n37207;
  assign n37209 = n3476 & ~n37208;
  assign n37210 = ~n37200 & ~n37209;
  assign n37211 = n3374 & ~n37210;
  assign n37212 = ~n37195 & ~n37211;
  assign n37213 = ~n3655 & ~n37212;
  assign n37214 = ~n37186 & ~n37213;
  assign n37215 = n3652 & ~n37214;
  assign n37216 = n3492 & ~n36624;
  assign n37217 = n3492 & ~n37216;
  assign n37218 = n3485 & ~n37217;
  assign n37219 = n3485 & ~n37218;
  assign n37220 = ~n3476 & ~n37219;
  assign n37221 = ~n8525 & ~n37218;
  assign n37222 = n3476 & ~n37221;
  assign n37223 = ~n37220 & ~n37222;
  assign n37224 = ~n3374 & ~n37223;
  assign n37225 = n3492 & ~n36695;
  assign n37226 = n3492 & ~n37225;
  assign n37227 = n3485 & ~n37226;
  assign n37228 = n3485 & ~n37227;
  assign n37229 = ~n3476 & ~n37228;
  assign n37230 = ~n3281 & ~n37089;
  assign n37231 = ~n3492 & ~n37230;
  assign n37232 = ~n37175 & ~n37231;
  assign n37233 = ~n3485 & ~n37232;
  assign n37234 = n3492 & ~n36780;
  assign n37235 = ~n34669 & ~n37234;
  assign n37236 = n3485 & ~n37235;
  assign n37237 = ~n37233 & ~n37236;
  assign n37238 = n3476 & ~n37237;
  assign n37239 = ~n37229 & ~n37238;
  assign n37240 = n3374 & ~n37239;
  assign n37241 = ~n37224 & ~n37240;
  assign n37242 = n3655 & ~n37241;
  assign n37243 = n3492 & ~n36814;
  assign n37244 = n3492 & ~n37243;
  assign n37245 = n3485 & ~n37244;
  assign n37246 = n3485 & ~n37245;
  assign n37247 = ~n3476 & ~n37246;
  assign n37248 = ~n8525 & ~n37245;
  assign n37249 = n3476 & ~n37248;
  assign n37250 = ~n37247 & ~n37249;
  assign n37251 = ~n3374 & ~n37250;
  assign n37252 = n3492 & ~n36885;
  assign n37253 = n3492 & ~n37252;
  assign n37254 = n3485 & ~n37253;
  assign n37255 = n3485 & ~n37254;
  assign n37256 = ~n3476 & ~n37255;
  assign n37257 = ~n3281 & ~n37130;
  assign n37258 = ~n3492 & ~n37257;
  assign n37259 = ~n37175 & ~n37258;
  assign n37260 = ~n3485 & ~n37259;
  assign n37261 = n3492 & ~n36970;
  assign n37262 = ~n34669 & ~n37261;
  assign n37263 = n3485 & ~n37262;
  assign n37264 = ~n37260 & ~n37263;
  assign n37265 = n3476 & ~n37264;
  assign n37266 = ~n37256 & ~n37265;
  assign n37267 = n3374 & ~n37266;
  assign n37268 = ~n37251 & ~n37267;
  assign n37269 = ~n3655 & ~n37268;
  assign n37270 = ~n37242 & ~n37269;
  assign n37271 = ~n3652 & ~n37270;
  assign n37272 = ~n37215 & ~n37271;
  assign n37273 = n3368 & ~n37272;
  assign n37274 = ~n37158 & ~n37273;
  assign n37275 = ~n3362 & ~n37274;
  assign n37276 = ~n36987 & ~n37275;
  assign n37277 = n3359 & ~n37276;
  assign n37278 = ~n3485 & ~n37005;
  assign n37279 = ~n37011 & ~n37278;
  assign n37280 = n3476 & ~n37279;
  assign n37281 = ~n36992 & ~n37280;
  assign n37282 = ~n3374 & ~n37281;
  assign n37283 = ~n37023 & ~n37278;
  assign n37284 = n3476 & ~n37283;
  assign n37285 = ~n37020 & ~n37284;
  assign n37286 = n3374 & ~n37285;
  assign n37287 = ~n37282 & ~n37286;
  assign n37288 = n3655 & ~n37287;
  assign n37289 = ~n3485 & ~n37047;
  assign n37290 = ~n37052 & ~n37289;
  assign n37291 = n3476 & ~n37290;
  assign n37292 = ~n37034 & ~n37291;
  assign n37293 = ~n3374 & ~n37292;
  assign n37294 = ~n37064 & ~n37289;
  assign n37295 = n3476 & ~n37294;
  assign n37296 = ~n37061 & ~n37295;
  assign n37297 = n3374 & ~n37296;
  assign n37298 = ~n37293 & ~n37297;
  assign n37299 = ~n3655 & ~n37298;
  assign n37300 = ~n37288 & ~n37299;
  assign n37301 = n3652 & ~n37300;
  assign n37302 = ~n3485 & ~n37090;
  assign n37303 = ~n37095 & ~n37302;
  assign n37304 = n3476 & ~n37303;
  assign n37305 = ~n37077 & ~n37304;
  assign n37306 = ~n3374 & ~n37305;
  assign n37307 = ~n37107 & ~n37302;
  assign n37308 = n3476 & ~n37307;
  assign n37309 = ~n37104 & ~n37308;
  assign n37310 = n3374 & ~n37309;
  assign n37311 = ~n37306 & ~n37310;
  assign n37312 = n3655 & ~n37311;
  assign n37313 = ~n3485 & ~n37131;
  assign n37314 = ~n37136 & ~n37313;
  assign n37315 = n3476 & ~n37314;
  assign n37316 = ~n37118 & ~n37315;
  assign n37317 = ~n3374 & ~n37316;
  assign n37318 = ~n37148 & ~n37313;
  assign n37319 = n3476 & ~n37318;
  assign n37320 = ~n37145 & ~n37319;
  assign n37321 = n3374 & ~n37320;
  assign n37322 = ~n37317 & ~n37321;
  assign n37323 = ~n3655 & ~n37322;
  assign n37324 = ~n37312 & ~n37323;
  assign n37325 = ~n3652 & ~n37324;
  assign n37326 = ~n37301 & ~n37325;
  assign n37327 = ~n3368 & ~n37326;
  assign n37328 = ~n8689 & ~n37161;
  assign n37329 = n3476 & ~n37328;
  assign n37330 = ~n37163 & ~n37329;
  assign n37331 = ~n3374 & ~n37330;
  assign n37332 = ~n3485 & ~n37173;
  assign n37333 = ~n37180 & ~n37332;
  assign n37334 = n3476 & ~n37333;
  assign n37335 = ~n37172 & ~n37334;
  assign n37336 = n3374 & ~n37335;
  assign n37337 = ~n37331 & ~n37336;
  assign n37338 = n3655 & ~n37337;
  assign n37339 = ~n8689 & ~n37189;
  assign n37340 = n3476 & ~n37339;
  assign n37341 = ~n37191 & ~n37340;
  assign n37342 = ~n3374 & ~n37341;
  assign n37343 = ~n3485 & ~n37201;
  assign n37344 = ~n37207 & ~n37343;
  assign n37345 = n3476 & ~n37344;
  assign n37346 = ~n37200 & ~n37345;
  assign n37347 = n3374 & ~n37346;
  assign n37348 = ~n37342 & ~n37347;
  assign n37349 = ~n3655 & ~n37348;
  assign n37350 = ~n37338 & ~n37349;
  assign n37351 = n3652 & ~n37350;
  assign n37352 = ~n8689 & ~n37218;
  assign n37353 = n3476 & ~n37352;
  assign n37354 = ~n37220 & ~n37353;
  assign n37355 = ~n3374 & ~n37354;
  assign n37356 = ~n3485 & ~n37230;
  assign n37357 = ~n37236 & ~n37356;
  assign n37358 = n3476 & ~n37357;
  assign n37359 = ~n37229 & ~n37358;
  assign n37360 = n3374 & ~n37359;
  assign n37361 = ~n37355 & ~n37360;
  assign n37362 = n3655 & ~n37361;
  assign n37363 = ~n8689 & ~n37245;
  assign n37364 = n3476 & ~n37363;
  assign n37365 = ~n37247 & ~n37364;
  assign n37366 = ~n3374 & ~n37365;
  assign n37367 = ~n3485 & ~n37257;
  assign n37368 = ~n37263 & ~n37367;
  assign n37369 = n3476 & ~n37368;
  assign n37370 = ~n37256 & ~n37369;
  assign n37371 = n3374 & ~n37370;
  assign n37372 = ~n37366 & ~n37371;
  assign n37373 = ~n3655 & ~n37372;
  assign n37374 = ~n37362 & ~n37373;
  assign n37375 = ~n3652 & ~n37374;
  assign n37376 = ~n37351 & ~n37375;
  assign n37377 = n3368 & ~n37376;
  assign n37378 = ~n37327 & ~n37377;
  assign n37379 = n3362 & ~n37378;
  assign n37380 = n3378 & ~n34970;
  assign n37381 = ~n34022 & ~n34156;
  assign n37382 = ~controllable_hmaster1 & ~n37381;
  assign n37383 = ~n34155 & ~n37382;
  assign n37384 = i_hbusreq3 & ~n37383;
  assign n37385 = ~n34040 & ~n34156;
  assign n37386 = ~controllable_hmaster1 & ~n37385;
  assign n37387 = ~n34155 & ~n37386;
  assign n37388 = ~i_hbusreq3 & ~n37387;
  assign n37389 = ~n37384 & ~n37388;
  assign n37390 = controllable_hmaster2 & ~n37389;
  assign n37391 = ~n5161 & ~n37390;
  assign n37392 = ~controllable_hgrant3 & ~n37391;
  assign n37393 = ~n8750 & ~n37392;
  assign n37394 = controllable_nhgrant0 & ~n37393;
  assign n37395 = ~n8785 & ~n37394;
  assign n37396 = ~n3281 & ~n37395;
  assign n37397 = ~n3783 & ~n37396;
  assign n37398 = ~n3378 & ~n37397;
  assign n37399 = ~n37380 & ~n37398;
  assign n37400 = n3492 & ~n37399;
  assign n37401 = ~n3631 & ~n37400;
  assign n37402 = n3485 & ~n37401;
  assign n37403 = ~n3630 & ~n37402;
  assign n37404 = ~n3476 & ~n37403;
  assign n37405 = ~n37006 & ~n37400;
  assign n37406 = n3485 & ~n37405;
  assign n37407 = ~n37278 & ~n37406;
  assign n37408 = n3476 & ~n37407;
  assign n37409 = ~n37404 & ~n37408;
  assign n37410 = ~n3374 & ~n37409;
  assign n37411 = n3378 & ~n35102;
  assign n37412 = ~n34137 & ~n34156;
  assign n37413 = ~controllable_hmaster1 & ~n37412;
  assign n37414 = ~n34155 & ~n37413;
  assign n37415 = ~i_hbusreq3 & ~n37414;
  assign n37416 = ~n34160 & ~n37415;
  assign n37417 = controllable_hmaster2 & ~n37416;
  assign n37418 = ~n3850 & ~n34986;
  assign n37419 = ~controllable_hgrant2 & ~n37418;
  assign n37420 = ~n3410 & ~n37419;
  assign n37421 = controllable_hmaster0 & ~n37420;
  assign n37422 = ~n5288 & ~n37419;
  assign n37423 = ~controllable_hmaster0 & ~n37422;
  assign n37424 = ~n37421 & ~n37423;
  assign n37425 = controllable_hmaster1 & ~n37424;
  assign n37426 = ~n8822 & ~n34986;
  assign n37427 = ~controllable_hgrant2 & ~n37426;
  assign n37428 = ~n3410 & ~n37427;
  assign n37429 = controllable_hmaster0 & ~n37428;
  assign n37430 = ~controllable_hmaster0 & ~n37420;
  assign n37431 = ~n37429 & ~n37430;
  assign n37432 = ~controllable_hmaster1 & ~n37431;
  assign n37433 = ~n37425 & ~n37432;
  assign n37434 = i_hbusreq3 & ~n37433;
  assign n37435 = i_hbusreq2 & ~n37418;
  assign n37436 = ~n3884 & ~n35078;
  assign n37437 = ~i_hbusreq2 & ~n37436;
  assign n37438 = ~n37435 & ~n37437;
  assign n37439 = ~controllable_hgrant2 & ~n37438;
  assign n37440 = ~n3859 & ~n37439;
  assign n37441 = controllable_hmaster0 & ~n37440;
  assign n37442 = ~n5438 & ~n37439;
  assign n37443 = ~controllable_hmaster0 & ~n37442;
  assign n37444 = ~n37441 & ~n37443;
  assign n37445 = controllable_hmaster1 & ~n37444;
  assign n37446 = i_hbusreq2 & ~n37426;
  assign n37447 = ~n8854 & ~n35078;
  assign n37448 = ~i_hbusreq2 & ~n37447;
  assign n37449 = ~n37446 & ~n37448;
  assign n37450 = ~controllable_hgrant2 & ~n37449;
  assign n37451 = ~n3859 & ~n37450;
  assign n37452 = controllable_hmaster0 & ~n37451;
  assign n37453 = ~n8870 & ~n35392;
  assign n37454 = ~i_hbusreq2 & ~n37453;
  assign n37455 = ~n37435 & ~n37454;
  assign n37456 = ~controllable_hgrant2 & ~n37455;
  assign n37457 = ~n5461 & ~n37456;
  assign n37458 = ~controllable_hmaster0 & ~n37457;
  assign n37459 = ~n37452 & ~n37458;
  assign n37460 = ~controllable_hmaster1 & ~n37459;
  assign n37461 = ~n37445 & ~n37460;
  assign n37462 = ~i_hbusreq3 & ~n37461;
  assign n37463 = ~n37434 & ~n37462;
  assign n37464 = ~controllable_hmaster2 & ~n37463;
  assign n37465 = ~n37417 & ~n37464;
  assign n37466 = ~controllable_hgrant3 & ~n37465;
  assign n37467 = ~n8810 & ~n37466;
  assign n37468 = controllable_nhgrant0 & ~n37467;
  assign n37469 = ~n8902 & ~n37468;
  assign n37470 = ~n3281 & ~n37469;
  assign n37471 = ~n3950 & ~n37470;
  assign n37472 = ~n3378 & ~n37471;
  assign n37473 = ~n37411 & ~n37472;
  assign n37474 = n3492 & ~n37473;
  assign n37475 = ~n3631 & ~n37474;
  assign n37476 = n3485 & ~n37475;
  assign n37477 = ~n3630 & ~n37476;
  assign n37478 = ~n3476 & ~n37477;
  assign n37479 = n3378 & ~n35271;
  assign n37480 = controllable_hgrant4 & ~n9077;
  assign n37481 = ~n8950 & ~n37480;
  assign n37482 = ~i_hbusreq2 & ~n37481;
  assign n37483 = ~n35123 & ~n37482;
  assign n37484 = ~controllable_hgrant2 & ~n37483;
  assign n37485 = ~n8936 & ~n37484;
  assign n37486 = controllable_hmaster1 & ~n37485;
  assign n37487 = controllable_hmaster0 & ~n37485;
  assign n37488 = ~n8969 & ~n34214;
  assign n37489 = ~i_hbusreq2 & ~n37488;
  assign n37490 = ~n35131 & ~n37489;
  assign n37491 = ~controllable_hgrant2 & ~n37490;
  assign n37492 = ~n5862 & ~n37491;
  assign n37493 = ~controllable_hmaster0 & ~n37492;
  assign n37494 = ~n37487 & ~n37493;
  assign n37495 = ~controllable_hmaster1 & ~n37494;
  assign n37496 = ~n37486 & ~n37495;
  assign n37497 = ~i_hbusreq3 & ~n37496;
  assign n37498 = ~n35122 & ~n37497;
  assign n37499 = controllable_hmaster2 & ~n37498;
  assign n37500 = ~n5621 & ~n35144;
  assign n37501 = ~controllable_hgrant2 & ~n37500;
  assign n37502 = ~n5616 & ~n37501;
  assign n37503 = controllable_hmaster0 & ~n37502;
  assign n37504 = ~n5686 & ~n37501;
  assign n37505 = ~controllable_hmaster0 & ~n37504;
  assign n37506 = ~n37503 & ~n37505;
  assign n37507 = controllable_hmaster1 & ~n37506;
  assign n37508 = ~n8987 & ~n35144;
  assign n37509 = ~controllable_hgrant2 & ~n37508;
  assign n37510 = ~n5616 & ~n37509;
  assign n37511 = controllable_hmaster0 & ~n37510;
  assign n37512 = ~controllable_hmaster0 & ~n37502;
  assign n37513 = ~n37511 & ~n37512;
  assign n37514 = ~controllable_hmaster1 & ~n37513;
  assign n37515 = ~n37507 & ~n37514;
  assign n37516 = i_hbusreq3 & ~n37515;
  assign n37517 = i_hbusreq2 & ~n37500;
  assign n37518 = ~n8969 & ~n35234;
  assign n37519 = ~i_hbusreq2 & ~n37518;
  assign n37520 = ~n37517 & ~n37519;
  assign n37521 = ~controllable_hgrant2 & ~n37520;
  assign n37522 = ~n5862 & ~n37521;
  assign n37523 = controllable_hmaster0 & ~n37522;
  assign n37524 = ~n5950 & ~n37521;
  assign n37525 = ~controllable_hmaster0 & ~n37524;
  assign n37526 = ~n37523 & ~n37525;
  assign n37527 = controllable_hmaster1 & ~n37526;
  assign n37528 = i_hbusreq2 & ~n37508;
  assign n37529 = ~n9024 & ~n35234;
  assign n37530 = ~i_hbusreq2 & ~n37529;
  assign n37531 = ~n37528 & ~n37530;
  assign n37532 = ~controllable_hgrant2 & ~n37531;
  assign n37533 = ~n5862 & ~n37532;
  assign n37534 = controllable_hmaster0 & ~n37533;
  assign n37535 = ~n9038 & ~n35252;
  assign n37536 = ~i_hbusreq2 & ~n37535;
  assign n37537 = ~n37517 & ~n37536;
  assign n37538 = ~controllable_hgrant2 & ~n37537;
  assign n37539 = ~n5981 & ~n37538;
  assign n37540 = ~controllable_hmaster0 & ~n37539;
  assign n37541 = ~n37534 & ~n37540;
  assign n37542 = ~controllable_hmaster1 & ~n37541;
  assign n37543 = ~n37527 & ~n37542;
  assign n37544 = ~i_hbusreq3 & ~n37543;
  assign n37545 = ~n37516 & ~n37544;
  assign n37546 = ~controllable_hmaster2 & ~n37545;
  assign n37547 = ~n37499 & ~n37546;
  assign n37548 = ~controllable_hgrant3 & ~n37547;
  assign n37549 = ~n8935 & ~n37548;
  assign n37550 = controllable_nhgrant0 & ~n37549;
  assign n37551 = ~n9096 & ~n37550;
  assign n37552 = ~n3281 & ~n37551;
  assign n37553 = ~n4089 & ~n37552;
  assign n37554 = ~n3378 & ~n37553;
  assign n37555 = ~n37479 & ~n37554;
  assign n37556 = n3492 & ~n37555;
  assign n37557 = ~n37006 & ~n37556;
  assign n37558 = n3485 & ~n37557;
  assign n37559 = ~n37278 & ~n37558;
  assign n37560 = n3476 & ~n37559;
  assign n37561 = ~n37478 & ~n37560;
  assign n37562 = n3374 & ~n37561;
  assign n37563 = ~n37410 & ~n37562;
  assign n37564 = n3655 & ~n37563;
  assign n37565 = n3378 & ~n35312;
  assign n37566 = ~n9112 & ~n34055;
  assign n37567 = ~controllable_hgrant2 & ~n37566;
  assign n37568 = ~n3410 & ~n37567;
  assign n37569 = controllable_hmaster1 & ~n37568;
  assign n37570 = controllable_hmaster0 & ~n37568;
  assign n37571 = ~n34022 & ~n37570;
  assign n37572 = ~controllable_hmaster1 & ~n37571;
  assign n37573 = ~n37569 & ~n37572;
  assign n37574 = i_hbusreq3 & ~n37573;
  assign n37575 = ~n34040 & ~n37570;
  assign n37576 = ~controllable_hmaster1 & ~n37575;
  assign n37577 = ~n37569 & ~n37576;
  assign n37578 = ~i_hbusreq3 & ~n37577;
  assign n37579 = ~n37574 & ~n37578;
  assign n37580 = controllable_hmaster2 & ~n37579;
  assign n37581 = ~n6188 & ~n37580;
  assign n37582 = ~controllable_hgrant3 & ~n37581;
  assign n37583 = ~n8750 & ~n37582;
  assign n37584 = controllable_nhgrant0 & ~n37583;
  assign n37585 = ~n8785 & ~n37584;
  assign n37586 = ~n3281 & ~n37585;
  assign n37587 = ~n3783 & ~n37586;
  assign n37588 = ~n3378 & ~n37587;
  assign n37589 = ~n37565 & ~n37588;
  assign n37590 = n3492 & ~n37589;
  assign n37591 = ~n3631 & ~n37590;
  assign n37592 = n3485 & ~n37591;
  assign n37593 = ~n3630 & ~n37592;
  assign n37594 = ~n3476 & ~n37593;
  assign n37595 = ~n37048 & ~n37590;
  assign n37596 = n3485 & ~n37595;
  assign n37597 = ~n37289 & ~n37596;
  assign n37598 = n3476 & ~n37597;
  assign n37599 = ~n37594 & ~n37598;
  assign n37600 = ~n3374 & ~n37599;
  assign n37601 = n3378 & ~n35411;
  assign n37602 = ~n34309 & ~n37570;
  assign n37603 = ~controllable_hmaster1 & ~n37602;
  assign n37604 = ~n37569 & ~n37603;
  assign n37605 = i_hbusreq3 & ~n37604;
  assign n37606 = ~n34320 & ~n37570;
  assign n37607 = ~controllable_hmaster1 & ~n37606;
  assign n37608 = ~n37569 & ~n37607;
  assign n37609 = ~i_hbusreq3 & ~n37608;
  assign n37610 = ~n37605 & ~n37609;
  assign n37611 = controllable_hmaster2 & ~n37610;
  assign n37612 = ~n4182 & ~n34986;
  assign n37613 = ~controllable_hgrant2 & ~n37612;
  assign n37614 = ~n3410 & ~n37613;
  assign n37615 = controllable_hmaster0 & ~n37614;
  assign n37616 = ~n5288 & ~n37613;
  assign n37617 = ~controllable_hmaster0 & ~n37616;
  assign n37618 = ~n37615 & ~n37617;
  assign n37619 = controllable_hmaster1 & ~n37618;
  assign n37620 = ~n9170 & ~n34986;
  assign n37621 = ~controllable_hgrant2 & ~n37620;
  assign n37622 = ~n3410 & ~n37621;
  assign n37623 = controllable_hmaster0 & ~n37622;
  assign n37624 = ~controllable_hmaster0 & ~n37614;
  assign n37625 = ~n37623 & ~n37624;
  assign n37626 = ~controllable_hmaster1 & ~n37625;
  assign n37627 = ~n37619 & ~n37626;
  assign n37628 = i_hbusreq3 & ~n37627;
  assign n37629 = i_hbusreq2 & ~n37612;
  assign n37630 = ~n4204 & ~n35078;
  assign n37631 = ~i_hbusreq2 & ~n37630;
  assign n37632 = ~n37629 & ~n37631;
  assign n37633 = ~controllable_hgrant2 & ~n37632;
  assign n37634 = ~n3859 & ~n37633;
  assign n37635 = controllable_hmaster0 & ~n37634;
  assign n37636 = ~n5438 & ~n37633;
  assign n37637 = ~controllable_hmaster0 & ~n37636;
  assign n37638 = ~n37635 & ~n37637;
  assign n37639 = controllable_hmaster1 & ~n37638;
  assign n37640 = i_hbusreq2 & ~n37620;
  assign n37641 = ~n9204 & ~n35078;
  assign n37642 = ~i_hbusreq2 & ~n37641;
  assign n37643 = ~n37640 & ~n37642;
  assign n37644 = ~controllable_hgrant2 & ~n37643;
  assign n37645 = ~n3859 & ~n37644;
  assign n37646 = controllable_hmaster0 & ~n37645;
  assign n37647 = ~n9220 & ~n35392;
  assign n37648 = ~i_hbusreq2 & ~n37647;
  assign n37649 = ~n37629 & ~n37648;
  assign n37650 = ~controllable_hgrant2 & ~n37649;
  assign n37651 = ~n5461 & ~n37650;
  assign n37652 = ~controllable_hmaster0 & ~n37651;
  assign n37653 = ~n37646 & ~n37652;
  assign n37654 = ~controllable_hmaster1 & ~n37653;
  assign n37655 = ~n37639 & ~n37654;
  assign n37656 = ~i_hbusreq3 & ~n37655;
  assign n37657 = ~n37628 & ~n37656;
  assign n37658 = ~controllable_hmaster2 & ~n37657;
  assign n37659 = ~n37611 & ~n37658;
  assign n37660 = ~controllable_hgrant3 & ~n37659;
  assign n37661 = ~n8810 & ~n37660;
  assign n37662 = controllable_nhgrant0 & ~n37661;
  assign n37663 = ~n8902 & ~n37662;
  assign n37664 = ~n3281 & ~n37663;
  assign n37665 = ~n3950 & ~n37664;
  assign n37666 = ~n3378 & ~n37665;
  assign n37667 = ~n37601 & ~n37666;
  assign n37668 = n3492 & ~n37667;
  assign n37669 = ~n3631 & ~n37668;
  assign n37670 = n3485 & ~n37669;
  assign n37671 = ~n3630 & ~n37670;
  assign n37672 = ~n3476 & ~n37671;
  assign n37673 = n3378 & ~n35535;
  assign n37674 = ~n9248 & ~n34239;
  assign n37675 = ~controllable_hgrant2 & ~n37674;
  assign n37676 = ~n5616 & ~n37675;
  assign n37677 = controllable_hmaster1 & ~n37676;
  assign n37678 = controllable_hmaster0 & ~n37676;
  assign n37679 = ~n35456 & ~n37678;
  assign n37680 = ~controllable_hmaster1 & ~n37679;
  assign n37681 = ~n37677 & ~n37680;
  assign n37682 = i_hbusreq3 & ~n37681;
  assign n37683 = i_hbusreq2 & ~n37674;
  assign n37684 = ~n9270 & ~n37480;
  assign n37685 = ~i_hbusreq2 & ~n37684;
  assign n37686 = ~n37683 & ~n37685;
  assign n37687 = ~controllable_hgrant2 & ~n37686;
  assign n37688 = ~n8936 & ~n37687;
  assign n37689 = controllable_hmaster1 & ~n37688;
  assign n37690 = controllable_hmaster0 & ~n37688;
  assign n37691 = ~n9287 & ~n34214;
  assign n37692 = ~i_hbusreq2 & ~n37691;
  assign n37693 = ~n35469 & ~n37692;
  assign n37694 = ~controllable_hgrant2 & ~n37693;
  assign n37695 = ~n5862 & ~n37694;
  assign n37696 = ~controllable_hmaster0 & ~n37695;
  assign n37697 = ~n37690 & ~n37696;
  assign n37698 = ~controllable_hmaster1 & ~n37697;
  assign n37699 = ~n37689 & ~n37698;
  assign n37700 = ~i_hbusreq3 & ~n37699;
  assign n37701 = ~n37682 & ~n37700;
  assign n37702 = controllable_hmaster2 & ~n37701;
  assign n37703 = ~n6403 & ~n35144;
  assign n37704 = ~controllable_hgrant2 & ~n37703;
  assign n37705 = ~n5616 & ~n37704;
  assign n37706 = controllable_hmaster0 & ~n37705;
  assign n37707 = ~n5686 & ~n37704;
  assign n37708 = ~controllable_hmaster0 & ~n37707;
  assign n37709 = ~n37706 & ~n37708;
  assign n37710 = controllable_hmaster1 & ~n37709;
  assign n37711 = ~n9305 & ~n35144;
  assign n37712 = ~controllable_hgrant2 & ~n37711;
  assign n37713 = ~n5616 & ~n37712;
  assign n37714 = controllable_hmaster0 & ~n37713;
  assign n37715 = ~controllable_hmaster0 & ~n37705;
  assign n37716 = ~n37714 & ~n37715;
  assign n37717 = ~controllable_hmaster1 & ~n37716;
  assign n37718 = ~n37710 & ~n37717;
  assign n37719 = i_hbusreq3 & ~n37718;
  assign n37720 = i_hbusreq2 & ~n37703;
  assign n37721 = ~n9287 & ~n35234;
  assign n37722 = ~i_hbusreq2 & ~n37721;
  assign n37723 = ~n37720 & ~n37722;
  assign n37724 = ~controllable_hgrant2 & ~n37723;
  assign n37725 = ~n5862 & ~n37724;
  assign n37726 = controllable_hmaster0 & ~n37725;
  assign n37727 = ~n5950 & ~n37724;
  assign n37728 = ~controllable_hmaster0 & ~n37727;
  assign n37729 = ~n37726 & ~n37728;
  assign n37730 = controllable_hmaster1 & ~n37729;
  assign n37731 = i_hbusreq2 & ~n37711;
  assign n37732 = ~n9340 & ~n35234;
  assign n37733 = ~i_hbusreq2 & ~n37732;
  assign n37734 = ~n37731 & ~n37733;
  assign n37735 = ~controllable_hgrant2 & ~n37734;
  assign n37736 = ~n5862 & ~n37735;
  assign n37737 = controllable_hmaster0 & ~n37736;
  assign n37738 = ~n9354 & ~n35252;
  assign n37739 = ~i_hbusreq2 & ~n37738;
  assign n37740 = ~n37720 & ~n37739;
  assign n37741 = ~controllable_hgrant2 & ~n37740;
  assign n37742 = ~n5981 & ~n37741;
  assign n37743 = ~controllable_hmaster0 & ~n37742;
  assign n37744 = ~n37737 & ~n37743;
  assign n37745 = ~controllable_hmaster1 & ~n37744;
  assign n37746 = ~n37730 & ~n37745;
  assign n37747 = ~i_hbusreq3 & ~n37746;
  assign n37748 = ~n37719 & ~n37747;
  assign n37749 = ~controllable_hmaster2 & ~n37748;
  assign n37750 = ~n37702 & ~n37749;
  assign n37751 = ~controllable_hgrant3 & ~n37750;
  assign n37752 = ~n8935 & ~n37751;
  assign n37753 = controllable_nhgrant0 & ~n37752;
  assign n37754 = ~n9096 & ~n37753;
  assign n37755 = ~n3281 & ~n37754;
  assign n37756 = ~n4089 & ~n37755;
  assign n37757 = ~n3378 & ~n37756;
  assign n37758 = ~n37673 & ~n37757;
  assign n37759 = n3492 & ~n37758;
  assign n37760 = ~n37048 & ~n37759;
  assign n37761 = n3485 & ~n37760;
  assign n37762 = ~n37289 & ~n37761;
  assign n37763 = n3476 & ~n37762;
  assign n37764 = ~n37672 & ~n37763;
  assign n37765 = n3374 & ~n37764;
  assign n37766 = ~n37600 & ~n37765;
  assign n37767 = ~n3655 & ~n37766;
  assign n37768 = ~n37564 & ~n37767;
  assign n37769 = n3652 & ~n37768;
  assign n37770 = n3378 & ~n35571;
  assign n37771 = ~n9388 & ~n34153;
  assign n37772 = controllable_hmaster1 & ~n37771;
  assign n37773 = controllable_hmaster0 & ~n37771;
  assign n37774 = ~n34022 & ~n37773;
  assign n37775 = ~controllable_hmaster1 & ~n37774;
  assign n37776 = ~n37772 & ~n37775;
  assign n37777 = i_hbusreq3 & ~n37776;
  assign n37778 = ~n34040 & ~n37773;
  assign n37779 = ~controllable_hmaster1 & ~n37778;
  assign n37780 = ~n37772 & ~n37779;
  assign n37781 = ~i_hbusreq3 & ~n37780;
  assign n37782 = ~n37777 & ~n37781;
  assign n37783 = controllable_hmaster2 & ~n37782;
  assign n37784 = ~n6657 & ~n37783;
  assign n37785 = ~controllable_hgrant3 & ~n37784;
  assign n37786 = ~n8750 & ~n37785;
  assign n37787 = controllable_nhgrant0 & ~n37786;
  assign n37788 = ~n8785 & ~n37787;
  assign n37789 = ~n3281 & ~n37788;
  assign n37790 = ~n3783 & ~n37789;
  assign n37791 = ~n3378 & ~n37790;
  assign n37792 = ~n37770 & ~n37791;
  assign n37793 = n3492 & ~n37792;
  assign n37794 = ~n3631 & ~n37793;
  assign n37795 = n3485 & ~n37794;
  assign n37796 = ~n3630 & ~n37795;
  assign n37797 = ~n3476 & ~n37796;
  assign n37798 = ~n37091 & ~n37793;
  assign n37799 = n3485 & ~n37798;
  assign n37800 = ~n37302 & ~n37799;
  assign n37801 = n3476 & ~n37800;
  assign n37802 = ~n37797 & ~n37801;
  assign n37803 = ~n3374 & ~n37802;
  assign n37804 = n3378 & ~n35644;
  assign n37805 = ~n34430 & ~n37773;
  assign n37806 = ~controllable_hmaster1 & ~n37805;
  assign n37807 = ~n37772 & ~n37806;
  assign n37808 = i_hbusreq3 & ~n37807;
  assign n37809 = ~n34436 & ~n37773;
  assign n37810 = ~controllable_hmaster1 & ~n37809;
  assign n37811 = ~n37772 & ~n37810;
  assign n37812 = ~i_hbusreq3 & ~n37811;
  assign n37813 = ~n37808 & ~n37812;
  assign n37814 = controllable_hmaster2 & ~n37813;
  assign n37815 = ~n4333 & ~n37419;
  assign n37816 = controllable_hmaster0 & ~n37815;
  assign n37817 = ~n6697 & ~n37419;
  assign n37818 = ~controllable_hmaster0 & ~n37817;
  assign n37819 = ~n37816 & ~n37818;
  assign n37820 = controllable_hmaster1 & ~n37819;
  assign n37821 = ~n4333 & ~n37427;
  assign n37822 = controllable_hmaster0 & ~n37821;
  assign n37823 = ~controllable_hmaster0 & ~n37815;
  assign n37824 = ~n37822 & ~n37823;
  assign n37825 = ~controllable_hmaster1 & ~n37824;
  assign n37826 = ~n37820 & ~n37825;
  assign n37827 = i_hbusreq3 & ~n37826;
  assign n37828 = ~n4340 & ~n37439;
  assign n37829 = controllable_hmaster0 & ~n37828;
  assign n37830 = ~n6710 & ~n37439;
  assign n37831 = ~controllable_hmaster0 & ~n37830;
  assign n37832 = ~n37829 & ~n37831;
  assign n37833 = controllable_hmaster1 & ~n37832;
  assign n37834 = ~n4340 & ~n37450;
  assign n37835 = controllable_hmaster0 & ~n37834;
  assign n37836 = ~n6947 & ~n37456;
  assign n37837 = ~controllable_hmaster0 & ~n37836;
  assign n37838 = ~n37835 & ~n37837;
  assign n37839 = ~controllable_hmaster1 & ~n37838;
  assign n37840 = ~n37833 & ~n37839;
  assign n37841 = ~i_hbusreq3 & ~n37840;
  assign n37842 = ~n37827 & ~n37841;
  assign n37843 = ~controllable_hmaster2 & ~n37842;
  assign n37844 = ~n37814 & ~n37843;
  assign n37845 = ~controllable_hgrant3 & ~n37844;
  assign n37846 = ~n8810 & ~n37845;
  assign n37847 = controllable_nhgrant0 & ~n37846;
  assign n37848 = ~n8902 & ~n37847;
  assign n37849 = ~n3281 & ~n37848;
  assign n37850 = ~n3950 & ~n37849;
  assign n37851 = ~n3378 & ~n37850;
  assign n37852 = ~n37804 & ~n37851;
  assign n37853 = n3492 & ~n37852;
  assign n37854 = ~n3631 & ~n37853;
  assign n37855 = n3485 & ~n37854;
  assign n37856 = ~n3630 & ~n37855;
  assign n37857 = ~n3476 & ~n37856;
  assign n37858 = n3378 & ~n35729;
  assign n37859 = ~n9477 & ~n35111;
  assign n37860 = controllable_hmaster1 & ~n37859;
  assign n37861 = controllable_hmaster0 & ~n37859;
  assign n37862 = ~n35678 & ~n37861;
  assign n37863 = ~controllable_hmaster1 & ~n37862;
  assign n37864 = ~n37860 & ~n37863;
  assign n37865 = i_hbusreq3 & ~n37864;
  assign n37866 = ~n9485 & ~n37484;
  assign n37867 = controllable_hmaster1 & ~n37866;
  assign n37868 = controllable_hmaster0 & ~n37866;
  assign n37869 = ~n6772 & ~n37491;
  assign n37870 = ~controllable_hmaster0 & ~n37869;
  assign n37871 = ~n37868 & ~n37870;
  assign n37872 = ~controllable_hmaster1 & ~n37871;
  assign n37873 = ~n37867 & ~n37872;
  assign n37874 = ~i_hbusreq3 & ~n37873;
  assign n37875 = ~n37865 & ~n37874;
  assign n37876 = controllable_hmaster2 & ~n37875;
  assign n37877 = ~n6762 & ~n37501;
  assign n37878 = controllable_hmaster0 & ~n37877;
  assign n37879 = ~n6786 & ~n37501;
  assign n37880 = ~controllable_hmaster0 & ~n37879;
  assign n37881 = ~n37878 & ~n37880;
  assign n37882 = controllable_hmaster1 & ~n37881;
  assign n37883 = ~n6762 & ~n37509;
  assign n37884 = controllable_hmaster0 & ~n37883;
  assign n37885 = ~controllable_hmaster0 & ~n37877;
  assign n37886 = ~n37884 & ~n37885;
  assign n37887 = ~controllable_hmaster1 & ~n37886;
  assign n37888 = ~n37882 & ~n37887;
  assign n37889 = i_hbusreq3 & ~n37888;
  assign n37890 = ~n6772 & ~n37521;
  assign n37891 = controllable_hmaster0 & ~n37890;
  assign n37892 = ~n6813 & ~n37521;
  assign n37893 = ~controllable_hmaster0 & ~n37892;
  assign n37894 = ~n37891 & ~n37893;
  assign n37895 = controllable_hmaster1 & ~n37894;
  assign n37896 = ~n6772 & ~n37532;
  assign n37897 = controllable_hmaster0 & ~n37896;
  assign n37898 = ~n6831 & ~n37538;
  assign n37899 = ~controllable_hmaster0 & ~n37898;
  assign n37900 = ~n37897 & ~n37899;
  assign n37901 = ~controllable_hmaster1 & ~n37900;
  assign n37902 = ~n37895 & ~n37901;
  assign n37903 = ~i_hbusreq3 & ~n37902;
  assign n37904 = ~n37889 & ~n37903;
  assign n37905 = ~controllable_hmaster2 & ~n37904;
  assign n37906 = ~n37876 & ~n37905;
  assign n37907 = ~controllable_hgrant3 & ~n37906;
  assign n37908 = ~n8935 & ~n37907;
  assign n37909 = controllable_nhgrant0 & ~n37908;
  assign n37910 = ~n9096 & ~n37909;
  assign n37911 = ~n3281 & ~n37910;
  assign n37912 = ~n4089 & ~n37911;
  assign n37913 = ~n3378 & ~n37912;
  assign n37914 = ~n37858 & ~n37913;
  assign n37915 = n3492 & ~n37914;
  assign n37916 = ~n37091 & ~n37915;
  assign n37917 = n3485 & ~n37916;
  assign n37918 = ~n37302 & ~n37917;
  assign n37919 = n3476 & ~n37918;
  assign n37920 = ~n37857 & ~n37919;
  assign n37921 = n3374 & ~n37920;
  assign n37922 = ~n37803 & ~n37921;
  assign n37923 = n3655 & ~n37922;
  assign n37924 = n3378 & ~n35763;
  assign n37925 = ~n9388 & ~n37567;
  assign n37926 = controllable_hmaster1 & ~n37925;
  assign n37927 = controllable_hmaster0 & ~n37925;
  assign n37928 = ~n34022 & ~n37927;
  assign n37929 = ~controllable_hmaster1 & ~n37928;
  assign n37930 = ~n37926 & ~n37929;
  assign n37931 = i_hbusreq3 & ~n37930;
  assign n37932 = ~n34040 & ~n37927;
  assign n37933 = ~controllable_hmaster1 & ~n37932;
  assign n37934 = ~n37926 & ~n37933;
  assign n37935 = ~i_hbusreq3 & ~n37934;
  assign n37936 = ~n37931 & ~n37935;
  assign n37937 = controllable_hmaster2 & ~n37936;
  assign n37938 = ~n6887 & ~n37937;
  assign n37939 = ~controllable_hgrant3 & ~n37938;
  assign n37940 = ~n8750 & ~n37939;
  assign n37941 = controllable_nhgrant0 & ~n37940;
  assign n37942 = ~n8785 & ~n37941;
  assign n37943 = ~n3281 & ~n37942;
  assign n37944 = ~n3783 & ~n37943;
  assign n37945 = ~n3378 & ~n37944;
  assign n37946 = ~n37924 & ~n37945;
  assign n37947 = n3492 & ~n37946;
  assign n37948 = ~n3631 & ~n37947;
  assign n37949 = n3485 & ~n37948;
  assign n37950 = ~n3630 & ~n37949;
  assign n37951 = ~n3476 & ~n37950;
  assign n37952 = ~n37132 & ~n37947;
  assign n37953 = n3485 & ~n37952;
  assign n37954 = ~n37313 & ~n37953;
  assign n37955 = n3476 & ~n37954;
  assign n37956 = ~n37951 & ~n37955;
  assign n37957 = ~n3374 & ~n37956;
  assign n37958 = n3378 & ~n35836;
  assign n37959 = ~n34530 & ~n37927;
  assign n37960 = ~controllable_hmaster1 & ~n37959;
  assign n37961 = ~n37926 & ~n37960;
  assign n37962 = i_hbusreq3 & ~n37961;
  assign n37963 = ~n34536 & ~n37927;
  assign n37964 = ~controllable_hmaster1 & ~n37963;
  assign n37965 = ~n37926 & ~n37964;
  assign n37966 = ~i_hbusreq3 & ~n37965;
  assign n37967 = ~n37962 & ~n37966;
  assign n37968 = controllable_hmaster2 & ~n37967;
  assign n37969 = ~n4333 & ~n37613;
  assign n37970 = controllable_hmaster0 & ~n37969;
  assign n37971 = ~n6697 & ~n37613;
  assign n37972 = ~controllable_hmaster0 & ~n37971;
  assign n37973 = ~n37970 & ~n37972;
  assign n37974 = controllable_hmaster1 & ~n37973;
  assign n37975 = ~n4333 & ~n37621;
  assign n37976 = controllable_hmaster0 & ~n37975;
  assign n37977 = ~controllable_hmaster0 & ~n37969;
  assign n37978 = ~n37976 & ~n37977;
  assign n37979 = ~controllable_hmaster1 & ~n37978;
  assign n37980 = ~n37974 & ~n37979;
  assign n37981 = i_hbusreq3 & ~n37980;
  assign n37982 = ~n4340 & ~n37633;
  assign n37983 = controllable_hmaster0 & ~n37982;
  assign n37984 = ~n6710 & ~n37633;
  assign n37985 = ~controllable_hmaster0 & ~n37984;
  assign n37986 = ~n37983 & ~n37985;
  assign n37987 = controllable_hmaster1 & ~n37986;
  assign n37988 = ~n4340 & ~n37644;
  assign n37989 = controllable_hmaster0 & ~n37988;
  assign n37990 = ~n6947 & ~n37650;
  assign n37991 = ~controllable_hmaster0 & ~n37990;
  assign n37992 = ~n37989 & ~n37991;
  assign n37993 = ~controllable_hmaster1 & ~n37992;
  assign n37994 = ~n37987 & ~n37993;
  assign n37995 = ~i_hbusreq3 & ~n37994;
  assign n37996 = ~n37981 & ~n37995;
  assign n37997 = ~controllable_hmaster2 & ~n37996;
  assign n37998 = ~n37968 & ~n37997;
  assign n37999 = ~controllable_hgrant3 & ~n37998;
  assign n38000 = ~n8810 & ~n37999;
  assign n38001 = controllable_nhgrant0 & ~n38000;
  assign n38002 = ~n8902 & ~n38001;
  assign n38003 = ~n3281 & ~n38002;
  assign n38004 = ~n3950 & ~n38003;
  assign n38005 = ~n3378 & ~n38004;
  assign n38006 = ~n37958 & ~n38005;
  assign n38007 = n3492 & ~n38006;
  assign n38008 = ~n3631 & ~n38007;
  assign n38009 = n3485 & ~n38008;
  assign n38010 = ~n3630 & ~n38009;
  assign n38011 = ~n3476 & ~n38010;
  assign n38012 = n3378 & ~n35921;
  assign n38013 = ~n9477 & ~n37675;
  assign n38014 = controllable_hmaster1 & ~n38013;
  assign n38015 = controllable_hmaster0 & ~n38013;
  assign n38016 = ~n35870 & ~n38015;
  assign n38017 = ~controllable_hmaster1 & ~n38016;
  assign n38018 = ~n38014 & ~n38017;
  assign n38019 = i_hbusreq3 & ~n38018;
  assign n38020 = ~n9485 & ~n37687;
  assign n38021 = controllable_hmaster1 & ~n38020;
  assign n38022 = controllable_hmaster0 & ~n38020;
  assign n38023 = ~n6772 & ~n37694;
  assign n38024 = ~controllable_hmaster0 & ~n38023;
  assign n38025 = ~n38022 & ~n38024;
  assign n38026 = ~controllable_hmaster1 & ~n38025;
  assign n38027 = ~n38021 & ~n38026;
  assign n38028 = ~i_hbusreq3 & ~n38027;
  assign n38029 = ~n38019 & ~n38028;
  assign n38030 = controllable_hmaster2 & ~n38029;
  assign n38031 = ~n6762 & ~n37704;
  assign n38032 = controllable_hmaster0 & ~n38031;
  assign n38033 = ~n6786 & ~n37704;
  assign n38034 = ~controllable_hmaster0 & ~n38033;
  assign n38035 = ~n38032 & ~n38034;
  assign n38036 = controllable_hmaster1 & ~n38035;
  assign n38037 = ~n6762 & ~n37712;
  assign n38038 = controllable_hmaster0 & ~n38037;
  assign n38039 = ~controllable_hmaster0 & ~n38031;
  assign n38040 = ~n38038 & ~n38039;
  assign n38041 = ~controllable_hmaster1 & ~n38040;
  assign n38042 = ~n38036 & ~n38041;
  assign n38043 = i_hbusreq3 & ~n38042;
  assign n38044 = ~n6772 & ~n37724;
  assign n38045 = controllable_hmaster0 & ~n38044;
  assign n38046 = ~n6813 & ~n37724;
  assign n38047 = ~controllable_hmaster0 & ~n38046;
  assign n38048 = ~n38045 & ~n38047;
  assign n38049 = controllable_hmaster1 & ~n38048;
  assign n38050 = ~n6772 & ~n37735;
  assign n38051 = controllable_hmaster0 & ~n38050;
  assign n38052 = ~n6831 & ~n37741;
  assign n38053 = ~controllable_hmaster0 & ~n38052;
  assign n38054 = ~n38051 & ~n38053;
  assign n38055 = ~controllable_hmaster1 & ~n38054;
  assign n38056 = ~n38049 & ~n38055;
  assign n38057 = ~i_hbusreq3 & ~n38056;
  assign n38058 = ~n38043 & ~n38057;
  assign n38059 = ~controllable_hmaster2 & ~n38058;
  assign n38060 = ~n38030 & ~n38059;
  assign n38061 = ~controllable_hgrant3 & ~n38060;
  assign n38062 = ~n8935 & ~n38061;
  assign n38063 = controllable_nhgrant0 & ~n38062;
  assign n38064 = ~n9096 & ~n38063;
  assign n38065 = ~n3281 & ~n38064;
  assign n38066 = ~n4089 & ~n38065;
  assign n38067 = ~n3378 & ~n38066;
  assign n38068 = ~n38012 & ~n38067;
  assign n38069 = n3492 & ~n38068;
  assign n38070 = ~n37132 & ~n38069;
  assign n38071 = n3485 & ~n38070;
  assign n38072 = ~n37313 & ~n38071;
  assign n38073 = n3476 & ~n38072;
  assign n38074 = ~n38011 & ~n38073;
  assign n38075 = n3374 & ~n38074;
  assign n38076 = ~n37957 & ~n38075;
  assign n38077 = ~n3655 & ~n38076;
  assign n38078 = ~n37923 & ~n38077;
  assign n38079 = ~n3652 & ~n38078;
  assign n38080 = ~n37769 & ~n38079;
  assign n38081 = ~n3368 & ~n38080;
  assign n38082 = n3378 & ~n36000;
  assign n38083 = ~n3497 & ~n35937;
  assign n38084 = ~controllable_hgrant2 & ~n38083;
  assign n38085 = ~n3410 & ~n38084;
  assign n38086 = controllable_hmaster1 & ~n38085;
  assign n38087 = controllable_hmaster0 & ~n38085;
  assign n38088 = controllable_hmaster0 & ~n38087;
  assign n38089 = ~controllable_hmaster1 & ~n38088;
  assign n38090 = ~n38086 & ~n38089;
  assign n38091 = i_hbusreq3 & ~n38090;
  assign n38092 = i_hbusreq2 & ~n38083;
  assign n38093 = controllable_hgrant4 & ~n4629;
  assign n38094 = ~n9718 & ~n38093;
  assign n38095 = ~i_hbusreq2 & ~n38094;
  assign n38096 = ~n38092 & ~n38095;
  assign n38097 = ~controllable_hgrant2 & ~n38096;
  assign n38098 = ~n4562 & ~n38097;
  assign n38099 = controllable_hmaster1 & ~n38098;
  assign n38100 = controllable_hmaster0 & ~n38098;
  assign n38101 = controllable_hmaster0 & ~n38100;
  assign n38102 = ~controllable_hmaster1 & ~n38101;
  assign n38103 = ~n38099 & ~n38102;
  assign n38104 = ~i_hbusreq3 & ~n38103;
  assign n38105 = ~n38091 & ~n38104;
  assign n38106 = controllable_hmaster2 & ~n38105;
  assign n38107 = controllable_hmaster2 & ~n38106;
  assign n38108 = ~controllable_hgrant3 & ~n38107;
  assign n38109 = ~n9708 & ~n38108;
  assign n38110 = controllable_nhgrant0 & ~n38109;
  assign n38111 = ~n9753 & ~n38110;
  assign n38112 = ~n3281 & ~n38111;
  assign n38113 = ~n3281 & ~n38112;
  assign n38114 = ~n3378 & ~n38113;
  assign n38115 = ~n38082 & ~n38114;
  assign n38116 = n3492 & ~n38115;
  assign n38117 = n3492 & ~n38116;
  assign n38118 = n3485 & ~n38117;
  assign n38119 = n3485 & ~n38118;
  assign n38120 = ~n3476 & ~n38119;
  assign n38121 = ~n8523 & ~n38116;
  assign n38122 = n3485 & ~n38121;
  assign n38123 = ~n8689 & ~n38122;
  assign n38124 = n3476 & ~n38123;
  assign n38125 = ~n38120 & ~n38124;
  assign n38126 = ~n3374 & ~n38125;
  assign n38127 = n3378 & ~n36132;
  assign n38128 = ~n34637 & ~n38087;
  assign n38129 = ~controllable_hmaster1 & ~n38128;
  assign n38130 = ~n38086 & ~n38129;
  assign n38131 = i_hbusreq3 & ~n38130;
  assign n38132 = ~n34649 & ~n38100;
  assign n38133 = ~controllable_hmaster1 & ~n38132;
  assign n38134 = ~n38099 & ~n38133;
  assign n38135 = ~i_hbusreq3 & ~n38134;
  assign n38136 = ~n38131 & ~n38135;
  assign n38137 = controllable_hmaster2 & ~n38136;
  assign n38138 = ~n3850 & ~n35937;
  assign n38139 = ~controllable_hgrant2 & ~n38138;
  assign n38140 = ~n3410 & ~n38139;
  assign n38141 = controllable_hmaster0 & ~n38140;
  assign n38142 = ~n5288 & ~n38139;
  assign n38143 = ~controllable_hmaster0 & ~n38142;
  assign n38144 = ~n38141 & ~n38143;
  assign n38145 = controllable_hmaster1 & ~n38144;
  assign n38146 = ~n8822 & ~n35937;
  assign n38147 = ~controllable_hgrant2 & ~n38146;
  assign n38148 = ~n3410 & ~n38147;
  assign n38149 = controllable_hmaster0 & ~n38148;
  assign n38150 = ~controllable_hmaster0 & ~n38140;
  assign n38151 = ~n38149 & ~n38150;
  assign n38152 = ~controllable_hmaster1 & ~n38151;
  assign n38153 = ~n38145 & ~n38152;
  assign n38154 = i_hbusreq3 & ~n38153;
  assign n38155 = i_hbusreq2 & ~n38138;
  assign n38156 = ~n4585 & ~n38093;
  assign n38157 = ~i_hbusreq2 & ~n38156;
  assign n38158 = ~n38155 & ~n38157;
  assign n38159 = ~controllable_hgrant2 & ~n38158;
  assign n38160 = ~n4562 & ~n38159;
  assign n38161 = controllable_hmaster0 & ~n38160;
  assign n38162 = ~n9803 & ~n38159;
  assign n38163 = ~controllable_hmaster0 & ~n38162;
  assign n38164 = ~n38161 & ~n38163;
  assign n38165 = controllable_hmaster1 & ~n38164;
  assign n38166 = i_hbusreq2 & ~n38146;
  assign n38167 = ~n9820 & ~n38093;
  assign n38168 = ~i_hbusreq2 & ~n38167;
  assign n38169 = ~n38166 & ~n38168;
  assign n38170 = ~controllable_hgrant2 & ~n38169;
  assign n38171 = ~n4562 & ~n38170;
  assign n38172 = controllable_hmaster0 & ~n38171;
  assign n38173 = ~n38150 & ~n38172;
  assign n38174 = ~controllable_hmaster1 & ~n38173;
  assign n38175 = ~n38165 & ~n38174;
  assign n38176 = ~i_hbusreq3 & ~n38175;
  assign n38177 = ~n38154 & ~n38176;
  assign n38178 = ~controllable_hmaster2 & ~n38177;
  assign n38179 = ~n38137 & ~n38178;
  assign n38180 = ~controllable_hgrant3 & ~n38179;
  assign n38181 = ~n9790 & ~n38180;
  assign n38182 = controllable_nhgrant0 & ~n38181;
  assign n38183 = ~n9861 & ~n38182;
  assign n38184 = ~n3281 & ~n38183;
  assign n38185 = ~n3281 & ~n38184;
  assign n38186 = ~n3378 & ~n38185;
  assign n38187 = ~n38127 & ~n38186;
  assign n38188 = n3492 & ~n38187;
  assign n38189 = n3492 & ~n38188;
  assign n38190 = n3485 & ~n38189;
  assign n38191 = n3485 & ~n38190;
  assign n38192 = ~n3476 & ~n38191;
  assign n38193 = ~n9873 & ~n36143;
  assign n38194 = ~controllable_hgrant2 & ~n38193;
  assign n38195 = ~n5616 & ~n38194;
  assign n38196 = controllable_hmaster1 & ~n38195;
  assign n38197 = controllable_hmaster0 & ~n38195;
  assign n38198 = ~n5621 & ~n34682;
  assign n38199 = ~controllable_hgrant2 & ~n38198;
  assign n38200 = ~n5616 & ~n38199;
  assign n38201 = ~controllable_hmaster0 & ~n38200;
  assign n38202 = ~n38197 & ~n38201;
  assign n38203 = ~controllable_hmaster1 & ~n38202;
  assign n38204 = ~n38196 & ~n38203;
  assign n38205 = i_hbusreq3 & ~n38204;
  assign n38206 = i_hbusreq2 & ~n38193;
  assign n38207 = ~n9895 & ~n36254;
  assign n38208 = ~i_hbusreq2 & ~n38207;
  assign n38209 = ~n38206 & ~n38208;
  assign n38210 = ~controllable_hgrant2 & ~n38209;
  assign n38211 = ~n5862 & ~n38210;
  assign n38212 = controllable_hmaster1 & ~n38211;
  assign n38213 = controllable_hmaster0 & ~n38211;
  assign n38214 = i_hbusreq2 & ~n38198;
  assign n38215 = ~n9910 & ~n34712;
  assign n38216 = ~i_hbusreq2 & ~n38215;
  assign n38217 = ~n38214 & ~n38216;
  assign n38218 = ~controllable_hgrant2 & ~n38217;
  assign n38219 = ~n7507 & ~n38218;
  assign n38220 = ~controllable_hmaster0 & ~n38219;
  assign n38221 = ~n38213 & ~n38220;
  assign n38222 = ~controllable_hmaster1 & ~n38221;
  assign n38223 = ~n38212 & ~n38222;
  assign n38224 = ~i_hbusreq3 & ~n38223;
  assign n38225 = ~n38205 & ~n38224;
  assign n38226 = controllable_hmaster2 & ~n38225;
  assign n38227 = ~n5911 & ~n36143;
  assign n38228 = ~controllable_hgrant2 & ~n38227;
  assign n38229 = ~n5616 & ~n38228;
  assign n38230 = controllable_hmaster0 & ~n38229;
  assign n38231 = ~n5686 & ~n38228;
  assign n38232 = ~controllable_hmaster0 & ~n38231;
  assign n38233 = ~n38230 & ~n38232;
  assign n38234 = controllable_hmaster1 & ~n38233;
  assign n38235 = ~n5921 & ~n36143;
  assign n38236 = ~controllable_hgrant2 & ~n38235;
  assign n38237 = ~n5616 & ~n38236;
  assign n38238 = controllable_hmaster0 & ~n38237;
  assign n38239 = ~controllable_hmaster0 & ~n38229;
  assign n38240 = ~n38238 & ~n38239;
  assign n38241 = ~controllable_hmaster1 & ~n38240;
  assign n38242 = ~n38234 & ~n38241;
  assign n38243 = i_hbusreq3 & ~n38242;
  assign n38244 = i_hbusreq2 & ~n38227;
  assign n38245 = ~n5943 & ~n36254;
  assign n38246 = ~i_hbusreq2 & ~n38245;
  assign n38247 = ~n38244 & ~n38246;
  assign n38248 = ~controllable_hgrant2 & ~n38247;
  assign n38249 = ~n5862 & ~n38248;
  assign n38250 = controllable_hmaster0 & ~n38249;
  assign n38251 = ~n5950 & ~n38248;
  assign n38252 = ~controllable_hmaster0 & ~n38251;
  assign n38253 = ~n38250 & ~n38252;
  assign n38254 = controllable_hmaster1 & ~n38253;
  assign n38255 = i_hbusreq2 & ~n38235;
  assign n38256 = ~n5974 & ~n36254;
  assign n38257 = ~i_hbusreq2 & ~n38256;
  assign n38258 = ~n38255 & ~n38257;
  assign n38259 = ~controllable_hgrant2 & ~n38258;
  assign n38260 = ~n5862 & ~n38259;
  assign n38261 = controllable_hmaster0 & ~n38260;
  assign n38262 = ~n5990 & ~n36315;
  assign n38263 = ~i_hbusreq2 & ~n38262;
  assign n38264 = ~n38244 & ~n38263;
  assign n38265 = ~controllable_hgrant2 & ~n38264;
  assign n38266 = ~n5981 & ~n38265;
  assign n38267 = ~controllable_hmaster0 & ~n38266;
  assign n38268 = ~n38261 & ~n38267;
  assign n38269 = ~controllable_hmaster1 & ~n38268;
  assign n38270 = ~n38254 & ~n38269;
  assign n38271 = ~i_hbusreq3 & ~n38270;
  assign n38272 = ~n38243 & ~n38271;
  assign n38273 = ~controllable_hmaster2 & ~n38272;
  assign n38274 = ~n38226 & ~n38273;
  assign n38275 = ~controllable_hgrant3 & ~n38274;
  assign n38276 = ~n7457 & ~n38275;
  assign n38277 = controllable_nhgrant0 & ~n38276;
  assign n38278 = ~n10071 & ~n38277;
  assign n38279 = ~n3281 & ~n38278;
  assign n38280 = ~n3281 & ~n38279;
  assign n38281 = n3378 & ~n38280;
  assign n38282 = ~n5621 & ~n36143;
  assign n38283 = ~controllable_hgrant2 & ~n38282;
  assign n38284 = ~n5616 & ~n38283;
  assign n38285 = controllable_hmaster1 & ~n38284;
  assign n38286 = controllable_hmaster0 & ~n38284;
  assign n38287 = ~n38201 & ~n38286;
  assign n38288 = ~controllable_hmaster1 & ~n38287;
  assign n38289 = ~n38285 & ~n38288;
  assign n38290 = i_hbusreq3 & ~n38289;
  assign n38291 = i_hbusreq2 & ~n38282;
  assign n38292 = i_hlock4 & ~n11030;
  assign n38293 = ~i_hlock4 & ~n11040;
  assign n38294 = ~n38292 & ~n38293;
  assign n38295 = ~i_hbusreq4 & ~n38294;
  assign n38296 = ~n36158 & ~n38295;
  assign n38297 = controllable_hgrant4 & ~n38296;
  assign n38298 = ~n10120 & ~n38297;
  assign n38299 = ~i_hbusreq2 & ~n38298;
  assign n38300 = ~n38291 & ~n38299;
  assign n38301 = ~controllable_hgrant2 & ~n38300;
  assign n38302 = ~n10111 & ~n38301;
  assign n38303 = controllable_hmaster1 & ~n38302;
  assign n38304 = controllable_hmaster0 & ~n38302;
  assign n38305 = ~n10133 & ~n34712;
  assign n38306 = ~i_hbusreq2 & ~n38305;
  assign n38307 = ~n38214 & ~n38306;
  assign n38308 = ~controllable_hgrant2 & ~n38307;
  assign n38309 = ~n10111 & ~n38308;
  assign n38310 = ~controllable_hmaster0 & ~n38309;
  assign n38311 = ~n38304 & ~n38310;
  assign n38312 = ~controllable_hmaster1 & ~n38311;
  assign n38313 = ~n38303 & ~n38312;
  assign n38314 = ~i_hbusreq3 & ~n38313;
  assign n38315 = ~n38290 & ~n38314;
  assign n38316 = controllable_hmaster2 & ~n38315;
  assign n38317 = ~n5686 & ~n38283;
  assign n38318 = ~controllable_hmaster0 & ~n38317;
  assign n38319 = ~n38286 & ~n38318;
  assign n38320 = controllable_hmaster1 & ~n38319;
  assign n38321 = ~n8987 & ~n36143;
  assign n38322 = ~controllable_hgrant2 & ~n38321;
  assign n38323 = ~n5616 & ~n38322;
  assign n38324 = controllable_hmaster0 & ~n38323;
  assign n38325 = ~controllable_hmaster0 & ~n38284;
  assign n38326 = ~n38324 & ~n38325;
  assign n38327 = ~controllable_hmaster1 & ~n38326;
  assign n38328 = ~n38320 & ~n38327;
  assign n38329 = i_hbusreq3 & ~n38328;
  assign n38330 = ~n10133 & ~n38297;
  assign n38331 = ~i_hbusreq2 & ~n38330;
  assign n38332 = ~n38291 & ~n38331;
  assign n38333 = ~controllable_hgrant2 & ~n38332;
  assign n38334 = ~n10111 & ~n38333;
  assign n38335 = controllable_hmaster0 & ~n38334;
  assign n38336 = ~n10152 & ~n38333;
  assign n38337 = ~controllable_hmaster0 & ~n38336;
  assign n38338 = ~n38335 & ~n38337;
  assign n38339 = controllable_hmaster1 & ~n38338;
  assign n38340 = i_hbusreq2 & ~n38321;
  assign n38341 = ~n10169 & ~n38297;
  assign n38342 = ~i_hbusreq2 & ~n38341;
  assign n38343 = ~n38340 & ~n38342;
  assign n38344 = ~controllable_hgrant2 & ~n38343;
  assign n38345 = ~n10111 & ~n38344;
  assign n38346 = controllable_hmaster0 & ~n38345;
  assign n38347 = i_hlock4 & ~n11118;
  assign n38348 = ~n36141 & ~n38347;
  assign n38349 = ~i_hbusreq4 & ~n38348;
  assign n38350 = ~n36158 & ~n38349;
  assign n38351 = controllable_hgrant4 & ~n38350;
  assign n38352 = ~n10180 & ~n38351;
  assign n38353 = ~i_hbusreq2 & ~n38352;
  assign n38354 = ~n38291 & ~n38353;
  assign n38355 = ~controllable_hgrant2 & ~n38354;
  assign n38356 = ~n5616 & ~n38355;
  assign n38357 = ~controllable_hmaster0 & ~n38356;
  assign n38358 = ~n38346 & ~n38357;
  assign n38359 = ~controllable_hmaster1 & ~n38358;
  assign n38360 = ~n38339 & ~n38359;
  assign n38361 = ~i_hbusreq3 & ~n38360;
  assign n38362 = ~n38329 & ~n38361;
  assign n38363 = ~controllable_hmaster2 & ~n38362;
  assign n38364 = ~n38316 & ~n38363;
  assign n38365 = ~controllable_hgrant3 & ~n38364;
  assign n38366 = ~n10110 & ~n38365;
  assign n38367 = controllable_nhgrant0 & ~n38366;
  assign n38368 = ~n10240 & ~n38367;
  assign n38369 = ~n3281 & ~n38368;
  assign n38370 = ~n3281 & ~n38369;
  assign n38371 = ~n3378 & ~n38370;
  assign n38372 = ~n38281 & ~n38371;
  assign n38373 = n3492 & ~n38372;
  assign n38374 = ~n37174 & ~n38373;
  assign n38375 = n3485 & ~n38374;
  assign n38376 = ~n37332 & ~n38375;
  assign n38377 = n3476 & ~n38376;
  assign n38378 = ~n38192 & ~n38377;
  assign n38379 = n3374 & ~n38378;
  assign n38380 = ~n38126 & ~n38379;
  assign n38381 = n3655 & ~n38380;
  assign n38382 = n3378 & ~n36375;
  assign n38383 = ~n10257 & ~n35937;
  assign n38384 = ~controllable_hgrant2 & ~n38383;
  assign n38385 = ~n3410 & ~n38384;
  assign n38386 = controllable_hmaster1 & ~n38385;
  assign n38387 = controllable_hmaster0 & ~n38385;
  assign n38388 = controllable_hmaster0 & ~n38387;
  assign n38389 = ~controllable_hmaster1 & ~n38388;
  assign n38390 = ~n38386 & ~n38389;
  assign n38391 = i_hbusreq3 & ~n38390;
  assign n38392 = i_hbusreq2 & ~n38383;
  assign n38393 = ~n10278 & ~n38093;
  assign n38394 = ~i_hbusreq2 & ~n38393;
  assign n38395 = ~n38392 & ~n38394;
  assign n38396 = ~controllable_hgrant2 & ~n38395;
  assign n38397 = ~n4562 & ~n38396;
  assign n38398 = controllable_hmaster1 & ~n38397;
  assign n38399 = controllable_hmaster0 & ~n38397;
  assign n38400 = controllable_hmaster0 & ~n38399;
  assign n38401 = ~controllable_hmaster1 & ~n38400;
  assign n38402 = ~n38398 & ~n38401;
  assign n38403 = ~i_hbusreq3 & ~n38402;
  assign n38404 = ~n38391 & ~n38403;
  assign n38405 = controllable_hmaster2 & ~n38404;
  assign n38406 = controllable_hmaster2 & ~n38405;
  assign n38407 = ~controllable_hgrant3 & ~n38406;
  assign n38408 = ~n9708 & ~n38407;
  assign n38409 = controllable_nhgrant0 & ~n38408;
  assign n38410 = ~n9753 & ~n38409;
  assign n38411 = ~n3281 & ~n38410;
  assign n38412 = ~n3281 & ~n38411;
  assign n38413 = ~n3378 & ~n38412;
  assign n38414 = ~n38382 & ~n38413;
  assign n38415 = n3492 & ~n38414;
  assign n38416 = n3492 & ~n38415;
  assign n38417 = n3485 & ~n38416;
  assign n38418 = n3485 & ~n38417;
  assign n38419 = ~n3476 & ~n38418;
  assign n38420 = ~n8523 & ~n38415;
  assign n38421 = n3485 & ~n38420;
  assign n38422 = ~n8689 & ~n38421;
  assign n38423 = n3476 & ~n38422;
  assign n38424 = ~n38419 & ~n38423;
  assign n38425 = ~n3374 & ~n38424;
  assign n38426 = n3378 & ~n36464;
  assign n38427 = ~n34748 & ~n38387;
  assign n38428 = ~controllable_hmaster1 & ~n38427;
  assign n38429 = ~n38386 & ~n38428;
  assign n38430 = i_hbusreq3 & ~n38429;
  assign n38431 = ~n34759 & ~n38399;
  assign n38432 = ~controllable_hmaster1 & ~n38431;
  assign n38433 = ~n38398 & ~n38432;
  assign n38434 = ~i_hbusreq3 & ~n38433;
  assign n38435 = ~n38430 & ~n38434;
  assign n38436 = controllable_hmaster2 & ~n38435;
  assign n38437 = ~n4701 & ~n35937;
  assign n38438 = ~controllable_hgrant2 & ~n38437;
  assign n38439 = ~n3410 & ~n38438;
  assign n38440 = controllable_hmaster0 & ~n38439;
  assign n38441 = ~n5288 & ~n38438;
  assign n38442 = ~controllable_hmaster0 & ~n38441;
  assign n38443 = ~n38440 & ~n38442;
  assign n38444 = controllable_hmaster1 & ~n38443;
  assign n38445 = ~n10332 & ~n35937;
  assign n38446 = ~controllable_hgrant2 & ~n38445;
  assign n38447 = ~n3410 & ~n38446;
  assign n38448 = controllable_hmaster0 & ~n38447;
  assign n38449 = ~controllable_hmaster0 & ~n38439;
  assign n38450 = ~n38448 & ~n38449;
  assign n38451 = ~controllable_hmaster1 & ~n38450;
  assign n38452 = ~n38444 & ~n38451;
  assign n38453 = i_hbusreq3 & ~n38452;
  assign n38454 = i_hbusreq2 & ~n38437;
  assign n38455 = ~n4723 & ~n38093;
  assign n38456 = ~i_hbusreq2 & ~n38455;
  assign n38457 = ~n38454 & ~n38456;
  assign n38458 = ~controllable_hgrant2 & ~n38457;
  assign n38459 = ~n4562 & ~n38458;
  assign n38460 = controllable_hmaster0 & ~n38459;
  assign n38461 = ~n9803 & ~n38458;
  assign n38462 = ~controllable_hmaster0 & ~n38461;
  assign n38463 = ~n38460 & ~n38462;
  assign n38464 = controllable_hmaster1 & ~n38463;
  assign n38465 = i_hbusreq2 & ~n38445;
  assign n38466 = ~n10370 & ~n38093;
  assign n38467 = ~i_hbusreq2 & ~n38466;
  assign n38468 = ~n38465 & ~n38467;
  assign n38469 = ~controllable_hgrant2 & ~n38468;
  assign n38470 = ~n4562 & ~n38469;
  assign n38471 = controllable_hmaster0 & ~n38470;
  assign n38472 = ~n38449 & ~n38471;
  assign n38473 = ~controllable_hmaster1 & ~n38472;
  assign n38474 = ~n38464 & ~n38473;
  assign n38475 = ~i_hbusreq3 & ~n38474;
  assign n38476 = ~n38453 & ~n38475;
  assign n38477 = ~controllable_hmaster2 & ~n38476;
  assign n38478 = ~n38436 & ~n38477;
  assign n38479 = ~controllable_hgrant3 & ~n38478;
  assign n38480 = ~n9790 & ~n38479;
  assign n38481 = controllable_nhgrant0 & ~n38480;
  assign n38482 = ~n9861 & ~n38481;
  assign n38483 = ~n3281 & ~n38482;
  assign n38484 = ~n3281 & ~n38483;
  assign n38485 = ~n3378 & ~n38484;
  assign n38486 = ~n38426 & ~n38485;
  assign n38487 = n3492 & ~n38486;
  assign n38488 = n3492 & ~n38487;
  assign n38489 = n3485 & ~n38488;
  assign n38490 = n3485 & ~n38489;
  assign n38491 = ~n3476 & ~n38490;
  assign n38492 = ~n10404 & ~n36143;
  assign n38493 = ~controllable_hgrant2 & ~n38492;
  assign n38494 = ~n5616 & ~n38493;
  assign n38495 = controllable_hmaster1 & ~n38494;
  assign n38496 = controllable_hmaster0 & ~n38494;
  assign n38497 = ~n10412 & ~n34682;
  assign n38498 = ~controllable_hgrant2 & ~n38497;
  assign n38499 = ~n5616 & ~n38498;
  assign n38500 = ~controllable_hmaster0 & ~n38499;
  assign n38501 = ~n38496 & ~n38500;
  assign n38502 = ~controllable_hmaster1 & ~n38501;
  assign n38503 = ~n38495 & ~n38502;
  assign n38504 = i_hbusreq3 & ~n38503;
  assign n38505 = i_hbusreq2 & ~n38492;
  assign n38506 = ~n10443 & ~n36254;
  assign n38507 = ~i_hbusreq2 & ~n38506;
  assign n38508 = ~n38505 & ~n38507;
  assign n38509 = ~controllable_hgrant2 & ~n38508;
  assign n38510 = ~n5862 & ~n38509;
  assign n38511 = controllable_hmaster1 & ~n38510;
  assign n38512 = controllable_hmaster0 & ~n38510;
  assign n38513 = i_hbusreq2 & ~n38497;
  assign n38514 = ~n10468 & ~n34712;
  assign n38515 = ~i_hbusreq2 & ~n38514;
  assign n38516 = ~n38513 & ~n38515;
  assign n38517 = ~controllable_hgrant2 & ~n38516;
  assign n38518 = ~n7507 & ~n38517;
  assign n38519 = ~controllable_hmaster0 & ~n38518;
  assign n38520 = ~n38512 & ~n38519;
  assign n38521 = ~controllable_hmaster1 & ~n38520;
  assign n38522 = ~n38511 & ~n38521;
  assign n38523 = ~i_hbusreq3 & ~n38522;
  assign n38524 = ~n38504 & ~n38523;
  assign n38525 = controllable_hmaster2 & ~n38524;
  assign n38526 = ~n10483 & ~n36143;
  assign n38527 = ~controllable_hgrant2 & ~n38526;
  assign n38528 = ~n5616 & ~n38527;
  assign n38529 = controllable_hmaster0 & ~n38528;
  assign n38530 = ~n5686 & ~n38527;
  assign n38531 = ~controllable_hmaster0 & ~n38530;
  assign n38532 = ~n38529 & ~n38531;
  assign n38533 = controllable_hmaster1 & ~n38532;
  assign n38534 = ~n10498 & ~n36143;
  assign n38535 = ~controllable_hgrant2 & ~n38534;
  assign n38536 = ~n5616 & ~n38535;
  assign n38537 = controllable_hmaster0 & ~n38536;
  assign n38538 = ~controllable_hmaster0 & ~n38528;
  assign n38539 = ~n38537 & ~n38538;
  assign n38540 = ~controllable_hmaster1 & ~n38539;
  assign n38541 = ~n38533 & ~n38540;
  assign n38542 = i_hbusreq3 & ~n38541;
  assign n38543 = i_hbusreq2 & ~n38526;
  assign n38544 = ~n10521 & ~n36254;
  assign n38545 = ~i_hbusreq2 & ~n38544;
  assign n38546 = ~n38543 & ~n38545;
  assign n38547 = ~controllable_hgrant2 & ~n38546;
  assign n38548 = ~n5862 & ~n38547;
  assign n38549 = controllable_hmaster0 & ~n38548;
  assign n38550 = ~n5950 & ~n38547;
  assign n38551 = ~controllable_hmaster0 & ~n38550;
  assign n38552 = ~n38549 & ~n38551;
  assign n38553 = controllable_hmaster1 & ~n38552;
  assign n38554 = i_hbusreq2 & ~n38534;
  assign n38555 = ~n10552 & ~n36254;
  assign n38556 = ~i_hbusreq2 & ~n38555;
  assign n38557 = ~n38554 & ~n38556;
  assign n38558 = ~controllable_hgrant2 & ~n38557;
  assign n38559 = ~n5862 & ~n38558;
  assign n38560 = controllable_hmaster0 & ~n38559;
  assign n38561 = ~n10567 & ~n36315;
  assign n38562 = ~i_hbusreq2 & ~n38561;
  assign n38563 = ~n38543 & ~n38562;
  assign n38564 = ~controllable_hgrant2 & ~n38563;
  assign n38565 = ~n5981 & ~n38564;
  assign n38566 = ~controllable_hmaster0 & ~n38565;
  assign n38567 = ~n38560 & ~n38566;
  assign n38568 = ~controllable_hmaster1 & ~n38567;
  assign n38569 = ~n38553 & ~n38568;
  assign n38570 = ~i_hbusreq3 & ~n38569;
  assign n38571 = ~n38542 & ~n38570;
  assign n38572 = ~controllable_hmaster2 & ~n38571;
  assign n38573 = ~n38525 & ~n38572;
  assign n38574 = ~controllable_hgrant3 & ~n38573;
  assign n38575 = ~n7457 & ~n38574;
  assign n38576 = controllable_nhgrant0 & ~n38575;
  assign n38577 = ~n10071 & ~n38576;
  assign n38578 = ~n3281 & ~n38577;
  assign n38579 = ~n3281 & ~n38578;
  assign n38580 = n3378 & ~n38579;
  assign n38581 = ~n10412 & ~n36143;
  assign n38582 = ~controllable_hgrant2 & ~n38581;
  assign n38583 = ~n5616 & ~n38582;
  assign n38584 = controllable_hmaster1 & ~n38583;
  assign n38585 = controllable_hmaster0 & ~n38583;
  assign n38586 = ~n38500 & ~n38585;
  assign n38587 = ~controllable_hmaster1 & ~n38586;
  assign n38588 = ~n38584 & ~n38587;
  assign n38589 = i_hbusreq3 & ~n38588;
  assign n38590 = i_hbusreq2 & ~n38581;
  assign n38591 = ~n10607 & ~n38297;
  assign n38592 = ~i_hbusreq2 & ~n38591;
  assign n38593 = ~n38590 & ~n38592;
  assign n38594 = ~controllable_hgrant2 & ~n38593;
  assign n38595 = ~n10111 & ~n38594;
  assign n38596 = controllable_hmaster1 & ~n38595;
  assign n38597 = controllable_hmaster0 & ~n38595;
  assign n38598 = ~n10620 & ~n34712;
  assign n38599 = ~i_hbusreq2 & ~n38598;
  assign n38600 = ~n38513 & ~n38599;
  assign n38601 = ~controllable_hgrant2 & ~n38600;
  assign n38602 = ~n10111 & ~n38601;
  assign n38603 = ~controllable_hmaster0 & ~n38602;
  assign n38604 = ~n38597 & ~n38603;
  assign n38605 = ~controllable_hmaster1 & ~n38604;
  assign n38606 = ~n38596 & ~n38605;
  assign n38607 = ~i_hbusreq3 & ~n38606;
  assign n38608 = ~n38589 & ~n38607;
  assign n38609 = controllable_hmaster2 & ~n38608;
  assign n38610 = ~n5686 & ~n38582;
  assign n38611 = ~controllable_hmaster0 & ~n38610;
  assign n38612 = ~n38585 & ~n38611;
  assign n38613 = controllable_hmaster1 & ~n38612;
  assign n38614 = ~n10638 & ~n36143;
  assign n38615 = ~controllable_hgrant2 & ~n38614;
  assign n38616 = ~n5616 & ~n38615;
  assign n38617 = controllable_hmaster0 & ~n38616;
  assign n38618 = ~controllable_hmaster0 & ~n38583;
  assign n38619 = ~n38617 & ~n38618;
  assign n38620 = ~controllable_hmaster1 & ~n38619;
  assign n38621 = ~n38613 & ~n38620;
  assign n38622 = i_hbusreq3 & ~n38621;
  assign n38623 = ~n10620 & ~n38297;
  assign n38624 = ~i_hbusreq2 & ~n38623;
  assign n38625 = ~n38590 & ~n38624;
  assign n38626 = ~controllable_hgrant2 & ~n38625;
  assign n38627 = ~n10111 & ~n38626;
  assign n38628 = controllable_hmaster0 & ~n38627;
  assign n38629 = ~n10152 & ~n38626;
  assign n38630 = ~controllable_hmaster0 & ~n38629;
  assign n38631 = ~n38628 & ~n38630;
  assign n38632 = controllable_hmaster1 & ~n38631;
  assign n38633 = i_hbusreq2 & ~n38614;
  assign n38634 = ~n10674 & ~n38297;
  assign n38635 = ~i_hbusreq2 & ~n38634;
  assign n38636 = ~n38633 & ~n38635;
  assign n38637 = ~controllable_hgrant2 & ~n38636;
  assign n38638 = ~n10111 & ~n38637;
  assign n38639 = controllable_hmaster0 & ~n38638;
  assign n38640 = ~n10685 & ~n38351;
  assign n38641 = ~i_hbusreq2 & ~n38640;
  assign n38642 = ~n38590 & ~n38641;
  assign n38643 = ~controllable_hgrant2 & ~n38642;
  assign n38644 = ~n5616 & ~n38643;
  assign n38645 = ~controllable_hmaster0 & ~n38644;
  assign n38646 = ~n38639 & ~n38645;
  assign n38647 = ~controllable_hmaster1 & ~n38646;
  assign n38648 = ~n38632 & ~n38647;
  assign n38649 = ~i_hbusreq3 & ~n38648;
  assign n38650 = ~n38622 & ~n38649;
  assign n38651 = ~controllable_hmaster2 & ~n38650;
  assign n38652 = ~n38609 & ~n38651;
  assign n38653 = ~controllable_hgrant3 & ~n38652;
  assign n38654 = ~n10110 & ~n38653;
  assign n38655 = controllable_nhgrant0 & ~n38654;
  assign n38656 = ~n10240 & ~n38655;
  assign n38657 = ~n3281 & ~n38656;
  assign n38658 = ~n3281 & ~n38657;
  assign n38659 = ~n3378 & ~n38658;
  assign n38660 = ~n38580 & ~n38659;
  assign n38661 = n3492 & ~n38660;
  assign n38662 = ~n37202 & ~n38661;
  assign n38663 = n3485 & ~n38662;
  assign n38664 = ~n37343 & ~n38663;
  assign n38665 = n3476 & ~n38664;
  assign n38666 = ~n38491 & ~n38665;
  assign n38667 = n3374 & ~n38666;
  assign n38668 = ~n38425 & ~n38667;
  assign n38669 = ~n3655 & ~n38668;
  assign n38670 = ~n38381 & ~n38669;
  assign n38671 = n3652 & ~n38670;
  assign n38672 = n3378 & ~n36624;
  assign n38673 = ~n4787 & ~n38084;
  assign n38674 = controllable_hmaster1 & ~n38673;
  assign n38675 = controllable_hmaster0 & ~n38673;
  assign n38676 = controllable_hmaster0 & ~n38675;
  assign n38677 = ~controllable_hmaster1 & ~n38676;
  assign n38678 = ~n38674 & ~n38677;
  assign n38679 = i_hbusreq3 & ~n38678;
  assign n38680 = ~n4794 & ~n38097;
  assign n38681 = controllable_hmaster1 & ~n38680;
  assign n38682 = controllable_hmaster0 & ~n38680;
  assign n38683 = controllable_hmaster0 & ~n38682;
  assign n38684 = ~controllable_hmaster1 & ~n38683;
  assign n38685 = ~n38681 & ~n38684;
  assign n38686 = ~i_hbusreq3 & ~n38685;
  assign n38687 = ~n38679 & ~n38686;
  assign n38688 = controllable_hmaster2 & ~n38687;
  assign n38689 = controllable_hmaster2 & ~n38688;
  assign n38690 = ~controllable_hgrant3 & ~n38689;
  assign n38691 = ~n9708 & ~n38690;
  assign n38692 = controllable_nhgrant0 & ~n38691;
  assign n38693 = ~n9753 & ~n38692;
  assign n38694 = ~n3281 & ~n38693;
  assign n38695 = ~n3281 & ~n38694;
  assign n38696 = ~n3378 & ~n38695;
  assign n38697 = ~n38672 & ~n38696;
  assign n38698 = n3492 & ~n38697;
  assign n38699 = n3492 & ~n38698;
  assign n38700 = n3485 & ~n38699;
  assign n38701 = n3485 & ~n38700;
  assign n38702 = ~n3476 & ~n38701;
  assign n38703 = ~n8523 & ~n38698;
  assign n38704 = n3485 & ~n38703;
  assign n38705 = ~n8689 & ~n38704;
  assign n38706 = n3476 & ~n38705;
  assign n38707 = ~n38702 & ~n38706;
  assign n38708 = ~n3374 & ~n38707;
  assign n38709 = n3378 & ~n36695;
  assign n38710 = ~n34818 & ~n38675;
  assign n38711 = ~controllable_hmaster1 & ~n38710;
  assign n38712 = ~n38674 & ~n38711;
  assign n38713 = i_hbusreq3 & ~n38712;
  assign n38714 = ~n34824 & ~n38682;
  assign n38715 = ~controllable_hmaster1 & ~n38714;
  assign n38716 = ~n38681 & ~n38715;
  assign n38717 = ~i_hbusreq3 & ~n38716;
  assign n38718 = ~n38713 & ~n38717;
  assign n38719 = controllable_hmaster2 & ~n38718;
  assign n38720 = ~n4787 & ~n38139;
  assign n38721 = controllable_hmaster0 & ~n38720;
  assign n38722 = ~n10768 & ~n38139;
  assign n38723 = ~controllable_hmaster0 & ~n38722;
  assign n38724 = ~n38721 & ~n38723;
  assign n38725 = controllable_hmaster1 & ~n38724;
  assign n38726 = ~n4787 & ~n38147;
  assign n38727 = controllable_hmaster0 & ~n38726;
  assign n38728 = ~controllable_hmaster0 & ~n38720;
  assign n38729 = ~n38727 & ~n38728;
  assign n38730 = ~controllable_hmaster1 & ~n38729;
  assign n38731 = ~n38725 & ~n38730;
  assign n38732 = i_hbusreq3 & ~n38731;
  assign n38733 = ~n4794 & ~n38159;
  assign n38734 = controllable_hmaster0 & ~n38733;
  assign n38735 = ~n10782 & ~n38159;
  assign n38736 = ~controllable_hmaster0 & ~n38735;
  assign n38737 = ~n38734 & ~n38736;
  assign n38738 = controllable_hmaster1 & ~n38737;
  assign n38739 = ~n4794 & ~n38170;
  assign n38740 = controllable_hmaster0 & ~n38739;
  assign n38741 = ~n38728 & ~n38740;
  assign n38742 = ~controllable_hmaster1 & ~n38741;
  assign n38743 = ~n38738 & ~n38742;
  assign n38744 = ~i_hbusreq3 & ~n38743;
  assign n38745 = ~n38732 & ~n38744;
  assign n38746 = ~controllable_hmaster2 & ~n38745;
  assign n38747 = ~n38719 & ~n38746;
  assign n38748 = ~controllable_hgrant3 & ~n38747;
  assign n38749 = ~n9790 & ~n38748;
  assign n38750 = controllable_nhgrant0 & ~n38749;
  assign n38751 = ~n9861 & ~n38750;
  assign n38752 = ~n3281 & ~n38751;
  assign n38753 = ~n3281 & ~n38752;
  assign n38754 = ~n3378 & ~n38753;
  assign n38755 = ~n38709 & ~n38754;
  assign n38756 = n3492 & ~n38755;
  assign n38757 = n3492 & ~n38756;
  assign n38758 = n3485 & ~n38757;
  assign n38759 = n3485 & ~n38758;
  assign n38760 = ~n3476 & ~n38759;
  assign n38761 = ~n10816 & ~n38194;
  assign n38762 = controllable_hmaster1 & ~n38761;
  assign n38763 = controllable_hmaster0 & ~n38761;
  assign n38764 = ~n10827 & ~n38199;
  assign n38765 = ~controllable_hmaster0 & ~n38764;
  assign n38766 = ~n38763 & ~n38765;
  assign n38767 = ~controllable_hmaster1 & ~n38766;
  assign n38768 = ~n38762 & ~n38767;
  assign n38769 = i_hbusreq3 & ~n38768;
  assign n38770 = ~n10870 & ~n38210;
  assign n38771 = controllable_hmaster1 & ~n38770;
  assign n38772 = controllable_hmaster0 & ~n38770;
  assign n38773 = ~n10904 & ~n38218;
  assign n38774 = ~controllable_hmaster0 & ~n38773;
  assign n38775 = ~n38772 & ~n38774;
  assign n38776 = ~controllable_hmaster1 & ~n38775;
  assign n38777 = ~n38771 & ~n38776;
  assign n38778 = ~i_hbusreq3 & ~n38777;
  assign n38779 = ~n38769 & ~n38778;
  assign n38780 = controllable_hmaster2 & ~n38779;
  assign n38781 = ~n10816 & ~n38228;
  assign n38782 = controllable_hmaster0 & ~n38781;
  assign n38783 = ~n10922 & ~n38228;
  assign n38784 = ~controllable_hmaster0 & ~n38783;
  assign n38785 = ~n38782 & ~n38784;
  assign n38786 = controllable_hmaster1 & ~n38785;
  assign n38787 = ~n10816 & ~n38236;
  assign n38788 = controllable_hmaster0 & ~n38787;
  assign n38789 = ~controllable_hmaster0 & ~n38781;
  assign n38790 = ~n38788 & ~n38789;
  assign n38791 = ~controllable_hmaster1 & ~n38790;
  assign n38792 = ~n38786 & ~n38791;
  assign n38793 = i_hbusreq3 & ~n38792;
  assign n38794 = ~n10870 & ~n38248;
  assign n38795 = controllable_hmaster0 & ~n38794;
  assign n38796 = ~n10972 & ~n38248;
  assign n38797 = ~controllable_hmaster0 & ~n38796;
  assign n38798 = ~n38795 & ~n38797;
  assign n38799 = controllable_hmaster1 & ~n38798;
  assign n38800 = ~n10870 & ~n38259;
  assign n38801 = controllable_hmaster0 & ~n38800;
  assign n38802 = ~n11002 & ~n38265;
  assign n38803 = ~controllable_hmaster0 & ~n38802;
  assign n38804 = ~n38801 & ~n38803;
  assign n38805 = ~controllable_hmaster1 & ~n38804;
  assign n38806 = ~n38799 & ~n38805;
  assign n38807 = ~i_hbusreq3 & ~n38806;
  assign n38808 = ~n38793 & ~n38807;
  assign n38809 = ~controllable_hmaster2 & ~n38808;
  assign n38810 = ~n38780 & ~n38809;
  assign n38811 = ~controllable_hgrant3 & ~n38810;
  assign n38812 = ~n7457 & ~n38811;
  assign n38813 = controllable_nhgrant0 & ~n38812;
  assign n38814 = ~n10071 & ~n38813;
  assign n38815 = ~n3281 & ~n38814;
  assign n38816 = ~n3281 & ~n38815;
  assign n38817 = n3378 & ~n38816;
  assign n38818 = ~n10827 & ~n38283;
  assign n38819 = controllable_hmaster1 & ~n38818;
  assign n38820 = controllable_hmaster0 & ~n38818;
  assign n38821 = ~n38765 & ~n38820;
  assign n38822 = ~controllable_hmaster1 & ~n38821;
  assign n38823 = ~n38819 & ~n38822;
  assign n38824 = i_hbusreq3 & ~n38823;
  assign n38825 = ~n11049 & ~n38301;
  assign n38826 = controllable_hmaster1 & ~n38825;
  assign n38827 = controllable_hmaster0 & ~n38825;
  assign n38828 = ~n11049 & ~n38308;
  assign n38829 = ~controllable_hmaster0 & ~n38828;
  assign n38830 = ~n38827 & ~n38829;
  assign n38831 = ~controllable_hmaster1 & ~n38830;
  assign n38832 = ~n38826 & ~n38831;
  assign n38833 = ~i_hbusreq3 & ~n38832;
  assign n38834 = ~n38824 & ~n38833;
  assign n38835 = controllable_hmaster2 & ~n38834;
  assign n38836 = ~n11066 & ~n38283;
  assign n38837 = ~controllable_hmaster0 & ~n38836;
  assign n38838 = ~n38820 & ~n38837;
  assign n38839 = controllable_hmaster1 & ~n38838;
  assign n38840 = ~n10827 & ~n38322;
  assign n38841 = controllable_hmaster0 & ~n38840;
  assign n38842 = ~controllable_hmaster0 & ~n38818;
  assign n38843 = ~n38841 & ~n38842;
  assign n38844 = ~controllable_hmaster1 & ~n38843;
  assign n38845 = ~n38839 & ~n38844;
  assign n38846 = i_hbusreq3 & ~n38845;
  assign n38847 = ~n11049 & ~n38333;
  assign n38848 = controllable_hmaster0 & ~n38847;
  assign n38849 = ~n11110 & ~n38333;
  assign n38850 = ~controllable_hmaster0 & ~n38849;
  assign n38851 = ~n38848 & ~n38850;
  assign n38852 = controllable_hmaster1 & ~n38851;
  assign n38853 = ~n11049 & ~n38344;
  assign n38854 = controllable_hmaster0 & ~n38853;
  assign n38855 = ~n11127 & ~n38355;
  assign n38856 = ~controllable_hmaster0 & ~n38855;
  assign n38857 = ~n38854 & ~n38856;
  assign n38858 = ~controllable_hmaster1 & ~n38857;
  assign n38859 = ~n38852 & ~n38858;
  assign n38860 = ~i_hbusreq3 & ~n38859;
  assign n38861 = ~n38846 & ~n38860;
  assign n38862 = ~controllable_hmaster2 & ~n38861;
  assign n38863 = ~n38835 & ~n38862;
  assign n38864 = ~controllable_hgrant3 & ~n38863;
  assign n38865 = ~n10110 & ~n38864;
  assign n38866 = controllable_nhgrant0 & ~n38865;
  assign n38867 = ~n10240 & ~n38866;
  assign n38868 = ~n3281 & ~n38867;
  assign n38869 = ~n3281 & ~n38868;
  assign n38870 = ~n3378 & ~n38869;
  assign n38871 = ~n38817 & ~n38870;
  assign n38872 = n3492 & ~n38871;
  assign n38873 = ~n37231 & ~n38872;
  assign n38874 = n3485 & ~n38873;
  assign n38875 = ~n37356 & ~n38874;
  assign n38876 = n3476 & ~n38875;
  assign n38877 = ~n38760 & ~n38876;
  assign n38878 = n3374 & ~n38877;
  assign n38879 = ~n38708 & ~n38878;
  assign n38880 = n3655 & ~n38879;
  assign n38881 = n3378 & ~n36814;
  assign n38882 = ~n4787 & ~n38384;
  assign n38883 = controllable_hmaster1 & ~n38882;
  assign n38884 = controllable_hmaster0 & ~n38882;
  assign n38885 = controllable_hmaster0 & ~n38884;
  assign n38886 = ~controllable_hmaster1 & ~n38885;
  assign n38887 = ~n38883 & ~n38886;
  assign n38888 = i_hbusreq3 & ~n38887;
  assign n38889 = ~n4794 & ~n38396;
  assign n38890 = controllable_hmaster1 & ~n38889;
  assign n38891 = controllable_hmaster0 & ~n38889;
  assign n38892 = controllable_hmaster0 & ~n38891;
  assign n38893 = ~controllable_hmaster1 & ~n38892;
  assign n38894 = ~n38890 & ~n38893;
  assign n38895 = ~i_hbusreq3 & ~n38894;
  assign n38896 = ~n38888 & ~n38895;
  assign n38897 = controllable_hmaster2 & ~n38896;
  assign n38898 = controllable_hmaster2 & ~n38897;
  assign n38899 = ~controllable_hgrant3 & ~n38898;
  assign n38900 = ~n9708 & ~n38899;
  assign n38901 = controllable_nhgrant0 & ~n38900;
  assign n38902 = ~n9753 & ~n38901;
  assign n38903 = ~n3281 & ~n38902;
  assign n38904 = ~n3281 & ~n38903;
  assign n38905 = ~n3378 & ~n38904;
  assign n38906 = ~n38881 & ~n38905;
  assign n38907 = n3492 & ~n38906;
  assign n38908 = n3492 & ~n38907;
  assign n38909 = n3485 & ~n38908;
  assign n38910 = n3485 & ~n38909;
  assign n38911 = ~n3476 & ~n38910;
  assign n38912 = ~n8523 & ~n38907;
  assign n38913 = n3485 & ~n38912;
  assign n38914 = ~n8689 & ~n38913;
  assign n38915 = n3476 & ~n38914;
  assign n38916 = ~n38911 & ~n38915;
  assign n38917 = ~n3374 & ~n38916;
  assign n38918 = n3378 & ~n36885;
  assign n38919 = ~n34874 & ~n38884;
  assign n38920 = ~controllable_hmaster1 & ~n38919;
  assign n38921 = ~n38883 & ~n38920;
  assign n38922 = i_hbusreq3 & ~n38921;
  assign n38923 = ~n34880 & ~n38891;
  assign n38924 = ~controllable_hmaster1 & ~n38923;
  assign n38925 = ~n38890 & ~n38924;
  assign n38926 = ~i_hbusreq3 & ~n38925;
  assign n38927 = ~n38922 & ~n38926;
  assign n38928 = controllable_hmaster2 & ~n38927;
  assign n38929 = ~n4787 & ~n38438;
  assign n38930 = controllable_hmaster0 & ~n38929;
  assign n38931 = ~n10768 & ~n38438;
  assign n38932 = ~controllable_hmaster0 & ~n38931;
  assign n38933 = ~n38930 & ~n38932;
  assign n38934 = controllable_hmaster1 & ~n38933;
  assign n38935 = ~n4787 & ~n38446;
  assign n38936 = controllable_hmaster0 & ~n38935;
  assign n38937 = ~controllable_hmaster0 & ~n38929;
  assign n38938 = ~n38936 & ~n38937;
  assign n38939 = ~controllable_hmaster1 & ~n38938;
  assign n38940 = ~n38934 & ~n38939;
  assign n38941 = i_hbusreq3 & ~n38940;
  assign n38942 = ~n4794 & ~n38458;
  assign n38943 = controllable_hmaster0 & ~n38942;
  assign n38944 = ~n10782 & ~n38458;
  assign n38945 = ~controllable_hmaster0 & ~n38944;
  assign n38946 = ~n38943 & ~n38945;
  assign n38947 = controllable_hmaster1 & ~n38946;
  assign n38948 = ~n4794 & ~n38469;
  assign n38949 = controllable_hmaster0 & ~n38948;
  assign n38950 = ~n38937 & ~n38949;
  assign n38951 = ~controllable_hmaster1 & ~n38950;
  assign n38952 = ~n38947 & ~n38951;
  assign n38953 = ~i_hbusreq3 & ~n38952;
  assign n38954 = ~n38941 & ~n38953;
  assign n38955 = ~controllable_hmaster2 & ~n38954;
  assign n38956 = ~n38928 & ~n38955;
  assign n38957 = ~controllable_hgrant3 & ~n38956;
  assign n38958 = ~n9790 & ~n38957;
  assign n38959 = controllable_nhgrant0 & ~n38958;
  assign n38960 = ~n9861 & ~n38959;
  assign n38961 = ~n3281 & ~n38960;
  assign n38962 = ~n3281 & ~n38961;
  assign n38963 = ~n3378 & ~n38962;
  assign n38964 = ~n38918 & ~n38963;
  assign n38965 = n3492 & ~n38964;
  assign n38966 = n3492 & ~n38965;
  assign n38967 = n3485 & ~n38966;
  assign n38968 = n3485 & ~n38967;
  assign n38969 = ~n3476 & ~n38968;
  assign n38970 = ~n10816 & ~n38493;
  assign n38971 = controllable_hmaster1 & ~n38970;
  assign n38972 = controllable_hmaster0 & ~n38970;
  assign n38973 = ~n10827 & ~n38498;
  assign n38974 = ~controllable_hmaster0 & ~n38973;
  assign n38975 = ~n38972 & ~n38974;
  assign n38976 = ~controllable_hmaster1 & ~n38975;
  assign n38977 = ~n38971 & ~n38976;
  assign n38978 = i_hbusreq3 & ~n38977;
  assign n38979 = ~n10870 & ~n38509;
  assign n38980 = controllable_hmaster1 & ~n38979;
  assign n38981 = controllable_hmaster0 & ~n38979;
  assign n38982 = ~n10904 & ~n38517;
  assign n38983 = ~controllable_hmaster0 & ~n38982;
  assign n38984 = ~n38981 & ~n38983;
  assign n38985 = ~controllable_hmaster1 & ~n38984;
  assign n38986 = ~n38980 & ~n38985;
  assign n38987 = ~i_hbusreq3 & ~n38986;
  assign n38988 = ~n38978 & ~n38987;
  assign n38989 = controllable_hmaster2 & ~n38988;
  assign n38990 = ~n10816 & ~n38527;
  assign n38991 = controllable_hmaster0 & ~n38990;
  assign n38992 = ~n10922 & ~n38527;
  assign n38993 = ~controllable_hmaster0 & ~n38992;
  assign n38994 = ~n38991 & ~n38993;
  assign n38995 = controllable_hmaster1 & ~n38994;
  assign n38996 = ~n10816 & ~n38535;
  assign n38997 = controllable_hmaster0 & ~n38996;
  assign n38998 = ~controllable_hmaster0 & ~n38990;
  assign n38999 = ~n38997 & ~n38998;
  assign n39000 = ~controllable_hmaster1 & ~n38999;
  assign n39001 = ~n38995 & ~n39000;
  assign n39002 = i_hbusreq3 & ~n39001;
  assign n39003 = ~n10870 & ~n38547;
  assign n39004 = controllable_hmaster0 & ~n39003;
  assign n39005 = ~n10972 & ~n38547;
  assign n39006 = ~controllable_hmaster0 & ~n39005;
  assign n39007 = ~n39004 & ~n39006;
  assign n39008 = controllable_hmaster1 & ~n39007;
  assign n39009 = ~n10870 & ~n38558;
  assign n39010 = controllable_hmaster0 & ~n39009;
  assign n39011 = ~n11002 & ~n38564;
  assign n39012 = ~controllable_hmaster0 & ~n39011;
  assign n39013 = ~n39010 & ~n39012;
  assign n39014 = ~controllable_hmaster1 & ~n39013;
  assign n39015 = ~n39008 & ~n39014;
  assign n39016 = ~i_hbusreq3 & ~n39015;
  assign n39017 = ~n39002 & ~n39016;
  assign n39018 = ~controllable_hmaster2 & ~n39017;
  assign n39019 = ~n38989 & ~n39018;
  assign n39020 = ~controllable_hgrant3 & ~n39019;
  assign n39021 = ~n7457 & ~n39020;
  assign n39022 = controllable_nhgrant0 & ~n39021;
  assign n39023 = ~n10071 & ~n39022;
  assign n39024 = ~n3281 & ~n39023;
  assign n39025 = ~n3281 & ~n39024;
  assign n39026 = n3378 & ~n39025;
  assign n39027 = ~n10827 & ~n38582;
  assign n39028 = controllable_hmaster1 & ~n39027;
  assign n39029 = controllable_hmaster0 & ~n39027;
  assign n39030 = ~n38974 & ~n39029;
  assign n39031 = ~controllable_hmaster1 & ~n39030;
  assign n39032 = ~n39028 & ~n39031;
  assign n39033 = i_hbusreq3 & ~n39032;
  assign n39034 = ~n11049 & ~n38594;
  assign n39035 = controllable_hmaster1 & ~n39034;
  assign n39036 = controllable_hmaster0 & ~n39034;
  assign n39037 = ~n11049 & ~n38601;
  assign n39038 = ~controllable_hmaster0 & ~n39037;
  assign n39039 = ~n39036 & ~n39038;
  assign n39040 = ~controllable_hmaster1 & ~n39039;
  assign n39041 = ~n39035 & ~n39040;
  assign n39042 = ~i_hbusreq3 & ~n39041;
  assign n39043 = ~n39033 & ~n39042;
  assign n39044 = controllable_hmaster2 & ~n39043;
  assign n39045 = ~n11066 & ~n38582;
  assign n39046 = ~controllable_hmaster0 & ~n39045;
  assign n39047 = ~n39029 & ~n39046;
  assign n39048 = controllable_hmaster1 & ~n39047;
  assign n39049 = ~n10827 & ~n38615;
  assign n39050 = controllable_hmaster0 & ~n39049;
  assign n39051 = ~controllable_hmaster0 & ~n39027;
  assign n39052 = ~n39050 & ~n39051;
  assign n39053 = ~controllable_hmaster1 & ~n39052;
  assign n39054 = ~n39048 & ~n39053;
  assign n39055 = i_hbusreq3 & ~n39054;
  assign n39056 = ~n11049 & ~n38626;
  assign n39057 = controllable_hmaster0 & ~n39056;
  assign n39058 = ~n11110 & ~n38626;
  assign n39059 = ~controllable_hmaster0 & ~n39058;
  assign n39060 = ~n39057 & ~n39059;
  assign n39061 = controllable_hmaster1 & ~n39060;
  assign n39062 = ~n11049 & ~n38637;
  assign n39063 = controllable_hmaster0 & ~n39062;
  assign n39064 = ~n11127 & ~n38643;
  assign n39065 = ~controllable_hmaster0 & ~n39064;
  assign n39066 = ~n39063 & ~n39065;
  assign n39067 = ~controllable_hmaster1 & ~n39066;
  assign n39068 = ~n39061 & ~n39067;
  assign n39069 = ~i_hbusreq3 & ~n39068;
  assign n39070 = ~n39055 & ~n39069;
  assign n39071 = ~controllable_hmaster2 & ~n39070;
  assign n39072 = ~n39044 & ~n39071;
  assign n39073 = ~controllable_hgrant3 & ~n39072;
  assign n39074 = ~n10110 & ~n39073;
  assign n39075 = controllable_nhgrant0 & ~n39074;
  assign n39076 = ~n10240 & ~n39075;
  assign n39077 = ~n3281 & ~n39076;
  assign n39078 = ~n3281 & ~n39077;
  assign n39079 = ~n3378 & ~n39078;
  assign n39080 = ~n39026 & ~n39079;
  assign n39081 = n3492 & ~n39080;
  assign n39082 = ~n37258 & ~n39081;
  assign n39083 = n3485 & ~n39082;
  assign n39084 = ~n37367 & ~n39083;
  assign n39085 = n3476 & ~n39084;
  assign n39086 = ~n38969 & ~n39085;
  assign n39087 = n3374 & ~n39086;
  assign n39088 = ~n38917 & ~n39087;
  assign n39089 = ~n3655 & ~n39088;
  assign n39090 = ~n38880 & ~n39089;
  assign n39091 = ~n3652 & ~n39090;
  assign n39092 = ~n38671 & ~n39091;
  assign n39093 = n3368 & ~n39092;
  assign n39094 = ~n38081 & ~n39093;
  assign n39095 = ~n3362 & ~n39094;
  assign n39096 = ~n37379 & ~n39095;
  assign n39097 = ~n3359 & ~n39096;
  assign n39098 = ~n37277 & ~n39097;
  assign n39099 = ~n3356 & ~n39098;
  assign n39100 = ~n34938 & ~n39099;
  assign n39101 = n3345 & ~n39100;
  assign n39102 = ~n3649 & ~n39101;
  assign n39103 = ~n3341 & ~n39102;
  assign n39104 = controllable_hmaster0 & ~n37421;
  assign n39105 = controllable_hmaster1 & ~n39104;
  assign n39106 = controllable_hmaster1 & ~n39105;
  assign n39107 = i_hbusreq3 & ~n39106;
  assign n39108 = controllable_hmaster0 & ~n37441;
  assign n39109 = controllable_hmaster1 & ~n39108;
  assign n39110 = controllable_hmaster1 & ~n39109;
  assign n39111 = ~i_hbusreq3 & ~n39110;
  assign n39112 = ~n39107 & ~n39111;
  assign n39113 = ~controllable_hmaster2 & ~n39112;
  assign n39114 = ~controllable_hmaster2 & ~n39113;
  assign n39115 = ~controllable_hgrant3 & ~n39114;
  assign n39116 = ~n11460 & ~n39115;
  assign n39117 = controllable_nhgrant0 & ~n39116;
  assign n39118 = ~n11496 & ~n39117;
  assign n39119 = ~n3281 & ~n39118;
  assign n39120 = ~n3281 & ~n39119;
  assign n39121 = n3378 & ~n39120;
  assign n39122 = ~n3530 & ~n39113;
  assign n39123 = ~controllable_hgrant3 & ~n39122;
  assign n39124 = ~n11502 & ~n39123;
  assign n39125 = controllable_nhgrant0 & ~n39124;
  assign n39126 = ~n11512 & ~n39125;
  assign n39127 = ~n3281 & ~n39126;
  assign n39128 = ~n3950 & ~n39127;
  assign n39129 = ~n3378 & ~n39128;
  assign n39130 = ~n39121 & ~n39129;
  assign n39131 = n3492 & ~n39130;
  assign n39132 = ~n3493 & ~n39131;
  assign n39133 = n3485 & ~n39132;
  assign n39134 = ~n3486 & ~n39133;
  assign n39135 = ~n3476 & ~n39134;
  assign n39136 = ~n11553 & ~n39115;
  assign n39137 = controllable_nhgrant0 & ~n39136;
  assign n39138 = ~n11496 & ~n39137;
  assign n39139 = ~n3281 & ~n39138;
  assign n39140 = ~n3281 & ~n39139;
  assign n39141 = n3378 & ~n39140;
  assign n39142 = ~n3545 & ~n34986;
  assign n39143 = ~controllable_hgrant2 & ~n39142;
  assign n39144 = ~n3410 & ~n39143;
  assign n39145 = controllable_hmaster0 & ~n39144;
  assign n39146 = ~n3556 & ~n39145;
  assign n39147 = controllable_hmaster1 & ~n39146;
  assign n39148 = ~n11581 & ~n39147;
  assign n39149 = i_hbusreq3 & ~n39148;
  assign n39150 = i_hbusreq2 & ~n39142;
  assign n39151 = ~n4134 & ~n35078;
  assign n39152 = ~i_hbusreq2 & ~n39151;
  assign n39153 = ~n39150 & ~n39152;
  assign n39154 = ~controllable_hgrant2 & ~n39153;
  assign n39155 = ~n3859 & ~n39154;
  assign n39156 = controllable_hmaster0 & ~n39155;
  assign n39157 = ~n3596 & ~n39156;
  assign n39158 = controllable_hmaster1 & ~n39157;
  assign n39159 = ~n11592 & ~n39158;
  assign n39160 = ~i_hbusreq3 & ~n39159;
  assign n39161 = ~n39149 & ~n39160;
  assign n39162 = ~controllable_hmaster2 & ~n39161;
  assign n39163 = ~n3602 & ~n39162;
  assign n39164 = ~controllable_hgrant3 & ~n39163;
  assign n39165 = ~n11579 & ~n39164;
  assign n39166 = controllable_nhgrant0 & ~n39165;
  assign n39167 = ~n11512 & ~n39166;
  assign n39168 = ~n3281 & ~n39167;
  assign n39169 = ~n4089 & ~n39168;
  assign n39170 = ~n3378 & ~n39169;
  assign n39171 = ~n39141 & ~n39170;
  assign n39172 = n3492 & ~n39171;
  assign n39173 = ~n3493 & ~n39172;
  assign n39174 = n3485 & ~n39173;
  assign n39175 = ~n3486 & ~n39174;
  assign n39176 = n3476 & ~n39175;
  assign n39177 = ~n39135 & ~n39176;
  assign n39178 = n3374 & ~n39177;
  assign n39179 = ~n11449 & ~n39178;
  assign n39180 = n3655 & ~n39179;
  assign n39181 = controllable_hmaster0 & ~n37615;
  assign n39182 = controllable_hmaster1 & ~n39181;
  assign n39183 = controllable_hmaster1 & ~n39182;
  assign n39184 = i_hbusreq3 & ~n39183;
  assign n39185 = controllable_hmaster0 & ~n37635;
  assign n39186 = controllable_hmaster1 & ~n39185;
  assign n39187 = controllable_hmaster1 & ~n39186;
  assign n39188 = ~i_hbusreq3 & ~n39187;
  assign n39189 = ~n39184 & ~n39188;
  assign n39190 = ~controllable_hmaster2 & ~n39189;
  assign n39191 = ~controllable_hmaster2 & ~n39190;
  assign n39192 = ~controllable_hgrant3 & ~n39191;
  assign n39193 = ~n11460 & ~n39192;
  assign n39194 = controllable_nhgrant0 & ~n39193;
  assign n39195 = ~n11496 & ~n39194;
  assign n39196 = ~n3281 & ~n39195;
  assign n39197 = ~n3281 & ~n39196;
  assign n39198 = n3378 & ~n39197;
  assign n39199 = ~n3530 & ~n39190;
  assign n39200 = ~controllable_hgrant3 & ~n39199;
  assign n39201 = ~n11502 & ~n39200;
  assign n39202 = controllable_nhgrant0 & ~n39201;
  assign n39203 = ~n11512 & ~n39202;
  assign n39204 = ~n3281 & ~n39203;
  assign n39205 = ~n3950 & ~n39204;
  assign n39206 = ~n3378 & ~n39205;
  assign n39207 = ~n39198 & ~n39206;
  assign n39208 = n3492 & ~n39207;
  assign n39209 = ~n3493 & ~n39208;
  assign n39210 = n3485 & ~n39209;
  assign n39211 = ~n3486 & ~n39210;
  assign n39212 = ~n3476 & ~n39211;
  assign n39213 = ~n11553 & ~n39192;
  assign n39214 = controllable_nhgrant0 & ~n39213;
  assign n39215 = ~n11496 & ~n39214;
  assign n39216 = ~n3281 & ~n39215;
  assign n39217 = ~n3281 & ~n39216;
  assign n39218 = n3378 & ~n39217;
  assign n39219 = ~n4279 & ~n34986;
  assign n39220 = ~controllable_hgrant2 & ~n39219;
  assign n39221 = ~n3410 & ~n39220;
  assign n39222 = controllable_hmaster0 & ~n39221;
  assign n39223 = ~n3556 & ~n39222;
  assign n39224 = controllable_hmaster1 & ~n39223;
  assign n39225 = ~n11581 & ~n39224;
  assign n39226 = i_hbusreq3 & ~n39225;
  assign n39227 = i_hbusreq2 & ~n39219;
  assign n39228 = ~n4300 & ~n35078;
  assign n39229 = ~i_hbusreq2 & ~n39228;
  assign n39230 = ~n39227 & ~n39229;
  assign n39231 = ~controllable_hgrant2 & ~n39230;
  assign n39232 = ~n3859 & ~n39231;
  assign n39233 = controllable_hmaster0 & ~n39232;
  assign n39234 = ~n3596 & ~n39233;
  assign n39235 = controllable_hmaster1 & ~n39234;
  assign n39236 = ~n11592 & ~n39235;
  assign n39237 = ~i_hbusreq3 & ~n39236;
  assign n39238 = ~n39226 & ~n39237;
  assign n39239 = ~controllable_hmaster2 & ~n39238;
  assign n39240 = ~n3602 & ~n39239;
  assign n39241 = ~controllable_hgrant3 & ~n39240;
  assign n39242 = ~n11579 & ~n39241;
  assign n39243 = controllable_nhgrant0 & ~n39242;
  assign n39244 = ~n11512 & ~n39243;
  assign n39245 = ~n3281 & ~n39244;
  assign n39246 = ~n4089 & ~n39245;
  assign n39247 = ~n3378 & ~n39246;
  assign n39248 = ~n39218 & ~n39247;
  assign n39249 = n3492 & ~n39248;
  assign n39250 = ~n3493 & ~n39249;
  assign n39251 = n3485 & ~n39250;
  assign n39252 = ~n3486 & ~n39251;
  assign n39253 = n3476 & ~n39252;
  assign n39254 = ~n39212 & ~n39253;
  assign n39255 = n3374 & ~n39254;
  assign n39256 = ~n11449 & ~n39255;
  assign n39257 = ~n3655 & ~n39256;
  assign n39258 = ~n39180 & ~n39257;
  assign n39259 = n3652 & ~n39258;
  assign n39260 = controllable_hmaster0 & ~n37816;
  assign n39261 = controllable_hmaster1 & ~n39260;
  assign n39262 = controllable_hmaster1 & ~n39261;
  assign n39263 = i_hbusreq3 & ~n39262;
  assign n39264 = controllable_hmaster0 & ~n37829;
  assign n39265 = controllable_hmaster1 & ~n39264;
  assign n39266 = controllable_hmaster1 & ~n39265;
  assign n39267 = ~i_hbusreq3 & ~n39266;
  assign n39268 = ~n39263 & ~n39267;
  assign n39269 = ~controllable_hmaster2 & ~n39268;
  assign n39270 = ~controllable_hmaster2 & ~n39269;
  assign n39271 = ~controllable_hgrant3 & ~n39270;
  assign n39272 = ~n11460 & ~n39271;
  assign n39273 = controllable_nhgrant0 & ~n39272;
  assign n39274 = ~n11496 & ~n39273;
  assign n39275 = ~n3281 & ~n39274;
  assign n39276 = ~n3281 & ~n39275;
  assign n39277 = n3378 & ~n39276;
  assign n39278 = ~n3530 & ~n39269;
  assign n39279 = ~controllable_hgrant3 & ~n39278;
  assign n39280 = ~n11502 & ~n39279;
  assign n39281 = controllable_nhgrant0 & ~n39280;
  assign n39282 = ~n11512 & ~n39281;
  assign n39283 = ~n3281 & ~n39282;
  assign n39284 = ~n3950 & ~n39283;
  assign n39285 = ~n3378 & ~n39284;
  assign n39286 = ~n39277 & ~n39285;
  assign n39287 = n3492 & ~n39286;
  assign n39288 = ~n3493 & ~n39287;
  assign n39289 = n3485 & ~n39288;
  assign n39290 = ~n3486 & ~n39289;
  assign n39291 = ~n3476 & ~n39290;
  assign n39292 = ~n11553 & ~n39271;
  assign n39293 = controllable_nhgrant0 & ~n39292;
  assign n39294 = ~n11496 & ~n39293;
  assign n39295 = ~n3281 & ~n39294;
  assign n39296 = ~n3281 & ~n39295;
  assign n39297 = n3378 & ~n39296;
  assign n39298 = ~n4333 & ~n39143;
  assign n39299 = controllable_hmaster0 & ~n39298;
  assign n39300 = ~n3556 & ~n39299;
  assign n39301 = controllable_hmaster1 & ~n39300;
  assign n39302 = ~n11581 & ~n39301;
  assign n39303 = i_hbusreq3 & ~n39302;
  assign n39304 = ~n4340 & ~n39154;
  assign n39305 = controllable_hmaster0 & ~n39304;
  assign n39306 = ~n3596 & ~n39305;
  assign n39307 = controllable_hmaster1 & ~n39306;
  assign n39308 = ~n11592 & ~n39307;
  assign n39309 = ~i_hbusreq3 & ~n39308;
  assign n39310 = ~n39303 & ~n39309;
  assign n39311 = ~controllable_hmaster2 & ~n39310;
  assign n39312 = ~n3602 & ~n39311;
  assign n39313 = ~controllable_hgrant3 & ~n39312;
  assign n39314 = ~n11579 & ~n39313;
  assign n39315 = controllable_nhgrant0 & ~n39314;
  assign n39316 = ~n11512 & ~n39315;
  assign n39317 = ~n3281 & ~n39316;
  assign n39318 = ~n4089 & ~n39317;
  assign n39319 = ~n3378 & ~n39318;
  assign n39320 = ~n39297 & ~n39319;
  assign n39321 = n3492 & ~n39320;
  assign n39322 = ~n3493 & ~n39321;
  assign n39323 = n3485 & ~n39322;
  assign n39324 = ~n3486 & ~n39323;
  assign n39325 = n3476 & ~n39324;
  assign n39326 = ~n39291 & ~n39325;
  assign n39327 = n3374 & ~n39326;
  assign n39328 = ~n11449 & ~n39327;
  assign n39329 = n3655 & ~n39328;
  assign n39330 = controllable_hmaster0 & ~n37970;
  assign n39331 = controllable_hmaster1 & ~n39330;
  assign n39332 = controllable_hmaster1 & ~n39331;
  assign n39333 = i_hbusreq3 & ~n39332;
  assign n39334 = controllable_hmaster0 & ~n37983;
  assign n39335 = controllable_hmaster1 & ~n39334;
  assign n39336 = controllable_hmaster1 & ~n39335;
  assign n39337 = ~i_hbusreq3 & ~n39336;
  assign n39338 = ~n39333 & ~n39337;
  assign n39339 = ~controllable_hmaster2 & ~n39338;
  assign n39340 = ~controllable_hmaster2 & ~n39339;
  assign n39341 = ~controllable_hgrant3 & ~n39340;
  assign n39342 = ~n11460 & ~n39341;
  assign n39343 = controllable_nhgrant0 & ~n39342;
  assign n39344 = ~n11496 & ~n39343;
  assign n39345 = ~n3281 & ~n39344;
  assign n39346 = ~n3281 & ~n39345;
  assign n39347 = n3378 & ~n39346;
  assign n39348 = ~n3530 & ~n39339;
  assign n39349 = ~controllable_hgrant3 & ~n39348;
  assign n39350 = ~n11502 & ~n39349;
  assign n39351 = controllable_nhgrant0 & ~n39350;
  assign n39352 = ~n11512 & ~n39351;
  assign n39353 = ~n3281 & ~n39352;
  assign n39354 = ~n3950 & ~n39353;
  assign n39355 = ~n3378 & ~n39354;
  assign n39356 = ~n39347 & ~n39355;
  assign n39357 = n3492 & ~n39356;
  assign n39358 = ~n3493 & ~n39357;
  assign n39359 = n3485 & ~n39358;
  assign n39360 = ~n3486 & ~n39359;
  assign n39361 = ~n3476 & ~n39360;
  assign n39362 = ~n11553 & ~n39341;
  assign n39363 = controllable_nhgrant0 & ~n39362;
  assign n39364 = ~n11496 & ~n39363;
  assign n39365 = ~n3281 & ~n39364;
  assign n39366 = ~n3281 & ~n39365;
  assign n39367 = n3378 & ~n39366;
  assign n39368 = ~n4333 & ~n39220;
  assign n39369 = controllable_hmaster0 & ~n39368;
  assign n39370 = ~n3556 & ~n39369;
  assign n39371 = controllable_hmaster1 & ~n39370;
  assign n39372 = ~n11581 & ~n39371;
  assign n39373 = i_hbusreq3 & ~n39372;
  assign n39374 = ~n4340 & ~n39231;
  assign n39375 = controllable_hmaster0 & ~n39374;
  assign n39376 = ~n3596 & ~n39375;
  assign n39377 = controllable_hmaster1 & ~n39376;
  assign n39378 = ~n11592 & ~n39377;
  assign n39379 = ~i_hbusreq3 & ~n39378;
  assign n39380 = ~n39373 & ~n39379;
  assign n39381 = ~controllable_hmaster2 & ~n39380;
  assign n39382 = ~n3602 & ~n39381;
  assign n39383 = ~controllable_hgrant3 & ~n39382;
  assign n39384 = ~n11579 & ~n39383;
  assign n39385 = controllable_nhgrant0 & ~n39384;
  assign n39386 = ~n11512 & ~n39385;
  assign n39387 = ~n3281 & ~n39386;
  assign n39388 = ~n4089 & ~n39387;
  assign n39389 = ~n3378 & ~n39388;
  assign n39390 = ~n39367 & ~n39389;
  assign n39391 = n3492 & ~n39390;
  assign n39392 = ~n3493 & ~n39391;
  assign n39393 = n3485 & ~n39392;
  assign n39394 = ~n3486 & ~n39393;
  assign n39395 = n3476 & ~n39394;
  assign n39396 = ~n39361 & ~n39395;
  assign n39397 = n3374 & ~n39396;
  assign n39398 = ~n11449 & ~n39397;
  assign n39399 = ~n3655 & ~n39398;
  assign n39400 = ~n39329 & ~n39399;
  assign n39401 = ~n3652 & ~n39400;
  assign n39402 = ~n39259 & ~n39401;
  assign n39403 = ~n3368 & ~n39402;
  assign n39404 = controllable_hmaster0 & ~n38141;
  assign n39405 = controllable_hmaster1 & ~n39404;
  assign n39406 = controllable_hmaster1 & ~n39405;
  assign n39407 = i_hbusreq3 & ~n39406;
  assign n39408 = controllable_hmaster0 & ~n38161;
  assign n39409 = controllable_hmaster1 & ~n39408;
  assign n39410 = controllable_hmaster1 & ~n39409;
  assign n39411 = ~i_hbusreq3 & ~n39410;
  assign n39412 = ~n39407 & ~n39411;
  assign n39413 = ~controllable_hmaster2 & ~n39412;
  assign n39414 = ~controllable_hmaster2 & ~n39413;
  assign n39415 = ~controllable_hgrant3 & ~n39414;
  assign n39416 = ~n11845 & ~n39415;
  assign n39417 = controllable_nhgrant0 & ~n39416;
  assign n39418 = ~n11874 & ~n39417;
  assign n39419 = ~n3281 & ~n39418;
  assign n39420 = ~n3281 & ~n39419;
  assign n39421 = n3492 & ~n39420;
  assign n39422 = n3492 & ~n39421;
  assign n39423 = n3485 & ~n39422;
  assign n39424 = n3485 & ~n39423;
  assign n39425 = ~n3476 & ~n39424;
  assign n39426 = ~n11891 & ~n39415;
  assign n39427 = controllable_nhgrant0 & ~n39426;
  assign n39428 = ~n11874 & ~n39427;
  assign n39429 = ~n3281 & ~n39428;
  assign n39430 = ~n3281 & ~n39429;
  assign n39431 = n3492 & ~n39430;
  assign n39432 = n3492 & ~n39431;
  assign n39433 = n3485 & ~n39432;
  assign n39434 = n3485 & ~n39433;
  assign n39435 = n3476 & ~n39434;
  assign n39436 = ~n39425 & ~n39435;
  assign n39437 = n3374 & ~n39436;
  assign n39438 = n3374 & ~n39437;
  assign n39439 = n3655 & ~n39438;
  assign n39440 = controllable_hmaster0 & ~n38440;
  assign n39441 = controllable_hmaster1 & ~n39440;
  assign n39442 = controllable_hmaster1 & ~n39441;
  assign n39443 = i_hbusreq3 & ~n39442;
  assign n39444 = controllable_hmaster0 & ~n38460;
  assign n39445 = controllable_hmaster1 & ~n39444;
  assign n39446 = controllable_hmaster1 & ~n39445;
  assign n39447 = ~i_hbusreq3 & ~n39446;
  assign n39448 = ~n39443 & ~n39447;
  assign n39449 = ~controllable_hmaster2 & ~n39448;
  assign n39450 = ~controllable_hmaster2 & ~n39449;
  assign n39451 = ~controllable_hgrant3 & ~n39450;
  assign n39452 = ~n11845 & ~n39451;
  assign n39453 = controllable_nhgrant0 & ~n39452;
  assign n39454 = ~n11874 & ~n39453;
  assign n39455 = ~n3281 & ~n39454;
  assign n39456 = ~n3281 & ~n39455;
  assign n39457 = n3492 & ~n39456;
  assign n39458 = n3492 & ~n39457;
  assign n39459 = n3485 & ~n39458;
  assign n39460 = n3485 & ~n39459;
  assign n39461 = ~n3476 & ~n39460;
  assign n39462 = ~n11891 & ~n39451;
  assign n39463 = controllable_nhgrant0 & ~n39462;
  assign n39464 = ~n11874 & ~n39463;
  assign n39465 = ~n3281 & ~n39464;
  assign n39466 = ~n3281 & ~n39465;
  assign n39467 = n3492 & ~n39466;
  assign n39468 = n3492 & ~n39467;
  assign n39469 = n3485 & ~n39468;
  assign n39470 = n3485 & ~n39469;
  assign n39471 = n3476 & ~n39470;
  assign n39472 = ~n39461 & ~n39471;
  assign n39473 = n3374 & ~n39472;
  assign n39474 = n3374 & ~n39473;
  assign n39475 = ~n3655 & ~n39474;
  assign n39476 = ~n39439 & ~n39475;
  assign n39477 = n3652 & ~n39476;
  assign n39478 = controllable_hmaster0 & ~n38721;
  assign n39479 = controllable_hmaster1 & ~n39478;
  assign n39480 = controllable_hmaster1 & ~n39479;
  assign n39481 = i_hbusreq3 & ~n39480;
  assign n39482 = controllable_hmaster0 & ~n38734;
  assign n39483 = controllable_hmaster1 & ~n39482;
  assign n39484 = controllable_hmaster1 & ~n39483;
  assign n39485 = ~i_hbusreq3 & ~n39484;
  assign n39486 = ~n39481 & ~n39485;
  assign n39487 = ~controllable_hmaster2 & ~n39486;
  assign n39488 = ~controllable_hmaster2 & ~n39487;
  assign n39489 = ~controllable_hgrant3 & ~n39488;
  assign n39490 = ~n11845 & ~n39489;
  assign n39491 = controllable_nhgrant0 & ~n39490;
  assign n39492 = ~n11874 & ~n39491;
  assign n39493 = ~n3281 & ~n39492;
  assign n39494 = ~n3281 & ~n39493;
  assign n39495 = n3492 & ~n39494;
  assign n39496 = n3492 & ~n39495;
  assign n39497 = n3485 & ~n39496;
  assign n39498 = n3485 & ~n39497;
  assign n39499 = ~n3476 & ~n39498;
  assign n39500 = ~n11891 & ~n39489;
  assign n39501 = controllable_nhgrant0 & ~n39500;
  assign n39502 = ~n11874 & ~n39501;
  assign n39503 = ~n3281 & ~n39502;
  assign n39504 = ~n3281 & ~n39503;
  assign n39505 = n3492 & ~n39504;
  assign n39506 = n3492 & ~n39505;
  assign n39507 = n3485 & ~n39506;
  assign n39508 = n3485 & ~n39507;
  assign n39509 = n3476 & ~n39508;
  assign n39510 = ~n39499 & ~n39509;
  assign n39511 = n3374 & ~n39510;
  assign n39512 = n3374 & ~n39511;
  assign n39513 = n3655 & ~n39512;
  assign n39514 = controllable_hmaster0 & ~n38930;
  assign n39515 = controllable_hmaster1 & ~n39514;
  assign n39516 = controllable_hmaster1 & ~n39515;
  assign n39517 = i_hbusreq3 & ~n39516;
  assign n39518 = controllable_hmaster0 & ~n38943;
  assign n39519 = controllable_hmaster1 & ~n39518;
  assign n39520 = controllable_hmaster1 & ~n39519;
  assign n39521 = ~i_hbusreq3 & ~n39520;
  assign n39522 = ~n39517 & ~n39521;
  assign n39523 = ~controllable_hmaster2 & ~n39522;
  assign n39524 = ~controllable_hmaster2 & ~n39523;
  assign n39525 = ~controllable_hgrant3 & ~n39524;
  assign n39526 = ~n11845 & ~n39525;
  assign n39527 = controllable_nhgrant0 & ~n39526;
  assign n39528 = ~n11874 & ~n39527;
  assign n39529 = ~n3281 & ~n39528;
  assign n39530 = ~n3281 & ~n39529;
  assign n39531 = n3492 & ~n39530;
  assign n39532 = n3492 & ~n39531;
  assign n39533 = n3485 & ~n39532;
  assign n39534 = n3485 & ~n39533;
  assign n39535 = ~n3476 & ~n39534;
  assign n39536 = ~n11891 & ~n39525;
  assign n39537 = controllable_nhgrant0 & ~n39536;
  assign n39538 = ~n11874 & ~n39537;
  assign n39539 = ~n3281 & ~n39538;
  assign n39540 = ~n3281 & ~n39539;
  assign n39541 = n3492 & ~n39540;
  assign n39542 = n3492 & ~n39541;
  assign n39543 = n3485 & ~n39542;
  assign n39544 = n3485 & ~n39543;
  assign n39545 = n3476 & ~n39544;
  assign n39546 = ~n39535 & ~n39545;
  assign n39547 = n3374 & ~n39546;
  assign n39548 = n3374 & ~n39547;
  assign n39549 = ~n3655 & ~n39548;
  assign n39550 = ~n39513 & ~n39549;
  assign n39551 = ~n3652 & ~n39550;
  assign n39552 = ~n39477 & ~n39551;
  assign n39553 = n3368 & ~n39552;
  assign n39554 = ~n39403 & ~n39553;
  assign n39555 = ~n3362 & ~n39554;
  assign n39556 = ~n3362 & ~n39555;
  assign n39557 = ~n3359 & ~n39556;
  assign n39558 = ~n3359 & ~n39557;
  assign n39559 = n3356 & ~n39558;
  assign n39560 = ~n5041 & ~n34986;
  assign n39561 = ~controllable_hgrant2 & ~n39560;
  assign n39562 = ~n3410 & ~n39561;
  assign n39563 = controllable_hmaster1 & ~n39562;
  assign n39564 = controllable_hmaster0 & ~n39562;
  assign n39565 = ~n34022 & ~n39564;
  assign n39566 = ~controllable_hmaster1 & ~n39565;
  assign n39567 = ~n39563 & ~n39566;
  assign n39568 = i_hbusreq3 & ~n39567;
  assign n39569 = i_hbusreq2 & ~n39560;
  assign n39570 = ~n5064 & ~n35078;
  assign n39571 = ~i_hbusreq2 & ~n39570;
  assign n39572 = ~n39569 & ~n39571;
  assign n39573 = ~controllable_hgrant2 & ~n39572;
  assign n39574 = ~n3859 & ~n39573;
  assign n39575 = controllable_hmaster1 & ~n39574;
  assign n39576 = controllable_hmaster0 & ~n39574;
  assign n39577 = ~n34040 & ~n39576;
  assign n39578 = ~controllable_hmaster1 & ~n39577;
  assign n39579 = ~n39575 & ~n39578;
  assign n39580 = ~i_hbusreq3 & ~n39579;
  assign n39581 = ~n39568 & ~n39580;
  assign n39582 = controllable_hmaster2 & ~n39581;
  assign n39583 = ~n5161 & ~n39582;
  assign n39584 = ~controllable_hgrant3 & ~n39583;
  assign n39585 = ~n5037 & ~n39584;
  assign n39586 = controllable_nhgrant0 & ~n39585;
  assign n39587 = ~n5245 & ~n39586;
  assign n39588 = ~n3281 & ~n39587;
  assign n39589 = ~n3783 & ~n39588;
  assign n39590 = ~n3378 & ~n39589;
  assign n39591 = ~n12026 & ~n39590;
  assign n39592 = n3492 & ~n39591;
  assign n39593 = ~n3631 & ~n39592;
  assign n39594 = n3485 & ~n39593;
  assign n39595 = ~n3630 & ~n39594;
  assign n39596 = ~n3374 & ~n39595;
  assign n39597 = ~n5291 & ~n37421;
  assign n39598 = controllable_hmaster1 & ~n39597;
  assign n39599 = ~n5305 & ~n39598;
  assign n39600 = i_hbusreq3 & ~n39599;
  assign n39601 = ~n5311 & ~n37441;
  assign n39602 = controllable_hmaster1 & ~n39601;
  assign n39603 = ~n5334 & ~n39602;
  assign n39604 = ~i_hbusreq3 & ~n39603;
  assign n39605 = ~n39600 & ~n39604;
  assign n39606 = ~controllable_hmaster2 & ~n39605;
  assign n39607 = ~n12065 & ~n39606;
  assign n39608 = ~controllable_hgrant3 & ~n39607;
  assign n39609 = ~n12041 & ~n39608;
  assign n39610 = controllable_nhgrant0 & ~n39609;
  assign n39611 = ~n12101 & ~n39610;
  assign n39612 = ~n3281 & ~n39611;
  assign n39613 = ~n3950 & ~n39612;
  assign n39614 = n3378 & ~n39613;
  assign n39615 = ~n3497 & ~n34986;
  assign n39616 = ~controllable_hgrant2 & ~n39615;
  assign n39617 = ~n3410 & ~n39616;
  assign n39618 = controllable_hmaster1 & ~n39617;
  assign n39619 = controllable_hmaster0 & ~n39617;
  assign n39620 = ~n3906 & ~n34121;
  assign n39621 = ~controllable_hgrant2 & ~n39620;
  assign n39622 = ~n3410 & ~n39621;
  assign n39623 = ~controllable_hmaster0 & ~n39622;
  assign n39624 = ~n39619 & ~n39623;
  assign n39625 = ~controllable_hmaster1 & ~n39624;
  assign n39626 = ~n39618 & ~n39625;
  assign n39627 = i_hbusreq3 & ~n39626;
  assign n39628 = i_hbusreq2 & ~n39615;
  assign n39629 = ~n5410 & ~n35078;
  assign n39630 = ~i_hbusreq2 & ~n39629;
  assign n39631 = ~n39628 & ~n39630;
  assign n39632 = ~controllable_hgrant2 & ~n39631;
  assign n39633 = ~n3859 & ~n39632;
  assign n39634 = controllable_hmaster1 & ~n39633;
  assign n39635 = controllable_hmaster0 & ~n39633;
  assign n39636 = i_hbusreq2 & ~n39620;
  assign n39637 = ~n3929 & ~n34131;
  assign n39638 = ~i_hbusreq2 & ~n39637;
  assign n39639 = ~n39636 & ~n39638;
  assign n39640 = ~controllable_hgrant2 & ~n39639;
  assign n39641 = ~n3859 & ~n39640;
  assign n39642 = ~controllable_hmaster0 & ~n39641;
  assign n39643 = ~n39635 & ~n39642;
  assign n39644 = ~controllable_hmaster1 & ~n39643;
  assign n39645 = ~n39634 & ~n39644;
  assign n39646 = ~i_hbusreq3 & ~n39645;
  assign n39647 = ~n39627 & ~n39646;
  assign n39648 = controllable_hmaster2 & ~n39647;
  assign n39649 = ~n35055 & ~n37421;
  assign n39650 = controllable_hmaster1 & ~n39649;
  assign n39651 = ~n35064 & ~n39650;
  assign n39652 = i_hbusreq3 & ~n39651;
  assign n39653 = ~n35074 & ~n37441;
  assign n39654 = controllable_hmaster1 & ~n39653;
  assign n39655 = ~n35091 & ~n39654;
  assign n39656 = ~i_hbusreq3 & ~n39655;
  assign n39657 = ~n39652 & ~n39656;
  assign n39658 = ~controllable_hmaster2 & ~n39657;
  assign n39659 = ~n39648 & ~n39658;
  assign n39660 = ~controllable_hgrant3 & ~n39659;
  assign n39661 = ~n5402 & ~n39660;
  assign n39662 = controllable_nhgrant0 & ~n39661;
  assign n39663 = ~n5534 & ~n39662;
  assign n39664 = ~n3281 & ~n39663;
  assign n39665 = ~n3950 & ~n39664;
  assign n39666 = ~n3378 & ~n39665;
  assign n39667 = ~n39614 & ~n39666;
  assign n39668 = n3492 & ~n39667;
  assign n39669 = ~n3631 & ~n39668;
  assign n39670 = n3485 & ~n39669;
  assign n39671 = ~n3630 & ~n39670;
  assign n39672 = ~n3476 & ~n39671;
  assign n39673 = controllable_hgrant4 & ~n5759;
  assign n39674 = ~n5621 & ~n39673;
  assign n39675 = ~controllable_hgrant2 & ~n39674;
  assign n39676 = ~n5616 & ~n39675;
  assign n39677 = controllable_hmaster0 & ~n39676;
  assign n39678 = ~n5688 & ~n39677;
  assign n39679 = controllable_hmaster1 & ~n39678;
  assign n39680 = ~n5704 & ~n39679;
  assign n39681 = i_hbusreq3 & ~n39680;
  assign n39682 = i_hbusreq2 & ~n39674;
  assign n39683 = controllable_hgrant4 & ~n5780;
  assign n39684 = ~n5667 & ~n39683;
  assign n39685 = ~i_hbusreq2 & ~n39684;
  assign n39686 = ~n39682 & ~n39685;
  assign n39687 = ~controllable_hgrant2 & ~n39686;
  assign n39688 = ~n5657 & ~n39687;
  assign n39689 = controllable_hmaster0 & ~n39688;
  assign n39690 = ~n12210 & ~n39689;
  assign n39691 = controllable_hmaster1 & ~n39690;
  assign n39692 = ~n12222 & ~n39691;
  assign n39693 = ~i_hbusreq3 & ~n39692;
  assign n39694 = ~n39681 & ~n39693;
  assign n39695 = ~controllable_hmaster2 & ~n39694;
  assign n39696 = ~n12193 & ~n39695;
  assign n39697 = ~controllable_hgrant3 & ~n39696;
  assign n39698 = ~n12163 & ~n39697;
  assign n39699 = controllable_nhgrant0 & ~n39698;
  assign n39700 = ~n12249 & ~n39699;
  assign n39701 = ~n3281 & ~n39700;
  assign n39702 = ~n4089 & ~n39701;
  assign n39703 = n3378 & ~n39702;
  assign n39704 = controllable_hmaster1 & ~n37502;
  assign n39705 = ~n5911 & ~n34195;
  assign n39706 = ~controllable_hgrant2 & ~n39705;
  assign n39707 = ~n5616 & ~n39706;
  assign n39708 = ~controllable_hmaster0 & ~n39707;
  assign n39709 = ~n37503 & ~n39708;
  assign n39710 = ~controllable_hmaster1 & ~n39709;
  assign n39711 = ~n39704 & ~n39710;
  assign n39712 = i_hbusreq3 & ~n39711;
  assign n39713 = ~n5877 & ~n35234;
  assign n39714 = ~i_hbusreq2 & ~n39713;
  assign n39715 = ~n37517 & ~n39714;
  assign n39716 = ~controllable_hgrant2 & ~n39715;
  assign n39717 = ~n5862 & ~n39716;
  assign n39718 = controllable_hmaster1 & ~n39717;
  assign n39719 = controllable_hmaster0 & ~n39717;
  assign n39720 = i_hbusreq2 & ~n39705;
  assign n39721 = ~n5943 & ~n34214;
  assign n39722 = ~i_hbusreq2 & ~n39721;
  assign n39723 = ~n39720 & ~n39722;
  assign n39724 = ~controllable_hgrant2 & ~n39723;
  assign n39725 = ~n5862 & ~n39724;
  assign n39726 = ~controllable_hmaster0 & ~n39725;
  assign n39727 = ~n39719 & ~n39726;
  assign n39728 = ~controllable_hmaster1 & ~n39727;
  assign n39729 = ~n39718 & ~n39728;
  assign n39730 = ~i_hbusreq3 & ~n39729;
  assign n39731 = ~n39712 & ~n39730;
  assign n39732 = controllable_hmaster2 & ~n39731;
  assign n39733 = ~n35221 & ~n37503;
  assign n39734 = controllable_hmaster1 & ~n39733;
  assign n39735 = ~n35230 & ~n39734;
  assign n39736 = i_hbusreq3 & ~n39735;
  assign n39737 = ~n5897 & ~n35234;
  assign n39738 = ~i_hbusreq2 & ~n39737;
  assign n39739 = ~n37517 & ~n39738;
  assign n39740 = ~controllable_hgrant2 & ~n39739;
  assign n39741 = ~n5862 & ~n39740;
  assign n39742 = controllable_hmaster0 & ~n39741;
  assign n39743 = ~n35242 & ~n39742;
  assign n39744 = controllable_hmaster1 & ~n39743;
  assign n39745 = ~n35260 & ~n39744;
  assign n39746 = ~i_hbusreq3 & ~n39745;
  assign n39747 = ~n39736 & ~n39746;
  assign n39748 = ~controllable_hmaster2 & ~n39747;
  assign n39749 = ~n39732 & ~n39748;
  assign n39750 = ~controllable_hgrant3 & ~n39749;
  assign n39751 = ~n5861 & ~n39750;
  assign n39752 = controllable_nhgrant0 & ~n39751;
  assign n39753 = ~n6082 & ~n39752;
  assign n39754 = ~n3281 & ~n39753;
  assign n39755 = ~n4089 & ~n39754;
  assign n39756 = ~n3378 & ~n39755;
  assign n39757 = ~n39703 & ~n39756;
  assign n39758 = n3492 & ~n39757;
  assign n39759 = ~n3631 & ~n39758;
  assign n39760 = n3485 & ~n39759;
  assign n39761 = ~n3630 & ~n39760;
  assign n39762 = n3476 & ~n39761;
  assign n39763 = ~n39672 & ~n39762;
  assign n39764 = n3374 & ~n39763;
  assign n39765 = ~n39596 & ~n39764;
  assign n39766 = n3655 & ~n39765;
  assign n39767 = ~n6100 & ~n34986;
  assign n39768 = ~controllable_hgrant2 & ~n39767;
  assign n39769 = ~n3410 & ~n39768;
  assign n39770 = controllable_hmaster1 & ~n39769;
  assign n39771 = controllable_hmaster0 & ~n39769;
  assign n39772 = ~n34022 & ~n39771;
  assign n39773 = ~controllable_hmaster1 & ~n39772;
  assign n39774 = ~n39770 & ~n39773;
  assign n39775 = i_hbusreq3 & ~n39774;
  assign n39776 = i_hbusreq2 & ~n39767;
  assign n39777 = ~n6123 & ~n35078;
  assign n39778 = ~i_hbusreq2 & ~n39777;
  assign n39779 = ~n39776 & ~n39778;
  assign n39780 = ~controllable_hgrant2 & ~n39779;
  assign n39781 = ~n3859 & ~n39780;
  assign n39782 = controllable_hmaster1 & ~n39781;
  assign n39783 = controllable_hmaster0 & ~n39781;
  assign n39784 = ~n34040 & ~n39783;
  assign n39785 = ~controllable_hmaster1 & ~n39784;
  assign n39786 = ~n39782 & ~n39785;
  assign n39787 = ~i_hbusreq3 & ~n39786;
  assign n39788 = ~n39775 & ~n39787;
  assign n39789 = controllable_hmaster2 & ~n39788;
  assign n39790 = ~n6188 & ~n39789;
  assign n39791 = ~controllable_hgrant3 & ~n39790;
  assign n39792 = ~n5037 & ~n39791;
  assign n39793 = controllable_nhgrant0 & ~n39792;
  assign n39794 = ~n5245 & ~n39793;
  assign n39795 = ~n3281 & ~n39794;
  assign n39796 = ~n3783 & ~n39795;
  assign n39797 = ~n3378 & ~n39796;
  assign n39798 = ~n12026 & ~n39797;
  assign n39799 = n3492 & ~n39798;
  assign n39800 = ~n3631 & ~n39799;
  assign n39801 = n3485 & ~n39800;
  assign n39802 = ~n3630 & ~n39801;
  assign n39803 = ~n3374 & ~n39802;
  assign n39804 = ~n5291 & ~n37615;
  assign n39805 = controllable_hmaster1 & ~n39804;
  assign n39806 = ~n5305 & ~n39805;
  assign n39807 = i_hbusreq3 & ~n39806;
  assign n39808 = ~n5311 & ~n37635;
  assign n39809 = controllable_hmaster1 & ~n39808;
  assign n39810 = ~n5334 & ~n39809;
  assign n39811 = ~i_hbusreq3 & ~n39810;
  assign n39812 = ~n39807 & ~n39811;
  assign n39813 = ~controllable_hmaster2 & ~n39812;
  assign n39814 = ~n12065 & ~n39813;
  assign n39815 = ~controllable_hgrant3 & ~n39814;
  assign n39816 = ~n12041 & ~n39815;
  assign n39817 = controllable_nhgrant0 & ~n39816;
  assign n39818 = ~n12101 & ~n39817;
  assign n39819 = ~n3281 & ~n39818;
  assign n39820 = ~n3950 & ~n39819;
  assign n39821 = n3378 & ~n39820;
  assign n39822 = ~n6212 & ~n34986;
  assign n39823 = ~controllable_hgrant2 & ~n39822;
  assign n39824 = ~n3410 & ~n39823;
  assign n39825 = controllable_hmaster1 & ~n39824;
  assign n39826 = controllable_hmaster0 & ~n39824;
  assign n39827 = ~n6250 & ~n34121;
  assign n39828 = ~controllable_hgrant2 & ~n39827;
  assign n39829 = ~n3410 & ~n39828;
  assign n39830 = ~controllable_hmaster0 & ~n39829;
  assign n39831 = ~n39826 & ~n39830;
  assign n39832 = ~controllable_hmaster1 & ~n39831;
  assign n39833 = ~n39825 & ~n39832;
  assign n39834 = i_hbusreq3 & ~n39833;
  assign n39835 = i_hbusreq2 & ~n39822;
  assign n39836 = ~n6233 & ~n35078;
  assign n39837 = ~i_hbusreq2 & ~n39836;
  assign n39838 = ~n39835 & ~n39837;
  assign n39839 = ~controllable_hgrant2 & ~n39838;
  assign n39840 = ~n3859 & ~n39839;
  assign n39841 = controllable_hmaster1 & ~n39840;
  assign n39842 = controllable_hmaster0 & ~n39840;
  assign n39843 = i_hbusreq2 & ~n39827;
  assign n39844 = ~n6287 & ~n34131;
  assign n39845 = ~i_hbusreq2 & ~n39844;
  assign n39846 = ~n39843 & ~n39845;
  assign n39847 = ~controllable_hgrant2 & ~n39846;
  assign n39848 = ~n3859 & ~n39847;
  assign n39849 = ~controllable_hmaster0 & ~n39848;
  assign n39850 = ~n39842 & ~n39849;
  assign n39851 = ~controllable_hmaster1 & ~n39850;
  assign n39852 = ~n39841 & ~n39851;
  assign n39853 = ~i_hbusreq3 & ~n39852;
  assign n39854 = ~n39834 & ~n39853;
  assign n39855 = controllable_hmaster2 & ~n39854;
  assign n39856 = ~n35362 & ~n37615;
  assign n39857 = controllable_hmaster1 & ~n39856;
  assign n39858 = ~n35371 & ~n39857;
  assign n39859 = i_hbusreq3 & ~n39858;
  assign n39860 = ~n35382 & ~n37635;
  assign n39861 = controllable_hmaster1 & ~n39860;
  assign n39862 = ~n35400 & ~n39861;
  assign n39863 = ~i_hbusreq3 & ~n39862;
  assign n39864 = ~n39859 & ~n39863;
  assign n39865 = ~controllable_hmaster2 & ~n39864;
  assign n39866 = ~n39855 & ~n39865;
  assign n39867 = ~controllable_hgrant3 & ~n39866;
  assign n39868 = ~n5402 & ~n39867;
  assign n39869 = controllable_nhgrant0 & ~n39868;
  assign n39870 = ~n5534 & ~n39869;
  assign n39871 = ~n3281 & ~n39870;
  assign n39872 = ~n3950 & ~n39871;
  assign n39873 = ~n3378 & ~n39872;
  assign n39874 = ~n39821 & ~n39873;
  assign n39875 = n3492 & ~n39874;
  assign n39876 = ~n3631 & ~n39875;
  assign n39877 = n3485 & ~n39876;
  assign n39878 = ~n3630 & ~n39877;
  assign n39879 = ~n3476 & ~n39878;
  assign n39880 = ~n6359 & ~n39673;
  assign n39881 = ~controllable_hgrant2 & ~n39880;
  assign n39882 = ~n5616 & ~n39881;
  assign n39883 = controllable_hmaster0 & ~n39882;
  assign n39884 = ~n5688 & ~n39883;
  assign n39885 = controllable_hmaster1 & ~n39884;
  assign n39886 = ~n5704 & ~n39885;
  assign n39887 = i_hbusreq3 & ~n39886;
  assign n39888 = i_hbusreq2 & ~n39880;
  assign n39889 = ~n6380 & ~n39683;
  assign n39890 = ~i_hbusreq2 & ~n39889;
  assign n39891 = ~n39888 & ~n39890;
  assign n39892 = ~controllable_hgrant2 & ~n39891;
  assign n39893 = ~n5657 & ~n39892;
  assign n39894 = controllable_hmaster0 & ~n39893;
  assign n39895 = ~n12210 & ~n39894;
  assign n39896 = controllable_hmaster1 & ~n39895;
  assign n39897 = ~n12222 & ~n39896;
  assign n39898 = ~i_hbusreq3 & ~n39897;
  assign n39899 = ~n39887 & ~n39898;
  assign n39900 = ~controllable_hmaster2 & ~n39899;
  assign n39901 = ~n12193 & ~n39900;
  assign n39902 = ~controllable_hgrant3 & ~n39901;
  assign n39903 = ~n12163 & ~n39902;
  assign n39904 = controllable_nhgrant0 & ~n39903;
  assign n39905 = ~n12249 & ~n39904;
  assign n39906 = ~n3281 & ~n39905;
  assign n39907 = ~n4089 & ~n39906;
  assign n39908 = n3378 & ~n39907;
  assign n39909 = controllable_hmaster1 & ~n37705;
  assign n39910 = ~n6465 & ~n34195;
  assign n39911 = ~controllable_hgrant2 & ~n39910;
  assign n39912 = ~n5616 & ~n39911;
  assign n39913 = ~controllable_hmaster0 & ~n39912;
  assign n39914 = ~n37706 & ~n39913;
  assign n39915 = ~controllable_hmaster1 & ~n39914;
  assign n39916 = ~n39909 & ~n39915;
  assign n39917 = i_hbusreq3 & ~n39916;
  assign n39918 = ~n6433 & ~n35234;
  assign n39919 = ~i_hbusreq2 & ~n39918;
  assign n39920 = ~n37720 & ~n39919;
  assign n39921 = ~controllable_hgrant2 & ~n39920;
  assign n39922 = ~n5862 & ~n39921;
  assign n39923 = controllable_hmaster1 & ~n39922;
  assign n39924 = controllable_hmaster0 & ~n39922;
  assign n39925 = i_hbusreq2 & ~n39910;
  assign n39926 = ~n6498 & ~n34214;
  assign n39927 = ~i_hbusreq2 & ~n39926;
  assign n39928 = ~n39925 & ~n39927;
  assign n39929 = ~controllable_hgrant2 & ~n39928;
  assign n39930 = ~n5862 & ~n39929;
  assign n39931 = ~controllable_hmaster0 & ~n39930;
  assign n39932 = ~n39924 & ~n39931;
  assign n39933 = ~controllable_hmaster1 & ~n39932;
  assign n39934 = ~n39923 & ~n39933;
  assign n39935 = ~i_hbusreq3 & ~n39934;
  assign n39936 = ~n39917 & ~n39935;
  assign n39937 = controllable_hmaster2 & ~n39936;
  assign n39938 = ~n35487 & ~n37706;
  assign n39939 = controllable_hmaster1 & ~n39938;
  assign n39940 = ~n35496 & ~n39939;
  assign n39941 = i_hbusreq3 & ~n39940;
  assign n39942 = ~n6451 & ~n35234;
  assign n39943 = ~i_hbusreq2 & ~n39942;
  assign n39944 = ~n37720 & ~n39943;
  assign n39945 = ~controllable_hgrant2 & ~n39944;
  assign n39946 = ~n5862 & ~n39945;
  assign n39947 = controllable_hmaster0 & ~n39946;
  assign n39948 = ~n35507 & ~n39947;
  assign n39949 = controllable_hmaster1 & ~n39948;
  assign n39950 = ~n35524 & ~n39949;
  assign n39951 = ~i_hbusreq3 & ~n39950;
  assign n39952 = ~n39941 & ~n39951;
  assign n39953 = ~controllable_hmaster2 & ~n39952;
  assign n39954 = ~n39937 & ~n39953;
  assign n39955 = ~controllable_hgrant3 & ~n39954;
  assign n39956 = ~n5861 & ~n39955;
  assign n39957 = controllable_nhgrant0 & ~n39956;
  assign n39958 = ~n6082 & ~n39957;
  assign n39959 = ~n3281 & ~n39958;
  assign n39960 = ~n4089 & ~n39959;
  assign n39961 = ~n3378 & ~n39960;
  assign n39962 = ~n39908 & ~n39961;
  assign n39963 = n3492 & ~n39962;
  assign n39964 = ~n3631 & ~n39963;
  assign n39965 = n3485 & ~n39964;
  assign n39966 = ~n3630 & ~n39965;
  assign n39967 = n3476 & ~n39966;
  assign n39968 = ~n39879 & ~n39967;
  assign n39969 = n3374 & ~n39968;
  assign n39970 = ~n39803 & ~n39969;
  assign n39971 = ~n3655 & ~n39970;
  assign n39972 = ~n39766 & ~n39971;
  assign n39973 = n3652 & ~n39972;
  assign n39974 = ~n4333 & ~n39561;
  assign n39975 = controllable_hmaster1 & ~n39974;
  assign n39976 = controllable_hmaster0 & ~n39974;
  assign n39977 = ~n34022 & ~n39976;
  assign n39978 = ~controllable_hmaster1 & ~n39977;
  assign n39979 = ~n39975 & ~n39978;
  assign n39980 = i_hbusreq3 & ~n39979;
  assign n39981 = ~n4340 & ~n39573;
  assign n39982 = controllable_hmaster1 & ~n39981;
  assign n39983 = controllable_hmaster0 & ~n39981;
  assign n39984 = ~n34040 & ~n39983;
  assign n39985 = ~controllable_hmaster1 & ~n39984;
  assign n39986 = ~n39982 & ~n39985;
  assign n39987 = ~i_hbusreq3 & ~n39986;
  assign n39988 = ~n39980 & ~n39987;
  assign n39989 = controllable_hmaster2 & ~n39988;
  assign n39990 = ~n6657 & ~n39989;
  assign n39991 = ~controllable_hgrant3 & ~n39990;
  assign n39992 = ~n5037 & ~n39991;
  assign n39993 = controllable_nhgrant0 & ~n39992;
  assign n39994 = ~n5245 & ~n39993;
  assign n39995 = ~n3281 & ~n39994;
  assign n39996 = ~n3783 & ~n39995;
  assign n39997 = ~n3378 & ~n39996;
  assign n39998 = ~n12026 & ~n39997;
  assign n39999 = n3492 & ~n39998;
  assign n40000 = ~n3631 & ~n39999;
  assign n40001 = n3485 & ~n40000;
  assign n40002 = ~n3630 & ~n40001;
  assign n40003 = ~n3374 & ~n40002;
  assign n40004 = ~n5291 & ~n37816;
  assign n40005 = controllable_hmaster1 & ~n40004;
  assign n40006 = ~n5305 & ~n40005;
  assign n40007 = i_hbusreq3 & ~n40006;
  assign n40008 = ~n5311 & ~n37829;
  assign n40009 = controllable_hmaster1 & ~n40008;
  assign n40010 = ~n5334 & ~n40009;
  assign n40011 = ~i_hbusreq3 & ~n40010;
  assign n40012 = ~n40007 & ~n40011;
  assign n40013 = ~controllable_hmaster2 & ~n40012;
  assign n40014 = ~n12065 & ~n40013;
  assign n40015 = ~controllable_hgrant3 & ~n40014;
  assign n40016 = ~n12041 & ~n40015;
  assign n40017 = controllable_nhgrant0 & ~n40016;
  assign n40018 = ~n12101 & ~n40017;
  assign n40019 = ~n3281 & ~n40018;
  assign n40020 = ~n3950 & ~n40019;
  assign n40021 = n3378 & ~n40020;
  assign n40022 = ~n4333 & ~n39616;
  assign n40023 = controllable_hmaster1 & ~n40022;
  assign n40024 = controllable_hmaster0 & ~n40022;
  assign n40025 = ~n4333 & ~n39621;
  assign n40026 = ~controllable_hmaster0 & ~n40025;
  assign n40027 = ~n40024 & ~n40026;
  assign n40028 = ~controllable_hmaster1 & ~n40027;
  assign n40029 = ~n40023 & ~n40028;
  assign n40030 = i_hbusreq3 & ~n40029;
  assign n40031 = ~n4340 & ~n39632;
  assign n40032 = controllable_hmaster1 & ~n40031;
  assign n40033 = controllable_hmaster0 & ~n40031;
  assign n40034 = ~n4340 & ~n39640;
  assign n40035 = ~controllable_hmaster0 & ~n40034;
  assign n40036 = ~n40033 & ~n40035;
  assign n40037 = ~controllable_hmaster1 & ~n40036;
  assign n40038 = ~n40032 & ~n40037;
  assign n40039 = ~i_hbusreq3 & ~n40038;
  assign n40040 = ~n40030 & ~n40039;
  assign n40041 = controllable_hmaster2 & ~n40040;
  assign n40042 = ~n35612 & ~n37816;
  assign n40043 = controllable_hmaster1 & ~n40042;
  assign n40044 = ~n35619 & ~n40043;
  assign n40045 = i_hbusreq3 & ~n40044;
  assign n40046 = ~n35625 & ~n37829;
  assign n40047 = controllable_hmaster1 & ~n40046;
  assign n40048 = ~n35633 & ~n40047;
  assign n40049 = ~i_hbusreq3 & ~n40048;
  assign n40050 = ~n40045 & ~n40049;
  assign n40051 = ~controllable_hmaster2 & ~n40050;
  assign n40052 = ~n40041 & ~n40051;
  assign n40053 = ~controllable_hgrant3 & ~n40052;
  assign n40054 = ~n5402 & ~n40053;
  assign n40055 = controllable_nhgrant0 & ~n40054;
  assign n40056 = ~n5534 & ~n40055;
  assign n40057 = ~n3281 & ~n40056;
  assign n40058 = ~n3950 & ~n40057;
  assign n40059 = ~n3378 & ~n40058;
  assign n40060 = ~n40021 & ~n40059;
  assign n40061 = n3492 & ~n40060;
  assign n40062 = ~n3631 & ~n40061;
  assign n40063 = n3485 & ~n40062;
  assign n40064 = ~n3630 & ~n40063;
  assign n40065 = ~n3476 & ~n40064;
  assign n40066 = ~n6738 & ~n39675;
  assign n40067 = controllable_hmaster0 & ~n40066;
  assign n40068 = ~n5688 & ~n40067;
  assign n40069 = controllable_hmaster1 & ~n40068;
  assign n40070 = ~n5704 & ~n40069;
  assign n40071 = i_hbusreq3 & ~n40070;
  assign n40072 = ~n6745 & ~n39687;
  assign n40073 = controllable_hmaster0 & ~n40072;
  assign n40074 = ~n12210 & ~n40073;
  assign n40075 = controllable_hmaster1 & ~n40074;
  assign n40076 = ~n12222 & ~n40075;
  assign n40077 = ~i_hbusreq3 & ~n40076;
  assign n40078 = ~n40071 & ~n40077;
  assign n40079 = ~controllable_hmaster2 & ~n40078;
  assign n40080 = ~n12193 & ~n40079;
  assign n40081 = ~controllable_hgrant3 & ~n40080;
  assign n40082 = ~n12163 & ~n40081;
  assign n40083 = controllable_nhgrant0 & ~n40082;
  assign n40084 = ~n12249 & ~n40083;
  assign n40085 = ~n3281 & ~n40084;
  assign n40086 = ~n4089 & ~n40085;
  assign n40087 = n3378 & ~n40086;
  assign n40088 = controllable_hmaster1 & ~n37877;
  assign n40089 = ~n6762 & ~n39706;
  assign n40090 = ~controllable_hmaster0 & ~n40089;
  assign n40091 = ~n37878 & ~n40090;
  assign n40092 = ~controllable_hmaster1 & ~n40091;
  assign n40093 = ~n40088 & ~n40092;
  assign n40094 = i_hbusreq3 & ~n40093;
  assign n40095 = ~n6772 & ~n39716;
  assign n40096 = controllable_hmaster1 & ~n40095;
  assign n40097 = controllable_hmaster0 & ~n40095;
  assign n40098 = ~n6772 & ~n39724;
  assign n40099 = ~controllable_hmaster0 & ~n40098;
  assign n40100 = ~n40097 & ~n40099;
  assign n40101 = ~controllable_hmaster1 & ~n40100;
  assign n40102 = ~n40096 & ~n40101;
  assign n40103 = ~i_hbusreq3 & ~n40102;
  assign n40104 = ~n40094 & ~n40103;
  assign n40105 = controllable_hmaster2 & ~n40104;
  assign n40106 = ~n35697 & ~n37878;
  assign n40107 = controllable_hmaster1 & ~n40106;
  assign n40108 = ~n35704 & ~n40107;
  assign n40109 = i_hbusreq3 & ~n40108;
  assign n40110 = ~n6772 & ~n39740;
  assign n40111 = controllable_hmaster0 & ~n40110;
  assign n40112 = ~n35710 & ~n40111;
  assign n40113 = controllable_hmaster1 & ~n40112;
  assign n40114 = ~n35718 & ~n40113;
  assign n40115 = ~i_hbusreq3 & ~n40114;
  assign n40116 = ~n40109 & ~n40115;
  assign n40117 = ~controllable_hmaster2 & ~n40116;
  assign n40118 = ~n40105 & ~n40117;
  assign n40119 = ~controllable_hgrant3 & ~n40118;
  assign n40120 = ~n5861 & ~n40119;
  assign n40121 = controllable_nhgrant0 & ~n40120;
  assign n40122 = ~n6082 & ~n40121;
  assign n40123 = ~n3281 & ~n40122;
  assign n40124 = ~n4089 & ~n40123;
  assign n40125 = ~n3378 & ~n40124;
  assign n40126 = ~n40087 & ~n40125;
  assign n40127 = n3492 & ~n40126;
  assign n40128 = ~n3631 & ~n40127;
  assign n40129 = n3485 & ~n40128;
  assign n40130 = ~n3630 & ~n40129;
  assign n40131 = n3476 & ~n40130;
  assign n40132 = ~n40065 & ~n40131;
  assign n40133 = n3374 & ~n40132;
  assign n40134 = ~n40003 & ~n40133;
  assign n40135 = n3655 & ~n40134;
  assign n40136 = ~n4333 & ~n39768;
  assign n40137 = controllable_hmaster1 & ~n40136;
  assign n40138 = controllable_hmaster0 & ~n40136;
  assign n40139 = ~n34022 & ~n40138;
  assign n40140 = ~controllable_hmaster1 & ~n40139;
  assign n40141 = ~n40137 & ~n40140;
  assign n40142 = i_hbusreq3 & ~n40141;
  assign n40143 = ~n4340 & ~n39780;
  assign n40144 = controllable_hmaster1 & ~n40143;
  assign n40145 = controllable_hmaster0 & ~n40143;
  assign n40146 = ~n34040 & ~n40145;
  assign n40147 = ~controllable_hmaster1 & ~n40146;
  assign n40148 = ~n40144 & ~n40147;
  assign n40149 = ~i_hbusreq3 & ~n40148;
  assign n40150 = ~n40142 & ~n40149;
  assign n40151 = controllable_hmaster2 & ~n40150;
  assign n40152 = ~n6887 & ~n40151;
  assign n40153 = ~controllable_hgrant3 & ~n40152;
  assign n40154 = ~n5037 & ~n40153;
  assign n40155 = controllable_nhgrant0 & ~n40154;
  assign n40156 = ~n5245 & ~n40155;
  assign n40157 = ~n3281 & ~n40156;
  assign n40158 = ~n3783 & ~n40157;
  assign n40159 = ~n3378 & ~n40158;
  assign n40160 = ~n12026 & ~n40159;
  assign n40161 = n3492 & ~n40160;
  assign n40162 = ~n3631 & ~n40161;
  assign n40163 = n3485 & ~n40162;
  assign n40164 = ~n3630 & ~n40163;
  assign n40165 = ~n3374 & ~n40164;
  assign n40166 = ~n5291 & ~n37970;
  assign n40167 = controllable_hmaster1 & ~n40166;
  assign n40168 = ~n5305 & ~n40167;
  assign n40169 = i_hbusreq3 & ~n40168;
  assign n40170 = ~n5311 & ~n37983;
  assign n40171 = controllable_hmaster1 & ~n40170;
  assign n40172 = ~n5334 & ~n40171;
  assign n40173 = ~i_hbusreq3 & ~n40172;
  assign n40174 = ~n40169 & ~n40173;
  assign n40175 = ~controllable_hmaster2 & ~n40174;
  assign n40176 = ~n12065 & ~n40175;
  assign n40177 = ~controllable_hgrant3 & ~n40176;
  assign n40178 = ~n12041 & ~n40177;
  assign n40179 = controllable_nhgrant0 & ~n40178;
  assign n40180 = ~n12101 & ~n40179;
  assign n40181 = ~n3281 & ~n40180;
  assign n40182 = ~n3950 & ~n40181;
  assign n40183 = n3378 & ~n40182;
  assign n40184 = ~n4333 & ~n39823;
  assign n40185 = controllable_hmaster1 & ~n40184;
  assign n40186 = controllable_hmaster0 & ~n40184;
  assign n40187 = ~n4333 & ~n39828;
  assign n40188 = ~controllable_hmaster0 & ~n40187;
  assign n40189 = ~n40186 & ~n40188;
  assign n40190 = ~controllable_hmaster1 & ~n40189;
  assign n40191 = ~n40185 & ~n40190;
  assign n40192 = i_hbusreq3 & ~n40191;
  assign n40193 = ~n4340 & ~n39839;
  assign n40194 = controllable_hmaster1 & ~n40193;
  assign n40195 = controllable_hmaster0 & ~n40193;
  assign n40196 = ~n4340 & ~n39847;
  assign n40197 = ~controllable_hmaster0 & ~n40196;
  assign n40198 = ~n40195 & ~n40197;
  assign n40199 = ~controllable_hmaster1 & ~n40198;
  assign n40200 = ~n40194 & ~n40199;
  assign n40201 = ~i_hbusreq3 & ~n40200;
  assign n40202 = ~n40192 & ~n40201;
  assign n40203 = controllable_hmaster2 & ~n40202;
  assign n40204 = ~n35804 & ~n37970;
  assign n40205 = controllable_hmaster1 & ~n40204;
  assign n40206 = ~n35811 & ~n40205;
  assign n40207 = i_hbusreq3 & ~n40206;
  assign n40208 = ~n35817 & ~n37983;
  assign n40209 = controllable_hmaster1 & ~n40208;
  assign n40210 = ~n35825 & ~n40209;
  assign n40211 = ~i_hbusreq3 & ~n40210;
  assign n40212 = ~n40207 & ~n40211;
  assign n40213 = ~controllable_hmaster2 & ~n40212;
  assign n40214 = ~n40203 & ~n40213;
  assign n40215 = ~controllable_hgrant3 & ~n40214;
  assign n40216 = ~n5402 & ~n40215;
  assign n40217 = controllable_nhgrant0 & ~n40216;
  assign n40218 = ~n5534 & ~n40217;
  assign n40219 = ~n3281 & ~n40218;
  assign n40220 = ~n3950 & ~n40219;
  assign n40221 = ~n3378 & ~n40220;
  assign n40222 = ~n40183 & ~n40221;
  assign n40223 = n3492 & ~n40222;
  assign n40224 = ~n3631 & ~n40223;
  assign n40225 = n3485 & ~n40224;
  assign n40226 = ~n3630 & ~n40225;
  assign n40227 = ~n3476 & ~n40226;
  assign n40228 = ~n6738 & ~n39881;
  assign n40229 = controllable_hmaster0 & ~n40228;
  assign n40230 = ~n5688 & ~n40229;
  assign n40231 = controllable_hmaster1 & ~n40230;
  assign n40232 = ~n5704 & ~n40231;
  assign n40233 = i_hbusreq3 & ~n40232;
  assign n40234 = ~n6745 & ~n39892;
  assign n40235 = controllable_hmaster0 & ~n40234;
  assign n40236 = ~n12210 & ~n40235;
  assign n40237 = controllable_hmaster1 & ~n40236;
  assign n40238 = ~n12222 & ~n40237;
  assign n40239 = ~i_hbusreq3 & ~n40238;
  assign n40240 = ~n40233 & ~n40239;
  assign n40241 = ~controllable_hmaster2 & ~n40240;
  assign n40242 = ~n12193 & ~n40241;
  assign n40243 = ~controllable_hgrant3 & ~n40242;
  assign n40244 = ~n12163 & ~n40243;
  assign n40245 = controllable_nhgrant0 & ~n40244;
  assign n40246 = ~n12249 & ~n40245;
  assign n40247 = ~n3281 & ~n40246;
  assign n40248 = ~n4089 & ~n40247;
  assign n40249 = n3378 & ~n40248;
  assign n40250 = controllable_hmaster1 & ~n38031;
  assign n40251 = ~n6762 & ~n39911;
  assign n40252 = ~controllable_hmaster0 & ~n40251;
  assign n40253 = ~n38032 & ~n40252;
  assign n40254 = ~controllable_hmaster1 & ~n40253;
  assign n40255 = ~n40250 & ~n40254;
  assign n40256 = i_hbusreq3 & ~n40255;
  assign n40257 = ~n6772 & ~n39921;
  assign n40258 = controllable_hmaster1 & ~n40257;
  assign n40259 = controllable_hmaster0 & ~n40257;
  assign n40260 = ~n6772 & ~n39929;
  assign n40261 = ~controllable_hmaster0 & ~n40260;
  assign n40262 = ~n40259 & ~n40261;
  assign n40263 = ~controllable_hmaster1 & ~n40262;
  assign n40264 = ~n40258 & ~n40263;
  assign n40265 = ~i_hbusreq3 & ~n40264;
  assign n40266 = ~n40256 & ~n40265;
  assign n40267 = controllable_hmaster2 & ~n40266;
  assign n40268 = ~n35889 & ~n38032;
  assign n40269 = controllable_hmaster1 & ~n40268;
  assign n40270 = ~n35896 & ~n40269;
  assign n40271 = i_hbusreq3 & ~n40270;
  assign n40272 = ~n6772 & ~n39945;
  assign n40273 = controllable_hmaster0 & ~n40272;
  assign n40274 = ~n35902 & ~n40273;
  assign n40275 = controllable_hmaster1 & ~n40274;
  assign n40276 = ~n35910 & ~n40275;
  assign n40277 = ~i_hbusreq3 & ~n40276;
  assign n40278 = ~n40271 & ~n40277;
  assign n40279 = ~controllable_hmaster2 & ~n40278;
  assign n40280 = ~n40267 & ~n40279;
  assign n40281 = ~controllable_hgrant3 & ~n40280;
  assign n40282 = ~n5861 & ~n40281;
  assign n40283 = controllable_nhgrant0 & ~n40282;
  assign n40284 = ~n6082 & ~n40283;
  assign n40285 = ~n3281 & ~n40284;
  assign n40286 = ~n4089 & ~n40285;
  assign n40287 = ~n3378 & ~n40286;
  assign n40288 = ~n40249 & ~n40287;
  assign n40289 = n3492 & ~n40288;
  assign n40290 = ~n3631 & ~n40289;
  assign n40291 = n3485 & ~n40290;
  assign n40292 = ~n3630 & ~n40291;
  assign n40293 = n3476 & ~n40292;
  assign n40294 = ~n40227 & ~n40293;
  assign n40295 = n3374 & ~n40294;
  assign n40296 = ~n40165 & ~n40295;
  assign n40297 = ~n3655 & ~n40296;
  assign n40298 = ~n40135 & ~n40297;
  assign n40299 = ~n3652 & ~n40298;
  assign n40300 = ~n39973 & ~n40299;
  assign n40301 = ~n3368 & ~n40300;
  assign n40302 = controllable_hmaster0 & ~n39564;
  assign n40303 = ~controllable_hmaster1 & ~n40302;
  assign n40304 = ~n39563 & ~n40303;
  assign n40305 = i_hbusreq3 & ~n40304;
  assign n40306 = controllable_hmaster0 & ~n39576;
  assign n40307 = ~controllable_hmaster1 & ~n40306;
  assign n40308 = ~n39575 & ~n40307;
  assign n40309 = ~i_hbusreq3 & ~n40308;
  assign n40310 = ~n40305 & ~n40309;
  assign n40311 = controllable_hmaster2 & ~n40310;
  assign n40312 = controllable_hmaster2 & ~n40311;
  assign n40313 = ~controllable_hgrant3 & ~n40312;
  assign n40314 = ~n7090 & ~n40313;
  assign n40315 = controllable_nhgrant0 & ~n40314;
  assign n40316 = ~n7118 & ~n40315;
  assign n40317 = ~n3281 & ~n40316;
  assign n40318 = ~n3281 & ~n40317;
  assign n40319 = ~n3378 & ~n40318;
  assign n40320 = ~n7082 & ~n40319;
  assign n40321 = n3492 & ~n40320;
  assign n40322 = n3492 & ~n40321;
  assign n40323 = n3485 & ~n40322;
  assign n40324 = n3485 & ~n40323;
  assign n40325 = ~n3374 & ~n40324;
  assign n40326 = ~n5291 & ~n38141;
  assign n40327 = controllable_hmaster1 & ~n40326;
  assign n40328 = ~n5305 & ~n40327;
  assign n40329 = i_hbusreq3 & ~n40328;
  assign n40330 = ~n5311 & ~n38161;
  assign n40331 = controllable_hmaster1 & ~n40330;
  assign n40332 = ~n5334 & ~n40331;
  assign n40333 = ~i_hbusreq3 & ~n40332;
  assign n40334 = ~n40329 & ~n40333;
  assign n40335 = ~controllable_hmaster2 & ~n40334;
  assign n40336 = ~n12741 & ~n40335;
  assign n40337 = ~controllable_hgrant3 & ~n40336;
  assign n40338 = ~n12731 & ~n40337;
  assign n40339 = controllable_nhgrant0 & ~n40338;
  assign n40340 = ~n12773 & ~n40339;
  assign n40341 = ~n3281 & ~n40340;
  assign n40342 = ~n3281 & ~n40341;
  assign n40343 = n3378 & ~n40342;
  assign n40344 = ~n39564 & ~n39623;
  assign n40345 = ~controllable_hmaster1 & ~n40344;
  assign n40346 = ~n39563 & ~n40345;
  assign n40347 = i_hbusreq3 & ~n40346;
  assign n40348 = ~n39576 & ~n39642;
  assign n40349 = ~controllable_hmaster1 & ~n40348;
  assign n40350 = ~n39575 & ~n40349;
  assign n40351 = ~i_hbusreq3 & ~n40350;
  assign n40352 = ~n40347 & ~n40351;
  assign n40353 = controllable_hmaster2 & ~n40352;
  assign n40354 = ~n35055 & ~n38141;
  assign n40355 = controllable_hmaster1 & ~n40354;
  assign n40356 = ~n35064 & ~n40355;
  assign n40357 = i_hbusreq3 & ~n40356;
  assign n40358 = ~n35074 & ~n38161;
  assign n40359 = controllable_hmaster1 & ~n40358;
  assign n40360 = ~n35091 & ~n40359;
  assign n40361 = ~i_hbusreq3 & ~n40360;
  assign n40362 = ~n40357 & ~n40361;
  assign n40363 = ~controllable_hmaster2 & ~n40362;
  assign n40364 = ~n40353 & ~n40363;
  assign n40365 = ~controllable_hgrant3 & ~n40364;
  assign n40366 = ~n12785 & ~n40365;
  assign n40367 = controllable_nhgrant0 & ~n40366;
  assign n40368 = ~n12827 & ~n40367;
  assign n40369 = ~n3281 & ~n40368;
  assign n40370 = ~n3281 & ~n40369;
  assign n40371 = ~n3378 & ~n40370;
  assign n40372 = ~n40343 & ~n40371;
  assign n40373 = n3492 & ~n40372;
  assign n40374 = n3492 & ~n40373;
  assign n40375 = n3485 & ~n40374;
  assign n40376 = n3485 & ~n40375;
  assign n40377 = ~n3476 & ~n40376;
  assign n40378 = controllable_hgrant4 & ~n7394;
  assign n40379 = ~n7255 & ~n40378;
  assign n40380 = ~controllable_hgrant2 & ~n40379;
  assign n40381 = ~n5616 & ~n40380;
  assign n40382 = controllable_hmaster0 & ~n40381;
  assign n40383 = ~n7328 & ~n40382;
  assign n40384 = controllable_hmaster1 & ~n40383;
  assign n40385 = ~n7342 & ~n40384;
  assign n40386 = i_hbusreq3 & ~n40385;
  assign n40387 = i_hbusreq2 & ~n40379;
  assign n40388 = controllable_hgrant4 & ~n7415;
  assign n40389 = ~n7308 & ~n40388;
  assign n40390 = ~i_hbusreq2 & ~n40389;
  assign n40391 = ~n40387 & ~n40390;
  assign n40392 = ~controllable_hgrant2 & ~n40391;
  assign n40393 = ~n7290 & ~n40392;
  assign n40394 = controllable_hmaster0 & ~n40393;
  assign n40395 = ~n12906 & ~n40394;
  assign n40396 = controllable_hmaster1 & ~n40395;
  assign n40397 = ~n12918 & ~n40396;
  assign n40398 = ~i_hbusreq3 & ~n40397;
  assign n40399 = ~n40386 & ~n40398;
  assign n40400 = ~controllable_hmaster2 & ~n40399;
  assign n40401 = ~n12884 & ~n40400;
  assign n40402 = ~controllable_hgrant3 & ~n40401;
  assign n40403 = ~n12856 & ~n40402;
  assign n40404 = controllable_nhgrant0 & ~n40403;
  assign n40405 = ~n12942 & ~n40404;
  assign n40406 = ~n3281 & ~n40405;
  assign n40407 = ~n3281 & ~n40406;
  assign n40408 = n3378 & ~n40407;
  assign n40409 = ~n7461 & ~n35144;
  assign n40410 = ~controllable_hgrant2 & ~n40409;
  assign n40411 = ~n5616 & ~n40410;
  assign n40412 = controllable_hmaster1 & ~n40411;
  assign n40413 = controllable_hmaster0 & ~n40411;
  assign n40414 = ~n7535 & ~n34195;
  assign n40415 = ~controllable_hgrant2 & ~n40414;
  assign n40416 = ~n5616 & ~n40415;
  assign n40417 = ~controllable_hmaster0 & ~n40416;
  assign n40418 = ~n40413 & ~n40417;
  assign n40419 = ~controllable_hmaster1 & ~n40418;
  assign n40420 = ~n40412 & ~n40419;
  assign n40421 = i_hbusreq3 & ~n40420;
  assign n40422 = i_hbusreq2 & ~n40409;
  assign n40423 = ~n7499 & ~n35234;
  assign n40424 = ~i_hbusreq2 & ~n40423;
  assign n40425 = ~n40422 & ~n40424;
  assign n40426 = ~controllable_hgrant2 & ~n40425;
  assign n40427 = ~n5862 & ~n40426;
  assign n40428 = controllable_hmaster1 & ~n40427;
  assign n40429 = controllable_hmaster0 & ~n40427;
  assign n40430 = i_hbusreq2 & ~n40414;
  assign n40431 = ~n7568 & ~n34214;
  assign n40432 = ~i_hbusreq2 & ~n40431;
  assign n40433 = ~n40430 & ~n40432;
  assign n40434 = ~controllable_hgrant2 & ~n40433;
  assign n40435 = ~n5862 & ~n40434;
  assign n40436 = ~controllable_hmaster0 & ~n40435;
  assign n40437 = ~n40429 & ~n40436;
  assign n40438 = ~controllable_hmaster1 & ~n40437;
  assign n40439 = ~n40428 & ~n40438;
  assign n40440 = ~i_hbusreq3 & ~n40439;
  assign n40441 = ~n40421 & ~n40440;
  assign n40442 = controllable_hmaster2 & ~n40441;
  assign n40443 = controllable_hgrant4 & ~n7631;
  assign n40444 = ~n7470 & ~n40443;
  assign n40445 = ~controllable_hgrant2 & ~n40444;
  assign n40446 = ~n5616 & ~n40445;
  assign n40447 = controllable_hmaster0 & ~n40446;
  assign n40448 = ~n7535 & ~n35144;
  assign n40449 = ~controllable_hgrant2 & ~n40448;
  assign n40450 = ~n5686 & ~n40449;
  assign n40451 = ~controllable_hmaster0 & ~n40450;
  assign n40452 = ~n40447 & ~n40451;
  assign n40453 = controllable_hmaster1 & ~n40452;
  assign n40454 = ~n7547 & ~n35144;
  assign n40455 = ~controllable_hgrant2 & ~n40454;
  assign n40456 = ~n5616 & ~n40455;
  assign n40457 = controllable_hmaster0 & ~n40456;
  assign n40458 = ~n5616 & ~n40449;
  assign n40459 = ~controllable_hmaster0 & ~n40458;
  assign n40460 = ~n40457 & ~n40459;
  assign n40461 = ~controllable_hmaster1 & ~n40460;
  assign n40462 = ~n40453 & ~n40461;
  assign n40463 = i_hbusreq3 & ~n40462;
  assign n40464 = i_hbusreq2 & ~n40444;
  assign n40465 = controllable_hgrant4 & ~n7651;
  assign n40466 = ~n7521 & ~n40465;
  assign n40467 = ~i_hbusreq2 & ~n40466;
  assign n40468 = ~n40464 & ~n40467;
  assign n40469 = ~controllable_hgrant2 & ~n40468;
  assign n40470 = ~n7507 & ~n40469;
  assign n40471 = controllable_hmaster0 & ~n40470;
  assign n40472 = i_hbusreq2 & ~n40448;
  assign n40473 = ~n7568 & ~n35234;
  assign n40474 = ~i_hbusreq2 & ~n40473;
  assign n40475 = ~n40472 & ~n40474;
  assign n40476 = ~controllable_hgrant2 & ~n40475;
  assign n40477 = ~n5950 & ~n40476;
  assign n40478 = ~controllable_hmaster0 & ~n40477;
  assign n40479 = ~n40471 & ~n40478;
  assign n40480 = controllable_hmaster1 & ~n40479;
  assign n40481 = i_hbusreq2 & ~n40454;
  assign n40482 = ~n7592 & ~n35234;
  assign n40483 = ~i_hbusreq2 & ~n40482;
  assign n40484 = ~n40481 & ~n40483;
  assign n40485 = ~controllable_hgrant2 & ~n40484;
  assign n40486 = ~n5862 & ~n40485;
  assign n40487 = controllable_hmaster0 & ~n40486;
  assign n40488 = ~n7614 & ~n35252;
  assign n40489 = ~i_hbusreq2 & ~n40488;
  assign n40490 = ~n40472 & ~n40489;
  assign n40491 = ~controllable_hgrant2 & ~n40490;
  assign n40492 = ~n5981 & ~n40491;
  assign n40493 = ~controllable_hmaster0 & ~n40492;
  assign n40494 = ~n40487 & ~n40493;
  assign n40495 = ~controllable_hmaster1 & ~n40494;
  assign n40496 = ~n40480 & ~n40495;
  assign n40497 = ~i_hbusreq3 & ~n40496;
  assign n40498 = ~n40463 & ~n40497;
  assign n40499 = ~controllable_hmaster2 & ~n40498;
  assign n40500 = ~n40442 & ~n40499;
  assign n40501 = ~controllable_hgrant3 & ~n40500;
  assign n40502 = ~n12974 & ~n40501;
  assign n40503 = controllable_nhgrant0 & ~n40502;
  assign n40504 = ~n13064 & ~n40503;
  assign n40505 = ~n3281 & ~n40504;
  assign n40506 = ~n3281 & ~n40505;
  assign n40507 = ~n3378 & ~n40506;
  assign n40508 = ~n40408 & ~n40507;
  assign n40509 = n3492 & ~n40508;
  assign n40510 = n3492 & ~n40509;
  assign n40511 = n3485 & ~n40510;
  assign n40512 = n3485 & ~n40511;
  assign n40513 = n3476 & ~n40512;
  assign n40514 = ~n40377 & ~n40513;
  assign n40515 = n3374 & ~n40514;
  assign n40516 = ~n40325 & ~n40515;
  assign n40517 = n3655 & ~n40516;
  assign n40518 = controllable_hmaster0 & ~n39771;
  assign n40519 = ~controllable_hmaster1 & ~n40518;
  assign n40520 = ~n39770 & ~n40519;
  assign n40521 = i_hbusreq3 & ~n40520;
  assign n40522 = controllable_hmaster0 & ~n39783;
  assign n40523 = ~controllable_hmaster1 & ~n40522;
  assign n40524 = ~n39782 & ~n40523;
  assign n40525 = ~i_hbusreq3 & ~n40524;
  assign n40526 = ~n40521 & ~n40525;
  assign n40527 = controllable_hmaster2 & ~n40526;
  assign n40528 = controllable_hmaster2 & ~n40527;
  assign n40529 = ~controllable_hgrant3 & ~n40528;
  assign n40530 = ~n7090 & ~n40529;
  assign n40531 = controllable_nhgrant0 & ~n40530;
  assign n40532 = ~n7118 & ~n40531;
  assign n40533 = ~n3281 & ~n40532;
  assign n40534 = ~n3281 & ~n40533;
  assign n40535 = ~n3378 & ~n40534;
  assign n40536 = ~n7082 & ~n40535;
  assign n40537 = n3492 & ~n40536;
  assign n40538 = n3492 & ~n40537;
  assign n40539 = n3485 & ~n40538;
  assign n40540 = n3485 & ~n40539;
  assign n40541 = ~n3374 & ~n40540;
  assign n40542 = ~n5291 & ~n38440;
  assign n40543 = controllable_hmaster1 & ~n40542;
  assign n40544 = ~n5305 & ~n40543;
  assign n40545 = i_hbusreq3 & ~n40544;
  assign n40546 = ~n5311 & ~n38460;
  assign n40547 = controllable_hmaster1 & ~n40546;
  assign n40548 = ~n5334 & ~n40547;
  assign n40549 = ~i_hbusreq3 & ~n40548;
  assign n40550 = ~n40545 & ~n40549;
  assign n40551 = ~controllable_hmaster2 & ~n40550;
  assign n40552 = ~n12741 & ~n40551;
  assign n40553 = ~controllable_hgrant3 & ~n40552;
  assign n40554 = ~n12731 & ~n40553;
  assign n40555 = controllable_nhgrant0 & ~n40554;
  assign n40556 = ~n12773 & ~n40555;
  assign n40557 = ~n3281 & ~n40556;
  assign n40558 = ~n3281 & ~n40557;
  assign n40559 = n3378 & ~n40558;
  assign n40560 = ~n39771 & ~n39830;
  assign n40561 = ~controllable_hmaster1 & ~n40560;
  assign n40562 = ~n39770 & ~n40561;
  assign n40563 = i_hbusreq3 & ~n40562;
  assign n40564 = ~n39783 & ~n39849;
  assign n40565 = ~controllable_hmaster1 & ~n40564;
  assign n40566 = ~n39782 & ~n40565;
  assign n40567 = ~i_hbusreq3 & ~n40566;
  assign n40568 = ~n40563 & ~n40567;
  assign n40569 = controllable_hmaster2 & ~n40568;
  assign n40570 = ~n35362 & ~n38440;
  assign n40571 = controllable_hmaster1 & ~n40570;
  assign n40572 = ~n35371 & ~n40571;
  assign n40573 = i_hbusreq3 & ~n40572;
  assign n40574 = ~n35382 & ~n38460;
  assign n40575 = controllable_hmaster1 & ~n40574;
  assign n40576 = ~n35400 & ~n40575;
  assign n40577 = ~i_hbusreq3 & ~n40576;
  assign n40578 = ~n40573 & ~n40577;
  assign n40579 = ~controllable_hmaster2 & ~n40578;
  assign n40580 = ~n40569 & ~n40579;
  assign n40581 = ~controllable_hgrant3 & ~n40580;
  assign n40582 = ~n12785 & ~n40581;
  assign n40583 = controllable_nhgrant0 & ~n40582;
  assign n40584 = ~n12827 & ~n40583;
  assign n40585 = ~n3281 & ~n40584;
  assign n40586 = ~n3281 & ~n40585;
  assign n40587 = ~n3378 & ~n40586;
  assign n40588 = ~n40559 & ~n40587;
  assign n40589 = n3492 & ~n40588;
  assign n40590 = n3492 & ~n40589;
  assign n40591 = n3485 & ~n40590;
  assign n40592 = n3485 & ~n40591;
  assign n40593 = ~n3476 & ~n40592;
  assign n40594 = ~n7750 & ~n40378;
  assign n40595 = ~controllable_hgrant2 & ~n40594;
  assign n40596 = ~n5616 & ~n40595;
  assign n40597 = controllable_hmaster0 & ~n40596;
  assign n40598 = ~n7328 & ~n40597;
  assign n40599 = controllable_hmaster1 & ~n40598;
  assign n40600 = ~n7342 & ~n40599;
  assign n40601 = i_hbusreq3 & ~n40600;
  assign n40602 = i_hbusreq2 & ~n40594;
  assign n40603 = ~n7771 & ~n40388;
  assign n40604 = ~i_hbusreq2 & ~n40603;
  assign n40605 = ~n40602 & ~n40604;
  assign n40606 = ~controllable_hgrant2 & ~n40605;
  assign n40607 = ~n7290 & ~n40606;
  assign n40608 = controllable_hmaster0 & ~n40607;
  assign n40609 = ~n12906 & ~n40608;
  assign n40610 = controllable_hmaster1 & ~n40609;
  assign n40611 = ~n12918 & ~n40610;
  assign n40612 = ~i_hbusreq3 & ~n40611;
  assign n40613 = ~n40601 & ~n40612;
  assign n40614 = ~controllable_hmaster2 & ~n40613;
  assign n40615 = ~n12884 & ~n40614;
  assign n40616 = ~controllable_hgrant3 & ~n40615;
  assign n40617 = ~n12856 & ~n40616;
  assign n40618 = controllable_nhgrant0 & ~n40617;
  assign n40619 = ~n12942 & ~n40618;
  assign n40620 = ~n3281 & ~n40619;
  assign n40621 = ~n3281 & ~n40620;
  assign n40622 = n3378 & ~n40621;
  assign n40623 = ~n7794 & ~n35144;
  assign n40624 = ~controllable_hgrant2 & ~n40623;
  assign n40625 = ~n5616 & ~n40624;
  assign n40626 = controllable_hmaster1 & ~n40625;
  assign n40627 = controllable_hmaster0 & ~n40625;
  assign n40628 = ~n7859 & ~n34195;
  assign n40629 = ~controllable_hgrant2 & ~n40628;
  assign n40630 = ~n5616 & ~n40629;
  assign n40631 = ~controllable_hmaster0 & ~n40630;
  assign n40632 = ~n40627 & ~n40631;
  assign n40633 = ~controllable_hmaster1 & ~n40632;
  assign n40634 = ~n40626 & ~n40633;
  assign n40635 = i_hbusreq3 & ~n40634;
  assign n40636 = i_hbusreq2 & ~n40623;
  assign n40637 = ~n7824 & ~n35234;
  assign n40638 = ~i_hbusreq2 & ~n40637;
  assign n40639 = ~n40636 & ~n40638;
  assign n40640 = ~controllable_hgrant2 & ~n40639;
  assign n40641 = ~n5862 & ~n40640;
  assign n40642 = controllable_hmaster1 & ~n40641;
  assign n40643 = controllable_hmaster0 & ~n40641;
  assign n40644 = i_hbusreq2 & ~n40628;
  assign n40645 = ~n7891 & ~n34214;
  assign n40646 = ~i_hbusreq2 & ~n40645;
  assign n40647 = ~n40644 & ~n40646;
  assign n40648 = ~controllable_hgrant2 & ~n40647;
  assign n40649 = ~n5862 & ~n40648;
  assign n40650 = ~controllable_hmaster0 & ~n40649;
  assign n40651 = ~n40643 & ~n40650;
  assign n40652 = ~controllable_hmaster1 & ~n40651;
  assign n40653 = ~n40642 & ~n40652;
  assign n40654 = ~i_hbusreq3 & ~n40653;
  assign n40655 = ~n40635 & ~n40654;
  assign n40656 = controllable_hmaster2 & ~n40655;
  assign n40657 = ~n7802 & ~n40443;
  assign n40658 = ~controllable_hgrant2 & ~n40657;
  assign n40659 = ~n5616 & ~n40658;
  assign n40660 = controllable_hmaster0 & ~n40659;
  assign n40661 = ~n7859 & ~n35144;
  assign n40662 = ~controllable_hgrant2 & ~n40661;
  assign n40663 = ~n5686 & ~n40662;
  assign n40664 = ~controllable_hmaster0 & ~n40663;
  assign n40665 = ~n40660 & ~n40664;
  assign n40666 = controllable_hmaster1 & ~n40665;
  assign n40667 = ~n7870 & ~n35144;
  assign n40668 = ~controllable_hgrant2 & ~n40667;
  assign n40669 = ~n5616 & ~n40668;
  assign n40670 = controllable_hmaster0 & ~n40669;
  assign n40671 = ~n5616 & ~n40662;
  assign n40672 = ~controllable_hmaster0 & ~n40671;
  assign n40673 = ~n40670 & ~n40672;
  assign n40674 = ~controllable_hmaster1 & ~n40673;
  assign n40675 = ~n40666 & ~n40674;
  assign n40676 = i_hbusreq3 & ~n40675;
  assign n40677 = i_hbusreq2 & ~n40657;
  assign n40678 = ~n7845 & ~n40465;
  assign n40679 = ~i_hbusreq2 & ~n40678;
  assign n40680 = ~n40677 & ~n40679;
  assign n40681 = ~controllable_hgrant2 & ~n40680;
  assign n40682 = ~n7507 & ~n40681;
  assign n40683 = controllable_hmaster0 & ~n40682;
  assign n40684 = i_hbusreq2 & ~n40661;
  assign n40685 = ~n7891 & ~n35234;
  assign n40686 = ~i_hbusreq2 & ~n40685;
  assign n40687 = ~n40684 & ~n40686;
  assign n40688 = ~controllable_hgrant2 & ~n40687;
  assign n40689 = ~n5950 & ~n40688;
  assign n40690 = ~controllable_hmaster0 & ~n40689;
  assign n40691 = ~n40683 & ~n40690;
  assign n40692 = controllable_hmaster1 & ~n40691;
  assign n40693 = i_hbusreq2 & ~n40667;
  assign n40694 = ~n7916 & ~n35234;
  assign n40695 = ~i_hbusreq2 & ~n40694;
  assign n40696 = ~n40693 & ~n40695;
  assign n40697 = ~controllable_hgrant2 & ~n40696;
  assign n40698 = ~n5862 & ~n40697;
  assign n40699 = controllable_hmaster0 & ~n40698;
  assign n40700 = ~n7930 & ~n35252;
  assign n40701 = ~i_hbusreq2 & ~n40700;
  assign n40702 = ~n40684 & ~n40701;
  assign n40703 = ~controllable_hgrant2 & ~n40702;
  assign n40704 = ~n5981 & ~n40703;
  assign n40705 = ~controllable_hmaster0 & ~n40704;
  assign n40706 = ~n40699 & ~n40705;
  assign n40707 = ~controllable_hmaster1 & ~n40706;
  assign n40708 = ~n40692 & ~n40707;
  assign n40709 = ~i_hbusreq3 & ~n40708;
  assign n40710 = ~n40676 & ~n40709;
  assign n40711 = ~controllable_hmaster2 & ~n40710;
  assign n40712 = ~n40656 & ~n40711;
  assign n40713 = ~controllable_hgrant3 & ~n40712;
  assign n40714 = ~n12974 & ~n40713;
  assign n40715 = controllable_nhgrant0 & ~n40714;
  assign n40716 = ~n13064 & ~n40715;
  assign n40717 = ~n3281 & ~n40716;
  assign n40718 = ~n3281 & ~n40717;
  assign n40719 = ~n3378 & ~n40718;
  assign n40720 = ~n40622 & ~n40719;
  assign n40721 = n3492 & ~n40720;
  assign n40722 = n3492 & ~n40721;
  assign n40723 = n3485 & ~n40722;
  assign n40724 = n3485 & ~n40723;
  assign n40725 = n3476 & ~n40724;
  assign n40726 = ~n40593 & ~n40725;
  assign n40727 = n3374 & ~n40726;
  assign n40728 = ~n40541 & ~n40727;
  assign n40729 = ~n3655 & ~n40728;
  assign n40730 = ~n40517 & ~n40729;
  assign n40731 = n3652 & ~n40730;
  assign n40732 = controllable_hmaster0 & ~n39976;
  assign n40733 = ~controllable_hmaster1 & ~n40732;
  assign n40734 = ~n39975 & ~n40733;
  assign n40735 = i_hbusreq3 & ~n40734;
  assign n40736 = controllable_hmaster0 & ~n39983;
  assign n40737 = ~controllable_hmaster1 & ~n40736;
  assign n40738 = ~n39982 & ~n40737;
  assign n40739 = ~i_hbusreq3 & ~n40738;
  assign n40740 = ~n40735 & ~n40739;
  assign n40741 = controllable_hmaster2 & ~n40740;
  assign n40742 = controllable_hmaster2 & ~n40741;
  assign n40743 = ~controllable_hgrant3 & ~n40742;
  assign n40744 = ~n7090 & ~n40743;
  assign n40745 = controllable_nhgrant0 & ~n40744;
  assign n40746 = ~n7118 & ~n40745;
  assign n40747 = ~n3281 & ~n40746;
  assign n40748 = ~n3281 & ~n40747;
  assign n40749 = ~n3378 & ~n40748;
  assign n40750 = ~n7082 & ~n40749;
  assign n40751 = n3492 & ~n40750;
  assign n40752 = n3492 & ~n40751;
  assign n40753 = n3485 & ~n40752;
  assign n40754 = n3485 & ~n40753;
  assign n40755 = ~n3374 & ~n40754;
  assign n40756 = ~n5291 & ~n38721;
  assign n40757 = controllable_hmaster1 & ~n40756;
  assign n40758 = ~n5305 & ~n40757;
  assign n40759 = i_hbusreq3 & ~n40758;
  assign n40760 = ~n5311 & ~n38734;
  assign n40761 = controllable_hmaster1 & ~n40760;
  assign n40762 = ~n5334 & ~n40761;
  assign n40763 = ~i_hbusreq3 & ~n40762;
  assign n40764 = ~n40759 & ~n40763;
  assign n40765 = ~controllable_hmaster2 & ~n40764;
  assign n40766 = ~n12741 & ~n40765;
  assign n40767 = ~controllable_hgrant3 & ~n40766;
  assign n40768 = ~n12731 & ~n40767;
  assign n40769 = controllable_nhgrant0 & ~n40768;
  assign n40770 = ~n12773 & ~n40769;
  assign n40771 = ~n3281 & ~n40770;
  assign n40772 = ~n3281 & ~n40771;
  assign n40773 = n3378 & ~n40772;
  assign n40774 = ~n39976 & ~n40026;
  assign n40775 = ~controllable_hmaster1 & ~n40774;
  assign n40776 = ~n39975 & ~n40775;
  assign n40777 = i_hbusreq3 & ~n40776;
  assign n40778 = ~n39983 & ~n40035;
  assign n40779 = ~controllable_hmaster1 & ~n40778;
  assign n40780 = ~n39982 & ~n40779;
  assign n40781 = ~i_hbusreq3 & ~n40780;
  assign n40782 = ~n40777 & ~n40781;
  assign n40783 = controllable_hmaster2 & ~n40782;
  assign n40784 = ~n35612 & ~n38721;
  assign n40785 = controllable_hmaster1 & ~n40784;
  assign n40786 = ~n35619 & ~n40785;
  assign n40787 = i_hbusreq3 & ~n40786;
  assign n40788 = ~n35625 & ~n38734;
  assign n40789 = controllable_hmaster1 & ~n40788;
  assign n40790 = ~n35633 & ~n40789;
  assign n40791 = ~i_hbusreq3 & ~n40790;
  assign n40792 = ~n40787 & ~n40791;
  assign n40793 = ~controllable_hmaster2 & ~n40792;
  assign n40794 = ~n40783 & ~n40793;
  assign n40795 = ~controllable_hgrant3 & ~n40794;
  assign n40796 = ~n12785 & ~n40795;
  assign n40797 = controllable_nhgrant0 & ~n40796;
  assign n40798 = ~n12827 & ~n40797;
  assign n40799 = ~n3281 & ~n40798;
  assign n40800 = ~n3281 & ~n40799;
  assign n40801 = ~n3378 & ~n40800;
  assign n40802 = ~n40773 & ~n40801;
  assign n40803 = n3492 & ~n40802;
  assign n40804 = n3492 & ~n40803;
  assign n40805 = n3485 & ~n40804;
  assign n40806 = n3485 & ~n40805;
  assign n40807 = ~n3476 & ~n40806;
  assign n40808 = ~n8029 & ~n40380;
  assign n40809 = controllable_hmaster0 & ~n40808;
  assign n40810 = ~n7328 & ~n40809;
  assign n40811 = controllable_hmaster1 & ~n40810;
  assign n40812 = ~n7342 & ~n40811;
  assign n40813 = i_hbusreq3 & ~n40812;
  assign n40814 = ~n8036 & ~n40392;
  assign n40815 = controllable_hmaster0 & ~n40814;
  assign n40816 = ~n12906 & ~n40815;
  assign n40817 = controllable_hmaster1 & ~n40816;
  assign n40818 = ~n12918 & ~n40817;
  assign n40819 = ~i_hbusreq3 & ~n40818;
  assign n40820 = ~n40813 & ~n40819;
  assign n40821 = ~controllable_hmaster2 & ~n40820;
  assign n40822 = ~n12884 & ~n40821;
  assign n40823 = ~controllable_hgrant3 & ~n40822;
  assign n40824 = ~n12856 & ~n40823;
  assign n40825 = controllable_nhgrant0 & ~n40824;
  assign n40826 = ~n12942 & ~n40825;
  assign n40827 = ~n3281 & ~n40826;
  assign n40828 = ~n3281 & ~n40827;
  assign n40829 = n3378 & ~n40828;
  assign n40830 = ~n6762 & ~n40410;
  assign n40831 = controllable_hmaster1 & ~n40830;
  assign n40832 = controllable_hmaster0 & ~n40830;
  assign n40833 = ~n6762 & ~n40415;
  assign n40834 = ~controllable_hmaster0 & ~n40833;
  assign n40835 = ~n40832 & ~n40834;
  assign n40836 = ~controllable_hmaster1 & ~n40835;
  assign n40837 = ~n40831 & ~n40836;
  assign n40838 = i_hbusreq3 & ~n40837;
  assign n40839 = ~n6772 & ~n40426;
  assign n40840 = controllable_hmaster1 & ~n40839;
  assign n40841 = controllable_hmaster0 & ~n40839;
  assign n40842 = ~n6772 & ~n40434;
  assign n40843 = ~controllable_hmaster0 & ~n40842;
  assign n40844 = ~n40841 & ~n40843;
  assign n40845 = ~controllable_hmaster1 & ~n40844;
  assign n40846 = ~n40840 & ~n40845;
  assign n40847 = ~i_hbusreq3 & ~n40846;
  assign n40848 = ~n40838 & ~n40847;
  assign n40849 = controllable_hmaster2 & ~n40848;
  assign n40850 = ~n8056 & ~n40445;
  assign n40851 = controllable_hmaster0 & ~n40850;
  assign n40852 = ~n6786 & ~n40449;
  assign n40853 = ~controllable_hmaster0 & ~n40852;
  assign n40854 = ~n40851 & ~n40853;
  assign n40855 = controllable_hmaster1 & ~n40854;
  assign n40856 = ~n6762 & ~n40455;
  assign n40857 = controllable_hmaster0 & ~n40856;
  assign n40858 = ~n6762 & ~n40449;
  assign n40859 = ~controllable_hmaster0 & ~n40858;
  assign n40860 = ~n40857 & ~n40859;
  assign n40861 = ~controllable_hmaster1 & ~n40860;
  assign n40862 = ~n40855 & ~n40861;
  assign n40863 = i_hbusreq3 & ~n40862;
  assign n40864 = ~n8066 & ~n40469;
  assign n40865 = controllable_hmaster0 & ~n40864;
  assign n40866 = ~n6813 & ~n40476;
  assign n40867 = ~controllable_hmaster0 & ~n40866;
  assign n40868 = ~n40865 & ~n40867;
  assign n40869 = controllable_hmaster1 & ~n40868;
  assign n40870 = ~n6772 & ~n40485;
  assign n40871 = controllable_hmaster0 & ~n40870;
  assign n40872 = ~n6831 & ~n40491;
  assign n40873 = ~controllable_hmaster0 & ~n40872;
  assign n40874 = ~n40871 & ~n40873;
  assign n40875 = ~controllable_hmaster1 & ~n40874;
  assign n40876 = ~n40869 & ~n40875;
  assign n40877 = ~i_hbusreq3 & ~n40876;
  assign n40878 = ~n40863 & ~n40877;
  assign n40879 = ~controllable_hmaster2 & ~n40878;
  assign n40880 = ~n40849 & ~n40879;
  assign n40881 = ~controllable_hgrant3 & ~n40880;
  assign n40882 = ~n12974 & ~n40881;
  assign n40883 = controllable_nhgrant0 & ~n40882;
  assign n40884 = ~n13064 & ~n40883;
  assign n40885 = ~n3281 & ~n40884;
  assign n40886 = ~n3281 & ~n40885;
  assign n40887 = ~n3378 & ~n40886;
  assign n40888 = ~n40829 & ~n40887;
  assign n40889 = n3492 & ~n40888;
  assign n40890 = n3492 & ~n40889;
  assign n40891 = n3485 & ~n40890;
  assign n40892 = n3485 & ~n40891;
  assign n40893 = n3476 & ~n40892;
  assign n40894 = ~n40807 & ~n40893;
  assign n40895 = n3374 & ~n40894;
  assign n40896 = ~n40755 & ~n40895;
  assign n40897 = n3655 & ~n40896;
  assign n40898 = controllable_hmaster0 & ~n40138;
  assign n40899 = ~controllable_hmaster1 & ~n40898;
  assign n40900 = ~n40137 & ~n40899;
  assign n40901 = i_hbusreq3 & ~n40900;
  assign n40902 = controllable_hmaster0 & ~n40145;
  assign n40903 = ~controllable_hmaster1 & ~n40902;
  assign n40904 = ~n40144 & ~n40903;
  assign n40905 = ~i_hbusreq3 & ~n40904;
  assign n40906 = ~n40901 & ~n40905;
  assign n40907 = controllable_hmaster2 & ~n40906;
  assign n40908 = controllable_hmaster2 & ~n40907;
  assign n40909 = ~controllable_hgrant3 & ~n40908;
  assign n40910 = ~n7090 & ~n40909;
  assign n40911 = controllable_nhgrant0 & ~n40910;
  assign n40912 = ~n7118 & ~n40911;
  assign n40913 = ~n3281 & ~n40912;
  assign n40914 = ~n3281 & ~n40913;
  assign n40915 = ~n3378 & ~n40914;
  assign n40916 = ~n7082 & ~n40915;
  assign n40917 = n3492 & ~n40916;
  assign n40918 = n3492 & ~n40917;
  assign n40919 = n3485 & ~n40918;
  assign n40920 = n3485 & ~n40919;
  assign n40921 = ~n3374 & ~n40920;
  assign n40922 = ~n5291 & ~n38930;
  assign n40923 = controllable_hmaster1 & ~n40922;
  assign n40924 = ~n5305 & ~n40923;
  assign n40925 = i_hbusreq3 & ~n40924;
  assign n40926 = ~n5311 & ~n38943;
  assign n40927 = controllable_hmaster1 & ~n40926;
  assign n40928 = ~n5334 & ~n40927;
  assign n40929 = ~i_hbusreq3 & ~n40928;
  assign n40930 = ~n40925 & ~n40929;
  assign n40931 = ~controllable_hmaster2 & ~n40930;
  assign n40932 = ~n12741 & ~n40931;
  assign n40933 = ~controllable_hgrant3 & ~n40932;
  assign n40934 = ~n12731 & ~n40933;
  assign n40935 = controllable_nhgrant0 & ~n40934;
  assign n40936 = ~n12773 & ~n40935;
  assign n40937 = ~n3281 & ~n40936;
  assign n40938 = ~n3281 & ~n40937;
  assign n40939 = n3378 & ~n40938;
  assign n40940 = ~n40138 & ~n40188;
  assign n40941 = ~controllable_hmaster1 & ~n40940;
  assign n40942 = ~n40137 & ~n40941;
  assign n40943 = i_hbusreq3 & ~n40942;
  assign n40944 = ~n40145 & ~n40197;
  assign n40945 = ~controllable_hmaster1 & ~n40944;
  assign n40946 = ~n40144 & ~n40945;
  assign n40947 = ~i_hbusreq3 & ~n40946;
  assign n40948 = ~n40943 & ~n40947;
  assign n40949 = controllable_hmaster2 & ~n40948;
  assign n40950 = ~n35804 & ~n38930;
  assign n40951 = controllable_hmaster1 & ~n40950;
  assign n40952 = ~n35811 & ~n40951;
  assign n40953 = i_hbusreq3 & ~n40952;
  assign n40954 = ~n35817 & ~n38943;
  assign n40955 = controllable_hmaster1 & ~n40954;
  assign n40956 = ~n35825 & ~n40955;
  assign n40957 = ~i_hbusreq3 & ~n40956;
  assign n40958 = ~n40953 & ~n40957;
  assign n40959 = ~controllable_hmaster2 & ~n40958;
  assign n40960 = ~n40949 & ~n40959;
  assign n40961 = ~controllable_hgrant3 & ~n40960;
  assign n40962 = ~n12785 & ~n40961;
  assign n40963 = controllable_nhgrant0 & ~n40962;
  assign n40964 = ~n12827 & ~n40963;
  assign n40965 = ~n3281 & ~n40964;
  assign n40966 = ~n3281 & ~n40965;
  assign n40967 = ~n3378 & ~n40966;
  assign n40968 = ~n40939 & ~n40967;
  assign n40969 = n3492 & ~n40968;
  assign n40970 = n3492 & ~n40969;
  assign n40971 = n3485 & ~n40970;
  assign n40972 = n3485 & ~n40971;
  assign n40973 = ~n3476 & ~n40972;
  assign n40974 = ~n8029 & ~n40595;
  assign n40975 = controllable_hmaster0 & ~n40974;
  assign n40976 = ~n7328 & ~n40975;
  assign n40977 = controllable_hmaster1 & ~n40976;
  assign n40978 = ~n7342 & ~n40977;
  assign n40979 = i_hbusreq3 & ~n40978;
  assign n40980 = ~n8036 & ~n40606;
  assign n40981 = controllable_hmaster0 & ~n40980;
  assign n40982 = ~n12906 & ~n40981;
  assign n40983 = controllable_hmaster1 & ~n40982;
  assign n40984 = ~n12918 & ~n40983;
  assign n40985 = ~i_hbusreq3 & ~n40984;
  assign n40986 = ~n40979 & ~n40985;
  assign n40987 = ~controllable_hmaster2 & ~n40986;
  assign n40988 = ~n12884 & ~n40987;
  assign n40989 = ~controllable_hgrant3 & ~n40988;
  assign n40990 = ~n12856 & ~n40989;
  assign n40991 = controllable_nhgrant0 & ~n40990;
  assign n40992 = ~n12942 & ~n40991;
  assign n40993 = ~n3281 & ~n40992;
  assign n40994 = ~n3281 & ~n40993;
  assign n40995 = n3378 & ~n40994;
  assign n40996 = ~n6762 & ~n40624;
  assign n40997 = controllable_hmaster1 & ~n40996;
  assign n40998 = controllable_hmaster0 & ~n40996;
  assign n40999 = ~n6762 & ~n40629;
  assign n41000 = ~controllable_hmaster0 & ~n40999;
  assign n41001 = ~n40998 & ~n41000;
  assign n41002 = ~controllable_hmaster1 & ~n41001;
  assign n41003 = ~n40997 & ~n41002;
  assign n41004 = i_hbusreq3 & ~n41003;
  assign n41005 = ~n6772 & ~n40640;
  assign n41006 = controllable_hmaster1 & ~n41005;
  assign n41007 = controllable_hmaster0 & ~n41005;
  assign n41008 = ~n6772 & ~n40648;
  assign n41009 = ~controllable_hmaster0 & ~n41008;
  assign n41010 = ~n41007 & ~n41009;
  assign n41011 = ~controllable_hmaster1 & ~n41010;
  assign n41012 = ~n41006 & ~n41011;
  assign n41013 = ~i_hbusreq3 & ~n41012;
  assign n41014 = ~n41004 & ~n41013;
  assign n41015 = controllable_hmaster2 & ~n41014;
  assign n41016 = ~n8056 & ~n40658;
  assign n41017 = controllable_hmaster0 & ~n41016;
  assign n41018 = ~n6786 & ~n40662;
  assign n41019 = ~controllable_hmaster0 & ~n41018;
  assign n41020 = ~n41017 & ~n41019;
  assign n41021 = controllable_hmaster1 & ~n41020;
  assign n41022 = ~n6762 & ~n40668;
  assign n41023 = controllable_hmaster0 & ~n41022;
  assign n41024 = ~n6762 & ~n40662;
  assign n41025 = ~controllable_hmaster0 & ~n41024;
  assign n41026 = ~n41023 & ~n41025;
  assign n41027 = ~controllable_hmaster1 & ~n41026;
  assign n41028 = ~n41021 & ~n41027;
  assign n41029 = i_hbusreq3 & ~n41028;
  assign n41030 = ~n8066 & ~n40681;
  assign n41031 = controllable_hmaster0 & ~n41030;
  assign n41032 = ~n6813 & ~n40688;
  assign n41033 = ~controllable_hmaster0 & ~n41032;
  assign n41034 = ~n41031 & ~n41033;
  assign n41035 = controllable_hmaster1 & ~n41034;
  assign n41036 = ~n6772 & ~n40697;
  assign n41037 = controllable_hmaster0 & ~n41036;
  assign n41038 = ~n6831 & ~n40703;
  assign n41039 = ~controllable_hmaster0 & ~n41038;
  assign n41040 = ~n41037 & ~n41039;
  assign n41041 = ~controllable_hmaster1 & ~n41040;
  assign n41042 = ~n41035 & ~n41041;
  assign n41043 = ~i_hbusreq3 & ~n41042;
  assign n41044 = ~n41029 & ~n41043;
  assign n41045 = ~controllable_hmaster2 & ~n41044;
  assign n41046 = ~n41015 & ~n41045;
  assign n41047 = ~controllable_hgrant3 & ~n41046;
  assign n41048 = ~n12974 & ~n41047;
  assign n41049 = controllable_nhgrant0 & ~n41048;
  assign n41050 = ~n13064 & ~n41049;
  assign n41051 = ~n3281 & ~n41050;
  assign n41052 = ~n3281 & ~n41051;
  assign n41053 = ~n3378 & ~n41052;
  assign n41054 = ~n40995 & ~n41053;
  assign n41055 = n3492 & ~n41054;
  assign n41056 = n3492 & ~n41055;
  assign n41057 = n3485 & ~n41056;
  assign n41058 = n3485 & ~n41057;
  assign n41059 = n3476 & ~n41058;
  assign n41060 = ~n40973 & ~n41059;
  assign n41061 = n3374 & ~n41060;
  assign n41062 = ~n40921 & ~n41061;
  assign n41063 = ~n3655 & ~n41062;
  assign n41064 = ~n40897 & ~n41063;
  assign n41065 = ~n3652 & ~n41064;
  assign n41066 = ~n40731 & ~n41065;
  assign n41067 = n3368 & ~n41066;
  assign n41068 = ~n40301 & ~n41067;
  assign n41069 = n3362 & ~n41068;
  assign n41070 = n3492 & ~n39589;
  assign n41071 = ~n3631 & ~n41070;
  assign n41072 = n3485 & ~n41071;
  assign n41073 = ~n3630 & ~n41072;
  assign n41074 = ~n3476 & ~n41073;
  assign n41075 = ~n8310 & ~n37006;
  assign n41076 = ~n3485 & ~n41075;
  assign n41077 = ~n41072 & ~n41076;
  assign n41078 = n3476 & ~n41077;
  assign n41079 = ~n41074 & ~n41078;
  assign n41080 = ~n3374 & ~n41079;
  assign n41081 = n3492 & ~n39665;
  assign n41082 = ~n3631 & ~n41081;
  assign n41083 = n3485 & ~n41082;
  assign n41084 = ~n3630 & ~n41083;
  assign n41085 = ~n3476 & ~n41084;
  assign n41086 = n3492 & ~n39755;
  assign n41087 = ~n3631 & ~n41086;
  assign n41088 = n3485 & ~n41087;
  assign n41089 = ~n41076 & ~n41088;
  assign n41090 = n3476 & ~n41089;
  assign n41091 = ~n41085 & ~n41090;
  assign n41092 = n3374 & ~n41091;
  assign n41093 = ~n41080 & ~n41092;
  assign n41094 = n3655 & ~n41093;
  assign n41095 = n3492 & ~n39796;
  assign n41096 = ~n3631 & ~n41095;
  assign n41097 = n3485 & ~n41096;
  assign n41098 = ~n3630 & ~n41097;
  assign n41099 = ~n3476 & ~n41098;
  assign n41100 = ~n8310 & ~n37048;
  assign n41101 = ~n3485 & ~n41100;
  assign n41102 = ~n41097 & ~n41101;
  assign n41103 = n3476 & ~n41102;
  assign n41104 = ~n41099 & ~n41103;
  assign n41105 = ~n3374 & ~n41104;
  assign n41106 = n3492 & ~n39872;
  assign n41107 = ~n3631 & ~n41106;
  assign n41108 = n3485 & ~n41107;
  assign n41109 = ~n3630 & ~n41108;
  assign n41110 = ~n3476 & ~n41109;
  assign n41111 = n3492 & ~n39960;
  assign n41112 = ~n3631 & ~n41111;
  assign n41113 = n3485 & ~n41112;
  assign n41114 = ~n41101 & ~n41113;
  assign n41115 = n3476 & ~n41114;
  assign n41116 = ~n41110 & ~n41115;
  assign n41117 = n3374 & ~n41116;
  assign n41118 = ~n41105 & ~n41117;
  assign n41119 = ~n3655 & ~n41118;
  assign n41120 = ~n41094 & ~n41119;
  assign n41121 = n3652 & ~n41120;
  assign n41122 = n3492 & ~n39996;
  assign n41123 = ~n3631 & ~n41122;
  assign n41124 = n3485 & ~n41123;
  assign n41125 = ~n3630 & ~n41124;
  assign n41126 = ~n3476 & ~n41125;
  assign n41127 = ~n8310 & ~n37091;
  assign n41128 = ~n3485 & ~n41127;
  assign n41129 = ~n41124 & ~n41128;
  assign n41130 = n3476 & ~n41129;
  assign n41131 = ~n41126 & ~n41130;
  assign n41132 = ~n3374 & ~n41131;
  assign n41133 = n3492 & ~n40058;
  assign n41134 = ~n3631 & ~n41133;
  assign n41135 = n3485 & ~n41134;
  assign n41136 = ~n3630 & ~n41135;
  assign n41137 = ~n3476 & ~n41136;
  assign n41138 = n3492 & ~n40124;
  assign n41139 = ~n3631 & ~n41138;
  assign n41140 = n3485 & ~n41139;
  assign n41141 = ~n41128 & ~n41140;
  assign n41142 = n3476 & ~n41141;
  assign n41143 = ~n41137 & ~n41142;
  assign n41144 = n3374 & ~n41143;
  assign n41145 = ~n41132 & ~n41144;
  assign n41146 = n3655 & ~n41145;
  assign n41147 = n3492 & ~n40158;
  assign n41148 = ~n3631 & ~n41147;
  assign n41149 = n3485 & ~n41148;
  assign n41150 = ~n3630 & ~n41149;
  assign n41151 = ~n3476 & ~n41150;
  assign n41152 = ~n8310 & ~n37132;
  assign n41153 = ~n3485 & ~n41152;
  assign n41154 = ~n41149 & ~n41153;
  assign n41155 = n3476 & ~n41154;
  assign n41156 = ~n41151 & ~n41155;
  assign n41157 = ~n3374 & ~n41156;
  assign n41158 = n3492 & ~n40220;
  assign n41159 = ~n3631 & ~n41158;
  assign n41160 = n3485 & ~n41159;
  assign n41161 = ~n3630 & ~n41160;
  assign n41162 = ~n3476 & ~n41161;
  assign n41163 = n3492 & ~n40286;
  assign n41164 = ~n3631 & ~n41163;
  assign n41165 = n3485 & ~n41164;
  assign n41166 = ~n41153 & ~n41165;
  assign n41167 = n3476 & ~n41166;
  assign n41168 = ~n41162 & ~n41167;
  assign n41169 = n3374 & ~n41168;
  assign n41170 = ~n41157 & ~n41169;
  assign n41171 = ~n3655 & ~n41170;
  assign n41172 = ~n41146 & ~n41171;
  assign n41173 = ~n3652 & ~n41172;
  assign n41174 = ~n41121 & ~n41173;
  assign n41175 = ~n3368 & ~n41174;
  assign n41176 = n3492 & ~n40318;
  assign n41177 = n3492 & ~n41176;
  assign n41178 = n3485 & ~n41177;
  assign n41179 = n3485 & ~n41178;
  assign n41180 = ~n3476 & ~n41179;
  assign n41181 = ~n8525 & ~n41178;
  assign n41182 = n3476 & ~n41181;
  assign n41183 = ~n41180 & ~n41182;
  assign n41184 = ~n3374 & ~n41183;
  assign n41185 = n3492 & ~n40370;
  assign n41186 = n3492 & ~n41185;
  assign n41187 = n3485 & ~n41186;
  assign n41188 = n3485 & ~n41187;
  assign n41189 = ~n3476 & ~n41188;
  assign n41190 = ~n3492 & ~n37174;
  assign n41191 = ~n3485 & ~n41190;
  assign n41192 = n3492 & ~n40506;
  assign n41193 = n3492 & ~n41192;
  assign n41194 = n3485 & ~n41193;
  assign n41195 = ~n41191 & ~n41194;
  assign n41196 = n3476 & ~n41195;
  assign n41197 = ~n41189 & ~n41196;
  assign n41198 = n3374 & ~n41197;
  assign n41199 = ~n41184 & ~n41198;
  assign n41200 = n3655 & ~n41199;
  assign n41201 = n3492 & ~n40534;
  assign n41202 = n3492 & ~n41201;
  assign n41203 = n3485 & ~n41202;
  assign n41204 = n3485 & ~n41203;
  assign n41205 = ~n3476 & ~n41204;
  assign n41206 = ~n8525 & ~n41203;
  assign n41207 = n3476 & ~n41206;
  assign n41208 = ~n41205 & ~n41207;
  assign n41209 = ~n3374 & ~n41208;
  assign n41210 = n3492 & ~n40586;
  assign n41211 = n3492 & ~n41210;
  assign n41212 = n3485 & ~n41211;
  assign n41213 = n3485 & ~n41212;
  assign n41214 = ~n3476 & ~n41213;
  assign n41215 = ~n3492 & ~n37202;
  assign n41216 = ~n3485 & ~n41215;
  assign n41217 = n3492 & ~n40718;
  assign n41218 = n3492 & ~n41217;
  assign n41219 = n3485 & ~n41218;
  assign n41220 = ~n41216 & ~n41219;
  assign n41221 = n3476 & ~n41220;
  assign n41222 = ~n41214 & ~n41221;
  assign n41223 = n3374 & ~n41222;
  assign n41224 = ~n41209 & ~n41223;
  assign n41225 = ~n3655 & ~n41224;
  assign n41226 = ~n41200 & ~n41225;
  assign n41227 = n3652 & ~n41226;
  assign n41228 = n3492 & ~n40748;
  assign n41229 = n3492 & ~n41228;
  assign n41230 = n3485 & ~n41229;
  assign n41231 = n3485 & ~n41230;
  assign n41232 = ~n3476 & ~n41231;
  assign n41233 = ~n8525 & ~n41230;
  assign n41234 = n3476 & ~n41233;
  assign n41235 = ~n41232 & ~n41234;
  assign n41236 = ~n3374 & ~n41235;
  assign n41237 = n3492 & ~n40800;
  assign n41238 = n3492 & ~n41237;
  assign n41239 = n3485 & ~n41238;
  assign n41240 = n3485 & ~n41239;
  assign n41241 = ~n3476 & ~n41240;
  assign n41242 = ~n3492 & ~n37231;
  assign n41243 = ~n3485 & ~n41242;
  assign n41244 = n3492 & ~n40886;
  assign n41245 = n3492 & ~n41244;
  assign n41246 = n3485 & ~n41245;
  assign n41247 = ~n41243 & ~n41246;
  assign n41248 = n3476 & ~n41247;
  assign n41249 = ~n41241 & ~n41248;
  assign n41250 = n3374 & ~n41249;
  assign n41251 = ~n41236 & ~n41250;
  assign n41252 = n3655 & ~n41251;
  assign n41253 = n3492 & ~n40914;
  assign n41254 = n3492 & ~n41253;
  assign n41255 = n3485 & ~n41254;
  assign n41256 = n3485 & ~n41255;
  assign n41257 = ~n3476 & ~n41256;
  assign n41258 = ~n8525 & ~n41255;
  assign n41259 = n3476 & ~n41258;
  assign n41260 = ~n41257 & ~n41259;
  assign n41261 = ~n3374 & ~n41260;
  assign n41262 = n3492 & ~n40966;
  assign n41263 = n3492 & ~n41262;
  assign n41264 = n3485 & ~n41263;
  assign n41265 = n3485 & ~n41264;
  assign n41266 = ~n3476 & ~n41265;
  assign n41267 = ~n3492 & ~n37258;
  assign n41268 = ~n3485 & ~n41267;
  assign n41269 = n3492 & ~n41052;
  assign n41270 = n3492 & ~n41269;
  assign n41271 = n3485 & ~n41270;
  assign n41272 = ~n41268 & ~n41271;
  assign n41273 = n3476 & ~n41272;
  assign n41274 = ~n41266 & ~n41273;
  assign n41275 = n3374 & ~n41274;
  assign n41276 = ~n41261 & ~n41275;
  assign n41277 = ~n3655 & ~n41276;
  assign n41278 = ~n41252 & ~n41277;
  assign n41279 = ~n3652 & ~n41278;
  assign n41280 = ~n41227 & ~n41279;
  assign n41281 = n3368 & ~n41280;
  assign n41282 = ~n41175 & ~n41281;
  assign n41283 = ~n3362 & ~n41282;
  assign n41284 = ~n41069 & ~n41283;
  assign n41285 = n3359 & ~n41284;
  assign n41286 = ~n37278 & ~n41072;
  assign n41287 = n3476 & ~n41286;
  assign n41288 = ~n41074 & ~n41287;
  assign n41289 = ~n3374 & ~n41288;
  assign n41290 = ~n37278 & ~n41088;
  assign n41291 = n3476 & ~n41290;
  assign n41292 = ~n41085 & ~n41291;
  assign n41293 = n3374 & ~n41292;
  assign n41294 = ~n41289 & ~n41293;
  assign n41295 = n3655 & ~n41294;
  assign n41296 = ~n37289 & ~n41097;
  assign n41297 = n3476 & ~n41296;
  assign n41298 = ~n41099 & ~n41297;
  assign n41299 = ~n3374 & ~n41298;
  assign n41300 = ~n37289 & ~n41113;
  assign n41301 = n3476 & ~n41300;
  assign n41302 = ~n41110 & ~n41301;
  assign n41303 = n3374 & ~n41302;
  assign n41304 = ~n41299 & ~n41303;
  assign n41305 = ~n3655 & ~n41304;
  assign n41306 = ~n41295 & ~n41305;
  assign n41307 = n3652 & ~n41306;
  assign n41308 = ~n37302 & ~n41124;
  assign n41309 = n3476 & ~n41308;
  assign n41310 = ~n41126 & ~n41309;
  assign n41311 = ~n3374 & ~n41310;
  assign n41312 = ~n37302 & ~n41140;
  assign n41313 = n3476 & ~n41312;
  assign n41314 = ~n41137 & ~n41313;
  assign n41315 = n3374 & ~n41314;
  assign n41316 = ~n41311 & ~n41315;
  assign n41317 = n3655 & ~n41316;
  assign n41318 = ~n37313 & ~n41149;
  assign n41319 = n3476 & ~n41318;
  assign n41320 = ~n41151 & ~n41319;
  assign n41321 = ~n3374 & ~n41320;
  assign n41322 = ~n37313 & ~n41165;
  assign n41323 = n3476 & ~n41322;
  assign n41324 = ~n41162 & ~n41323;
  assign n41325 = n3374 & ~n41324;
  assign n41326 = ~n41321 & ~n41325;
  assign n41327 = ~n3655 & ~n41326;
  assign n41328 = ~n41317 & ~n41327;
  assign n41329 = ~n3652 & ~n41328;
  assign n41330 = ~n41307 & ~n41329;
  assign n41331 = ~n3368 & ~n41330;
  assign n41332 = ~n8689 & ~n41178;
  assign n41333 = n3476 & ~n41332;
  assign n41334 = ~n41180 & ~n41333;
  assign n41335 = ~n3374 & ~n41334;
  assign n41336 = ~n37332 & ~n41194;
  assign n41337 = n3476 & ~n41336;
  assign n41338 = ~n41189 & ~n41337;
  assign n41339 = n3374 & ~n41338;
  assign n41340 = ~n41335 & ~n41339;
  assign n41341 = n3655 & ~n41340;
  assign n41342 = ~n8689 & ~n41203;
  assign n41343 = n3476 & ~n41342;
  assign n41344 = ~n41205 & ~n41343;
  assign n41345 = ~n3374 & ~n41344;
  assign n41346 = ~n37343 & ~n41219;
  assign n41347 = n3476 & ~n41346;
  assign n41348 = ~n41214 & ~n41347;
  assign n41349 = n3374 & ~n41348;
  assign n41350 = ~n41345 & ~n41349;
  assign n41351 = ~n3655 & ~n41350;
  assign n41352 = ~n41341 & ~n41351;
  assign n41353 = n3652 & ~n41352;
  assign n41354 = ~n8689 & ~n41230;
  assign n41355 = n3476 & ~n41354;
  assign n41356 = ~n41232 & ~n41355;
  assign n41357 = ~n3374 & ~n41356;
  assign n41358 = ~n37356 & ~n41246;
  assign n41359 = n3476 & ~n41358;
  assign n41360 = ~n41241 & ~n41359;
  assign n41361 = n3374 & ~n41360;
  assign n41362 = ~n41357 & ~n41361;
  assign n41363 = n3655 & ~n41362;
  assign n41364 = ~n8689 & ~n41255;
  assign n41365 = n3476 & ~n41364;
  assign n41366 = ~n41257 & ~n41365;
  assign n41367 = ~n3374 & ~n41366;
  assign n41368 = ~n37367 & ~n41271;
  assign n41369 = n3476 & ~n41368;
  assign n41370 = ~n41266 & ~n41369;
  assign n41371 = n3374 & ~n41370;
  assign n41372 = ~n41367 & ~n41371;
  assign n41373 = ~n3655 & ~n41372;
  assign n41374 = ~n41363 & ~n41373;
  assign n41375 = ~n3652 & ~n41374;
  assign n41376 = ~n41353 & ~n41375;
  assign n41377 = n3368 & ~n41376;
  assign n41378 = ~n41331 & ~n41377;
  assign n41379 = n3362 & ~n41378;
  assign n41380 = n3378 & ~n39589;
  assign n41381 = ~n37398 & ~n41380;
  assign n41382 = n3492 & ~n41381;
  assign n41383 = ~n3631 & ~n41382;
  assign n41384 = n3485 & ~n41383;
  assign n41385 = ~n3630 & ~n41384;
  assign n41386 = ~n3476 & ~n41385;
  assign n41387 = ~n37006 & ~n41382;
  assign n41388 = n3485 & ~n41387;
  assign n41389 = ~n37278 & ~n41388;
  assign n41390 = n3476 & ~n41389;
  assign n41391 = ~n41386 & ~n41390;
  assign n41392 = ~n3374 & ~n41391;
  assign n41393 = n3378 & ~n39665;
  assign n41394 = ~n37472 & ~n41393;
  assign n41395 = n3492 & ~n41394;
  assign n41396 = ~n3631 & ~n41395;
  assign n41397 = n3485 & ~n41396;
  assign n41398 = ~n3630 & ~n41397;
  assign n41399 = ~n3476 & ~n41398;
  assign n41400 = n3378 & ~n39755;
  assign n41401 = ~n37554 & ~n41400;
  assign n41402 = n3492 & ~n41401;
  assign n41403 = ~n37006 & ~n41402;
  assign n41404 = n3485 & ~n41403;
  assign n41405 = ~n37278 & ~n41404;
  assign n41406 = n3476 & ~n41405;
  assign n41407 = ~n41399 & ~n41406;
  assign n41408 = n3374 & ~n41407;
  assign n41409 = ~n41392 & ~n41408;
  assign n41410 = n3655 & ~n41409;
  assign n41411 = n3378 & ~n39796;
  assign n41412 = ~n37588 & ~n41411;
  assign n41413 = n3492 & ~n41412;
  assign n41414 = ~n3631 & ~n41413;
  assign n41415 = n3485 & ~n41414;
  assign n41416 = ~n3630 & ~n41415;
  assign n41417 = ~n3476 & ~n41416;
  assign n41418 = ~n37048 & ~n41413;
  assign n41419 = n3485 & ~n41418;
  assign n41420 = ~n37289 & ~n41419;
  assign n41421 = n3476 & ~n41420;
  assign n41422 = ~n41417 & ~n41421;
  assign n41423 = ~n3374 & ~n41422;
  assign n41424 = n3378 & ~n39872;
  assign n41425 = ~n37666 & ~n41424;
  assign n41426 = n3492 & ~n41425;
  assign n41427 = ~n3631 & ~n41426;
  assign n41428 = n3485 & ~n41427;
  assign n41429 = ~n3630 & ~n41428;
  assign n41430 = ~n3476 & ~n41429;
  assign n41431 = n3378 & ~n39960;
  assign n41432 = ~n37757 & ~n41431;
  assign n41433 = n3492 & ~n41432;
  assign n41434 = ~n37048 & ~n41433;
  assign n41435 = n3485 & ~n41434;
  assign n41436 = ~n37289 & ~n41435;
  assign n41437 = n3476 & ~n41436;
  assign n41438 = ~n41430 & ~n41437;
  assign n41439 = n3374 & ~n41438;
  assign n41440 = ~n41423 & ~n41439;
  assign n41441 = ~n3655 & ~n41440;
  assign n41442 = ~n41410 & ~n41441;
  assign n41443 = n3652 & ~n41442;
  assign n41444 = n3378 & ~n39996;
  assign n41445 = ~n37791 & ~n41444;
  assign n41446 = n3492 & ~n41445;
  assign n41447 = ~n3631 & ~n41446;
  assign n41448 = n3485 & ~n41447;
  assign n41449 = ~n3630 & ~n41448;
  assign n41450 = ~n3476 & ~n41449;
  assign n41451 = ~n37091 & ~n41446;
  assign n41452 = n3485 & ~n41451;
  assign n41453 = ~n37302 & ~n41452;
  assign n41454 = n3476 & ~n41453;
  assign n41455 = ~n41450 & ~n41454;
  assign n41456 = ~n3374 & ~n41455;
  assign n41457 = n3378 & ~n40058;
  assign n41458 = ~n37851 & ~n41457;
  assign n41459 = n3492 & ~n41458;
  assign n41460 = ~n3631 & ~n41459;
  assign n41461 = n3485 & ~n41460;
  assign n41462 = ~n3630 & ~n41461;
  assign n41463 = ~n3476 & ~n41462;
  assign n41464 = n3378 & ~n40124;
  assign n41465 = ~n37913 & ~n41464;
  assign n41466 = n3492 & ~n41465;
  assign n41467 = ~n37091 & ~n41466;
  assign n41468 = n3485 & ~n41467;
  assign n41469 = ~n37302 & ~n41468;
  assign n41470 = n3476 & ~n41469;
  assign n41471 = ~n41463 & ~n41470;
  assign n41472 = n3374 & ~n41471;
  assign n41473 = ~n41456 & ~n41472;
  assign n41474 = n3655 & ~n41473;
  assign n41475 = n3378 & ~n40158;
  assign n41476 = ~n37945 & ~n41475;
  assign n41477 = n3492 & ~n41476;
  assign n41478 = ~n3631 & ~n41477;
  assign n41479 = n3485 & ~n41478;
  assign n41480 = ~n3630 & ~n41479;
  assign n41481 = ~n3476 & ~n41480;
  assign n41482 = ~n37132 & ~n41477;
  assign n41483 = n3485 & ~n41482;
  assign n41484 = ~n37313 & ~n41483;
  assign n41485 = n3476 & ~n41484;
  assign n41486 = ~n41481 & ~n41485;
  assign n41487 = ~n3374 & ~n41486;
  assign n41488 = n3378 & ~n40220;
  assign n41489 = ~n38005 & ~n41488;
  assign n41490 = n3492 & ~n41489;
  assign n41491 = ~n3631 & ~n41490;
  assign n41492 = n3485 & ~n41491;
  assign n41493 = ~n3630 & ~n41492;
  assign n41494 = ~n3476 & ~n41493;
  assign n41495 = n3378 & ~n40286;
  assign n41496 = ~n38067 & ~n41495;
  assign n41497 = n3492 & ~n41496;
  assign n41498 = ~n37132 & ~n41497;
  assign n41499 = n3485 & ~n41498;
  assign n41500 = ~n37313 & ~n41499;
  assign n41501 = n3476 & ~n41500;
  assign n41502 = ~n41494 & ~n41501;
  assign n41503 = n3374 & ~n41502;
  assign n41504 = ~n41487 & ~n41503;
  assign n41505 = ~n3655 & ~n41504;
  assign n41506 = ~n41474 & ~n41505;
  assign n41507 = ~n3652 & ~n41506;
  assign n41508 = ~n41443 & ~n41507;
  assign n41509 = ~n3368 & ~n41508;
  assign n41510 = n3378 & ~n40318;
  assign n41511 = ~n38114 & ~n41510;
  assign n41512 = n3492 & ~n41511;
  assign n41513 = n3492 & ~n41512;
  assign n41514 = n3485 & ~n41513;
  assign n41515 = n3485 & ~n41514;
  assign n41516 = ~n3476 & ~n41515;
  assign n41517 = ~n8523 & ~n41512;
  assign n41518 = n3485 & ~n41517;
  assign n41519 = ~n8689 & ~n41518;
  assign n41520 = n3476 & ~n41519;
  assign n41521 = ~n41516 & ~n41520;
  assign n41522 = ~n3374 & ~n41521;
  assign n41523 = n3378 & ~n40370;
  assign n41524 = ~n38186 & ~n41523;
  assign n41525 = n3492 & ~n41524;
  assign n41526 = n3492 & ~n41525;
  assign n41527 = n3485 & ~n41526;
  assign n41528 = n3485 & ~n41527;
  assign n41529 = ~n3476 & ~n41528;
  assign n41530 = i_hlock4 & ~n9955;
  assign n41531 = ~i_hlock4 & ~n9959;
  assign n41532 = ~n41530 & ~n41531;
  assign n41533 = controllable_hgrant4 & ~n41532;
  assign n41534 = ~n9873 & ~n41533;
  assign n41535 = ~controllable_hgrant2 & ~n41534;
  assign n41536 = ~n5616 & ~n41535;
  assign n41537 = controllable_hmaster1 & ~n41536;
  assign n41538 = controllable_hmaster0 & ~n41536;
  assign n41539 = i_hlock4 & ~n10029;
  assign n41540 = ~i_hlock4 & ~n10033;
  assign n41541 = ~n41539 & ~n41540;
  assign n41542 = controllable_hgrant4 & ~n41541;
  assign n41543 = ~n5911 & ~n41542;
  assign n41544 = ~controllable_hgrant2 & ~n41543;
  assign n41545 = ~n5616 & ~n41544;
  assign n41546 = ~controllable_hmaster0 & ~n41545;
  assign n41547 = ~n41538 & ~n41546;
  assign n41548 = ~controllable_hmaster1 & ~n41547;
  assign n41549 = ~n41537 & ~n41548;
  assign n41550 = i_hbusreq3 & ~n41549;
  assign n41551 = i_hbusreq2 & ~n41534;
  assign n41552 = i_hbusreq4 & ~n41532;
  assign n41553 = i_hlock4 & ~n10847;
  assign n41554 = ~i_hlock4 & ~n10861;
  assign n41555 = ~n41553 & ~n41554;
  assign n41556 = ~i_hbusreq4 & ~n41555;
  assign n41557 = ~n41552 & ~n41556;
  assign n41558 = controllable_hgrant4 & ~n41557;
  assign n41559 = ~n9895 & ~n41558;
  assign n41560 = ~i_hbusreq2 & ~n41559;
  assign n41561 = ~n41551 & ~n41560;
  assign n41562 = ~controllable_hgrant2 & ~n41561;
  assign n41563 = ~n5862 & ~n41562;
  assign n41564 = controllable_hmaster1 & ~n41563;
  assign n41565 = controllable_hmaster0 & ~n41563;
  assign n41566 = i_hbusreq2 & ~n41543;
  assign n41567 = i_hbusreq4 & ~n41541;
  assign n41568 = i_hlock4 & ~n10949;
  assign n41569 = ~i_hlock4 & ~n10963;
  assign n41570 = ~n41568 & ~n41569;
  assign n41571 = ~i_hbusreq4 & ~n41570;
  assign n41572 = ~n41567 & ~n41571;
  assign n41573 = controllable_hgrant4 & ~n41572;
  assign n41574 = ~n5943 & ~n41573;
  assign n41575 = ~i_hbusreq2 & ~n41574;
  assign n41576 = ~n41566 & ~n41575;
  assign n41577 = ~controllable_hgrant2 & ~n41576;
  assign n41578 = ~n5862 & ~n41577;
  assign n41579 = ~controllable_hmaster0 & ~n41578;
  assign n41580 = ~n41565 & ~n41579;
  assign n41581 = ~controllable_hmaster1 & ~n41580;
  assign n41582 = ~n41564 & ~n41581;
  assign n41583 = ~i_hbusreq3 & ~n41582;
  assign n41584 = ~n41550 & ~n41583;
  assign n41585 = controllable_hmaster2 & ~n41584;
  assign n41586 = ~n5911 & ~n41533;
  assign n41587 = ~controllable_hgrant2 & ~n41586;
  assign n41588 = ~n5686 & ~n41587;
  assign n41589 = ~controllable_hmaster0 & ~n41588;
  assign n41590 = ~n38286 & ~n41589;
  assign n41591 = controllable_hmaster1 & ~n41590;
  assign n41592 = ~n5921 & ~n41533;
  assign n41593 = ~controllable_hgrant2 & ~n41592;
  assign n41594 = ~n5616 & ~n41593;
  assign n41595 = controllable_hmaster0 & ~n41594;
  assign n41596 = ~n5616 & ~n41587;
  assign n41597 = ~controllable_hmaster0 & ~n41596;
  assign n41598 = ~n41595 & ~n41597;
  assign n41599 = ~controllable_hmaster1 & ~n41598;
  assign n41600 = ~n41591 & ~n41599;
  assign n41601 = i_hbusreq3 & ~n41600;
  assign n41602 = i_hlock4 & ~n10883;
  assign n41603 = ~i_hlock4 & ~n10895;
  assign n41604 = ~n41602 & ~n41603;
  assign n41605 = ~i_hbusreq4 & ~n41604;
  assign n41606 = ~n36158 & ~n41605;
  assign n41607 = controllable_hgrant4 & ~n41606;
  assign n41608 = ~n9910 & ~n41607;
  assign n41609 = ~i_hbusreq2 & ~n41608;
  assign n41610 = ~n38291 & ~n41609;
  assign n41611 = ~controllable_hgrant2 & ~n41610;
  assign n41612 = ~n7507 & ~n41611;
  assign n41613 = controllable_hmaster0 & ~n41612;
  assign n41614 = i_hbusreq2 & ~n41586;
  assign n41615 = ~n5943 & ~n41558;
  assign n41616 = ~i_hbusreq2 & ~n41615;
  assign n41617 = ~n41614 & ~n41616;
  assign n41618 = ~controllable_hgrant2 & ~n41617;
  assign n41619 = ~n5950 & ~n41618;
  assign n41620 = ~controllable_hmaster0 & ~n41619;
  assign n41621 = ~n41613 & ~n41620;
  assign n41622 = controllable_hmaster1 & ~n41621;
  assign n41623 = i_hbusreq2 & ~n41592;
  assign n41624 = ~n5974 & ~n41558;
  assign n41625 = ~i_hbusreq2 & ~n41624;
  assign n41626 = ~n41623 & ~n41625;
  assign n41627 = ~controllable_hgrant2 & ~n41626;
  assign n41628 = ~n5862 & ~n41627;
  assign n41629 = controllable_hmaster0 & ~n41628;
  assign n41630 = i_hlock4 & ~n10983;
  assign n41631 = ~i_hlock4 & ~n10993;
  assign n41632 = ~n41630 & ~n41631;
  assign n41633 = ~i_hbusreq4 & ~n41632;
  assign n41634 = ~n41552 & ~n41633;
  assign n41635 = controllable_hgrant4 & ~n41634;
  assign n41636 = ~n5990 & ~n41635;
  assign n41637 = ~i_hbusreq2 & ~n41636;
  assign n41638 = ~n41614 & ~n41637;
  assign n41639 = ~controllable_hgrant2 & ~n41638;
  assign n41640 = ~n5981 & ~n41639;
  assign n41641 = ~controllable_hmaster0 & ~n41640;
  assign n41642 = ~n41629 & ~n41641;
  assign n41643 = ~controllable_hmaster1 & ~n41642;
  assign n41644 = ~n41622 & ~n41643;
  assign n41645 = ~i_hbusreq3 & ~n41644;
  assign n41646 = ~n41601 & ~n41645;
  assign n41647 = ~controllable_hmaster2 & ~n41646;
  assign n41648 = ~n41585 & ~n41647;
  assign n41649 = ~controllable_hgrant3 & ~n41648;
  assign n41650 = ~n12974 & ~n41649;
  assign n41651 = controllable_nhgrant0 & ~n41650;
  assign n41652 = ~n13845 & ~n41651;
  assign n41653 = ~n3281 & ~n41652;
  assign n41654 = ~n3281 & ~n41653;
  assign n41655 = n3378 & ~n41654;
  assign n41656 = ~n38371 & ~n41655;
  assign n41657 = n3492 & ~n41656;
  assign n41658 = ~n37174 & ~n41657;
  assign n41659 = n3485 & ~n41658;
  assign n41660 = ~n37332 & ~n41659;
  assign n41661 = n3476 & ~n41660;
  assign n41662 = ~n41529 & ~n41661;
  assign n41663 = n3374 & ~n41662;
  assign n41664 = ~n41522 & ~n41663;
  assign n41665 = n3655 & ~n41664;
  assign n41666 = n3378 & ~n40534;
  assign n41667 = ~n38413 & ~n41666;
  assign n41668 = n3492 & ~n41667;
  assign n41669 = n3492 & ~n41668;
  assign n41670 = n3485 & ~n41669;
  assign n41671 = n3485 & ~n41670;
  assign n41672 = ~n3476 & ~n41671;
  assign n41673 = ~n8523 & ~n41668;
  assign n41674 = n3485 & ~n41673;
  assign n41675 = ~n8689 & ~n41674;
  assign n41676 = n3476 & ~n41675;
  assign n41677 = ~n41672 & ~n41676;
  assign n41678 = ~n3374 & ~n41677;
  assign n41679 = n3378 & ~n40586;
  assign n41680 = ~n38485 & ~n41679;
  assign n41681 = n3492 & ~n41680;
  assign n41682 = n3492 & ~n41681;
  assign n41683 = n3485 & ~n41682;
  assign n41684 = n3485 & ~n41683;
  assign n41685 = ~n3476 & ~n41684;
  assign n41686 = ~n10404 & ~n41533;
  assign n41687 = ~controllable_hgrant2 & ~n41686;
  assign n41688 = ~n5616 & ~n41687;
  assign n41689 = controllable_hmaster1 & ~n41688;
  assign n41690 = controllable_hmaster0 & ~n41688;
  assign n41691 = ~n10483 & ~n41542;
  assign n41692 = ~controllable_hgrant2 & ~n41691;
  assign n41693 = ~n5616 & ~n41692;
  assign n41694 = ~controllable_hmaster0 & ~n41693;
  assign n41695 = ~n41690 & ~n41694;
  assign n41696 = ~controllable_hmaster1 & ~n41695;
  assign n41697 = ~n41689 & ~n41696;
  assign n41698 = i_hbusreq3 & ~n41697;
  assign n41699 = i_hbusreq2 & ~n41686;
  assign n41700 = ~n10443 & ~n41558;
  assign n41701 = ~i_hbusreq2 & ~n41700;
  assign n41702 = ~n41699 & ~n41701;
  assign n41703 = ~controllable_hgrant2 & ~n41702;
  assign n41704 = ~n5862 & ~n41703;
  assign n41705 = controllable_hmaster1 & ~n41704;
  assign n41706 = controllable_hmaster0 & ~n41704;
  assign n41707 = i_hbusreq2 & ~n41691;
  assign n41708 = ~n10521 & ~n41573;
  assign n41709 = ~i_hbusreq2 & ~n41708;
  assign n41710 = ~n41707 & ~n41709;
  assign n41711 = ~controllable_hgrant2 & ~n41710;
  assign n41712 = ~n5862 & ~n41711;
  assign n41713 = ~controllable_hmaster0 & ~n41712;
  assign n41714 = ~n41706 & ~n41713;
  assign n41715 = ~controllable_hmaster1 & ~n41714;
  assign n41716 = ~n41705 & ~n41715;
  assign n41717 = ~i_hbusreq3 & ~n41716;
  assign n41718 = ~n41698 & ~n41717;
  assign n41719 = controllable_hmaster2 & ~n41718;
  assign n41720 = ~n10483 & ~n41533;
  assign n41721 = ~controllable_hgrant2 & ~n41720;
  assign n41722 = ~n5686 & ~n41721;
  assign n41723 = ~controllable_hmaster0 & ~n41722;
  assign n41724 = ~n38585 & ~n41723;
  assign n41725 = controllable_hmaster1 & ~n41724;
  assign n41726 = ~n10498 & ~n41533;
  assign n41727 = ~controllable_hgrant2 & ~n41726;
  assign n41728 = ~n5616 & ~n41727;
  assign n41729 = controllable_hmaster0 & ~n41728;
  assign n41730 = ~n5616 & ~n41721;
  assign n41731 = ~controllable_hmaster0 & ~n41730;
  assign n41732 = ~n41729 & ~n41731;
  assign n41733 = ~controllable_hmaster1 & ~n41732;
  assign n41734 = ~n41725 & ~n41733;
  assign n41735 = i_hbusreq3 & ~n41734;
  assign n41736 = ~n10468 & ~n41607;
  assign n41737 = ~i_hbusreq2 & ~n41736;
  assign n41738 = ~n38590 & ~n41737;
  assign n41739 = ~controllable_hgrant2 & ~n41738;
  assign n41740 = ~n7507 & ~n41739;
  assign n41741 = controllable_hmaster0 & ~n41740;
  assign n41742 = i_hbusreq2 & ~n41720;
  assign n41743 = ~n10521 & ~n41558;
  assign n41744 = ~i_hbusreq2 & ~n41743;
  assign n41745 = ~n41742 & ~n41744;
  assign n41746 = ~controllable_hgrant2 & ~n41745;
  assign n41747 = ~n5950 & ~n41746;
  assign n41748 = ~controllable_hmaster0 & ~n41747;
  assign n41749 = ~n41741 & ~n41748;
  assign n41750 = controllable_hmaster1 & ~n41749;
  assign n41751 = i_hbusreq2 & ~n41726;
  assign n41752 = ~n10552 & ~n41558;
  assign n41753 = ~i_hbusreq2 & ~n41752;
  assign n41754 = ~n41751 & ~n41753;
  assign n41755 = ~controllable_hgrant2 & ~n41754;
  assign n41756 = ~n5862 & ~n41755;
  assign n41757 = controllable_hmaster0 & ~n41756;
  assign n41758 = ~n10567 & ~n41635;
  assign n41759 = ~i_hbusreq2 & ~n41758;
  assign n41760 = ~n41742 & ~n41759;
  assign n41761 = ~controllable_hgrant2 & ~n41760;
  assign n41762 = ~n5981 & ~n41761;
  assign n41763 = ~controllable_hmaster0 & ~n41762;
  assign n41764 = ~n41757 & ~n41763;
  assign n41765 = ~controllable_hmaster1 & ~n41764;
  assign n41766 = ~n41750 & ~n41765;
  assign n41767 = ~i_hbusreq3 & ~n41766;
  assign n41768 = ~n41735 & ~n41767;
  assign n41769 = ~controllable_hmaster2 & ~n41768;
  assign n41770 = ~n41719 & ~n41769;
  assign n41771 = ~controllable_hgrant3 & ~n41770;
  assign n41772 = ~n12974 & ~n41771;
  assign n41773 = controllable_nhgrant0 & ~n41772;
  assign n41774 = ~n13845 & ~n41773;
  assign n41775 = ~n3281 & ~n41774;
  assign n41776 = ~n3281 & ~n41775;
  assign n41777 = n3378 & ~n41776;
  assign n41778 = ~n38659 & ~n41777;
  assign n41779 = n3492 & ~n41778;
  assign n41780 = ~n37202 & ~n41779;
  assign n41781 = n3485 & ~n41780;
  assign n41782 = ~n37343 & ~n41781;
  assign n41783 = n3476 & ~n41782;
  assign n41784 = ~n41685 & ~n41783;
  assign n41785 = n3374 & ~n41784;
  assign n41786 = ~n41678 & ~n41785;
  assign n41787 = ~n3655 & ~n41786;
  assign n41788 = ~n41665 & ~n41787;
  assign n41789 = n3652 & ~n41788;
  assign n41790 = n3378 & ~n40748;
  assign n41791 = ~n38696 & ~n41790;
  assign n41792 = n3492 & ~n41791;
  assign n41793 = n3492 & ~n41792;
  assign n41794 = n3485 & ~n41793;
  assign n41795 = n3485 & ~n41794;
  assign n41796 = ~n3476 & ~n41795;
  assign n41797 = ~n8523 & ~n41792;
  assign n41798 = n3485 & ~n41797;
  assign n41799 = ~n8689 & ~n41798;
  assign n41800 = n3476 & ~n41799;
  assign n41801 = ~n41796 & ~n41800;
  assign n41802 = ~n3374 & ~n41801;
  assign n41803 = n3378 & ~n40800;
  assign n41804 = ~n38754 & ~n41803;
  assign n41805 = n3492 & ~n41804;
  assign n41806 = n3492 & ~n41805;
  assign n41807 = n3485 & ~n41806;
  assign n41808 = n3485 & ~n41807;
  assign n41809 = ~n3476 & ~n41808;
  assign n41810 = ~n10816 & ~n41535;
  assign n41811 = controllable_hmaster1 & ~n41810;
  assign n41812 = controllable_hmaster0 & ~n41810;
  assign n41813 = ~n10816 & ~n41544;
  assign n41814 = ~controllable_hmaster0 & ~n41813;
  assign n41815 = ~n41812 & ~n41814;
  assign n41816 = ~controllable_hmaster1 & ~n41815;
  assign n41817 = ~n41811 & ~n41816;
  assign n41818 = i_hbusreq3 & ~n41817;
  assign n41819 = ~n10870 & ~n41562;
  assign n41820 = controllable_hmaster1 & ~n41819;
  assign n41821 = controllable_hmaster0 & ~n41819;
  assign n41822 = ~n10870 & ~n41577;
  assign n41823 = ~controllable_hmaster0 & ~n41822;
  assign n41824 = ~n41821 & ~n41823;
  assign n41825 = ~controllable_hmaster1 & ~n41824;
  assign n41826 = ~n41820 & ~n41825;
  assign n41827 = ~i_hbusreq3 & ~n41826;
  assign n41828 = ~n41818 & ~n41827;
  assign n41829 = controllable_hmaster2 & ~n41828;
  assign n41830 = ~n10922 & ~n41587;
  assign n41831 = ~controllable_hmaster0 & ~n41830;
  assign n41832 = ~n38820 & ~n41831;
  assign n41833 = controllable_hmaster1 & ~n41832;
  assign n41834 = ~n10816 & ~n41593;
  assign n41835 = controllable_hmaster0 & ~n41834;
  assign n41836 = ~n10816 & ~n41587;
  assign n41837 = ~controllable_hmaster0 & ~n41836;
  assign n41838 = ~n41835 & ~n41837;
  assign n41839 = ~controllable_hmaster1 & ~n41838;
  assign n41840 = ~n41833 & ~n41839;
  assign n41841 = i_hbusreq3 & ~n41840;
  assign n41842 = ~n10904 & ~n41611;
  assign n41843 = controllable_hmaster0 & ~n41842;
  assign n41844 = ~n10972 & ~n41618;
  assign n41845 = ~controllable_hmaster0 & ~n41844;
  assign n41846 = ~n41843 & ~n41845;
  assign n41847 = controllable_hmaster1 & ~n41846;
  assign n41848 = ~n10870 & ~n41627;
  assign n41849 = controllable_hmaster0 & ~n41848;
  assign n41850 = ~n11002 & ~n41639;
  assign n41851 = ~controllable_hmaster0 & ~n41850;
  assign n41852 = ~n41849 & ~n41851;
  assign n41853 = ~controllable_hmaster1 & ~n41852;
  assign n41854 = ~n41847 & ~n41853;
  assign n41855 = ~i_hbusreq3 & ~n41854;
  assign n41856 = ~n41841 & ~n41855;
  assign n41857 = ~controllable_hmaster2 & ~n41856;
  assign n41858 = ~n41829 & ~n41857;
  assign n41859 = ~controllable_hgrant3 & ~n41858;
  assign n41860 = ~n12974 & ~n41859;
  assign n41861 = controllable_nhgrant0 & ~n41860;
  assign n41862 = ~n13845 & ~n41861;
  assign n41863 = ~n3281 & ~n41862;
  assign n41864 = ~n3281 & ~n41863;
  assign n41865 = n3378 & ~n41864;
  assign n41866 = ~n38870 & ~n41865;
  assign n41867 = n3492 & ~n41866;
  assign n41868 = ~n37231 & ~n41867;
  assign n41869 = n3485 & ~n41868;
  assign n41870 = ~n37356 & ~n41869;
  assign n41871 = n3476 & ~n41870;
  assign n41872 = ~n41809 & ~n41871;
  assign n41873 = n3374 & ~n41872;
  assign n41874 = ~n41802 & ~n41873;
  assign n41875 = n3655 & ~n41874;
  assign n41876 = n3378 & ~n40914;
  assign n41877 = ~n38905 & ~n41876;
  assign n41878 = n3492 & ~n41877;
  assign n41879 = n3492 & ~n41878;
  assign n41880 = n3485 & ~n41879;
  assign n41881 = n3485 & ~n41880;
  assign n41882 = ~n3476 & ~n41881;
  assign n41883 = ~n8523 & ~n41878;
  assign n41884 = n3485 & ~n41883;
  assign n41885 = ~n8689 & ~n41884;
  assign n41886 = n3476 & ~n41885;
  assign n41887 = ~n41882 & ~n41886;
  assign n41888 = ~n3374 & ~n41887;
  assign n41889 = n3378 & ~n40966;
  assign n41890 = ~n38963 & ~n41889;
  assign n41891 = n3492 & ~n41890;
  assign n41892 = n3492 & ~n41891;
  assign n41893 = n3485 & ~n41892;
  assign n41894 = n3485 & ~n41893;
  assign n41895 = ~n3476 & ~n41894;
  assign n41896 = ~n10816 & ~n41687;
  assign n41897 = controllable_hmaster1 & ~n41896;
  assign n41898 = controllable_hmaster0 & ~n41896;
  assign n41899 = ~n10816 & ~n41692;
  assign n41900 = ~controllable_hmaster0 & ~n41899;
  assign n41901 = ~n41898 & ~n41900;
  assign n41902 = ~controllable_hmaster1 & ~n41901;
  assign n41903 = ~n41897 & ~n41902;
  assign n41904 = i_hbusreq3 & ~n41903;
  assign n41905 = ~n10870 & ~n41703;
  assign n41906 = controllable_hmaster1 & ~n41905;
  assign n41907 = controllable_hmaster0 & ~n41905;
  assign n41908 = ~n10870 & ~n41711;
  assign n41909 = ~controllable_hmaster0 & ~n41908;
  assign n41910 = ~n41907 & ~n41909;
  assign n41911 = ~controllable_hmaster1 & ~n41910;
  assign n41912 = ~n41906 & ~n41911;
  assign n41913 = ~i_hbusreq3 & ~n41912;
  assign n41914 = ~n41904 & ~n41913;
  assign n41915 = controllable_hmaster2 & ~n41914;
  assign n41916 = ~n10922 & ~n41721;
  assign n41917 = ~controllable_hmaster0 & ~n41916;
  assign n41918 = ~n39029 & ~n41917;
  assign n41919 = controllable_hmaster1 & ~n41918;
  assign n41920 = ~n10816 & ~n41727;
  assign n41921 = controllable_hmaster0 & ~n41920;
  assign n41922 = ~n10816 & ~n41721;
  assign n41923 = ~controllable_hmaster0 & ~n41922;
  assign n41924 = ~n41921 & ~n41923;
  assign n41925 = ~controllable_hmaster1 & ~n41924;
  assign n41926 = ~n41919 & ~n41925;
  assign n41927 = i_hbusreq3 & ~n41926;
  assign n41928 = ~n10904 & ~n41739;
  assign n41929 = controllable_hmaster0 & ~n41928;
  assign n41930 = ~n10972 & ~n41746;
  assign n41931 = ~controllable_hmaster0 & ~n41930;
  assign n41932 = ~n41929 & ~n41931;
  assign n41933 = controllable_hmaster1 & ~n41932;
  assign n41934 = ~n10870 & ~n41755;
  assign n41935 = controllable_hmaster0 & ~n41934;
  assign n41936 = ~n11002 & ~n41761;
  assign n41937 = ~controllable_hmaster0 & ~n41936;
  assign n41938 = ~n41935 & ~n41937;
  assign n41939 = ~controllable_hmaster1 & ~n41938;
  assign n41940 = ~n41933 & ~n41939;
  assign n41941 = ~i_hbusreq3 & ~n41940;
  assign n41942 = ~n41927 & ~n41941;
  assign n41943 = ~controllable_hmaster2 & ~n41942;
  assign n41944 = ~n41915 & ~n41943;
  assign n41945 = ~controllable_hgrant3 & ~n41944;
  assign n41946 = ~n12974 & ~n41945;
  assign n41947 = controllable_nhgrant0 & ~n41946;
  assign n41948 = ~n13845 & ~n41947;
  assign n41949 = ~n3281 & ~n41948;
  assign n41950 = ~n3281 & ~n41949;
  assign n41951 = n3378 & ~n41950;
  assign n41952 = ~n39079 & ~n41951;
  assign n41953 = n3492 & ~n41952;
  assign n41954 = ~n37258 & ~n41953;
  assign n41955 = n3485 & ~n41954;
  assign n41956 = ~n37367 & ~n41955;
  assign n41957 = n3476 & ~n41956;
  assign n41958 = ~n41895 & ~n41957;
  assign n41959 = n3374 & ~n41958;
  assign n41960 = ~n41888 & ~n41959;
  assign n41961 = ~n3655 & ~n41960;
  assign n41962 = ~n41875 & ~n41961;
  assign n41963 = ~n3652 & ~n41962;
  assign n41964 = ~n41789 & ~n41963;
  assign n41965 = n3368 & ~n41964;
  assign n41966 = ~n41509 & ~n41965;
  assign n41967 = ~n3362 & ~n41966;
  assign n41968 = ~n41379 & ~n41967;
  assign n41969 = ~n3359 & ~n41968;
  assign n41970 = ~n41285 & ~n41969;
  assign n41971 = ~n3356 & ~n41970;
  assign n41972 = ~n39559 & ~n41971;
  assign n41973 = ~n3345 & ~n41972;
  assign n41974 = ~controllable_hmaster0 & ~n37423;
  assign n41975 = controllable_hmaster1 & ~n41974;
  assign n41976 = controllable_hmaster1 & ~n41975;
  assign n41977 = i_hbusreq3 & ~n41976;
  assign n41978 = ~controllable_hmaster0 & ~n37443;
  assign n41979 = controllable_hmaster1 & ~n41978;
  assign n41980 = controllable_hmaster1 & ~n41979;
  assign n41981 = ~i_hbusreq3 & ~n41980;
  assign n41982 = ~n41977 & ~n41981;
  assign n41983 = ~controllable_hmaster2 & ~n41982;
  assign n41984 = ~controllable_hmaster2 & ~n41983;
  assign n41985 = ~controllable_hgrant3 & ~n41984;
  assign n41986 = ~n14140 & ~n41985;
  assign n41987 = controllable_nhgrant0 & ~n41986;
  assign n41988 = ~n14166 & ~n41987;
  assign n41989 = ~n3281 & ~n41988;
  assign n41990 = ~n3281 & ~n41989;
  assign n41991 = n3378 & ~n41990;
  assign n41992 = ~n3530 & ~n41983;
  assign n41993 = ~controllable_hgrant3 & ~n41992;
  assign n41994 = ~n14172 & ~n41993;
  assign n41995 = controllable_nhgrant0 & ~n41994;
  assign n41996 = ~n14180 & ~n41995;
  assign n41997 = ~n3281 & ~n41996;
  assign n41998 = ~n3950 & ~n41997;
  assign n41999 = ~n3378 & ~n41998;
  assign n42000 = ~n41991 & ~n41999;
  assign n42001 = n3492 & ~n42000;
  assign n42002 = ~n3493 & ~n42001;
  assign n42003 = n3485 & ~n42002;
  assign n42004 = ~n3486 & ~n42003;
  assign n42005 = ~n3476 & ~n42004;
  assign n42006 = ~n5686 & ~n37419;
  assign n42007 = ~controllable_hmaster0 & ~n42006;
  assign n42008 = ~n14199 & ~n42007;
  assign n42009 = controllable_hmaster1 & ~n42008;
  assign n42010 = ~n14204 & ~n42009;
  assign n42011 = i_hbusreq3 & ~n42010;
  assign n42012 = ~n5950 & ~n37439;
  assign n42013 = ~controllable_hmaster0 & ~n42012;
  assign n42014 = ~n14207 & ~n42013;
  assign n42015 = controllable_hmaster1 & ~n42014;
  assign n42016 = ~n14212 & ~n42015;
  assign n42017 = ~i_hbusreq3 & ~n42016;
  assign n42018 = ~n42011 & ~n42017;
  assign n42019 = ~controllable_hmaster2 & ~n42018;
  assign n42020 = ~n14198 & ~n42019;
  assign n42021 = ~controllable_hgrant3 & ~n42020;
  assign n42022 = ~n14140 & ~n42021;
  assign n42023 = controllable_nhgrant0 & ~n42022;
  assign n42024 = ~n14166 & ~n42023;
  assign n42025 = ~n3281 & ~n42024;
  assign n42026 = ~n3281 & ~n42025;
  assign n42027 = n3378 & ~n42026;
  assign n42028 = ~n5686 & ~n39143;
  assign n42029 = ~controllable_hmaster0 & ~n42028;
  assign n42030 = ~n14246 & ~n42029;
  assign n42031 = controllable_hmaster1 & ~n42030;
  assign n42032 = ~n14251 & ~n42031;
  assign n42033 = i_hbusreq3 & ~n42032;
  assign n42034 = ~n5950 & ~n39154;
  assign n42035 = ~controllable_hmaster0 & ~n42034;
  assign n42036 = ~n14254 & ~n42035;
  assign n42037 = controllable_hmaster1 & ~n42036;
  assign n42038 = ~n14259 & ~n42037;
  assign n42039 = ~i_hbusreq3 & ~n42038;
  assign n42040 = ~n42033 & ~n42039;
  assign n42041 = ~controllable_hmaster2 & ~n42040;
  assign n42042 = ~n14245 & ~n42041;
  assign n42043 = ~controllable_hgrant3 & ~n42042;
  assign n42044 = ~n14172 & ~n42043;
  assign n42045 = controllable_nhgrant0 & ~n42044;
  assign n42046 = ~n14180 & ~n42045;
  assign n42047 = ~n3281 & ~n42046;
  assign n42048 = ~n4089 & ~n42047;
  assign n42049 = ~n3378 & ~n42048;
  assign n42050 = ~n42027 & ~n42049;
  assign n42051 = n3492 & ~n42050;
  assign n42052 = ~n3493 & ~n42051;
  assign n42053 = n3485 & ~n42052;
  assign n42054 = ~n3486 & ~n42053;
  assign n42055 = n3476 & ~n42054;
  assign n42056 = ~n42005 & ~n42055;
  assign n42057 = n3374 & ~n42056;
  assign n42058 = ~n14130 & ~n42057;
  assign n42059 = n3655 & ~n42058;
  assign n42060 = ~controllable_hmaster0 & ~n37617;
  assign n42061 = controllable_hmaster1 & ~n42060;
  assign n42062 = controllable_hmaster1 & ~n42061;
  assign n42063 = i_hbusreq3 & ~n42062;
  assign n42064 = ~controllable_hmaster0 & ~n37637;
  assign n42065 = controllable_hmaster1 & ~n42064;
  assign n42066 = controllable_hmaster1 & ~n42065;
  assign n42067 = ~i_hbusreq3 & ~n42066;
  assign n42068 = ~n42063 & ~n42067;
  assign n42069 = ~controllable_hmaster2 & ~n42068;
  assign n42070 = ~controllable_hmaster2 & ~n42069;
  assign n42071 = ~controllable_hgrant3 & ~n42070;
  assign n42072 = ~n14140 & ~n42071;
  assign n42073 = controllable_nhgrant0 & ~n42072;
  assign n42074 = ~n14166 & ~n42073;
  assign n42075 = ~n3281 & ~n42074;
  assign n42076 = ~n3281 & ~n42075;
  assign n42077 = n3378 & ~n42076;
  assign n42078 = ~n3530 & ~n42069;
  assign n42079 = ~controllable_hgrant3 & ~n42078;
  assign n42080 = ~n14172 & ~n42079;
  assign n42081 = controllable_nhgrant0 & ~n42080;
  assign n42082 = ~n14180 & ~n42081;
  assign n42083 = ~n3281 & ~n42082;
  assign n42084 = ~n3950 & ~n42083;
  assign n42085 = ~n3378 & ~n42084;
  assign n42086 = ~n42077 & ~n42085;
  assign n42087 = n3492 & ~n42086;
  assign n42088 = ~n3493 & ~n42087;
  assign n42089 = n3485 & ~n42088;
  assign n42090 = ~n3486 & ~n42089;
  assign n42091 = ~n3476 & ~n42090;
  assign n42092 = ~n5686 & ~n37613;
  assign n42093 = ~controllable_hmaster0 & ~n42092;
  assign n42094 = ~n14199 & ~n42093;
  assign n42095 = controllable_hmaster1 & ~n42094;
  assign n42096 = ~n14204 & ~n42095;
  assign n42097 = i_hbusreq3 & ~n42096;
  assign n42098 = ~n5950 & ~n37633;
  assign n42099 = ~controllable_hmaster0 & ~n42098;
  assign n42100 = ~n14207 & ~n42099;
  assign n42101 = controllable_hmaster1 & ~n42100;
  assign n42102 = ~n14212 & ~n42101;
  assign n42103 = ~i_hbusreq3 & ~n42102;
  assign n42104 = ~n42097 & ~n42103;
  assign n42105 = ~controllable_hmaster2 & ~n42104;
  assign n42106 = ~n14198 & ~n42105;
  assign n42107 = ~controllable_hgrant3 & ~n42106;
  assign n42108 = ~n14140 & ~n42107;
  assign n42109 = controllable_nhgrant0 & ~n42108;
  assign n42110 = ~n14166 & ~n42109;
  assign n42111 = ~n3281 & ~n42110;
  assign n42112 = ~n3281 & ~n42111;
  assign n42113 = n3378 & ~n42112;
  assign n42114 = ~n5686 & ~n39220;
  assign n42115 = ~controllable_hmaster0 & ~n42114;
  assign n42116 = ~n14246 & ~n42115;
  assign n42117 = controllable_hmaster1 & ~n42116;
  assign n42118 = ~n14251 & ~n42117;
  assign n42119 = i_hbusreq3 & ~n42118;
  assign n42120 = ~n5950 & ~n39231;
  assign n42121 = ~controllable_hmaster0 & ~n42120;
  assign n42122 = ~n14254 & ~n42121;
  assign n42123 = controllable_hmaster1 & ~n42122;
  assign n42124 = ~n14259 & ~n42123;
  assign n42125 = ~i_hbusreq3 & ~n42124;
  assign n42126 = ~n42119 & ~n42125;
  assign n42127 = ~controllable_hmaster2 & ~n42126;
  assign n42128 = ~n14245 & ~n42127;
  assign n42129 = ~controllable_hgrant3 & ~n42128;
  assign n42130 = ~n14172 & ~n42129;
  assign n42131 = controllable_nhgrant0 & ~n42130;
  assign n42132 = ~n14180 & ~n42131;
  assign n42133 = ~n3281 & ~n42132;
  assign n42134 = ~n4089 & ~n42133;
  assign n42135 = ~n3378 & ~n42134;
  assign n42136 = ~n42113 & ~n42135;
  assign n42137 = n3492 & ~n42136;
  assign n42138 = ~n3493 & ~n42137;
  assign n42139 = n3485 & ~n42138;
  assign n42140 = ~n3486 & ~n42139;
  assign n42141 = n3476 & ~n42140;
  assign n42142 = ~n42091 & ~n42141;
  assign n42143 = n3374 & ~n42142;
  assign n42144 = ~n14130 & ~n42143;
  assign n42145 = ~n3655 & ~n42144;
  assign n42146 = ~n42059 & ~n42145;
  assign n42147 = n3652 & ~n42146;
  assign n42148 = ~controllable_hmaster0 & ~n37818;
  assign n42149 = controllable_hmaster1 & ~n42148;
  assign n42150 = controllable_hmaster1 & ~n42149;
  assign n42151 = i_hbusreq3 & ~n42150;
  assign n42152 = ~controllable_hmaster0 & ~n37831;
  assign n42153 = controllable_hmaster1 & ~n42152;
  assign n42154 = controllable_hmaster1 & ~n42153;
  assign n42155 = ~i_hbusreq3 & ~n42154;
  assign n42156 = ~n42151 & ~n42155;
  assign n42157 = ~controllable_hmaster2 & ~n42156;
  assign n42158 = ~controllable_hmaster2 & ~n42157;
  assign n42159 = ~controllable_hgrant3 & ~n42158;
  assign n42160 = ~n14140 & ~n42159;
  assign n42161 = controllable_nhgrant0 & ~n42160;
  assign n42162 = ~n14166 & ~n42161;
  assign n42163 = ~n3281 & ~n42162;
  assign n42164 = ~n3281 & ~n42163;
  assign n42165 = n3378 & ~n42164;
  assign n42166 = ~n14470 & ~n42157;
  assign n42167 = ~controllable_hgrant3 & ~n42166;
  assign n42168 = ~n14172 & ~n42167;
  assign n42169 = controllable_nhgrant0 & ~n42168;
  assign n42170 = ~n14180 & ~n42169;
  assign n42171 = ~n3281 & ~n42170;
  assign n42172 = ~n3950 & ~n42171;
  assign n42173 = ~n3378 & ~n42172;
  assign n42174 = ~n42165 & ~n42173;
  assign n42175 = n3492 & ~n42174;
  assign n42176 = ~n3493 & ~n42175;
  assign n42177 = n3485 & ~n42176;
  assign n42178 = ~n3486 & ~n42177;
  assign n42179 = ~n3476 & ~n42178;
  assign n42180 = ~n6786 & ~n37419;
  assign n42181 = ~controllable_hmaster0 & ~n42180;
  assign n42182 = ~n14511 & ~n42181;
  assign n42183 = controllable_hmaster1 & ~n42182;
  assign n42184 = ~n14516 & ~n42183;
  assign n42185 = i_hbusreq3 & ~n42184;
  assign n42186 = ~n6813 & ~n37439;
  assign n42187 = ~controllable_hmaster0 & ~n42186;
  assign n42188 = ~n14519 & ~n42187;
  assign n42189 = controllable_hmaster1 & ~n42188;
  assign n42190 = ~n14524 & ~n42189;
  assign n42191 = ~i_hbusreq3 & ~n42190;
  assign n42192 = ~n42185 & ~n42191;
  assign n42193 = ~controllable_hmaster2 & ~n42192;
  assign n42194 = ~n14510 & ~n42193;
  assign n42195 = ~controllable_hgrant3 & ~n42194;
  assign n42196 = ~n14140 & ~n42195;
  assign n42197 = controllable_nhgrant0 & ~n42196;
  assign n42198 = ~n14166 & ~n42197;
  assign n42199 = ~n3281 & ~n42198;
  assign n42200 = ~n3281 & ~n42199;
  assign n42201 = n3378 & ~n42200;
  assign n42202 = ~n6786 & ~n39143;
  assign n42203 = ~controllable_hmaster0 & ~n42202;
  assign n42204 = ~n14571 & ~n42203;
  assign n42205 = controllable_hmaster1 & ~n42204;
  assign n42206 = ~n14576 & ~n42205;
  assign n42207 = i_hbusreq3 & ~n42206;
  assign n42208 = ~n6813 & ~n39154;
  assign n42209 = ~controllable_hmaster0 & ~n42208;
  assign n42210 = ~n14579 & ~n42209;
  assign n42211 = controllable_hmaster1 & ~n42210;
  assign n42212 = ~n14584 & ~n42211;
  assign n42213 = ~i_hbusreq3 & ~n42212;
  assign n42214 = ~n42207 & ~n42213;
  assign n42215 = ~controllable_hmaster2 & ~n42214;
  assign n42216 = ~n14570 & ~n42215;
  assign n42217 = ~controllable_hgrant3 & ~n42216;
  assign n42218 = ~n14172 & ~n42217;
  assign n42219 = controllable_nhgrant0 & ~n42218;
  assign n42220 = ~n14180 & ~n42219;
  assign n42221 = ~n3281 & ~n42220;
  assign n42222 = ~n4089 & ~n42221;
  assign n42223 = ~n3378 & ~n42222;
  assign n42224 = ~n42201 & ~n42223;
  assign n42225 = n3492 & ~n42224;
  assign n42226 = ~n14433 & ~n42225;
  assign n42227 = n3485 & ~n42226;
  assign n42228 = ~n14432 & ~n42227;
  assign n42229 = n3476 & ~n42228;
  assign n42230 = ~n42179 & ~n42229;
  assign n42231 = n3374 & ~n42230;
  assign n42232 = ~n14439 & ~n42231;
  assign n42233 = n3655 & ~n42232;
  assign n42234 = ~controllable_hmaster0 & ~n37972;
  assign n42235 = controllable_hmaster1 & ~n42234;
  assign n42236 = controllable_hmaster1 & ~n42235;
  assign n42237 = i_hbusreq3 & ~n42236;
  assign n42238 = ~controllable_hmaster0 & ~n37985;
  assign n42239 = controllable_hmaster1 & ~n42238;
  assign n42240 = controllable_hmaster1 & ~n42239;
  assign n42241 = ~i_hbusreq3 & ~n42240;
  assign n42242 = ~n42237 & ~n42241;
  assign n42243 = ~controllable_hmaster2 & ~n42242;
  assign n42244 = ~controllable_hmaster2 & ~n42243;
  assign n42245 = ~controllable_hgrant3 & ~n42244;
  assign n42246 = ~n14140 & ~n42245;
  assign n42247 = controllable_nhgrant0 & ~n42246;
  assign n42248 = ~n14166 & ~n42247;
  assign n42249 = ~n3281 & ~n42248;
  assign n42250 = ~n3281 & ~n42249;
  assign n42251 = n3378 & ~n42250;
  assign n42252 = ~n14470 & ~n42243;
  assign n42253 = ~controllable_hgrant3 & ~n42252;
  assign n42254 = ~n14172 & ~n42253;
  assign n42255 = controllable_nhgrant0 & ~n42254;
  assign n42256 = ~n14180 & ~n42255;
  assign n42257 = ~n3281 & ~n42256;
  assign n42258 = ~n3950 & ~n42257;
  assign n42259 = ~n3378 & ~n42258;
  assign n42260 = ~n42251 & ~n42259;
  assign n42261 = n3492 & ~n42260;
  assign n42262 = ~n3493 & ~n42261;
  assign n42263 = n3485 & ~n42262;
  assign n42264 = ~n3486 & ~n42263;
  assign n42265 = ~n3476 & ~n42264;
  assign n42266 = ~n6786 & ~n37613;
  assign n42267 = ~controllable_hmaster0 & ~n42266;
  assign n42268 = ~n14511 & ~n42267;
  assign n42269 = controllable_hmaster1 & ~n42268;
  assign n42270 = ~n14516 & ~n42269;
  assign n42271 = i_hbusreq3 & ~n42270;
  assign n42272 = ~n6813 & ~n37633;
  assign n42273 = ~controllable_hmaster0 & ~n42272;
  assign n42274 = ~n14519 & ~n42273;
  assign n42275 = controllable_hmaster1 & ~n42274;
  assign n42276 = ~n14524 & ~n42275;
  assign n42277 = ~i_hbusreq3 & ~n42276;
  assign n42278 = ~n42271 & ~n42277;
  assign n42279 = ~controllable_hmaster2 & ~n42278;
  assign n42280 = ~n14510 & ~n42279;
  assign n42281 = ~controllable_hgrant3 & ~n42280;
  assign n42282 = ~n14140 & ~n42281;
  assign n42283 = controllable_nhgrant0 & ~n42282;
  assign n42284 = ~n14166 & ~n42283;
  assign n42285 = ~n3281 & ~n42284;
  assign n42286 = ~n3281 & ~n42285;
  assign n42287 = n3378 & ~n42286;
  assign n42288 = ~n6786 & ~n39220;
  assign n42289 = ~controllable_hmaster0 & ~n42288;
  assign n42290 = ~n14571 & ~n42289;
  assign n42291 = controllable_hmaster1 & ~n42290;
  assign n42292 = ~n14576 & ~n42291;
  assign n42293 = i_hbusreq3 & ~n42292;
  assign n42294 = ~n6813 & ~n39231;
  assign n42295 = ~controllable_hmaster0 & ~n42294;
  assign n42296 = ~n14579 & ~n42295;
  assign n42297 = controllable_hmaster1 & ~n42296;
  assign n42298 = ~n14584 & ~n42297;
  assign n42299 = ~i_hbusreq3 & ~n42298;
  assign n42300 = ~n42293 & ~n42299;
  assign n42301 = ~controllable_hmaster2 & ~n42300;
  assign n42302 = ~n14570 & ~n42301;
  assign n42303 = ~controllable_hgrant3 & ~n42302;
  assign n42304 = ~n14172 & ~n42303;
  assign n42305 = controllable_nhgrant0 & ~n42304;
  assign n42306 = ~n14180 & ~n42305;
  assign n42307 = ~n3281 & ~n42306;
  assign n42308 = ~n4089 & ~n42307;
  assign n42309 = ~n3378 & ~n42308;
  assign n42310 = ~n42287 & ~n42309;
  assign n42311 = n3492 & ~n42310;
  assign n42312 = ~n14433 & ~n42311;
  assign n42313 = n3485 & ~n42312;
  assign n42314 = ~n14432 & ~n42313;
  assign n42315 = n3476 & ~n42314;
  assign n42316 = ~n42265 & ~n42315;
  assign n42317 = n3374 & ~n42316;
  assign n42318 = ~n14439 & ~n42317;
  assign n42319 = ~n3655 & ~n42318;
  assign n42320 = ~n42233 & ~n42319;
  assign n42321 = ~n3652 & ~n42320;
  assign n42322 = ~n42147 & ~n42321;
  assign n42323 = ~n3368 & ~n42322;
  assign n42324 = ~controllable_hmaster0 & ~n38143;
  assign n42325 = controllable_hmaster1 & ~n42324;
  assign n42326 = controllable_hmaster1 & ~n42325;
  assign n42327 = i_hbusreq3 & ~n42326;
  assign n42328 = ~controllable_hmaster0 & ~n38163;
  assign n42329 = controllable_hmaster1 & ~n42328;
  assign n42330 = controllable_hmaster1 & ~n42329;
  assign n42331 = ~i_hbusreq3 & ~n42330;
  assign n42332 = ~n42327 & ~n42331;
  assign n42333 = ~controllable_hmaster2 & ~n42332;
  assign n42334 = ~controllable_hmaster2 & ~n42333;
  assign n42335 = ~controllable_hgrant3 & ~n42334;
  assign n42336 = ~n14703 & ~n42335;
  assign n42337 = controllable_nhgrant0 & ~n42336;
  assign n42338 = ~n14725 & ~n42337;
  assign n42339 = ~n3281 & ~n42338;
  assign n42340 = ~n3281 & ~n42339;
  assign n42341 = n3492 & ~n42340;
  assign n42342 = n3492 & ~n42341;
  assign n42343 = n3485 & ~n42342;
  assign n42344 = n3485 & ~n42343;
  assign n42345 = ~n3476 & ~n42344;
  assign n42346 = ~n5686 & ~n38139;
  assign n42347 = ~controllable_hmaster0 & ~n42346;
  assign n42348 = ~n14199 & ~n42347;
  assign n42349 = controllable_hmaster1 & ~n42348;
  assign n42350 = ~n14204 & ~n42349;
  assign n42351 = i_hbusreq3 & ~n42350;
  assign n42352 = ~n10152 & ~n38159;
  assign n42353 = ~controllable_hmaster0 & ~n42352;
  assign n42354 = ~n14199 & ~n42353;
  assign n42355 = controllable_hmaster1 & ~n42354;
  assign n42356 = ~n14204 & ~n42355;
  assign n42357 = ~i_hbusreq3 & ~n42356;
  assign n42358 = ~n42351 & ~n42357;
  assign n42359 = ~controllable_hmaster2 & ~n42358;
  assign n42360 = ~n14734 & ~n42359;
  assign n42361 = ~controllable_hgrant3 & ~n42360;
  assign n42362 = ~n14703 & ~n42361;
  assign n42363 = controllable_nhgrant0 & ~n42362;
  assign n42364 = ~n14725 & ~n42363;
  assign n42365 = ~n3281 & ~n42364;
  assign n42366 = ~n3281 & ~n42365;
  assign n42367 = n3492 & ~n42366;
  assign n42368 = n3492 & ~n42367;
  assign n42369 = n3485 & ~n42368;
  assign n42370 = n3485 & ~n42369;
  assign n42371 = n3476 & ~n42370;
  assign n42372 = ~n42345 & ~n42371;
  assign n42373 = n3374 & ~n42372;
  assign n42374 = n3374 & ~n42373;
  assign n42375 = n3655 & ~n42374;
  assign n42376 = ~controllable_hmaster0 & ~n38442;
  assign n42377 = controllable_hmaster1 & ~n42376;
  assign n42378 = controllable_hmaster1 & ~n42377;
  assign n42379 = i_hbusreq3 & ~n42378;
  assign n42380 = ~controllable_hmaster0 & ~n38462;
  assign n42381 = controllable_hmaster1 & ~n42380;
  assign n42382 = controllable_hmaster1 & ~n42381;
  assign n42383 = ~i_hbusreq3 & ~n42382;
  assign n42384 = ~n42379 & ~n42383;
  assign n42385 = ~controllable_hmaster2 & ~n42384;
  assign n42386 = ~controllable_hmaster2 & ~n42385;
  assign n42387 = ~controllable_hgrant3 & ~n42386;
  assign n42388 = ~n14703 & ~n42387;
  assign n42389 = controllable_nhgrant0 & ~n42388;
  assign n42390 = ~n14725 & ~n42389;
  assign n42391 = ~n3281 & ~n42390;
  assign n42392 = ~n3281 & ~n42391;
  assign n42393 = n3492 & ~n42392;
  assign n42394 = n3492 & ~n42393;
  assign n42395 = n3485 & ~n42394;
  assign n42396 = n3485 & ~n42395;
  assign n42397 = ~n3476 & ~n42396;
  assign n42398 = ~n5686 & ~n38438;
  assign n42399 = ~controllable_hmaster0 & ~n42398;
  assign n42400 = ~n14199 & ~n42399;
  assign n42401 = controllable_hmaster1 & ~n42400;
  assign n42402 = ~n14204 & ~n42401;
  assign n42403 = i_hbusreq3 & ~n42402;
  assign n42404 = ~n10152 & ~n38458;
  assign n42405 = ~controllable_hmaster0 & ~n42404;
  assign n42406 = ~n14199 & ~n42405;
  assign n42407 = controllable_hmaster1 & ~n42406;
  assign n42408 = ~n14204 & ~n42407;
  assign n42409 = ~i_hbusreq3 & ~n42408;
  assign n42410 = ~n42403 & ~n42409;
  assign n42411 = ~controllable_hmaster2 & ~n42410;
  assign n42412 = ~n14734 & ~n42411;
  assign n42413 = ~controllable_hgrant3 & ~n42412;
  assign n42414 = ~n14703 & ~n42413;
  assign n42415 = controllable_nhgrant0 & ~n42414;
  assign n42416 = ~n14725 & ~n42415;
  assign n42417 = ~n3281 & ~n42416;
  assign n42418 = ~n3281 & ~n42417;
  assign n42419 = n3492 & ~n42418;
  assign n42420 = n3492 & ~n42419;
  assign n42421 = n3485 & ~n42420;
  assign n42422 = n3485 & ~n42421;
  assign n42423 = n3476 & ~n42422;
  assign n42424 = ~n42397 & ~n42423;
  assign n42425 = n3374 & ~n42424;
  assign n42426 = n3374 & ~n42425;
  assign n42427 = ~n3655 & ~n42426;
  assign n42428 = ~n42375 & ~n42427;
  assign n42429 = n3652 & ~n42428;
  assign n42430 = ~controllable_hmaster0 & ~n38723;
  assign n42431 = controllable_hmaster1 & ~n42430;
  assign n42432 = controllable_hmaster1 & ~n42431;
  assign n42433 = i_hbusreq3 & ~n42432;
  assign n42434 = ~controllable_hmaster0 & ~n38736;
  assign n42435 = controllable_hmaster1 & ~n42434;
  assign n42436 = controllable_hmaster1 & ~n42435;
  assign n42437 = ~i_hbusreq3 & ~n42436;
  assign n42438 = ~n42433 & ~n42437;
  assign n42439 = ~controllable_hmaster2 & ~n42438;
  assign n42440 = ~controllable_hmaster2 & ~n42439;
  assign n42441 = ~controllable_hgrant3 & ~n42440;
  assign n42442 = ~n14703 & ~n42441;
  assign n42443 = controllable_nhgrant0 & ~n42442;
  assign n42444 = ~n14725 & ~n42443;
  assign n42445 = ~n3281 & ~n42444;
  assign n42446 = ~n3281 & ~n42445;
  assign n42447 = n3492 & ~n42446;
  assign n42448 = n3492 & ~n42447;
  assign n42449 = n3485 & ~n42448;
  assign n42450 = n3485 & ~n42449;
  assign n42451 = ~n3476 & ~n42450;
  assign n42452 = ~n11066 & ~n38139;
  assign n42453 = ~controllable_hmaster0 & ~n42452;
  assign n42454 = ~n14863 & ~n42453;
  assign n42455 = controllable_hmaster1 & ~n42454;
  assign n42456 = ~n14868 & ~n42455;
  assign n42457 = i_hbusreq3 & ~n42456;
  assign n42458 = ~n11110 & ~n38159;
  assign n42459 = ~controllable_hmaster0 & ~n42458;
  assign n42460 = ~n14871 & ~n42459;
  assign n42461 = controllable_hmaster1 & ~n42460;
  assign n42462 = ~n14876 & ~n42461;
  assign n42463 = ~i_hbusreq3 & ~n42462;
  assign n42464 = ~n42457 & ~n42463;
  assign n42465 = ~controllable_hmaster2 & ~n42464;
  assign n42466 = ~n14862 & ~n42465;
  assign n42467 = ~controllable_hgrant3 & ~n42466;
  assign n42468 = ~n14703 & ~n42467;
  assign n42469 = controllable_nhgrant0 & ~n42468;
  assign n42470 = ~n14725 & ~n42469;
  assign n42471 = ~n3281 & ~n42470;
  assign n42472 = ~n3281 & ~n42471;
  assign n42473 = n3492 & ~n42472;
  assign n42474 = ~n14836 & ~n42473;
  assign n42475 = n3485 & ~n42474;
  assign n42476 = ~n14835 & ~n42475;
  assign n42477 = n3476 & ~n42476;
  assign n42478 = ~n42451 & ~n42477;
  assign n42479 = n3374 & ~n42478;
  assign n42480 = n3374 & ~n42479;
  assign n42481 = n3655 & ~n42480;
  assign n42482 = ~controllable_hmaster0 & ~n38932;
  assign n42483 = controllable_hmaster1 & ~n42482;
  assign n42484 = controllable_hmaster1 & ~n42483;
  assign n42485 = i_hbusreq3 & ~n42484;
  assign n42486 = ~controllable_hmaster0 & ~n38945;
  assign n42487 = controllable_hmaster1 & ~n42486;
  assign n42488 = controllable_hmaster1 & ~n42487;
  assign n42489 = ~i_hbusreq3 & ~n42488;
  assign n42490 = ~n42485 & ~n42489;
  assign n42491 = ~controllable_hmaster2 & ~n42490;
  assign n42492 = ~controllable_hmaster2 & ~n42491;
  assign n42493 = ~controllable_hgrant3 & ~n42492;
  assign n42494 = ~n14703 & ~n42493;
  assign n42495 = controllable_nhgrant0 & ~n42494;
  assign n42496 = ~n14725 & ~n42495;
  assign n42497 = ~n3281 & ~n42496;
  assign n42498 = ~n3281 & ~n42497;
  assign n42499 = n3492 & ~n42498;
  assign n42500 = n3492 & ~n42499;
  assign n42501 = n3485 & ~n42500;
  assign n42502 = n3485 & ~n42501;
  assign n42503 = ~n3476 & ~n42502;
  assign n42504 = ~n11066 & ~n38438;
  assign n42505 = ~controllable_hmaster0 & ~n42504;
  assign n42506 = ~n14863 & ~n42505;
  assign n42507 = controllable_hmaster1 & ~n42506;
  assign n42508 = ~n14868 & ~n42507;
  assign n42509 = i_hbusreq3 & ~n42508;
  assign n42510 = ~n11110 & ~n38458;
  assign n42511 = ~controllable_hmaster0 & ~n42510;
  assign n42512 = ~n14871 & ~n42511;
  assign n42513 = controllable_hmaster1 & ~n42512;
  assign n42514 = ~n14876 & ~n42513;
  assign n42515 = ~i_hbusreq3 & ~n42514;
  assign n42516 = ~n42509 & ~n42515;
  assign n42517 = ~controllable_hmaster2 & ~n42516;
  assign n42518 = ~n14862 & ~n42517;
  assign n42519 = ~controllable_hgrant3 & ~n42518;
  assign n42520 = ~n14703 & ~n42519;
  assign n42521 = controllable_nhgrant0 & ~n42520;
  assign n42522 = ~n14725 & ~n42521;
  assign n42523 = ~n3281 & ~n42522;
  assign n42524 = ~n3281 & ~n42523;
  assign n42525 = n3492 & ~n42524;
  assign n42526 = ~n14836 & ~n42525;
  assign n42527 = n3485 & ~n42526;
  assign n42528 = ~n14835 & ~n42527;
  assign n42529 = n3476 & ~n42528;
  assign n42530 = ~n42503 & ~n42529;
  assign n42531 = n3374 & ~n42530;
  assign n42532 = n3374 & ~n42531;
  assign n42533 = ~n3655 & ~n42532;
  assign n42534 = ~n42481 & ~n42533;
  assign n42535 = ~n3652 & ~n42534;
  assign n42536 = ~n42429 & ~n42535;
  assign n42537 = n3368 & ~n42536;
  assign n42538 = ~n42323 & ~n42537;
  assign n42539 = ~n3362 & ~n42538;
  assign n42540 = ~n3362 & ~n42539;
  assign n42541 = ~n3359 & ~n42540;
  assign n42542 = ~n3359 & ~n42541;
  assign n42543 = n3356 & ~n42542;
  assign n42544 = ~n14959 & ~n39590;
  assign n42545 = n3492 & ~n42544;
  assign n42546 = ~n3631 & ~n42545;
  assign n42547 = n3485 & ~n42546;
  assign n42548 = ~n3630 & ~n42547;
  assign n42549 = ~n3374 & ~n42548;
  assign n42550 = ~n3382 & ~n37423;
  assign n42551 = controllable_hmaster1 & ~n42550;
  assign n42552 = ~n5305 & ~n42551;
  assign n42553 = i_hbusreq3 & ~n42552;
  assign n42554 = ~n3401 & ~n37443;
  assign n42555 = controllable_hmaster1 & ~n42554;
  assign n42556 = ~n5334 & ~n42555;
  assign n42557 = ~i_hbusreq3 & ~n42556;
  assign n42558 = ~n42553 & ~n42557;
  assign n42559 = ~controllable_hmaster2 & ~n42558;
  assign n42560 = ~n12065 & ~n42559;
  assign n42561 = ~controllable_hgrant3 & ~n42560;
  assign n42562 = ~n14973 & ~n42561;
  assign n42563 = controllable_nhgrant0 & ~n42562;
  assign n42564 = ~n15006 & ~n42563;
  assign n42565 = ~n3281 & ~n42564;
  assign n42566 = ~n3950 & ~n42565;
  assign n42567 = n3378 & ~n42566;
  assign n42568 = ~n35053 & ~n37423;
  assign n42569 = controllable_hmaster1 & ~n42568;
  assign n42570 = ~n35064 & ~n42569;
  assign n42571 = i_hbusreq3 & ~n42570;
  assign n42572 = ~n35072 & ~n37443;
  assign n42573 = controllable_hmaster1 & ~n42572;
  assign n42574 = ~n35091 & ~n42573;
  assign n42575 = ~i_hbusreq3 & ~n42574;
  assign n42576 = ~n42571 & ~n42575;
  assign n42577 = ~controllable_hmaster2 & ~n42576;
  assign n42578 = ~n39648 & ~n42577;
  assign n42579 = ~controllable_hgrant3 & ~n42578;
  assign n42580 = ~n5402 & ~n42579;
  assign n42581 = controllable_nhgrant0 & ~n42580;
  assign n42582 = ~n5534 & ~n42581;
  assign n42583 = ~n3281 & ~n42582;
  assign n42584 = ~n3950 & ~n42583;
  assign n42585 = ~n3378 & ~n42584;
  assign n42586 = ~n42567 & ~n42585;
  assign n42587 = n3492 & ~n42586;
  assign n42588 = ~n3631 & ~n42587;
  assign n42589 = n3485 & ~n42588;
  assign n42590 = ~n3630 & ~n42589;
  assign n42591 = ~n3476 & ~n42590;
  assign n42592 = ~n5686 & ~n39675;
  assign n42593 = ~controllable_hmaster0 & ~n42592;
  assign n42594 = ~n5685 & ~n42593;
  assign n42595 = controllable_hmaster1 & ~n42594;
  assign n42596 = ~n5704 & ~n42595;
  assign n42597 = i_hbusreq3 & ~n42596;
  assign n42598 = ~n5950 & ~n39687;
  assign n42599 = ~controllable_hmaster0 & ~n42598;
  assign n42600 = ~n15059 & ~n42599;
  assign n42601 = controllable_hmaster1 & ~n42600;
  assign n42602 = ~n15068 & ~n42601;
  assign n42603 = ~i_hbusreq3 & ~n42602;
  assign n42604 = ~n42597 & ~n42603;
  assign n42605 = ~controllable_hmaster2 & ~n42604;
  assign n42606 = ~n15053 & ~n42605;
  assign n42607 = ~controllable_hgrant3 & ~n42606;
  assign n42608 = ~n15042 & ~n42607;
  assign n42609 = controllable_nhgrant0 & ~n42608;
  assign n42610 = ~n15088 & ~n42609;
  assign n42611 = ~n3281 & ~n42610;
  assign n42612 = ~n4089 & ~n42611;
  assign n42613 = n3378 & ~n42612;
  assign n42614 = ~n35219 & ~n37505;
  assign n42615 = controllable_hmaster1 & ~n42614;
  assign n42616 = ~n35230 & ~n42615;
  assign n42617 = i_hbusreq3 & ~n42616;
  assign n42618 = ~n5950 & ~n39740;
  assign n42619 = ~controllable_hmaster0 & ~n42618;
  assign n42620 = ~n35240 & ~n42619;
  assign n42621 = controllable_hmaster1 & ~n42620;
  assign n42622 = ~n35260 & ~n42621;
  assign n42623 = ~i_hbusreq3 & ~n42622;
  assign n42624 = ~n42617 & ~n42623;
  assign n42625 = ~controllable_hmaster2 & ~n42624;
  assign n42626 = ~n39732 & ~n42625;
  assign n42627 = ~controllable_hgrant3 & ~n42626;
  assign n42628 = ~n5861 & ~n42627;
  assign n42629 = controllable_nhgrant0 & ~n42628;
  assign n42630 = ~n6082 & ~n42629;
  assign n42631 = ~n3281 & ~n42630;
  assign n42632 = ~n4089 & ~n42631;
  assign n42633 = ~n3378 & ~n42632;
  assign n42634 = ~n42613 & ~n42633;
  assign n42635 = n3492 & ~n42634;
  assign n42636 = ~n3631 & ~n42635;
  assign n42637 = n3485 & ~n42636;
  assign n42638 = ~n3630 & ~n42637;
  assign n42639 = n3476 & ~n42638;
  assign n42640 = ~n42591 & ~n42639;
  assign n42641 = n3374 & ~n42640;
  assign n42642 = ~n42549 & ~n42641;
  assign n42643 = n3655 & ~n42642;
  assign n42644 = ~n14959 & ~n39797;
  assign n42645 = n3492 & ~n42644;
  assign n42646 = ~n3631 & ~n42645;
  assign n42647 = n3485 & ~n42646;
  assign n42648 = ~n3630 & ~n42647;
  assign n42649 = ~n3374 & ~n42648;
  assign n42650 = ~n3382 & ~n37617;
  assign n42651 = controllable_hmaster1 & ~n42650;
  assign n42652 = ~n5305 & ~n42651;
  assign n42653 = i_hbusreq3 & ~n42652;
  assign n42654 = ~n3401 & ~n37637;
  assign n42655 = controllable_hmaster1 & ~n42654;
  assign n42656 = ~n5334 & ~n42655;
  assign n42657 = ~i_hbusreq3 & ~n42656;
  assign n42658 = ~n42653 & ~n42657;
  assign n42659 = ~controllable_hmaster2 & ~n42658;
  assign n42660 = ~n12065 & ~n42659;
  assign n42661 = ~controllable_hgrant3 & ~n42660;
  assign n42662 = ~n14973 & ~n42661;
  assign n42663 = controllable_nhgrant0 & ~n42662;
  assign n42664 = ~n15006 & ~n42663;
  assign n42665 = ~n3281 & ~n42664;
  assign n42666 = ~n3950 & ~n42665;
  assign n42667 = n3378 & ~n42666;
  assign n42668 = ~n35360 & ~n37617;
  assign n42669 = controllable_hmaster1 & ~n42668;
  assign n42670 = ~n35371 & ~n42669;
  assign n42671 = i_hbusreq3 & ~n42670;
  assign n42672 = ~n35380 & ~n37637;
  assign n42673 = controllable_hmaster1 & ~n42672;
  assign n42674 = ~n35400 & ~n42673;
  assign n42675 = ~i_hbusreq3 & ~n42674;
  assign n42676 = ~n42671 & ~n42675;
  assign n42677 = ~controllable_hmaster2 & ~n42676;
  assign n42678 = ~n39855 & ~n42677;
  assign n42679 = ~controllable_hgrant3 & ~n42678;
  assign n42680 = ~n5402 & ~n42679;
  assign n42681 = controllable_nhgrant0 & ~n42680;
  assign n42682 = ~n5534 & ~n42681;
  assign n42683 = ~n3281 & ~n42682;
  assign n42684 = ~n3950 & ~n42683;
  assign n42685 = ~n3378 & ~n42684;
  assign n42686 = ~n42667 & ~n42685;
  assign n42687 = n3492 & ~n42686;
  assign n42688 = ~n3631 & ~n42687;
  assign n42689 = n3485 & ~n42688;
  assign n42690 = ~n3630 & ~n42689;
  assign n42691 = ~n3476 & ~n42690;
  assign n42692 = ~n5686 & ~n39881;
  assign n42693 = ~controllable_hmaster0 & ~n42692;
  assign n42694 = ~n5685 & ~n42693;
  assign n42695 = controllable_hmaster1 & ~n42694;
  assign n42696 = ~n5704 & ~n42695;
  assign n42697 = i_hbusreq3 & ~n42696;
  assign n42698 = ~n5950 & ~n39892;
  assign n42699 = ~controllable_hmaster0 & ~n42698;
  assign n42700 = ~n15059 & ~n42699;
  assign n42701 = controllable_hmaster1 & ~n42700;
  assign n42702 = ~n15068 & ~n42701;
  assign n42703 = ~i_hbusreq3 & ~n42702;
  assign n42704 = ~n42697 & ~n42703;
  assign n42705 = ~controllable_hmaster2 & ~n42704;
  assign n42706 = ~n15053 & ~n42705;
  assign n42707 = ~controllable_hgrant3 & ~n42706;
  assign n42708 = ~n15042 & ~n42707;
  assign n42709 = controllable_nhgrant0 & ~n42708;
  assign n42710 = ~n15088 & ~n42709;
  assign n42711 = ~n3281 & ~n42710;
  assign n42712 = ~n4089 & ~n42711;
  assign n42713 = n3378 & ~n42712;
  assign n42714 = ~n35485 & ~n37708;
  assign n42715 = controllable_hmaster1 & ~n42714;
  assign n42716 = ~n35496 & ~n42715;
  assign n42717 = i_hbusreq3 & ~n42716;
  assign n42718 = ~n5950 & ~n39945;
  assign n42719 = ~controllable_hmaster0 & ~n42718;
  assign n42720 = ~n35505 & ~n42719;
  assign n42721 = controllable_hmaster1 & ~n42720;
  assign n42722 = ~n35524 & ~n42721;
  assign n42723 = ~i_hbusreq3 & ~n42722;
  assign n42724 = ~n42717 & ~n42723;
  assign n42725 = ~controllable_hmaster2 & ~n42724;
  assign n42726 = ~n39937 & ~n42725;
  assign n42727 = ~controllable_hgrant3 & ~n42726;
  assign n42728 = ~n5861 & ~n42727;
  assign n42729 = controllable_nhgrant0 & ~n42728;
  assign n42730 = ~n6082 & ~n42729;
  assign n42731 = ~n3281 & ~n42730;
  assign n42732 = ~n4089 & ~n42731;
  assign n42733 = ~n3378 & ~n42732;
  assign n42734 = ~n42713 & ~n42733;
  assign n42735 = n3492 & ~n42734;
  assign n42736 = ~n3631 & ~n42735;
  assign n42737 = n3485 & ~n42736;
  assign n42738 = ~n3630 & ~n42737;
  assign n42739 = n3476 & ~n42738;
  assign n42740 = ~n42691 & ~n42739;
  assign n42741 = n3374 & ~n42740;
  assign n42742 = ~n42649 & ~n42741;
  assign n42743 = ~n3655 & ~n42742;
  assign n42744 = ~n42643 & ~n42743;
  assign n42745 = n3652 & ~n42744;
  assign n42746 = ~n9388 & ~n39561;
  assign n42747 = controllable_hmaster1 & ~n42746;
  assign n42748 = controllable_hmaster0 & ~n42746;
  assign n42749 = ~n34022 & ~n42748;
  assign n42750 = ~controllable_hmaster1 & ~n42749;
  assign n42751 = ~n42747 & ~n42750;
  assign n42752 = i_hbusreq3 & ~n42751;
  assign n42753 = ~n15233 & ~n39573;
  assign n42754 = controllable_hmaster1 & ~n42753;
  assign n42755 = controllable_hmaster0 & ~n42753;
  assign n42756 = ~n34040 & ~n42755;
  assign n42757 = ~controllable_hmaster1 & ~n42756;
  assign n42758 = ~n42754 & ~n42757;
  assign n42759 = ~i_hbusreq3 & ~n42758;
  assign n42760 = ~n42752 & ~n42759;
  assign n42761 = controllable_hmaster2 & ~n42760;
  assign n42762 = ~n6657 & ~n42761;
  assign n42763 = ~controllable_hgrant3 & ~n42762;
  assign n42764 = ~n5037 & ~n42763;
  assign n42765 = controllable_nhgrant0 & ~n42764;
  assign n42766 = ~n5245 & ~n42765;
  assign n42767 = ~n3281 & ~n42766;
  assign n42768 = ~n3783 & ~n42767;
  assign n42769 = ~n3378 & ~n42768;
  assign n42770 = ~n15225 & ~n42769;
  assign n42771 = n3492 & ~n42770;
  assign n42772 = ~n3631 & ~n42771;
  assign n42773 = n3485 & ~n42772;
  assign n42774 = ~n3630 & ~n42773;
  assign n42775 = ~n3476 & ~n42774;
  assign n42776 = ~n15258 & ~n42771;
  assign n42777 = n3485 & ~n42776;
  assign n42778 = ~n15257 & ~n42777;
  assign n42779 = n3476 & ~n42778;
  assign n42780 = ~n42775 & ~n42779;
  assign n42781 = ~n3374 & ~n42780;
  assign n42782 = ~n15289 & ~n37818;
  assign n42783 = controllable_hmaster1 & ~n42782;
  assign n42784 = ~n15296 & ~n42783;
  assign n42785 = i_hbusreq3 & ~n42784;
  assign n42786 = ~n15300 & ~n37831;
  assign n42787 = controllable_hmaster1 & ~n42786;
  assign n42788 = ~n15307 & ~n42787;
  assign n42789 = ~i_hbusreq3 & ~n42788;
  assign n42790 = ~n42785 & ~n42789;
  assign n42791 = ~controllable_hmaster2 & ~n42790;
  assign n42792 = ~n15287 & ~n42791;
  assign n42793 = ~controllable_hgrant3 & ~n42792;
  assign n42794 = ~n14973 & ~n42793;
  assign n42795 = controllable_nhgrant0 & ~n42794;
  assign n42796 = ~n15006 & ~n42795;
  assign n42797 = ~n3281 & ~n42796;
  assign n42798 = ~n3950 & ~n42797;
  assign n42799 = n3378 & ~n42798;
  assign n42800 = ~n9388 & ~n39616;
  assign n42801 = controllable_hmaster1 & ~n42800;
  assign n42802 = controllable_hmaster0 & ~n42800;
  assign n42803 = ~n40026 & ~n42802;
  assign n42804 = ~controllable_hmaster1 & ~n42803;
  assign n42805 = ~n42801 & ~n42804;
  assign n42806 = i_hbusreq3 & ~n42805;
  assign n42807 = ~n15233 & ~n39632;
  assign n42808 = controllable_hmaster1 & ~n42807;
  assign n42809 = controllable_hmaster0 & ~n42807;
  assign n42810 = ~n40035 & ~n42809;
  assign n42811 = ~controllable_hmaster1 & ~n42810;
  assign n42812 = ~n42808 & ~n42811;
  assign n42813 = ~i_hbusreq3 & ~n42812;
  assign n42814 = ~n42806 & ~n42813;
  assign n42815 = controllable_hmaster2 & ~n42814;
  assign n42816 = ~n35610 & ~n37818;
  assign n42817 = controllable_hmaster1 & ~n42816;
  assign n42818 = ~n35619 & ~n42817;
  assign n42819 = i_hbusreq3 & ~n42818;
  assign n42820 = ~n35623 & ~n37831;
  assign n42821 = controllable_hmaster1 & ~n42820;
  assign n42822 = ~n35633 & ~n42821;
  assign n42823 = ~i_hbusreq3 & ~n42822;
  assign n42824 = ~n42819 & ~n42823;
  assign n42825 = ~controllable_hmaster2 & ~n42824;
  assign n42826 = ~n42815 & ~n42825;
  assign n42827 = ~controllable_hgrant3 & ~n42826;
  assign n42828 = ~n5402 & ~n42827;
  assign n42829 = controllable_nhgrant0 & ~n42828;
  assign n42830 = ~n5534 & ~n42829;
  assign n42831 = ~n3281 & ~n42830;
  assign n42832 = ~n3950 & ~n42831;
  assign n42833 = ~n3378 & ~n42832;
  assign n42834 = ~n42799 & ~n42833;
  assign n42835 = n3492 & ~n42834;
  assign n42836 = ~n3631 & ~n42835;
  assign n42837 = n3485 & ~n42836;
  assign n42838 = ~n3630 & ~n42837;
  assign n42839 = ~n3476 & ~n42838;
  assign n42840 = ~n6786 & ~n39675;
  assign n42841 = ~controllable_hmaster0 & ~n42840;
  assign n42842 = ~n15387 & ~n42841;
  assign n42843 = controllable_hmaster1 & ~n42842;
  assign n42844 = ~n15394 & ~n42843;
  assign n42845 = i_hbusreq3 & ~n42844;
  assign n42846 = ~n6813 & ~n39687;
  assign n42847 = ~controllable_hmaster0 & ~n42846;
  assign n42848 = ~n15398 & ~n42847;
  assign n42849 = controllable_hmaster1 & ~n42848;
  assign n42850 = ~n15407 & ~n42849;
  assign n42851 = ~i_hbusreq3 & ~n42850;
  assign n42852 = ~n42845 & ~n42851;
  assign n42853 = ~controllable_hmaster2 & ~n42852;
  assign n42854 = ~n15385 & ~n42853;
  assign n42855 = ~controllable_hgrant3 & ~n42854;
  assign n42856 = ~n15042 & ~n42855;
  assign n42857 = controllable_nhgrant0 & ~n42856;
  assign n42858 = ~n15088 & ~n42857;
  assign n42859 = ~n3281 & ~n42858;
  assign n42860 = ~n4089 & ~n42859;
  assign n42861 = n3378 & ~n42860;
  assign n42862 = ~n9477 & ~n37501;
  assign n42863 = controllable_hmaster1 & ~n42862;
  assign n42864 = controllable_hmaster0 & ~n42862;
  assign n42865 = ~n40090 & ~n42864;
  assign n42866 = ~controllable_hmaster1 & ~n42865;
  assign n42867 = ~n42863 & ~n42866;
  assign n42868 = i_hbusreq3 & ~n42867;
  assign n42869 = ~n15433 & ~n39716;
  assign n42870 = controllable_hmaster1 & ~n42869;
  assign n42871 = controllable_hmaster0 & ~n42869;
  assign n42872 = ~n40099 & ~n42871;
  assign n42873 = ~controllable_hmaster1 & ~n42872;
  assign n42874 = ~n42870 & ~n42873;
  assign n42875 = ~i_hbusreq3 & ~n42874;
  assign n42876 = ~n42868 & ~n42875;
  assign n42877 = controllable_hmaster2 & ~n42876;
  assign n42878 = ~n35695 & ~n37880;
  assign n42879 = controllable_hmaster1 & ~n42878;
  assign n42880 = ~n35704 & ~n42879;
  assign n42881 = i_hbusreq3 & ~n42880;
  assign n42882 = ~n6813 & ~n39740;
  assign n42883 = ~controllable_hmaster0 & ~n42882;
  assign n42884 = ~n35708 & ~n42883;
  assign n42885 = controllable_hmaster1 & ~n42884;
  assign n42886 = ~n35718 & ~n42885;
  assign n42887 = ~i_hbusreq3 & ~n42886;
  assign n42888 = ~n42881 & ~n42887;
  assign n42889 = ~controllable_hmaster2 & ~n42888;
  assign n42890 = ~n42877 & ~n42889;
  assign n42891 = ~controllable_hgrant3 & ~n42890;
  assign n42892 = ~n5861 & ~n42891;
  assign n42893 = controllable_nhgrant0 & ~n42892;
  assign n42894 = ~n6082 & ~n42893;
  assign n42895 = ~n3281 & ~n42894;
  assign n42896 = ~n4089 & ~n42895;
  assign n42897 = ~n3378 & ~n42896;
  assign n42898 = ~n42861 & ~n42897;
  assign n42899 = n3492 & ~n42898;
  assign n42900 = ~n15258 & ~n42899;
  assign n42901 = n3485 & ~n42900;
  assign n42902 = ~n15257 & ~n42901;
  assign n42903 = n3476 & ~n42902;
  assign n42904 = ~n42839 & ~n42903;
  assign n42905 = n3374 & ~n42904;
  assign n42906 = ~n42781 & ~n42905;
  assign n42907 = n3655 & ~n42906;
  assign n42908 = ~n9388 & ~n39768;
  assign n42909 = controllable_hmaster1 & ~n42908;
  assign n42910 = controllable_hmaster0 & ~n42908;
  assign n42911 = ~n34022 & ~n42910;
  assign n42912 = ~controllable_hmaster1 & ~n42911;
  assign n42913 = ~n42909 & ~n42912;
  assign n42914 = i_hbusreq3 & ~n42913;
  assign n42915 = ~n15233 & ~n39780;
  assign n42916 = controllable_hmaster1 & ~n42915;
  assign n42917 = controllable_hmaster0 & ~n42915;
  assign n42918 = ~n34040 & ~n42917;
  assign n42919 = ~controllable_hmaster1 & ~n42918;
  assign n42920 = ~n42916 & ~n42919;
  assign n42921 = ~i_hbusreq3 & ~n42920;
  assign n42922 = ~n42914 & ~n42921;
  assign n42923 = controllable_hmaster2 & ~n42922;
  assign n42924 = ~n6887 & ~n42923;
  assign n42925 = ~controllable_hgrant3 & ~n42924;
  assign n42926 = ~n5037 & ~n42925;
  assign n42927 = controllable_nhgrant0 & ~n42926;
  assign n42928 = ~n5245 & ~n42927;
  assign n42929 = ~n3281 & ~n42928;
  assign n42930 = ~n3783 & ~n42929;
  assign n42931 = ~n3378 & ~n42930;
  assign n42932 = ~n15225 & ~n42931;
  assign n42933 = n3492 & ~n42932;
  assign n42934 = ~n3631 & ~n42933;
  assign n42935 = n3485 & ~n42934;
  assign n42936 = ~n3630 & ~n42935;
  assign n42937 = ~n3476 & ~n42936;
  assign n42938 = ~n15258 & ~n42933;
  assign n42939 = n3485 & ~n42938;
  assign n42940 = ~n15257 & ~n42939;
  assign n42941 = n3476 & ~n42940;
  assign n42942 = ~n42937 & ~n42941;
  assign n42943 = ~n3374 & ~n42942;
  assign n42944 = ~n15289 & ~n37972;
  assign n42945 = controllable_hmaster1 & ~n42944;
  assign n42946 = ~n15296 & ~n42945;
  assign n42947 = i_hbusreq3 & ~n42946;
  assign n42948 = ~n15300 & ~n37985;
  assign n42949 = controllable_hmaster1 & ~n42948;
  assign n42950 = ~n15307 & ~n42949;
  assign n42951 = ~i_hbusreq3 & ~n42950;
  assign n42952 = ~n42947 & ~n42951;
  assign n42953 = ~controllable_hmaster2 & ~n42952;
  assign n42954 = ~n15287 & ~n42953;
  assign n42955 = ~controllable_hgrant3 & ~n42954;
  assign n42956 = ~n14973 & ~n42955;
  assign n42957 = controllable_nhgrant0 & ~n42956;
  assign n42958 = ~n15006 & ~n42957;
  assign n42959 = ~n3281 & ~n42958;
  assign n42960 = ~n3950 & ~n42959;
  assign n42961 = n3378 & ~n42960;
  assign n42962 = ~n9388 & ~n39823;
  assign n42963 = controllable_hmaster1 & ~n42962;
  assign n42964 = controllable_hmaster0 & ~n42962;
  assign n42965 = ~n40188 & ~n42964;
  assign n42966 = ~controllable_hmaster1 & ~n42965;
  assign n42967 = ~n42963 & ~n42966;
  assign n42968 = i_hbusreq3 & ~n42967;
  assign n42969 = ~n15233 & ~n39839;
  assign n42970 = controllable_hmaster1 & ~n42969;
  assign n42971 = controllable_hmaster0 & ~n42969;
  assign n42972 = ~n40197 & ~n42971;
  assign n42973 = ~controllable_hmaster1 & ~n42972;
  assign n42974 = ~n42970 & ~n42973;
  assign n42975 = ~i_hbusreq3 & ~n42974;
  assign n42976 = ~n42968 & ~n42975;
  assign n42977 = controllable_hmaster2 & ~n42976;
  assign n42978 = ~n35802 & ~n37972;
  assign n42979 = controllable_hmaster1 & ~n42978;
  assign n42980 = ~n35811 & ~n42979;
  assign n42981 = i_hbusreq3 & ~n42980;
  assign n42982 = ~n35815 & ~n37985;
  assign n42983 = controllable_hmaster1 & ~n42982;
  assign n42984 = ~n35825 & ~n42983;
  assign n42985 = ~i_hbusreq3 & ~n42984;
  assign n42986 = ~n42981 & ~n42985;
  assign n42987 = ~controllable_hmaster2 & ~n42986;
  assign n42988 = ~n42977 & ~n42987;
  assign n42989 = ~controllable_hgrant3 & ~n42988;
  assign n42990 = ~n5402 & ~n42989;
  assign n42991 = controllable_nhgrant0 & ~n42990;
  assign n42992 = ~n5534 & ~n42991;
  assign n42993 = ~n3281 & ~n42992;
  assign n42994 = ~n3950 & ~n42993;
  assign n42995 = ~n3378 & ~n42994;
  assign n42996 = ~n42961 & ~n42995;
  assign n42997 = n3492 & ~n42996;
  assign n42998 = ~n3631 & ~n42997;
  assign n42999 = n3485 & ~n42998;
  assign n43000 = ~n3630 & ~n42999;
  assign n43001 = ~n3476 & ~n43000;
  assign n43002 = ~n6786 & ~n39881;
  assign n43003 = ~controllable_hmaster0 & ~n43002;
  assign n43004 = ~n15387 & ~n43003;
  assign n43005 = controllable_hmaster1 & ~n43004;
  assign n43006 = ~n15394 & ~n43005;
  assign n43007 = i_hbusreq3 & ~n43006;
  assign n43008 = ~n6813 & ~n39892;
  assign n43009 = ~controllable_hmaster0 & ~n43008;
  assign n43010 = ~n15398 & ~n43009;
  assign n43011 = controllable_hmaster1 & ~n43010;
  assign n43012 = ~n15407 & ~n43011;
  assign n43013 = ~i_hbusreq3 & ~n43012;
  assign n43014 = ~n43007 & ~n43013;
  assign n43015 = ~controllable_hmaster2 & ~n43014;
  assign n43016 = ~n15385 & ~n43015;
  assign n43017 = ~controllable_hgrant3 & ~n43016;
  assign n43018 = ~n15042 & ~n43017;
  assign n43019 = controllable_nhgrant0 & ~n43018;
  assign n43020 = ~n15088 & ~n43019;
  assign n43021 = ~n3281 & ~n43020;
  assign n43022 = ~n4089 & ~n43021;
  assign n43023 = n3378 & ~n43022;
  assign n43024 = ~n9477 & ~n37704;
  assign n43025 = controllable_hmaster1 & ~n43024;
  assign n43026 = controllable_hmaster0 & ~n43024;
  assign n43027 = ~n40252 & ~n43026;
  assign n43028 = ~controllable_hmaster1 & ~n43027;
  assign n43029 = ~n43025 & ~n43028;
  assign n43030 = i_hbusreq3 & ~n43029;
  assign n43031 = ~n15433 & ~n39921;
  assign n43032 = controllable_hmaster1 & ~n43031;
  assign n43033 = controllable_hmaster0 & ~n43031;
  assign n43034 = ~n40261 & ~n43033;
  assign n43035 = ~controllable_hmaster1 & ~n43034;
  assign n43036 = ~n43032 & ~n43035;
  assign n43037 = ~i_hbusreq3 & ~n43036;
  assign n43038 = ~n43030 & ~n43037;
  assign n43039 = controllable_hmaster2 & ~n43038;
  assign n43040 = ~n35887 & ~n38034;
  assign n43041 = controllable_hmaster1 & ~n43040;
  assign n43042 = ~n35896 & ~n43041;
  assign n43043 = i_hbusreq3 & ~n43042;
  assign n43044 = ~n6813 & ~n39945;
  assign n43045 = ~controllable_hmaster0 & ~n43044;
  assign n43046 = ~n35900 & ~n43045;
  assign n43047 = controllable_hmaster1 & ~n43046;
  assign n43048 = ~n35910 & ~n43047;
  assign n43049 = ~i_hbusreq3 & ~n43048;
  assign n43050 = ~n43043 & ~n43049;
  assign n43051 = ~controllable_hmaster2 & ~n43050;
  assign n43052 = ~n43039 & ~n43051;
  assign n43053 = ~controllable_hgrant3 & ~n43052;
  assign n43054 = ~n5861 & ~n43053;
  assign n43055 = controllable_nhgrant0 & ~n43054;
  assign n43056 = ~n6082 & ~n43055;
  assign n43057 = ~n3281 & ~n43056;
  assign n43058 = ~n4089 & ~n43057;
  assign n43059 = ~n3378 & ~n43058;
  assign n43060 = ~n43023 & ~n43059;
  assign n43061 = n3492 & ~n43060;
  assign n43062 = ~n15258 & ~n43061;
  assign n43063 = n3485 & ~n43062;
  assign n43064 = ~n15257 & ~n43063;
  assign n43065 = n3476 & ~n43064;
  assign n43066 = ~n43001 & ~n43065;
  assign n43067 = n3374 & ~n43066;
  assign n43068 = ~n42943 & ~n43067;
  assign n43069 = ~n3655 & ~n43068;
  assign n43070 = ~n42907 & ~n43069;
  assign n43071 = ~n3652 & ~n43070;
  assign n43072 = ~n42745 & ~n43071;
  assign n43073 = ~n3368 & ~n43072;
  assign n43074 = ~n3382 & ~n38143;
  assign n43075 = controllable_hmaster1 & ~n43074;
  assign n43076 = ~n5305 & ~n43075;
  assign n43077 = i_hbusreq3 & ~n43076;
  assign n43078 = ~n3401 & ~n38163;
  assign n43079 = controllable_hmaster1 & ~n43078;
  assign n43080 = ~n5334 & ~n43079;
  assign n43081 = ~i_hbusreq3 & ~n43080;
  assign n43082 = ~n43077 & ~n43081;
  assign n43083 = ~controllable_hmaster2 & ~n43082;
  assign n43084 = ~n12741 & ~n43083;
  assign n43085 = ~controllable_hgrant3 & ~n43084;
  assign n43086 = ~n15646 & ~n43085;
  assign n43087 = controllable_nhgrant0 & ~n43086;
  assign n43088 = ~n15675 & ~n43087;
  assign n43089 = ~n3281 & ~n43088;
  assign n43090 = ~n3281 & ~n43089;
  assign n43091 = n3378 & ~n43090;
  assign n43092 = ~n35053 & ~n38143;
  assign n43093 = controllable_hmaster1 & ~n43092;
  assign n43094 = ~n35064 & ~n43093;
  assign n43095 = i_hbusreq3 & ~n43094;
  assign n43096 = ~n35072 & ~n38163;
  assign n43097 = controllable_hmaster1 & ~n43096;
  assign n43098 = ~n35091 & ~n43097;
  assign n43099 = ~i_hbusreq3 & ~n43098;
  assign n43100 = ~n43095 & ~n43099;
  assign n43101 = ~controllable_hmaster2 & ~n43100;
  assign n43102 = ~n40353 & ~n43101;
  assign n43103 = ~controllable_hgrant3 & ~n43102;
  assign n43104 = ~n15687 & ~n43103;
  assign n43105 = controllable_nhgrant0 & ~n43104;
  assign n43106 = ~n15716 & ~n43105;
  assign n43107 = ~n3281 & ~n43106;
  assign n43108 = ~n3281 & ~n43107;
  assign n43109 = ~n3378 & ~n43108;
  assign n43110 = ~n43091 & ~n43109;
  assign n43111 = n3492 & ~n43110;
  assign n43112 = n3492 & ~n43111;
  assign n43113 = n3485 & ~n43112;
  assign n43114 = n3485 & ~n43113;
  assign n43115 = ~n3476 & ~n43114;
  assign n43116 = ~n5686 & ~n40380;
  assign n43117 = ~controllable_hmaster0 & ~n43116;
  assign n43118 = ~n7326 & ~n43117;
  assign n43119 = controllable_hmaster1 & ~n43118;
  assign n43120 = ~n7342 & ~n43119;
  assign n43121 = i_hbusreq3 & ~n43120;
  assign n43122 = ~n10152 & ~n40392;
  assign n43123 = ~controllable_hmaster0 & ~n43122;
  assign n43124 = ~n15754 & ~n43123;
  assign n43125 = controllable_hmaster1 & ~n43124;
  assign n43126 = ~n15763 & ~n43125;
  assign n43127 = ~i_hbusreq3 & ~n43126;
  assign n43128 = ~n43121 & ~n43127;
  assign n43129 = ~controllable_hmaster2 & ~n43128;
  assign n43130 = ~n15746 & ~n43129;
  assign n43131 = ~controllable_hgrant3 & ~n43130;
  assign n43132 = ~n15734 & ~n43131;
  assign n43133 = controllable_nhgrant0 & ~n43132;
  assign n43134 = ~n15783 & ~n43133;
  assign n43135 = ~n3281 & ~n43134;
  assign n43136 = ~n3281 & ~n43135;
  assign n43137 = n3378 & ~n43136;
  assign n43138 = ~n15796 & ~n40426;
  assign n43139 = controllable_hmaster1 & ~n43138;
  assign n43140 = controllable_hmaster0 & ~n43138;
  assign n43141 = ~n15796 & ~n40434;
  assign n43142 = ~controllable_hmaster0 & ~n43141;
  assign n43143 = ~n43140 & ~n43142;
  assign n43144 = ~controllable_hmaster1 & ~n43143;
  assign n43145 = ~n43139 & ~n43144;
  assign n43146 = ~i_hbusreq3 & ~n43145;
  assign n43147 = ~n40421 & ~n43146;
  assign n43148 = controllable_hmaster2 & ~n43147;
  assign n43149 = controllable_hmaster0 & ~n40458;
  assign n43150 = ~n5686 & ~n40445;
  assign n43151 = ~controllable_hmaster0 & ~n43150;
  assign n43152 = ~n43149 & ~n43151;
  assign n43153 = controllable_hmaster1 & ~n43152;
  assign n43154 = ~n40461 & ~n43153;
  assign n43155 = i_hbusreq3 & ~n43154;
  assign n43156 = ~n15796 & ~n40476;
  assign n43157 = controllable_hmaster0 & ~n43156;
  assign n43158 = ~n10152 & ~n40469;
  assign n43159 = ~controllable_hmaster0 & ~n43158;
  assign n43160 = ~n43157 & ~n43159;
  assign n43161 = controllable_hmaster1 & ~n43160;
  assign n43162 = ~n15796 & ~n40485;
  assign n43163 = controllable_hmaster0 & ~n43162;
  assign n43164 = ~n15822 & ~n40491;
  assign n43165 = ~controllable_hmaster0 & ~n43164;
  assign n43166 = ~n43163 & ~n43165;
  assign n43167 = ~controllable_hmaster1 & ~n43166;
  assign n43168 = ~n43161 & ~n43167;
  assign n43169 = ~i_hbusreq3 & ~n43168;
  assign n43170 = ~n43155 & ~n43169;
  assign n43171 = ~controllable_hmaster2 & ~n43170;
  assign n43172 = ~n43148 & ~n43171;
  assign n43173 = ~controllable_hgrant3 & ~n43172;
  assign n43174 = ~n15795 & ~n43173;
  assign n43175 = controllable_nhgrant0 & ~n43174;
  assign n43176 = ~n15846 & ~n43175;
  assign n43177 = ~n3281 & ~n43176;
  assign n43178 = ~n3281 & ~n43177;
  assign n43179 = ~n3378 & ~n43178;
  assign n43180 = ~n43137 & ~n43179;
  assign n43181 = n3492 & ~n43180;
  assign n43182 = n3492 & ~n43181;
  assign n43183 = n3485 & ~n43182;
  assign n43184 = n3485 & ~n43183;
  assign n43185 = n3476 & ~n43184;
  assign n43186 = ~n43115 & ~n43185;
  assign n43187 = n3374 & ~n43186;
  assign n43188 = ~n40325 & ~n43187;
  assign n43189 = n3655 & ~n43188;
  assign n43190 = ~n3382 & ~n38442;
  assign n43191 = controllable_hmaster1 & ~n43190;
  assign n43192 = ~n5305 & ~n43191;
  assign n43193 = i_hbusreq3 & ~n43192;
  assign n43194 = ~n3401 & ~n38462;
  assign n43195 = controllable_hmaster1 & ~n43194;
  assign n43196 = ~n5334 & ~n43195;
  assign n43197 = ~i_hbusreq3 & ~n43196;
  assign n43198 = ~n43193 & ~n43197;
  assign n43199 = ~controllable_hmaster2 & ~n43198;
  assign n43200 = ~n12741 & ~n43199;
  assign n43201 = ~controllable_hgrant3 & ~n43200;
  assign n43202 = ~n15646 & ~n43201;
  assign n43203 = controllable_nhgrant0 & ~n43202;
  assign n43204 = ~n15675 & ~n43203;
  assign n43205 = ~n3281 & ~n43204;
  assign n43206 = ~n3281 & ~n43205;
  assign n43207 = n3378 & ~n43206;
  assign n43208 = ~n35360 & ~n38442;
  assign n43209 = controllable_hmaster1 & ~n43208;
  assign n43210 = ~n35371 & ~n43209;
  assign n43211 = i_hbusreq3 & ~n43210;
  assign n43212 = ~n35380 & ~n38462;
  assign n43213 = controllable_hmaster1 & ~n43212;
  assign n43214 = ~n35400 & ~n43213;
  assign n43215 = ~i_hbusreq3 & ~n43214;
  assign n43216 = ~n43211 & ~n43215;
  assign n43217 = ~controllable_hmaster2 & ~n43216;
  assign n43218 = ~n40569 & ~n43217;
  assign n43219 = ~controllable_hgrant3 & ~n43218;
  assign n43220 = ~n15687 & ~n43219;
  assign n43221 = controllable_nhgrant0 & ~n43220;
  assign n43222 = ~n15716 & ~n43221;
  assign n43223 = ~n3281 & ~n43222;
  assign n43224 = ~n3281 & ~n43223;
  assign n43225 = ~n3378 & ~n43224;
  assign n43226 = ~n43207 & ~n43225;
  assign n43227 = n3492 & ~n43226;
  assign n43228 = n3492 & ~n43227;
  assign n43229 = n3485 & ~n43228;
  assign n43230 = n3485 & ~n43229;
  assign n43231 = ~n3476 & ~n43230;
  assign n43232 = ~n5686 & ~n40595;
  assign n43233 = ~controllable_hmaster0 & ~n43232;
  assign n43234 = ~n7326 & ~n43233;
  assign n43235 = controllable_hmaster1 & ~n43234;
  assign n43236 = ~n7342 & ~n43235;
  assign n43237 = i_hbusreq3 & ~n43236;
  assign n43238 = ~n10152 & ~n40606;
  assign n43239 = ~controllable_hmaster0 & ~n43238;
  assign n43240 = ~n15754 & ~n43239;
  assign n43241 = controllable_hmaster1 & ~n43240;
  assign n43242 = ~n15763 & ~n43241;
  assign n43243 = ~i_hbusreq3 & ~n43242;
  assign n43244 = ~n43237 & ~n43243;
  assign n43245 = ~controllable_hmaster2 & ~n43244;
  assign n43246 = ~n15746 & ~n43245;
  assign n43247 = ~controllable_hgrant3 & ~n43246;
  assign n43248 = ~n15734 & ~n43247;
  assign n43249 = controllable_nhgrant0 & ~n43248;
  assign n43250 = ~n15783 & ~n43249;
  assign n43251 = ~n3281 & ~n43250;
  assign n43252 = ~n3281 & ~n43251;
  assign n43253 = n3378 & ~n43252;
  assign n43254 = ~n15796 & ~n40640;
  assign n43255 = controllable_hmaster1 & ~n43254;
  assign n43256 = controllable_hmaster0 & ~n43254;
  assign n43257 = ~n15796 & ~n40648;
  assign n43258 = ~controllable_hmaster0 & ~n43257;
  assign n43259 = ~n43256 & ~n43258;
  assign n43260 = ~controllable_hmaster1 & ~n43259;
  assign n43261 = ~n43255 & ~n43260;
  assign n43262 = ~i_hbusreq3 & ~n43261;
  assign n43263 = ~n40635 & ~n43262;
  assign n43264 = controllable_hmaster2 & ~n43263;
  assign n43265 = controllable_hmaster0 & ~n40671;
  assign n43266 = ~n5686 & ~n40658;
  assign n43267 = ~controllable_hmaster0 & ~n43266;
  assign n43268 = ~n43265 & ~n43267;
  assign n43269 = controllable_hmaster1 & ~n43268;
  assign n43270 = ~n40674 & ~n43269;
  assign n43271 = i_hbusreq3 & ~n43270;
  assign n43272 = ~n15796 & ~n40688;
  assign n43273 = controllable_hmaster0 & ~n43272;
  assign n43274 = ~n10152 & ~n40681;
  assign n43275 = ~controllable_hmaster0 & ~n43274;
  assign n43276 = ~n43273 & ~n43275;
  assign n43277 = controllable_hmaster1 & ~n43276;
  assign n43278 = ~n15796 & ~n40697;
  assign n43279 = controllable_hmaster0 & ~n43278;
  assign n43280 = ~n15822 & ~n40703;
  assign n43281 = ~controllable_hmaster0 & ~n43280;
  assign n43282 = ~n43279 & ~n43281;
  assign n43283 = ~controllable_hmaster1 & ~n43282;
  assign n43284 = ~n43277 & ~n43283;
  assign n43285 = ~i_hbusreq3 & ~n43284;
  assign n43286 = ~n43271 & ~n43285;
  assign n43287 = ~controllable_hmaster2 & ~n43286;
  assign n43288 = ~n43264 & ~n43287;
  assign n43289 = ~controllable_hgrant3 & ~n43288;
  assign n43290 = ~n15795 & ~n43289;
  assign n43291 = controllable_nhgrant0 & ~n43290;
  assign n43292 = ~n15846 & ~n43291;
  assign n43293 = ~n3281 & ~n43292;
  assign n43294 = ~n3281 & ~n43293;
  assign n43295 = ~n3378 & ~n43294;
  assign n43296 = ~n43253 & ~n43295;
  assign n43297 = n3492 & ~n43296;
  assign n43298 = n3492 & ~n43297;
  assign n43299 = n3485 & ~n43298;
  assign n43300 = n3485 & ~n43299;
  assign n43301 = n3476 & ~n43300;
  assign n43302 = ~n43231 & ~n43301;
  assign n43303 = n3374 & ~n43302;
  assign n43304 = ~n40541 & ~n43303;
  assign n43305 = ~n3655 & ~n43304;
  assign n43306 = ~n43189 & ~n43305;
  assign n43307 = n3652 & ~n43306;
  assign n43308 = ~n4787 & ~n39561;
  assign n43309 = controllable_hmaster1 & ~n43308;
  assign n43310 = controllable_hmaster0 & ~n43308;
  assign n43311 = controllable_hmaster0 & ~n43310;
  assign n43312 = ~controllable_hmaster1 & ~n43311;
  assign n43313 = ~n43309 & ~n43312;
  assign n43314 = i_hbusreq3 & ~n43313;
  assign n43315 = ~n16031 & ~n39573;
  assign n43316 = controllable_hmaster1 & ~n43315;
  assign n43317 = controllable_hmaster0 & ~n43315;
  assign n43318 = controllable_hmaster0 & ~n43317;
  assign n43319 = ~controllable_hmaster1 & ~n43318;
  assign n43320 = ~n43316 & ~n43319;
  assign n43321 = ~i_hbusreq3 & ~n43320;
  assign n43322 = ~n43314 & ~n43321;
  assign n43323 = controllable_hmaster2 & ~n43322;
  assign n43324 = controllable_hmaster2 & ~n43323;
  assign n43325 = ~controllable_hgrant3 & ~n43324;
  assign n43326 = ~n7090 & ~n43325;
  assign n43327 = controllable_nhgrant0 & ~n43326;
  assign n43328 = ~n7118 & ~n43327;
  assign n43329 = ~n3281 & ~n43328;
  assign n43330 = ~n3281 & ~n43329;
  assign n43331 = ~n3378 & ~n43330;
  assign n43332 = ~n16013 & ~n43331;
  assign n43333 = n3492 & ~n43332;
  assign n43334 = n3492 & ~n43333;
  assign n43335 = n3485 & ~n43334;
  assign n43336 = n3485 & ~n43335;
  assign n43337 = ~n3374 & ~n43336;
  assign n43338 = ~n16070 & ~n38723;
  assign n43339 = controllable_hmaster1 & ~n43338;
  assign n43340 = ~n16077 & ~n43339;
  assign n43341 = i_hbusreq3 & ~n43340;
  assign n43342 = ~n16081 & ~n38736;
  assign n43343 = controllable_hmaster1 & ~n43342;
  assign n43344 = ~n16088 & ~n43343;
  assign n43345 = ~i_hbusreq3 & ~n43344;
  assign n43346 = ~n43341 & ~n43345;
  assign n43347 = ~controllable_hmaster2 & ~n43346;
  assign n43348 = ~n16068 & ~n43347;
  assign n43349 = ~controllable_hgrant3 & ~n43348;
  assign n43350 = ~n15646 & ~n43349;
  assign n43351 = controllable_nhgrant0 & ~n43350;
  assign n43352 = ~n15675 & ~n43351;
  assign n43353 = ~n3281 & ~n43352;
  assign n43354 = ~n3281 & ~n43353;
  assign n43355 = n3378 & ~n43354;
  assign n43356 = ~n4787 & ~n39621;
  assign n43357 = ~controllable_hmaster0 & ~n43356;
  assign n43358 = ~n43310 & ~n43357;
  assign n43359 = ~controllable_hmaster1 & ~n43358;
  assign n43360 = ~n43309 & ~n43359;
  assign n43361 = i_hbusreq3 & ~n43360;
  assign n43362 = ~n16031 & ~n39640;
  assign n43363 = ~controllable_hmaster0 & ~n43362;
  assign n43364 = ~n43317 & ~n43363;
  assign n43365 = ~controllable_hmaster1 & ~n43364;
  assign n43366 = ~n43316 & ~n43365;
  assign n43367 = ~i_hbusreq3 & ~n43366;
  assign n43368 = ~n43361 & ~n43367;
  assign n43369 = controllable_hmaster2 & ~n43368;
  assign n43370 = ~n4787 & ~n35051;
  assign n43371 = controllable_hmaster0 & ~n43370;
  assign n43372 = ~n38723 & ~n43371;
  assign n43373 = controllable_hmaster1 & ~n43372;
  assign n43374 = ~n4787 & ~n35059;
  assign n43375 = controllable_hmaster0 & ~n43374;
  assign n43376 = ~controllable_hmaster0 & ~n43370;
  assign n43377 = ~n43375 & ~n43376;
  assign n43378 = ~controllable_hmaster1 & ~n43377;
  assign n43379 = ~n43373 & ~n43378;
  assign n43380 = i_hbusreq3 & ~n43379;
  assign n43381 = ~n16031 & ~n35070;
  assign n43382 = controllable_hmaster0 & ~n43381;
  assign n43383 = ~n38736 & ~n43382;
  assign n43384 = controllable_hmaster1 & ~n43383;
  assign n43385 = ~n16031 & ~n35082;
  assign n43386 = controllable_hmaster0 & ~n43385;
  assign n43387 = ~n16145 & ~n35087;
  assign n43388 = ~controllable_hmaster0 & ~n43387;
  assign n43389 = ~n43386 & ~n43388;
  assign n43390 = ~controllable_hmaster1 & ~n43389;
  assign n43391 = ~n43384 & ~n43390;
  assign n43392 = ~i_hbusreq3 & ~n43391;
  assign n43393 = ~n43380 & ~n43392;
  assign n43394 = ~controllable_hmaster2 & ~n43393;
  assign n43395 = ~n43369 & ~n43394;
  assign n43396 = ~controllable_hgrant3 & ~n43395;
  assign n43397 = ~n15687 & ~n43396;
  assign n43398 = controllable_nhgrant0 & ~n43397;
  assign n43399 = ~n15716 & ~n43398;
  assign n43400 = ~n3281 & ~n43399;
  assign n43401 = ~n3281 & ~n43400;
  assign n43402 = ~n3378 & ~n43401;
  assign n43403 = ~n43355 & ~n43402;
  assign n43404 = n3492 & ~n43403;
  assign n43405 = n3492 & ~n43404;
  assign n43406 = n3485 & ~n43405;
  assign n43407 = n3485 & ~n43406;
  assign n43408 = ~n3476 & ~n43407;
  assign n43409 = ~n11066 & ~n40380;
  assign n43410 = ~controllable_hmaster0 & ~n43409;
  assign n43411 = ~n16209 & ~n43410;
  assign n43412 = controllable_hmaster1 & ~n43411;
  assign n43413 = ~n16218 & ~n43412;
  assign n43414 = i_hbusreq3 & ~n43413;
  assign n43415 = ~n11110 & ~n40392;
  assign n43416 = ~controllable_hmaster0 & ~n43415;
  assign n43417 = ~n16222 & ~n43416;
  assign n43418 = controllable_hmaster1 & ~n43417;
  assign n43419 = ~n16231 & ~n43418;
  assign n43420 = ~i_hbusreq3 & ~n43419;
  assign n43421 = ~n43414 & ~n43420;
  assign n43422 = ~controllable_hmaster2 & ~n43421;
  assign n43423 = ~n16207 & ~n43422;
  assign n43424 = ~controllable_hgrant3 & ~n43423;
  assign n43425 = ~n15734 & ~n43424;
  assign n43426 = controllable_nhgrant0 & ~n43425;
  assign n43427 = ~n15783 & ~n43426;
  assign n43428 = ~n3281 & ~n43427;
  assign n43429 = ~n3281 & ~n43428;
  assign n43430 = n3378 & ~n43429;
  assign n43431 = ~n10827 & ~n40410;
  assign n43432 = controllable_hmaster1 & ~n43431;
  assign n43433 = controllable_hmaster0 & ~n43431;
  assign n43434 = ~n10827 & ~n40415;
  assign n43435 = ~controllable_hmaster0 & ~n43434;
  assign n43436 = ~n43433 & ~n43435;
  assign n43437 = ~controllable_hmaster1 & ~n43436;
  assign n43438 = ~n43432 & ~n43437;
  assign n43439 = i_hbusreq3 & ~n43438;
  assign n43440 = ~n16274 & ~n40426;
  assign n43441 = controllable_hmaster1 & ~n43440;
  assign n43442 = controllable_hmaster0 & ~n43440;
  assign n43443 = ~n16274 & ~n40434;
  assign n43444 = ~controllable_hmaster0 & ~n43443;
  assign n43445 = ~n43442 & ~n43444;
  assign n43446 = ~controllable_hmaster1 & ~n43445;
  assign n43447 = ~n43441 & ~n43446;
  assign n43448 = ~i_hbusreq3 & ~n43447;
  assign n43449 = ~n43439 & ~n43448;
  assign n43450 = controllable_hmaster2 & ~n43449;
  assign n43451 = ~n10827 & ~n40449;
  assign n43452 = controllable_hmaster0 & ~n43451;
  assign n43453 = ~n11066 & ~n40445;
  assign n43454 = ~controllable_hmaster0 & ~n43453;
  assign n43455 = ~n43452 & ~n43454;
  assign n43456 = controllable_hmaster1 & ~n43455;
  assign n43457 = ~n10827 & ~n40455;
  assign n43458 = controllable_hmaster0 & ~n43457;
  assign n43459 = ~controllable_hmaster0 & ~n43451;
  assign n43460 = ~n43458 & ~n43459;
  assign n43461 = ~controllable_hmaster1 & ~n43460;
  assign n43462 = ~n43456 & ~n43461;
  assign n43463 = i_hbusreq3 & ~n43462;
  assign n43464 = ~n16274 & ~n40476;
  assign n43465 = controllable_hmaster0 & ~n43464;
  assign n43466 = ~n11110 & ~n40469;
  assign n43467 = ~controllable_hmaster0 & ~n43466;
  assign n43468 = ~n43465 & ~n43467;
  assign n43469 = controllable_hmaster1 & ~n43468;
  assign n43470 = ~n16274 & ~n40485;
  assign n43471 = controllable_hmaster0 & ~n43470;
  assign n43472 = ~n16330 & ~n40491;
  assign n43473 = ~controllable_hmaster0 & ~n43472;
  assign n43474 = ~n43471 & ~n43473;
  assign n43475 = ~controllable_hmaster1 & ~n43474;
  assign n43476 = ~n43469 & ~n43475;
  assign n43477 = ~i_hbusreq3 & ~n43476;
  assign n43478 = ~n43463 & ~n43477;
  assign n43479 = ~controllable_hmaster2 & ~n43478;
  assign n43480 = ~n43450 & ~n43479;
  assign n43481 = ~controllable_hgrant3 & ~n43480;
  assign n43482 = ~n15795 & ~n43481;
  assign n43483 = controllable_nhgrant0 & ~n43482;
  assign n43484 = ~n15846 & ~n43483;
  assign n43485 = ~n3281 & ~n43484;
  assign n43486 = ~n3281 & ~n43485;
  assign n43487 = ~n3378 & ~n43486;
  assign n43488 = ~n43430 & ~n43487;
  assign n43489 = n3492 & ~n43488;
  assign n43490 = ~n14836 & ~n43489;
  assign n43491 = n3485 & ~n43490;
  assign n43492 = ~n14835 & ~n43491;
  assign n43493 = n3476 & ~n43492;
  assign n43494 = ~n43408 & ~n43493;
  assign n43495 = n3374 & ~n43494;
  assign n43496 = ~n43337 & ~n43495;
  assign n43497 = n3655 & ~n43496;
  assign n43498 = ~n4787 & ~n39768;
  assign n43499 = controllable_hmaster1 & ~n43498;
  assign n43500 = controllable_hmaster0 & ~n43498;
  assign n43501 = controllable_hmaster0 & ~n43500;
  assign n43502 = ~controllable_hmaster1 & ~n43501;
  assign n43503 = ~n43499 & ~n43502;
  assign n43504 = i_hbusreq3 & ~n43503;
  assign n43505 = ~n16031 & ~n39780;
  assign n43506 = controllable_hmaster1 & ~n43505;
  assign n43507 = controllable_hmaster0 & ~n43505;
  assign n43508 = controllable_hmaster0 & ~n43507;
  assign n43509 = ~controllable_hmaster1 & ~n43508;
  assign n43510 = ~n43506 & ~n43509;
  assign n43511 = ~i_hbusreq3 & ~n43510;
  assign n43512 = ~n43504 & ~n43511;
  assign n43513 = controllable_hmaster2 & ~n43512;
  assign n43514 = controllable_hmaster2 & ~n43513;
  assign n43515 = ~controllable_hgrant3 & ~n43514;
  assign n43516 = ~n7090 & ~n43515;
  assign n43517 = controllable_nhgrant0 & ~n43516;
  assign n43518 = ~n7118 & ~n43517;
  assign n43519 = ~n3281 & ~n43518;
  assign n43520 = ~n3281 & ~n43519;
  assign n43521 = ~n3378 & ~n43520;
  assign n43522 = ~n16013 & ~n43521;
  assign n43523 = n3492 & ~n43522;
  assign n43524 = n3492 & ~n43523;
  assign n43525 = n3485 & ~n43524;
  assign n43526 = n3485 & ~n43525;
  assign n43527 = ~n3374 & ~n43526;
  assign n43528 = ~n16070 & ~n38932;
  assign n43529 = controllable_hmaster1 & ~n43528;
  assign n43530 = ~n16077 & ~n43529;
  assign n43531 = i_hbusreq3 & ~n43530;
  assign n43532 = ~n16081 & ~n38945;
  assign n43533 = controllable_hmaster1 & ~n43532;
  assign n43534 = ~n16088 & ~n43533;
  assign n43535 = ~i_hbusreq3 & ~n43534;
  assign n43536 = ~n43531 & ~n43535;
  assign n43537 = ~controllable_hmaster2 & ~n43536;
  assign n43538 = ~n16068 & ~n43537;
  assign n43539 = ~controllable_hgrant3 & ~n43538;
  assign n43540 = ~n15646 & ~n43539;
  assign n43541 = controllable_nhgrant0 & ~n43540;
  assign n43542 = ~n15675 & ~n43541;
  assign n43543 = ~n3281 & ~n43542;
  assign n43544 = ~n3281 & ~n43543;
  assign n43545 = n3378 & ~n43544;
  assign n43546 = ~n4787 & ~n39828;
  assign n43547 = ~controllable_hmaster0 & ~n43546;
  assign n43548 = ~n43500 & ~n43547;
  assign n43549 = ~controllable_hmaster1 & ~n43548;
  assign n43550 = ~n43499 & ~n43549;
  assign n43551 = i_hbusreq3 & ~n43550;
  assign n43552 = ~n16031 & ~n39847;
  assign n43553 = ~controllable_hmaster0 & ~n43552;
  assign n43554 = ~n43507 & ~n43553;
  assign n43555 = ~controllable_hmaster1 & ~n43554;
  assign n43556 = ~n43506 & ~n43555;
  assign n43557 = ~i_hbusreq3 & ~n43556;
  assign n43558 = ~n43551 & ~n43557;
  assign n43559 = controllable_hmaster2 & ~n43558;
  assign n43560 = ~n4787 & ~n35358;
  assign n43561 = controllable_hmaster0 & ~n43560;
  assign n43562 = ~n38932 & ~n43561;
  assign n43563 = controllable_hmaster1 & ~n43562;
  assign n43564 = ~n4787 & ~n35366;
  assign n43565 = controllable_hmaster0 & ~n43564;
  assign n43566 = ~controllable_hmaster0 & ~n43560;
  assign n43567 = ~n43565 & ~n43566;
  assign n43568 = ~controllable_hmaster1 & ~n43567;
  assign n43569 = ~n43563 & ~n43568;
  assign n43570 = i_hbusreq3 & ~n43569;
  assign n43571 = ~n16031 & ~n35378;
  assign n43572 = controllable_hmaster0 & ~n43571;
  assign n43573 = ~n38945 & ~n43572;
  assign n43574 = controllable_hmaster1 & ~n43573;
  assign n43575 = ~n16031 & ~n35389;
  assign n43576 = controllable_hmaster0 & ~n43575;
  assign n43577 = ~n16145 & ~n35396;
  assign n43578 = ~controllable_hmaster0 & ~n43577;
  assign n43579 = ~n43576 & ~n43578;
  assign n43580 = ~controllable_hmaster1 & ~n43579;
  assign n43581 = ~n43574 & ~n43580;
  assign n43582 = ~i_hbusreq3 & ~n43581;
  assign n43583 = ~n43570 & ~n43582;
  assign n43584 = ~controllable_hmaster2 & ~n43583;
  assign n43585 = ~n43559 & ~n43584;
  assign n43586 = ~controllable_hgrant3 & ~n43585;
  assign n43587 = ~n15687 & ~n43586;
  assign n43588 = controllable_nhgrant0 & ~n43587;
  assign n43589 = ~n15716 & ~n43588;
  assign n43590 = ~n3281 & ~n43589;
  assign n43591 = ~n3281 & ~n43590;
  assign n43592 = ~n3378 & ~n43591;
  assign n43593 = ~n43545 & ~n43592;
  assign n43594 = n3492 & ~n43593;
  assign n43595 = n3492 & ~n43594;
  assign n43596 = n3485 & ~n43595;
  assign n43597 = n3485 & ~n43596;
  assign n43598 = ~n3476 & ~n43597;
  assign n43599 = ~n11066 & ~n40595;
  assign n43600 = ~controllable_hmaster0 & ~n43599;
  assign n43601 = ~n16209 & ~n43600;
  assign n43602 = controllable_hmaster1 & ~n43601;
  assign n43603 = ~n16218 & ~n43602;
  assign n43604 = i_hbusreq3 & ~n43603;
  assign n43605 = ~n11110 & ~n40606;
  assign n43606 = ~controllable_hmaster0 & ~n43605;
  assign n43607 = ~n16222 & ~n43606;
  assign n43608 = controllable_hmaster1 & ~n43607;
  assign n43609 = ~n16231 & ~n43608;
  assign n43610 = ~i_hbusreq3 & ~n43609;
  assign n43611 = ~n43604 & ~n43610;
  assign n43612 = ~controllable_hmaster2 & ~n43611;
  assign n43613 = ~n16207 & ~n43612;
  assign n43614 = ~controllable_hgrant3 & ~n43613;
  assign n43615 = ~n15734 & ~n43614;
  assign n43616 = controllable_nhgrant0 & ~n43615;
  assign n43617 = ~n15783 & ~n43616;
  assign n43618 = ~n3281 & ~n43617;
  assign n43619 = ~n3281 & ~n43618;
  assign n43620 = n3378 & ~n43619;
  assign n43621 = ~n10827 & ~n40624;
  assign n43622 = controllable_hmaster1 & ~n43621;
  assign n43623 = controllable_hmaster0 & ~n43621;
  assign n43624 = ~n10827 & ~n40629;
  assign n43625 = ~controllable_hmaster0 & ~n43624;
  assign n43626 = ~n43623 & ~n43625;
  assign n43627 = ~controllable_hmaster1 & ~n43626;
  assign n43628 = ~n43622 & ~n43627;
  assign n43629 = i_hbusreq3 & ~n43628;
  assign n43630 = ~n16274 & ~n40640;
  assign n43631 = controllable_hmaster1 & ~n43630;
  assign n43632 = controllable_hmaster0 & ~n43630;
  assign n43633 = ~n16274 & ~n40648;
  assign n43634 = ~controllable_hmaster0 & ~n43633;
  assign n43635 = ~n43632 & ~n43634;
  assign n43636 = ~controllable_hmaster1 & ~n43635;
  assign n43637 = ~n43631 & ~n43636;
  assign n43638 = ~i_hbusreq3 & ~n43637;
  assign n43639 = ~n43629 & ~n43638;
  assign n43640 = controllable_hmaster2 & ~n43639;
  assign n43641 = ~n10827 & ~n40662;
  assign n43642 = controllable_hmaster0 & ~n43641;
  assign n43643 = ~n11066 & ~n40658;
  assign n43644 = ~controllable_hmaster0 & ~n43643;
  assign n43645 = ~n43642 & ~n43644;
  assign n43646 = controllable_hmaster1 & ~n43645;
  assign n43647 = ~n10827 & ~n40668;
  assign n43648 = controllable_hmaster0 & ~n43647;
  assign n43649 = ~controllable_hmaster0 & ~n43641;
  assign n43650 = ~n43648 & ~n43649;
  assign n43651 = ~controllable_hmaster1 & ~n43650;
  assign n43652 = ~n43646 & ~n43651;
  assign n43653 = i_hbusreq3 & ~n43652;
  assign n43654 = ~n16274 & ~n40688;
  assign n43655 = controllable_hmaster0 & ~n43654;
  assign n43656 = ~n11110 & ~n40681;
  assign n43657 = ~controllable_hmaster0 & ~n43656;
  assign n43658 = ~n43655 & ~n43657;
  assign n43659 = controllable_hmaster1 & ~n43658;
  assign n43660 = ~n16274 & ~n40697;
  assign n43661 = controllable_hmaster0 & ~n43660;
  assign n43662 = ~n16330 & ~n40703;
  assign n43663 = ~controllable_hmaster0 & ~n43662;
  assign n43664 = ~n43661 & ~n43663;
  assign n43665 = ~controllable_hmaster1 & ~n43664;
  assign n43666 = ~n43659 & ~n43665;
  assign n43667 = ~i_hbusreq3 & ~n43666;
  assign n43668 = ~n43653 & ~n43667;
  assign n43669 = ~controllable_hmaster2 & ~n43668;
  assign n43670 = ~n43640 & ~n43669;
  assign n43671 = ~controllable_hgrant3 & ~n43670;
  assign n43672 = ~n15795 & ~n43671;
  assign n43673 = controllable_nhgrant0 & ~n43672;
  assign n43674 = ~n15846 & ~n43673;
  assign n43675 = ~n3281 & ~n43674;
  assign n43676 = ~n3281 & ~n43675;
  assign n43677 = ~n3378 & ~n43676;
  assign n43678 = ~n43620 & ~n43677;
  assign n43679 = n3492 & ~n43678;
  assign n43680 = ~n14836 & ~n43679;
  assign n43681 = n3485 & ~n43680;
  assign n43682 = ~n14835 & ~n43681;
  assign n43683 = n3476 & ~n43682;
  assign n43684 = ~n43598 & ~n43683;
  assign n43685 = n3374 & ~n43684;
  assign n43686 = ~n43527 & ~n43685;
  assign n43687 = ~n3655 & ~n43686;
  assign n43688 = ~n43497 & ~n43687;
  assign n43689 = ~n3652 & ~n43688;
  assign n43690 = ~n43307 & ~n43689;
  assign n43691 = n3368 & ~n43690;
  assign n43692 = ~n43073 & ~n43691;
  assign n43693 = n3362 & ~n43692;
  assign n43694 = n3492 & ~n42584;
  assign n43695 = ~n3631 & ~n43694;
  assign n43696 = n3485 & ~n43695;
  assign n43697 = ~n3630 & ~n43696;
  assign n43698 = ~n3476 & ~n43697;
  assign n43699 = n3492 & ~n42632;
  assign n43700 = ~n3631 & ~n43699;
  assign n43701 = n3485 & ~n43700;
  assign n43702 = ~n41076 & ~n43701;
  assign n43703 = n3476 & ~n43702;
  assign n43704 = ~n43698 & ~n43703;
  assign n43705 = n3374 & ~n43704;
  assign n43706 = ~n41080 & ~n43705;
  assign n43707 = n3655 & ~n43706;
  assign n43708 = n3492 & ~n42684;
  assign n43709 = ~n3631 & ~n43708;
  assign n43710 = n3485 & ~n43709;
  assign n43711 = ~n3630 & ~n43710;
  assign n43712 = ~n3476 & ~n43711;
  assign n43713 = n3492 & ~n42732;
  assign n43714 = ~n3631 & ~n43713;
  assign n43715 = n3485 & ~n43714;
  assign n43716 = ~n41101 & ~n43715;
  assign n43717 = n3476 & ~n43716;
  assign n43718 = ~n43712 & ~n43717;
  assign n43719 = n3374 & ~n43718;
  assign n43720 = ~n41105 & ~n43719;
  assign n43721 = ~n3655 & ~n43720;
  assign n43722 = ~n43707 & ~n43721;
  assign n43723 = n3652 & ~n43722;
  assign n43724 = n3492 & ~n42768;
  assign n43725 = ~n3631 & ~n43724;
  assign n43726 = n3485 & ~n43725;
  assign n43727 = ~n3630 & ~n43726;
  assign n43728 = ~n3476 & ~n43727;
  assign n43729 = ~n16588 & ~n37091;
  assign n43730 = ~n3485 & ~n43729;
  assign n43731 = ~n15258 & ~n43724;
  assign n43732 = n3485 & ~n43731;
  assign n43733 = ~n43730 & ~n43732;
  assign n43734 = n3476 & ~n43733;
  assign n43735 = ~n43728 & ~n43734;
  assign n43736 = ~n3374 & ~n43735;
  assign n43737 = n3492 & ~n42832;
  assign n43738 = ~n3631 & ~n43737;
  assign n43739 = n3485 & ~n43738;
  assign n43740 = ~n3630 & ~n43739;
  assign n43741 = ~n3476 & ~n43740;
  assign n43742 = n3492 & ~n42896;
  assign n43743 = ~n15258 & ~n43742;
  assign n43744 = n3485 & ~n43743;
  assign n43745 = ~n43730 & ~n43744;
  assign n43746 = n3476 & ~n43745;
  assign n43747 = ~n43741 & ~n43746;
  assign n43748 = n3374 & ~n43747;
  assign n43749 = ~n43736 & ~n43748;
  assign n43750 = n3655 & ~n43749;
  assign n43751 = n3492 & ~n42930;
  assign n43752 = ~n3631 & ~n43751;
  assign n43753 = n3485 & ~n43752;
  assign n43754 = ~n3630 & ~n43753;
  assign n43755 = ~n3476 & ~n43754;
  assign n43756 = ~n16588 & ~n37132;
  assign n43757 = ~n3485 & ~n43756;
  assign n43758 = ~n15258 & ~n43751;
  assign n43759 = n3485 & ~n43758;
  assign n43760 = ~n43757 & ~n43759;
  assign n43761 = n3476 & ~n43760;
  assign n43762 = ~n43755 & ~n43761;
  assign n43763 = ~n3374 & ~n43762;
  assign n43764 = n3492 & ~n42994;
  assign n43765 = ~n3631 & ~n43764;
  assign n43766 = n3485 & ~n43765;
  assign n43767 = ~n3630 & ~n43766;
  assign n43768 = ~n3476 & ~n43767;
  assign n43769 = n3492 & ~n43058;
  assign n43770 = ~n15258 & ~n43769;
  assign n43771 = n3485 & ~n43770;
  assign n43772 = ~n43757 & ~n43771;
  assign n43773 = n3476 & ~n43772;
  assign n43774 = ~n43768 & ~n43773;
  assign n43775 = n3374 & ~n43774;
  assign n43776 = ~n43763 & ~n43775;
  assign n43777 = ~n3655 & ~n43776;
  assign n43778 = ~n43750 & ~n43777;
  assign n43779 = ~n3652 & ~n43778;
  assign n43780 = ~n43723 & ~n43779;
  assign n43781 = ~n3368 & ~n43780;
  assign n43782 = n3492 & ~n43108;
  assign n43783 = n3492 & ~n43782;
  assign n43784 = n3485 & ~n43783;
  assign n43785 = n3485 & ~n43784;
  assign n43786 = ~n3476 & ~n43785;
  assign n43787 = n3492 & ~n43178;
  assign n43788 = n3492 & ~n43787;
  assign n43789 = n3485 & ~n43788;
  assign n43790 = ~n41191 & ~n43789;
  assign n43791 = n3476 & ~n43790;
  assign n43792 = ~n43786 & ~n43791;
  assign n43793 = n3374 & ~n43792;
  assign n43794 = ~n41184 & ~n43793;
  assign n43795 = n3655 & ~n43794;
  assign n43796 = n3492 & ~n43224;
  assign n43797 = n3492 & ~n43796;
  assign n43798 = n3485 & ~n43797;
  assign n43799 = n3485 & ~n43798;
  assign n43800 = ~n3476 & ~n43799;
  assign n43801 = n3492 & ~n43294;
  assign n43802 = n3492 & ~n43801;
  assign n43803 = n3485 & ~n43802;
  assign n43804 = ~n41216 & ~n43803;
  assign n43805 = n3476 & ~n43804;
  assign n43806 = ~n43800 & ~n43805;
  assign n43807 = n3374 & ~n43806;
  assign n43808 = ~n41209 & ~n43807;
  assign n43809 = ~n3655 & ~n43808;
  assign n43810 = ~n43795 & ~n43809;
  assign n43811 = n3652 & ~n43810;
  assign n43812 = n3492 & ~n43330;
  assign n43813 = n3492 & ~n43812;
  assign n43814 = n3485 & ~n43813;
  assign n43815 = n3485 & ~n43814;
  assign n43816 = ~n3476 & ~n43815;
  assign n43817 = ~n8525 & ~n43814;
  assign n43818 = n3476 & ~n43817;
  assign n43819 = ~n43816 & ~n43818;
  assign n43820 = ~n3374 & ~n43819;
  assign n43821 = n3492 & ~n43401;
  assign n43822 = n3492 & ~n43821;
  assign n43823 = n3485 & ~n43822;
  assign n43824 = n3485 & ~n43823;
  assign n43825 = ~n3476 & ~n43824;
  assign n43826 = ~n16686 & ~n37231;
  assign n43827 = ~n3485 & ~n43826;
  assign n43828 = n3492 & ~n43486;
  assign n43829 = ~n14836 & ~n43828;
  assign n43830 = n3485 & ~n43829;
  assign n43831 = ~n43827 & ~n43830;
  assign n43832 = n3476 & ~n43831;
  assign n43833 = ~n43825 & ~n43832;
  assign n43834 = n3374 & ~n43833;
  assign n43835 = ~n43820 & ~n43834;
  assign n43836 = n3655 & ~n43835;
  assign n43837 = n3492 & ~n43520;
  assign n43838 = n3492 & ~n43837;
  assign n43839 = n3485 & ~n43838;
  assign n43840 = n3485 & ~n43839;
  assign n43841 = ~n3476 & ~n43840;
  assign n43842 = ~n8525 & ~n43839;
  assign n43843 = n3476 & ~n43842;
  assign n43844 = ~n43841 & ~n43843;
  assign n43845 = ~n3374 & ~n43844;
  assign n43846 = n3492 & ~n43591;
  assign n43847 = n3492 & ~n43846;
  assign n43848 = n3485 & ~n43847;
  assign n43849 = n3485 & ~n43848;
  assign n43850 = ~n3476 & ~n43849;
  assign n43851 = ~n16686 & ~n37258;
  assign n43852 = ~n3485 & ~n43851;
  assign n43853 = n3492 & ~n43676;
  assign n43854 = ~n14836 & ~n43853;
  assign n43855 = n3485 & ~n43854;
  assign n43856 = ~n43852 & ~n43855;
  assign n43857 = n3476 & ~n43856;
  assign n43858 = ~n43850 & ~n43857;
  assign n43859 = n3374 & ~n43858;
  assign n43860 = ~n43845 & ~n43859;
  assign n43861 = ~n3655 & ~n43860;
  assign n43862 = ~n43836 & ~n43861;
  assign n43863 = ~n3652 & ~n43862;
  assign n43864 = ~n43811 & ~n43863;
  assign n43865 = n3368 & ~n43864;
  assign n43866 = ~n43781 & ~n43865;
  assign n43867 = ~n3362 & ~n43866;
  assign n43868 = ~n43693 & ~n43867;
  assign n43869 = n3359 & ~n43868;
  assign n43870 = ~n37278 & ~n43701;
  assign n43871 = n3476 & ~n43870;
  assign n43872 = ~n43698 & ~n43871;
  assign n43873 = n3374 & ~n43872;
  assign n43874 = ~n41289 & ~n43873;
  assign n43875 = n3655 & ~n43874;
  assign n43876 = ~n37289 & ~n43715;
  assign n43877 = n3476 & ~n43876;
  assign n43878 = ~n43712 & ~n43877;
  assign n43879 = n3374 & ~n43878;
  assign n43880 = ~n41299 & ~n43879;
  assign n43881 = ~n3655 & ~n43880;
  assign n43882 = ~n43875 & ~n43881;
  assign n43883 = n3652 & ~n43882;
  assign n43884 = ~n37302 & ~n43732;
  assign n43885 = n3476 & ~n43884;
  assign n43886 = ~n43728 & ~n43885;
  assign n43887 = ~n3374 & ~n43886;
  assign n43888 = ~n37302 & ~n43744;
  assign n43889 = n3476 & ~n43888;
  assign n43890 = ~n43741 & ~n43889;
  assign n43891 = n3374 & ~n43890;
  assign n43892 = ~n43887 & ~n43891;
  assign n43893 = n3655 & ~n43892;
  assign n43894 = ~n37313 & ~n43759;
  assign n43895 = n3476 & ~n43894;
  assign n43896 = ~n43755 & ~n43895;
  assign n43897 = ~n3374 & ~n43896;
  assign n43898 = ~n37313 & ~n43771;
  assign n43899 = n3476 & ~n43898;
  assign n43900 = ~n43768 & ~n43899;
  assign n43901 = n3374 & ~n43900;
  assign n43902 = ~n43897 & ~n43901;
  assign n43903 = ~n3655 & ~n43902;
  assign n43904 = ~n43893 & ~n43903;
  assign n43905 = ~n3652 & ~n43904;
  assign n43906 = ~n43883 & ~n43905;
  assign n43907 = ~n3368 & ~n43906;
  assign n43908 = ~n37332 & ~n43789;
  assign n43909 = n3476 & ~n43908;
  assign n43910 = ~n43786 & ~n43909;
  assign n43911 = n3374 & ~n43910;
  assign n43912 = ~n41335 & ~n43911;
  assign n43913 = n3655 & ~n43912;
  assign n43914 = ~n37343 & ~n43803;
  assign n43915 = n3476 & ~n43914;
  assign n43916 = ~n43800 & ~n43915;
  assign n43917 = n3374 & ~n43916;
  assign n43918 = ~n41345 & ~n43917;
  assign n43919 = ~n3655 & ~n43918;
  assign n43920 = ~n43913 & ~n43919;
  assign n43921 = n3652 & ~n43920;
  assign n43922 = ~n8689 & ~n43814;
  assign n43923 = n3476 & ~n43922;
  assign n43924 = ~n43816 & ~n43923;
  assign n43925 = ~n3374 & ~n43924;
  assign n43926 = ~n37356 & ~n43830;
  assign n43927 = n3476 & ~n43926;
  assign n43928 = ~n43825 & ~n43927;
  assign n43929 = n3374 & ~n43928;
  assign n43930 = ~n43925 & ~n43929;
  assign n43931 = n3655 & ~n43930;
  assign n43932 = ~n8689 & ~n43839;
  assign n43933 = n3476 & ~n43932;
  assign n43934 = ~n43841 & ~n43933;
  assign n43935 = ~n3374 & ~n43934;
  assign n43936 = ~n37367 & ~n43855;
  assign n43937 = n3476 & ~n43936;
  assign n43938 = ~n43850 & ~n43937;
  assign n43939 = n3374 & ~n43938;
  assign n43940 = ~n43935 & ~n43939;
  assign n43941 = ~n3655 & ~n43940;
  assign n43942 = ~n43931 & ~n43941;
  assign n43943 = ~n3652 & ~n43942;
  assign n43944 = ~n43921 & ~n43943;
  assign n43945 = n3368 & ~n43944;
  assign n43946 = ~n43907 & ~n43945;
  assign n43947 = n3362 & ~n43946;
  assign n43948 = n3378 & ~n42584;
  assign n43949 = ~n37472 & ~n43948;
  assign n43950 = n3492 & ~n43949;
  assign n43951 = ~n3631 & ~n43950;
  assign n43952 = n3485 & ~n43951;
  assign n43953 = ~n3630 & ~n43952;
  assign n43954 = ~n3476 & ~n43953;
  assign n43955 = n3378 & ~n42632;
  assign n43956 = ~n37554 & ~n43955;
  assign n43957 = n3492 & ~n43956;
  assign n43958 = ~n37006 & ~n43957;
  assign n43959 = n3485 & ~n43958;
  assign n43960 = ~n37278 & ~n43959;
  assign n43961 = n3476 & ~n43960;
  assign n43962 = ~n43954 & ~n43961;
  assign n43963 = n3374 & ~n43962;
  assign n43964 = ~n41392 & ~n43963;
  assign n43965 = n3655 & ~n43964;
  assign n43966 = n3378 & ~n42684;
  assign n43967 = ~n37666 & ~n43966;
  assign n43968 = n3492 & ~n43967;
  assign n43969 = ~n3631 & ~n43968;
  assign n43970 = n3485 & ~n43969;
  assign n43971 = ~n3630 & ~n43970;
  assign n43972 = ~n3476 & ~n43971;
  assign n43973 = n3378 & ~n42732;
  assign n43974 = ~n37757 & ~n43973;
  assign n43975 = n3492 & ~n43974;
  assign n43976 = ~n37048 & ~n43975;
  assign n43977 = n3485 & ~n43976;
  assign n43978 = ~n37289 & ~n43977;
  assign n43979 = n3476 & ~n43978;
  assign n43980 = ~n43972 & ~n43979;
  assign n43981 = n3374 & ~n43980;
  assign n43982 = ~n41423 & ~n43981;
  assign n43983 = ~n3655 & ~n43982;
  assign n43984 = ~n43965 & ~n43983;
  assign n43985 = n3652 & ~n43984;
  assign n43986 = n3378 & ~n42768;
  assign n43987 = ~n37791 & ~n43986;
  assign n43988 = n3492 & ~n43987;
  assign n43989 = ~n3631 & ~n43988;
  assign n43990 = n3485 & ~n43989;
  assign n43991 = ~n3630 & ~n43990;
  assign n43992 = ~n3476 & ~n43991;
  assign n43993 = ~n37091 & ~n43988;
  assign n43994 = n3485 & ~n43993;
  assign n43995 = ~n37302 & ~n43994;
  assign n43996 = n3476 & ~n43995;
  assign n43997 = ~n43992 & ~n43996;
  assign n43998 = ~n3374 & ~n43997;
  assign n43999 = n3378 & ~n42832;
  assign n44000 = ~n37851 & ~n43999;
  assign n44001 = n3492 & ~n44000;
  assign n44002 = ~n3631 & ~n44001;
  assign n44003 = n3485 & ~n44002;
  assign n44004 = ~n3630 & ~n44003;
  assign n44005 = ~n3476 & ~n44004;
  assign n44006 = n3378 & ~n42896;
  assign n44007 = ~n37913 & ~n44006;
  assign n44008 = n3492 & ~n44007;
  assign n44009 = ~n37091 & ~n44008;
  assign n44010 = n3485 & ~n44009;
  assign n44011 = ~n37302 & ~n44010;
  assign n44012 = n3476 & ~n44011;
  assign n44013 = ~n44005 & ~n44012;
  assign n44014 = n3374 & ~n44013;
  assign n44015 = ~n43998 & ~n44014;
  assign n44016 = n3655 & ~n44015;
  assign n44017 = n3378 & ~n42930;
  assign n44018 = ~n37945 & ~n44017;
  assign n44019 = n3492 & ~n44018;
  assign n44020 = ~n3631 & ~n44019;
  assign n44021 = n3485 & ~n44020;
  assign n44022 = ~n3630 & ~n44021;
  assign n44023 = ~n3476 & ~n44022;
  assign n44024 = ~n37132 & ~n44019;
  assign n44025 = n3485 & ~n44024;
  assign n44026 = ~n37313 & ~n44025;
  assign n44027 = n3476 & ~n44026;
  assign n44028 = ~n44023 & ~n44027;
  assign n44029 = ~n3374 & ~n44028;
  assign n44030 = n3378 & ~n42994;
  assign n44031 = ~n38005 & ~n44030;
  assign n44032 = n3492 & ~n44031;
  assign n44033 = ~n3631 & ~n44032;
  assign n44034 = n3485 & ~n44033;
  assign n44035 = ~n3630 & ~n44034;
  assign n44036 = ~n3476 & ~n44035;
  assign n44037 = n3378 & ~n43058;
  assign n44038 = ~n38067 & ~n44037;
  assign n44039 = n3492 & ~n44038;
  assign n44040 = ~n37132 & ~n44039;
  assign n44041 = n3485 & ~n44040;
  assign n44042 = ~n37313 & ~n44041;
  assign n44043 = n3476 & ~n44042;
  assign n44044 = ~n44036 & ~n44043;
  assign n44045 = n3374 & ~n44044;
  assign n44046 = ~n44029 & ~n44045;
  assign n44047 = ~n3655 & ~n44046;
  assign n44048 = ~n44016 & ~n44047;
  assign n44049 = ~n3652 & ~n44048;
  assign n44050 = ~n43985 & ~n44049;
  assign n44051 = ~n3368 & ~n44050;
  assign n44052 = n3378 & ~n43108;
  assign n44053 = ~n38186 & ~n44052;
  assign n44054 = n3492 & ~n44053;
  assign n44055 = n3492 & ~n44054;
  assign n44056 = n3485 & ~n44055;
  assign n44057 = n3485 & ~n44056;
  assign n44058 = ~n3476 & ~n44057;
  assign n44059 = ~n15796 & ~n41562;
  assign n44060 = controllable_hmaster1 & ~n44059;
  assign n44061 = controllable_hmaster0 & ~n44059;
  assign n44062 = ~n15796 & ~n41577;
  assign n44063 = ~controllable_hmaster0 & ~n44062;
  assign n44064 = ~n44061 & ~n44063;
  assign n44065 = ~controllable_hmaster1 & ~n44064;
  assign n44066 = ~n44060 & ~n44065;
  assign n44067 = ~i_hbusreq3 & ~n44066;
  assign n44068 = ~n41550 & ~n44067;
  assign n44069 = controllable_hmaster2 & ~n44068;
  assign n44070 = controllable_hmaster0 & ~n41596;
  assign n44071 = ~n38318 & ~n44070;
  assign n44072 = controllable_hmaster1 & ~n44071;
  assign n44073 = ~n41599 & ~n44072;
  assign n44074 = i_hbusreq3 & ~n44073;
  assign n44075 = ~n15796 & ~n41618;
  assign n44076 = controllable_hmaster0 & ~n44075;
  assign n44077 = ~n10152 & ~n41611;
  assign n44078 = ~controllable_hmaster0 & ~n44077;
  assign n44079 = ~n44076 & ~n44078;
  assign n44080 = controllable_hmaster1 & ~n44079;
  assign n44081 = ~n15796 & ~n41627;
  assign n44082 = controllable_hmaster0 & ~n44081;
  assign n44083 = ~n15822 & ~n41639;
  assign n44084 = ~controllable_hmaster0 & ~n44083;
  assign n44085 = ~n44082 & ~n44084;
  assign n44086 = ~controllable_hmaster1 & ~n44085;
  assign n44087 = ~n44080 & ~n44086;
  assign n44088 = ~i_hbusreq3 & ~n44087;
  assign n44089 = ~n44074 & ~n44088;
  assign n44090 = ~controllable_hmaster2 & ~n44089;
  assign n44091 = ~n44069 & ~n44090;
  assign n44092 = ~controllable_hgrant3 & ~n44091;
  assign n44093 = ~n15795 & ~n44092;
  assign n44094 = controllable_nhgrant0 & ~n44093;
  assign n44095 = ~n16962 & ~n44094;
  assign n44096 = ~n3281 & ~n44095;
  assign n44097 = ~n3281 & ~n44096;
  assign n44098 = n3378 & ~n44097;
  assign n44099 = ~n38371 & ~n44098;
  assign n44100 = n3492 & ~n44099;
  assign n44101 = ~n37174 & ~n44100;
  assign n44102 = n3485 & ~n44101;
  assign n44103 = ~n37332 & ~n44102;
  assign n44104 = n3476 & ~n44103;
  assign n44105 = ~n44058 & ~n44104;
  assign n44106 = n3374 & ~n44105;
  assign n44107 = ~n41522 & ~n44106;
  assign n44108 = n3655 & ~n44107;
  assign n44109 = n3378 & ~n43224;
  assign n44110 = ~n38485 & ~n44109;
  assign n44111 = n3492 & ~n44110;
  assign n44112 = n3492 & ~n44111;
  assign n44113 = n3485 & ~n44112;
  assign n44114 = n3485 & ~n44113;
  assign n44115 = ~n3476 & ~n44114;
  assign n44116 = ~n15796 & ~n41703;
  assign n44117 = controllable_hmaster1 & ~n44116;
  assign n44118 = controllable_hmaster0 & ~n44116;
  assign n44119 = ~n15796 & ~n41711;
  assign n44120 = ~controllable_hmaster0 & ~n44119;
  assign n44121 = ~n44118 & ~n44120;
  assign n44122 = ~controllable_hmaster1 & ~n44121;
  assign n44123 = ~n44117 & ~n44122;
  assign n44124 = ~i_hbusreq3 & ~n44123;
  assign n44125 = ~n41698 & ~n44124;
  assign n44126 = controllable_hmaster2 & ~n44125;
  assign n44127 = controllable_hmaster0 & ~n41730;
  assign n44128 = ~n38611 & ~n44127;
  assign n44129 = controllable_hmaster1 & ~n44128;
  assign n44130 = ~n41733 & ~n44129;
  assign n44131 = i_hbusreq3 & ~n44130;
  assign n44132 = ~n15796 & ~n41746;
  assign n44133 = controllable_hmaster0 & ~n44132;
  assign n44134 = ~n10152 & ~n41739;
  assign n44135 = ~controllable_hmaster0 & ~n44134;
  assign n44136 = ~n44133 & ~n44135;
  assign n44137 = controllable_hmaster1 & ~n44136;
  assign n44138 = ~n15796 & ~n41755;
  assign n44139 = controllable_hmaster0 & ~n44138;
  assign n44140 = ~n15822 & ~n41761;
  assign n44141 = ~controllable_hmaster0 & ~n44140;
  assign n44142 = ~n44139 & ~n44141;
  assign n44143 = ~controllable_hmaster1 & ~n44142;
  assign n44144 = ~n44137 & ~n44143;
  assign n44145 = ~i_hbusreq3 & ~n44144;
  assign n44146 = ~n44131 & ~n44145;
  assign n44147 = ~controllable_hmaster2 & ~n44146;
  assign n44148 = ~n44126 & ~n44147;
  assign n44149 = ~controllable_hgrant3 & ~n44148;
  assign n44150 = ~n15795 & ~n44149;
  assign n44151 = controllable_nhgrant0 & ~n44150;
  assign n44152 = ~n16962 & ~n44151;
  assign n44153 = ~n3281 & ~n44152;
  assign n44154 = ~n3281 & ~n44153;
  assign n44155 = n3378 & ~n44154;
  assign n44156 = ~n38659 & ~n44155;
  assign n44157 = n3492 & ~n44156;
  assign n44158 = ~n37202 & ~n44157;
  assign n44159 = n3485 & ~n44158;
  assign n44160 = ~n37343 & ~n44159;
  assign n44161 = n3476 & ~n44160;
  assign n44162 = ~n44115 & ~n44161;
  assign n44163 = n3374 & ~n44162;
  assign n44164 = ~n41678 & ~n44163;
  assign n44165 = ~n3655 & ~n44164;
  assign n44166 = ~n44108 & ~n44165;
  assign n44167 = n3652 & ~n44166;
  assign n44168 = n3378 & ~n43330;
  assign n44169 = ~n38696 & ~n44168;
  assign n44170 = n3492 & ~n44169;
  assign n44171 = n3492 & ~n44170;
  assign n44172 = n3485 & ~n44171;
  assign n44173 = n3485 & ~n44172;
  assign n44174 = ~n3476 & ~n44173;
  assign n44175 = ~n8523 & ~n44170;
  assign n44176 = n3485 & ~n44175;
  assign n44177 = ~n8689 & ~n44176;
  assign n44178 = n3476 & ~n44177;
  assign n44179 = ~n44174 & ~n44178;
  assign n44180 = ~n3374 & ~n44179;
  assign n44181 = n3378 & ~n43401;
  assign n44182 = ~n38754 & ~n44181;
  assign n44183 = n3492 & ~n44182;
  assign n44184 = n3492 & ~n44183;
  assign n44185 = n3485 & ~n44184;
  assign n44186 = n3485 & ~n44185;
  assign n44187 = ~n3476 & ~n44186;
  assign n44188 = ~n10827 & ~n41535;
  assign n44189 = controllable_hmaster1 & ~n44188;
  assign n44190 = controllable_hmaster0 & ~n44188;
  assign n44191 = ~n10827 & ~n41544;
  assign n44192 = ~controllable_hmaster0 & ~n44191;
  assign n44193 = ~n44190 & ~n44192;
  assign n44194 = ~controllable_hmaster1 & ~n44193;
  assign n44195 = ~n44189 & ~n44194;
  assign n44196 = i_hbusreq3 & ~n44195;
  assign n44197 = ~n16274 & ~n41562;
  assign n44198 = controllable_hmaster1 & ~n44197;
  assign n44199 = controllable_hmaster0 & ~n44197;
  assign n44200 = ~n16274 & ~n41577;
  assign n44201 = ~controllable_hmaster0 & ~n44200;
  assign n44202 = ~n44199 & ~n44201;
  assign n44203 = ~controllable_hmaster1 & ~n44202;
  assign n44204 = ~n44198 & ~n44203;
  assign n44205 = ~i_hbusreq3 & ~n44204;
  assign n44206 = ~n44196 & ~n44205;
  assign n44207 = controllable_hmaster2 & ~n44206;
  assign n44208 = ~n10827 & ~n41587;
  assign n44209 = controllable_hmaster0 & ~n44208;
  assign n44210 = ~n38837 & ~n44209;
  assign n44211 = controllable_hmaster1 & ~n44210;
  assign n44212 = ~n10827 & ~n41593;
  assign n44213 = controllable_hmaster0 & ~n44212;
  assign n44214 = ~controllable_hmaster0 & ~n44208;
  assign n44215 = ~n44213 & ~n44214;
  assign n44216 = ~controllable_hmaster1 & ~n44215;
  assign n44217 = ~n44211 & ~n44216;
  assign n44218 = i_hbusreq3 & ~n44217;
  assign n44219 = ~n16274 & ~n41618;
  assign n44220 = controllable_hmaster0 & ~n44219;
  assign n44221 = ~n11110 & ~n41611;
  assign n44222 = ~controllable_hmaster0 & ~n44221;
  assign n44223 = ~n44220 & ~n44222;
  assign n44224 = controllable_hmaster1 & ~n44223;
  assign n44225 = ~n16274 & ~n41627;
  assign n44226 = controllable_hmaster0 & ~n44225;
  assign n44227 = ~n16330 & ~n41639;
  assign n44228 = ~controllable_hmaster0 & ~n44227;
  assign n44229 = ~n44226 & ~n44228;
  assign n44230 = ~controllable_hmaster1 & ~n44229;
  assign n44231 = ~n44224 & ~n44230;
  assign n44232 = ~i_hbusreq3 & ~n44231;
  assign n44233 = ~n44218 & ~n44232;
  assign n44234 = ~controllable_hmaster2 & ~n44233;
  assign n44235 = ~n44207 & ~n44234;
  assign n44236 = ~controllable_hgrant3 & ~n44235;
  assign n44237 = ~n15795 & ~n44236;
  assign n44238 = controllable_nhgrant0 & ~n44237;
  assign n44239 = ~n16962 & ~n44238;
  assign n44240 = ~n3281 & ~n44239;
  assign n44241 = ~n3281 & ~n44240;
  assign n44242 = n3378 & ~n44241;
  assign n44243 = ~n38870 & ~n44242;
  assign n44244 = n3492 & ~n44243;
  assign n44245 = ~n37231 & ~n44244;
  assign n44246 = n3485 & ~n44245;
  assign n44247 = ~n37356 & ~n44246;
  assign n44248 = n3476 & ~n44247;
  assign n44249 = ~n44187 & ~n44248;
  assign n44250 = n3374 & ~n44249;
  assign n44251 = ~n44180 & ~n44250;
  assign n44252 = n3655 & ~n44251;
  assign n44253 = n3378 & ~n43520;
  assign n44254 = ~n38905 & ~n44253;
  assign n44255 = n3492 & ~n44254;
  assign n44256 = n3492 & ~n44255;
  assign n44257 = n3485 & ~n44256;
  assign n44258 = n3485 & ~n44257;
  assign n44259 = ~n3476 & ~n44258;
  assign n44260 = ~n8523 & ~n44255;
  assign n44261 = n3485 & ~n44260;
  assign n44262 = ~n8689 & ~n44261;
  assign n44263 = n3476 & ~n44262;
  assign n44264 = ~n44259 & ~n44263;
  assign n44265 = ~n3374 & ~n44264;
  assign n44266 = n3378 & ~n43591;
  assign n44267 = ~n38963 & ~n44266;
  assign n44268 = n3492 & ~n44267;
  assign n44269 = n3492 & ~n44268;
  assign n44270 = n3485 & ~n44269;
  assign n44271 = n3485 & ~n44270;
  assign n44272 = ~n3476 & ~n44271;
  assign n44273 = ~n10827 & ~n41687;
  assign n44274 = controllable_hmaster1 & ~n44273;
  assign n44275 = controllable_hmaster0 & ~n44273;
  assign n44276 = ~n10827 & ~n41692;
  assign n44277 = ~controllable_hmaster0 & ~n44276;
  assign n44278 = ~n44275 & ~n44277;
  assign n44279 = ~controllable_hmaster1 & ~n44278;
  assign n44280 = ~n44274 & ~n44279;
  assign n44281 = i_hbusreq3 & ~n44280;
  assign n44282 = ~n16274 & ~n41703;
  assign n44283 = controllable_hmaster1 & ~n44282;
  assign n44284 = controllable_hmaster0 & ~n44282;
  assign n44285 = ~n16274 & ~n41711;
  assign n44286 = ~controllable_hmaster0 & ~n44285;
  assign n44287 = ~n44284 & ~n44286;
  assign n44288 = ~controllable_hmaster1 & ~n44287;
  assign n44289 = ~n44283 & ~n44288;
  assign n44290 = ~i_hbusreq3 & ~n44289;
  assign n44291 = ~n44281 & ~n44290;
  assign n44292 = controllable_hmaster2 & ~n44291;
  assign n44293 = ~n10827 & ~n41721;
  assign n44294 = controllable_hmaster0 & ~n44293;
  assign n44295 = ~n39046 & ~n44294;
  assign n44296 = controllable_hmaster1 & ~n44295;
  assign n44297 = ~n10827 & ~n41727;
  assign n44298 = controllable_hmaster0 & ~n44297;
  assign n44299 = ~controllable_hmaster0 & ~n44293;
  assign n44300 = ~n44298 & ~n44299;
  assign n44301 = ~controllable_hmaster1 & ~n44300;
  assign n44302 = ~n44296 & ~n44301;
  assign n44303 = i_hbusreq3 & ~n44302;
  assign n44304 = ~n16274 & ~n41746;
  assign n44305 = controllable_hmaster0 & ~n44304;
  assign n44306 = ~n11110 & ~n41739;
  assign n44307 = ~controllable_hmaster0 & ~n44306;
  assign n44308 = ~n44305 & ~n44307;
  assign n44309 = controllable_hmaster1 & ~n44308;
  assign n44310 = ~n16274 & ~n41755;
  assign n44311 = controllable_hmaster0 & ~n44310;
  assign n44312 = ~n16330 & ~n41761;
  assign n44313 = ~controllable_hmaster0 & ~n44312;
  assign n44314 = ~n44311 & ~n44313;
  assign n44315 = ~controllable_hmaster1 & ~n44314;
  assign n44316 = ~n44309 & ~n44315;
  assign n44317 = ~i_hbusreq3 & ~n44316;
  assign n44318 = ~n44303 & ~n44317;
  assign n44319 = ~controllable_hmaster2 & ~n44318;
  assign n44320 = ~n44292 & ~n44319;
  assign n44321 = ~controllable_hgrant3 & ~n44320;
  assign n44322 = ~n15795 & ~n44321;
  assign n44323 = controllable_nhgrant0 & ~n44322;
  assign n44324 = ~n16962 & ~n44323;
  assign n44325 = ~n3281 & ~n44324;
  assign n44326 = ~n3281 & ~n44325;
  assign n44327 = n3378 & ~n44326;
  assign n44328 = ~n39079 & ~n44327;
  assign n44329 = n3492 & ~n44328;
  assign n44330 = ~n37258 & ~n44329;
  assign n44331 = n3485 & ~n44330;
  assign n44332 = ~n37367 & ~n44331;
  assign n44333 = n3476 & ~n44332;
  assign n44334 = ~n44272 & ~n44333;
  assign n44335 = n3374 & ~n44334;
  assign n44336 = ~n44265 & ~n44335;
  assign n44337 = ~n3655 & ~n44336;
  assign n44338 = ~n44252 & ~n44337;
  assign n44339 = ~n3652 & ~n44338;
  assign n44340 = ~n44167 & ~n44339;
  assign n44341 = n3368 & ~n44340;
  assign n44342 = ~n44051 & ~n44341;
  assign n44343 = ~n3362 & ~n44342;
  assign n44344 = ~n43947 & ~n44343;
  assign n44345 = ~n3359 & ~n44344;
  assign n44346 = ~n43869 & ~n44345;
  assign n44347 = ~n3356 & ~n44346;
  assign n44348 = ~n42543 & ~n44347;
  assign n44349 = n3345 & ~n44348;
  assign n44350 = ~n41973 & ~n44349;
  assign n44351 = n3341 & ~n44350;
  assign n44352 = ~n39103 & ~n44351;
  assign n44353 = ~n3337 & ~n44352;
  assign n44354 = controllable_hmaster0 & ~n37429;
  assign n44355 = ~controllable_hmaster1 & ~n44354;
  assign n44356 = ~controllable_hmaster1 & ~n44355;
  assign n44357 = i_hbusreq3 & ~n44356;
  assign n44358 = controllable_hmaster0 & ~n37452;
  assign n44359 = ~controllable_hmaster1 & ~n44358;
  assign n44360 = ~controllable_hmaster1 & ~n44359;
  assign n44361 = ~i_hbusreq3 & ~n44360;
  assign n44362 = ~n44357 & ~n44361;
  assign n44363 = ~controllable_hmaster2 & ~n44362;
  assign n44364 = ~controllable_hmaster2 & ~n44363;
  assign n44365 = ~controllable_hgrant3 & ~n44364;
  assign n44366 = ~n17276 & ~n44365;
  assign n44367 = controllable_nhgrant0 & ~n44366;
  assign n44368 = ~n17300 & ~n44367;
  assign n44369 = ~n3281 & ~n44368;
  assign n44370 = ~n3281 & ~n44369;
  assign n44371 = n3378 & ~n44370;
  assign n44372 = ~n3530 & ~n44363;
  assign n44373 = ~controllable_hgrant3 & ~n44372;
  assign n44374 = ~n17306 & ~n44373;
  assign n44375 = controllable_nhgrant0 & ~n44374;
  assign n44376 = ~n17314 & ~n44375;
  assign n44377 = ~n3281 & ~n44376;
  assign n44378 = ~n3950 & ~n44377;
  assign n44379 = ~n3378 & ~n44378;
  assign n44380 = ~n44371 & ~n44379;
  assign n44381 = n3492 & ~n44380;
  assign n44382 = ~n3493 & ~n44381;
  assign n44383 = n3485 & ~n44382;
  assign n44384 = ~n3486 & ~n44383;
  assign n44385 = ~n3476 & ~n44384;
  assign n44386 = ~n17365 & ~n34986;
  assign n44387 = ~controllable_hgrant2 & ~n44386;
  assign n44388 = ~n3410 & ~n44387;
  assign n44389 = controllable_hmaster0 & ~n44388;
  assign n44390 = ~n17370 & ~n44389;
  assign n44391 = ~controllable_hmaster1 & ~n44390;
  assign n44392 = ~n17360 & ~n44391;
  assign n44393 = i_hbusreq3 & ~n44392;
  assign n44394 = i_hbusreq2 & ~n44386;
  assign n44395 = ~n17391 & ~n35078;
  assign n44396 = ~i_hbusreq2 & ~n44395;
  assign n44397 = ~n44394 & ~n44396;
  assign n44398 = ~controllable_hgrant2 & ~n44397;
  assign n44399 = ~n3859 & ~n44398;
  assign n44400 = controllable_hmaster0 & ~n44399;
  assign n44401 = ~n17398 & ~n44400;
  assign n44402 = ~controllable_hmaster1 & ~n44401;
  assign n44403 = ~n17375 & ~n44402;
  assign n44404 = ~i_hbusreq3 & ~n44403;
  assign n44405 = ~n44393 & ~n44404;
  assign n44406 = ~controllable_hmaster2 & ~n44405;
  assign n44407 = ~n17359 & ~n44406;
  assign n44408 = ~controllable_hgrant3 & ~n44407;
  assign n44409 = ~n17276 & ~n44408;
  assign n44410 = controllable_nhgrant0 & ~n44409;
  assign n44411 = ~n17300 & ~n44410;
  assign n44412 = ~n3281 & ~n44411;
  assign n44413 = ~n3281 & ~n44412;
  assign n44414 = n3378 & ~n44413;
  assign n44415 = ~n8987 & ~n34986;
  assign n44416 = ~controllable_hgrant2 & ~n44415;
  assign n44417 = ~n3410 & ~n44416;
  assign n44418 = controllable_hmaster0 & ~n44417;
  assign n44419 = ~n17423 & ~n44418;
  assign n44420 = ~controllable_hmaster1 & ~n44419;
  assign n44421 = ~n17474 & ~n44420;
  assign n44422 = i_hbusreq3 & ~n44421;
  assign n44423 = i_hbusreq2 & ~n44415;
  assign n44424 = ~n17499 & ~n35078;
  assign n44425 = ~i_hbusreq2 & ~n44424;
  assign n44426 = ~n44423 & ~n44425;
  assign n44427 = ~controllable_hgrant2 & ~n44426;
  assign n44428 = ~n3859 & ~n44427;
  assign n44429 = controllable_hmaster0 & ~n44428;
  assign n44430 = ~n17467 & ~n44429;
  assign n44431 = ~controllable_hmaster1 & ~n44430;
  assign n44432 = ~n17483 & ~n44431;
  assign n44433 = ~i_hbusreq3 & ~n44432;
  assign n44434 = ~n44422 & ~n44433;
  assign n44435 = ~controllable_hmaster2 & ~n44434;
  assign n44436 = ~n17473 & ~n44435;
  assign n44437 = ~controllable_hgrant3 & ~n44436;
  assign n44438 = ~n17306 & ~n44437;
  assign n44439 = controllable_nhgrant0 & ~n44438;
  assign n44440 = ~n17314 & ~n44439;
  assign n44441 = ~n3281 & ~n44440;
  assign n44442 = ~n4089 & ~n44441;
  assign n44443 = ~n3378 & ~n44442;
  assign n44444 = ~n44414 & ~n44443;
  assign n44445 = n3492 & ~n44444;
  assign n44446 = ~n3493 & ~n44445;
  assign n44447 = n3485 & ~n44446;
  assign n44448 = ~n3486 & ~n44447;
  assign n44449 = n3476 & ~n44448;
  assign n44450 = ~n44385 & ~n44449;
  assign n44451 = n3374 & ~n44450;
  assign n44452 = ~n17268 & ~n44451;
  assign n44453 = n3655 & ~n44452;
  assign n44454 = controllable_hmaster0 & ~n37623;
  assign n44455 = ~controllable_hmaster1 & ~n44454;
  assign n44456 = ~controllable_hmaster1 & ~n44455;
  assign n44457 = i_hbusreq3 & ~n44456;
  assign n44458 = controllable_hmaster0 & ~n37646;
  assign n44459 = ~controllable_hmaster1 & ~n44458;
  assign n44460 = ~controllable_hmaster1 & ~n44459;
  assign n44461 = ~i_hbusreq3 & ~n44460;
  assign n44462 = ~n44457 & ~n44461;
  assign n44463 = ~controllable_hmaster2 & ~n44462;
  assign n44464 = ~controllable_hmaster2 & ~n44463;
  assign n44465 = ~controllable_hgrant3 & ~n44464;
  assign n44466 = ~n17276 & ~n44465;
  assign n44467 = controllable_nhgrant0 & ~n44466;
  assign n44468 = ~n17300 & ~n44467;
  assign n44469 = ~n3281 & ~n44468;
  assign n44470 = ~n3281 & ~n44469;
  assign n44471 = n3378 & ~n44470;
  assign n44472 = ~n17664 & ~n44463;
  assign n44473 = ~controllable_hgrant3 & ~n44472;
  assign n44474 = ~n17306 & ~n44473;
  assign n44475 = controllable_nhgrant0 & ~n44474;
  assign n44476 = ~n17314 & ~n44475;
  assign n44477 = ~n3281 & ~n44476;
  assign n44478 = ~n3950 & ~n44477;
  assign n44479 = ~n3378 & ~n44478;
  assign n44480 = ~n44471 & ~n44479;
  assign n44481 = n3492 & ~n44480;
  assign n44482 = ~n3493 & ~n44481;
  assign n44483 = n3485 & ~n44482;
  assign n44484 = ~n3486 & ~n44483;
  assign n44485 = ~n3476 & ~n44484;
  assign n44486 = ~n17712 & ~n34986;
  assign n44487 = ~controllable_hgrant2 & ~n44486;
  assign n44488 = ~n3410 & ~n44487;
  assign n44489 = controllable_hmaster0 & ~n44488;
  assign n44490 = ~n17717 & ~n44489;
  assign n44491 = ~controllable_hmaster1 & ~n44490;
  assign n44492 = ~n17709 & ~n44491;
  assign n44493 = i_hbusreq3 & ~n44492;
  assign n44494 = i_hbusreq2 & ~n44486;
  assign n44495 = ~n17738 & ~n35078;
  assign n44496 = ~i_hbusreq2 & ~n44495;
  assign n44497 = ~n44494 & ~n44496;
  assign n44498 = ~controllable_hgrant2 & ~n44497;
  assign n44499 = ~n3859 & ~n44498;
  assign n44500 = controllable_hmaster0 & ~n44499;
  assign n44501 = ~n17745 & ~n44500;
  assign n44502 = ~controllable_hmaster1 & ~n44501;
  assign n44503 = ~n17722 & ~n44502;
  assign n44504 = ~i_hbusreq3 & ~n44503;
  assign n44505 = ~n44493 & ~n44504;
  assign n44506 = ~controllable_hmaster2 & ~n44505;
  assign n44507 = ~n17708 & ~n44506;
  assign n44508 = ~controllable_hgrant3 & ~n44507;
  assign n44509 = ~n17276 & ~n44508;
  assign n44510 = controllable_nhgrant0 & ~n44509;
  assign n44511 = ~n17300 & ~n44510;
  assign n44512 = ~n3281 & ~n44511;
  assign n44513 = ~n3281 & ~n44512;
  assign n44514 = n3378 & ~n44513;
  assign n44515 = ~n9305 & ~n34986;
  assign n44516 = ~controllable_hgrant2 & ~n44515;
  assign n44517 = ~n3410 & ~n44516;
  assign n44518 = controllable_hmaster0 & ~n44517;
  assign n44519 = ~n17770 & ~n44518;
  assign n44520 = ~controllable_hmaster1 & ~n44519;
  assign n44521 = ~n17820 & ~n44520;
  assign n44522 = i_hbusreq3 & ~n44521;
  assign n44523 = i_hbusreq2 & ~n44515;
  assign n44524 = ~n17843 & ~n35078;
  assign n44525 = ~i_hbusreq2 & ~n44524;
  assign n44526 = ~n44523 & ~n44525;
  assign n44527 = ~controllable_hgrant2 & ~n44526;
  assign n44528 = ~n3859 & ~n44527;
  assign n44529 = controllable_hmaster0 & ~n44528;
  assign n44530 = ~n17813 & ~n44529;
  assign n44531 = ~controllable_hmaster1 & ~n44530;
  assign n44532 = ~n17829 & ~n44531;
  assign n44533 = ~i_hbusreq3 & ~n44532;
  assign n44534 = ~n44522 & ~n44533;
  assign n44535 = ~controllable_hmaster2 & ~n44534;
  assign n44536 = ~n17819 & ~n44535;
  assign n44537 = ~controllable_hgrant3 & ~n44536;
  assign n44538 = ~n17306 & ~n44537;
  assign n44539 = controllable_nhgrant0 & ~n44538;
  assign n44540 = ~n17314 & ~n44539;
  assign n44541 = ~n3281 & ~n44540;
  assign n44542 = ~n4089 & ~n44541;
  assign n44543 = ~n3378 & ~n44542;
  assign n44544 = ~n44514 & ~n44543;
  assign n44545 = n3492 & ~n44544;
  assign n44546 = ~n17612 & ~n44545;
  assign n44547 = n3485 & ~n44546;
  assign n44548 = ~n17611 & ~n44547;
  assign n44549 = n3476 & ~n44548;
  assign n44550 = ~n44485 & ~n44549;
  assign n44551 = n3374 & ~n44550;
  assign n44552 = ~n17618 & ~n44551;
  assign n44553 = ~n3655 & ~n44552;
  assign n44554 = ~n44453 & ~n44553;
  assign n44555 = n3652 & ~n44554;
  assign n44556 = controllable_hmaster0 & ~n37822;
  assign n44557 = ~controllable_hmaster1 & ~n44556;
  assign n44558 = ~controllable_hmaster1 & ~n44557;
  assign n44559 = i_hbusreq3 & ~n44558;
  assign n44560 = controllable_hmaster0 & ~n37835;
  assign n44561 = ~controllable_hmaster1 & ~n44560;
  assign n44562 = ~controllable_hmaster1 & ~n44561;
  assign n44563 = ~i_hbusreq3 & ~n44562;
  assign n44564 = ~n44559 & ~n44563;
  assign n44565 = ~controllable_hmaster2 & ~n44564;
  assign n44566 = ~controllable_hmaster2 & ~n44565;
  assign n44567 = ~controllable_hgrant3 & ~n44566;
  assign n44568 = ~n17276 & ~n44567;
  assign n44569 = controllable_nhgrant0 & ~n44568;
  assign n44570 = ~n17300 & ~n44569;
  assign n44571 = ~n3281 & ~n44570;
  assign n44572 = ~n3281 & ~n44571;
  assign n44573 = n3378 & ~n44572;
  assign n44574 = ~n3530 & ~n44565;
  assign n44575 = ~controllable_hgrant3 & ~n44574;
  assign n44576 = ~n17306 & ~n44575;
  assign n44577 = controllable_nhgrant0 & ~n44576;
  assign n44578 = ~n17314 & ~n44577;
  assign n44579 = ~n3281 & ~n44578;
  assign n44580 = ~n3950 & ~n44579;
  assign n44581 = ~n3378 & ~n44580;
  assign n44582 = ~n44573 & ~n44581;
  assign n44583 = n3492 & ~n44582;
  assign n44584 = ~n3493 & ~n44583;
  assign n44585 = n3485 & ~n44584;
  assign n44586 = ~n3486 & ~n44585;
  assign n44587 = ~n3476 & ~n44586;
  assign n44588 = ~n4333 & ~n44387;
  assign n44589 = controllable_hmaster0 & ~n44588;
  assign n44590 = ~n17370 & ~n44589;
  assign n44591 = ~controllable_hmaster1 & ~n44590;
  assign n44592 = ~n17360 & ~n44591;
  assign n44593 = i_hbusreq3 & ~n44592;
  assign n44594 = ~n4340 & ~n44398;
  assign n44595 = controllable_hmaster0 & ~n44594;
  assign n44596 = ~n17398 & ~n44595;
  assign n44597 = ~controllable_hmaster1 & ~n44596;
  assign n44598 = ~n17375 & ~n44597;
  assign n44599 = ~i_hbusreq3 & ~n44598;
  assign n44600 = ~n44593 & ~n44599;
  assign n44601 = ~controllable_hmaster2 & ~n44600;
  assign n44602 = ~n17359 & ~n44601;
  assign n44603 = ~controllable_hgrant3 & ~n44602;
  assign n44604 = ~n17276 & ~n44603;
  assign n44605 = controllable_nhgrant0 & ~n44604;
  assign n44606 = ~n17300 & ~n44605;
  assign n44607 = ~n3281 & ~n44606;
  assign n44608 = ~n3281 & ~n44607;
  assign n44609 = n3378 & ~n44608;
  assign n44610 = ~n4333 & ~n44416;
  assign n44611 = controllable_hmaster0 & ~n44610;
  assign n44612 = ~n17423 & ~n44611;
  assign n44613 = ~controllable_hmaster1 & ~n44612;
  assign n44614 = ~n17474 & ~n44613;
  assign n44615 = i_hbusreq3 & ~n44614;
  assign n44616 = ~n4340 & ~n44427;
  assign n44617 = controllable_hmaster0 & ~n44616;
  assign n44618 = ~n17467 & ~n44617;
  assign n44619 = ~controllable_hmaster1 & ~n44618;
  assign n44620 = ~n17483 & ~n44619;
  assign n44621 = ~i_hbusreq3 & ~n44620;
  assign n44622 = ~n44615 & ~n44621;
  assign n44623 = ~controllable_hmaster2 & ~n44622;
  assign n44624 = ~n17473 & ~n44623;
  assign n44625 = ~controllable_hgrant3 & ~n44624;
  assign n44626 = ~n17306 & ~n44625;
  assign n44627 = controllable_nhgrant0 & ~n44626;
  assign n44628 = ~n17314 & ~n44627;
  assign n44629 = ~n3281 & ~n44628;
  assign n44630 = ~n4089 & ~n44629;
  assign n44631 = ~n3378 & ~n44630;
  assign n44632 = ~n44609 & ~n44631;
  assign n44633 = n3492 & ~n44632;
  assign n44634 = ~n3493 & ~n44633;
  assign n44635 = n3485 & ~n44634;
  assign n44636 = ~n3486 & ~n44635;
  assign n44637 = n3476 & ~n44636;
  assign n44638 = ~n44587 & ~n44637;
  assign n44639 = n3374 & ~n44638;
  assign n44640 = ~n17268 & ~n44639;
  assign n44641 = n3655 & ~n44640;
  assign n44642 = controllable_hmaster0 & ~n37976;
  assign n44643 = ~controllable_hmaster1 & ~n44642;
  assign n44644 = ~controllable_hmaster1 & ~n44643;
  assign n44645 = i_hbusreq3 & ~n44644;
  assign n44646 = controllable_hmaster0 & ~n37989;
  assign n44647 = ~controllable_hmaster1 & ~n44646;
  assign n44648 = ~controllable_hmaster1 & ~n44647;
  assign n44649 = ~i_hbusreq3 & ~n44648;
  assign n44650 = ~n44645 & ~n44649;
  assign n44651 = ~controllable_hmaster2 & ~n44650;
  assign n44652 = ~controllable_hmaster2 & ~n44651;
  assign n44653 = ~controllable_hgrant3 & ~n44652;
  assign n44654 = ~n17276 & ~n44653;
  assign n44655 = controllable_nhgrant0 & ~n44654;
  assign n44656 = ~n17300 & ~n44655;
  assign n44657 = ~n3281 & ~n44656;
  assign n44658 = ~n3281 & ~n44657;
  assign n44659 = n3378 & ~n44658;
  assign n44660 = ~n17664 & ~n44651;
  assign n44661 = ~controllable_hgrant3 & ~n44660;
  assign n44662 = ~n17306 & ~n44661;
  assign n44663 = controllable_nhgrant0 & ~n44662;
  assign n44664 = ~n17314 & ~n44663;
  assign n44665 = ~n3281 & ~n44664;
  assign n44666 = ~n3950 & ~n44665;
  assign n44667 = ~n3378 & ~n44666;
  assign n44668 = ~n44659 & ~n44667;
  assign n44669 = n3492 & ~n44668;
  assign n44670 = ~n3493 & ~n44669;
  assign n44671 = n3485 & ~n44670;
  assign n44672 = ~n3486 & ~n44671;
  assign n44673 = ~n3476 & ~n44672;
  assign n44674 = ~n4333 & ~n44487;
  assign n44675 = controllable_hmaster0 & ~n44674;
  assign n44676 = ~n17717 & ~n44675;
  assign n44677 = ~controllable_hmaster1 & ~n44676;
  assign n44678 = ~n17709 & ~n44677;
  assign n44679 = i_hbusreq3 & ~n44678;
  assign n44680 = ~n4340 & ~n44498;
  assign n44681 = controllable_hmaster0 & ~n44680;
  assign n44682 = ~n17745 & ~n44681;
  assign n44683 = ~controllable_hmaster1 & ~n44682;
  assign n44684 = ~n17722 & ~n44683;
  assign n44685 = ~i_hbusreq3 & ~n44684;
  assign n44686 = ~n44679 & ~n44685;
  assign n44687 = ~controllable_hmaster2 & ~n44686;
  assign n44688 = ~n17708 & ~n44687;
  assign n44689 = ~controllable_hgrant3 & ~n44688;
  assign n44690 = ~n17276 & ~n44689;
  assign n44691 = controllable_nhgrant0 & ~n44690;
  assign n44692 = ~n17300 & ~n44691;
  assign n44693 = ~n3281 & ~n44692;
  assign n44694 = ~n3281 & ~n44693;
  assign n44695 = n3378 & ~n44694;
  assign n44696 = ~n4333 & ~n44516;
  assign n44697 = controllable_hmaster0 & ~n44696;
  assign n44698 = ~n17770 & ~n44697;
  assign n44699 = ~controllable_hmaster1 & ~n44698;
  assign n44700 = ~n17820 & ~n44699;
  assign n44701 = i_hbusreq3 & ~n44700;
  assign n44702 = ~n4340 & ~n44527;
  assign n44703 = controllable_hmaster0 & ~n44702;
  assign n44704 = ~n17813 & ~n44703;
  assign n44705 = ~controllable_hmaster1 & ~n44704;
  assign n44706 = ~n17829 & ~n44705;
  assign n44707 = ~i_hbusreq3 & ~n44706;
  assign n44708 = ~n44701 & ~n44707;
  assign n44709 = ~controllable_hmaster2 & ~n44708;
  assign n44710 = ~n17819 & ~n44709;
  assign n44711 = ~controllable_hgrant3 & ~n44710;
  assign n44712 = ~n17306 & ~n44711;
  assign n44713 = controllable_nhgrant0 & ~n44712;
  assign n44714 = ~n17314 & ~n44713;
  assign n44715 = ~n3281 & ~n44714;
  assign n44716 = ~n4089 & ~n44715;
  assign n44717 = ~n3378 & ~n44716;
  assign n44718 = ~n44695 & ~n44717;
  assign n44719 = n3492 & ~n44718;
  assign n44720 = ~n17612 & ~n44719;
  assign n44721 = n3485 & ~n44720;
  assign n44722 = ~n17611 & ~n44721;
  assign n44723 = n3476 & ~n44722;
  assign n44724 = ~n44673 & ~n44723;
  assign n44725 = n3374 & ~n44724;
  assign n44726 = ~n17618 & ~n44725;
  assign n44727 = ~n3655 & ~n44726;
  assign n44728 = ~n44641 & ~n44727;
  assign n44729 = ~n3652 & ~n44728;
  assign n44730 = ~n44555 & ~n44729;
  assign n44731 = ~n3368 & ~n44730;
  assign n44732 = controllable_hmaster0 & ~n38149;
  assign n44733 = ~controllable_hmaster1 & ~n44732;
  assign n44734 = ~controllable_hmaster1 & ~n44733;
  assign n44735 = i_hbusreq3 & ~n44734;
  assign n44736 = controllable_hmaster0 & ~n38172;
  assign n44737 = ~controllable_hmaster1 & ~n44736;
  assign n44738 = ~controllable_hmaster1 & ~n44737;
  assign n44739 = ~i_hbusreq3 & ~n44738;
  assign n44740 = ~n44735 & ~n44739;
  assign n44741 = ~controllable_hmaster2 & ~n44740;
  assign n44742 = ~controllable_hmaster2 & ~n44741;
  assign n44743 = ~controllable_hgrant3 & ~n44742;
  assign n44744 = ~n18057 & ~n44743;
  assign n44745 = controllable_nhgrant0 & ~n44744;
  assign n44746 = ~n18077 & ~n44745;
  assign n44747 = ~n3281 & ~n44746;
  assign n44748 = ~n3281 & ~n44747;
  assign n44749 = n3492 & ~n44748;
  assign n44750 = n3492 & ~n44749;
  assign n44751 = n3485 & ~n44750;
  assign n44752 = n3485 & ~n44751;
  assign n44753 = ~n3476 & ~n44752;
  assign n44754 = ~n17365 & ~n35937;
  assign n44755 = ~controllable_hgrant2 & ~n44754;
  assign n44756 = ~n3410 & ~n44755;
  assign n44757 = controllable_hmaster0 & ~n44756;
  assign n44758 = ~n17370 & ~n44757;
  assign n44759 = ~controllable_hmaster1 & ~n44758;
  assign n44760 = ~n17360 & ~n44759;
  assign n44761 = i_hbusreq3 & ~n44760;
  assign n44762 = i_hbusreq2 & ~n44754;
  assign n44763 = ~n18099 & ~n38093;
  assign n44764 = ~i_hbusreq2 & ~n44763;
  assign n44765 = ~n44762 & ~n44764;
  assign n44766 = ~controllable_hgrant2 & ~n44765;
  assign n44767 = ~n4562 & ~n44766;
  assign n44768 = controllable_hmaster0 & ~n44767;
  assign n44769 = ~n17370 & ~n44768;
  assign n44770 = ~controllable_hmaster1 & ~n44769;
  assign n44771 = ~n17360 & ~n44770;
  assign n44772 = ~i_hbusreq3 & ~n44771;
  assign n44773 = ~n44761 & ~n44772;
  assign n44774 = ~controllable_hmaster2 & ~n44773;
  assign n44775 = ~n18086 & ~n44774;
  assign n44776 = ~controllable_hgrant3 & ~n44775;
  assign n44777 = ~n18057 & ~n44776;
  assign n44778 = controllable_nhgrant0 & ~n44777;
  assign n44779 = ~n18077 & ~n44778;
  assign n44780 = ~n3281 & ~n44779;
  assign n44781 = ~n3281 & ~n44780;
  assign n44782 = n3492 & ~n44781;
  assign n44783 = n3492 & ~n44782;
  assign n44784 = n3485 & ~n44783;
  assign n44785 = n3485 & ~n44784;
  assign n44786 = n3476 & ~n44785;
  assign n44787 = ~n44753 & ~n44786;
  assign n44788 = n3374 & ~n44787;
  assign n44789 = n3374 & ~n44788;
  assign n44790 = n3655 & ~n44789;
  assign n44791 = controllable_hmaster0 & ~n38448;
  assign n44792 = ~controllable_hmaster1 & ~n44791;
  assign n44793 = ~controllable_hmaster1 & ~n44792;
  assign n44794 = i_hbusreq3 & ~n44793;
  assign n44795 = controllable_hmaster0 & ~n38471;
  assign n44796 = ~controllable_hmaster1 & ~n44795;
  assign n44797 = ~controllable_hmaster1 & ~n44796;
  assign n44798 = ~i_hbusreq3 & ~n44797;
  assign n44799 = ~n44794 & ~n44798;
  assign n44800 = ~controllable_hmaster2 & ~n44799;
  assign n44801 = ~controllable_hmaster2 & ~n44800;
  assign n44802 = ~controllable_hgrant3 & ~n44801;
  assign n44803 = ~n18057 & ~n44802;
  assign n44804 = controllable_nhgrant0 & ~n44803;
  assign n44805 = ~n18077 & ~n44804;
  assign n44806 = ~n3281 & ~n44805;
  assign n44807 = ~n3281 & ~n44806;
  assign n44808 = n3492 & ~n44807;
  assign n44809 = n3492 & ~n44808;
  assign n44810 = n3485 & ~n44809;
  assign n44811 = n3485 & ~n44810;
  assign n44812 = ~n3476 & ~n44811;
  assign n44813 = ~n18191 & ~n35937;
  assign n44814 = ~controllable_hgrant2 & ~n44813;
  assign n44815 = ~n3410 & ~n44814;
  assign n44816 = controllable_hmaster0 & ~n44815;
  assign n44817 = ~n18196 & ~n44816;
  assign n44818 = ~controllable_hmaster1 & ~n44817;
  assign n44819 = ~n18184 & ~n44818;
  assign n44820 = i_hbusreq3 & ~n44819;
  assign n44821 = i_hbusreq2 & ~n44813;
  assign n44822 = ~n18223 & ~n38093;
  assign n44823 = ~i_hbusreq2 & ~n44822;
  assign n44824 = ~n44821 & ~n44823;
  assign n44825 = ~controllable_hgrant2 & ~n44824;
  assign n44826 = ~n4562 & ~n44825;
  assign n44827 = controllable_hmaster0 & ~n44826;
  assign n44828 = ~n18230 & ~n44827;
  assign n44829 = ~controllable_hmaster1 & ~n44828;
  assign n44830 = ~n18201 & ~n44829;
  assign n44831 = ~i_hbusreq3 & ~n44830;
  assign n44832 = ~n44820 & ~n44831;
  assign n44833 = ~controllable_hmaster2 & ~n44832;
  assign n44834 = ~n18183 & ~n44833;
  assign n44835 = ~controllable_hgrant3 & ~n44834;
  assign n44836 = ~n18057 & ~n44835;
  assign n44837 = controllable_nhgrant0 & ~n44836;
  assign n44838 = ~n18077 & ~n44837;
  assign n44839 = ~n3281 & ~n44838;
  assign n44840 = ~n3281 & ~n44839;
  assign n44841 = n3492 & ~n44840;
  assign n44842 = ~n18151 & ~n44841;
  assign n44843 = n3485 & ~n44842;
  assign n44844 = ~n18150 & ~n44843;
  assign n44845 = n3476 & ~n44844;
  assign n44846 = ~n44812 & ~n44845;
  assign n44847 = n3374 & ~n44846;
  assign n44848 = n3374 & ~n44847;
  assign n44849 = ~n3655 & ~n44848;
  assign n44850 = ~n44790 & ~n44849;
  assign n44851 = n3652 & ~n44850;
  assign n44852 = controllable_hmaster0 & ~n38727;
  assign n44853 = ~controllable_hmaster1 & ~n44852;
  assign n44854 = ~controllable_hmaster1 & ~n44853;
  assign n44855 = i_hbusreq3 & ~n44854;
  assign n44856 = controllable_hmaster0 & ~n38740;
  assign n44857 = ~controllable_hmaster1 & ~n44856;
  assign n44858 = ~controllable_hmaster1 & ~n44857;
  assign n44859 = ~i_hbusreq3 & ~n44858;
  assign n44860 = ~n44855 & ~n44859;
  assign n44861 = ~controllable_hmaster2 & ~n44860;
  assign n44862 = ~controllable_hmaster2 & ~n44861;
  assign n44863 = ~controllable_hgrant3 & ~n44862;
  assign n44864 = ~n18057 & ~n44863;
  assign n44865 = controllable_nhgrant0 & ~n44864;
  assign n44866 = ~n18077 & ~n44865;
  assign n44867 = ~n3281 & ~n44866;
  assign n44868 = ~n3281 & ~n44867;
  assign n44869 = n3492 & ~n44868;
  assign n44870 = n3492 & ~n44869;
  assign n44871 = n3485 & ~n44870;
  assign n44872 = n3485 & ~n44871;
  assign n44873 = ~n3476 & ~n44872;
  assign n44874 = ~n4787 & ~n44755;
  assign n44875 = controllable_hmaster0 & ~n44874;
  assign n44876 = ~n17370 & ~n44875;
  assign n44877 = ~controllable_hmaster1 & ~n44876;
  assign n44878 = ~n17360 & ~n44877;
  assign n44879 = i_hbusreq3 & ~n44878;
  assign n44880 = ~n4794 & ~n44766;
  assign n44881 = controllable_hmaster0 & ~n44880;
  assign n44882 = ~n17370 & ~n44881;
  assign n44883 = ~controllable_hmaster1 & ~n44882;
  assign n44884 = ~n17360 & ~n44883;
  assign n44885 = ~i_hbusreq3 & ~n44884;
  assign n44886 = ~n44879 & ~n44885;
  assign n44887 = ~controllable_hmaster2 & ~n44886;
  assign n44888 = ~n18086 & ~n44887;
  assign n44889 = ~controllable_hgrant3 & ~n44888;
  assign n44890 = ~n18057 & ~n44889;
  assign n44891 = controllable_nhgrant0 & ~n44890;
  assign n44892 = ~n18077 & ~n44891;
  assign n44893 = ~n3281 & ~n44892;
  assign n44894 = ~n3281 & ~n44893;
  assign n44895 = n3492 & ~n44894;
  assign n44896 = n3492 & ~n44895;
  assign n44897 = n3485 & ~n44896;
  assign n44898 = n3485 & ~n44897;
  assign n44899 = n3476 & ~n44898;
  assign n44900 = ~n44873 & ~n44899;
  assign n44901 = n3374 & ~n44900;
  assign n44902 = n3374 & ~n44901;
  assign n44903 = n3655 & ~n44902;
  assign n44904 = controllable_hmaster0 & ~n38936;
  assign n44905 = ~controllable_hmaster1 & ~n44904;
  assign n44906 = ~controllable_hmaster1 & ~n44905;
  assign n44907 = i_hbusreq3 & ~n44906;
  assign n44908 = controllable_hmaster0 & ~n38949;
  assign n44909 = ~controllable_hmaster1 & ~n44908;
  assign n44910 = ~controllable_hmaster1 & ~n44909;
  assign n44911 = ~i_hbusreq3 & ~n44910;
  assign n44912 = ~n44907 & ~n44911;
  assign n44913 = ~controllable_hmaster2 & ~n44912;
  assign n44914 = ~controllable_hmaster2 & ~n44913;
  assign n44915 = ~controllable_hgrant3 & ~n44914;
  assign n44916 = ~n18057 & ~n44915;
  assign n44917 = controllable_nhgrant0 & ~n44916;
  assign n44918 = ~n18077 & ~n44917;
  assign n44919 = ~n3281 & ~n44918;
  assign n44920 = ~n3281 & ~n44919;
  assign n44921 = n3492 & ~n44920;
  assign n44922 = n3492 & ~n44921;
  assign n44923 = n3485 & ~n44922;
  assign n44924 = n3485 & ~n44923;
  assign n44925 = ~n3476 & ~n44924;
  assign n44926 = ~n4787 & ~n44814;
  assign n44927 = controllable_hmaster0 & ~n44926;
  assign n44928 = ~n18196 & ~n44927;
  assign n44929 = ~controllable_hmaster1 & ~n44928;
  assign n44930 = ~n18184 & ~n44929;
  assign n44931 = i_hbusreq3 & ~n44930;
  assign n44932 = ~n4794 & ~n44825;
  assign n44933 = controllable_hmaster0 & ~n44932;
  assign n44934 = ~n18230 & ~n44933;
  assign n44935 = ~controllable_hmaster1 & ~n44934;
  assign n44936 = ~n18201 & ~n44935;
  assign n44937 = ~i_hbusreq3 & ~n44936;
  assign n44938 = ~n44931 & ~n44937;
  assign n44939 = ~controllable_hmaster2 & ~n44938;
  assign n44940 = ~n18183 & ~n44939;
  assign n44941 = ~controllable_hgrant3 & ~n44940;
  assign n44942 = ~n18057 & ~n44941;
  assign n44943 = controllable_nhgrant0 & ~n44942;
  assign n44944 = ~n18077 & ~n44943;
  assign n44945 = ~n3281 & ~n44944;
  assign n44946 = ~n3281 & ~n44945;
  assign n44947 = n3492 & ~n44946;
  assign n44948 = ~n18151 & ~n44947;
  assign n44949 = n3485 & ~n44948;
  assign n44950 = ~n18150 & ~n44949;
  assign n44951 = n3476 & ~n44950;
  assign n44952 = ~n44925 & ~n44951;
  assign n44953 = n3374 & ~n44952;
  assign n44954 = n3374 & ~n44953;
  assign n44955 = ~n3655 & ~n44954;
  assign n44956 = ~n44903 & ~n44955;
  assign n44957 = ~n3652 & ~n44956;
  assign n44958 = ~n44851 & ~n44957;
  assign n44959 = n3368 & ~n44958;
  assign n44960 = ~n44731 & ~n44959;
  assign n44961 = ~n3362 & ~n44960;
  assign n44962 = ~n3362 & ~n44961;
  assign n44963 = ~n3359 & ~n44962;
  assign n44964 = ~n3359 & ~n44963;
  assign n44965 = n3356 & ~n44964;
  assign n44966 = ~n18369 & ~n39590;
  assign n44967 = n3492 & ~n44966;
  assign n44968 = ~n3631 & ~n44967;
  assign n44969 = n3485 & ~n44968;
  assign n44970 = ~n3630 & ~n44969;
  assign n44971 = ~n3374 & ~n44970;
  assign n44972 = ~n3821 & ~n37429;
  assign n44973 = ~controllable_hmaster1 & ~n44972;
  assign n44974 = ~n5293 & ~n44973;
  assign n44975 = i_hbusreq3 & ~n44974;
  assign n44976 = ~n5278 & ~n37452;
  assign n44977 = ~controllable_hmaster1 & ~n44976;
  assign n44978 = ~n5313 & ~n44977;
  assign n44979 = ~i_hbusreq3 & ~n44978;
  assign n44980 = ~n44975 & ~n44979;
  assign n44981 = ~controllable_hmaster2 & ~n44980;
  assign n44982 = ~n12065 & ~n44981;
  assign n44983 = ~controllable_hgrant3 & ~n44982;
  assign n44984 = ~n18382 & ~n44983;
  assign n44985 = controllable_nhgrant0 & ~n44984;
  assign n44986 = ~n18416 & ~n44985;
  assign n44987 = ~n3281 & ~n44986;
  assign n44988 = ~n3950 & ~n44987;
  assign n44989 = n3378 & ~n44988;
  assign n44990 = ~n35062 & ~n37429;
  assign n44991 = ~controllable_hmaster1 & ~n44990;
  assign n44992 = ~n35057 & ~n44991;
  assign n44993 = i_hbusreq3 & ~n44992;
  assign n44994 = ~n35089 & ~n37452;
  assign n44995 = ~controllable_hmaster1 & ~n44994;
  assign n44996 = ~n35076 & ~n44995;
  assign n44997 = ~i_hbusreq3 & ~n44996;
  assign n44998 = ~n44993 & ~n44997;
  assign n44999 = ~controllable_hmaster2 & ~n44998;
  assign n45000 = ~n39648 & ~n44999;
  assign n45001 = ~controllable_hgrant3 & ~n45000;
  assign n45002 = ~n5402 & ~n45001;
  assign n45003 = controllable_nhgrant0 & ~n45002;
  assign n45004 = ~n5534 & ~n45003;
  assign n45005 = ~n3281 & ~n45004;
  assign n45006 = ~n3950 & ~n45005;
  assign n45007 = ~n3378 & ~n45006;
  assign n45008 = ~n44989 & ~n45007;
  assign n45009 = n3492 & ~n45008;
  assign n45010 = ~n3631 & ~n45009;
  assign n45011 = n3485 & ~n45010;
  assign n45012 = ~n3630 & ~n45011;
  assign n45013 = ~n3476 & ~n45012;
  assign n45014 = ~n8987 & ~n39673;
  assign n45015 = ~controllable_hgrant2 & ~n45014;
  assign n45016 = ~n5616 & ~n45015;
  assign n45017 = controllable_hmaster0 & ~n45016;
  assign n45018 = ~n5702 & ~n45017;
  assign n45019 = ~controllable_hmaster1 & ~n45018;
  assign n45020 = ~n5690 & ~n45019;
  assign n45021 = i_hbusreq3 & ~n45020;
  assign n45022 = i_hbusreq2 & ~n45014;
  assign n45023 = ~n17499 & ~n39683;
  assign n45024 = ~i_hbusreq2 & ~n45023;
  assign n45025 = ~n45022 & ~n45024;
  assign n45026 = ~controllable_hgrant2 & ~n45025;
  assign n45027 = ~n5657 & ~n45026;
  assign n45028 = controllable_hmaster0 & ~n45027;
  assign n45029 = ~n18502 & ~n45028;
  assign n45030 = ~controllable_hmaster1 & ~n45029;
  assign n45031 = ~n18495 & ~n45030;
  assign n45032 = ~i_hbusreq3 & ~n45031;
  assign n45033 = ~n45021 & ~n45032;
  assign n45034 = ~controllable_hmaster2 & ~n45033;
  assign n45035 = ~n18481 & ~n45034;
  assign n45036 = ~controllable_hgrant3 & ~n45035;
  assign n45037 = ~n18453 & ~n45036;
  assign n45038 = controllable_nhgrant0 & ~n45037;
  assign n45039 = ~n18526 & ~n45038;
  assign n45040 = ~n3281 & ~n45039;
  assign n45041 = ~n4089 & ~n45040;
  assign n45042 = n3378 & ~n45041;
  assign n45043 = ~n35228 & ~n37511;
  assign n45044 = ~controllable_hmaster1 & ~n45043;
  assign n45045 = ~n35223 & ~n45044;
  assign n45046 = i_hbusreq3 & ~n45045;
  assign n45047 = ~n18540 & ~n35234;
  assign n45048 = ~i_hbusreq2 & ~n45047;
  assign n45049 = ~n37528 & ~n45048;
  assign n45050 = ~controllable_hgrant2 & ~n45049;
  assign n45051 = ~n5862 & ~n45050;
  assign n45052 = controllable_hmaster0 & ~n45051;
  assign n45053 = ~n35258 & ~n45052;
  assign n45054 = ~controllable_hmaster1 & ~n45053;
  assign n45055 = ~n35244 & ~n45054;
  assign n45056 = ~i_hbusreq3 & ~n45055;
  assign n45057 = ~n45046 & ~n45056;
  assign n45058 = ~controllable_hmaster2 & ~n45057;
  assign n45059 = ~n39732 & ~n45058;
  assign n45060 = ~controllable_hgrant3 & ~n45059;
  assign n45061 = ~n5861 & ~n45060;
  assign n45062 = controllable_nhgrant0 & ~n45061;
  assign n45063 = ~n6082 & ~n45062;
  assign n45064 = ~n3281 & ~n45063;
  assign n45065 = ~n4089 & ~n45064;
  assign n45066 = ~n3378 & ~n45065;
  assign n45067 = ~n45042 & ~n45066;
  assign n45068 = n3492 & ~n45067;
  assign n45069 = ~n3631 & ~n45068;
  assign n45070 = n3485 & ~n45069;
  assign n45071 = ~n3630 & ~n45070;
  assign n45072 = n3476 & ~n45071;
  assign n45073 = ~n45013 & ~n45072;
  assign n45074 = n3374 & ~n45073;
  assign n45075 = ~n44971 & ~n45074;
  assign n45076 = n3655 & ~n45075;
  assign n45077 = ~n18578 & ~n34986;
  assign n45078 = ~controllable_hgrant2 & ~n45077;
  assign n45079 = ~n3410 & ~n45078;
  assign n45080 = controllable_hmaster1 & ~n45079;
  assign n45081 = controllable_hmaster0 & ~n45079;
  assign n45082 = ~n34022 & ~n45081;
  assign n45083 = ~controllable_hmaster1 & ~n45082;
  assign n45084 = ~n45080 & ~n45083;
  assign n45085 = i_hbusreq3 & ~n45084;
  assign n45086 = i_hbusreq2 & ~n45077;
  assign n45087 = ~n18601 & ~n35078;
  assign n45088 = ~i_hbusreq2 & ~n45087;
  assign n45089 = ~n45086 & ~n45088;
  assign n45090 = ~controllable_hgrant2 & ~n45089;
  assign n45091 = ~n3859 & ~n45090;
  assign n45092 = controllable_hmaster1 & ~n45091;
  assign n45093 = controllable_hmaster0 & ~n45091;
  assign n45094 = ~n34040 & ~n45093;
  assign n45095 = ~controllable_hmaster1 & ~n45094;
  assign n45096 = ~n45092 & ~n45095;
  assign n45097 = ~i_hbusreq3 & ~n45096;
  assign n45098 = ~n45085 & ~n45097;
  assign n45099 = controllable_hmaster2 & ~n45098;
  assign n45100 = ~n6188 & ~n45099;
  assign n45101 = ~controllable_hgrant3 & ~n45100;
  assign n45102 = ~n5037 & ~n45101;
  assign n45103 = controllable_nhgrant0 & ~n45102;
  assign n45104 = ~n5245 & ~n45103;
  assign n45105 = ~n3281 & ~n45104;
  assign n45106 = ~n3783 & ~n45105;
  assign n45107 = ~n3378 & ~n45106;
  assign n45108 = ~n18571 & ~n45107;
  assign n45109 = n3492 & ~n45108;
  assign n45110 = ~n3631 & ~n45109;
  assign n45111 = n3485 & ~n45110;
  assign n45112 = ~n3630 & ~n45111;
  assign n45113 = ~n3476 & ~n45112;
  assign n45114 = ~n18630 & ~n45109;
  assign n45115 = n3485 & ~n45114;
  assign n45116 = ~n18629 & ~n45115;
  assign n45117 = n3476 & ~n45116;
  assign n45118 = ~n45113 & ~n45117;
  assign n45119 = ~n3374 & ~n45118;
  assign n45120 = ~n18679 & ~n37623;
  assign n45121 = ~controllable_hmaster1 & ~n45120;
  assign n45122 = ~n18678 & ~n45121;
  assign n45123 = i_hbusreq3 & ~n45122;
  assign n45124 = ~n18695 & ~n37646;
  assign n45125 = ~controllable_hmaster1 & ~n45124;
  assign n45126 = ~n18694 & ~n45125;
  assign n45127 = ~i_hbusreq3 & ~n45126;
  assign n45128 = ~n45123 & ~n45127;
  assign n45129 = ~controllable_hmaster2 & ~n45128;
  assign n45130 = ~n18670 & ~n45129;
  assign n45131 = ~controllable_hgrant3 & ~n45130;
  assign n45132 = ~n18382 & ~n45131;
  assign n45133 = controllable_nhgrant0 & ~n45132;
  assign n45134 = ~n18416 & ~n45133;
  assign n45135 = ~n3281 & ~n45134;
  assign n45136 = ~n3950 & ~n45135;
  assign n45137 = n3378 & ~n45136;
  assign n45138 = ~n9112 & ~n34986;
  assign n45139 = ~controllable_hgrant2 & ~n45138;
  assign n45140 = ~n3410 & ~n45139;
  assign n45141 = controllable_hmaster1 & ~n45140;
  assign n45142 = controllable_hmaster0 & ~n45140;
  assign n45143 = ~n39830 & ~n45142;
  assign n45144 = ~controllable_hmaster1 & ~n45143;
  assign n45145 = ~n45141 & ~n45144;
  assign n45146 = i_hbusreq3 & ~n45145;
  assign n45147 = i_hbusreq2 & ~n45138;
  assign n45148 = ~n18721 & ~n35078;
  assign n45149 = ~i_hbusreq2 & ~n45148;
  assign n45150 = ~n45147 & ~n45149;
  assign n45151 = ~controllable_hgrant2 & ~n45150;
  assign n45152 = ~n3859 & ~n45151;
  assign n45153 = controllable_hmaster1 & ~n45152;
  assign n45154 = controllable_hmaster0 & ~n45152;
  assign n45155 = ~n39849 & ~n45154;
  assign n45156 = ~controllable_hmaster1 & ~n45155;
  assign n45157 = ~n45153 & ~n45156;
  assign n45158 = ~i_hbusreq3 & ~n45157;
  assign n45159 = ~n45146 & ~n45158;
  assign n45160 = controllable_hmaster2 & ~n45159;
  assign n45161 = ~n35369 & ~n37623;
  assign n45162 = ~controllable_hmaster1 & ~n45161;
  assign n45163 = ~n35364 & ~n45162;
  assign n45164 = i_hbusreq3 & ~n45163;
  assign n45165 = ~n35398 & ~n37646;
  assign n45166 = ~controllable_hmaster1 & ~n45165;
  assign n45167 = ~n35384 & ~n45166;
  assign n45168 = ~i_hbusreq3 & ~n45167;
  assign n45169 = ~n45164 & ~n45168;
  assign n45170 = ~controllable_hmaster2 & ~n45169;
  assign n45171 = ~n45160 & ~n45170;
  assign n45172 = ~controllable_hgrant3 & ~n45171;
  assign n45173 = ~n5402 & ~n45172;
  assign n45174 = controllable_nhgrant0 & ~n45173;
  assign n45175 = ~n5534 & ~n45174;
  assign n45176 = ~n3281 & ~n45175;
  assign n45177 = ~n3950 & ~n45176;
  assign n45178 = ~n3378 & ~n45177;
  assign n45179 = ~n45137 & ~n45178;
  assign n45180 = n3492 & ~n45179;
  assign n45181 = ~n3631 & ~n45180;
  assign n45182 = n3485 & ~n45181;
  assign n45183 = ~n3630 & ~n45182;
  assign n45184 = ~n3476 & ~n45183;
  assign n45185 = ~n9305 & ~n39673;
  assign n45186 = ~controllable_hgrant2 & ~n45185;
  assign n45187 = ~n5616 & ~n45186;
  assign n45188 = controllable_hmaster0 & ~n45187;
  assign n45189 = ~n18809 & ~n45188;
  assign n45190 = ~controllable_hmaster1 & ~n45189;
  assign n45191 = ~n18808 & ~n45190;
  assign n45192 = i_hbusreq3 & ~n45191;
  assign n45193 = i_hbusreq2 & ~n45185;
  assign n45194 = ~n17843 & ~n39683;
  assign n45195 = ~i_hbusreq2 & ~n45194;
  assign n45196 = ~n45193 & ~n45195;
  assign n45197 = ~controllable_hgrant2 & ~n45196;
  assign n45198 = ~n5657 & ~n45197;
  assign n45199 = controllable_hmaster0 & ~n45198;
  assign n45200 = ~n18831 & ~n45199;
  assign n45201 = ~controllable_hmaster1 & ~n45200;
  assign n45202 = ~n18824 & ~n45201;
  assign n45203 = ~i_hbusreq3 & ~n45202;
  assign n45204 = ~n45192 & ~n45203;
  assign n45205 = ~controllable_hmaster2 & ~n45204;
  assign n45206 = ~n18800 & ~n45205;
  assign n45207 = ~controllable_hgrant3 & ~n45206;
  assign n45208 = ~n18453 & ~n45207;
  assign n45209 = controllable_nhgrant0 & ~n45208;
  assign n45210 = ~n18526 & ~n45209;
  assign n45211 = ~n3281 & ~n45210;
  assign n45212 = ~n4089 & ~n45211;
  assign n45213 = n3378 & ~n45212;
  assign n45214 = ~n9248 & ~n35144;
  assign n45215 = ~controllable_hgrant2 & ~n45214;
  assign n45216 = ~n5616 & ~n45215;
  assign n45217 = controllable_hmaster1 & ~n45216;
  assign n45218 = controllable_hmaster0 & ~n45216;
  assign n45219 = ~n39913 & ~n45218;
  assign n45220 = ~controllable_hmaster1 & ~n45219;
  assign n45221 = ~n45217 & ~n45220;
  assign n45222 = i_hbusreq3 & ~n45221;
  assign n45223 = i_hbusreq2 & ~n45214;
  assign n45224 = ~n18855 & ~n35234;
  assign n45225 = ~i_hbusreq2 & ~n45224;
  assign n45226 = ~n45223 & ~n45225;
  assign n45227 = ~controllable_hgrant2 & ~n45226;
  assign n45228 = ~n5862 & ~n45227;
  assign n45229 = controllable_hmaster1 & ~n45228;
  assign n45230 = controllable_hmaster0 & ~n45228;
  assign n45231 = ~n39931 & ~n45230;
  assign n45232 = ~controllable_hmaster1 & ~n45231;
  assign n45233 = ~n45229 & ~n45232;
  assign n45234 = ~i_hbusreq3 & ~n45233;
  assign n45235 = ~n45222 & ~n45234;
  assign n45236 = controllable_hmaster2 & ~n45235;
  assign n45237 = ~n35494 & ~n37714;
  assign n45238 = ~controllable_hmaster1 & ~n45237;
  assign n45239 = ~n35489 & ~n45238;
  assign n45240 = i_hbusreq3 & ~n45239;
  assign n45241 = ~n18878 & ~n35234;
  assign n45242 = ~i_hbusreq2 & ~n45241;
  assign n45243 = ~n37731 & ~n45242;
  assign n45244 = ~controllable_hgrant2 & ~n45243;
  assign n45245 = ~n5862 & ~n45244;
  assign n45246 = controllable_hmaster0 & ~n45245;
  assign n45247 = ~n35522 & ~n45246;
  assign n45248 = ~controllable_hmaster1 & ~n45247;
  assign n45249 = ~n35509 & ~n45248;
  assign n45250 = ~i_hbusreq3 & ~n45249;
  assign n45251 = ~n45240 & ~n45250;
  assign n45252 = ~controllable_hmaster2 & ~n45251;
  assign n45253 = ~n45236 & ~n45252;
  assign n45254 = ~controllable_hgrant3 & ~n45253;
  assign n45255 = ~n5861 & ~n45254;
  assign n45256 = controllable_nhgrant0 & ~n45255;
  assign n45257 = ~n6082 & ~n45256;
  assign n45258 = ~n3281 & ~n45257;
  assign n45259 = ~n4089 & ~n45258;
  assign n45260 = ~n3378 & ~n45259;
  assign n45261 = ~n45213 & ~n45260;
  assign n45262 = n3492 & ~n45261;
  assign n45263 = ~n18630 & ~n45262;
  assign n45264 = n3485 & ~n45263;
  assign n45265 = ~n18629 & ~n45264;
  assign n45266 = n3476 & ~n45265;
  assign n45267 = ~n45184 & ~n45266;
  assign n45268 = n3374 & ~n45267;
  assign n45269 = ~n45119 & ~n45268;
  assign n45270 = ~n3655 & ~n45269;
  assign n45271 = ~n45076 & ~n45270;
  assign n45272 = n3652 & ~n45271;
  assign n45273 = ~n18369 & ~n39997;
  assign n45274 = n3492 & ~n45273;
  assign n45275 = ~n3631 & ~n45274;
  assign n45276 = n3485 & ~n45275;
  assign n45277 = ~n3630 & ~n45276;
  assign n45278 = ~n3374 & ~n45277;
  assign n45279 = ~n3821 & ~n37822;
  assign n45280 = ~controllable_hmaster1 & ~n45279;
  assign n45281 = ~n5293 & ~n45280;
  assign n45282 = i_hbusreq3 & ~n45281;
  assign n45283 = ~n5278 & ~n37835;
  assign n45284 = ~controllable_hmaster1 & ~n45283;
  assign n45285 = ~n5313 & ~n45284;
  assign n45286 = ~i_hbusreq3 & ~n45285;
  assign n45287 = ~n45282 & ~n45286;
  assign n45288 = ~controllable_hmaster2 & ~n45287;
  assign n45289 = ~n12065 & ~n45288;
  assign n45290 = ~controllable_hgrant3 & ~n45289;
  assign n45291 = ~n18382 & ~n45290;
  assign n45292 = controllable_nhgrant0 & ~n45291;
  assign n45293 = ~n18416 & ~n45292;
  assign n45294 = ~n3281 & ~n45293;
  assign n45295 = ~n3950 & ~n45294;
  assign n45296 = n3378 & ~n45295;
  assign n45297 = ~n35617 & ~n37822;
  assign n45298 = ~controllable_hmaster1 & ~n45297;
  assign n45299 = ~n35614 & ~n45298;
  assign n45300 = i_hbusreq3 & ~n45299;
  assign n45301 = ~n35631 & ~n37835;
  assign n45302 = ~controllable_hmaster1 & ~n45301;
  assign n45303 = ~n35627 & ~n45302;
  assign n45304 = ~i_hbusreq3 & ~n45303;
  assign n45305 = ~n45300 & ~n45304;
  assign n45306 = ~controllable_hmaster2 & ~n45305;
  assign n45307 = ~n40041 & ~n45306;
  assign n45308 = ~controllable_hgrant3 & ~n45307;
  assign n45309 = ~n5402 & ~n45308;
  assign n45310 = controllable_nhgrant0 & ~n45309;
  assign n45311 = ~n5534 & ~n45310;
  assign n45312 = ~n3281 & ~n45311;
  assign n45313 = ~n3950 & ~n45312;
  assign n45314 = ~n3378 & ~n45313;
  assign n45315 = ~n45296 & ~n45314;
  assign n45316 = n3492 & ~n45315;
  assign n45317 = ~n3631 & ~n45316;
  assign n45318 = n3485 & ~n45317;
  assign n45319 = ~n3630 & ~n45318;
  assign n45320 = ~n3476 & ~n45319;
  assign n45321 = ~n6738 & ~n45015;
  assign n45322 = controllable_hmaster0 & ~n45321;
  assign n45323 = ~n5702 & ~n45322;
  assign n45324 = ~controllable_hmaster1 & ~n45323;
  assign n45325 = ~n5690 & ~n45324;
  assign n45326 = i_hbusreq3 & ~n45325;
  assign n45327 = ~n6745 & ~n45026;
  assign n45328 = controllable_hmaster0 & ~n45327;
  assign n45329 = ~n18502 & ~n45328;
  assign n45330 = ~controllable_hmaster1 & ~n45329;
  assign n45331 = ~n18495 & ~n45330;
  assign n45332 = ~i_hbusreq3 & ~n45331;
  assign n45333 = ~n45326 & ~n45332;
  assign n45334 = ~controllable_hmaster2 & ~n45333;
  assign n45335 = ~n18481 & ~n45334;
  assign n45336 = ~controllable_hgrant3 & ~n45335;
  assign n45337 = ~n18453 & ~n45336;
  assign n45338 = controllable_nhgrant0 & ~n45337;
  assign n45339 = ~n18526 & ~n45338;
  assign n45340 = ~n3281 & ~n45339;
  assign n45341 = ~n4089 & ~n45340;
  assign n45342 = n3378 & ~n45341;
  assign n45343 = ~n35702 & ~n37884;
  assign n45344 = ~controllable_hmaster1 & ~n45343;
  assign n45345 = ~n35699 & ~n45344;
  assign n45346 = i_hbusreq3 & ~n45345;
  assign n45347 = ~n6772 & ~n45050;
  assign n45348 = controllable_hmaster0 & ~n45347;
  assign n45349 = ~n35716 & ~n45348;
  assign n45350 = ~controllable_hmaster1 & ~n45349;
  assign n45351 = ~n35712 & ~n45350;
  assign n45352 = ~i_hbusreq3 & ~n45351;
  assign n45353 = ~n45346 & ~n45352;
  assign n45354 = ~controllable_hmaster2 & ~n45353;
  assign n45355 = ~n40105 & ~n45354;
  assign n45356 = ~controllable_hgrant3 & ~n45355;
  assign n45357 = ~n5861 & ~n45356;
  assign n45358 = controllable_nhgrant0 & ~n45357;
  assign n45359 = ~n6082 & ~n45358;
  assign n45360 = ~n3281 & ~n45359;
  assign n45361 = ~n4089 & ~n45360;
  assign n45362 = ~n3378 & ~n45361;
  assign n45363 = ~n45342 & ~n45362;
  assign n45364 = n3492 & ~n45363;
  assign n45365 = ~n3631 & ~n45364;
  assign n45366 = n3485 & ~n45365;
  assign n45367 = ~n3630 & ~n45366;
  assign n45368 = n3476 & ~n45367;
  assign n45369 = ~n45320 & ~n45368;
  assign n45370 = n3374 & ~n45369;
  assign n45371 = ~n45278 & ~n45370;
  assign n45372 = n3655 & ~n45371;
  assign n45373 = ~n4333 & ~n45078;
  assign n45374 = controllable_hmaster1 & ~n45373;
  assign n45375 = controllable_hmaster0 & ~n45373;
  assign n45376 = ~n34022 & ~n45375;
  assign n45377 = ~controllable_hmaster1 & ~n45376;
  assign n45378 = ~n45374 & ~n45377;
  assign n45379 = i_hbusreq3 & ~n45378;
  assign n45380 = ~n4340 & ~n45090;
  assign n45381 = controllable_hmaster1 & ~n45380;
  assign n45382 = controllable_hmaster0 & ~n45380;
  assign n45383 = ~n34040 & ~n45382;
  assign n45384 = ~controllable_hmaster1 & ~n45383;
  assign n45385 = ~n45381 & ~n45384;
  assign n45386 = ~i_hbusreq3 & ~n45385;
  assign n45387 = ~n45379 & ~n45386;
  assign n45388 = controllable_hmaster2 & ~n45387;
  assign n45389 = ~n6887 & ~n45388;
  assign n45390 = ~controllable_hgrant3 & ~n45389;
  assign n45391 = ~n5037 & ~n45390;
  assign n45392 = controllable_nhgrant0 & ~n45391;
  assign n45393 = ~n5245 & ~n45392;
  assign n45394 = ~n3281 & ~n45393;
  assign n45395 = ~n3783 & ~n45394;
  assign n45396 = ~n3378 & ~n45395;
  assign n45397 = ~n18571 & ~n45396;
  assign n45398 = n3492 & ~n45397;
  assign n45399 = ~n3631 & ~n45398;
  assign n45400 = n3485 & ~n45399;
  assign n45401 = ~n3630 & ~n45400;
  assign n45402 = ~n3476 & ~n45401;
  assign n45403 = ~n18630 & ~n45398;
  assign n45404 = n3485 & ~n45403;
  assign n45405 = ~n18629 & ~n45404;
  assign n45406 = n3476 & ~n45405;
  assign n45407 = ~n45402 & ~n45406;
  assign n45408 = ~n3374 & ~n45407;
  assign n45409 = ~n18679 & ~n37976;
  assign n45410 = ~controllable_hmaster1 & ~n45409;
  assign n45411 = ~n18678 & ~n45410;
  assign n45412 = i_hbusreq3 & ~n45411;
  assign n45413 = ~n18695 & ~n37989;
  assign n45414 = ~controllable_hmaster1 & ~n45413;
  assign n45415 = ~n18694 & ~n45414;
  assign n45416 = ~i_hbusreq3 & ~n45415;
  assign n45417 = ~n45412 & ~n45416;
  assign n45418 = ~controllable_hmaster2 & ~n45417;
  assign n45419 = ~n18670 & ~n45418;
  assign n45420 = ~controllable_hgrant3 & ~n45419;
  assign n45421 = ~n18382 & ~n45420;
  assign n45422 = controllable_nhgrant0 & ~n45421;
  assign n45423 = ~n18416 & ~n45422;
  assign n45424 = ~n3281 & ~n45423;
  assign n45425 = ~n3950 & ~n45424;
  assign n45426 = n3378 & ~n45425;
  assign n45427 = ~n4333 & ~n45139;
  assign n45428 = controllable_hmaster1 & ~n45427;
  assign n45429 = controllable_hmaster0 & ~n45427;
  assign n45430 = ~n40188 & ~n45429;
  assign n45431 = ~controllable_hmaster1 & ~n45430;
  assign n45432 = ~n45428 & ~n45431;
  assign n45433 = i_hbusreq3 & ~n45432;
  assign n45434 = ~n4340 & ~n45151;
  assign n45435 = controllable_hmaster1 & ~n45434;
  assign n45436 = controllable_hmaster0 & ~n45434;
  assign n45437 = ~n40197 & ~n45436;
  assign n45438 = ~controllable_hmaster1 & ~n45437;
  assign n45439 = ~n45435 & ~n45438;
  assign n45440 = ~i_hbusreq3 & ~n45439;
  assign n45441 = ~n45433 & ~n45440;
  assign n45442 = controllable_hmaster2 & ~n45441;
  assign n45443 = ~n35809 & ~n37976;
  assign n45444 = ~controllable_hmaster1 & ~n45443;
  assign n45445 = ~n35806 & ~n45444;
  assign n45446 = i_hbusreq3 & ~n45445;
  assign n45447 = ~n35823 & ~n37989;
  assign n45448 = ~controllable_hmaster1 & ~n45447;
  assign n45449 = ~n35819 & ~n45448;
  assign n45450 = ~i_hbusreq3 & ~n45449;
  assign n45451 = ~n45446 & ~n45450;
  assign n45452 = ~controllable_hmaster2 & ~n45451;
  assign n45453 = ~n45442 & ~n45452;
  assign n45454 = ~controllable_hgrant3 & ~n45453;
  assign n45455 = ~n5402 & ~n45454;
  assign n45456 = controllable_nhgrant0 & ~n45455;
  assign n45457 = ~n5534 & ~n45456;
  assign n45458 = ~n3281 & ~n45457;
  assign n45459 = ~n3950 & ~n45458;
  assign n45460 = ~n3378 & ~n45459;
  assign n45461 = ~n45426 & ~n45460;
  assign n45462 = n3492 & ~n45461;
  assign n45463 = ~n3631 & ~n45462;
  assign n45464 = n3485 & ~n45463;
  assign n45465 = ~n3630 & ~n45464;
  assign n45466 = ~n3476 & ~n45465;
  assign n45467 = ~n6738 & ~n45186;
  assign n45468 = controllable_hmaster0 & ~n45467;
  assign n45469 = ~n18809 & ~n45468;
  assign n45470 = ~controllable_hmaster1 & ~n45469;
  assign n45471 = ~n18808 & ~n45470;
  assign n45472 = i_hbusreq3 & ~n45471;
  assign n45473 = ~n6745 & ~n45197;
  assign n45474 = controllable_hmaster0 & ~n45473;
  assign n45475 = ~n18831 & ~n45474;
  assign n45476 = ~controllable_hmaster1 & ~n45475;
  assign n45477 = ~n18824 & ~n45476;
  assign n45478 = ~i_hbusreq3 & ~n45477;
  assign n45479 = ~n45472 & ~n45478;
  assign n45480 = ~controllable_hmaster2 & ~n45479;
  assign n45481 = ~n18800 & ~n45480;
  assign n45482 = ~controllable_hgrant3 & ~n45481;
  assign n45483 = ~n18453 & ~n45482;
  assign n45484 = controllable_nhgrant0 & ~n45483;
  assign n45485 = ~n18526 & ~n45484;
  assign n45486 = ~n3281 & ~n45485;
  assign n45487 = ~n4089 & ~n45486;
  assign n45488 = n3378 & ~n45487;
  assign n45489 = ~n6762 & ~n45215;
  assign n45490 = controllable_hmaster1 & ~n45489;
  assign n45491 = controllable_hmaster0 & ~n45489;
  assign n45492 = ~n40252 & ~n45491;
  assign n45493 = ~controllable_hmaster1 & ~n45492;
  assign n45494 = ~n45490 & ~n45493;
  assign n45495 = i_hbusreq3 & ~n45494;
  assign n45496 = ~n6772 & ~n45227;
  assign n45497 = controllable_hmaster1 & ~n45496;
  assign n45498 = controllable_hmaster0 & ~n45496;
  assign n45499 = ~n40261 & ~n45498;
  assign n45500 = ~controllable_hmaster1 & ~n45499;
  assign n45501 = ~n45497 & ~n45500;
  assign n45502 = ~i_hbusreq3 & ~n45501;
  assign n45503 = ~n45495 & ~n45502;
  assign n45504 = controllable_hmaster2 & ~n45503;
  assign n45505 = ~n35894 & ~n38038;
  assign n45506 = ~controllable_hmaster1 & ~n45505;
  assign n45507 = ~n35891 & ~n45506;
  assign n45508 = i_hbusreq3 & ~n45507;
  assign n45509 = ~n6772 & ~n45244;
  assign n45510 = controllable_hmaster0 & ~n45509;
  assign n45511 = ~n35908 & ~n45510;
  assign n45512 = ~controllable_hmaster1 & ~n45511;
  assign n45513 = ~n35904 & ~n45512;
  assign n45514 = ~i_hbusreq3 & ~n45513;
  assign n45515 = ~n45508 & ~n45514;
  assign n45516 = ~controllable_hmaster2 & ~n45515;
  assign n45517 = ~n45504 & ~n45516;
  assign n45518 = ~controllable_hgrant3 & ~n45517;
  assign n45519 = ~n5861 & ~n45518;
  assign n45520 = controllable_nhgrant0 & ~n45519;
  assign n45521 = ~n6082 & ~n45520;
  assign n45522 = ~n3281 & ~n45521;
  assign n45523 = ~n4089 & ~n45522;
  assign n45524 = ~n3378 & ~n45523;
  assign n45525 = ~n45488 & ~n45524;
  assign n45526 = n3492 & ~n45525;
  assign n45527 = ~n18630 & ~n45526;
  assign n45528 = n3485 & ~n45527;
  assign n45529 = ~n18629 & ~n45528;
  assign n45530 = n3476 & ~n45529;
  assign n45531 = ~n45466 & ~n45530;
  assign n45532 = n3374 & ~n45531;
  assign n45533 = ~n45408 & ~n45532;
  assign n45534 = ~n3655 & ~n45533;
  assign n45535 = ~n45372 & ~n45534;
  assign n45536 = ~n3652 & ~n45535;
  assign n45537 = ~n45272 & ~n45536;
  assign n45538 = ~n3368 & ~n45537;
  assign n45539 = ~n3821 & ~n38149;
  assign n45540 = ~controllable_hmaster1 & ~n45539;
  assign n45541 = ~n5293 & ~n45540;
  assign n45542 = i_hbusreq3 & ~n45541;
  assign n45543 = ~n5278 & ~n38172;
  assign n45544 = ~controllable_hmaster1 & ~n45543;
  assign n45545 = ~n5313 & ~n45544;
  assign n45546 = ~i_hbusreq3 & ~n45545;
  assign n45547 = ~n45542 & ~n45546;
  assign n45548 = ~controllable_hmaster2 & ~n45547;
  assign n45549 = ~n12741 & ~n45548;
  assign n45550 = ~controllable_hgrant3 & ~n45549;
  assign n45551 = ~n19183 & ~n45550;
  assign n45552 = controllable_nhgrant0 & ~n45551;
  assign n45553 = ~n19213 & ~n45552;
  assign n45554 = ~n3281 & ~n45553;
  assign n45555 = ~n3281 & ~n45554;
  assign n45556 = n3378 & ~n45555;
  assign n45557 = ~n35062 & ~n38149;
  assign n45558 = ~controllable_hmaster1 & ~n45557;
  assign n45559 = ~n35057 & ~n45558;
  assign n45560 = i_hbusreq3 & ~n45559;
  assign n45561 = ~n35089 & ~n38172;
  assign n45562 = ~controllable_hmaster1 & ~n45561;
  assign n45563 = ~n35076 & ~n45562;
  assign n45564 = ~i_hbusreq3 & ~n45563;
  assign n45565 = ~n45560 & ~n45564;
  assign n45566 = ~controllable_hmaster2 & ~n45565;
  assign n45567 = ~n40353 & ~n45566;
  assign n45568 = ~controllable_hgrant3 & ~n45567;
  assign n45569 = ~n19225 & ~n45568;
  assign n45570 = controllable_nhgrant0 & ~n45569;
  assign n45571 = ~n19255 & ~n45570;
  assign n45572 = ~n3281 & ~n45571;
  assign n45573 = ~n3281 & ~n45572;
  assign n45574 = ~n3378 & ~n45573;
  assign n45575 = ~n45556 & ~n45574;
  assign n45576 = n3492 & ~n45575;
  assign n45577 = n3492 & ~n45576;
  assign n45578 = n3485 & ~n45577;
  assign n45579 = n3485 & ~n45578;
  assign n45580 = ~n3476 & ~n45579;
  assign n45581 = ~n19315 & ~n40378;
  assign n45582 = ~controllable_hgrant2 & ~n45581;
  assign n45583 = ~n5616 & ~n45582;
  assign n45584 = controllable_hmaster0 & ~n45583;
  assign n45585 = ~n7340 & ~n45584;
  assign n45586 = ~controllable_hmaster1 & ~n45585;
  assign n45587 = ~n7330 & ~n45586;
  assign n45588 = i_hbusreq3 & ~n45587;
  assign n45589 = i_hbusreq2 & ~n45581;
  assign n45590 = ~n19354 & ~n40388;
  assign n45591 = ~i_hbusreq2 & ~n45590;
  assign n45592 = ~n45589 & ~n45591;
  assign n45593 = ~controllable_hgrant2 & ~n45592;
  assign n45594 = ~n7290 & ~n45593;
  assign n45595 = controllable_hmaster0 & ~n45594;
  assign n45596 = ~n19361 & ~n45595;
  assign n45597 = ~controllable_hmaster1 & ~n45596;
  assign n45598 = ~n19333 & ~n45597;
  assign n45599 = ~i_hbusreq3 & ~n45598;
  assign n45600 = ~n45588 & ~n45599;
  assign n45601 = ~controllable_hmaster2 & ~n45600;
  assign n45602 = ~n19313 & ~n45601;
  assign n45603 = ~controllable_hgrant3 & ~n45602;
  assign n45604 = ~n19274 & ~n45603;
  assign n45605 = controllable_nhgrant0 & ~n45604;
  assign n45606 = ~n19385 & ~n45605;
  assign n45607 = ~n3281 & ~n45606;
  assign n45608 = ~n3281 & ~n45607;
  assign n45609 = n3378 & ~n45608;
  assign n45610 = ~n19408 & ~n35234;
  assign n45611 = ~i_hbusreq2 & ~n45610;
  assign n45612 = ~n40422 & ~n45611;
  assign n45613 = ~controllable_hgrant2 & ~n45612;
  assign n45614 = ~n5862 & ~n45613;
  assign n45615 = controllable_hmaster1 & ~n45614;
  assign n45616 = controllable_hmaster0 & ~n45614;
  assign n45617 = ~n19425 & ~n34214;
  assign n45618 = ~i_hbusreq2 & ~n45617;
  assign n45619 = ~n40430 & ~n45618;
  assign n45620 = ~controllable_hgrant2 & ~n45619;
  assign n45621 = ~n5862 & ~n45620;
  assign n45622 = ~controllable_hmaster0 & ~n45621;
  assign n45623 = ~n45616 & ~n45622;
  assign n45624 = ~controllable_hmaster1 & ~n45623;
  assign n45625 = ~n45615 & ~n45624;
  assign n45626 = ~i_hbusreq3 & ~n45625;
  assign n45627 = ~n40421 & ~n45626;
  assign n45628 = controllable_hmaster2 & ~n45627;
  assign n45629 = ~n40451 & ~n43149;
  assign n45630 = controllable_hmaster1 & ~n45629;
  assign n45631 = ~n19439 & ~n40443;
  assign n45632 = ~controllable_hgrant2 & ~n45631;
  assign n45633 = ~n5616 & ~n45632;
  assign n45634 = controllable_hmaster0 & ~n45633;
  assign n45635 = ~n40459 & ~n45634;
  assign n45636 = ~controllable_hmaster1 & ~n45635;
  assign n45637 = ~n45630 & ~n45636;
  assign n45638 = i_hbusreq3 & ~n45637;
  assign n45639 = ~n19425 & ~n35234;
  assign n45640 = ~i_hbusreq2 & ~n45639;
  assign n45641 = ~n40472 & ~n45640;
  assign n45642 = ~controllable_hgrant2 & ~n45641;
  assign n45643 = ~n5862 & ~n45642;
  assign n45644 = controllable_hmaster0 & ~n45643;
  assign n45645 = ~n5950 & ~n45642;
  assign n45646 = ~controllable_hmaster0 & ~n45645;
  assign n45647 = ~n45644 & ~n45646;
  assign n45648 = controllable_hmaster1 & ~n45647;
  assign n45649 = i_hbusreq2 & ~n45631;
  assign n45650 = ~n19471 & ~n40465;
  assign n45651 = ~i_hbusreq2 & ~n45650;
  assign n45652 = ~n45649 & ~n45651;
  assign n45653 = ~controllable_hgrant2 & ~n45652;
  assign n45654 = ~n7507 & ~n45653;
  assign n45655 = controllable_hmaster0 & ~n45654;
  assign n45656 = ~n19485 & ~n35252;
  assign n45657 = ~i_hbusreq2 & ~n45656;
  assign n45658 = ~n40472 & ~n45657;
  assign n45659 = ~controllable_hgrant2 & ~n45658;
  assign n45660 = ~n5981 & ~n45659;
  assign n45661 = ~controllable_hmaster0 & ~n45660;
  assign n45662 = ~n45655 & ~n45661;
  assign n45663 = ~controllable_hmaster1 & ~n45662;
  assign n45664 = ~n45648 & ~n45663;
  assign n45665 = ~i_hbusreq3 & ~n45664;
  assign n45666 = ~n45638 & ~n45665;
  assign n45667 = ~controllable_hmaster2 & ~n45666;
  assign n45668 = ~n45628 & ~n45667;
  assign n45669 = ~controllable_hgrant3 & ~n45668;
  assign n45670 = ~n19398 & ~n45669;
  assign n45671 = controllable_nhgrant0 & ~n45670;
  assign n45672 = ~n19515 & ~n45671;
  assign n45673 = ~n3281 & ~n45672;
  assign n45674 = ~n3281 & ~n45673;
  assign n45675 = ~n3378 & ~n45674;
  assign n45676 = ~n45609 & ~n45675;
  assign n45677 = n3492 & ~n45676;
  assign n45678 = n3492 & ~n45677;
  assign n45679 = n3485 & ~n45678;
  assign n45680 = n3485 & ~n45679;
  assign n45681 = n3476 & ~n45680;
  assign n45682 = ~n45580 & ~n45681;
  assign n45683 = n3374 & ~n45682;
  assign n45684 = ~n40325 & ~n45683;
  assign n45685 = n3655 & ~n45684;
  assign n45686 = ~n19580 & ~n34986;
  assign n45687 = ~controllable_hgrant2 & ~n45686;
  assign n45688 = ~n3410 & ~n45687;
  assign n45689 = controllable_hmaster1 & ~n45688;
  assign n45690 = controllable_hmaster0 & ~n45688;
  assign n45691 = controllable_hmaster0 & ~n45690;
  assign n45692 = ~controllable_hmaster1 & ~n45691;
  assign n45693 = ~n45689 & ~n45692;
  assign n45694 = i_hbusreq3 & ~n45693;
  assign n45695 = i_hbusreq2 & ~n45686;
  assign n45696 = ~n19603 & ~n35078;
  assign n45697 = ~i_hbusreq2 & ~n45696;
  assign n45698 = ~n45695 & ~n45697;
  assign n45699 = ~controllable_hgrant2 & ~n45698;
  assign n45700 = ~n3859 & ~n45699;
  assign n45701 = controllable_hmaster1 & ~n45700;
  assign n45702 = controllable_hmaster0 & ~n45700;
  assign n45703 = controllable_hmaster0 & ~n45702;
  assign n45704 = ~controllable_hmaster1 & ~n45703;
  assign n45705 = ~n45701 & ~n45704;
  assign n45706 = ~i_hbusreq3 & ~n45705;
  assign n45707 = ~n45694 & ~n45706;
  assign n45708 = controllable_hmaster2 & ~n45707;
  assign n45709 = controllable_hmaster2 & ~n45708;
  assign n45710 = ~controllable_hgrant3 & ~n45709;
  assign n45711 = ~n7090 & ~n45710;
  assign n45712 = controllable_nhgrant0 & ~n45711;
  assign n45713 = ~n7118 & ~n45712;
  assign n45714 = ~n3281 & ~n45713;
  assign n45715 = ~n3281 & ~n45714;
  assign n45716 = ~n3378 & ~n45715;
  assign n45717 = ~n19575 & ~n45716;
  assign n45718 = n3492 & ~n45717;
  assign n45719 = n3492 & ~n45718;
  assign n45720 = n3485 & ~n45719;
  assign n45721 = n3485 & ~n45720;
  assign n45722 = ~n3374 & ~n45721;
  assign n45723 = ~n19670 & ~n38448;
  assign n45724 = ~controllable_hmaster1 & ~n45723;
  assign n45725 = ~n19669 & ~n45724;
  assign n45726 = i_hbusreq3 & ~n45725;
  assign n45727 = ~n19686 & ~n38471;
  assign n45728 = ~controllable_hmaster1 & ~n45727;
  assign n45729 = ~n19685 & ~n45728;
  assign n45730 = ~i_hbusreq3 & ~n45729;
  assign n45731 = ~n45726 & ~n45730;
  assign n45732 = ~controllable_hmaster2 & ~n45731;
  assign n45733 = ~n19661 & ~n45732;
  assign n45734 = ~controllable_hgrant3 & ~n45733;
  assign n45735 = ~n19183 & ~n45734;
  assign n45736 = controllable_nhgrant0 & ~n45735;
  assign n45737 = ~n19213 & ~n45736;
  assign n45738 = ~n3281 & ~n45737;
  assign n45739 = ~n3281 & ~n45738;
  assign n45740 = n3378 & ~n45739;
  assign n45741 = ~n19705 & ~n34121;
  assign n45742 = ~controllable_hgrant2 & ~n45741;
  assign n45743 = ~n3410 & ~n45742;
  assign n45744 = ~controllable_hmaster0 & ~n45743;
  assign n45745 = ~n45690 & ~n45744;
  assign n45746 = ~controllable_hmaster1 & ~n45745;
  assign n45747 = ~n45689 & ~n45746;
  assign n45748 = i_hbusreq3 & ~n45747;
  assign n45749 = i_hbusreq2 & ~n45741;
  assign n45750 = ~n19727 & ~n34131;
  assign n45751 = ~i_hbusreq2 & ~n45750;
  assign n45752 = ~n45749 & ~n45751;
  assign n45753 = ~controllable_hgrant2 & ~n45752;
  assign n45754 = ~n3859 & ~n45753;
  assign n45755 = ~controllable_hmaster0 & ~n45754;
  assign n45756 = ~n45702 & ~n45755;
  assign n45757 = ~controllable_hmaster1 & ~n45756;
  assign n45758 = ~n45701 & ~n45757;
  assign n45759 = ~i_hbusreq3 & ~n45758;
  assign n45760 = ~n45748 & ~n45759;
  assign n45761 = controllable_hmaster2 & ~n45760;
  assign n45762 = ~n19705 & ~n34986;
  assign n45763 = ~controllable_hgrant2 & ~n45762;
  assign n45764 = ~n3410 & ~n45763;
  assign n45765 = controllable_hmaster0 & ~n45764;
  assign n45766 = ~n5288 & ~n45763;
  assign n45767 = ~controllable_hmaster0 & ~n45766;
  assign n45768 = ~n45765 & ~n45767;
  assign n45769 = controllable_hmaster1 & ~n45768;
  assign n45770 = ~controllable_hmaster0 & ~n45764;
  assign n45771 = ~n38448 & ~n45770;
  assign n45772 = ~controllable_hmaster1 & ~n45771;
  assign n45773 = ~n45769 & ~n45772;
  assign n45774 = i_hbusreq3 & ~n45773;
  assign n45775 = i_hbusreq2 & ~n45762;
  assign n45776 = ~n19727 & ~n35078;
  assign n45777 = ~i_hbusreq2 & ~n45776;
  assign n45778 = ~n45775 & ~n45777;
  assign n45779 = ~controllable_hgrant2 & ~n45778;
  assign n45780 = ~n3859 & ~n45779;
  assign n45781 = controllable_hmaster0 & ~n45780;
  assign n45782 = ~n5438 & ~n45779;
  assign n45783 = ~controllable_hmaster0 & ~n45782;
  assign n45784 = ~n45781 & ~n45783;
  assign n45785 = controllable_hmaster1 & ~n45784;
  assign n45786 = ~n19773 & ~n35392;
  assign n45787 = ~i_hbusreq2 & ~n45786;
  assign n45788 = ~n45775 & ~n45787;
  assign n45789 = ~controllable_hgrant2 & ~n45788;
  assign n45790 = ~n5461 & ~n45789;
  assign n45791 = ~controllable_hmaster0 & ~n45790;
  assign n45792 = ~n38471 & ~n45791;
  assign n45793 = ~controllable_hmaster1 & ~n45792;
  assign n45794 = ~n45785 & ~n45793;
  assign n45795 = ~i_hbusreq3 & ~n45794;
  assign n45796 = ~n45774 & ~n45795;
  assign n45797 = ~controllable_hmaster2 & ~n45796;
  assign n45798 = ~n45761 & ~n45797;
  assign n45799 = ~controllable_hgrant3 & ~n45798;
  assign n45800 = ~n19225 & ~n45799;
  assign n45801 = controllable_nhgrant0 & ~n45800;
  assign n45802 = ~n19255 & ~n45801;
  assign n45803 = ~n3281 & ~n45802;
  assign n45804 = ~n3281 & ~n45803;
  assign n45805 = ~n3378 & ~n45804;
  assign n45806 = ~n45740 & ~n45805;
  assign n45807 = n3492 & ~n45806;
  assign n45808 = n3492 & ~n45807;
  assign n45809 = n3485 & ~n45808;
  assign n45810 = n3485 & ~n45809;
  assign n45811 = ~n3476 & ~n45810;
  assign n45812 = ~n19892 & ~n40378;
  assign n45813 = ~controllable_hgrant2 & ~n45812;
  assign n45814 = ~n5616 & ~n45813;
  assign n45815 = controllable_hmaster0 & ~n45814;
  assign n45816 = ~n19897 & ~n45815;
  assign n45817 = ~controllable_hmaster1 & ~n45816;
  assign n45818 = ~n19885 & ~n45817;
  assign n45819 = i_hbusreq3 & ~n45818;
  assign n45820 = i_hbusreq2 & ~n45812;
  assign n45821 = ~n19934 & ~n40388;
  assign n45822 = ~i_hbusreq2 & ~n45821;
  assign n45823 = ~n45820 & ~n45822;
  assign n45824 = ~controllable_hgrant2 & ~n45823;
  assign n45825 = ~n7290 & ~n45824;
  assign n45826 = controllable_hmaster0 & ~n45825;
  assign n45827 = ~n19941 & ~n45826;
  assign n45828 = ~controllable_hmaster1 & ~n45827;
  assign n45829 = ~n19912 & ~n45828;
  assign n45830 = ~i_hbusreq3 & ~n45829;
  assign n45831 = ~n45819 & ~n45830;
  assign n45832 = ~controllable_hmaster2 & ~n45831;
  assign n45833 = ~n19877 & ~n45832;
  assign n45834 = ~controllable_hgrant3 & ~n45833;
  assign n45835 = ~n19274 & ~n45834;
  assign n45836 = controllable_nhgrant0 & ~n45835;
  assign n45837 = ~n19385 & ~n45836;
  assign n45838 = ~n3281 & ~n45837;
  assign n45839 = ~n3281 & ~n45838;
  assign n45840 = n3378 & ~n45839;
  assign n45841 = ~n19960 & ~n35144;
  assign n45842 = ~controllable_hgrant2 & ~n45841;
  assign n45843 = ~n5616 & ~n45842;
  assign n45844 = controllable_hmaster1 & ~n45843;
  assign n45845 = controllable_hmaster0 & ~n45843;
  assign n45846 = ~n19971 & ~n34195;
  assign n45847 = ~controllable_hgrant2 & ~n45846;
  assign n45848 = ~n5616 & ~n45847;
  assign n45849 = ~controllable_hmaster0 & ~n45848;
  assign n45850 = ~n45845 & ~n45849;
  assign n45851 = ~controllable_hmaster1 & ~n45850;
  assign n45852 = ~n45844 & ~n45851;
  assign n45853 = i_hbusreq3 & ~n45852;
  assign n45854 = i_hbusreq2 & ~n45841;
  assign n45855 = ~n19999 & ~n35234;
  assign n45856 = ~i_hbusreq2 & ~n45855;
  assign n45857 = ~n45854 & ~n45856;
  assign n45858 = ~controllable_hgrant2 & ~n45857;
  assign n45859 = ~n5862 & ~n45858;
  assign n45860 = controllable_hmaster1 & ~n45859;
  assign n45861 = controllable_hmaster0 & ~n45859;
  assign n45862 = i_hbusreq2 & ~n45846;
  assign n45863 = ~n20026 & ~n34214;
  assign n45864 = ~i_hbusreq2 & ~n45863;
  assign n45865 = ~n45862 & ~n45864;
  assign n45866 = ~controllable_hgrant2 & ~n45865;
  assign n45867 = ~n5862 & ~n45866;
  assign n45868 = ~controllable_hmaster0 & ~n45867;
  assign n45869 = ~n45861 & ~n45868;
  assign n45870 = ~controllable_hmaster1 & ~n45869;
  assign n45871 = ~n45860 & ~n45870;
  assign n45872 = ~i_hbusreq3 & ~n45871;
  assign n45873 = ~n45853 & ~n45872;
  assign n45874 = controllable_hmaster2 & ~n45873;
  assign n45875 = ~n19971 & ~n35144;
  assign n45876 = ~controllable_hgrant2 & ~n45875;
  assign n45877 = ~n5616 & ~n45876;
  assign n45878 = controllable_hmaster0 & ~n45877;
  assign n45879 = ~n5686 & ~n45876;
  assign n45880 = ~controllable_hmaster0 & ~n45879;
  assign n45881 = ~n45878 & ~n45880;
  assign n45882 = controllable_hmaster1 & ~n45881;
  assign n45883 = ~n20050 & ~n40443;
  assign n45884 = ~controllable_hgrant2 & ~n45883;
  assign n45885 = ~n5616 & ~n45884;
  assign n45886 = controllable_hmaster0 & ~n45885;
  assign n45887 = ~controllable_hmaster0 & ~n45877;
  assign n45888 = ~n45886 & ~n45887;
  assign n45889 = ~controllable_hmaster1 & ~n45888;
  assign n45890 = ~n45882 & ~n45889;
  assign n45891 = i_hbusreq3 & ~n45890;
  assign n45892 = i_hbusreq2 & ~n45875;
  assign n45893 = ~n20026 & ~n35234;
  assign n45894 = ~i_hbusreq2 & ~n45893;
  assign n45895 = ~n45892 & ~n45894;
  assign n45896 = ~controllable_hgrant2 & ~n45895;
  assign n45897 = ~n5862 & ~n45896;
  assign n45898 = controllable_hmaster0 & ~n45897;
  assign n45899 = ~n5950 & ~n45896;
  assign n45900 = ~controllable_hmaster0 & ~n45899;
  assign n45901 = ~n45898 & ~n45900;
  assign n45902 = controllable_hmaster1 & ~n45901;
  assign n45903 = i_hbusreq2 & ~n45883;
  assign n45904 = ~n20089 & ~n40465;
  assign n45905 = ~i_hbusreq2 & ~n45904;
  assign n45906 = ~n45903 & ~n45905;
  assign n45907 = ~controllable_hgrant2 & ~n45906;
  assign n45908 = ~n7507 & ~n45907;
  assign n45909 = controllable_hmaster0 & ~n45908;
  assign n45910 = ~n20104 & ~n35252;
  assign n45911 = ~i_hbusreq2 & ~n45910;
  assign n45912 = ~n45892 & ~n45911;
  assign n45913 = ~controllable_hgrant2 & ~n45912;
  assign n45914 = ~n5981 & ~n45913;
  assign n45915 = ~controllable_hmaster0 & ~n45914;
  assign n45916 = ~n45909 & ~n45915;
  assign n45917 = ~controllable_hmaster1 & ~n45916;
  assign n45918 = ~n45902 & ~n45917;
  assign n45919 = ~i_hbusreq3 & ~n45918;
  assign n45920 = ~n45891 & ~n45919;
  assign n45921 = ~controllable_hmaster2 & ~n45920;
  assign n45922 = ~n45874 & ~n45921;
  assign n45923 = ~controllable_hgrant3 & ~n45922;
  assign n45924 = ~n19398 & ~n45923;
  assign n45925 = controllable_nhgrant0 & ~n45924;
  assign n45926 = ~n19515 & ~n45925;
  assign n45927 = ~n3281 & ~n45926;
  assign n45928 = ~n3281 & ~n45927;
  assign n45929 = ~n3378 & ~n45928;
  assign n45930 = ~n45840 & ~n45929;
  assign n45931 = n3492 & ~n45930;
  assign n45932 = ~n18151 & ~n45931;
  assign n45933 = n3485 & ~n45932;
  assign n45934 = ~n18150 & ~n45933;
  assign n45935 = n3476 & ~n45934;
  assign n45936 = ~n45811 & ~n45935;
  assign n45937 = n3374 & ~n45936;
  assign n45938 = ~n45722 & ~n45937;
  assign n45939 = ~n3655 & ~n45938;
  assign n45940 = ~n45685 & ~n45939;
  assign n45941 = n3652 & ~n45940;
  assign n45942 = ~n3821 & ~n38727;
  assign n45943 = ~controllable_hmaster1 & ~n45942;
  assign n45944 = ~n5293 & ~n45943;
  assign n45945 = i_hbusreq3 & ~n45944;
  assign n45946 = ~n5278 & ~n38740;
  assign n45947 = ~controllable_hmaster1 & ~n45946;
  assign n45948 = ~n5313 & ~n45947;
  assign n45949 = ~i_hbusreq3 & ~n45948;
  assign n45950 = ~n45945 & ~n45949;
  assign n45951 = ~controllable_hmaster2 & ~n45950;
  assign n45952 = ~n12741 & ~n45951;
  assign n45953 = ~controllable_hgrant3 & ~n45952;
  assign n45954 = ~n19183 & ~n45953;
  assign n45955 = controllable_nhgrant0 & ~n45954;
  assign n45956 = ~n19213 & ~n45955;
  assign n45957 = ~n3281 & ~n45956;
  assign n45958 = ~n3281 & ~n45957;
  assign n45959 = n3378 & ~n45958;
  assign n45960 = ~n35617 & ~n38727;
  assign n45961 = ~controllable_hmaster1 & ~n45960;
  assign n45962 = ~n35614 & ~n45961;
  assign n45963 = i_hbusreq3 & ~n45962;
  assign n45964 = ~n35631 & ~n38740;
  assign n45965 = ~controllable_hmaster1 & ~n45964;
  assign n45966 = ~n35627 & ~n45965;
  assign n45967 = ~i_hbusreq3 & ~n45966;
  assign n45968 = ~n45963 & ~n45967;
  assign n45969 = ~controllable_hmaster2 & ~n45968;
  assign n45970 = ~n40783 & ~n45969;
  assign n45971 = ~controllable_hgrant3 & ~n45970;
  assign n45972 = ~n19225 & ~n45971;
  assign n45973 = controllable_nhgrant0 & ~n45972;
  assign n45974 = ~n19255 & ~n45973;
  assign n45975 = ~n3281 & ~n45974;
  assign n45976 = ~n3281 & ~n45975;
  assign n45977 = ~n3378 & ~n45976;
  assign n45978 = ~n45959 & ~n45977;
  assign n45979 = n3492 & ~n45978;
  assign n45980 = n3492 & ~n45979;
  assign n45981 = n3485 & ~n45980;
  assign n45982 = n3485 & ~n45981;
  assign n45983 = ~n3476 & ~n45982;
  assign n45984 = ~n8029 & ~n45582;
  assign n45985 = controllable_hmaster0 & ~n45984;
  assign n45986 = ~n7340 & ~n45985;
  assign n45987 = ~controllable_hmaster1 & ~n45986;
  assign n45988 = ~n7330 & ~n45987;
  assign n45989 = i_hbusreq3 & ~n45988;
  assign n45990 = ~n8036 & ~n45593;
  assign n45991 = controllable_hmaster0 & ~n45990;
  assign n45992 = ~n19361 & ~n45991;
  assign n45993 = ~controllable_hmaster1 & ~n45992;
  assign n45994 = ~n19333 & ~n45993;
  assign n45995 = ~i_hbusreq3 & ~n45994;
  assign n45996 = ~n45989 & ~n45995;
  assign n45997 = ~controllable_hmaster2 & ~n45996;
  assign n45998 = ~n19313 & ~n45997;
  assign n45999 = ~controllable_hgrant3 & ~n45998;
  assign n46000 = ~n19274 & ~n45999;
  assign n46001 = controllable_nhgrant0 & ~n46000;
  assign n46002 = ~n19385 & ~n46001;
  assign n46003 = ~n3281 & ~n46002;
  assign n46004 = ~n3281 & ~n46003;
  assign n46005 = n3378 & ~n46004;
  assign n46006 = ~n6772 & ~n45613;
  assign n46007 = controllable_hmaster1 & ~n46006;
  assign n46008 = controllable_hmaster0 & ~n46006;
  assign n46009 = ~n6772 & ~n45620;
  assign n46010 = ~controllable_hmaster0 & ~n46009;
  assign n46011 = ~n46008 & ~n46010;
  assign n46012 = ~controllable_hmaster1 & ~n46011;
  assign n46013 = ~n46007 & ~n46012;
  assign n46014 = ~i_hbusreq3 & ~n46013;
  assign n46015 = ~n40838 & ~n46014;
  assign n46016 = controllable_hmaster2 & ~n46015;
  assign n46017 = controllable_hmaster0 & ~n40858;
  assign n46018 = ~n40853 & ~n46017;
  assign n46019 = controllable_hmaster1 & ~n46018;
  assign n46020 = ~n8056 & ~n45632;
  assign n46021 = controllable_hmaster0 & ~n46020;
  assign n46022 = ~n40859 & ~n46021;
  assign n46023 = ~controllable_hmaster1 & ~n46022;
  assign n46024 = ~n46019 & ~n46023;
  assign n46025 = i_hbusreq3 & ~n46024;
  assign n46026 = ~n6772 & ~n45642;
  assign n46027 = controllable_hmaster0 & ~n46026;
  assign n46028 = ~n6813 & ~n45642;
  assign n46029 = ~controllable_hmaster0 & ~n46028;
  assign n46030 = ~n46027 & ~n46029;
  assign n46031 = controllable_hmaster1 & ~n46030;
  assign n46032 = ~n8066 & ~n45653;
  assign n46033 = controllable_hmaster0 & ~n46032;
  assign n46034 = ~n6831 & ~n45659;
  assign n46035 = ~controllable_hmaster0 & ~n46034;
  assign n46036 = ~n46033 & ~n46035;
  assign n46037 = ~controllable_hmaster1 & ~n46036;
  assign n46038 = ~n46031 & ~n46037;
  assign n46039 = ~i_hbusreq3 & ~n46038;
  assign n46040 = ~n46025 & ~n46039;
  assign n46041 = ~controllable_hmaster2 & ~n46040;
  assign n46042 = ~n46016 & ~n46041;
  assign n46043 = ~controllable_hgrant3 & ~n46042;
  assign n46044 = ~n19398 & ~n46043;
  assign n46045 = controllable_nhgrant0 & ~n46044;
  assign n46046 = ~n19515 & ~n46045;
  assign n46047 = ~n3281 & ~n46046;
  assign n46048 = ~n3281 & ~n46047;
  assign n46049 = ~n3378 & ~n46048;
  assign n46050 = ~n46005 & ~n46049;
  assign n46051 = n3492 & ~n46050;
  assign n46052 = n3492 & ~n46051;
  assign n46053 = n3485 & ~n46052;
  assign n46054 = n3485 & ~n46053;
  assign n46055 = n3476 & ~n46054;
  assign n46056 = ~n45983 & ~n46055;
  assign n46057 = n3374 & ~n46056;
  assign n46058 = ~n40755 & ~n46057;
  assign n46059 = n3655 & ~n46058;
  assign n46060 = ~n4333 & ~n45687;
  assign n46061 = controllable_hmaster1 & ~n46060;
  assign n46062 = controllable_hmaster0 & ~n46060;
  assign n46063 = controllable_hmaster0 & ~n46062;
  assign n46064 = ~controllable_hmaster1 & ~n46063;
  assign n46065 = ~n46061 & ~n46064;
  assign n46066 = i_hbusreq3 & ~n46065;
  assign n46067 = ~n4340 & ~n45699;
  assign n46068 = controllable_hmaster1 & ~n46067;
  assign n46069 = controllable_hmaster0 & ~n46067;
  assign n46070 = controllable_hmaster0 & ~n46069;
  assign n46071 = ~controllable_hmaster1 & ~n46070;
  assign n46072 = ~n46068 & ~n46071;
  assign n46073 = ~i_hbusreq3 & ~n46072;
  assign n46074 = ~n46066 & ~n46073;
  assign n46075 = controllable_hmaster2 & ~n46074;
  assign n46076 = controllable_hmaster2 & ~n46075;
  assign n46077 = ~controllable_hgrant3 & ~n46076;
  assign n46078 = ~n7090 & ~n46077;
  assign n46079 = controllable_nhgrant0 & ~n46078;
  assign n46080 = ~n7118 & ~n46079;
  assign n46081 = ~n3281 & ~n46080;
  assign n46082 = ~n3281 & ~n46081;
  assign n46083 = ~n3378 & ~n46082;
  assign n46084 = ~n19575 & ~n46083;
  assign n46085 = n3492 & ~n46084;
  assign n46086 = n3492 & ~n46085;
  assign n46087 = n3485 & ~n46086;
  assign n46088 = n3485 & ~n46087;
  assign n46089 = ~n3374 & ~n46088;
  assign n46090 = ~n19670 & ~n38936;
  assign n46091 = ~controllable_hmaster1 & ~n46090;
  assign n46092 = ~n19669 & ~n46091;
  assign n46093 = i_hbusreq3 & ~n46092;
  assign n46094 = ~n19686 & ~n38949;
  assign n46095 = ~controllable_hmaster1 & ~n46094;
  assign n46096 = ~n19685 & ~n46095;
  assign n46097 = ~i_hbusreq3 & ~n46096;
  assign n46098 = ~n46093 & ~n46097;
  assign n46099 = ~controllable_hmaster2 & ~n46098;
  assign n46100 = ~n19661 & ~n46099;
  assign n46101 = ~controllable_hgrant3 & ~n46100;
  assign n46102 = ~n19183 & ~n46101;
  assign n46103 = controllable_nhgrant0 & ~n46102;
  assign n46104 = ~n19213 & ~n46103;
  assign n46105 = ~n3281 & ~n46104;
  assign n46106 = ~n3281 & ~n46105;
  assign n46107 = n3378 & ~n46106;
  assign n46108 = ~n4333 & ~n45742;
  assign n46109 = ~controllable_hmaster0 & ~n46108;
  assign n46110 = ~n46062 & ~n46109;
  assign n46111 = ~controllable_hmaster1 & ~n46110;
  assign n46112 = ~n46061 & ~n46111;
  assign n46113 = i_hbusreq3 & ~n46112;
  assign n46114 = ~n4340 & ~n45753;
  assign n46115 = ~controllable_hmaster0 & ~n46114;
  assign n46116 = ~n46069 & ~n46115;
  assign n46117 = ~controllable_hmaster1 & ~n46116;
  assign n46118 = ~n46068 & ~n46117;
  assign n46119 = ~i_hbusreq3 & ~n46118;
  assign n46120 = ~n46113 & ~n46119;
  assign n46121 = controllable_hmaster2 & ~n46120;
  assign n46122 = ~n4333 & ~n45763;
  assign n46123 = controllable_hmaster0 & ~n46122;
  assign n46124 = ~n6697 & ~n45763;
  assign n46125 = ~controllable_hmaster0 & ~n46124;
  assign n46126 = ~n46123 & ~n46125;
  assign n46127 = controllable_hmaster1 & ~n46126;
  assign n46128 = ~controllable_hmaster0 & ~n46122;
  assign n46129 = ~n38936 & ~n46128;
  assign n46130 = ~controllable_hmaster1 & ~n46129;
  assign n46131 = ~n46127 & ~n46130;
  assign n46132 = i_hbusreq3 & ~n46131;
  assign n46133 = ~n4340 & ~n45779;
  assign n46134 = controllable_hmaster0 & ~n46133;
  assign n46135 = ~n6710 & ~n45779;
  assign n46136 = ~controllable_hmaster0 & ~n46135;
  assign n46137 = ~n46134 & ~n46136;
  assign n46138 = controllable_hmaster1 & ~n46137;
  assign n46139 = ~n6947 & ~n45789;
  assign n46140 = ~controllable_hmaster0 & ~n46139;
  assign n46141 = ~n38949 & ~n46140;
  assign n46142 = ~controllable_hmaster1 & ~n46141;
  assign n46143 = ~n46138 & ~n46142;
  assign n46144 = ~i_hbusreq3 & ~n46143;
  assign n46145 = ~n46132 & ~n46144;
  assign n46146 = ~controllable_hmaster2 & ~n46145;
  assign n46147 = ~n46121 & ~n46146;
  assign n46148 = ~controllable_hgrant3 & ~n46147;
  assign n46149 = ~n19225 & ~n46148;
  assign n46150 = controllable_nhgrant0 & ~n46149;
  assign n46151 = ~n19255 & ~n46150;
  assign n46152 = ~n3281 & ~n46151;
  assign n46153 = ~n3281 & ~n46152;
  assign n46154 = ~n3378 & ~n46153;
  assign n46155 = ~n46107 & ~n46154;
  assign n46156 = n3492 & ~n46155;
  assign n46157 = n3492 & ~n46156;
  assign n46158 = n3485 & ~n46157;
  assign n46159 = n3485 & ~n46158;
  assign n46160 = ~n3476 & ~n46159;
  assign n46161 = ~n8029 & ~n45813;
  assign n46162 = controllable_hmaster0 & ~n46161;
  assign n46163 = ~n19897 & ~n46162;
  assign n46164 = ~controllable_hmaster1 & ~n46163;
  assign n46165 = ~n19885 & ~n46164;
  assign n46166 = i_hbusreq3 & ~n46165;
  assign n46167 = ~n8036 & ~n45824;
  assign n46168 = controllable_hmaster0 & ~n46167;
  assign n46169 = ~n19941 & ~n46168;
  assign n46170 = ~controllable_hmaster1 & ~n46169;
  assign n46171 = ~n19912 & ~n46170;
  assign n46172 = ~i_hbusreq3 & ~n46171;
  assign n46173 = ~n46166 & ~n46172;
  assign n46174 = ~controllable_hmaster2 & ~n46173;
  assign n46175 = ~n19877 & ~n46174;
  assign n46176 = ~controllable_hgrant3 & ~n46175;
  assign n46177 = ~n19274 & ~n46176;
  assign n46178 = controllable_nhgrant0 & ~n46177;
  assign n46179 = ~n19385 & ~n46178;
  assign n46180 = ~n3281 & ~n46179;
  assign n46181 = ~n3281 & ~n46180;
  assign n46182 = n3378 & ~n46181;
  assign n46183 = ~n6762 & ~n45842;
  assign n46184 = controllable_hmaster1 & ~n46183;
  assign n46185 = controllable_hmaster0 & ~n46183;
  assign n46186 = ~n6762 & ~n45847;
  assign n46187 = ~controllable_hmaster0 & ~n46186;
  assign n46188 = ~n46185 & ~n46187;
  assign n46189 = ~controllable_hmaster1 & ~n46188;
  assign n46190 = ~n46184 & ~n46189;
  assign n46191 = i_hbusreq3 & ~n46190;
  assign n46192 = ~n6772 & ~n45858;
  assign n46193 = controllable_hmaster1 & ~n46192;
  assign n46194 = controllable_hmaster0 & ~n46192;
  assign n46195 = ~n6772 & ~n45866;
  assign n46196 = ~controllable_hmaster0 & ~n46195;
  assign n46197 = ~n46194 & ~n46196;
  assign n46198 = ~controllable_hmaster1 & ~n46197;
  assign n46199 = ~n46193 & ~n46198;
  assign n46200 = ~i_hbusreq3 & ~n46199;
  assign n46201 = ~n46191 & ~n46200;
  assign n46202 = controllable_hmaster2 & ~n46201;
  assign n46203 = ~n6762 & ~n45876;
  assign n46204 = controllable_hmaster0 & ~n46203;
  assign n46205 = ~n6786 & ~n45876;
  assign n46206 = ~controllable_hmaster0 & ~n46205;
  assign n46207 = ~n46204 & ~n46206;
  assign n46208 = controllable_hmaster1 & ~n46207;
  assign n46209 = ~n8056 & ~n45884;
  assign n46210 = controllable_hmaster0 & ~n46209;
  assign n46211 = ~controllable_hmaster0 & ~n46203;
  assign n46212 = ~n46210 & ~n46211;
  assign n46213 = ~controllable_hmaster1 & ~n46212;
  assign n46214 = ~n46208 & ~n46213;
  assign n46215 = i_hbusreq3 & ~n46214;
  assign n46216 = ~n6772 & ~n45896;
  assign n46217 = controllable_hmaster0 & ~n46216;
  assign n46218 = ~n6813 & ~n45896;
  assign n46219 = ~controllable_hmaster0 & ~n46218;
  assign n46220 = ~n46217 & ~n46219;
  assign n46221 = controllable_hmaster1 & ~n46220;
  assign n46222 = ~n8066 & ~n45907;
  assign n46223 = controllable_hmaster0 & ~n46222;
  assign n46224 = ~n6831 & ~n45913;
  assign n46225 = ~controllable_hmaster0 & ~n46224;
  assign n46226 = ~n46223 & ~n46225;
  assign n46227 = ~controllable_hmaster1 & ~n46226;
  assign n46228 = ~n46221 & ~n46227;
  assign n46229 = ~i_hbusreq3 & ~n46228;
  assign n46230 = ~n46215 & ~n46229;
  assign n46231 = ~controllable_hmaster2 & ~n46230;
  assign n46232 = ~n46202 & ~n46231;
  assign n46233 = ~controllable_hgrant3 & ~n46232;
  assign n46234 = ~n19398 & ~n46233;
  assign n46235 = controllable_nhgrant0 & ~n46234;
  assign n46236 = ~n19515 & ~n46235;
  assign n46237 = ~n3281 & ~n46236;
  assign n46238 = ~n3281 & ~n46237;
  assign n46239 = ~n3378 & ~n46238;
  assign n46240 = ~n46182 & ~n46239;
  assign n46241 = n3492 & ~n46240;
  assign n46242 = ~n18151 & ~n46241;
  assign n46243 = n3485 & ~n46242;
  assign n46244 = ~n18150 & ~n46243;
  assign n46245 = n3476 & ~n46244;
  assign n46246 = ~n46160 & ~n46245;
  assign n46247 = n3374 & ~n46246;
  assign n46248 = ~n46089 & ~n46247;
  assign n46249 = ~n3655 & ~n46248;
  assign n46250 = ~n46059 & ~n46249;
  assign n46251 = ~n3652 & ~n46250;
  assign n46252 = ~n45941 & ~n46251;
  assign n46253 = n3368 & ~n46252;
  assign n46254 = ~n45538 & ~n46253;
  assign n46255 = n3362 & ~n46254;
  assign n46256 = n3492 & ~n45006;
  assign n46257 = ~n3631 & ~n46256;
  assign n46258 = n3485 & ~n46257;
  assign n46259 = ~n3630 & ~n46258;
  assign n46260 = ~n3476 & ~n46259;
  assign n46261 = n3492 & ~n45065;
  assign n46262 = ~n3631 & ~n46261;
  assign n46263 = n3485 & ~n46262;
  assign n46264 = ~n41076 & ~n46263;
  assign n46265 = n3476 & ~n46264;
  assign n46266 = ~n46260 & ~n46265;
  assign n46267 = n3374 & ~n46266;
  assign n46268 = ~n41080 & ~n46267;
  assign n46269 = n3655 & ~n46268;
  assign n46270 = n3492 & ~n45106;
  assign n46271 = ~n3631 & ~n46270;
  assign n46272 = n3485 & ~n46271;
  assign n46273 = ~n3630 & ~n46272;
  assign n46274 = ~n3476 & ~n46273;
  assign n46275 = ~n20467 & ~n37048;
  assign n46276 = ~n3485 & ~n46275;
  assign n46277 = ~n18630 & ~n46270;
  assign n46278 = n3485 & ~n46277;
  assign n46279 = ~n46276 & ~n46278;
  assign n46280 = n3476 & ~n46279;
  assign n46281 = ~n46274 & ~n46280;
  assign n46282 = ~n3374 & ~n46281;
  assign n46283 = n3492 & ~n45177;
  assign n46284 = ~n3631 & ~n46283;
  assign n46285 = n3485 & ~n46284;
  assign n46286 = ~n3630 & ~n46285;
  assign n46287 = ~n3476 & ~n46286;
  assign n46288 = n3492 & ~n45259;
  assign n46289 = ~n18630 & ~n46288;
  assign n46290 = n3485 & ~n46289;
  assign n46291 = ~n46276 & ~n46290;
  assign n46292 = n3476 & ~n46291;
  assign n46293 = ~n46287 & ~n46292;
  assign n46294 = n3374 & ~n46293;
  assign n46295 = ~n46282 & ~n46294;
  assign n46296 = ~n3655 & ~n46295;
  assign n46297 = ~n46269 & ~n46296;
  assign n46298 = n3652 & ~n46297;
  assign n46299 = n3492 & ~n45313;
  assign n46300 = ~n3631 & ~n46299;
  assign n46301 = n3485 & ~n46300;
  assign n46302 = ~n3630 & ~n46301;
  assign n46303 = ~n3476 & ~n46302;
  assign n46304 = n3492 & ~n45361;
  assign n46305 = ~n3631 & ~n46304;
  assign n46306 = n3485 & ~n46305;
  assign n46307 = ~n41128 & ~n46306;
  assign n46308 = n3476 & ~n46307;
  assign n46309 = ~n46303 & ~n46308;
  assign n46310 = n3374 & ~n46309;
  assign n46311 = ~n41132 & ~n46310;
  assign n46312 = n3655 & ~n46311;
  assign n46313 = n3492 & ~n45395;
  assign n46314 = ~n3631 & ~n46313;
  assign n46315 = n3485 & ~n46314;
  assign n46316 = ~n3630 & ~n46315;
  assign n46317 = ~n3476 & ~n46316;
  assign n46318 = ~n20467 & ~n37132;
  assign n46319 = ~n3485 & ~n46318;
  assign n46320 = ~n18630 & ~n46313;
  assign n46321 = n3485 & ~n46320;
  assign n46322 = ~n46319 & ~n46321;
  assign n46323 = n3476 & ~n46322;
  assign n46324 = ~n46317 & ~n46323;
  assign n46325 = ~n3374 & ~n46324;
  assign n46326 = n3492 & ~n45459;
  assign n46327 = ~n3631 & ~n46326;
  assign n46328 = n3485 & ~n46327;
  assign n46329 = ~n3630 & ~n46328;
  assign n46330 = ~n3476 & ~n46329;
  assign n46331 = n3492 & ~n45523;
  assign n46332 = ~n18630 & ~n46331;
  assign n46333 = n3485 & ~n46332;
  assign n46334 = ~n46319 & ~n46333;
  assign n46335 = n3476 & ~n46334;
  assign n46336 = ~n46330 & ~n46335;
  assign n46337 = n3374 & ~n46336;
  assign n46338 = ~n46325 & ~n46337;
  assign n46339 = ~n3655 & ~n46338;
  assign n46340 = ~n46312 & ~n46339;
  assign n46341 = ~n3652 & ~n46340;
  assign n46342 = ~n46298 & ~n46341;
  assign n46343 = ~n3368 & ~n46342;
  assign n46344 = n3492 & ~n45573;
  assign n46345 = n3492 & ~n46344;
  assign n46346 = n3485 & ~n46345;
  assign n46347 = n3485 & ~n46346;
  assign n46348 = ~n3476 & ~n46347;
  assign n46349 = n3492 & ~n45674;
  assign n46350 = n3492 & ~n46349;
  assign n46351 = n3485 & ~n46350;
  assign n46352 = ~n41191 & ~n46351;
  assign n46353 = n3476 & ~n46352;
  assign n46354 = ~n46348 & ~n46353;
  assign n46355 = n3374 & ~n46354;
  assign n46356 = ~n41184 & ~n46355;
  assign n46357 = n3655 & ~n46356;
  assign n46358 = n3492 & ~n45715;
  assign n46359 = n3492 & ~n46358;
  assign n46360 = n3485 & ~n46359;
  assign n46361 = n3485 & ~n46360;
  assign n46362 = ~n3476 & ~n46361;
  assign n46363 = ~n8525 & ~n46360;
  assign n46364 = n3476 & ~n46363;
  assign n46365 = ~n46362 & ~n46364;
  assign n46366 = ~n3374 & ~n46365;
  assign n46367 = n3492 & ~n45804;
  assign n46368 = n3492 & ~n46367;
  assign n46369 = n3485 & ~n46368;
  assign n46370 = n3485 & ~n46369;
  assign n46371 = ~n3476 & ~n46370;
  assign n46372 = ~n20565 & ~n37202;
  assign n46373 = ~n3485 & ~n46372;
  assign n46374 = n3492 & ~n45928;
  assign n46375 = ~n18151 & ~n46374;
  assign n46376 = n3485 & ~n46375;
  assign n46377 = ~n46373 & ~n46376;
  assign n46378 = n3476 & ~n46377;
  assign n46379 = ~n46371 & ~n46378;
  assign n46380 = n3374 & ~n46379;
  assign n46381 = ~n46366 & ~n46380;
  assign n46382 = ~n3655 & ~n46381;
  assign n46383 = ~n46357 & ~n46382;
  assign n46384 = n3652 & ~n46383;
  assign n46385 = n3492 & ~n45976;
  assign n46386 = n3492 & ~n46385;
  assign n46387 = n3485 & ~n46386;
  assign n46388 = n3485 & ~n46387;
  assign n46389 = ~n3476 & ~n46388;
  assign n46390 = n3492 & ~n46048;
  assign n46391 = n3492 & ~n46390;
  assign n46392 = n3485 & ~n46391;
  assign n46393 = ~n41243 & ~n46392;
  assign n46394 = n3476 & ~n46393;
  assign n46395 = ~n46389 & ~n46394;
  assign n46396 = n3374 & ~n46395;
  assign n46397 = ~n41236 & ~n46396;
  assign n46398 = n3655 & ~n46397;
  assign n46399 = n3492 & ~n46082;
  assign n46400 = n3492 & ~n46399;
  assign n46401 = n3485 & ~n46400;
  assign n46402 = n3485 & ~n46401;
  assign n46403 = ~n3476 & ~n46402;
  assign n46404 = ~n8525 & ~n46401;
  assign n46405 = n3476 & ~n46404;
  assign n46406 = ~n46403 & ~n46405;
  assign n46407 = ~n3374 & ~n46406;
  assign n46408 = n3492 & ~n46153;
  assign n46409 = n3492 & ~n46408;
  assign n46410 = n3485 & ~n46409;
  assign n46411 = n3485 & ~n46410;
  assign n46412 = ~n3476 & ~n46411;
  assign n46413 = ~n20565 & ~n37258;
  assign n46414 = ~n3485 & ~n46413;
  assign n46415 = n3492 & ~n46238;
  assign n46416 = ~n18151 & ~n46415;
  assign n46417 = n3485 & ~n46416;
  assign n46418 = ~n46414 & ~n46417;
  assign n46419 = n3476 & ~n46418;
  assign n46420 = ~n46412 & ~n46419;
  assign n46421 = n3374 & ~n46420;
  assign n46422 = ~n46407 & ~n46421;
  assign n46423 = ~n3655 & ~n46422;
  assign n46424 = ~n46398 & ~n46423;
  assign n46425 = ~n3652 & ~n46424;
  assign n46426 = ~n46384 & ~n46425;
  assign n46427 = n3368 & ~n46426;
  assign n46428 = ~n46343 & ~n46427;
  assign n46429 = ~n3362 & ~n46428;
  assign n46430 = ~n46255 & ~n46429;
  assign n46431 = n3359 & ~n46430;
  assign n46432 = ~n37278 & ~n46263;
  assign n46433 = n3476 & ~n46432;
  assign n46434 = ~n46260 & ~n46433;
  assign n46435 = n3374 & ~n46434;
  assign n46436 = ~n41289 & ~n46435;
  assign n46437 = n3655 & ~n46436;
  assign n46438 = ~n37289 & ~n46278;
  assign n46439 = n3476 & ~n46438;
  assign n46440 = ~n46274 & ~n46439;
  assign n46441 = ~n3374 & ~n46440;
  assign n46442 = ~n37289 & ~n46290;
  assign n46443 = n3476 & ~n46442;
  assign n46444 = ~n46287 & ~n46443;
  assign n46445 = n3374 & ~n46444;
  assign n46446 = ~n46441 & ~n46445;
  assign n46447 = ~n3655 & ~n46446;
  assign n46448 = ~n46437 & ~n46447;
  assign n46449 = n3652 & ~n46448;
  assign n46450 = ~n37302 & ~n46306;
  assign n46451 = n3476 & ~n46450;
  assign n46452 = ~n46303 & ~n46451;
  assign n46453 = n3374 & ~n46452;
  assign n46454 = ~n41311 & ~n46453;
  assign n46455 = n3655 & ~n46454;
  assign n46456 = ~n37313 & ~n46321;
  assign n46457 = n3476 & ~n46456;
  assign n46458 = ~n46317 & ~n46457;
  assign n46459 = ~n3374 & ~n46458;
  assign n46460 = ~n37313 & ~n46333;
  assign n46461 = n3476 & ~n46460;
  assign n46462 = ~n46330 & ~n46461;
  assign n46463 = n3374 & ~n46462;
  assign n46464 = ~n46459 & ~n46463;
  assign n46465 = ~n3655 & ~n46464;
  assign n46466 = ~n46455 & ~n46465;
  assign n46467 = ~n3652 & ~n46466;
  assign n46468 = ~n46449 & ~n46467;
  assign n46469 = ~n3368 & ~n46468;
  assign n46470 = ~n37332 & ~n46351;
  assign n46471 = n3476 & ~n46470;
  assign n46472 = ~n46348 & ~n46471;
  assign n46473 = n3374 & ~n46472;
  assign n46474 = ~n41335 & ~n46473;
  assign n46475 = n3655 & ~n46474;
  assign n46476 = ~n8689 & ~n46360;
  assign n46477 = n3476 & ~n46476;
  assign n46478 = ~n46362 & ~n46477;
  assign n46479 = ~n3374 & ~n46478;
  assign n46480 = ~n37343 & ~n46376;
  assign n46481 = n3476 & ~n46480;
  assign n46482 = ~n46371 & ~n46481;
  assign n46483 = n3374 & ~n46482;
  assign n46484 = ~n46479 & ~n46483;
  assign n46485 = ~n3655 & ~n46484;
  assign n46486 = ~n46475 & ~n46485;
  assign n46487 = n3652 & ~n46486;
  assign n46488 = ~n37356 & ~n46392;
  assign n46489 = n3476 & ~n46488;
  assign n46490 = ~n46389 & ~n46489;
  assign n46491 = n3374 & ~n46490;
  assign n46492 = ~n41357 & ~n46491;
  assign n46493 = n3655 & ~n46492;
  assign n46494 = ~n8689 & ~n46401;
  assign n46495 = n3476 & ~n46494;
  assign n46496 = ~n46403 & ~n46495;
  assign n46497 = ~n3374 & ~n46496;
  assign n46498 = ~n37367 & ~n46417;
  assign n46499 = n3476 & ~n46498;
  assign n46500 = ~n46412 & ~n46499;
  assign n46501 = n3374 & ~n46500;
  assign n46502 = ~n46497 & ~n46501;
  assign n46503 = ~n3655 & ~n46502;
  assign n46504 = ~n46493 & ~n46503;
  assign n46505 = ~n3652 & ~n46504;
  assign n46506 = ~n46487 & ~n46505;
  assign n46507 = n3368 & ~n46506;
  assign n46508 = ~n46469 & ~n46507;
  assign n46509 = n3362 & ~n46508;
  assign n46510 = n3378 & ~n45006;
  assign n46511 = ~n37472 & ~n46510;
  assign n46512 = n3492 & ~n46511;
  assign n46513 = ~n3631 & ~n46512;
  assign n46514 = n3485 & ~n46513;
  assign n46515 = ~n3630 & ~n46514;
  assign n46516 = ~n3476 & ~n46515;
  assign n46517 = n3378 & ~n45065;
  assign n46518 = ~n37554 & ~n46517;
  assign n46519 = n3492 & ~n46518;
  assign n46520 = ~n37006 & ~n46519;
  assign n46521 = n3485 & ~n46520;
  assign n46522 = ~n37278 & ~n46521;
  assign n46523 = n3476 & ~n46522;
  assign n46524 = ~n46516 & ~n46523;
  assign n46525 = n3374 & ~n46524;
  assign n46526 = ~n41392 & ~n46525;
  assign n46527 = n3655 & ~n46526;
  assign n46528 = n3378 & ~n45106;
  assign n46529 = ~n37588 & ~n46528;
  assign n46530 = n3492 & ~n46529;
  assign n46531 = ~n3631 & ~n46530;
  assign n46532 = n3485 & ~n46531;
  assign n46533 = ~n3630 & ~n46532;
  assign n46534 = ~n3476 & ~n46533;
  assign n46535 = ~n37048 & ~n46530;
  assign n46536 = n3485 & ~n46535;
  assign n46537 = ~n37289 & ~n46536;
  assign n46538 = n3476 & ~n46537;
  assign n46539 = ~n46534 & ~n46538;
  assign n46540 = ~n3374 & ~n46539;
  assign n46541 = n3378 & ~n45177;
  assign n46542 = ~n37666 & ~n46541;
  assign n46543 = n3492 & ~n46542;
  assign n46544 = ~n3631 & ~n46543;
  assign n46545 = n3485 & ~n46544;
  assign n46546 = ~n3630 & ~n46545;
  assign n46547 = ~n3476 & ~n46546;
  assign n46548 = n3378 & ~n45259;
  assign n46549 = ~n37757 & ~n46548;
  assign n46550 = n3492 & ~n46549;
  assign n46551 = ~n37048 & ~n46550;
  assign n46552 = n3485 & ~n46551;
  assign n46553 = ~n37289 & ~n46552;
  assign n46554 = n3476 & ~n46553;
  assign n46555 = ~n46547 & ~n46554;
  assign n46556 = n3374 & ~n46555;
  assign n46557 = ~n46540 & ~n46556;
  assign n46558 = ~n3655 & ~n46557;
  assign n46559 = ~n46527 & ~n46558;
  assign n46560 = n3652 & ~n46559;
  assign n46561 = n3378 & ~n45313;
  assign n46562 = ~n37851 & ~n46561;
  assign n46563 = n3492 & ~n46562;
  assign n46564 = ~n3631 & ~n46563;
  assign n46565 = n3485 & ~n46564;
  assign n46566 = ~n3630 & ~n46565;
  assign n46567 = ~n3476 & ~n46566;
  assign n46568 = n3378 & ~n45361;
  assign n46569 = ~n37913 & ~n46568;
  assign n46570 = n3492 & ~n46569;
  assign n46571 = ~n37091 & ~n46570;
  assign n46572 = n3485 & ~n46571;
  assign n46573 = ~n37302 & ~n46572;
  assign n46574 = n3476 & ~n46573;
  assign n46575 = ~n46567 & ~n46574;
  assign n46576 = n3374 & ~n46575;
  assign n46577 = ~n41456 & ~n46576;
  assign n46578 = n3655 & ~n46577;
  assign n46579 = n3378 & ~n45395;
  assign n46580 = ~n37945 & ~n46579;
  assign n46581 = n3492 & ~n46580;
  assign n46582 = ~n3631 & ~n46581;
  assign n46583 = n3485 & ~n46582;
  assign n46584 = ~n3630 & ~n46583;
  assign n46585 = ~n3476 & ~n46584;
  assign n46586 = ~n37132 & ~n46581;
  assign n46587 = n3485 & ~n46586;
  assign n46588 = ~n37313 & ~n46587;
  assign n46589 = n3476 & ~n46588;
  assign n46590 = ~n46585 & ~n46589;
  assign n46591 = ~n3374 & ~n46590;
  assign n46592 = n3378 & ~n45459;
  assign n46593 = ~n38005 & ~n46592;
  assign n46594 = n3492 & ~n46593;
  assign n46595 = ~n3631 & ~n46594;
  assign n46596 = n3485 & ~n46595;
  assign n46597 = ~n3630 & ~n46596;
  assign n46598 = ~n3476 & ~n46597;
  assign n46599 = n3378 & ~n45523;
  assign n46600 = ~n38067 & ~n46599;
  assign n46601 = n3492 & ~n46600;
  assign n46602 = ~n37132 & ~n46601;
  assign n46603 = n3485 & ~n46602;
  assign n46604 = ~n37313 & ~n46603;
  assign n46605 = n3476 & ~n46604;
  assign n46606 = ~n46598 & ~n46605;
  assign n46607 = n3374 & ~n46606;
  assign n46608 = ~n46591 & ~n46607;
  assign n46609 = ~n3655 & ~n46608;
  assign n46610 = ~n46578 & ~n46609;
  assign n46611 = ~n3652 & ~n46610;
  assign n46612 = ~n46560 & ~n46611;
  assign n46613 = ~n3368 & ~n46612;
  assign n46614 = n3378 & ~n45573;
  assign n46615 = ~n38186 & ~n46614;
  assign n46616 = n3492 & ~n46615;
  assign n46617 = n3492 & ~n46616;
  assign n46618 = n3485 & ~n46617;
  assign n46619 = n3485 & ~n46618;
  assign n46620 = ~n3476 & ~n46619;
  assign n46621 = ~n20822 & ~n41558;
  assign n46622 = ~i_hbusreq2 & ~n46621;
  assign n46623 = ~n41551 & ~n46622;
  assign n46624 = ~controllable_hgrant2 & ~n46623;
  assign n46625 = ~n5862 & ~n46624;
  assign n46626 = controllable_hmaster1 & ~n46625;
  assign n46627 = controllable_hmaster0 & ~n46625;
  assign n46628 = ~n20837 & ~n41573;
  assign n46629 = ~i_hbusreq2 & ~n46628;
  assign n46630 = ~n41566 & ~n46629;
  assign n46631 = ~controllable_hgrant2 & ~n46630;
  assign n46632 = ~n5862 & ~n46631;
  assign n46633 = ~controllable_hmaster0 & ~n46632;
  assign n46634 = ~n46627 & ~n46633;
  assign n46635 = ~controllable_hmaster1 & ~n46634;
  assign n46636 = ~n46626 & ~n46635;
  assign n46637 = ~i_hbusreq3 & ~n46636;
  assign n46638 = ~n41550 & ~n46637;
  assign n46639 = controllable_hmaster2 & ~n46638;
  assign n46640 = ~n41589 & ~n44070;
  assign n46641 = controllable_hmaster1 & ~n46640;
  assign n46642 = ~n38324 & ~n41597;
  assign n46643 = ~controllable_hmaster1 & ~n46642;
  assign n46644 = ~n46641 & ~n46643;
  assign n46645 = i_hbusreq3 & ~n46644;
  assign n46646 = ~n20837 & ~n41558;
  assign n46647 = ~i_hbusreq2 & ~n46646;
  assign n46648 = ~n41614 & ~n46647;
  assign n46649 = ~controllable_hgrant2 & ~n46648;
  assign n46650 = ~n5862 & ~n46649;
  assign n46651 = controllable_hmaster0 & ~n46650;
  assign n46652 = ~n5950 & ~n46649;
  assign n46653 = ~controllable_hmaster0 & ~n46652;
  assign n46654 = ~n46651 & ~n46653;
  assign n46655 = controllable_hmaster1 & ~n46654;
  assign n46656 = ~n20871 & ~n41607;
  assign n46657 = ~i_hbusreq2 & ~n46656;
  assign n46658 = ~n38340 & ~n46657;
  assign n46659 = ~controllable_hgrant2 & ~n46658;
  assign n46660 = ~n7507 & ~n46659;
  assign n46661 = controllable_hmaster0 & ~n46660;
  assign n46662 = ~n20885 & ~n41635;
  assign n46663 = ~i_hbusreq2 & ~n46662;
  assign n46664 = ~n41614 & ~n46663;
  assign n46665 = ~controllable_hgrant2 & ~n46664;
  assign n46666 = ~n5981 & ~n46665;
  assign n46667 = ~controllable_hmaster0 & ~n46666;
  assign n46668 = ~n46661 & ~n46667;
  assign n46669 = ~controllable_hmaster1 & ~n46668;
  assign n46670 = ~n46655 & ~n46669;
  assign n46671 = ~i_hbusreq3 & ~n46670;
  assign n46672 = ~n46645 & ~n46671;
  assign n46673 = ~controllable_hmaster2 & ~n46672;
  assign n46674 = ~n46639 & ~n46673;
  assign n46675 = ~controllable_hgrant3 & ~n46674;
  assign n46676 = ~n19398 & ~n46675;
  assign n46677 = controllable_nhgrant0 & ~n46676;
  assign n46678 = ~n20915 & ~n46677;
  assign n46679 = ~n3281 & ~n46678;
  assign n46680 = ~n3281 & ~n46679;
  assign n46681 = n3378 & ~n46680;
  assign n46682 = ~n38371 & ~n46681;
  assign n46683 = n3492 & ~n46682;
  assign n46684 = ~n37174 & ~n46683;
  assign n46685 = n3485 & ~n46684;
  assign n46686 = ~n37332 & ~n46685;
  assign n46687 = n3476 & ~n46686;
  assign n46688 = ~n46620 & ~n46687;
  assign n46689 = n3374 & ~n46688;
  assign n46690 = ~n41522 & ~n46689;
  assign n46691 = n3655 & ~n46690;
  assign n46692 = n3378 & ~n45715;
  assign n46693 = ~n38413 & ~n46692;
  assign n46694 = n3492 & ~n46693;
  assign n46695 = n3492 & ~n46694;
  assign n46696 = n3485 & ~n46695;
  assign n46697 = n3485 & ~n46696;
  assign n46698 = ~n3476 & ~n46697;
  assign n46699 = ~n8523 & ~n46694;
  assign n46700 = n3485 & ~n46699;
  assign n46701 = ~n8689 & ~n46700;
  assign n46702 = n3476 & ~n46701;
  assign n46703 = ~n46698 & ~n46702;
  assign n46704 = ~n3374 & ~n46703;
  assign n46705 = n3378 & ~n45804;
  assign n46706 = ~n38485 & ~n46705;
  assign n46707 = n3492 & ~n46706;
  assign n46708 = n3492 & ~n46707;
  assign n46709 = n3485 & ~n46708;
  assign n46710 = n3485 & ~n46709;
  assign n46711 = ~n3476 & ~n46710;
  assign n46712 = ~n20951 & ~n41533;
  assign n46713 = ~controllable_hgrant2 & ~n46712;
  assign n46714 = ~n5616 & ~n46713;
  assign n46715 = controllable_hmaster1 & ~n46714;
  assign n46716 = controllable_hmaster0 & ~n46714;
  assign n46717 = ~n20958 & ~n41542;
  assign n46718 = ~controllable_hgrant2 & ~n46717;
  assign n46719 = ~n5616 & ~n46718;
  assign n46720 = ~controllable_hmaster0 & ~n46719;
  assign n46721 = ~n46716 & ~n46720;
  assign n46722 = ~controllable_hmaster1 & ~n46721;
  assign n46723 = ~n46715 & ~n46722;
  assign n46724 = i_hbusreq3 & ~n46723;
  assign n46725 = i_hbusreq2 & ~n46712;
  assign n46726 = ~n20983 & ~n41558;
  assign n46727 = ~i_hbusreq2 & ~n46726;
  assign n46728 = ~n46725 & ~n46727;
  assign n46729 = ~controllable_hgrant2 & ~n46728;
  assign n46730 = ~n5862 & ~n46729;
  assign n46731 = controllable_hmaster1 & ~n46730;
  assign n46732 = controllable_hmaster0 & ~n46730;
  assign n46733 = i_hbusreq2 & ~n46717;
  assign n46734 = ~n21003 & ~n41573;
  assign n46735 = ~i_hbusreq2 & ~n46734;
  assign n46736 = ~n46733 & ~n46735;
  assign n46737 = ~controllable_hgrant2 & ~n46736;
  assign n46738 = ~n5862 & ~n46737;
  assign n46739 = ~controllable_hmaster0 & ~n46738;
  assign n46740 = ~n46732 & ~n46739;
  assign n46741 = ~controllable_hmaster1 & ~n46740;
  assign n46742 = ~n46731 & ~n46741;
  assign n46743 = ~i_hbusreq3 & ~n46742;
  assign n46744 = ~n46724 & ~n46743;
  assign n46745 = controllable_hmaster2 & ~n46744;
  assign n46746 = ~n20958 & ~n41533;
  assign n46747 = ~controllable_hgrant2 & ~n46746;
  assign n46748 = ~n5616 & ~n46747;
  assign n46749 = controllable_hmaster0 & ~n46748;
  assign n46750 = ~n5686 & ~n46747;
  assign n46751 = ~controllable_hmaster0 & ~n46750;
  assign n46752 = ~n46749 & ~n46751;
  assign n46753 = controllable_hmaster1 & ~n46752;
  assign n46754 = ~controllable_hmaster0 & ~n46748;
  assign n46755 = ~n38617 & ~n46754;
  assign n46756 = ~controllable_hmaster1 & ~n46755;
  assign n46757 = ~n46753 & ~n46756;
  assign n46758 = i_hbusreq3 & ~n46757;
  assign n46759 = i_hbusreq2 & ~n46746;
  assign n46760 = ~n21003 & ~n41558;
  assign n46761 = ~i_hbusreq2 & ~n46760;
  assign n46762 = ~n46759 & ~n46761;
  assign n46763 = ~controllable_hgrant2 & ~n46762;
  assign n46764 = ~n5862 & ~n46763;
  assign n46765 = controllable_hmaster0 & ~n46764;
  assign n46766 = ~n5950 & ~n46763;
  assign n46767 = ~controllable_hmaster0 & ~n46766;
  assign n46768 = ~n46765 & ~n46767;
  assign n46769 = controllable_hmaster1 & ~n46768;
  assign n46770 = ~n21051 & ~n41607;
  assign n46771 = ~i_hbusreq2 & ~n46770;
  assign n46772 = ~n38633 & ~n46771;
  assign n46773 = ~controllable_hgrant2 & ~n46772;
  assign n46774 = ~n7507 & ~n46773;
  assign n46775 = controllable_hmaster0 & ~n46774;
  assign n46776 = ~n21065 & ~n41635;
  assign n46777 = ~i_hbusreq2 & ~n46776;
  assign n46778 = ~n46759 & ~n46777;
  assign n46779 = ~controllable_hgrant2 & ~n46778;
  assign n46780 = ~n5981 & ~n46779;
  assign n46781 = ~controllable_hmaster0 & ~n46780;
  assign n46782 = ~n46775 & ~n46781;
  assign n46783 = ~controllable_hmaster1 & ~n46782;
  assign n46784 = ~n46769 & ~n46783;
  assign n46785 = ~i_hbusreq3 & ~n46784;
  assign n46786 = ~n46758 & ~n46785;
  assign n46787 = ~controllable_hmaster2 & ~n46786;
  assign n46788 = ~n46745 & ~n46787;
  assign n46789 = ~controllable_hgrant3 & ~n46788;
  assign n46790 = ~n19398 & ~n46789;
  assign n46791 = controllable_nhgrant0 & ~n46790;
  assign n46792 = ~n20915 & ~n46791;
  assign n46793 = ~n3281 & ~n46792;
  assign n46794 = ~n3281 & ~n46793;
  assign n46795 = n3378 & ~n46794;
  assign n46796 = ~n38659 & ~n46795;
  assign n46797 = n3492 & ~n46796;
  assign n46798 = ~n37202 & ~n46797;
  assign n46799 = n3485 & ~n46798;
  assign n46800 = ~n37343 & ~n46799;
  assign n46801 = n3476 & ~n46800;
  assign n46802 = ~n46711 & ~n46801;
  assign n46803 = n3374 & ~n46802;
  assign n46804 = ~n46704 & ~n46803;
  assign n46805 = ~n3655 & ~n46804;
  assign n46806 = ~n46691 & ~n46805;
  assign n46807 = n3652 & ~n46806;
  assign n46808 = n3378 & ~n45976;
  assign n46809 = ~n38754 & ~n46808;
  assign n46810 = n3492 & ~n46809;
  assign n46811 = n3492 & ~n46810;
  assign n46812 = n3485 & ~n46811;
  assign n46813 = n3485 & ~n46812;
  assign n46814 = ~n3476 & ~n46813;
  assign n46815 = ~n10870 & ~n46624;
  assign n46816 = controllable_hmaster1 & ~n46815;
  assign n46817 = controllable_hmaster0 & ~n46815;
  assign n46818 = ~n10870 & ~n46631;
  assign n46819 = ~controllable_hmaster0 & ~n46818;
  assign n46820 = ~n46817 & ~n46819;
  assign n46821 = ~controllable_hmaster1 & ~n46820;
  assign n46822 = ~n46816 & ~n46821;
  assign n46823 = ~i_hbusreq3 & ~n46822;
  assign n46824 = ~n41818 & ~n46823;
  assign n46825 = controllable_hmaster2 & ~n46824;
  assign n46826 = controllable_hmaster0 & ~n41836;
  assign n46827 = ~n41831 & ~n46826;
  assign n46828 = controllable_hmaster1 & ~n46827;
  assign n46829 = ~n38841 & ~n41837;
  assign n46830 = ~controllable_hmaster1 & ~n46829;
  assign n46831 = ~n46828 & ~n46830;
  assign n46832 = i_hbusreq3 & ~n46831;
  assign n46833 = ~n10870 & ~n46649;
  assign n46834 = controllable_hmaster0 & ~n46833;
  assign n46835 = ~n10972 & ~n46649;
  assign n46836 = ~controllable_hmaster0 & ~n46835;
  assign n46837 = ~n46834 & ~n46836;
  assign n46838 = controllable_hmaster1 & ~n46837;
  assign n46839 = ~n10904 & ~n46659;
  assign n46840 = controllable_hmaster0 & ~n46839;
  assign n46841 = ~n11002 & ~n46665;
  assign n46842 = ~controllable_hmaster0 & ~n46841;
  assign n46843 = ~n46840 & ~n46842;
  assign n46844 = ~controllable_hmaster1 & ~n46843;
  assign n46845 = ~n46838 & ~n46844;
  assign n46846 = ~i_hbusreq3 & ~n46845;
  assign n46847 = ~n46832 & ~n46846;
  assign n46848 = ~controllable_hmaster2 & ~n46847;
  assign n46849 = ~n46825 & ~n46848;
  assign n46850 = ~controllable_hgrant3 & ~n46849;
  assign n46851 = ~n19398 & ~n46850;
  assign n46852 = controllable_nhgrant0 & ~n46851;
  assign n46853 = ~n20915 & ~n46852;
  assign n46854 = ~n3281 & ~n46853;
  assign n46855 = ~n3281 & ~n46854;
  assign n46856 = n3378 & ~n46855;
  assign n46857 = ~n38870 & ~n46856;
  assign n46858 = n3492 & ~n46857;
  assign n46859 = ~n37231 & ~n46858;
  assign n46860 = n3485 & ~n46859;
  assign n46861 = ~n37356 & ~n46860;
  assign n46862 = n3476 & ~n46861;
  assign n46863 = ~n46814 & ~n46862;
  assign n46864 = n3374 & ~n46863;
  assign n46865 = ~n41802 & ~n46864;
  assign n46866 = n3655 & ~n46865;
  assign n46867 = n3378 & ~n46082;
  assign n46868 = ~n38905 & ~n46867;
  assign n46869 = n3492 & ~n46868;
  assign n46870 = n3492 & ~n46869;
  assign n46871 = n3485 & ~n46870;
  assign n46872 = n3485 & ~n46871;
  assign n46873 = ~n3476 & ~n46872;
  assign n46874 = ~n8523 & ~n46869;
  assign n46875 = n3485 & ~n46874;
  assign n46876 = ~n8689 & ~n46875;
  assign n46877 = n3476 & ~n46876;
  assign n46878 = ~n46873 & ~n46877;
  assign n46879 = ~n3374 & ~n46878;
  assign n46880 = n3378 & ~n46153;
  assign n46881 = ~n38963 & ~n46880;
  assign n46882 = n3492 & ~n46881;
  assign n46883 = n3492 & ~n46882;
  assign n46884 = n3485 & ~n46883;
  assign n46885 = n3485 & ~n46884;
  assign n46886 = ~n3476 & ~n46885;
  assign n46887 = ~n10816 & ~n46713;
  assign n46888 = controllable_hmaster1 & ~n46887;
  assign n46889 = controllable_hmaster0 & ~n46887;
  assign n46890 = ~n10816 & ~n46718;
  assign n46891 = ~controllable_hmaster0 & ~n46890;
  assign n46892 = ~n46889 & ~n46891;
  assign n46893 = ~controllable_hmaster1 & ~n46892;
  assign n46894 = ~n46888 & ~n46893;
  assign n46895 = i_hbusreq3 & ~n46894;
  assign n46896 = ~n10870 & ~n46729;
  assign n46897 = controllable_hmaster1 & ~n46896;
  assign n46898 = controllable_hmaster0 & ~n46896;
  assign n46899 = ~n10870 & ~n46737;
  assign n46900 = ~controllable_hmaster0 & ~n46899;
  assign n46901 = ~n46898 & ~n46900;
  assign n46902 = ~controllable_hmaster1 & ~n46901;
  assign n46903 = ~n46897 & ~n46902;
  assign n46904 = ~i_hbusreq3 & ~n46903;
  assign n46905 = ~n46895 & ~n46904;
  assign n46906 = controllable_hmaster2 & ~n46905;
  assign n46907 = ~n10816 & ~n46747;
  assign n46908 = controllable_hmaster0 & ~n46907;
  assign n46909 = ~n10922 & ~n46747;
  assign n46910 = ~controllable_hmaster0 & ~n46909;
  assign n46911 = ~n46908 & ~n46910;
  assign n46912 = controllable_hmaster1 & ~n46911;
  assign n46913 = ~controllable_hmaster0 & ~n46907;
  assign n46914 = ~n39050 & ~n46913;
  assign n46915 = ~controllable_hmaster1 & ~n46914;
  assign n46916 = ~n46912 & ~n46915;
  assign n46917 = i_hbusreq3 & ~n46916;
  assign n46918 = ~n10870 & ~n46763;
  assign n46919 = controllable_hmaster0 & ~n46918;
  assign n46920 = ~n10972 & ~n46763;
  assign n46921 = ~controllable_hmaster0 & ~n46920;
  assign n46922 = ~n46919 & ~n46921;
  assign n46923 = controllable_hmaster1 & ~n46922;
  assign n46924 = ~n10904 & ~n46773;
  assign n46925 = controllable_hmaster0 & ~n46924;
  assign n46926 = ~n11002 & ~n46779;
  assign n46927 = ~controllable_hmaster0 & ~n46926;
  assign n46928 = ~n46925 & ~n46927;
  assign n46929 = ~controllable_hmaster1 & ~n46928;
  assign n46930 = ~n46923 & ~n46929;
  assign n46931 = ~i_hbusreq3 & ~n46930;
  assign n46932 = ~n46917 & ~n46931;
  assign n46933 = ~controllable_hmaster2 & ~n46932;
  assign n46934 = ~n46906 & ~n46933;
  assign n46935 = ~controllable_hgrant3 & ~n46934;
  assign n46936 = ~n19398 & ~n46935;
  assign n46937 = controllable_nhgrant0 & ~n46936;
  assign n46938 = ~n20915 & ~n46937;
  assign n46939 = ~n3281 & ~n46938;
  assign n46940 = ~n3281 & ~n46939;
  assign n46941 = n3378 & ~n46940;
  assign n46942 = ~n39079 & ~n46941;
  assign n46943 = n3492 & ~n46942;
  assign n46944 = ~n37258 & ~n46943;
  assign n46945 = n3485 & ~n46944;
  assign n46946 = ~n37367 & ~n46945;
  assign n46947 = n3476 & ~n46946;
  assign n46948 = ~n46886 & ~n46947;
  assign n46949 = n3374 & ~n46948;
  assign n46950 = ~n46879 & ~n46949;
  assign n46951 = ~n3655 & ~n46950;
  assign n46952 = ~n46866 & ~n46951;
  assign n46953 = ~n3652 & ~n46952;
  assign n46954 = ~n46807 & ~n46953;
  assign n46955 = n3368 & ~n46954;
  assign n46956 = ~n46613 & ~n46955;
  assign n46957 = ~n3362 & ~n46956;
  assign n46958 = ~n46509 & ~n46957;
  assign n46959 = ~n3359 & ~n46958;
  assign n46960 = ~n46431 & ~n46959;
  assign n46961 = ~n3356 & ~n46960;
  assign n46962 = ~n44965 & ~n46961;
  assign n46963 = ~n3345 & ~n46962;
  assign n46964 = ~controllable_hmaster0 & ~n37430;
  assign n46965 = ~controllable_hmaster1 & ~n46964;
  assign n46966 = ~controllable_hmaster1 & ~n46965;
  assign n46967 = i_hbusreq3 & ~n46966;
  assign n46968 = ~controllable_hmaster0 & ~n37458;
  assign n46969 = ~controllable_hmaster1 & ~n46968;
  assign n46970 = ~controllable_hmaster1 & ~n46969;
  assign n46971 = ~i_hbusreq3 & ~n46970;
  assign n46972 = ~n46967 & ~n46971;
  assign n46973 = ~controllable_hmaster2 & ~n46972;
  assign n46974 = ~controllable_hmaster2 & ~n46973;
  assign n46975 = ~controllable_hgrant3 & ~n46974;
  assign n46976 = ~n21304 & ~n46975;
  assign n46977 = controllable_nhgrant0 & ~n46976;
  assign n46978 = ~n21332 & ~n46977;
  assign n46979 = ~n3281 & ~n46978;
  assign n46980 = ~n3281 & ~n46979;
  assign n46981 = n3378 & ~n46980;
  assign n46982 = ~n21339 & ~n46973;
  assign n46983 = ~controllable_hgrant3 & ~n46982;
  assign n46984 = ~n21338 & ~n46983;
  assign n46985 = controllable_nhgrant0 & ~n46984;
  assign n46986 = ~n21347 & ~n46985;
  assign n46987 = ~n3281 & ~n46986;
  assign n46988 = ~n3950 & ~n46987;
  assign n46989 = ~n3378 & ~n46988;
  assign n46990 = ~n46981 & ~n46989;
  assign n46991 = n3492 & ~n46990;
  assign n46992 = ~n3493 & ~n46991;
  assign n46993 = n3485 & ~n46992;
  assign n46994 = ~n3486 & ~n46993;
  assign n46995 = ~n3476 & ~n46994;
  assign n46996 = ~n21383 & ~n46977;
  assign n46997 = ~n3281 & ~n46996;
  assign n46998 = ~n3281 & ~n46997;
  assign n46999 = n3378 & ~n46998;
  assign n47000 = ~controllable_hmaster0 & ~n39144;
  assign n47001 = ~n21412 & ~n47000;
  assign n47002 = ~controllable_hmaster1 & ~n47001;
  assign n47003 = ~n21411 & ~n47002;
  assign n47004 = i_hbusreq3 & ~n47003;
  assign n47005 = ~n21429 & ~n35392;
  assign n47006 = ~i_hbusreq2 & ~n47005;
  assign n47007 = ~n39150 & ~n47006;
  assign n47008 = ~controllable_hgrant2 & ~n47007;
  assign n47009 = ~n5461 & ~n47008;
  assign n47010 = ~controllable_hmaster0 & ~n47009;
  assign n47011 = ~n21419 & ~n47010;
  assign n47012 = ~controllable_hmaster1 & ~n47011;
  assign n47013 = ~n21418 & ~n47012;
  assign n47014 = ~i_hbusreq3 & ~n47013;
  assign n47015 = ~n47004 & ~n47014;
  assign n47016 = ~controllable_hmaster2 & ~n47015;
  assign n47017 = ~n21410 & ~n47016;
  assign n47018 = ~controllable_hgrant3 & ~n47017;
  assign n47019 = ~n21338 & ~n47018;
  assign n47020 = controllable_nhgrant0 & ~n47019;
  assign n47021 = ~n21461 & ~n47020;
  assign n47022 = ~n3281 & ~n47021;
  assign n47023 = ~n4089 & ~n47022;
  assign n47024 = ~n3378 & ~n47023;
  assign n47025 = ~n46999 & ~n47024;
  assign n47026 = n3492 & ~n47025;
  assign n47027 = ~n21290 & ~n47026;
  assign n47028 = n3485 & ~n47027;
  assign n47029 = ~n21289 & ~n47028;
  assign n47030 = n3476 & ~n47029;
  assign n47031 = ~n46995 & ~n47030;
  assign n47032 = n3374 & ~n47031;
  assign n47033 = ~n21296 & ~n47032;
  assign n47034 = n3655 & ~n47033;
  assign n47035 = ~controllable_hmaster0 & ~n37624;
  assign n47036 = ~controllable_hmaster1 & ~n47035;
  assign n47037 = ~controllable_hmaster1 & ~n47036;
  assign n47038 = i_hbusreq3 & ~n47037;
  assign n47039 = ~controllable_hmaster0 & ~n37652;
  assign n47040 = ~controllable_hmaster1 & ~n47039;
  assign n47041 = ~controllable_hmaster1 & ~n47040;
  assign n47042 = ~i_hbusreq3 & ~n47041;
  assign n47043 = ~n47038 & ~n47042;
  assign n47044 = ~controllable_hmaster2 & ~n47043;
  assign n47045 = ~controllable_hmaster2 & ~n47044;
  assign n47046 = ~controllable_hgrant3 & ~n47045;
  assign n47047 = ~n21304 & ~n47046;
  assign n47048 = controllable_nhgrant0 & ~n47047;
  assign n47049 = ~n21332 & ~n47048;
  assign n47050 = ~n3281 & ~n47049;
  assign n47051 = ~n3281 & ~n47050;
  assign n47052 = n3378 & ~n47051;
  assign n47053 = ~n21339 & ~n47044;
  assign n47054 = ~controllable_hgrant3 & ~n47053;
  assign n47055 = ~n21338 & ~n47054;
  assign n47056 = controllable_nhgrant0 & ~n47055;
  assign n47057 = ~n21347 & ~n47056;
  assign n47058 = ~n3281 & ~n47057;
  assign n47059 = ~n3950 & ~n47058;
  assign n47060 = ~n3378 & ~n47059;
  assign n47061 = ~n47052 & ~n47060;
  assign n47062 = n3492 & ~n47061;
  assign n47063 = ~n3493 & ~n47062;
  assign n47064 = n3485 & ~n47063;
  assign n47065 = ~n3486 & ~n47064;
  assign n47066 = ~n3476 & ~n47065;
  assign n47067 = ~n21383 & ~n47048;
  assign n47068 = ~n3281 & ~n47067;
  assign n47069 = ~n3281 & ~n47068;
  assign n47070 = n3378 & ~n47069;
  assign n47071 = ~controllable_hmaster0 & ~n39221;
  assign n47072 = ~n21412 & ~n47071;
  assign n47073 = ~controllable_hmaster1 & ~n47072;
  assign n47074 = ~n21411 & ~n47073;
  assign n47075 = i_hbusreq3 & ~n47074;
  assign n47076 = ~n21526 & ~n35392;
  assign n47077 = ~i_hbusreq2 & ~n47076;
  assign n47078 = ~n39227 & ~n47077;
  assign n47079 = ~controllable_hgrant2 & ~n47078;
  assign n47080 = ~n5461 & ~n47079;
  assign n47081 = ~controllable_hmaster0 & ~n47080;
  assign n47082 = ~n21419 & ~n47081;
  assign n47083 = ~controllable_hmaster1 & ~n47082;
  assign n47084 = ~n21418 & ~n47083;
  assign n47085 = ~i_hbusreq3 & ~n47084;
  assign n47086 = ~n47075 & ~n47085;
  assign n47087 = ~controllable_hmaster2 & ~n47086;
  assign n47088 = ~n21410 & ~n47087;
  assign n47089 = ~controllable_hgrant3 & ~n47088;
  assign n47090 = ~n21338 & ~n47089;
  assign n47091 = controllable_nhgrant0 & ~n47090;
  assign n47092 = ~n21461 & ~n47091;
  assign n47093 = ~n3281 & ~n47092;
  assign n47094 = ~n4089 & ~n47093;
  assign n47095 = ~n3378 & ~n47094;
  assign n47096 = ~n47070 & ~n47095;
  assign n47097 = n3492 & ~n47096;
  assign n47098 = ~n21290 & ~n47097;
  assign n47099 = n3485 & ~n47098;
  assign n47100 = ~n21289 & ~n47099;
  assign n47101 = n3476 & ~n47100;
  assign n47102 = ~n47066 & ~n47101;
  assign n47103 = n3374 & ~n47102;
  assign n47104 = ~n21296 & ~n47103;
  assign n47105 = ~n3655 & ~n47104;
  assign n47106 = ~n47034 & ~n47105;
  assign n47107 = n3652 & ~n47106;
  assign n47108 = ~controllable_hmaster0 & ~n37823;
  assign n47109 = ~controllable_hmaster1 & ~n47108;
  assign n47110 = ~controllable_hmaster1 & ~n47109;
  assign n47111 = i_hbusreq3 & ~n47110;
  assign n47112 = ~controllable_hmaster0 & ~n37837;
  assign n47113 = ~controllable_hmaster1 & ~n47112;
  assign n47114 = ~controllable_hmaster1 & ~n47113;
  assign n47115 = ~i_hbusreq3 & ~n47114;
  assign n47116 = ~n47111 & ~n47115;
  assign n47117 = ~controllable_hmaster2 & ~n47116;
  assign n47118 = ~controllable_hmaster2 & ~n47117;
  assign n47119 = ~controllable_hgrant3 & ~n47118;
  assign n47120 = ~n21304 & ~n47119;
  assign n47121 = controllable_nhgrant0 & ~n47120;
  assign n47122 = ~n21332 & ~n47121;
  assign n47123 = ~n3281 & ~n47122;
  assign n47124 = ~n3281 & ~n47123;
  assign n47125 = n3378 & ~n47124;
  assign n47126 = ~n21339 & ~n47117;
  assign n47127 = ~controllable_hgrant3 & ~n47126;
  assign n47128 = ~n21338 & ~n47127;
  assign n47129 = controllable_nhgrant0 & ~n47128;
  assign n47130 = ~n21347 & ~n47129;
  assign n47131 = ~n3281 & ~n47130;
  assign n47132 = ~n3950 & ~n47131;
  assign n47133 = ~n3378 & ~n47132;
  assign n47134 = ~n47125 & ~n47133;
  assign n47135 = n3492 & ~n47134;
  assign n47136 = ~n3493 & ~n47135;
  assign n47137 = n3485 & ~n47136;
  assign n47138 = ~n3486 & ~n47137;
  assign n47139 = ~n3476 & ~n47138;
  assign n47140 = ~n21383 & ~n47121;
  assign n47141 = ~n3281 & ~n47140;
  assign n47142 = ~n3281 & ~n47141;
  assign n47143 = n3378 & ~n47142;
  assign n47144 = ~controllable_hmaster0 & ~n39298;
  assign n47145 = ~n21412 & ~n47144;
  assign n47146 = ~controllable_hmaster1 & ~n47145;
  assign n47147 = ~n21411 & ~n47146;
  assign n47148 = i_hbusreq3 & ~n47147;
  assign n47149 = ~n6947 & ~n47008;
  assign n47150 = ~controllable_hmaster0 & ~n47149;
  assign n47151 = ~n21419 & ~n47150;
  assign n47152 = ~controllable_hmaster1 & ~n47151;
  assign n47153 = ~n21418 & ~n47152;
  assign n47154 = ~i_hbusreq3 & ~n47153;
  assign n47155 = ~n47148 & ~n47154;
  assign n47156 = ~controllable_hmaster2 & ~n47155;
  assign n47157 = ~n21410 & ~n47156;
  assign n47158 = ~controllable_hgrant3 & ~n47157;
  assign n47159 = ~n21338 & ~n47158;
  assign n47160 = controllable_nhgrant0 & ~n47159;
  assign n47161 = ~n21461 & ~n47160;
  assign n47162 = ~n3281 & ~n47161;
  assign n47163 = ~n4089 & ~n47162;
  assign n47164 = ~n3378 & ~n47163;
  assign n47165 = ~n47143 & ~n47164;
  assign n47166 = n3492 & ~n47165;
  assign n47167 = ~n21290 & ~n47166;
  assign n47168 = n3485 & ~n47167;
  assign n47169 = ~n21289 & ~n47168;
  assign n47170 = n3476 & ~n47169;
  assign n47171 = ~n47139 & ~n47170;
  assign n47172 = n3374 & ~n47171;
  assign n47173 = ~n21296 & ~n47172;
  assign n47174 = n3655 & ~n47173;
  assign n47175 = ~controllable_hmaster0 & ~n37977;
  assign n47176 = ~controllable_hmaster1 & ~n47175;
  assign n47177 = ~controllable_hmaster1 & ~n47176;
  assign n47178 = i_hbusreq3 & ~n47177;
  assign n47179 = ~controllable_hmaster0 & ~n37991;
  assign n47180 = ~controllable_hmaster1 & ~n47179;
  assign n47181 = ~controllable_hmaster1 & ~n47180;
  assign n47182 = ~i_hbusreq3 & ~n47181;
  assign n47183 = ~n47178 & ~n47182;
  assign n47184 = ~controllable_hmaster2 & ~n47183;
  assign n47185 = ~controllable_hmaster2 & ~n47184;
  assign n47186 = ~controllable_hgrant3 & ~n47185;
  assign n47187 = ~n21304 & ~n47186;
  assign n47188 = controllable_nhgrant0 & ~n47187;
  assign n47189 = ~n21332 & ~n47188;
  assign n47190 = ~n3281 & ~n47189;
  assign n47191 = ~n3281 & ~n47190;
  assign n47192 = n3378 & ~n47191;
  assign n47193 = ~n21339 & ~n47184;
  assign n47194 = ~controllable_hgrant3 & ~n47193;
  assign n47195 = ~n21338 & ~n47194;
  assign n47196 = controllable_nhgrant0 & ~n47195;
  assign n47197 = ~n21347 & ~n47196;
  assign n47198 = ~n3281 & ~n47197;
  assign n47199 = ~n3950 & ~n47198;
  assign n47200 = ~n3378 & ~n47199;
  assign n47201 = ~n47192 & ~n47200;
  assign n47202 = n3492 & ~n47201;
  assign n47203 = ~n3493 & ~n47202;
  assign n47204 = n3485 & ~n47203;
  assign n47205 = ~n3486 & ~n47204;
  assign n47206 = ~n3476 & ~n47205;
  assign n47207 = ~n21383 & ~n47188;
  assign n47208 = ~n3281 & ~n47207;
  assign n47209 = ~n3281 & ~n47208;
  assign n47210 = n3378 & ~n47209;
  assign n47211 = ~controllable_hmaster0 & ~n39368;
  assign n47212 = ~n21412 & ~n47211;
  assign n47213 = ~controllable_hmaster1 & ~n47212;
  assign n47214 = ~n21411 & ~n47213;
  assign n47215 = i_hbusreq3 & ~n47214;
  assign n47216 = ~n6947 & ~n47079;
  assign n47217 = ~controllable_hmaster0 & ~n47216;
  assign n47218 = ~n21419 & ~n47217;
  assign n47219 = ~controllable_hmaster1 & ~n47218;
  assign n47220 = ~n21418 & ~n47219;
  assign n47221 = ~i_hbusreq3 & ~n47220;
  assign n47222 = ~n47215 & ~n47221;
  assign n47223 = ~controllable_hmaster2 & ~n47222;
  assign n47224 = ~n21410 & ~n47223;
  assign n47225 = ~controllable_hgrant3 & ~n47224;
  assign n47226 = ~n21338 & ~n47225;
  assign n47227 = controllable_nhgrant0 & ~n47226;
  assign n47228 = ~n21461 & ~n47227;
  assign n47229 = ~n3281 & ~n47228;
  assign n47230 = ~n4089 & ~n47229;
  assign n47231 = ~n3378 & ~n47230;
  assign n47232 = ~n47210 & ~n47231;
  assign n47233 = n3492 & ~n47232;
  assign n47234 = ~n21290 & ~n47233;
  assign n47235 = n3485 & ~n47234;
  assign n47236 = ~n21289 & ~n47235;
  assign n47237 = n3476 & ~n47236;
  assign n47238 = ~n47206 & ~n47237;
  assign n47239 = n3374 & ~n47238;
  assign n47240 = ~n21296 & ~n47239;
  assign n47241 = ~n3655 & ~n47240;
  assign n47242 = ~n47174 & ~n47241;
  assign n47243 = ~n3652 & ~n47242;
  assign n47244 = ~n47107 & ~n47243;
  assign n47245 = ~n3368 & ~n47244;
  assign n47246 = ~controllable_hmaster0 & ~n38150;
  assign n47247 = ~controllable_hmaster1 & ~n47246;
  assign n47248 = ~controllable_hmaster1 & ~n47247;
  assign n47249 = ~controllable_hmaster2 & ~n47248;
  assign n47250 = ~controllable_hmaster2 & ~n47249;
  assign n47251 = ~controllable_hgrant3 & ~n47250;
  assign n47252 = ~n21699 & ~n47251;
  assign n47253 = controllable_nhgrant0 & ~n47252;
  assign n47254 = ~n21712 & ~n47253;
  assign n47255 = ~n3281 & ~n47254;
  assign n47256 = ~n3281 & ~n47255;
  assign n47257 = n3492 & ~n47256;
  assign n47258 = n3492 & ~n47257;
  assign n47259 = n3485 & ~n47258;
  assign n47260 = n3485 & ~n47259;
  assign n47261 = ~n3476 & ~n47260;
  assign n47262 = ~n21740 & ~n47253;
  assign n47263 = ~n3281 & ~n47262;
  assign n47264 = ~n3281 & ~n47263;
  assign n47265 = n3492 & ~n47264;
  assign n47266 = ~n21722 & ~n47265;
  assign n47267 = n3485 & ~n47266;
  assign n47268 = ~n21721 & ~n47267;
  assign n47269 = n3476 & ~n47268;
  assign n47270 = ~n47261 & ~n47269;
  assign n47271 = n3374 & ~n47270;
  assign n47272 = n3374 & ~n47271;
  assign n47273 = n3655 & ~n47272;
  assign n47274 = ~controllable_hmaster0 & ~n38449;
  assign n47275 = ~controllable_hmaster1 & ~n47274;
  assign n47276 = ~controllable_hmaster1 & ~n47275;
  assign n47277 = ~controllable_hmaster2 & ~n47276;
  assign n47278 = ~controllable_hmaster2 & ~n47277;
  assign n47279 = ~controllable_hgrant3 & ~n47278;
  assign n47280 = ~n21699 & ~n47279;
  assign n47281 = controllable_nhgrant0 & ~n47280;
  assign n47282 = ~n21712 & ~n47281;
  assign n47283 = ~n3281 & ~n47282;
  assign n47284 = ~n3281 & ~n47283;
  assign n47285 = n3492 & ~n47284;
  assign n47286 = n3492 & ~n47285;
  assign n47287 = n3485 & ~n47286;
  assign n47288 = n3485 & ~n47287;
  assign n47289 = ~n3476 & ~n47288;
  assign n47290 = ~n21740 & ~n47281;
  assign n47291 = ~n3281 & ~n47290;
  assign n47292 = ~n3281 & ~n47291;
  assign n47293 = n3492 & ~n47292;
  assign n47294 = ~n21722 & ~n47293;
  assign n47295 = n3485 & ~n47294;
  assign n47296 = ~n21721 & ~n47295;
  assign n47297 = n3476 & ~n47296;
  assign n47298 = ~n47289 & ~n47297;
  assign n47299 = n3374 & ~n47298;
  assign n47300 = n3374 & ~n47299;
  assign n47301 = ~n3655 & ~n47300;
  assign n47302 = ~n47273 & ~n47301;
  assign n47303 = n3652 & ~n47302;
  assign n47304 = ~controllable_hmaster0 & ~n38728;
  assign n47305 = ~controllable_hmaster1 & ~n47304;
  assign n47306 = ~controllable_hmaster1 & ~n47305;
  assign n47307 = ~controllable_hmaster2 & ~n47306;
  assign n47308 = ~controllable_hmaster2 & ~n47307;
  assign n47309 = ~controllable_hgrant3 & ~n47308;
  assign n47310 = ~n21699 & ~n47309;
  assign n47311 = controllable_nhgrant0 & ~n47310;
  assign n47312 = ~n21712 & ~n47311;
  assign n47313 = ~n3281 & ~n47312;
  assign n47314 = ~n3281 & ~n47313;
  assign n47315 = n3492 & ~n47314;
  assign n47316 = n3492 & ~n47315;
  assign n47317 = n3485 & ~n47316;
  assign n47318 = n3485 & ~n47317;
  assign n47319 = ~n3476 & ~n47318;
  assign n47320 = ~n21740 & ~n47311;
  assign n47321 = ~n3281 & ~n47320;
  assign n47322 = ~n3281 & ~n47321;
  assign n47323 = n3492 & ~n47322;
  assign n47324 = ~n21722 & ~n47323;
  assign n47325 = n3485 & ~n47324;
  assign n47326 = ~n21721 & ~n47325;
  assign n47327 = n3476 & ~n47326;
  assign n47328 = ~n47319 & ~n47327;
  assign n47329 = n3374 & ~n47328;
  assign n47330 = n3374 & ~n47329;
  assign n47331 = n3655 & ~n47330;
  assign n47332 = ~controllable_hmaster0 & ~n38937;
  assign n47333 = ~controllable_hmaster1 & ~n47332;
  assign n47334 = ~controllable_hmaster1 & ~n47333;
  assign n47335 = ~controllable_hmaster2 & ~n47334;
  assign n47336 = ~controllable_hmaster2 & ~n47335;
  assign n47337 = ~controllable_hgrant3 & ~n47336;
  assign n47338 = ~n21699 & ~n47337;
  assign n47339 = controllable_nhgrant0 & ~n47338;
  assign n47340 = ~n21712 & ~n47339;
  assign n47341 = ~n3281 & ~n47340;
  assign n47342 = ~n3281 & ~n47341;
  assign n47343 = n3492 & ~n47342;
  assign n47344 = n3492 & ~n47343;
  assign n47345 = n3485 & ~n47344;
  assign n47346 = n3485 & ~n47345;
  assign n47347 = ~n3476 & ~n47346;
  assign n47348 = ~n21740 & ~n47339;
  assign n47349 = ~n3281 & ~n47348;
  assign n47350 = ~n3281 & ~n47349;
  assign n47351 = n3492 & ~n47350;
  assign n47352 = ~n21722 & ~n47351;
  assign n47353 = n3485 & ~n47352;
  assign n47354 = ~n21721 & ~n47353;
  assign n47355 = n3476 & ~n47354;
  assign n47356 = ~n47347 & ~n47355;
  assign n47357 = n3374 & ~n47356;
  assign n47358 = n3374 & ~n47357;
  assign n47359 = ~n3655 & ~n47358;
  assign n47360 = ~n47331 & ~n47359;
  assign n47361 = ~n3652 & ~n47360;
  assign n47362 = ~n47303 & ~n47361;
  assign n47363 = n3368 & ~n47362;
  assign n47364 = ~n47245 & ~n47363;
  assign n47365 = ~n3362 & ~n47364;
  assign n47366 = ~n3362 & ~n47365;
  assign n47367 = ~n3359 & ~n47366;
  assign n47368 = ~n3359 & ~n47367;
  assign n47369 = n3356 & ~n47368;
  assign n47370 = ~n34040 & ~n39564;
  assign n47371 = ~controllable_hmaster1 & ~n47370;
  assign n47372 = ~n39563 & ~n47371;
  assign n47373 = ~i_hbusreq3 & ~n47372;
  assign n47374 = ~n39568 & ~n47373;
  assign n47375 = controllable_hmaster2 & ~n47374;
  assign n47376 = ~n5161 & ~n47375;
  assign n47377 = ~controllable_hgrant3 & ~n47376;
  assign n47378 = ~n8750 & ~n47377;
  assign n47379 = controllable_nhgrant0 & ~n47378;
  assign n47380 = ~n8785 & ~n47379;
  assign n47381 = ~n3281 & ~n47380;
  assign n47382 = ~n3783 & ~n47381;
  assign n47383 = ~n3378 & ~n47382;
  assign n47384 = ~n21849 & ~n47383;
  assign n47385 = n3492 & ~n47384;
  assign n47386 = ~n3631 & ~n47385;
  assign n47387 = n3485 & ~n47386;
  assign n47388 = ~n3630 & ~n47387;
  assign n47389 = ~n3476 & ~n47388;
  assign n47390 = ~n8309 & ~n47385;
  assign n47391 = n3485 & ~n47390;
  assign n47392 = ~n8639 & ~n47391;
  assign n47393 = n3476 & ~n47392;
  assign n47394 = ~n47389 & ~n47393;
  assign n47395 = ~n3374 & ~n47394;
  assign n47396 = ~n5303 & ~n37430;
  assign n47397 = ~controllable_hmaster1 & ~n47396;
  assign n47398 = ~n5293 & ~n47397;
  assign n47399 = i_hbusreq3 & ~n47398;
  assign n47400 = ~n21911 & ~n37458;
  assign n47401 = ~controllable_hmaster1 & ~n47400;
  assign n47402 = ~n21897 & ~n47401;
  assign n47403 = ~i_hbusreq3 & ~n47402;
  assign n47404 = ~n47399 & ~n47403;
  assign n47405 = ~controllable_hmaster2 & ~n47404;
  assign n47406 = ~n21888 & ~n47405;
  assign n47407 = ~controllable_hgrant3 & ~n47406;
  assign n47408 = ~n8810 & ~n47407;
  assign n47409 = controllable_nhgrant0 & ~n47408;
  assign n47410 = ~n8902 & ~n47409;
  assign n47411 = ~n3281 & ~n47410;
  assign n47412 = ~n3950 & ~n47411;
  assign n47413 = n3378 & ~n47412;
  assign n47414 = ~n39619 & ~n39642;
  assign n47415 = ~controllable_hmaster1 & ~n47414;
  assign n47416 = ~n39618 & ~n47415;
  assign n47417 = ~i_hbusreq3 & ~n47416;
  assign n47418 = ~n39627 & ~n47417;
  assign n47419 = controllable_hmaster2 & ~n47418;
  assign n47420 = ~n35061 & ~n37430;
  assign n47421 = ~controllable_hmaster1 & ~n47420;
  assign n47422 = ~n35057 & ~n47421;
  assign n47423 = i_hbusreq3 & ~n47422;
  assign n47424 = ~n35084 & ~n37458;
  assign n47425 = ~controllable_hmaster1 & ~n47424;
  assign n47426 = ~n35076 & ~n47425;
  assign n47427 = ~i_hbusreq3 & ~n47426;
  assign n47428 = ~n47423 & ~n47427;
  assign n47429 = ~controllable_hmaster2 & ~n47428;
  assign n47430 = ~n47419 & ~n47429;
  assign n47431 = ~controllable_hgrant3 & ~n47430;
  assign n47432 = ~n8810 & ~n47431;
  assign n47433 = controllable_nhgrant0 & ~n47432;
  assign n47434 = ~n8902 & ~n47433;
  assign n47435 = ~n3281 & ~n47434;
  assign n47436 = ~n3950 & ~n47435;
  assign n47437 = ~n3378 & ~n47436;
  assign n47438 = ~n47413 & ~n47437;
  assign n47439 = n3492 & ~n47438;
  assign n47440 = ~n3631 & ~n47439;
  assign n47441 = n3485 & ~n47440;
  assign n47442 = ~n3630 & ~n47441;
  assign n47443 = ~n3476 & ~n47442;
  assign n47444 = ~controllable_hmaster0 & ~n39676;
  assign n47445 = ~n5701 & ~n47444;
  assign n47446 = ~controllable_hmaster1 & ~n47445;
  assign n47447 = ~n5690 & ~n47446;
  assign n47448 = i_hbusreq3 & ~n47447;
  assign n47449 = controllable_hgrant4 & ~n22378;
  assign n47450 = ~n9038 & ~n47449;
  assign n47451 = ~i_hbusreq2 & ~n47450;
  assign n47452 = ~n39682 & ~n47451;
  assign n47453 = ~controllable_hgrant2 & ~n47452;
  assign n47454 = ~n5981 & ~n47453;
  assign n47455 = ~controllable_hmaster0 & ~n47454;
  assign n47456 = ~n22007 & ~n47455;
  assign n47457 = ~controllable_hmaster1 & ~n47456;
  assign n47458 = ~n21991 & ~n47457;
  assign n47459 = ~i_hbusreq3 & ~n47458;
  assign n47460 = ~n47448 & ~n47459;
  assign n47461 = ~controllable_hmaster2 & ~n47460;
  assign n47462 = ~n21977 & ~n47461;
  assign n47463 = ~controllable_hgrant3 & ~n47462;
  assign n47464 = ~n8935 & ~n47463;
  assign n47465 = controllable_nhgrant0 & ~n47464;
  assign n47466 = ~n9096 & ~n47465;
  assign n47467 = ~n3281 & ~n47466;
  assign n47468 = ~n4089 & ~n47467;
  assign n47469 = n3378 & ~n47468;
  assign n47470 = controllable_hgrant4 & ~n22406;
  assign n47471 = ~n8950 & ~n47470;
  assign n47472 = ~i_hbusreq2 & ~n47471;
  assign n47473 = ~n37517 & ~n47472;
  assign n47474 = ~controllable_hgrant2 & ~n47473;
  assign n47475 = ~n8936 & ~n47474;
  assign n47476 = controllable_hmaster1 & ~n47475;
  assign n47477 = controllable_hmaster0 & ~n47475;
  assign n47478 = ~n22029 & ~n34214;
  assign n47479 = ~i_hbusreq2 & ~n47478;
  assign n47480 = ~n39720 & ~n47479;
  assign n47481 = ~controllable_hgrant2 & ~n47480;
  assign n47482 = ~n5862 & ~n47481;
  assign n47483 = ~controllable_hmaster0 & ~n47482;
  assign n47484 = ~n47477 & ~n47483;
  assign n47485 = ~controllable_hmaster1 & ~n47484;
  assign n47486 = ~n47476 & ~n47485;
  assign n47487 = ~i_hbusreq3 & ~n47486;
  assign n47488 = ~n39712 & ~n47487;
  assign n47489 = controllable_hmaster2 & ~n47488;
  assign n47490 = ~n35227 & ~n37512;
  assign n47491 = ~controllable_hmaster1 & ~n47490;
  assign n47492 = ~n35223 & ~n47491;
  assign n47493 = i_hbusreq3 & ~n47492;
  assign n47494 = ~n22029 & ~n35234;
  assign n47495 = ~i_hbusreq2 & ~n47494;
  assign n47496 = ~n35233 & ~n47495;
  assign n47497 = ~controllable_hgrant2 & ~n47496;
  assign n47498 = ~n5862 & ~n47497;
  assign n47499 = controllable_hmaster0 & ~n47498;
  assign n47500 = ~n5950 & ~n47497;
  assign n47501 = ~controllable_hmaster0 & ~n47500;
  assign n47502 = ~n47499 & ~n47501;
  assign n47503 = controllable_hmaster1 & ~n47502;
  assign n47504 = ~n22063 & ~n35234;
  assign n47505 = ~i_hbusreq2 & ~n47504;
  assign n47506 = ~n35245 & ~n47505;
  assign n47507 = ~controllable_hgrant2 & ~n47506;
  assign n47508 = ~n5862 & ~n47507;
  assign n47509 = controllable_hmaster0 & ~n47508;
  assign n47510 = ~n37540 & ~n47509;
  assign n47511 = ~controllable_hmaster1 & ~n47510;
  assign n47512 = ~n47503 & ~n47511;
  assign n47513 = ~i_hbusreq3 & ~n47512;
  assign n47514 = ~n47493 & ~n47513;
  assign n47515 = ~controllable_hmaster2 & ~n47514;
  assign n47516 = ~n47489 & ~n47515;
  assign n47517 = ~controllable_hgrant3 & ~n47516;
  assign n47518 = ~n8935 & ~n47517;
  assign n47519 = controllable_nhgrant0 & ~n47518;
  assign n47520 = ~n9096 & ~n47519;
  assign n47521 = ~n3281 & ~n47520;
  assign n47522 = ~n4089 & ~n47521;
  assign n47523 = ~n3378 & ~n47522;
  assign n47524 = ~n47469 & ~n47523;
  assign n47525 = n3492 & ~n47524;
  assign n47526 = ~n8309 & ~n47525;
  assign n47527 = n3485 & ~n47526;
  assign n47528 = ~n8639 & ~n47527;
  assign n47529 = n3476 & ~n47528;
  assign n47530 = ~n47443 & ~n47529;
  assign n47531 = n3374 & ~n47530;
  assign n47532 = ~n47395 & ~n47531;
  assign n47533 = n3655 & ~n47532;
  assign n47534 = ~n34040 & ~n39771;
  assign n47535 = ~controllable_hmaster1 & ~n47534;
  assign n47536 = ~n39770 & ~n47535;
  assign n47537 = ~i_hbusreq3 & ~n47536;
  assign n47538 = ~n39775 & ~n47537;
  assign n47539 = controllable_hmaster2 & ~n47538;
  assign n47540 = ~n6188 & ~n47539;
  assign n47541 = ~controllable_hgrant3 & ~n47540;
  assign n47542 = ~n8750 & ~n47541;
  assign n47543 = controllable_nhgrant0 & ~n47542;
  assign n47544 = ~n8785 & ~n47543;
  assign n47545 = ~n3281 & ~n47544;
  assign n47546 = ~n3783 & ~n47545;
  assign n47547 = ~n3378 & ~n47546;
  assign n47548 = ~n21849 & ~n47547;
  assign n47549 = n3492 & ~n47548;
  assign n47550 = ~n3631 & ~n47549;
  assign n47551 = n3485 & ~n47550;
  assign n47552 = ~n3630 & ~n47551;
  assign n47553 = ~n3476 & ~n47552;
  assign n47554 = ~n8309 & ~n47549;
  assign n47555 = n3485 & ~n47554;
  assign n47556 = ~n8639 & ~n47555;
  assign n47557 = n3476 & ~n47556;
  assign n47558 = ~n47553 & ~n47557;
  assign n47559 = ~n3374 & ~n47558;
  assign n47560 = ~n5303 & ~n37624;
  assign n47561 = ~controllable_hmaster1 & ~n47560;
  assign n47562 = ~n5293 & ~n47561;
  assign n47563 = i_hbusreq3 & ~n47562;
  assign n47564 = ~n21911 & ~n37652;
  assign n47565 = ~controllable_hmaster1 & ~n47564;
  assign n47566 = ~n21897 & ~n47565;
  assign n47567 = ~i_hbusreq3 & ~n47566;
  assign n47568 = ~n47563 & ~n47567;
  assign n47569 = ~controllable_hmaster2 & ~n47568;
  assign n47570 = ~n21888 & ~n47569;
  assign n47571 = ~controllable_hgrant3 & ~n47570;
  assign n47572 = ~n8810 & ~n47571;
  assign n47573 = controllable_nhgrant0 & ~n47572;
  assign n47574 = ~n8902 & ~n47573;
  assign n47575 = ~n3281 & ~n47574;
  assign n47576 = ~n3950 & ~n47575;
  assign n47577 = n3378 & ~n47576;
  assign n47578 = ~n39826 & ~n39849;
  assign n47579 = ~controllable_hmaster1 & ~n47578;
  assign n47580 = ~n39825 & ~n47579;
  assign n47581 = ~i_hbusreq3 & ~n47580;
  assign n47582 = ~n39834 & ~n47581;
  assign n47583 = controllable_hmaster2 & ~n47582;
  assign n47584 = ~n35368 & ~n37624;
  assign n47585 = ~controllable_hmaster1 & ~n47584;
  assign n47586 = ~n35364 & ~n47585;
  assign n47587 = i_hbusreq3 & ~n47586;
  assign n47588 = ~n35391 & ~n37652;
  assign n47589 = ~controllable_hmaster1 & ~n47588;
  assign n47590 = ~n35384 & ~n47589;
  assign n47591 = ~i_hbusreq3 & ~n47590;
  assign n47592 = ~n47587 & ~n47591;
  assign n47593 = ~controllable_hmaster2 & ~n47592;
  assign n47594 = ~n47583 & ~n47593;
  assign n47595 = ~controllable_hgrant3 & ~n47594;
  assign n47596 = ~n8810 & ~n47595;
  assign n47597 = controllable_nhgrant0 & ~n47596;
  assign n47598 = ~n8902 & ~n47597;
  assign n47599 = ~n3281 & ~n47598;
  assign n47600 = ~n3950 & ~n47599;
  assign n47601 = ~n3378 & ~n47600;
  assign n47602 = ~n47577 & ~n47601;
  assign n47603 = n3492 & ~n47602;
  assign n47604 = ~n3631 & ~n47603;
  assign n47605 = n3485 & ~n47604;
  assign n47606 = ~n3630 & ~n47605;
  assign n47607 = ~n3476 & ~n47606;
  assign n47608 = ~controllable_hmaster0 & ~n39882;
  assign n47609 = ~n5701 & ~n47608;
  assign n47610 = ~controllable_hmaster1 & ~n47609;
  assign n47611 = ~n5690 & ~n47610;
  assign n47612 = i_hbusreq3 & ~n47611;
  assign n47613 = ~n22182 & ~n47449;
  assign n47614 = ~i_hbusreq2 & ~n47613;
  assign n47615 = ~n39888 & ~n47614;
  assign n47616 = ~controllable_hgrant2 & ~n47615;
  assign n47617 = ~n5981 & ~n47616;
  assign n47618 = ~controllable_hmaster0 & ~n47617;
  assign n47619 = ~n22007 & ~n47618;
  assign n47620 = ~controllable_hmaster1 & ~n47619;
  assign n47621 = ~n21991 & ~n47620;
  assign n47622 = ~i_hbusreq3 & ~n47621;
  assign n47623 = ~n47612 & ~n47622;
  assign n47624 = ~controllable_hmaster2 & ~n47623;
  assign n47625 = ~n21977 & ~n47624;
  assign n47626 = ~controllable_hgrant3 & ~n47625;
  assign n47627 = ~n8935 & ~n47626;
  assign n47628 = controllable_nhgrant0 & ~n47627;
  assign n47629 = ~n9096 & ~n47628;
  assign n47630 = ~n3281 & ~n47629;
  assign n47631 = ~n4089 & ~n47630;
  assign n47632 = n3378 & ~n47631;
  assign n47633 = ~n22210 & ~n47470;
  assign n47634 = ~i_hbusreq2 & ~n47633;
  assign n47635 = ~n37720 & ~n47634;
  assign n47636 = ~controllable_hgrant2 & ~n47635;
  assign n47637 = ~n8936 & ~n47636;
  assign n47638 = controllable_hmaster1 & ~n47637;
  assign n47639 = controllable_hmaster0 & ~n47637;
  assign n47640 = ~n22225 & ~n34214;
  assign n47641 = ~i_hbusreq2 & ~n47640;
  assign n47642 = ~n39925 & ~n47641;
  assign n47643 = ~controllable_hgrant2 & ~n47642;
  assign n47644 = ~n5862 & ~n47643;
  assign n47645 = ~controllable_hmaster0 & ~n47644;
  assign n47646 = ~n47639 & ~n47645;
  assign n47647 = ~controllable_hmaster1 & ~n47646;
  assign n47648 = ~n47638 & ~n47647;
  assign n47649 = ~i_hbusreq3 & ~n47648;
  assign n47650 = ~n39917 & ~n47649;
  assign n47651 = controllable_hmaster2 & ~n47650;
  assign n47652 = ~n35493 & ~n37715;
  assign n47653 = ~controllable_hmaster1 & ~n47652;
  assign n47654 = ~n35489 & ~n47653;
  assign n47655 = i_hbusreq3 & ~n47654;
  assign n47656 = ~n22225 & ~n35234;
  assign n47657 = ~i_hbusreq2 & ~n47656;
  assign n47658 = ~n35499 & ~n47657;
  assign n47659 = ~controllable_hgrant2 & ~n47658;
  assign n47660 = ~n5862 & ~n47659;
  assign n47661 = controllable_hmaster0 & ~n47660;
  assign n47662 = ~n5950 & ~n47659;
  assign n47663 = ~controllable_hmaster0 & ~n47662;
  assign n47664 = ~n47661 & ~n47663;
  assign n47665 = controllable_hmaster1 & ~n47664;
  assign n47666 = ~n22259 & ~n35234;
  assign n47667 = ~i_hbusreq2 & ~n47666;
  assign n47668 = ~n35510 & ~n47667;
  assign n47669 = ~controllable_hgrant2 & ~n47668;
  assign n47670 = ~n5862 & ~n47669;
  assign n47671 = controllable_hmaster0 & ~n47670;
  assign n47672 = ~n37743 & ~n47671;
  assign n47673 = ~controllable_hmaster1 & ~n47672;
  assign n47674 = ~n47665 & ~n47673;
  assign n47675 = ~i_hbusreq3 & ~n47674;
  assign n47676 = ~n47655 & ~n47675;
  assign n47677 = ~controllable_hmaster2 & ~n47676;
  assign n47678 = ~n47651 & ~n47677;
  assign n47679 = ~controllable_hgrant3 & ~n47678;
  assign n47680 = ~n8935 & ~n47679;
  assign n47681 = controllable_nhgrant0 & ~n47680;
  assign n47682 = ~n9096 & ~n47681;
  assign n47683 = ~n3281 & ~n47682;
  assign n47684 = ~n4089 & ~n47683;
  assign n47685 = ~n3378 & ~n47684;
  assign n47686 = ~n47632 & ~n47685;
  assign n47687 = n3492 & ~n47686;
  assign n47688 = ~n8309 & ~n47687;
  assign n47689 = n3485 & ~n47688;
  assign n47690 = ~n8639 & ~n47689;
  assign n47691 = n3476 & ~n47690;
  assign n47692 = ~n47607 & ~n47691;
  assign n47693 = n3374 & ~n47692;
  assign n47694 = ~n47559 & ~n47693;
  assign n47695 = ~n3655 & ~n47694;
  assign n47696 = ~n47533 & ~n47695;
  assign n47697 = n3652 & ~n47696;
  assign n47698 = ~n34040 & ~n39976;
  assign n47699 = ~controllable_hmaster1 & ~n47698;
  assign n47700 = ~n39975 & ~n47699;
  assign n47701 = ~i_hbusreq3 & ~n47700;
  assign n47702 = ~n39980 & ~n47701;
  assign n47703 = controllable_hmaster2 & ~n47702;
  assign n47704 = ~n6657 & ~n47703;
  assign n47705 = ~controllable_hgrant3 & ~n47704;
  assign n47706 = ~n8750 & ~n47705;
  assign n47707 = controllable_nhgrant0 & ~n47706;
  assign n47708 = ~n8785 & ~n47707;
  assign n47709 = ~n3281 & ~n47708;
  assign n47710 = ~n3783 & ~n47709;
  assign n47711 = ~n3378 & ~n47710;
  assign n47712 = ~n21849 & ~n47711;
  assign n47713 = n3492 & ~n47712;
  assign n47714 = ~n3631 & ~n47713;
  assign n47715 = n3485 & ~n47714;
  assign n47716 = ~n3630 & ~n47715;
  assign n47717 = ~n3476 & ~n47716;
  assign n47718 = ~n8309 & ~n47713;
  assign n47719 = n3485 & ~n47718;
  assign n47720 = ~n8639 & ~n47719;
  assign n47721 = n3476 & ~n47720;
  assign n47722 = ~n47717 & ~n47721;
  assign n47723 = ~n3374 & ~n47722;
  assign n47724 = ~n5303 & ~n37823;
  assign n47725 = ~controllable_hmaster1 & ~n47724;
  assign n47726 = ~n5293 & ~n47725;
  assign n47727 = i_hbusreq3 & ~n47726;
  assign n47728 = ~n21911 & ~n37837;
  assign n47729 = ~controllable_hmaster1 & ~n47728;
  assign n47730 = ~n21897 & ~n47729;
  assign n47731 = ~i_hbusreq3 & ~n47730;
  assign n47732 = ~n47727 & ~n47731;
  assign n47733 = ~controllable_hmaster2 & ~n47732;
  assign n47734 = ~n21888 & ~n47733;
  assign n47735 = ~controllable_hgrant3 & ~n47734;
  assign n47736 = ~n8810 & ~n47735;
  assign n47737 = controllable_nhgrant0 & ~n47736;
  assign n47738 = ~n8902 & ~n47737;
  assign n47739 = ~n3281 & ~n47738;
  assign n47740 = ~n3950 & ~n47739;
  assign n47741 = n3378 & ~n47740;
  assign n47742 = ~n40024 & ~n40035;
  assign n47743 = ~controllable_hmaster1 & ~n47742;
  assign n47744 = ~n40023 & ~n47743;
  assign n47745 = ~i_hbusreq3 & ~n47744;
  assign n47746 = ~n40030 & ~n47745;
  assign n47747 = controllable_hmaster2 & ~n47746;
  assign n47748 = ~n35616 & ~n37823;
  assign n47749 = ~controllable_hmaster1 & ~n47748;
  assign n47750 = ~n35614 & ~n47749;
  assign n47751 = i_hbusreq3 & ~n47750;
  assign n47752 = ~n35629 & ~n37837;
  assign n47753 = ~controllable_hmaster1 & ~n47752;
  assign n47754 = ~n35627 & ~n47753;
  assign n47755 = ~i_hbusreq3 & ~n47754;
  assign n47756 = ~n47751 & ~n47755;
  assign n47757 = ~controllable_hmaster2 & ~n47756;
  assign n47758 = ~n47747 & ~n47757;
  assign n47759 = ~controllable_hgrant3 & ~n47758;
  assign n47760 = ~n8810 & ~n47759;
  assign n47761 = controllable_nhgrant0 & ~n47760;
  assign n47762 = ~n8902 & ~n47761;
  assign n47763 = ~n3281 & ~n47762;
  assign n47764 = ~n3950 & ~n47763;
  assign n47765 = ~n3378 & ~n47764;
  assign n47766 = ~n47741 & ~n47765;
  assign n47767 = n3492 & ~n47766;
  assign n47768 = ~n3631 & ~n47767;
  assign n47769 = n3485 & ~n47768;
  assign n47770 = ~n3630 & ~n47769;
  assign n47771 = ~n3476 & ~n47770;
  assign n47772 = ~controllable_hmaster0 & ~n40066;
  assign n47773 = ~n5701 & ~n47772;
  assign n47774 = ~controllable_hmaster1 & ~n47773;
  assign n47775 = ~n5690 & ~n47774;
  assign n47776 = i_hbusreq3 & ~n47775;
  assign n47777 = ~n22383 & ~n47453;
  assign n47778 = ~controllable_hmaster0 & ~n47777;
  assign n47779 = ~n22007 & ~n47778;
  assign n47780 = ~controllable_hmaster1 & ~n47779;
  assign n47781 = ~n21991 & ~n47780;
  assign n47782 = ~i_hbusreq3 & ~n47781;
  assign n47783 = ~n47776 & ~n47782;
  assign n47784 = ~controllable_hmaster2 & ~n47783;
  assign n47785 = ~n21977 & ~n47784;
  assign n47786 = ~controllable_hgrant3 & ~n47785;
  assign n47787 = ~n8935 & ~n47786;
  assign n47788 = controllable_nhgrant0 & ~n47787;
  assign n47789 = ~n9096 & ~n47788;
  assign n47790 = ~n3281 & ~n47789;
  assign n47791 = ~n4089 & ~n47790;
  assign n47792 = n3378 & ~n47791;
  assign n47793 = ~n22411 & ~n47474;
  assign n47794 = controllable_hmaster1 & ~n47793;
  assign n47795 = controllable_hmaster0 & ~n47793;
  assign n47796 = ~n6772 & ~n47481;
  assign n47797 = ~controllable_hmaster0 & ~n47796;
  assign n47798 = ~n47795 & ~n47797;
  assign n47799 = ~controllable_hmaster1 & ~n47798;
  assign n47800 = ~n47794 & ~n47799;
  assign n47801 = ~i_hbusreq3 & ~n47800;
  assign n47802 = ~n40094 & ~n47801;
  assign n47803 = controllable_hmaster2 & ~n47802;
  assign n47804 = ~n35701 & ~n37885;
  assign n47805 = ~controllable_hmaster1 & ~n47804;
  assign n47806 = ~n35699 & ~n47805;
  assign n47807 = i_hbusreq3 & ~n47806;
  assign n47808 = ~n6772 & ~n47497;
  assign n47809 = controllable_hmaster0 & ~n47808;
  assign n47810 = ~n6813 & ~n47497;
  assign n47811 = ~controllable_hmaster0 & ~n47810;
  assign n47812 = ~n47809 & ~n47811;
  assign n47813 = controllable_hmaster1 & ~n47812;
  assign n47814 = ~n6772 & ~n47507;
  assign n47815 = controllable_hmaster0 & ~n47814;
  assign n47816 = ~n37899 & ~n47815;
  assign n47817 = ~controllable_hmaster1 & ~n47816;
  assign n47818 = ~n47813 & ~n47817;
  assign n47819 = ~i_hbusreq3 & ~n47818;
  assign n47820 = ~n47807 & ~n47819;
  assign n47821 = ~controllable_hmaster2 & ~n47820;
  assign n47822 = ~n47803 & ~n47821;
  assign n47823 = ~controllable_hgrant3 & ~n47822;
  assign n47824 = ~n8935 & ~n47823;
  assign n47825 = controllable_nhgrant0 & ~n47824;
  assign n47826 = ~n9096 & ~n47825;
  assign n47827 = ~n3281 & ~n47826;
  assign n47828 = ~n4089 & ~n47827;
  assign n47829 = ~n3378 & ~n47828;
  assign n47830 = ~n47792 & ~n47829;
  assign n47831 = n3492 & ~n47830;
  assign n47832 = ~n8309 & ~n47831;
  assign n47833 = n3485 & ~n47832;
  assign n47834 = ~n8639 & ~n47833;
  assign n47835 = n3476 & ~n47834;
  assign n47836 = ~n47771 & ~n47835;
  assign n47837 = n3374 & ~n47836;
  assign n47838 = ~n47723 & ~n47837;
  assign n47839 = n3655 & ~n47838;
  assign n47840 = ~n34040 & ~n40138;
  assign n47841 = ~controllable_hmaster1 & ~n47840;
  assign n47842 = ~n40137 & ~n47841;
  assign n47843 = ~i_hbusreq3 & ~n47842;
  assign n47844 = ~n40142 & ~n47843;
  assign n47845 = controllable_hmaster2 & ~n47844;
  assign n47846 = ~n6887 & ~n47845;
  assign n47847 = ~controllable_hgrant3 & ~n47846;
  assign n47848 = ~n8750 & ~n47847;
  assign n47849 = controllable_nhgrant0 & ~n47848;
  assign n47850 = ~n8785 & ~n47849;
  assign n47851 = ~n3281 & ~n47850;
  assign n47852 = ~n3783 & ~n47851;
  assign n47853 = ~n3378 & ~n47852;
  assign n47854 = ~n21849 & ~n47853;
  assign n47855 = n3492 & ~n47854;
  assign n47856 = ~n3631 & ~n47855;
  assign n47857 = n3485 & ~n47856;
  assign n47858 = ~n3630 & ~n47857;
  assign n47859 = ~n3476 & ~n47858;
  assign n47860 = ~n8309 & ~n47855;
  assign n47861 = n3485 & ~n47860;
  assign n47862 = ~n8639 & ~n47861;
  assign n47863 = n3476 & ~n47862;
  assign n47864 = ~n47859 & ~n47863;
  assign n47865 = ~n3374 & ~n47864;
  assign n47866 = ~n5303 & ~n37977;
  assign n47867 = ~controllable_hmaster1 & ~n47866;
  assign n47868 = ~n5293 & ~n47867;
  assign n47869 = i_hbusreq3 & ~n47868;
  assign n47870 = ~n21911 & ~n37991;
  assign n47871 = ~controllable_hmaster1 & ~n47870;
  assign n47872 = ~n21897 & ~n47871;
  assign n47873 = ~i_hbusreq3 & ~n47872;
  assign n47874 = ~n47869 & ~n47873;
  assign n47875 = ~controllable_hmaster2 & ~n47874;
  assign n47876 = ~n21888 & ~n47875;
  assign n47877 = ~controllable_hgrant3 & ~n47876;
  assign n47878 = ~n8810 & ~n47877;
  assign n47879 = controllable_nhgrant0 & ~n47878;
  assign n47880 = ~n8902 & ~n47879;
  assign n47881 = ~n3281 & ~n47880;
  assign n47882 = ~n3950 & ~n47881;
  assign n47883 = n3378 & ~n47882;
  assign n47884 = ~n40186 & ~n40197;
  assign n47885 = ~controllable_hmaster1 & ~n47884;
  assign n47886 = ~n40185 & ~n47885;
  assign n47887 = ~i_hbusreq3 & ~n47886;
  assign n47888 = ~n40192 & ~n47887;
  assign n47889 = controllable_hmaster2 & ~n47888;
  assign n47890 = ~n35808 & ~n37977;
  assign n47891 = ~controllable_hmaster1 & ~n47890;
  assign n47892 = ~n35806 & ~n47891;
  assign n47893 = i_hbusreq3 & ~n47892;
  assign n47894 = ~n35821 & ~n37991;
  assign n47895 = ~controllable_hmaster1 & ~n47894;
  assign n47896 = ~n35819 & ~n47895;
  assign n47897 = ~i_hbusreq3 & ~n47896;
  assign n47898 = ~n47893 & ~n47897;
  assign n47899 = ~controllable_hmaster2 & ~n47898;
  assign n47900 = ~n47889 & ~n47899;
  assign n47901 = ~controllable_hgrant3 & ~n47900;
  assign n47902 = ~n8810 & ~n47901;
  assign n47903 = controllable_nhgrant0 & ~n47902;
  assign n47904 = ~n8902 & ~n47903;
  assign n47905 = ~n3281 & ~n47904;
  assign n47906 = ~n3950 & ~n47905;
  assign n47907 = ~n3378 & ~n47906;
  assign n47908 = ~n47883 & ~n47907;
  assign n47909 = n3492 & ~n47908;
  assign n47910 = ~n3631 & ~n47909;
  assign n47911 = n3485 & ~n47910;
  assign n47912 = ~n3630 & ~n47911;
  assign n47913 = ~n3476 & ~n47912;
  assign n47914 = ~controllable_hmaster0 & ~n40228;
  assign n47915 = ~n5701 & ~n47914;
  assign n47916 = ~controllable_hmaster1 & ~n47915;
  assign n47917 = ~n5690 & ~n47916;
  assign n47918 = i_hbusreq3 & ~n47917;
  assign n47919 = ~n22383 & ~n47616;
  assign n47920 = ~controllable_hmaster0 & ~n47919;
  assign n47921 = ~n22007 & ~n47920;
  assign n47922 = ~controllable_hmaster1 & ~n47921;
  assign n47923 = ~n21991 & ~n47922;
  assign n47924 = ~i_hbusreq3 & ~n47923;
  assign n47925 = ~n47918 & ~n47924;
  assign n47926 = ~controllable_hmaster2 & ~n47925;
  assign n47927 = ~n21977 & ~n47926;
  assign n47928 = ~controllable_hgrant3 & ~n47927;
  assign n47929 = ~n8935 & ~n47928;
  assign n47930 = controllable_nhgrant0 & ~n47929;
  assign n47931 = ~n9096 & ~n47930;
  assign n47932 = ~n3281 & ~n47931;
  assign n47933 = ~n4089 & ~n47932;
  assign n47934 = n3378 & ~n47933;
  assign n47935 = ~n22411 & ~n47636;
  assign n47936 = controllable_hmaster1 & ~n47935;
  assign n47937 = controllable_hmaster0 & ~n47935;
  assign n47938 = ~n6772 & ~n47643;
  assign n47939 = ~controllable_hmaster0 & ~n47938;
  assign n47940 = ~n47937 & ~n47939;
  assign n47941 = ~controllable_hmaster1 & ~n47940;
  assign n47942 = ~n47936 & ~n47941;
  assign n47943 = ~i_hbusreq3 & ~n47942;
  assign n47944 = ~n40256 & ~n47943;
  assign n47945 = controllable_hmaster2 & ~n47944;
  assign n47946 = ~n35893 & ~n38039;
  assign n47947 = ~controllable_hmaster1 & ~n47946;
  assign n47948 = ~n35891 & ~n47947;
  assign n47949 = i_hbusreq3 & ~n47948;
  assign n47950 = ~n6772 & ~n47659;
  assign n47951 = controllable_hmaster0 & ~n47950;
  assign n47952 = ~n6813 & ~n47659;
  assign n47953 = ~controllable_hmaster0 & ~n47952;
  assign n47954 = ~n47951 & ~n47953;
  assign n47955 = controllable_hmaster1 & ~n47954;
  assign n47956 = ~n6772 & ~n47669;
  assign n47957 = controllable_hmaster0 & ~n47956;
  assign n47958 = ~n38053 & ~n47957;
  assign n47959 = ~controllable_hmaster1 & ~n47958;
  assign n47960 = ~n47955 & ~n47959;
  assign n47961 = ~i_hbusreq3 & ~n47960;
  assign n47962 = ~n47949 & ~n47961;
  assign n47963 = ~controllable_hmaster2 & ~n47962;
  assign n47964 = ~n47945 & ~n47963;
  assign n47965 = ~controllable_hgrant3 & ~n47964;
  assign n47966 = ~n8935 & ~n47965;
  assign n47967 = controllable_nhgrant0 & ~n47966;
  assign n47968 = ~n9096 & ~n47967;
  assign n47969 = ~n3281 & ~n47968;
  assign n47970 = ~n4089 & ~n47969;
  assign n47971 = ~n3378 & ~n47970;
  assign n47972 = ~n47934 & ~n47971;
  assign n47973 = n3492 & ~n47972;
  assign n47974 = ~n8309 & ~n47973;
  assign n47975 = n3485 & ~n47974;
  assign n47976 = ~n8639 & ~n47975;
  assign n47977 = n3476 & ~n47976;
  assign n47978 = ~n47913 & ~n47977;
  assign n47979 = n3374 & ~n47978;
  assign n47980 = ~n47865 & ~n47979;
  assign n47981 = ~n3655 & ~n47980;
  assign n47982 = ~n47839 & ~n47981;
  assign n47983 = ~n3652 & ~n47982;
  assign n47984 = ~n47697 & ~n47983;
  assign n47985 = ~n3368 & ~n47984;
  assign n47986 = controllable_hgrant4 & ~n22710;
  assign n47987 = ~n22628 & ~n47986;
  assign n47988 = ~i_hbusreq2 & ~n47987;
  assign n47989 = ~n39569 & ~n47988;
  assign n47990 = ~controllable_hgrant2 & ~n47989;
  assign n47991 = ~n4562 & ~n47990;
  assign n47992 = controllable_hmaster1 & ~n47991;
  assign n47993 = controllable_hmaster0 & ~n47991;
  assign n47994 = controllable_hmaster0 & ~n47993;
  assign n47995 = ~controllable_hmaster1 & ~n47994;
  assign n47996 = ~n47992 & ~n47995;
  assign n47997 = ~i_hbusreq3 & ~n47996;
  assign n47998 = ~n40305 & ~n47997;
  assign n47999 = controllable_hmaster2 & ~n47998;
  assign n48000 = controllable_hmaster2 & ~n47999;
  assign n48001 = ~controllable_hgrant3 & ~n48000;
  assign n48002 = ~n9708 & ~n48001;
  assign n48003 = controllable_nhgrant0 & ~n48002;
  assign n48004 = ~n9753 & ~n48003;
  assign n48005 = ~n3281 & ~n48004;
  assign n48006 = ~n3281 & ~n48005;
  assign n48007 = ~n3378 & ~n48006;
  assign n48008 = ~n22618 & ~n48007;
  assign n48009 = n3492 & ~n48008;
  assign n48010 = n3492 & ~n48009;
  assign n48011 = n3485 & ~n48010;
  assign n48012 = n3485 & ~n48011;
  assign n48013 = ~n3374 & ~n48012;
  assign n48014 = ~n5303 & ~n38150;
  assign n48015 = ~controllable_hmaster1 & ~n48014;
  assign n48016 = ~n5293 & ~n48015;
  assign n48017 = i_hbusreq3 & ~n48016;
  assign n48018 = ~n22687 & ~n38150;
  assign n48019 = ~controllable_hmaster1 & ~n48018;
  assign n48020 = ~n22673 & ~n48019;
  assign n48021 = ~i_hbusreq3 & ~n48020;
  assign n48022 = ~n48017 & ~n48021;
  assign n48023 = ~controllable_hmaster2 & ~n48022;
  assign n48024 = ~n22668 & ~n48023;
  assign n48025 = ~controllable_hgrant3 & ~n48024;
  assign n48026 = ~n9790 & ~n48025;
  assign n48027 = controllable_nhgrant0 & ~n48026;
  assign n48028 = ~n9861 & ~n48027;
  assign n48029 = ~n3281 & ~n48028;
  assign n48030 = ~n3281 & ~n48029;
  assign n48031 = n3378 & ~n48030;
  assign n48032 = controllable_hgrant4 & ~n22627;
  assign n48033 = ~n22711 & ~n48032;
  assign n48034 = ~i_hbusreq2 & ~n48033;
  assign n48035 = ~n39636 & ~n48034;
  assign n48036 = ~controllable_hgrant2 & ~n48035;
  assign n48037 = ~n4562 & ~n48036;
  assign n48038 = ~controllable_hmaster0 & ~n48037;
  assign n48039 = ~n47993 & ~n48038;
  assign n48040 = ~controllable_hmaster1 & ~n48039;
  assign n48041 = ~n47992 & ~n48040;
  assign n48042 = ~i_hbusreq3 & ~n48041;
  assign n48043 = ~n40347 & ~n48042;
  assign n48044 = controllable_hmaster2 & ~n48043;
  assign n48045 = ~n35061 & ~n38150;
  assign n48046 = ~controllable_hmaster1 & ~n48045;
  assign n48047 = ~n35057 & ~n48046;
  assign n48048 = i_hbusreq3 & ~n48047;
  assign n48049 = ~i_hbusreq2 & ~n22710;
  assign n48050 = ~n35067 & ~n48049;
  assign n48051 = ~controllable_hgrant2 & ~n48050;
  assign n48052 = ~n4562 & ~n48051;
  assign n48053 = controllable_hmaster0 & ~n48052;
  assign n48054 = ~n9803 & ~n48051;
  assign n48055 = ~controllable_hmaster0 & ~n48054;
  assign n48056 = ~n48053 & ~n48055;
  assign n48057 = controllable_hmaster1 & ~n48056;
  assign n48058 = ~n22741 & ~n47986;
  assign n48059 = ~i_hbusreq2 & ~n48058;
  assign n48060 = ~n35077 & ~n48059;
  assign n48061 = ~controllable_hgrant2 & ~n48060;
  assign n48062 = ~n4562 & ~n48061;
  assign n48063 = controllable_hmaster0 & ~n48062;
  assign n48064 = ~n38150 & ~n48063;
  assign n48065 = ~controllable_hmaster1 & ~n48064;
  assign n48066 = ~n48057 & ~n48065;
  assign n48067 = ~i_hbusreq3 & ~n48066;
  assign n48068 = ~n48048 & ~n48067;
  assign n48069 = ~controllable_hmaster2 & ~n48068;
  assign n48070 = ~n48044 & ~n48069;
  assign n48071 = ~controllable_hgrant3 & ~n48070;
  assign n48072 = ~n9790 & ~n48071;
  assign n48073 = controllable_nhgrant0 & ~n48072;
  assign n48074 = ~n9861 & ~n48073;
  assign n48075 = ~n3281 & ~n48074;
  assign n48076 = ~n3281 & ~n48075;
  assign n48077 = ~n3378 & ~n48076;
  assign n48078 = ~n48031 & ~n48077;
  assign n48079 = n3492 & ~n48078;
  assign n48080 = n3492 & ~n48079;
  assign n48081 = n3485 & ~n48080;
  assign n48082 = n3485 & ~n48081;
  assign n48083 = ~n3476 & ~n48082;
  assign n48084 = ~controllable_hmaster0 & ~n40381;
  assign n48085 = ~n7339 & ~n48084;
  assign n48086 = ~controllable_hmaster1 & ~n48085;
  assign n48087 = ~n7330 & ~n48086;
  assign n48088 = i_hbusreq3 & ~n48087;
  assign n48089 = ~n22842 & ~n48084;
  assign n48090 = ~controllable_hmaster1 & ~n48089;
  assign n48091 = ~n22823 & ~n48090;
  assign n48092 = ~i_hbusreq3 & ~n48091;
  assign n48093 = ~n48088 & ~n48092;
  assign n48094 = ~controllable_hmaster2 & ~n48093;
  assign n48095 = ~n22808 & ~n48094;
  assign n48096 = ~controllable_hgrant3 & ~n48095;
  assign n48097 = ~n10110 & ~n48096;
  assign n48098 = controllable_nhgrant0 & ~n48097;
  assign n48099 = ~n10240 & ~n48098;
  assign n48100 = ~n3281 & ~n48099;
  assign n48101 = ~n3281 & ~n48100;
  assign n48102 = n3378 & ~n48101;
  assign n48103 = controllable_hgrant4 & ~n23297;
  assign n48104 = ~n22866 & ~n48103;
  assign n48105 = ~i_hbusreq2 & ~n48104;
  assign n48106 = ~n40422 & ~n48105;
  assign n48107 = ~controllable_hgrant2 & ~n48106;
  assign n48108 = ~n10111 & ~n48107;
  assign n48109 = controllable_hmaster1 & ~n48108;
  assign n48110 = controllable_hmaster0 & ~n48108;
  assign n48111 = controllable_hgrant4 & ~n23329;
  assign n48112 = ~n22881 & ~n48111;
  assign n48113 = ~i_hbusreq2 & ~n48112;
  assign n48114 = ~n40430 & ~n48113;
  assign n48115 = ~controllable_hgrant2 & ~n48114;
  assign n48116 = ~n10111 & ~n48115;
  assign n48117 = ~controllable_hmaster0 & ~n48116;
  assign n48118 = ~n48110 & ~n48117;
  assign n48119 = ~controllable_hmaster1 & ~n48118;
  assign n48120 = ~n48109 & ~n48119;
  assign n48121 = ~i_hbusreq3 & ~n48120;
  assign n48122 = ~n40421 & ~n48121;
  assign n48123 = controllable_hmaster2 & ~n48122;
  assign n48124 = ~controllable_hmaster0 & ~n40446;
  assign n48125 = ~n40457 & ~n48124;
  assign n48126 = ~controllable_hmaster1 & ~n48125;
  assign n48127 = ~n45630 & ~n48126;
  assign n48128 = i_hbusreq3 & ~n48127;
  assign n48129 = ~n22881 & ~n48103;
  assign n48130 = ~i_hbusreq2 & ~n48129;
  assign n48131 = ~n40472 & ~n48130;
  assign n48132 = ~controllable_hgrant2 & ~n48131;
  assign n48133 = ~n10111 & ~n48132;
  assign n48134 = controllable_hmaster0 & ~n48133;
  assign n48135 = ~n10152 & ~n48132;
  assign n48136 = ~controllable_hmaster0 & ~n48135;
  assign n48137 = ~n48134 & ~n48136;
  assign n48138 = controllable_hmaster1 & ~n48137;
  assign n48139 = ~n22918 & ~n48103;
  assign n48140 = ~i_hbusreq2 & ~n48139;
  assign n48141 = ~n40481 & ~n48140;
  assign n48142 = ~controllable_hgrant2 & ~n48141;
  assign n48143 = ~n10111 & ~n48142;
  assign n48144 = controllable_hmaster0 & ~n48143;
  assign n48145 = ~n48124 & ~n48144;
  assign n48146 = ~controllable_hmaster1 & ~n48145;
  assign n48147 = ~n48138 & ~n48146;
  assign n48148 = ~i_hbusreq3 & ~n48147;
  assign n48149 = ~n48128 & ~n48148;
  assign n48150 = ~controllable_hmaster2 & ~n48149;
  assign n48151 = ~n48123 & ~n48150;
  assign n48152 = ~controllable_hgrant3 & ~n48151;
  assign n48153 = ~n10110 & ~n48152;
  assign n48154 = controllable_nhgrant0 & ~n48153;
  assign n48155 = ~n10240 & ~n48154;
  assign n48156 = ~n3281 & ~n48155;
  assign n48157 = ~n3281 & ~n48156;
  assign n48158 = ~n3378 & ~n48157;
  assign n48159 = ~n48102 & ~n48158;
  assign n48160 = n3492 & ~n48159;
  assign n48161 = ~n21722 & ~n48160;
  assign n48162 = n3485 & ~n48161;
  assign n48163 = ~n21721 & ~n48162;
  assign n48164 = n3476 & ~n48163;
  assign n48165 = ~n48083 & ~n48164;
  assign n48166 = n3374 & ~n48165;
  assign n48167 = ~n48013 & ~n48166;
  assign n48168 = n3655 & ~n48167;
  assign n48169 = ~n22958 & ~n47986;
  assign n48170 = ~i_hbusreq2 & ~n48169;
  assign n48171 = ~n39776 & ~n48170;
  assign n48172 = ~controllable_hgrant2 & ~n48171;
  assign n48173 = ~n4562 & ~n48172;
  assign n48174 = controllable_hmaster1 & ~n48173;
  assign n48175 = controllable_hmaster0 & ~n48173;
  assign n48176 = controllable_hmaster0 & ~n48175;
  assign n48177 = ~controllable_hmaster1 & ~n48176;
  assign n48178 = ~n48174 & ~n48177;
  assign n48179 = ~i_hbusreq3 & ~n48178;
  assign n48180 = ~n40521 & ~n48179;
  assign n48181 = controllable_hmaster2 & ~n48180;
  assign n48182 = controllable_hmaster2 & ~n48181;
  assign n48183 = ~controllable_hgrant3 & ~n48182;
  assign n48184 = ~n9708 & ~n48183;
  assign n48185 = controllable_nhgrant0 & ~n48184;
  assign n48186 = ~n9753 & ~n48185;
  assign n48187 = ~n3281 & ~n48186;
  assign n48188 = ~n3281 & ~n48187;
  assign n48189 = ~n3378 & ~n48188;
  assign n48190 = ~n22618 & ~n48189;
  assign n48191 = n3492 & ~n48190;
  assign n48192 = n3492 & ~n48191;
  assign n48193 = n3485 & ~n48192;
  assign n48194 = n3485 & ~n48193;
  assign n48195 = ~n3374 & ~n48194;
  assign n48196 = ~n5303 & ~n38449;
  assign n48197 = ~controllable_hmaster1 & ~n48196;
  assign n48198 = ~n5293 & ~n48197;
  assign n48199 = i_hbusreq3 & ~n48198;
  assign n48200 = ~n22687 & ~n38449;
  assign n48201 = ~controllable_hmaster1 & ~n48200;
  assign n48202 = ~n22673 & ~n48201;
  assign n48203 = ~i_hbusreq3 & ~n48202;
  assign n48204 = ~n48199 & ~n48203;
  assign n48205 = ~controllable_hmaster2 & ~n48204;
  assign n48206 = ~n22668 & ~n48205;
  assign n48207 = ~controllable_hgrant3 & ~n48206;
  assign n48208 = ~n9790 & ~n48207;
  assign n48209 = controllable_nhgrant0 & ~n48208;
  assign n48210 = ~n9861 & ~n48209;
  assign n48211 = ~n3281 & ~n48210;
  assign n48212 = ~n3281 & ~n48211;
  assign n48213 = n3378 & ~n48212;
  assign n48214 = ~n23013 & ~n48032;
  assign n48215 = ~i_hbusreq2 & ~n48214;
  assign n48216 = ~n39843 & ~n48215;
  assign n48217 = ~controllable_hgrant2 & ~n48216;
  assign n48218 = ~n4562 & ~n48217;
  assign n48219 = ~controllable_hmaster0 & ~n48218;
  assign n48220 = ~n48175 & ~n48219;
  assign n48221 = ~controllable_hmaster1 & ~n48220;
  assign n48222 = ~n48174 & ~n48221;
  assign n48223 = ~i_hbusreq3 & ~n48222;
  assign n48224 = ~n40563 & ~n48223;
  assign n48225 = controllable_hmaster2 & ~n48224;
  assign n48226 = ~n35368 & ~n38449;
  assign n48227 = ~controllable_hmaster1 & ~n48226;
  assign n48228 = ~n35364 & ~n48227;
  assign n48229 = i_hbusreq3 & ~n48228;
  assign n48230 = ~n23013 & ~n47986;
  assign n48231 = ~i_hbusreq2 & ~n48230;
  assign n48232 = ~n35374 & ~n48231;
  assign n48233 = ~controllable_hgrant2 & ~n48232;
  assign n48234 = ~n4562 & ~n48233;
  assign n48235 = controllable_hmaster0 & ~n48234;
  assign n48236 = ~n9803 & ~n48233;
  assign n48237 = ~controllable_hmaster0 & ~n48236;
  assign n48238 = ~n48235 & ~n48237;
  assign n48239 = controllable_hmaster1 & ~n48238;
  assign n48240 = ~n23049 & ~n47986;
  assign n48241 = ~i_hbusreq2 & ~n48240;
  assign n48242 = ~n35385 & ~n48241;
  assign n48243 = ~controllable_hgrant2 & ~n48242;
  assign n48244 = ~n4562 & ~n48243;
  assign n48245 = controllable_hmaster0 & ~n48244;
  assign n48246 = ~n38449 & ~n48245;
  assign n48247 = ~controllable_hmaster1 & ~n48246;
  assign n48248 = ~n48239 & ~n48247;
  assign n48249 = ~i_hbusreq3 & ~n48248;
  assign n48250 = ~n48229 & ~n48249;
  assign n48251 = ~controllable_hmaster2 & ~n48250;
  assign n48252 = ~n48225 & ~n48251;
  assign n48253 = ~controllable_hgrant3 & ~n48252;
  assign n48254 = ~n9790 & ~n48253;
  assign n48255 = controllable_nhgrant0 & ~n48254;
  assign n48256 = ~n9861 & ~n48255;
  assign n48257 = ~n3281 & ~n48256;
  assign n48258 = ~n3281 & ~n48257;
  assign n48259 = ~n3378 & ~n48258;
  assign n48260 = ~n48213 & ~n48259;
  assign n48261 = n3492 & ~n48260;
  assign n48262 = n3492 & ~n48261;
  assign n48263 = n3485 & ~n48262;
  assign n48264 = n3485 & ~n48263;
  assign n48265 = ~n3476 & ~n48264;
  assign n48266 = ~controllable_hmaster0 & ~n40596;
  assign n48267 = ~n7339 & ~n48266;
  assign n48268 = ~controllable_hmaster1 & ~n48267;
  assign n48269 = ~n7330 & ~n48268;
  assign n48270 = i_hbusreq3 & ~n48269;
  assign n48271 = ~n22842 & ~n48266;
  assign n48272 = ~controllable_hmaster1 & ~n48271;
  assign n48273 = ~n22823 & ~n48272;
  assign n48274 = ~i_hbusreq3 & ~n48273;
  assign n48275 = ~n48270 & ~n48274;
  assign n48276 = ~controllable_hmaster2 & ~n48275;
  assign n48277 = ~n22808 & ~n48276;
  assign n48278 = ~controllable_hgrant3 & ~n48277;
  assign n48279 = ~n10110 & ~n48278;
  assign n48280 = controllable_nhgrant0 & ~n48279;
  assign n48281 = ~n10240 & ~n48280;
  assign n48282 = ~n3281 & ~n48281;
  assign n48283 = ~n3281 & ~n48282;
  assign n48284 = n3378 & ~n48283;
  assign n48285 = ~n23104 & ~n48103;
  assign n48286 = ~i_hbusreq2 & ~n48285;
  assign n48287 = ~n40636 & ~n48286;
  assign n48288 = ~controllable_hgrant2 & ~n48287;
  assign n48289 = ~n10111 & ~n48288;
  assign n48290 = controllable_hmaster1 & ~n48289;
  assign n48291 = controllable_hmaster0 & ~n48289;
  assign n48292 = ~n23119 & ~n48111;
  assign n48293 = ~i_hbusreq2 & ~n48292;
  assign n48294 = ~n40644 & ~n48293;
  assign n48295 = ~controllable_hgrant2 & ~n48294;
  assign n48296 = ~n10111 & ~n48295;
  assign n48297 = ~controllable_hmaster0 & ~n48296;
  assign n48298 = ~n48291 & ~n48297;
  assign n48299 = ~controllable_hmaster1 & ~n48298;
  assign n48300 = ~n48290 & ~n48299;
  assign n48301 = ~i_hbusreq3 & ~n48300;
  assign n48302 = ~n40635 & ~n48301;
  assign n48303 = controllable_hmaster2 & ~n48302;
  assign n48304 = ~n40664 & ~n43265;
  assign n48305 = controllable_hmaster1 & ~n48304;
  assign n48306 = ~controllable_hmaster0 & ~n40659;
  assign n48307 = ~n40670 & ~n48306;
  assign n48308 = ~controllable_hmaster1 & ~n48307;
  assign n48309 = ~n48305 & ~n48308;
  assign n48310 = i_hbusreq3 & ~n48309;
  assign n48311 = ~n23119 & ~n48103;
  assign n48312 = ~i_hbusreq2 & ~n48311;
  assign n48313 = ~n40684 & ~n48312;
  assign n48314 = ~controllable_hgrant2 & ~n48313;
  assign n48315 = ~n10111 & ~n48314;
  assign n48316 = controllable_hmaster0 & ~n48315;
  assign n48317 = ~n10152 & ~n48314;
  assign n48318 = ~controllable_hmaster0 & ~n48317;
  assign n48319 = ~n48316 & ~n48318;
  assign n48320 = controllable_hmaster1 & ~n48319;
  assign n48321 = ~n23157 & ~n48103;
  assign n48322 = ~i_hbusreq2 & ~n48321;
  assign n48323 = ~n40693 & ~n48322;
  assign n48324 = ~controllable_hgrant2 & ~n48323;
  assign n48325 = ~n10111 & ~n48324;
  assign n48326 = controllable_hmaster0 & ~n48325;
  assign n48327 = ~n48306 & ~n48326;
  assign n48328 = ~controllable_hmaster1 & ~n48327;
  assign n48329 = ~n48320 & ~n48328;
  assign n48330 = ~i_hbusreq3 & ~n48329;
  assign n48331 = ~n48310 & ~n48330;
  assign n48332 = ~controllable_hmaster2 & ~n48331;
  assign n48333 = ~n48303 & ~n48332;
  assign n48334 = ~controllable_hgrant3 & ~n48333;
  assign n48335 = ~n10110 & ~n48334;
  assign n48336 = controllable_nhgrant0 & ~n48335;
  assign n48337 = ~n10240 & ~n48336;
  assign n48338 = ~n3281 & ~n48337;
  assign n48339 = ~n3281 & ~n48338;
  assign n48340 = ~n3378 & ~n48339;
  assign n48341 = ~n48284 & ~n48340;
  assign n48342 = n3492 & ~n48341;
  assign n48343 = ~n21722 & ~n48342;
  assign n48344 = n3485 & ~n48343;
  assign n48345 = ~n21721 & ~n48344;
  assign n48346 = n3476 & ~n48345;
  assign n48347 = ~n48265 & ~n48346;
  assign n48348 = n3374 & ~n48347;
  assign n48349 = ~n48195 & ~n48348;
  assign n48350 = ~n3655 & ~n48349;
  assign n48351 = ~n48168 & ~n48350;
  assign n48352 = n3652 & ~n48351;
  assign n48353 = ~n23190 & ~n47990;
  assign n48354 = controllable_hmaster1 & ~n48353;
  assign n48355 = controllable_hmaster0 & ~n48353;
  assign n48356 = controllable_hmaster0 & ~n48355;
  assign n48357 = ~controllable_hmaster1 & ~n48356;
  assign n48358 = ~n48354 & ~n48357;
  assign n48359 = ~i_hbusreq3 & ~n48358;
  assign n48360 = ~n40735 & ~n48359;
  assign n48361 = controllable_hmaster2 & ~n48360;
  assign n48362 = controllable_hmaster2 & ~n48361;
  assign n48363 = ~controllable_hgrant3 & ~n48362;
  assign n48364 = ~n9708 & ~n48363;
  assign n48365 = controllable_nhgrant0 & ~n48364;
  assign n48366 = ~n9753 & ~n48365;
  assign n48367 = ~n3281 & ~n48366;
  assign n48368 = ~n3281 & ~n48367;
  assign n48369 = ~n3378 & ~n48368;
  assign n48370 = ~n22618 & ~n48369;
  assign n48371 = n3492 & ~n48370;
  assign n48372 = n3492 & ~n48371;
  assign n48373 = n3485 & ~n48372;
  assign n48374 = n3485 & ~n48373;
  assign n48375 = ~n3374 & ~n48374;
  assign n48376 = ~n5303 & ~n38728;
  assign n48377 = ~controllable_hmaster1 & ~n48376;
  assign n48378 = ~n5293 & ~n48377;
  assign n48379 = i_hbusreq3 & ~n48378;
  assign n48380 = ~n22687 & ~n38728;
  assign n48381 = ~controllable_hmaster1 & ~n48380;
  assign n48382 = ~n22673 & ~n48381;
  assign n48383 = ~i_hbusreq3 & ~n48382;
  assign n48384 = ~n48379 & ~n48383;
  assign n48385 = ~controllable_hmaster2 & ~n48384;
  assign n48386 = ~n22668 & ~n48385;
  assign n48387 = ~controllable_hgrant3 & ~n48386;
  assign n48388 = ~n9790 & ~n48387;
  assign n48389 = controllable_nhgrant0 & ~n48388;
  assign n48390 = ~n9861 & ~n48389;
  assign n48391 = ~n3281 & ~n48390;
  assign n48392 = ~n3281 & ~n48391;
  assign n48393 = n3378 & ~n48392;
  assign n48394 = ~n23190 & ~n48036;
  assign n48395 = ~controllable_hmaster0 & ~n48394;
  assign n48396 = ~n48355 & ~n48395;
  assign n48397 = ~controllable_hmaster1 & ~n48396;
  assign n48398 = ~n48354 & ~n48397;
  assign n48399 = ~i_hbusreq3 & ~n48398;
  assign n48400 = ~n40777 & ~n48399;
  assign n48401 = controllable_hmaster2 & ~n48400;
  assign n48402 = ~n35616 & ~n38728;
  assign n48403 = ~controllable_hmaster1 & ~n48402;
  assign n48404 = ~n35614 & ~n48403;
  assign n48405 = i_hbusreq3 & ~n48404;
  assign n48406 = ~n23190 & ~n48051;
  assign n48407 = controllable_hmaster0 & ~n48406;
  assign n48408 = ~n23245 & ~n48051;
  assign n48409 = ~controllable_hmaster0 & ~n48408;
  assign n48410 = ~n48407 & ~n48409;
  assign n48411 = controllable_hmaster1 & ~n48410;
  assign n48412 = ~n23190 & ~n48061;
  assign n48413 = controllable_hmaster0 & ~n48412;
  assign n48414 = ~n38728 & ~n48413;
  assign n48415 = ~controllable_hmaster1 & ~n48414;
  assign n48416 = ~n48411 & ~n48415;
  assign n48417 = ~i_hbusreq3 & ~n48416;
  assign n48418 = ~n48405 & ~n48417;
  assign n48419 = ~controllable_hmaster2 & ~n48418;
  assign n48420 = ~n48401 & ~n48419;
  assign n48421 = ~controllable_hgrant3 & ~n48420;
  assign n48422 = ~n9790 & ~n48421;
  assign n48423 = controllable_nhgrant0 & ~n48422;
  assign n48424 = ~n9861 & ~n48423;
  assign n48425 = ~n3281 & ~n48424;
  assign n48426 = ~n3281 & ~n48425;
  assign n48427 = ~n3378 & ~n48426;
  assign n48428 = ~n48393 & ~n48427;
  assign n48429 = n3492 & ~n48428;
  assign n48430 = n3492 & ~n48429;
  assign n48431 = n3485 & ~n48430;
  assign n48432 = n3485 & ~n48431;
  assign n48433 = ~n3476 & ~n48432;
  assign n48434 = ~controllable_hmaster0 & ~n40808;
  assign n48435 = ~n7339 & ~n48434;
  assign n48436 = ~controllable_hmaster1 & ~n48435;
  assign n48437 = ~n7330 & ~n48436;
  assign n48438 = i_hbusreq3 & ~n48437;
  assign n48439 = ~n22842 & ~n48434;
  assign n48440 = ~controllable_hmaster1 & ~n48439;
  assign n48441 = ~n22823 & ~n48440;
  assign n48442 = ~i_hbusreq3 & ~n48441;
  assign n48443 = ~n48438 & ~n48442;
  assign n48444 = ~controllable_hmaster2 & ~n48443;
  assign n48445 = ~n22808 & ~n48444;
  assign n48446 = ~controllable_hgrant3 & ~n48445;
  assign n48447 = ~n10110 & ~n48446;
  assign n48448 = controllable_nhgrant0 & ~n48447;
  assign n48449 = ~n10240 & ~n48448;
  assign n48450 = ~n3281 & ~n48449;
  assign n48451 = ~n3281 & ~n48450;
  assign n48452 = n3378 & ~n48451;
  assign n48453 = ~n23302 & ~n48107;
  assign n48454 = controllable_hmaster1 & ~n48453;
  assign n48455 = controllable_hmaster0 & ~n48453;
  assign n48456 = ~n23302 & ~n48115;
  assign n48457 = ~controllable_hmaster0 & ~n48456;
  assign n48458 = ~n48455 & ~n48457;
  assign n48459 = ~controllable_hmaster1 & ~n48458;
  assign n48460 = ~n48454 & ~n48459;
  assign n48461 = ~i_hbusreq3 & ~n48460;
  assign n48462 = ~n40838 & ~n48461;
  assign n48463 = controllable_hmaster2 & ~n48462;
  assign n48464 = ~controllable_hmaster0 & ~n40850;
  assign n48465 = ~n40857 & ~n48464;
  assign n48466 = ~controllable_hmaster1 & ~n48465;
  assign n48467 = ~n46019 & ~n48466;
  assign n48468 = i_hbusreq3 & ~n48467;
  assign n48469 = ~n23302 & ~n48132;
  assign n48470 = controllable_hmaster0 & ~n48469;
  assign n48471 = ~n23334 & ~n48132;
  assign n48472 = ~controllable_hmaster0 & ~n48471;
  assign n48473 = ~n48470 & ~n48472;
  assign n48474 = controllable_hmaster1 & ~n48473;
  assign n48475 = ~n23302 & ~n48142;
  assign n48476 = controllable_hmaster0 & ~n48475;
  assign n48477 = ~n48464 & ~n48476;
  assign n48478 = ~controllable_hmaster1 & ~n48477;
  assign n48479 = ~n48474 & ~n48478;
  assign n48480 = ~i_hbusreq3 & ~n48479;
  assign n48481 = ~n48468 & ~n48480;
  assign n48482 = ~controllable_hmaster2 & ~n48481;
  assign n48483 = ~n48463 & ~n48482;
  assign n48484 = ~controllable_hgrant3 & ~n48483;
  assign n48485 = ~n10110 & ~n48484;
  assign n48486 = controllable_nhgrant0 & ~n48485;
  assign n48487 = ~n10240 & ~n48486;
  assign n48488 = ~n3281 & ~n48487;
  assign n48489 = ~n3281 & ~n48488;
  assign n48490 = ~n3378 & ~n48489;
  assign n48491 = ~n48452 & ~n48490;
  assign n48492 = n3492 & ~n48491;
  assign n48493 = ~n21722 & ~n48492;
  assign n48494 = n3485 & ~n48493;
  assign n48495 = ~n21721 & ~n48494;
  assign n48496 = n3476 & ~n48495;
  assign n48497 = ~n48433 & ~n48496;
  assign n48498 = n3374 & ~n48497;
  assign n48499 = ~n48375 & ~n48498;
  assign n48500 = n3655 & ~n48499;
  assign n48501 = ~n23190 & ~n48172;
  assign n48502 = controllable_hmaster1 & ~n48501;
  assign n48503 = controllable_hmaster0 & ~n48501;
  assign n48504 = controllable_hmaster0 & ~n48503;
  assign n48505 = ~controllable_hmaster1 & ~n48504;
  assign n48506 = ~n48502 & ~n48505;
  assign n48507 = ~i_hbusreq3 & ~n48506;
  assign n48508 = ~n40901 & ~n48507;
  assign n48509 = controllable_hmaster2 & ~n48508;
  assign n48510 = controllable_hmaster2 & ~n48509;
  assign n48511 = ~controllable_hgrant3 & ~n48510;
  assign n48512 = ~n9708 & ~n48511;
  assign n48513 = controllable_nhgrant0 & ~n48512;
  assign n48514 = ~n9753 & ~n48513;
  assign n48515 = ~n3281 & ~n48514;
  assign n48516 = ~n3281 & ~n48515;
  assign n48517 = ~n3378 & ~n48516;
  assign n48518 = ~n22618 & ~n48517;
  assign n48519 = n3492 & ~n48518;
  assign n48520 = n3492 & ~n48519;
  assign n48521 = n3485 & ~n48520;
  assign n48522 = n3485 & ~n48521;
  assign n48523 = ~n3374 & ~n48522;
  assign n48524 = ~n5303 & ~n38937;
  assign n48525 = ~controllable_hmaster1 & ~n48524;
  assign n48526 = ~n5293 & ~n48525;
  assign n48527 = i_hbusreq3 & ~n48526;
  assign n48528 = ~n22687 & ~n38937;
  assign n48529 = ~controllable_hmaster1 & ~n48528;
  assign n48530 = ~n22673 & ~n48529;
  assign n48531 = ~i_hbusreq3 & ~n48530;
  assign n48532 = ~n48527 & ~n48531;
  assign n48533 = ~controllable_hmaster2 & ~n48532;
  assign n48534 = ~n22668 & ~n48533;
  assign n48535 = ~controllable_hgrant3 & ~n48534;
  assign n48536 = ~n9790 & ~n48535;
  assign n48537 = controllable_nhgrant0 & ~n48536;
  assign n48538 = ~n9861 & ~n48537;
  assign n48539 = ~n3281 & ~n48538;
  assign n48540 = ~n3281 & ~n48539;
  assign n48541 = n3378 & ~n48540;
  assign n48542 = ~n23190 & ~n48217;
  assign n48543 = ~controllable_hmaster0 & ~n48542;
  assign n48544 = ~n48503 & ~n48543;
  assign n48545 = ~controllable_hmaster1 & ~n48544;
  assign n48546 = ~n48502 & ~n48545;
  assign n48547 = ~i_hbusreq3 & ~n48546;
  assign n48548 = ~n40943 & ~n48547;
  assign n48549 = controllable_hmaster2 & ~n48548;
  assign n48550 = ~n35808 & ~n38937;
  assign n48551 = ~controllable_hmaster1 & ~n48550;
  assign n48552 = ~n35806 & ~n48551;
  assign n48553 = i_hbusreq3 & ~n48552;
  assign n48554 = ~n23190 & ~n48233;
  assign n48555 = controllable_hmaster0 & ~n48554;
  assign n48556 = ~n23245 & ~n48233;
  assign n48557 = ~controllable_hmaster0 & ~n48556;
  assign n48558 = ~n48555 & ~n48557;
  assign n48559 = controllable_hmaster1 & ~n48558;
  assign n48560 = ~n23190 & ~n48243;
  assign n48561 = controllable_hmaster0 & ~n48560;
  assign n48562 = ~n38937 & ~n48561;
  assign n48563 = ~controllable_hmaster1 & ~n48562;
  assign n48564 = ~n48559 & ~n48563;
  assign n48565 = ~i_hbusreq3 & ~n48564;
  assign n48566 = ~n48553 & ~n48565;
  assign n48567 = ~controllable_hmaster2 & ~n48566;
  assign n48568 = ~n48549 & ~n48567;
  assign n48569 = ~controllable_hgrant3 & ~n48568;
  assign n48570 = ~n9790 & ~n48569;
  assign n48571 = controllable_nhgrant0 & ~n48570;
  assign n48572 = ~n9861 & ~n48571;
  assign n48573 = ~n3281 & ~n48572;
  assign n48574 = ~n3281 & ~n48573;
  assign n48575 = ~n3378 & ~n48574;
  assign n48576 = ~n48541 & ~n48575;
  assign n48577 = n3492 & ~n48576;
  assign n48578 = n3492 & ~n48577;
  assign n48579 = n3485 & ~n48578;
  assign n48580 = n3485 & ~n48579;
  assign n48581 = ~n3476 & ~n48580;
  assign n48582 = ~controllable_hmaster0 & ~n40974;
  assign n48583 = ~n7339 & ~n48582;
  assign n48584 = ~controllable_hmaster1 & ~n48583;
  assign n48585 = ~n7330 & ~n48584;
  assign n48586 = i_hbusreq3 & ~n48585;
  assign n48587 = ~n22842 & ~n48582;
  assign n48588 = ~controllable_hmaster1 & ~n48587;
  assign n48589 = ~n22823 & ~n48588;
  assign n48590 = ~i_hbusreq3 & ~n48589;
  assign n48591 = ~n48586 & ~n48590;
  assign n48592 = ~controllable_hmaster2 & ~n48591;
  assign n48593 = ~n22808 & ~n48592;
  assign n48594 = ~controllable_hgrant3 & ~n48593;
  assign n48595 = ~n10110 & ~n48594;
  assign n48596 = controllable_nhgrant0 & ~n48595;
  assign n48597 = ~n10240 & ~n48596;
  assign n48598 = ~n3281 & ~n48597;
  assign n48599 = ~n3281 & ~n48598;
  assign n48600 = n3378 & ~n48599;
  assign n48601 = ~n23302 & ~n48288;
  assign n48602 = controllable_hmaster1 & ~n48601;
  assign n48603 = controllable_hmaster0 & ~n48601;
  assign n48604 = ~n23302 & ~n48295;
  assign n48605 = ~controllable_hmaster0 & ~n48604;
  assign n48606 = ~n48603 & ~n48605;
  assign n48607 = ~controllable_hmaster1 & ~n48606;
  assign n48608 = ~n48602 & ~n48607;
  assign n48609 = ~i_hbusreq3 & ~n48608;
  assign n48610 = ~n41004 & ~n48609;
  assign n48611 = controllable_hmaster2 & ~n48610;
  assign n48612 = controllable_hmaster0 & ~n41024;
  assign n48613 = ~n41019 & ~n48612;
  assign n48614 = controllable_hmaster1 & ~n48613;
  assign n48615 = ~controllable_hmaster0 & ~n41016;
  assign n48616 = ~n41023 & ~n48615;
  assign n48617 = ~controllable_hmaster1 & ~n48616;
  assign n48618 = ~n48614 & ~n48617;
  assign n48619 = i_hbusreq3 & ~n48618;
  assign n48620 = ~n23302 & ~n48314;
  assign n48621 = controllable_hmaster0 & ~n48620;
  assign n48622 = ~n23334 & ~n48314;
  assign n48623 = ~controllable_hmaster0 & ~n48622;
  assign n48624 = ~n48621 & ~n48623;
  assign n48625 = controllable_hmaster1 & ~n48624;
  assign n48626 = ~n23302 & ~n48324;
  assign n48627 = controllable_hmaster0 & ~n48626;
  assign n48628 = ~n48615 & ~n48627;
  assign n48629 = ~controllable_hmaster1 & ~n48628;
  assign n48630 = ~n48625 & ~n48629;
  assign n48631 = ~i_hbusreq3 & ~n48630;
  assign n48632 = ~n48619 & ~n48631;
  assign n48633 = ~controllable_hmaster2 & ~n48632;
  assign n48634 = ~n48611 & ~n48633;
  assign n48635 = ~controllable_hgrant3 & ~n48634;
  assign n48636 = ~n10110 & ~n48635;
  assign n48637 = controllable_nhgrant0 & ~n48636;
  assign n48638 = ~n10240 & ~n48637;
  assign n48639 = ~n3281 & ~n48638;
  assign n48640 = ~n3281 & ~n48639;
  assign n48641 = ~n3378 & ~n48640;
  assign n48642 = ~n48600 & ~n48641;
  assign n48643 = n3492 & ~n48642;
  assign n48644 = ~n21722 & ~n48643;
  assign n48645 = n3485 & ~n48644;
  assign n48646 = ~n21721 & ~n48645;
  assign n48647 = n3476 & ~n48646;
  assign n48648 = ~n48581 & ~n48647;
  assign n48649 = n3374 & ~n48648;
  assign n48650 = ~n48523 & ~n48649;
  assign n48651 = ~n3655 & ~n48650;
  assign n48652 = ~n48500 & ~n48651;
  assign n48653 = ~n3652 & ~n48652;
  assign n48654 = ~n48352 & ~n48653;
  assign n48655 = n3368 & ~n48654;
  assign n48656 = ~n47985 & ~n48655;
  assign n48657 = n3362 & ~n48656;
  assign n48658 = n3492 & ~n47382;
  assign n48659 = ~n3631 & ~n48658;
  assign n48660 = n3485 & ~n48659;
  assign n48661 = ~n3630 & ~n48660;
  assign n48662 = ~n3476 & ~n48661;
  assign n48663 = ~n23549 & ~n37006;
  assign n48664 = ~n3485 & ~n48663;
  assign n48665 = ~n8309 & ~n48658;
  assign n48666 = n3485 & ~n48665;
  assign n48667 = ~n48664 & ~n48666;
  assign n48668 = n3476 & ~n48667;
  assign n48669 = ~n48662 & ~n48668;
  assign n48670 = ~n3374 & ~n48669;
  assign n48671 = n3492 & ~n47436;
  assign n48672 = ~n3631 & ~n48671;
  assign n48673 = n3485 & ~n48672;
  assign n48674 = ~n3630 & ~n48673;
  assign n48675 = ~n3476 & ~n48674;
  assign n48676 = n3492 & ~n47522;
  assign n48677 = ~n8309 & ~n48676;
  assign n48678 = n3485 & ~n48677;
  assign n48679 = ~n48664 & ~n48678;
  assign n48680 = n3476 & ~n48679;
  assign n48681 = ~n48675 & ~n48680;
  assign n48682 = n3374 & ~n48681;
  assign n48683 = ~n48670 & ~n48682;
  assign n48684 = n3655 & ~n48683;
  assign n48685 = n3492 & ~n47546;
  assign n48686 = ~n3631 & ~n48685;
  assign n48687 = n3485 & ~n48686;
  assign n48688 = ~n3630 & ~n48687;
  assign n48689 = ~n3476 & ~n48688;
  assign n48690 = ~n23549 & ~n37048;
  assign n48691 = ~n3485 & ~n48690;
  assign n48692 = ~n8309 & ~n48685;
  assign n48693 = n3485 & ~n48692;
  assign n48694 = ~n48691 & ~n48693;
  assign n48695 = n3476 & ~n48694;
  assign n48696 = ~n48689 & ~n48695;
  assign n48697 = ~n3374 & ~n48696;
  assign n48698 = n3492 & ~n47600;
  assign n48699 = ~n3631 & ~n48698;
  assign n48700 = n3485 & ~n48699;
  assign n48701 = ~n3630 & ~n48700;
  assign n48702 = ~n3476 & ~n48701;
  assign n48703 = n3492 & ~n47684;
  assign n48704 = ~n8309 & ~n48703;
  assign n48705 = n3485 & ~n48704;
  assign n48706 = ~n48691 & ~n48705;
  assign n48707 = n3476 & ~n48706;
  assign n48708 = ~n48702 & ~n48707;
  assign n48709 = n3374 & ~n48708;
  assign n48710 = ~n48697 & ~n48709;
  assign n48711 = ~n3655 & ~n48710;
  assign n48712 = ~n48684 & ~n48711;
  assign n48713 = n3652 & ~n48712;
  assign n48714 = n3492 & ~n47710;
  assign n48715 = ~n3631 & ~n48714;
  assign n48716 = n3485 & ~n48715;
  assign n48717 = ~n3630 & ~n48716;
  assign n48718 = ~n3476 & ~n48717;
  assign n48719 = ~n23549 & ~n37091;
  assign n48720 = ~n3485 & ~n48719;
  assign n48721 = ~n8309 & ~n48714;
  assign n48722 = n3485 & ~n48721;
  assign n48723 = ~n48720 & ~n48722;
  assign n48724 = n3476 & ~n48723;
  assign n48725 = ~n48718 & ~n48724;
  assign n48726 = ~n3374 & ~n48725;
  assign n48727 = n3492 & ~n47764;
  assign n48728 = ~n3631 & ~n48727;
  assign n48729 = n3485 & ~n48728;
  assign n48730 = ~n3630 & ~n48729;
  assign n48731 = ~n3476 & ~n48730;
  assign n48732 = n3492 & ~n47828;
  assign n48733 = ~n8309 & ~n48732;
  assign n48734 = n3485 & ~n48733;
  assign n48735 = ~n48720 & ~n48734;
  assign n48736 = n3476 & ~n48735;
  assign n48737 = ~n48731 & ~n48736;
  assign n48738 = n3374 & ~n48737;
  assign n48739 = ~n48726 & ~n48738;
  assign n48740 = n3655 & ~n48739;
  assign n48741 = n3492 & ~n47852;
  assign n48742 = ~n3631 & ~n48741;
  assign n48743 = n3485 & ~n48742;
  assign n48744 = ~n3630 & ~n48743;
  assign n48745 = ~n3476 & ~n48744;
  assign n48746 = ~n23549 & ~n37132;
  assign n48747 = ~n3485 & ~n48746;
  assign n48748 = ~n8309 & ~n48741;
  assign n48749 = n3485 & ~n48748;
  assign n48750 = ~n48747 & ~n48749;
  assign n48751 = n3476 & ~n48750;
  assign n48752 = ~n48745 & ~n48751;
  assign n48753 = ~n3374 & ~n48752;
  assign n48754 = n3492 & ~n47906;
  assign n48755 = ~n3631 & ~n48754;
  assign n48756 = n3485 & ~n48755;
  assign n48757 = ~n3630 & ~n48756;
  assign n48758 = ~n3476 & ~n48757;
  assign n48759 = n3492 & ~n47970;
  assign n48760 = ~n8309 & ~n48759;
  assign n48761 = n3485 & ~n48760;
  assign n48762 = ~n48747 & ~n48761;
  assign n48763 = n3476 & ~n48762;
  assign n48764 = ~n48758 & ~n48763;
  assign n48765 = n3374 & ~n48764;
  assign n48766 = ~n48753 & ~n48765;
  assign n48767 = ~n3655 & ~n48766;
  assign n48768 = ~n48740 & ~n48767;
  assign n48769 = ~n3652 & ~n48768;
  assign n48770 = ~n48713 & ~n48769;
  assign n48771 = ~n3368 & ~n48770;
  assign n48772 = n3492 & ~n48006;
  assign n48773 = n3492 & ~n48772;
  assign n48774 = n3485 & ~n48773;
  assign n48775 = n3485 & ~n48774;
  assign n48776 = ~n3476 & ~n48775;
  assign n48777 = ~n8525 & ~n48774;
  assign n48778 = n3476 & ~n48777;
  assign n48779 = ~n48776 & ~n48778;
  assign n48780 = ~n3374 & ~n48779;
  assign n48781 = n3492 & ~n48076;
  assign n48782 = n3492 & ~n48781;
  assign n48783 = n3485 & ~n48782;
  assign n48784 = n3485 & ~n48783;
  assign n48785 = ~n3476 & ~n48784;
  assign n48786 = ~n23646 & ~n37174;
  assign n48787 = ~n3485 & ~n48786;
  assign n48788 = n3492 & ~n48157;
  assign n48789 = ~n21722 & ~n48788;
  assign n48790 = n3485 & ~n48789;
  assign n48791 = ~n48787 & ~n48790;
  assign n48792 = n3476 & ~n48791;
  assign n48793 = ~n48785 & ~n48792;
  assign n48794 = n3374 & ~n48793;
  assign n48795 = ~n48780 & ~n48794;
  assign n48796 = n3655 & ~n48795;
  assign n48797 = n3492 & ~n48188;
  assign n48798 = n3492 & ~n48797;
  assign n48799 = n3485 & ~n48798;
  assign n48800 = n3485 & ~n48799;
  assign n48801 = ~n3476 & ~n48800;
  assign n48802 = ~n8525 & ~n48799;
  assign n48803 = n3476 & ~n48802;
  assign n48804 = ~n48801 & ~n48803;
  assign n48805 = ~n3374 & ~n48804;
  assign n48806 = n3492 & ~n48258;
  assign n48807 = n3492 & ~n48806;
  assign n48808 = n3485 & ~n48807;
  assign n48809 = n3485 & ~n48808;
  assign n48810 = ~n3476 & ~n48809;
  assign n48811 = ~n23646 & ~n37202;
  assign n48812 = ~n3485 & ~n48811;
  assign n48813 = n3492 & ~n48339;
  assign n48814 = ~n21722 & ~n48813;
  assign n48815 = n3485 & ~n48814;
  assign n48816 = ~n48812 & ~n48815;
  assign n48817 = n3476 & ~n48816;
  assign n48818 = ~n48810 & ~n48817;
  assign n48819 = n3374 & ~n48818;
  assign n48820 = ~n48805 & ~n48819;
  assign n48821 = ~n3655 & ~n48820;
  assign n48822 = ~n48796 & ~n48821;
  assign n48823 = n3652 & ~n48822;
  assign n48824 = n3492 & ~n48368;
  assign n48825 = n3492 & ~n48824;
  assign n48826 = n3485 & ~n48825;
  assign n48827 = n3485 & ~n48826;
  assign n48828 = ~n3476 & ~n48827;
  assign n48829 = ~n8525 & ~n48826;
  assign n48830 = n3476 & ~n48829;
  assign n48831 = ~n48828 & ~n48830;
  assign n48832 = ~n3374 & ~n48831;
  assign n48833 = n3492 & ~n48426;
  assign n48834 = n3492 & ~n48833;
  assign n48835 = n3485 & ~n48834;
  assign n48836 = n3485 & ~n48835;
  assign n48837 = ~n3476 & ~n48836;
  assign n48838 = ~n23646 & ~n37231;
  assign n48839 = ~n3485 & ~n48838;
  assign n48840 = n3492 & ~n48489;
  assign n48841 = ~n21722 & ~n48840;
  assign n48842 = n3485 & ~n48841;
  assign n48843 = ~n48839 & ~n48842;
  assign n48844 = n3476 & ~n48843;
  assign n48845 = ~n48837 & ~n48844;
  assign n48846 = n3374 & ~n48845;
  assign n48847 = ~n48832 & ~n48846;
  assign n48848 = n3655 & ~n48847;
  assign n48849 = n3492 & ~n48516;
  assign n48850 = n3492 & ~n48849;
  assign n48851 = n3485 & ~n48850;
  assign n48852 = n3485 & ~n48851;
  assign n48853 = ~n3476 & ~n48852;
  assign n48854 = ~n8525 & ~n48851;
  assign n48855 = n3476 & ~n48854;
  assign n48856 = ~n48853 & ~n48855;
  assign n48857 = ~n3374 & ~n48856;
  assign n48858 = n3492 & ~n48574;
  assign n48859 = n3492 & ~n48858;
  assign n48860 = n3485 & ~n48859;
  assign n48861 = n3485 & ~n48860;
  assign n48862 = ~n3476 & ~n48861;
  assign n48863 = ~n23646 & ~n37258;
  assign n48864 = ~n3485 & ~n48863;
  assign n48865 = n3492 & ~n48640;
  assign n48866 = ~n21722 & ~n48865;
  assign n48867 = n3485 & ~n48866;
  assign n48868 = ~n48864 & ~n48867;
  assign n48869 = n3476 & ~n48868;
  assign n48870 = ~n48862 & ~n48869;
  assign n48871 = n3374 & ~n48870;
  assign n48872 = ~n48857 & ~n48871;
  assign n48873 = ~n3655 & ~n48872;
  assign n48874 = ~n48848 & ~n48873;
  assign n48875 = ~n3652 & ~n48874;
  assign n48876 = ~n48823 & ~n48875;
  assign n48877 = n3368 & ~n48876;
  assign n48878 = ~n48771 & ~n48877;
  assign n48879 = ~n3362 & ~n48878;
  assign n48880 = ~n48657 & ~n48879;
  assign n48881 = n3359 & ~n48880;
  assign n48882 = ~n37278 & ~n48666;
  assign n48883 = n3476 & ~n48882;
  assign n48884 = ~n48662 & ~n48883;
  assign n48885 = ~n3374 & ~n48884;
  assign n48886 = ~n37278 & ~n48678;
  assign n48887 = n3476 & ~n48886;
  assign n48888 = ~n48675 & ~n48887;
  assign n48889 = n3374 & ~n48888;
  assign n48890 = ~n48885 & ~n48889;
  assign n48891 = n3655 & ~n48890;
  assign n48892 = ~n37289 & ~n48693;
  assign n48893 = n3476 & ~n48892;
  assign n48894 = ~n48689 & ~n48893;
  assign n48895 = ~n3374 & ~n48894;
  assign n48896 = ~n37289 & ~n48705;
  assign n48897 = n3476 & ~n48896;
  assign n48898 = ~n48702 & ~n48897;
  assign n48899 = n3374 & ~n48898;
  assign n48900 = ~n48895 & ~n48899;
  assign n48901 = ~n3655 & ~n48900;
  assign n48902 = ~n48891 & ~n48901;
  assign n48903 = n3652 & ~n48902;
  assign n48904 = ~n37302 & ~n48722;
  assign n48905 = n3476 & ~n48904;
  assign n48906 = ~n48718 & ~n48905;
  assign n48907 = ~n3374 & ~n48906;
  assign n48908 = ~n37302 & ~n48734;
  assign n48909 = n3476 & ~n48908;
  assign n48910 = ~n48731 & ~n48909;
  assign n48911 = n3374 & ~n48910;
  assign n48912 = ~n48907 & ~n48911;
  assign n48913 = n3655 & ~n48912;
  assign n48914 = ~n37313 & ~n48749;
  assign n48915 = n3476 & ~n48914;
  assign n48916 = ~n48745 & ~n48915;
  assign n48917 = ~n3374 & ~n48916;
  assign n48918 = ~n37313 & ~n48761;
  assign n48919 = n3476 & ~n48918;
  assign n48920 = ~n48758 & ~n48919;
  assign n48921 = n3374 & ~n48920;
  assign n48922 = ~n48917 & ~n48921;
  assign n48923 = ~n3655 & ~n48922;
  assign n48924 = ~n48913 & ~n48923;
  assign n48925 = ~n3652 & ~n48924;
  assign n48926 = ~n48903 & ~n48925;
  assign n48927 = ~n3368 & ~n48926;
  assign n48928 = ~n8689 & ~n48774;
  assign n48929 = n3476 & ~n48928;
  assign n48930 = ~n48776 & ~n48929;
  assign n48931 = ~n3374 & ~n48930;
  assign n48932 = ~n37332 & ~n48790;
  assign n48933 = n3476 & ~n48932;
  assign n48934 = ~n48785 & ~n48933;
  assign n48935 = n3374 & ~n48934;
  assign n48936 = ~n48931 & ~n48935;
  assign n48937 = n3655 & ~n48936;
  assign n48938 = ~n8689 & ~n48799;
  assign n48939 = n3476 & ~n48938;
  assign n48940 = ~n48801 & ~n48939;
  assign n48941 = ~n3374 & ~n48940;
  assign n48942 = ~n37343 & ~n48815;
  assign n48943 = n3476 & ~n48942;
  assign n48944 = ~n48810 & ~n48943;
  assign n48945 = n3374 & ~n48944;
  assign n48946 = ~n48941 & ~n48945;
  assign n48947 = ~n3655 & ~n48946;
  assign n48948 = ~n48937 & ~n48947;
  assign n48949 = n3652 & ~n48948;
  assign n48950 = ~n8689 & ~n48826;
  assign n48951 = n3476 & ~n48950;
  assign n48952 = ~n48828 & ~n48951;
  assign n48953 = ~n3374 & ~n48952;
  assign n48954 = ~n37356 & ~n48842;
  assign n48955 = n3476 & ~n48954;
  assign n48956 = ~n48837 & ~n48955;
  assign n48957 = n3374 & ~n48956;
  assign n48958 = ~n48953 & ~n48957;
  assign n48959 = n3655 & ~n48958;
  assign n48960 = ~n8689 & ~n48851;
  assign n48961 = n3476 & ~n48960;
  assign n48962 = ~n48853 & ~n48961;
  assign n48963 = ~n3374 & ~n48962;
  assign n48964 = ~n37367 & ~n48867;
  assign n48965 = n3476 & ~n48964;
  assign n48966 = ~n48862 & ~n48965;
  assign n48967 = n3374 & ~n48966;
  assign n48968 = ~n48963 & ~n48967;
  assign n48969 = ~n3655 & ~n48968;
  assign n48970 = ~n48959 & ~n48969;
  assign n48971 = ~n3652 & ~n48970;
  assign n48972 = ~n48949 & ~n48971;
  assign n48973 = n3368 & ~n48972;
  assign n48974 = ~n48927 & ~n48973;
  assign n48975 = n3362 & ~n48974;
  assign n48976 = n3378 & ~n47382;
  assign n48977 = ~n37398 & ~n48976;
  assign n48978 = n3492 & ~n48977;
  assign n48979 = ~n3631 & ~n48978;
  assign n48980 = n3485 & ~n48979;
  assign n48981 = ~n3630 & ~n48980;
  assign n48982 = ~n3476 & ~n48981;
  assign n48983 = ~n37006 & ~n48978;
  assign n48984 = n3485 & ~n48983;
  assign n48985 = ~n37278 & ~n48984;
  assign n48986 = n3476 & ~n48985;
  assign n48987 = ~n48982 & ~n48986;
  assign n48988 = ~n3374 & ~n48987;
  assign n48989 = n3378 & ~n47436;
  assign n48990 = ~n37472 & ~n48989;
  assign n48991 = n3492 & ~n48990;
  assign n48992 = ~n3631 & ~n48991;
  assign n48993 = n3485 & ~n48992;
  assign n48994 = ~n3630 & ~n48993;
  assign n48995 = ~n3476 & ~n48994;
  assign n48996 = n3378 & ~n47522;
  assign n48997 = ~n37554 & ~n48996;
  assign n48998 = n3492 & ~n48997;
  assign n48999 = ~n37006 & ~n48998;
  assign n49000 = n3485 & ~n48999;
  assign n49001 = ~n37278 & ~n49000;
  assign n49002 = n3476 & ~n49001;
  assign n49003 = ~n48995 & ~n49002;
  assign n49004 = n3374 & ~n49003;
  assign n49005 = ~n48988 & ~n49004;
  assign n49006 = n3655 & ~n49005;
  assign n49007 = n3378 & ~n47546;
  assign n49008 = ~n37588 & ~n49007;
  assign n49009 = n3492 & ~n49008;
  assign n49010 = ~n3631 & ~n49009;
  assign n49011 = n3485 & ~n49010;
  assign n49012 = ~n3630 & ~n49011;
  assign n49013 = ~n3476 & ~n49012;
  assign n49014 = ~n37048 & ~n49009;
  assign n49015 = n3485 & ~n49014;
  assign n49016 = ~n37289 & ~n49015;
  assign n49017 = n3476 & ~n49016;
  assign n49018 = ~n49013 & ~n49017;
  assign n49019 = ~n3374 & ~n49018;
  assign n49020 = n3378 & ~n47600;
  assign n49021 = ~n37666 & ~n49020;
  assign n49022 = n3492 & ~n49021;
  assign n49023 = ~n3631 & ~n49022;
  assign n49024 = n3485 & ~n49023;
  assign n49025 = ~n3630 & ~n49024;
  assign n49026 = ~n3476 & ~n49025;
  assign n49027 = n3378 & ~n47684;
  assign n49028 = ~n37757 & ~n49027;
  assign n49029 = n3492 & ~n49028;
  assign n49030 = ~n37048 & ~n49029;
  assign n49031 = n3485 & ~n49030;
  assign n49032 = ~n37289 & ~n49031;
  assign n49033 = n3476 & ~n49032;
  assign n49034 = ~n49026 & ~n49033;
  assign n49035 = n3374 & ~n49034;
  assign n49036 = ~n49019 & ~n49035;
  assign n49037 = ~n3655 & ~n49036;
  assign n49038 = ~n49006 & ~n49037;
  assign n49039 = n3652 & ~n49038;
  assign n49040 = n3378 & ~n47710;
  assign n49041 = ~n37791 & ~n49040;
  assign n49042 = n3492 & ~n49041;
  assign n49043 = ~n3631 & ~n49042;
  assign n49044 = n3485 & ~n49043;
  assign n49045 = ~n3630 & ~n49044;
  assign n49046 = ~n3476 & ~n49045;
  assign n49047 = ~n37091 & ~n49042;
  assign n49048 = n3485 & ~n49047;
  assign n49049 = ~n37302 & ~n49048;
  assign n49050 = n3476 & ~n49049;
  assign n49051 = ~n49046 & ~n49050;
  assign n49052 = ~n3374 & ~n49051;
  assign n49053 = n3378 & ~n47764;
  assign n49054 = ~n37851 & ~n49053;
  assign n49055 = n3492 & ~n49054;
  assign n49056 = ~n3631 & ~n49055;
  assign n49057 = n3485 & ~n49056;
  assign n49058 = ~n3630 & ~n49057;
  assign n49059 = ~n3476 & ~n49058;
  assign n49060 = n3378 & ~n47828;
  assign n49061 = ~n37913 & ~n49060;
  assign n49062 = n3492 & ~n49061;
  assign n49063 = ~n37091 & ~n49062;
  assign n49064 = n3485 & ~n49063;
  assign n49065 = ~n37302 & ~n49064;
  assign n49066 = n3476 & ~n49065;
  assign n49067 = ~n49059 & ~n49066;
  assign n49068 = n3374 & ~n49067;
  assign n49069 = ~n49052 & ~n49068;
  assign n49070 = n3655 & ~n49069;
  assign n49071 = n3378 & ~n47852;
  assign n49072 = ~n37945 & ~n49071;
  assign n49073 = n3492 & ~n49072;
  assign n49074 = ~n3631 & ~n49073;
  assign n49075 = n3485 & ~n49074;
  assign n49076 = ~n3630 & ~n49075;
  assign n49077 = ~n3476 & ~n49076;
  assign n49078 = ~n37132 & ~n49073;
  assign n49079 = n3485 & ~n49078;
  assign n49080 = ~n37313 & ~n49079;
  assign n49081 = n3476 & ~n49080;
  assign n49082 = ~n49077 & ~n49081;
  assign n49083 = ~n3374 & ~n49082;
  assign n49084 = n3378 & ~n47906;
  assign n49085 = ~n38005 & ~n49084;
  assign n49086 = n3492 & ~n49085;
  assign n49087 = ~n3631 & ~n49086;
  assign n49088 = n3485 & ~n49087;
  assign n49089 = ~n3630 & ~n49088;
  assign n49090 = ~n3476 & ~n49089;
  assign n49091 = n3378 & ~n47970;
  assign n49092 = ~n38067 & ~n49091;
  assign n49093 = n3492 & ~n49092;
  assign n49094 = ~n37132 & ~n49093;
  assign n49095 = n3485 & ~n49094;
  assign n49096 = ~n37313 & ~n49095;
  assign n49097 = n3476 & ~n49096;
  assign n49098 = ~n49090 & ~n49097;
  assign n49099 = n3374 & ~n49098;
  assign n49100 = ~n49083 & ~n49099;
  assign n49101 = ~n3655 & ~n49100;
  assign n49102 = ~n49070 & ~n49101;
  assign n49103 = ~n3652 & ~n49102;
  assign n49104 = ~n49039 & ~n49103;
  assign n49105 = ~n3368 & ~n49104;
  assign n49106 = n3378 & ~n48006;
  assign n49107 = ~n38114 & ~n49106;
  assign n49108 = n3492 & ~n49107;
  assign n49109 = n3492 & ~n49108;
  assign n49110 = n3485 & ~n49109;
  assign n49111 = n3485 & ~n49110;
  assign n49112 = ~n3476 & ~n49111;
  assign n49113 = ~n8523 & ~n49108;
  assign n49114 = n3485 & ~n49113;
  assign n49115 = ~n8689 & ~n49114;
  assign n49116 = n3476 & ~n49115;
  assign n49117 = ~n49112 & ~n49116;
  assign n49118 = ~n3374 & ~n49117;
  assign n49119 = n3378 & ~n48076;
  assign n49120 = ~n38186 & ~n49119;
  assign n49121 = n3492 & ~n49120;
  assign n49122 = n3492 & ~n49121;
  assign n49123 = n3485 & ~n49122;
  assign n49124 = n3485 & ~n49123;
  assign n49125 = ~n3476 & ~n49124;
  assign n49126 = i_hlock4 & ~n24195;
  assign n49127 = ~i_hlock4 & ~n24205;
  assign n49128 = ~n49126 & ~n49127;
  assign n49129 = ~i_hbusreq4 & ~n49128;
  assign n49130 = ~n41552 & ~n49129;
  assign n49131 = controllable_hgrant4 & ~n49130;
  assign n49132 = ~n23984 & ~n49131;
  assign n49133 = ~i_hbusreq2 & ~n49132;
  assign n49134 = ~n41551 & ~n49133;
  assign n49135 = ~controllable_hgrant2 & ~n49134;
  assign n49136 = ~n10111 & ~n49135;
  assign n49137 = controllable_hmaster1 & ~n49136;
  assign n49138 = controllable_hmaster0 & ~n49136;
  assign n49139 = i_hlock4 & ~n24236;
  assign n49140 = ~i_hlock4 & ~n24246;
  assign n49141 = ~n49139 & ~n49140;
  assign n49142 = ~i_hbusreq4 & ~n49141;
  assign n49143 = ~n41567 & ~n49142;
  assign n49144 = controllable_hgrant4 & ~n49143;
  assign n49145 = ~n23999 & ~n49144;
  assign n49146 = ~i_hbusreq2 & ~n49145;
  assign n49147 = ~n41566 & ~n49146;
  assign n49148 = ~controllable_hgrant2 & ~n49147;
  assign n49149 = ~n10111 & ~n49148;
  assign n49150 = ~controllable_hmaster0 & ~n49149;
  assign n49151 = ~n49138 & ~n49150;
  assign n49152 = ~controllable_hmaster1 & ~n49151;
  assign n49153 = ~n49137 & ~n49152;
  assign n49154 = ~i_hbusreq3 & ~n49153;
  assign n49155 = ~n41550 & ~n49154;
  assign n49156 = controllable_hmaster2 & ~n49155;
  assign n49157 = ~n38325 & ~n41595;
  assign n49158 = ~controllable_hmaster1 & ~n49157;
  assign n49159 = ~n46641 & ~n49158;
  assign n49160 = i_hbusreq3 & ~n49159;
  assign n49161 = ~n23999 & ~n49131;
  assign n49162 = ~i_hbusreq2 & ~n49161;
  assign n49163 = ~n41614 & ~n49162;
  assign n49164 = ~controllable_hgrant2 & ~n49163;
  assign n49165 = ~n10111 & ~n49164;
  assign n49166 = controllable_hmaster0 & ~n49165;
  assign n49167 = ~n10152 & ~n49164;
  assign n49168 = ~controllable_hmaster0 & ~n49167;
  assign n49169 = ~n49166 & ~n49168;
  assign n49170 = controllable_hmaster1 & ~n49169;
  assign n49171 = ~n24029 & ~n49131;
  assign n49172 = ~i_hbusreq2 & ~n49171;
  assign n49173 = ~n41623 & ~n49172;
  assign n49174 = ~controllable_hgrant2 & ~n49173;
  assign n49175 = ~n10111 & ~n49174;
  assign n49176 = controllable_hmaster0 & ~n49175;
  assign n49177 = ~n38357 & ~n49176;
  assign n49178 = ~controllable_hmaster1 & ~n49177;
  assign n49179 = ~n49170 & ~n49178;
  assign n49180 = ~i_hbusreq3 & ~n49179;
  assign n49181 = ~n49160 & ~n49180;
  assign n49182 = ~controllable_hmaster2 & ~n49181;
  assign n49183 = ~n49156 & ~n49182;
  assign n49184 = ~controllable_hgrant3 & ~n49183;
  assign n49185 = ~n10110 & ~n49184;
  assign n49186 = controllable_nhgrant0 & ~n49185;
  assign n49187 = ~n10240 & ~n49186;
  assign n49188 = ~n3281 & ~n49187;
  assign n49189 = ~n3281 & ~n49188;
  assign n49190 = n3378 & ~n49189;
  assign n49191 = ~n38371 & ~n49190;
  assign n49192 = n3492 & ~n49191;
  assign n49193 = ~n37174 & ~n49192;
  assign n49194 = n3485 & ~n49193;
  assign n49195 = ~n37332 & ~n49194;
  assign n49196 = n3476 & ~n49195;
  assign n49197 = ~n49125 & ~n49196;
  assign n49198 = n3374 & ~n49197;
  assign n49199 = ~n49118 & ~n49198;
  assign n49200 = n3655 & ~n49199;
  assign n49201 = n3378 & ~n48188;
  assign n49202 = ~n38413 & ~n49201;
  assign n49203 = n3492 & ~n49202;
  assign n49204 = n3492 & ~n49203;
  assign n49205 = n3485 & ~n49204;
  assign n49206 = n3485 & ~n49205;
  assign n49207 = ~n3476 & ~n49206;
  assign n49208 = ~n8523 & ~n49203;
  assign n49209 = n3485 & ~n49208;
  assign n49210 = ~n8689 & ~n49209;
  assign n49211 = n3476 & ~n49210;
  assign n49212 = ~n49207 & ~n49211;
  assign n49213 = ~n3374 & ~n49212;
  assign n49214 = n3378 & ~n48258;
  assign n49215 = ~n38485 & ~n49214;
  assign n49216 = n3492 & ~n49215;
  assign n49217 = n3492 & ~n49216;
  assign n49218 = n3485 & ~n49217;
  assign n49219 = n3485 & ~n49218;
  assign n49220 = ~n3476 & ~n49219;
  assign n49221 = ~n24088 & ~n49131;
  assign n49222 = ~i_hbusreq2 & ~n49221;
  assign n49223 = ~n41699 & ~n49222;
  assign n49224 = ~controllable_hgrant2 & ~n49223;
  assign n49225 = ~n10111 & ~n49224;
  assign n49226 = controllable_hmaster1 & ~n49225;
  assign n49227 = controllable_hmaster0 & ~n49225;
  assign n49228 = ~n24104 & ~n49144;
  assign n49229 = ~i_hbusreq2 & ~n49228;
  assign n49230 = ~n41707 & ~n49229;
  assign n49231 = ~controllable_hgrant2 & ~n49230;
  assign n49232 = ~n10111 & ~n49231;
  assign n49233 = ~controllable_hmaster0 & ~n49232;
  assign n49234 = ~n49227 & ~n49233;
  assign n49235 = ~controllable_hmaster1 & ~n49234;
  assign n49236 = ~n49226 & ~n49235;
  assign n49237 = ~i_hbusreq3 & ~n49236;
  assign n49238 = ~n41698 & ~n49237;
  assign n49239 = controllable_hmaster2 & ~n49238;
  assign n49240 = ~n41723 & ~n44127;
  assign n49241 = controllable_hmaster1 & ~n49240;
  assign n49242 = ~n38618 & ~n41729;
  assign n49243 = ~controllable_hmaster1 & ~n49242;
  assign n49244 = ~n49241 & ~n49243;
  assign n49245 = i_hbusreq3 & ~n49244;
  assign n49246 = ~n24104 & ~n49131;
  assign n49247 = ~i_hbusreq2 & ~n49246;
  assign n49248 = ~n41742 & ~n49247;
  assign n49249 = ~controllable_hgrant2 & ~n49248;
  assign n49250 = ~n10111 & ~n49249;
  assign n49251 = controllable_hmaster0 & ~n49250;
  assign n49252 = ~n10152 & ~n49249;
  assign n49253 = ~controllable_hmaster0 & ~n49252;
  assign n49254 = ~n49251 & ~n49253;
  assign n49255 = controllable_hmaster1 & ~n49254;
  assign n49256 = ~n24138 & ~n49131;
  assign n49257 = ~i_hbusreq2 & ~n49256;
  assign n49258 = ~n41751 & ~n49257;
  assign n49259 = ~controllable_hgrant2 & ~n49258;
  assign n49260 = ~n10111 & ~n49259;
  assign n49261 = controllable_hmaster0 & ~n49260;
  assign n49262 = ~n38645 & ~n49261;
  assign n49263 = ~controllable_hmaster1 & ~n49262;
  assign n49264 = ~n49255 & ~n49263;
  assign n49265 = ~i_hbusreq3 & ~n49264;
  assign n49266 = ~n49245 & ~n49265;
  assign n49267 = ~controllable_hmaster2 & ~n49266;
  assign n49268 = ~n49239 & ~n49267;
  assign n49269 = ~controllable_hgrant3 & ~n49268;
  assign n49270 = ~n10110 & ~n49269;
  assign n49271 = controllable_nhgrant0 & ~n49270;
  assign n49272 = ~n10240 & ~n49271;
  assign n49273 = ~n3281 & ~n49272;
  assign n49274 = ~n3281 & ~n49273;
  assign n49275 = n3378 & ~n49274;
  assign n49276 = ~n38659 & ~n49275;
  assign n49277 = n3492 & ~n49276;
  assign n49278 = ~n37202 & ~n49277;
  assign n49279 = n3485 & ~n49278;
  assign n49280 = ~n37343 & ~n49279;
  assign n49281 = n3476 & ~n49280;
  assign n49282 = ~n49220 & ~n49281;
  assign n49283 = n3374 & ~n49282;
  assign n49284 = ~n49213 & ~n49283;
  assign n49285 = ~n3655 & ~n49284;
  assign n49286 = ~n49200 & ~n49285;
  assign n49287 = n3652 & ~n49286;
  assign n49288 = n3378 & ~n48368;
  assign n49289 = ~n38696 & ~n49288;
  assign n49290 = n3492 & ~n49289;
  assign n49291 = n3492 & ~n49290;
  assign n49292 = n3485 & ~n49291;
  assign n49293 = n3485 & ~n49292;
  assign n49294 = ~n3476 & ~n49293;
  assign n49295 = ~n8523 & ~n49290;
  assign n49296 = n3485 & ~n49295;
  assign n49297 = ~n8689 & ~n49296;
  assign n49298 = n3476 & ~n49297;
  assign n49299 = ~n49294 & ~n49298;
  assign n49300 = ~n3374 & ~n49299;
  assign n49301 = n3378 & ~n48426;
  assign n49302 = ~n38754 & ~n49301;
  assign n49303 = n3492 & ~n49302;
  assign n49304 = n3492 & ~n49303;
  assign n49305 = n3485 & ~n49304;
  assign n49306 = n3485 & ~n49305;
  assign n49307 = ~n3476 & ~n49306;
  assign n49308 = ~n24214 & ~n49135;
  assign n49309 = controllable_hmaster1 & ~n49308;
  assign n49310 = controllable_hmaster0 & ~n49308;
  assign n49311 = ~n24214 & ~n49148;
  assign n49312 = ~controllable_hmaster0 & ~n49311;
  assign n49313 = ~n49310 & ~n49312;
  assign n49314 = ~controllable_hmaster1 & ~n49313;
  assign n49315 = ~n49309 & ~n49314;
  assign n49316 = ~i_hbusreq3 & ~n49315;
  assign n49317 = ~n41818 & ~n49316;
  assign n49318 = controllable_hmaster2 & ~n49317;
  assign n49319 = ~n38842 & ~n41835;
  assign n49320 = ~controllable_hmaster1 & ~n49319;
  assign n49321 = ~n46828 & ~n49320;
  assign n49322 = i_hbusreq3 & ~n49321;
  assign n49323 = ~n24214 & ~n49164;
  assign n49324 = controllable_hmaster0 & ~n49323;
  assign n49325 = ~n24255 & ~n49164;
  assign n49326 = ~controllable_hmaster0 & ~n49325;
  assign n49327 = ~n49324 & ~n49326;
  assign n49328 = controllable_hmaster1 & ~n49327;
  assign n49329 = ~n24214 & ~n49174;
  assign n49330 = controllable_hmaster0 & ~n49329;
  assign n49331 = ~n38856 & ~n49330;
  assign n49332 = ~controllable_hmaster1 & ~n49331;
  assign n49333 = ~n49328 & ~n49332;
  assign n49334 = ~i_hbusreq3 & ~n49333;
  assign n49335 = ~n49322 & ~n49334;
  assign n49336 = ~controllable_hmaster2 & ~n49335;
  assign n49337 = ~n49318 & ~n49336;
  assign n49338 = ~controllable_hgrant3 & ~n49337;
  assign n49339 = ~n10110 & ~n49338;
  assign n49340 = controllable_nhgrant0 & ~n49339;
  assign n49341 = ~n10240 & ~n49340;
  assign n49342 = ~n3281 & ~n49341;
  assign n49343 = ~n3281 & ~n49342;
  assign n49344 = n3378 & ~n49343;
  assign n49345 = ~n38870 & ~n49344;
  assign n49346 = n3492 & ~n49345;
  assign n49347 = ~n37231 & ~n49346;
  assign n49348 = n3485 & ~n49347;
  assign n49349 = ~n37356 & ~n49348;
  assign n49350 = n3476 & ~n49349;
  assign n49351 = ~n49307 & ~n49350;
  assign n49352 = n3374 & ~n49351;
  assign n49353 = ~n49300 & ~n49352;
  assign n49354 = n3655 & ~n49353;
  assign n49355 = n3378 & ~n48516;
  assign n49356 = ~n38905 & ~n49355;
  assign n49357 = n3492 & ~n49356;
  assign n49358 = n3492 & ~n49357;
  assign n49359 = n3485 & ~n49358;
  assign n49360 = n3485 & ~n49359;
  assign n49361 = ~n3476 & ~n49360;
  assign n49362 = ~n8523 & ~n49357;
  assign n49363 = n3485 & ~n49362;
  assign n49364 = ~n8689 & ~n49363;
  assign n49365 = n3476 & ~n49364;
  assign n49366 = ~n49361 & ~n49365;
  assign n49367 = ~n3374 & ~n49366;
  assign n49368 = n3378 & ~n48574;
  assign n49369 = ~n38963 & ~n49368;
  assign n49370 = n3492 & ~n49369;
  assign n49371 = n3492 & ~n49370;
  assign n49372 = n3485 & ~n49371;
  assign n49373 = n3485 & ~n49372;
  assign n49374 = ~n3476 & ~n49373;
  assign n49375 = ~n24214 & ~n49224;
  assign n49376 = controllable_hmaster1 & ~n49375;
  assign n49377 = controllable_hmaster0 & ~n49375;
  assign n49378 = ~n24214 & ~n49231;
  assign n49379 = ~controllable_hmaster0 & ~n49378;
  assign n49380 = ~n49377 & ~n49379;
  assign n49381 = ~controllable_hmaster1 & ~n49380;
  assign n49382 = ~n49376 & ~n49381;
  assign n49383 = ~i_hbusreq3 & ~n49382;
  assign n49384 = ~n41904 & ~n49383;
  assign n49385 = controllable_hmaster2 & ~n49384;
  assign n49386 = controllable_hmaster0 & ~n41922;
  assign n49387 = ~n41917 & ~n49386;
  assign n49388 = controllable_hmaster1 & ~n49387;
  assign n49389 = ~n39051 & ~n41921;
  assign n49390 = ~controllable_hmaster1 & ~n49389;
  assign n49391 = ~n49388 & ~n49390;
  assign n49392 = i_hbusreq3 & ~n49391;
  assign n49393 = ~n24214 & ~n49249;
  assign n49394 = controllable_hmaster0 & ~n49393;
  assign n49395 = ~n24255 & ~n49249;
  assign n49396 = ~controllable_hmaster0 & ~n49395;
  assign n49397 = ~n49394 & ~n49396;
  assign n49398 = controllable_hmaster1 & ~n49397;
  assign n49399 = ~n24214 & ~n49259;
  assign n49400 = controllable_hmaster0 & ~n49399;
  assign n49401 = ~n39065 & ~n49400;
  assign n49402 = ~controllable_hmaster1 & ~n49401;
  assign n49403 = ~n49398 & ~n49402;
  assign n49404 = ~i_hbusreq3 & ~n49403;
  assign n49405 = ~n49392 & ~n49404;
  assign n49406 = ~controllable_hmaster2 & ~n49405;
  assign n49407 = ~n49385 & ~n49406;
  assign n49408 = ~controllable_hgrant3 & ~n49407;
  assign n49409 = ~n10110 & ~n49408;
  assign n49410 = controllable_nhgrant0 & ~n49409;
  assign n49411 = ~n10240 & ~n49410;
  assign n49412 = ~n3281 & ~n49411;
  assign n49413 = ~n3281 & ~n49412;
  assign n49414 = n3378 & ~n49413;
  assign n49415 = ~n39079 & ~n49414;
  assign n49416 = n3492 & ~n49415;
  assign n49417 = ~n37258 & ~n49416;
  assign n49418 = n3485 & ~n49417;
  assign n49419 = ~n37367 & ~n49418;
  assign n49420 = n3476 & ~n49419;
  assign n49421 = ~n49374 & ~n49420;
  assign n49422 = n3374 & ~n49421;
  assign n49423 = ~n49367 & ~n49422;
  assign n49424 = ~n3655 & ~n49423;
  assign n49425 = ~n49354 & ~n49424;
  assign n49426 = ~n3652 & ~n49425;
  assign n49427 = ~n49287 & ~n49426;
  assign n49428 = n3368 & ~n49427;
  assign n49429 = ~n49105 & ~n49428;
  assign n49430 = ~n3362 & ~n49429;
  assign n49431 = ~n48975 & ~n49430;
  assign n49432 = ~n3359 & ~n49431;
  assign n49433 = ~n48881 & ~n49432;
  assign n49434 = ~n3356 & ~n49433;
  assign n49435 = ~n47369 & ~n49434;
  assign n49436 = n3345 & ~n49435;
  assign n49437 = ~n46963 & ~n49436;
  assign n49438 = ~n3341 & ~n49437;
  assign n49439 = controllable_hmaster0 & ~n34156;
  assign n49440 = ~controllable_hmaster1 & ~n49439;
  assign n49441 = ~n34155 & ~n49440;
  assign n49442 = controllable_hmaster2 & ~n49441;
  assign n49443 = controllable_hmaster2 & ~n49442;
  assign n49444 = ~controllable_hgrant3 & ~n49443;
  assign n49445 = ~n24368 & ~n49444;
  assign n49446 = controllable_nhgrant0 & ~n49445;
  assign n49447 = ~n24376 & ~n49446;
  assign n49448 = ~n3281 & ~n49447;
  assign n49449 = ~n3783 & ~n49448;
  assign n49450 = ~n3378 & ~n49449;
  assign n49451 = ~n3378 & ~n49450;
  assign n49452 = n3492 & ~n49451;
  assign n49453 = ~n3493 & ~n49452;
  assign n49454 = n3485 & ~n49453;
  assign n49455 = ~n3486 & ~n49454;
  assign n49456 = ~n3476 & ~n49455;
  assign n49457 = ~n3281 & ~n37396;
  assign n49458 = n3378 & ~n49457;
  assign n49459 = ~n37398 & ~n49458;
  assign n49460 = n3492 & ~n49459;
  assign n49461 = ~n3493 & ~n49460;
  assign n49462 = n3485 & ~n49461;
  assign n49463 = ~n3486 & ~n49462;
  assign n49464 = n3476 & ~n49463;
  assign n49465 = ~n49456 & ~n49464;
  assign n49466 = ~n3374 & ~n49465;
  assign n49467 = ~n3950 & ~n49448;
  assign n49468 = ~n3378 & ~n49467;
  assign n49469 = ~n3378 & ~n49468;
  assign n49470 = n3492 & ~n49469;
  assign n49471 = ~n3493 & ~n49470;
  assign n49472 = n3485 & ~n49471;
  assign n49473 = ~n3486 & ~n49472;
  assign n49474 = ~n3476 & ~n49473;
  assign n49475 = ~n3281 & ~n37552;
  assign n49476 = n3378 & ~n49475;
  assign n49477 = ~n37554 & ~n49476;
  assign n49478 = n3492 & ~n49477;
  assign n49479 = ~n3493 & ~n49478;
  assign n49480 = n3485 & ~n49479;
  assign n49481 = ~n3486 & ~n49480;
  assign n49482 = n3476 & ~n49481;
  assign n49483 = ~n49474 & ~n49482;
  assign n49484 = n3374 & ~n49483;
  assign n49485 = ~n49466 & ~n49484;
  assign n49486 = n3655 & ~n49485;
  assign n49487 = controllable_hmaster0 & ~n37570;
  assign n49488 = ~controllable_hmaster1 & ~n49487;
  assign n49489 = ~n37569 & ~n49488;
  assign n49490 = controllable_hmaster2 & ~n49489;
  assign n49491 = controllable_hmaster2 & ~n49490;
  assign n49492 = ~controllable_hgrant3 & ~n49491;
  assign n49493 = ~n24368 & ~n49492;
  assign n49494 = controllable_nhgrant0 & ~n49493;
  assign n49495 = ~n24376 & ~n49494;
  assign n49496 = ~n3281 & ~n49495;
  assign n49497 = ~n3783 & ~n49496;
  assign n49498 = ~n3378 & ~n49497;
  assign n49499 = ~n3378 & ~n49498;
  assign n49500 = n3492 & ~n49499;
  assign n49501 = ~n3493 & ~n49500;
  assign n49502 = n3485 & ~n49501;
  assign n49503 = ~n3486 & ~n49502;
  assign n49504 = ~n3476 & ~n49503;
  assign n49505 = ~n3281 & ~n37586;
  assign n49506 = n3378 & ~n49505;
  assign n49507 = ~n37588 & ~n49506;
  assign n49508 = n3492 & ~n49507;
  assign n49509 = ~n3493 & ~n49508;
  assign n49510 = n3485 & ~n49509;
  assign n49511 = ~n3486 & ~n49510;
  assign n49512 = n3476 & ~n49511;
  assign n49513 = ~n49504 & ~n49512;
  assign n49514 = ~n3374 & ~n49513;
  assign n49515 = ~n3950 & ~n49496;
  assign n49516 = ~n3378 & ~n49515;
  assign n49517 = ~n3378 & ~n49516;
  assign n49518 = n3492 & ~n49517;
  assign n49519 = ~n3493 & ~n49518;
  assign n49520 = n3485 & ~n49519;
  assign n49521 = ~n3486 & ~n49520;
  assign n49522 = ~n3476 & ~n49521;
  assign n49523 = ~n3281 & ~n37755;
  assign n49524 = n3378 & ~n49523;
  assign n49525 = ~n37757 & ~n49524;
  assign n49526 = n3492 & ~n49525;
  assign n49527 = ~n3493 & ~n49526;
  assign n49528 = n3485 & ~n49527;
  assign n49529 = ~n3486 & ~n49528;
  assign n49530 = n3476 & ~n49529;
  assign n49531 = ~n49522 & ~n49530;
  assign n49532 = n3374 & ~n49531;
  assign n49533 = ~n49514 & ~n49532;
  assign n49534 = ~n3655 & ~n49533;
  assign n49535 = ~n49486 & ~n49534;
  assign n49536 = n3652 & ~n49535;
  assign n49537 = controllable_hmaster0 & ~n37773;
  assign n49538 = ~controllable_hmaster1 & ~n49537;
  assign n49539 = ~n37772 & ~n49538;
  assign n49540 = controllable_hmaster2 & ~n49539;
  assign n49541 = controllable_hmaster2 & ~n49540;
  assign n49542 = ~controllable_hgrant3 & ~n49541;
  assign n49543 = ~n24368 & ~n49542;
  assign n49544 = controllable_nhgrant0 & ~n49543;
  assign n49545 = ~n24376 & ~n49544;
  assign n49546 = ~n3281 & ~n49545;
  assign n49547 = ~n3783 & ~n49546;
  assign n49548 = ~n3378 & ~n49547;
  assign n49549 = ~n3378 & ~n49548;
  assign n49550 = n3492 & ~n49549;
  assign n49551 = ~n3493 & ~n49550;
  assign n49552 = n3485 & ~n49551;
  assign n49553 = ~n3486 & ~n49552;
  assign n49554 = ~n3476 & ~n49553;
  assign n49555 = ~n3281 & ~n37789;
  assign n49556 = n3378 & ~n49555;
  assign n49557 = ~n37791 & ~n49556;
  assign n49558 = n3492 & ~n49557;
  assign n49559 = ~n3493 & ~n49558;
  assign n49560 = n3485 & ~n49559;
  assign n49561 = ~n3486 & ~n49560;
  assign n49562 = n3476 & ~n49561;
  assign n49563 = ~n49554 & ~n49562;
  assign n49564 = ~n3374 & ~n49563;
  assign n49565 = ~n3950 & ~n49546;
  assign n49566 = ~n3378 & ~n49565;
  assign n49567 = ~n3378 & ~n49566;
  assign n49568 = n3492 & ~n49567;
  assign n49569 = ~n3493 & ~n49568;
  assign n49570 = n3485 & ~n49569;
  assign n49571 = ~n3486 & ~n49570;
  assign n49572 = ~n3476 & ~n49571;
  assign n49573 = ~n3281 & ~n37911;
  assign n49574 = n3378 & ~n49573;
  assign n49575 = ~n37913 & ~n49574;
  assign n49576 = n3492 & ~n49575;
  assign n49577 = ~n3493 & ~n49576;
  assign n49578 = n3485 & ~n49577;
  assign n49579 = ~n3486 & ~n49578;
  assign n49580 = n3476 & ~n49579;
  assign n49581 = ~n49572 & ~n49580;
  assign n49582 = n3374 & ~n49581;
  assign n49583 = ~n49564 & ~n49582;
  assign n49584 = n3655 & ~n49583;
  assign n49585 = controllable_hmaster0 & ~n37927;
  assign n49586 = ~controllable_hmaster1 & ~n49585;
  assign n49587 = ~n37926 & ~n49586;
  assign n49588 = controllable_hmaster2 & ~n49587;
  assign n49589 = controllable_hmaster2 & ~n49588;
  assign n49590 = ~controllable_hgrant3 & ~n49589;
  assign n49591 = ~n24368 & ~n49590;
  assign n49592 = controllable_nhgrant0 & ~n49591;
  assign n49593 = ~n24376 & ~n49592;
  assign n49594 = ~n3281 & ~n49593;
  assign n49595 = ~n3783 & ~n49594;
  assign n49596 = ~n3378 & ~n49595;
  assign n49597 = ~n3378 & ~n49596;
  assign n49598 = n3492 & ~n49597;
  assign n49599 = ~n3493 & ~n49598;
  assign n49600 = n3485 & ~n49599;
  assign n49601 = ~n3486 & ~n49600;
  assign n49602 = ~n3476 & ~n49601;
  assign n49603 = ~n3281 & ~n37943;
  assign n49604 = n3378 & ~n49603;
  assign n49605 = ~n37945 & ~n49604;
  assign n49606 = n3492 & ~n49605;
  assign n49607 = ~n3493 & ~n49606;
  assign n49608 = n3485 & ~n49607;
  assign n49609 = ~n3486 & ~n49608;
  assign n49610 = n3476 & ~n49609;
  assign n49611 = ~n49602 & ~n49610;
  assign n49612 = ~n3374 & ~n49611;
  assign n49613 = ~n3950 & ~n49594;
  assign n49614 = ~n3378 & ~n49613;
  assign n49615 = ~n3378 & ~n49614;
  assign n49616 = n3492 & ~n49615;
  assign n49617 = ~n3493 & ~n49616;
  assign n49618 = n3485 & ~n49617;
  assign n49619 = ~n3486 & ~n49618;
  assign n49620 = ~n3476 & ~n49619;
  assign n49621 = ~n3281 & ~n38065;
  assign n49622 = n3378 & ~n49621;
  assign n49623 = ~n38067 & ~n49622;
  assign n49624 = n3492 & ~n49623;
  assign n49625 = ~n3493 & ~n49624;
  assign n49626 = n3485 & ~n49625;
  assign n49627 = ~n3486 & ~n49626;
  assign n49628 = n3476 & ~n49627;
  assign n49629 = ~n49620 & ~n49628;
  assign n49630 = n3374 & ~n49629;
  assign n49631 = ~n49612 & ~n49630;
  assign n49632 = ~n3655 & ~n49631;
  assign n49633 = ~n49584 & ~n49632;
  assign n49634 = ~n3652 & ~n49633;
  assign n49635 = ~n49536 & ~n49634;
  assign n49636 = ~n3368 & ~n49635;
  assign n49637 = n3492 & ~n38113;
  assign n49638 = n3492 & ~n49637;
  assign n49639 = n3485 & ~n49638;
  assign n49640 = n3485 & ~n49639;
  assign n49641 = n3476 & ~n49640;
  assign n49642 = n3476 & ~n49641;
  assign n49643 = ~n3374 & ~n49642;
  assign n49644 = n3492 & ~n38370;
  assign n49645 = n3492 & ~n49644;
  assign n49646 = n3485 & ~n49645;
  assign n49647 = n3485 & ~n49646;
  assign n49648 = n3476 & ~n49647;
  assign n49649 = n3476 & ~n49648;
  assign n49650 = n3374 & ~n49649;
  assign n49651 = ~n49643 & ~n49650;
  assign n49652 = n3655 & ~n49651;
  assign n49653 = n3492 & ~n38412;
  assign n49654 = n3492 & ~n49653;
  assign n49655 = n3485 & ~n49654;
  assign n49656 = n3485 & ~n49655;
  assign n49657 = n3476 & ~n49656;
  assign n49658 = n3476 & ~n49657;
  assign n49659 = ~n3374 & ~n49658;
  assign n49660 = n3492 & ~n38658;
  assign n49661 = n3492 & ~n49660;
  assign n49662 = n3485 & ~n49661;
  assign n49663 = n3485 & ~n49662;
  assign n49664 = n3476 & ~n49663;
  assign n49665 = n3476 & ~n49664;
  assign n49666 = n3374 & ~n49665;
  assign n49667 = ~n49659 & ~n49666;
  assign n49668 = ~n3655 & ~n49667;
  assign n49669 = ~n49652 & ~n49668;
  assign n49670 = n3652 & ~n49669;
  assign n49671 = n3492 & ~n38695;
  assign n49672 = n3492 & ~n49671;
  assign n49673 = n3485 & ~n49672;
  assign n49674 = n3485 & ~n49673;
  assign n49675 = n3476 & ~n49674;
  assign n49676 = n3476 & ~n49675;
  assign n49677 = ~n3374 & ~n49676;
  assign n49678 = n3492 & ~n38869;
  assign n49679 = n3492 & ~n49678;
  assign n49680 = n3485 & ~n49679;
  assign n49681 = n3485 & ~n49680;
  assign n49682 = n3476 & ~n49681;
  assign n49683 = n3476 & ~n49682;
  assign n49684 = n3374 & ~n49683;
  assign n49685 = ~n49677 & ~n49684;
  assign n49686 = n3655 & ~n49685;
  assign n49687 = n3492 & ~n38904;
  assign n49688 = n3492 & ~n49687;
  assign n49689 = n3485 & ~n49688;
  assign n49690 = n3485 & ~n49689;
  assign n49691 = n3476 & ~n49690;
  assign n49692 = n3476 & ~n49691;
  assign n49693 = ~n3374 & ~n49692;
  assign n49694 = n3492 & ~n39078;
  assign n49695 = n3492 & ~n49694;
  assign n49696 = n3485 & ~n49695;
  assign n49697 = n3485 & ~n49696;
  assign n49698 = n3476 & ~n49697;
  assign n49699 = n3476 & ~n49698;
  assign n49700 = n3374 & ~n49699;
  assign n49701 = ~n49693 & ~n49700;
  assign n49702 = ~n3655 & ~n49701;
  assign n49703 = ~n49686 & ~n49702;
  assign n49704 = ~n3652 & ~n49703;
  assign n49705 = ~n49670 & ~n49704;
  assign n49706 = n3368 & ~n49705;
  assign n49707 = ~n49636 & ~n49706;
  assign n49708 = ~n3362 & ~n49707;
  assign n49709 = ~n3362 & ~n49708;
  assign n49710 = ~n3359 & ~n49709;
  assign n49711 = ~n3359 & ~n49710;
  assign n49712 = n3356 & ~n49711;
  assign n49713 = n3492 & ~n37397;
  assign n49714 = ~n3631 & ~n49713;
  assign n49715 = n3485 & ~n49714;
  assign n49716 = ~n3630 & ~n49715;
  assign n49717 = ~n3374 & ~n49716;
  assign n49718 = n3492 & ~n37471;
  assign n49719 = ~n3631 & ~n49718;
  assign n49720 = n3485 & ~n49719;
  assign n49721 = ~n3630 & ~n49720;
  assign n49722 = ~n3476 & ~n49721;
  assign n49723 = n3492 & ~n37553;
  assign n49724 = ~n3631 & ~n49723;
  assign n49725 = n3485 & ~n49724;
  assign n49726 = ~n3630 & ~n49725;
  assign n49727 = n3476 & ~n49726;
  assign n49728 = ~n49722 & ~n49727;
  assign n49729 = n3374 & ~n49728;
  assign n49730 = ~n49717 & ~n49729;
  assign n49731 = n3655 & ~n49730;
  assign n49732 = n3492 & ~n37587;
  assign n49733 = ~n3631 & ~n49732;
  assign n49734 = n3485 & ~n49733;
  assign n49735 = ~n3630 & ~n49734;
  assign n49736 = ~n3374 & ~n49735;
  assign n49737 = n3492 & ~n37665;
  assign n49738 = ~n3631 & ~n49737;
  assign n49739 = n3485 & ~n49738;
  assign n49740 = ~n3630 & ~n49739;
  assign n49741 = ~n3476 & ~n49740;
  assign n49742 = n3492 & ~n37756;
  assign n49743 = ~n3631 & ~n49742;
  assign n49744 = n3485 & ~n49743;
  assign n49745 = ~n3630 & ~n49744;
  assign n49746 = n3476 & ~n49745;
  assign n49747 = ~n49741 & ~n49746;
  assign n49748 = n3374 & ~n49747;
  assign n49749 = ~n49736 & ~n49748;
  assign n49750 = ~n3655 & ~n49749;
  assign n49751 = ~n49731 & ~n49750;
  assign n49752 = n3652 & ~n49751;
  assign n49753 = n3492 & ~n37790;
  assign n49754 = ~n3631 & ~n49753;
  assign n49755 = n3485 & ~n49754;
  assign n49756 = ~n3630 & ~n49755;
  assign n49757 = ~n3374 & ~n49756;
  assign n49758 = n3492 & ~n37850;
  assign n49759 = ~n3631 & ~n49758;
  assign n49760 = n3485 & ~n49759;
  assign n49761 = ~n3630 & ~n49760;
  assign n49762 = ~n3476 & ~n49761;
  assign n49763 = n3492 & ~n37912;
  assign n49764 = ~n3631 & ~n49763;
  assign n49765 = n3485 & ~n49764;
  assign n49766 = ~n3630 & ~n49765;
  assign n49767 = n3476 & ~n49766;
  assign n49768 = ~n49762 & ~n49767;
  assign n49769 = n3374 & ~n49768;
  assign n49770 = ~n49757 & ~n49769;
  assign n49771 = n3655 & ~n49770;
  assign n49772 = n3492 & ~n37944;
  assign n49773 = ~n3631 & ~n49772;
  assign n49774 = n3485 & ~n49773;
  assign n49775 = ~n3630 & ~n49774;
  assign n49776 = ~n3374 & ~n49775;
  assign n49777 = n3492 & ~n38004;
  assign n49778 = ~n3631 & ~n49777;
  assign n49779 = n3485 & ~n49778;
  assign n49780 = ~n3630 & ~n49779;
  assign n49781 = ~n3476 & ~n49780;
  assign n49782 = n3492 & ~n38066;
  assign n49783 = ~n3631 & ~n49782;
  assign n49784 = n3485 & ~n49783;
  assign n49785 = ~n3630 & ~n49784;
  assign n49786 = n3476 & ~n49785;
  assign n49787 = ~n49781 & ~n49786;
  assign n49788 = n3374 & ~n49787;
  assign n49789 = ~n49776 & ~n49788;
  assign n49790 = ~n3655 & ~n49789;
  assign n49791 = ~n49771 & ~n49790;
  assign n49792 = ~n3652 & ~n49791;
  assign n49793 = ~n49752 & ~n49792;
  assign n49794 = ~n3368 & ~n49793;
  assign n49795 = ~n3374 & ~n49640;
  assign n49796 = n3492 & ~n38185;
  assign n49797 = n3492 & ~n49796;
  assign n49798 = n3485 & ~n49797;
  assign n49799 = n3485 & ~n49798;
  assign n49800 = ~n3476 & ~n49799;
  assign n49801 = ~n49648 & ~n49800;
  assign n49802 = n3374 & ~n49801;
  assign n49803 = ~n49795 & ~n49802;
  assign n49804 = n3655 & ~n49803;
  assign n49805 = ~n3374 & ~n49656;
  assign n49806 = n3492 & ~n38484;
  assign n49807 = n3492 & ~n49806;
  assign n49808 = n3485 & ~n49807;
  assign n49809 = n3485 & ~n49808;
  assign n49810 = ~n3476 & ~n49809;
  assign n49811 = ~n49664 & ~n49810;
  assign n49812 = n3374 & ~n49811;
  assign n49813 = ~n49805 & ~n49812;
  assign n49814 = ~n3655 & ~n49813;
  assign n49815 = ~n49804 & ~n49814;
  assign n49816 = n3652 & ~n49815;
  assign n49817 = ~n3374 & ~n49674;
  assign n49818 = n3492 & ~n38753;
  assign n49819 = n3492 & ~n49818;
  assign n49820 = n3485 & ~n49819;
  assign n49821 = n3485 & ~n49820;
  assign n49822 = ~n3476 & ~n49821;
  assign n49823 = ~n49682 & ~n49822;
  assign n49824 = n3374 & ~n49823;
  assign n49825 = ~n49817 & ~n49824;
  assign n49826 = n3655 & ~n49825;
  assign n49827 = ~n3374 & ~n49690;
  assign n49828 = n3492 & ~n38962;
  assign n49829 = n3492 & ~n49828;
  assign n49830 = n3485 & ~n49829;
  assign n49831 = n3485 & ~n49830;
  assign n49832 = ~n3476 & ~n49831;
  assign n49833 = ~n49698 & ~n49832;
  assign n49834 = n3374 & ~n49833;
  assign n49835 = ~n49827 & ~n49834;
  assign n49836 = ~n3655 & ~n49835;
  assign n49837 = ~n49826 & ~n49836;
  assign n49838 = ~n3652 & ~n49837;
  assign n49839 = ~n49816 & ~n49838;
  assign n49840 = n3368 & ~n49839;
  assign n49841 = ~n49794 & ~n49840;
  assign n49842 = n3362 & ~n49841;
  assign n49843 = ~n3476 & ~n49716;
  assign n49844 = ~n41076 & ~n49715;
  assign n49845 = n3476 & ~n49844;
  assign n49846 = ~n49843 & ~n49845;
  assign n49847 = ~n3374 & ~n49846;
  assign n49848 = ~n41076 & ~n49725;
  assign n49849 = n3476 & ~n49848;
  assign n49850 = ~n49722 & ~n49849;
  assign n49851 = n3374 & ~n49850;
  assign n49852 = ~n49847 & ~n49851;
  assign n49853 = n3655 & ~n49852;
  assign n49854 = ~n3476 & ~n49735;
  assign n49855 = ~n41101 & ~n49734;
  assign n49856 = n3476 & ~n49855;
  assign n49857 = ~n49854 & ~n49856;
  assign n49858 = ~n3374 & ~n49857;
  assign n49859 = ~n41101 & ~n49744;
  assign n49860 = n3476 & ~n49859;
  assign n49861 = ~n49741 & ~n49860;
  assign n49862 = n3374 & ~n49861;
  assign n49863 = ~n49858 & ~n49862;
  assign n49864 = ~n3655 & ~n49863;
  assign n49865 = ~n49853 & ~n49864;
  assign n49866 = n3652 & ~n49865;
  assign n49867 = ~n3476 & ~n49756;
  assign n49868 = ~n41128 & ~n49755;
  assign n49869 = n3476 & ~n49868;
  assign n49870 = ~n49867 & ~n49869;
  assign n49871 = ~n3374 & ~n49870;
  assign n49872 = ~n41128 & ~n49765;
  assign n49873 = n3476 & ~n49872;
  assign n49874 = ~n49762 & ~n49873;
  assign n49875 = n3374 & ~n49874;
  assign n49876 = ~n49871 & ~n49875;
  assign n49877 = n3655 & ~n49876;
  assign n49878 = ~n3476 & ~n49775;
  assign n49879 = ~n41153 & ~n49774;
  assign n49880 = n3476 & ~n49879;
  assign n49881 = ~n49878 & ~n49880;
  assign n49882 = ~n3374 & ~n49881;
  assign n49883 = ~n41153 & ~n49784;
  assign n49884 = n3476 & ~n49883;
  assign n49885 = ~n49781 & ~n49884;
  assign n49886 = n3374 & ~n49885;
  assign n49887 = ~n49882 & ~n49886;
  assign n49888 = ~n3655 & ~n49887;
  assign n49889 = ~n49877 & ~n49888;
  assign n49890 = ~n3652 & ~n49889;
  assign n49891 = ~n49866 & ~n49890;
  assign n49892 = ~n3368 & ~n49891;
  assign n49893 = ~n3476 & ~n49640;
  assign n49894 = ~n8525 & ~n49639;
  assign n49895 = n3476 & ~n49894;
  assign n49896 = ~n49893 & ~n49895;
  assign n49897 = ~n3374 & ~n49896;
  assign n49898 = ~n41191 & ~n49646;
  assign n49899 = n3476 & ~n49898;
  assign n49900 = ~n49800 & ~n49899;
  assign n49901 = n3374 & ~n49900;
  assign n49902 = ~n49897 & ~n49901;
  assign n49903 = n3655 & ~n49902;
  assign n49904 = ~n3476 & ~n49656;
  assign n49905 = ~n8525 & ~n49655;
  assign n49906 = n3476 & ~n49905;
  assign n49907 = ~n49904 & ~n49906;
  assign n49908 = ~n3374 & ~n49907;
  assign n49909 = ~n41216 & ~n49662;
  assign n49910 = n3476 & ~n49909;
  assign n49911 = ~n49810 & ~n49910;
  assign n49912 = n3374 & ~n49911;
  assign n49913 = ~n49908 & ~n49912;
  assign n49914 = ~n3655 & ~n49913;
  assign n49915 = ~n49903 & ~n49914;
  assign n49916 = n3652 & ~n49915;
  assign n49917 = ~n3476 & ~n49674;
  assign n49918 = ~n8525 & ~n49673;
  assign n49919 = n3476 & ~n49918;
  assign n49920 = ~n49917 & ~n49919;
  assign n49921 = ~n3374 & ~n49920;
  assign n49922 = ~n41243 & ~n49680;
  assign n49923 = n3476 & ~n49922;
  assign n49924 = ~n49822 & ~n49923;
  assign n49925 = n3374 & ~n49924;
  assign n49926 = ~n49921 & ~n49925;
  assign n49927 = n3655 & ~n49926;
  assign n49928 = ~n3476 & ~n49690;
  assign n49929 = ~n8525 & ~n49689;
  assign n49930 = n3476 & ~n49929;
  assign n49931 = ~n49928 & ~n49930;
  assign n49932 = ~n3374 & ~n49931;
  assign n49933 = ~n41268 & ~n49696;
  assign n49934 = n3476 & ~n49933;
  assign n49935 = ~n49832 & ~n49934;
  assign n49936 = n3374 & ~n49935;
  assign n49937 = ~n49932 & ~n49936;
  assign n49938 = ~n3655 & ~n49937;
  assign n49939 = ~n49927 & ~n49938;
  assign n49940 = ~n3652 & ~n49939;
  assign n49941 = ~n49916 & ~n49940;
  assign n49942 = n3368 & ~n49941;
  assign n49943 = ~n49892 & ~n49942;
  assign n49944 = ~n3362 & ~n49943;
  assign n49945 = ~n49842 & ~n49944;
  assign n49946 = n3359 & ~n49945;
  assign n49947 = ~n37278 & ~n49715;
  assign n49948 = n3476 & ~n49947;
  assign n49949 = ~n49843 & ~n49948;
  assign n49950 = ~n3374 & ~n49949;
  assign n49951 = ~n37278 & ~n49725;
  assign n49952 = n3476 & ~n49951;
  assign n49953 = ~n49722 & ~n49952;
  assign n49954 = n3374 & ~n49953;
  assign n49955 = ~n49950 & ~n49954;
  assign n49956 = n3655 & ~n49955;
  assign n49957 = ~n37289 & ~n49734;
  assign n49958 = n3476 & ~n49957;
  assign n49959 = ~n49854 & ~n49958;
  assign n49960 = ~n3374 & ~n49959;
  assign n49961 = ~n37289 & ~n49744;
  assign n49962 = n3476 & ~n49961;
  assign n49963 = ~n49741 & ~n49962;
  assign n49964 = n3374 & ~n49963;
  assign n49965 = ~n49960 & ~n49964;
  assign n49966 = ~n3655 & ~n49965;
  assign n49967 = ~n49956 & ~n49966;
  assign n49968 = n3652 & ~n49967;
  assign n49969 = ~n37302 & ~n49755;
  assign n49970 = n3476 & ~n49969;
  assign n49971 = ~n49867 & ~n49970;
  assign n49972 = ~n3374 & ~n49971;
  assign n49973 = ~n37302 & ~n49765;
  assign n49974 = n3476 & ~n49973;
  assign n49975 = ~n49762 & ~n49974;
  assign n49976 = n3374 & ~n49975;
  assign n49977 = ~n49972 & ~n49976;
  assign n49978 = n3655 & ~n49977;
  assign n49979 = ~n37313 & ~n49774;
  assign n49980 = n3476 & ~n49979;
  assign n49981 = ~n49878 & ~n49980;
  assign n49982 = ~n3374 & ~n49981;
  assign n49983 = ~n37313 & ~n49784;
  assign n49984 = n3476 & ~n49983;
  assign n49985 = ~n49781 & ~n49984;
  assign n49986 = n3374 & ~n49985;
  assign n49987 = ~n49982 & ~n49986;
  assign n49988 = ~n3655 & ~n49987;
  assign n49989 = ~n49978 & ~n49988;
  assign n49990 = ~n3652 & ~n49989;
  assign n49991 = ~n49968 & ~n49990;
  assign n49992 = ~n3368 & ~n49991;
  assign n49993 = ~n8689 & ~n49639;
  assign n49994 = n3476 & ~n49993;
  assign n49995 = ~n49893 & ~n49994;
  assign n49996 = ~n3374 & ~n49995;
  assign n49997 = ~n37332 & ~n49646;
  assign n49998 = n3476 & ~n49997;
  assign n49999 = ~n49800 & ~n49998;
  assign n50000 = n3374 & ~n49999;
  assign n50001 = ~n49996 & ~n50000;
  assign n50002 = n3655 & ~n50001;
  assign n50003 = ~n8689 & ~n49655;
  assign n50004 = n3476 & ~n50003;
  assign n50005 = ~n49904 & ~n50004;
  assign n50006 = ~n3374 & ~n50005;
  assign n50007 = ~n37343 & ~n49662;
  assign n50008 = n3476 & ~n50007;
  assign n50009 = ~n49810 & ~n50008;
  assign n50010 = n3374 & ~n50009;
  assign n50011 = ~n50006 & ~n50010;
  assign n50012 = ~n3655 & ~n50011;
  assign n50013 = ~n50002 & ~n50012;
  assign n50014 = n3652 & ~n50013;
  assign n50015 = ~n8689 & ~n49673;
  assign n50016 = n3476 & ~n50015;
  assign n50017 = ~n49917 & ~n50016;
  assign n50018 = ~n3374 & ~n50017;
  assign n50019 = ~n37356 & ~n49680;
  assign n50020 = n3476 & ~n50019;
  assign n50021 = ~n49822 & ~n50020;
  assign n50022 = n3374 & ~n50021;
  assign n50023 = ~n50018 & ~n50022;
  assign n50024 = n3655 & ~n50023;
  assign n50025 = ~n8689 & ~n49689;
  assign n50026 = n3476 & ~n50025;
  assign n50027 = ~n49928 & ~n50026;
  assign n50028 = ~n3374 & ~n50027;
  assign n50029 = ~n37367 & ~n49696;
  assign n50030 = n3476 & ~n50029;
  assign n50031 = ~n49832 & ~n50030;
  assign n50032 = n3374 & ~n50031;
  assign n50033 = ~n50028 & ~n50032;
  assign n50034 = ~n3655 & ~n50033;
  assign n50035 = ~n50024 & ~n50034;
  assign n50036 = ~n3652 & ~n50035;
  assign n50037 = ~n50014 & ~n50036;
  assign n50038 = n3368 & ~n50037;
  assign n50039 = ~n49992 & ~n50038;
  assign n50040 = n3362 & ~n50039;
  assign n50041 = ~n37006 & ~n49713;
  assign n50042 = n3485 & ~n50041;
  assign n50043 = ~n37278 & ~n50042;
  assign n50044 = n3476 & ~n50043;
  assign n50045 = ~n49843 & ~n50044;
  assign n50046 = ~n3374 & ~n50045;
  assign n50047 = ~n37006 & ~n49723;
  assign n50048 = n3485 & ~n50047;
  assign n50049 = ~n37278 & ~n50048;
  assign n50050 = n3476 & ~n50049;
  assign n50051 = ~n49722 & ~n50050;
  assign n50052 = n3374 & ~n50051;
  assign n50053 = ~n50046 & ~n50052;
  assign n50054 = n3655 & ~n50053;
  assign n50055 = ~n37048 & ~n49732;
  assign n50056 = n3485 & ~n50055;
  assign n50057 = ~n37289 & ~n50056;
  assign n50058 = n3476 & ~n50057;
  assign n50059 = ~n49854 & ~n50058;
  assign n50060 = ~n3374 & ~n50059;
  assign n50061 = ~n37048 & ~n49742;
  assign n50062 = n3485 & ~n50061;
  assign n50063 = ~n37289 & ~n50062;
  assign n50064 = n3476 & ~n50063;
  assign n50065 = ~n49741 & ~n50064;
  assign n50066 = n3374 & ~n50065;
  assign n50067 = ~n50060 & ~n50066;
  assign n50068 = ~n3655 & ~n50067;
  assign n50069 = ~n50054 & ~n50068;
  assign n50070 = n3652 & ~n50069;
  assign n50071 = ~n37091 & ~n49753;
  assign n50072 = n3485 & ~n50071;
  assign n50073 = ~n37302 & ~n50072;
  assign n50074 = n3476 & ~n50073;
  assign n50075 = ~n49867 & ~n50074;
  assign n50076 = ~n3374 & ~n50075;
  assign n50077 = ~n37091 & ~n49763;
  assign n50078 = n3485 & ~n50077;
  assign n50079 = ~n37302 & ~n50078;
  assign n50080 = n3476 & ~n50079;
  assign n50081 = ~n49762 & ~n50080;
  assign n50082 = n3374 & ~n50081;
  assign n50083 = ~n50076 & ~n50082;
  assign n50084 = n3655 & ~n50083;
  assign n50085 = ~n37132 & ~n49772;
  assign n50086 = n3485 & ~n50085;
  assign n50087 = ~n37313 & ~n50086;
  assign n50088 = n3476 & ~n50087;
  assign n50089 = ~n49878 & ~n50088;
  assign n50090 = ~n3374 & ~n50089;
  assign n50091 = ~n37132 & ~n49782;
  assign n50092 = n3485 & ~n50091;
  assign n50093 = ~n37313 & ~n50092;
  assign n50094 = n3476 & ~n50093;
  assign n50095 = ~n49781 & ~n50094;
  assign n50096 = n3374 & ~n50095;
  assign n50097 = ~n50090 & ~n50096;
  assign n50098 = ~n3655 & ~n50097;
  assign n50099 = ~n50084 & ~n50098;
  assign n50100 = ~n3652 & ~n50099;
  assign n50101 = ~n50070 & ~n50100;
  assign n50102 = ~n3368 & ~n50101;
  assign n50103 = ~n8523 & ~n49637;
  assign n50104 = n3485 & ~n50103;
  assign n50105 = ~n8689 & ~n50104;
  assign n50106 = n3476 & ~n50105;
  assign n50107 = ~n49893 & ~n50106;
  assign n50108 = ~n3374 & ~n50107;
  assign n50109 = ~n37174 & ~n49644;
  assign n50110 = n3485 & ~n50109;
  assign n50111 = ~n37332 & ~n50110;
  assign n50112 = n3476 & ~n50111;
  assign n50113 = ~n49800 & ~n50112;
  assign n50114 = n3374 & ~n50113;
  assign n50115 = ~n50108 & ~n50114;
  assign n50116 = n3655 & ~n50115;
  assign n50117 = ~n8523 & ~n49653;
  assign n50118 = n3485 & ~n50117;
  assign n50119 = ~n8689 & ~n50118;
  assign n50120 = n3476 & ~n50119;
  assign n50121 = ~n49904 & ~n50120;
  assign n50122 = ~n3374 & ~n50121;
  assign n50123 = ~n37202 & ~n49660;
  assign n50124 = n3485 & ~n50123;
  assign n50125 = ~n37343 & ~n50124;
  assign n50126 = n3476 & ~n50125;
  assign n50127 = ~n49810 & ~n50126;
  assign n50128 = n3374 & ~n50127;
  assign n50129 = ~n50122 & ~n50128;
  assign n50130 = ~n3655 & ~n50129;
  assign n50131 = ~n50116 & ~n50130;
  assign n50132 = n3652 & ~n50131;
  assign n50133 = ~n8523 & ~n49671;
  assign n50134 = n3485 & ~n50133;
  assign n50135 = ~n8689 & ~n50134;
  assign n50136 = n3476 & ~n50135;
  assign n50137 = ~n49917 & ~n50136;
  assign n50138 = ~n3374 & ~n50137;
  assign n50139 = ~n37231 & ~n49678;
  assign n50140 = n3485 & ~n50139;
  assign n50141 = ~n37356 & ~n50140;
  assign n50142 = n3476 & ~n50141;
  assign n50143 = ~n49822 & ~n50142;
  assign n50144 = n3374 & ~n50143;
  assign n50145 = ~n50138 & ~n50144;
  assign n50146 = n3655 & ~n50145;
  assign n50147 = ~n8523 & ~n49687;
  assign n50148 = n3485 & ~n50147;
  assign n50149 = ~n8689 & ~n50148;
  assign n50150 = n3476 & ~n50149;
  assign n50151 = ~n49928 & ~n50150;
  assign n50152 = ~n3374 & ~n50151;
  assign n50153 = ~n37258 & ~n49694;
  assign n50154 = n3485 & ~n50153;
  assign n50155 = ~n37367 & ~n50154;
  assign n50156 = n3476 & ~n50155;
  assign n50157 = ~n49832 & ~n50156;
  assign n50158 = n3374 & ~n50157;
  assign n50159 = ~n50152 & ~n50158;
  assign n50160 = ~n3655 & ~n50159;
  assign n50161 = ~n50146 & ~n50160;
  assign n50162 = ~n3652 & ~n50161;
  assign n50163 = ~n50132 & ~n50162;
  assign n50164 = n3368 & ~n50163;
  assign n50165 = ~n50102 & ~n50164;
  assign n50166 = ~n3362 & ~n50165;
  assign n50167 = ~n50040 & ~n50166;
  assign n50168 = ~n3359 & ~n50167;
  assign n50169 = ~n49946 & ~n50168;
  assign n50170 = ~n3356 & ~n50169;
  assign n50171 = ~n49712 & ~n50170;
  assign n50172 = ~n3345 & ~n50171;
  assign n50173 = ~n3378 & ~n37398;
  assign n50174 = n3492 & ~n50173;
  assign n50175 = ~n3493 & ~n50174;
  assign n50176 = n3485 & ~n50175;
  assign n50177 = ~n3486 & ~n50176;
  assign n50178 = ~n3476 & ~n50177;
  assign n50179 = ~n3378 & ~n37005;
  assign n50180 = ~n3378 & ~n50179;
  assign n50181 = ~n3485 & ~n50180;
  assign n50182 = ~n3492 & ~n50180;
  assign n50183 = ~n50174 & ~n50182;
  assign n50184 = n3485 & ~n50183;
  assign n50185 = ~n50181 & ~n50184;
  assign n50186 = n3476 & ~n50185;
  assign n50187 = ~n50178 & ~n50186;
  assign n50188 = ~n3374 & ~n50187;
  assign n50189 = ~n3281 & ~n37470;
  assign n50190 = n3378 & ~n50189;
  assign n50191 = ~n37472 & ~n50190;
  assign n50192 = n3492 & ~n50191;
  assign n50193 = ~n25115 & ~n50192;
  assign n50194 = n3485 & ~n50193;
  assign n50195 = ~n25114 & ~n50194;
  assign n50196 = ~n3476 & ~n50195;
  assign n50197 = n3378 & ~n37173;
  assign n50198 = ~n50179 & ~n50197;
  assign n50199 = ~n3485 & ~n50198;
  assign n50200 = ~n3492 & ~n50198;
  assign n50201 = ~n49478 & ~n50200;
  assign n50202 = n3485 & ~n50201;
  assign n50203 = ~n50199 & ~n50202;
  assign n50204 = n3476 & ~n50203;
  assign n50205 = ~n50196 & ~n50204;
  assign n50206 = n3374 & ~n50205;
  assign n50207 = ~n50188 & ~n50206;
  assign n50208 = n3655 & ~n50207;
  assign n50209 = ~n3378 & ~n37588;
  assign n50210 = n3492 & ~n50209;
  assign n50211 = ~n3493 & ~n50210;
  assign n50212 = n3485 & ~n50211;
  assign n50213 = ~n3486 & ~n50212;
  assign n50214 = ~n3476 & ~n50213;
  assign n50215 = ~n3378 & ~n37047;
  assign n50216 = ~n3378 & ~n50215;
  assign n50217 = ~n3485 & ~n50216;
  assign n50218 = ~n3492 & ~n50216;
  assign n50219 = ~n50210 & ~n50218;
  assign n50220 = n3485 & ~n50219;
  assign n50221 = ~n50217 & ~n50220;
  assign n50222 = n3476 & ~n50221;
  assign n50223 = ~n50214 & ~n50222;
  assign n50224 = ~n3374 & ~n50223;
  assign n50225 = ~n3281 & ~n37664;
  assign n50226 = n3378 & ~n50225;
  assign n50227 = ~n37666 & ~n50226;
  assign n50228 = n3492 & ~n50227;
  assign n50229 = ~n25115 & ~n50228;
  assign n50230 = n3485 & ~n50229;
  assign n50231 = ~n25114 & ~n50230;
  assign n50232 = ~n3476 & ~n50231;
  assign n50233 = n3378 & ~n37201;
  assign n50234 = ~n50215 & ~n50233;
  assign n50235 = ~n3485 & ~n50234;
  assign n50236 = ~n3492 & ~n50234;
  assign n50237 = ~n49526 & ~n50236;
  assign n50238 = n3485 & ~n50237;
  assign n50239 = ~n50235 & ~n50238;
  assign n50240 = n3476 & ~n50239;
  assign n50241 = ~n50232 & ~n50240;
  assign n50242 = n3374 & ~n50241;
  assign n50243 = ~n50224 & ~n50242;
  assign n50244 = ~n3655 & ~n50243;
  assign n50245 = ~n50208 & ~n50244;
  assign n50246 = n3652 & ~n50245;
  assign n50247 = ~n3378 & ~n37791;
  assign n50248 = n3492 & ~n50247;
  assign n50249 = ~n3493 & ~n50248;
  assign n50250 = n3485 & ~n50249;
  assign n50251 = ~n3486 & ~n50250;
  assign n50252 = ~n3476 & ~n50251;
  assign n50253 = ~n3378 & ~n37090;
  assign n50254 = ~n3378 & ~n50253;
  assign n50255 = ~n3485 & ~n50254;
  assign n50256 = ~n3492 & ~n50254;
  assign n50257 = ~n50248 & ~n50256;
  assign n50258 = n3485 & ~n50257;
  assign n50259 = ~n50255 & ~n50258;
  assign n50260 = n3476 & ~n50259;
  assign n50261 = ~n50252 & ~n50260;
  assign n50262 = ~n3374 & ~n50261;
  assign n50263 = ~n3281 & ~n37849;
  assign n50264 = n3378 & ~n50263;
  assign n50265 = ~n37851 & ~n50264;
  assign n50266 = n3492 & ~n50265;
  assign n50267 = ~n25115 & ~n50266;
  assign n50268 = n3485 & ~n50267;
  assign n50269 = ~n25114 & ~n50268;
  assign n50270 = ~n3476 & ~n50269;
  assign n50271 = n3378 & ~n37230;
  assign n50272 = ~n50253 & ~n50271;
  assign n50273 = ~n3485 & ~n50272;
  assign n50274 = ~n3492 & ~n50272;
  assign n50275 = ~n49576 & ~n50274;
  assign n50276 = n3485 & ~n50275;
  assign n50277 = ~n50273 & ~n50276;
  assign n50278 = n3476 & ~n50277;
  assign n50279 = ~n50270 & ~n50278;
  assign n50280 = n3374 & ~n50279;
  assign n50281 = ~n50262 & ~n50280;
  assign n50282 = n3655 & ~n50281;
  assign n50283 = ~n3378 & ~n37945;
  assign n50284 = n3492 & ~n50283;
  assign n50285 = ~n3493 & ~n50284;
  assign n50286 = n3485 & ~n50285;
  assign n50287 = ~n3486 & ~n50286;
  assign n50288 = ~n3476 & ~n50287;
  assign n50289 = ~n3378 & ~n37131;
  assign n50290 = ~n3378 & ~n50289;
  assign n50291 = ~n3485 & ~n50290;
  assign n50292 = ~n3492 & ~n50290;
  assign n50293 = ~n50284 & ~n50292;
  assign n50294 = n3485 & ~n50293;
  assign n50295 = ~n50291 & ~n50294;
  assign n50296 = n3476 & ~n50295;
  assign n50297 = ~n50288 & ~n50296;
  assign n50298 = ~n3374 & ~n50297;
  assign n50299 = ~n3281 & ~n38003;
  assign n50300 = n3378 & ~n50299;
  assign n50301 = ~n38005 & ~n50300;
  assign n50302 = n3492 & ~n50301;
  assign n50303 = ~n25115 & ~n50302;
  assign n50304 = n3485 & ~n50303;
  assign n50305 = ~n25114 & ~n50304;
  assign n50306 = ~n3476 & ~n50305;
  assign n50307 = n3378 & ~n37257;
  assign n50308 = ~n50289 & ~n50307;
  assign n50309 = ~n3485 & ~n50308;
  assign n50310 = ~n3492 & ~n50308;
  assign n50311 = ~n49624 & ~n50310;
  assign n50312 = n3485 & ~n50311;
  assign n50313 = ~n50309 & ~n50312;
  assign n50314 = n3476 & ~n50313;
  assign n50315 = ~n50306 & ~n50314;
  assign n50316 = n3374 & ~n50315;
  assign n50317 = ~n50298 & ~n50316;
  assign n50318 = ~n3655 & ~n50317;
  assign n50319 = ~n50282 & ~n50318;
  assign n50320 = ~n3652 & ~n50319;
  assign n50321 = ~n50246 & ~n50320;
  assign n50322 = ~n3368 & ~n50321;
  assign n50323 = ~n3378 & ~n38114;
  assign n50324 = n3492 & ~n50323;
  assign n50325 = n3492 & ~n50324;
  assign n50326 = n3485 & ~n50325;
  assign n50327 = n3485 & ~n50326;
  assign n50328 = ~n3476 & ~n50327;
  assign n50329 = ~n25259 & ~n50324;
  assign n50330 = n3485 & ~n50329;
  assign n50331 = ~n25258 & ~n50330;
  assign n50332 = n3476 & ~n50331;
  assign n50333 = ~n50328 & ~n50332;
  assign n50334 = ~n3374 & ~n50333;
  assign n50335 = ~n50114 & ~n50334;
  assign n50336 = n3655 & ~n50335;
  assign n50337 = ~n3378 & ~n38413;
  assign n50338 = n3492 & ~n50337;
  assign n50339 = n3492 & ~n50338;
  assign n50340 = n3485 & ~n50339;
  assign n50341 = n3485 & ~n50340;
  assign n50342 = ~n3476 & ~n50341;
  assign n50343 = ~n25259 & ~n50338;
  assign n50344 = n3485 & ~n50343;
  assign n50345 = ~n25258 & ~n50344;
  assign n50346 = n3476 & ~n50345;
  assign n50347 = ~n50342 & ~n50346;
  assign n50348 = ~n3374 & ~n50347;
  assign n50349 = ~n50128 & ~n50348;
  assign n50350 = ~n3655 & ~n50349;
  assign n50351 = ~n50336 & ~n50350;
  assign n50352 = n3652 & ~n50351;
  assign n50353 = ~n3378 & ~n38696;
  assign n50354 = n3492 & ~n50353;
  assign n50355 = n3492 & ~n50354;
  assign n50356 = n3485 & ~n50355;
  assign n50357 = n3485 & ~n50356;
  assign n50358 = ~n3476 & ~n50357;
  assign n50359 = ~n25259 & ~n50354;
  assign n50360 = n3485 & ~n50359;
  assign n50361 = ~n25258 & ~n50360;
  assign n50362 = n3476 & ~n50361;
  assign n50363 = ~n50358 & ~n50362;
  assign n50364 = ~n3374 & ~n50363;
  assign n50365 = ~n50144 & ~n50364;
  assign n50366 = n3655 & ~n50365;
  assign n50367 = ~n3378 & ~n38905;
  assign n50368 = n3492 & ~n50367;
  assign n50369 = n3492 & ~n50368;
  assign n50370 = n3485 & ~n50369;
  assign n50371 = n3485 & ~n50370;
  assign n50372 = ~n3476 & ~n50371;
  assign n50373 = ~n25259 & ~n50368;
  assign n50374 = n3485 & ~n50373;
  assign n50375 = ~n25258 & ~n50374;
  assign n50376 = n3476 & ~n50375;
  assign n50377 = ~n50372 & ~n50376;
  assign n50378 = ~n3374 & ~n50377;
  assign n50379 = ~n50158 & ~n50378;
  assign n50380 = ~n3655 & ~n50379;
  assign n50381 = ~n50366 & ~n50380;
  assign n50382 = ~n3652 & ~n50381;
  assign n50383 = ~n50352 & ~n50382;
  assign n50384 = n3368 & ~n50383;
  assign n50385 = ~n50322 & ~n50384;
  assign n50386 = ~n3362 & ~n50385;
  assign n50387 = ~n3362 & ~n50386;
  assign n50388 = ~n3359 & ~n50387;
  assign n50389 = ~n3359 & ~n50388;
  assign n50390 = n3356 & ~n50389;
  assign n50391 = ~n3356 & ~n50165;
  assign n50392 = ~n50390 & ~n50391;
  assign n50393 = n3345 & ~n50392;
  assign n50394 = ~n50172 & ~n50393;
  assign n50395 = n3341 & ~n50394;
  assign n50396 = ~n49438 & ~n50395;
  assign n50397 = n3337 & ~n50396;
  assign n50398 = ~n44353 & ~n50397;
  assign n50399 = n3280 & ~n50398;
  assign n50400 = ~n25331 & ~n34145;
  assign n50401 = controllable_nhgrant0 & ~n50400;
  assign n50402 = ~n3945 & ~n50401;
  assign n50403 = ~n3281 & ~n50402;
  assign n50404 = ~n3281 & ~n50403;
  assign n50405 = n3378 & ~n50404;
  assign n50406 = ~n25338 & ~n34176;
  assign n50407 = controllable_nhgrant0 & ~n50406;
  assign n50408 = ~n3987 & ~n50407;
  assign n50409 = ~n3281 & ~n50408;
  assign n50410 = ~n3950 & ~n50409;
  assign n50411 = ~n3378 & ~n50410;
  assign n50412 = ~n50405 & ~n50411;
  assign n50413 = n3492 & ~n50412;
  assign n50414 = ~n3493 & ~n50413;
  assign n50415 = n3485 & ~n50414;
  assign n50416 = ~n3486 & ~n50415;
  assign n50417 = ~n3476 & ~n50416;
  assign n50418 = ~n25331 & ~n34232;
  assign n50419 = controllable_nhgrant0 & ~n50418;
  assign n50420 = ~n3945 & ~n50419;
  assign n50421 = ~n3281 & ~n50420;
  assign n50422 = ~n3281 & ~n50421;
  assign n50423 = n3378 & ~n50422;
  assign n50424 = ~n25338 & ~n34289;
  assign n50425 = controllable_nhgrant0 & ~n50424;
  assign n50426 = ~n3987 & ~n50425;
  assign n50427 = ~n3281 & ~n50426;
  assign n50428 = ~n4089 & ~n50427;
  assign n50429 = ~n3378 & ~n50428;
  assign n50430 = ~n50423 & ~n50429;
  assign n50431 = n3492 & ~n50430;
  assign n50432 = ~n34114 & ~n50431;
  assign n50433 = n3485 & ~n50432;
  assign n50434 = ~n34113 & ~n50433;
  assign n50435 = n3476 & ~n50434;
  assign n50436 = ~n50417 & ~n50435;
  assign n50437 = n3374 & ~n50436;
  assign n50438 = ~n34120 & ~n50437;
  assign n50439 = n3655 & ~n50438;
  assign n50440 = ~n25331 & ~n34328;
  assign n50441 = controllable_nhgrant0 & ~n50440;
  assign n50442 = ~n3945 & ~n50441;
  assign n50443 = ~n3281 & ~n50442;
  assign n50444 = ~n3281 & ~n50443;
  assign n50445 = n3378 & ~n50444;
  assign n50446 = ~n25338 & ~n34346;
  assign n50447 = controllable_nhgrant0 & ~n50446;
  assign n50448 = ~n3987 & ~n50447;
  assign n50449 = ~n3281 & ~n50448;
  assign n50450 = ~n3950 & ~n50449;
  assign n50451 = ~n3378 & ~n50450;
  assign n50452 = ~n50445 & ~n50451;
  assign n50453 = n3492 & ~n50452;
  assign n50454 = ~n3493 & ~n50453;
  assign n50455 = n3485 & ~n50454;
  assign n50456 = ~n3486 & ~n50455;
  assign n50457 = ~n3476 & ~n50456;
  assign n50458 = ~n25331 & ~n34381;
  assign n50459 = controllable_nhgrant0 & ~n50458;
  assign n50460 = ~n3945 & ~n50459;
  assign n50461 = ~n3281 & ~n50460;
  assign n50462 = ~n3281 & ~n50461;
  assign n50463 = n3378 & ~n50462;
  assign n50464 = ~n25338 & ~n34410;
  assign n50465 = controllable_nhgrant0 & ~n50464;
  assign n50466 = ~n3987 & ~n50465;
  assign n50467 = ~n3281 & ~n50466;
  assign n50468 = ~n4089 & ~n50467;
  assign n50469 = ~n3378 & ~n50468;
  assign n50470 = ~n50463 & ~n50469;
  assign n50471 = n3492 & ~n50470;
  assign n50472 = ~n34114 & ~n50471;
  assign n50473 = n3485 & ~n50472;
  assign n50474 = ~n34113 & ~n50473;
  assign n50475 = n3476 & ~n50474;
  assign n50476 = ~n50457 & ~n50475;
  assign n50477 = n3374 & ~n50476;
  assign n50478 = ~n34120 & ~n50477;
  assign n50479 = ~n3655 & ~n50478;
  assign n50480 = ~n50439 & ~n50479;
  assign n50481 = n3652 & ~n50480;
  assign n50482 = ~n25331 & ~n34444;
  assign n50483 = controllable_nhgrant0 & ~n50482;
  assign n50484 = ~n3945 & ~n50483;
  assign n50485 = ~n3281 & ~n50484;
  assign n50486 = ~n3281 & ~n50485;
  assign n50487 = n3378 & ~n50486;
  assign n50488 = ~n25338 & ~n34462;
  assign n50489 = controllable_nhgrant0 & ~n50488;
  assign n50490 = ~n3987 & ~n50489;
  assign n50491 = ~n3281 & ~n50490;
  assign n50492 = ~n3950 & ~n50491;
  assign n50493 = ~n3378 & ~n50492;
  assign n50494 = ~n50487 & ~n50493;
  assign n50495 = n3492 & ~n50494;
  assign n50496 = ~n3493 & ~n50495;
  assign n50497 = n3485 & ~n50496;
  assign n50498 = ~n3486 & ~n50497;
  assign n50499 = ~n3476 & ~n50498;
  assign n50500 = ~n25331 & ~n34490;
  assign n50501 = controllable_nhgrant0 & ~n50500;
  assign n50502 = ~n3945 & ~n50501;
  assign n50503 = ~n3281 & ~n50502;
  assign n50504 = ~n3281 & ~n50503;
  assign n50505 = n3378 & ~n50504;
  assign n50506 = ~n25338 & ~n34512;
  assign n50507 = controllable_nhgrant0 & ~n50506;
  assign n50508 = ~n3987 & ~n50507;
  assign n50509 = ~n3281 & ~n50508;
  assign n50510 = ~n4089 & ~n50509;
  assign n50511 = ~n3378 & ~n50510;
  assign n50512 = ~n50505 & ~n50511;
  assign n50513 = n3492 & ~n50512;
  assign n50514 = ~n34114 & ~n50513;
  assign n50515 = n3485 & ~n50514;
  assign n50516 = ~n34113 & ~n50515;
  assign n50517 = n3476 & ~n50516;
  assign n50518 = ~n50499 & ~n50517;
  assign n50519 = n3374 & ~n50518;
  assign n50520 = ~n34120 & ~n50519;
  assign n50521 = n3655 & ~n50520;
  assign n50522 = ~n25331 & ~n34544;
  assign n50523 = controllable_nhgrant0 & ~n50522;
  assign n50524 = ~n3945 & ~n50523;
  assign n50525 = ~n3281 & ~n50524;
  assign n50526 = ~n3281 & ~n50525;
  assign n50527 = n3378 & ~n50526;
  assign n50528 = ~n25338 & ~n34562;
  assign n50529 = controllable_nhgrant0 & ~n50528;
  assign n50530 = ~n3987 & ~n50529;
  assign n50531 = ~n3281 & ~n50530;
  assign n50532 = ~n3950 & ~n50531;
  assign n50533 = ~n3378 & ~n50532;
  assign n50534 = ~n50527 & ~n50533;
  assign n50535 = n3492 & ~n50534;
  assign n50536 = ~n3493 & ~n50535;
  assign n50537 = n3485 & ~n50536;
  assign n50538 = ~n3486 & ~n50537;
  assign n50539 = ~n3476 & ~n50538;
  assign n50540 = ~n25331 & ~n34590;
  assign n50541 = controllable_nhgrant0 & ~n50540;
  assign n50542 = ~n3945 & ~n50541;
  assign n50543 = ~n3281 & ~n50542;
  assign n50544 = ~n3281 & ~n50543;
  assign n50545 = n3378 & ~n50544;
  assign n50546 = ~n25338 & ~n34612;
  assign n50547 = controllable_nhgrant0 & ~n50546;
  assign n50548 = ~n3987 & ~n50547;
  assign n50549 = ~n3281 & ~n50548;
  assign n50550 = ~n4089 & ~n50549;
  assign n50551 = ~n3378 & ~n50550;
  assign n50552 = ~n50545 & ~n50551;
  assign n50553 = n3492 & ~n50552;
  assign n50554 = ~n34114 & ~n50553;
  assign n50555 = n3485 & ~n50554;
  assign n50556 = ~n34113 & ~n50555;
  assign n50557 = n3476 & ~n50556;
  assign n50558 = ~n50539 & ~n50557;
  assign n50559 = n3374 & ~n50558;
  assign n50560 = ~n34120 & ~n50559;
  assign n50561 = ~n3655 & ~n50560;
  assign n50562 = ~n50521 & ~n50561;
  assign n50563 = ~n3652 & ~n50562;
  assign n50564 = ~n50481 & ~n50563;
  assign n50565 = ~n3368 & ~n50564;
  assign n50566 = ~n25499 & ~n34657;
  assign n50567 = controllable_nhgrant0 & ~n50566;
  assign n50568 = ~n4646 & ~n50567;
  assign n50569 = ~n3281 & ~n50568;
  assign n50570 = ~n3281 & ~n50569;
  assign n50571 = n3492 & ~n50570;
  assign n50572 = n3492 & ~n50571;
  assign n50573 = n3485 & ~n50572;
  assign n50574 = n3485 & ~n50573;
  assign n50575 = ~n3476 & ~n50574;
  assign n50576 = ~n25499 & ~n34730;
  assign n50577 = controllable_nhgrant0 & ~n50576;
  assign n50578 = ~n4646 & ~n50577;
  assign n50579 = ~n3281 & ~n50578;
  assign n50580 = ~n3281 & ~n50579;
  assign n50581 = n3492 & ~n50580;
  assign n50582 = ~n34669 & ~n50581;
  assign n50583 = n3485 & ~n50582;
  assign n50584 = ~n34668 & ~n50583;
  assign n50585 = n3476 & ~n50584;
  assign n50586 = ~n50575 & ~n50585;
  assign n50587 = n3374 & ~n50586;
  assign n50588 = n3374 & ~n50587;
  assign n50589 = n3655 & ~n50588;
  assign n50590 = ~n25499 & ~n34767;
  assign n50591 = controllable_nhgrant0 & ~n50590;
  assign n50592 = ~n4646 & ~n50591;
  assign n50593 = ~n3281 & ~n50592;
  assign n50594 = ~n3281 & ~n50593;
  assign n50595 = n3492 & ~n50594;
  assign n50596 = n3492 & ~n50595;
  assign n50597 = n3485 & ~n50596;
  assign n50598 = n3485 & ~n50597;
  assign n50599 = ~n3476 & ~n50598;
  assign n50600 = ~n25499 & ~n34800;
  assign n50601 = controllable_nhgrant0 & ~n50600;
  assign n50602 = ~n4646 & ~n50601;
  assign n50603 = ~n3281 & ~n50602;
  assign n50604 = ~n3281 & ~n50603;
  assign n50605 = n3492 & ~n50604;
  assign n50606 = ~n34669 & ~n50605;
  assign n50607 = n3485 & ~n50606;
  assign n50608 = ~n34668 & ~n50607;
  assign n50609 = n3476 & ~n50608;
  assign n50610 = ~n50599 & ~n50609;
  assign n50611 = n3374 & ~n50610;
  assign n50612 = n3374 & ~n50611;
  assign n50613 = ~n3655 & ~n50612;
  assign n50614 = ~n50589 & ~n50613;
  assign n50615 = n3652 & ~n50614;
  assign n50616 = ~n25499 & ~n34832;
  assign n50617 = controllable_nhgrant0 & ~n50616;
  assign n50618 = ~n4646 & ~n50617;
  assign n50619 = ~n3281 & ~n50618;
  assign n50620 = ~n3281 & ~n50619;
  assign n50621 = n3492 & ~n50620;
  assign n50622 = n3492 & ~n50621;
  assign n50623 = n3485 & ~n50622;
  assign n50624 = n3485 & ~n50623;
  assign n50625 = ~n3476 & ~n50624;
  assign n50626 = ~n25499 & ~n34858;
  assign n50627 = controllable_nhgrant0 & ~n50626;
  assign n50628 = ~n4646 & ~n50627;
  assign n50629 = ~n3281 & ~n50628;
  assign n50630 = ~n3281 & ~n50629;
  assign n50631 = n3492 & ~n50630;
  assign n50632 = ~n34669 & ~n50631;
  assign n50633 = n3485 & ~n50632;
  assign n50634 = ~n34668 & ~n50633;
  assign n50635 = n3476 & ~n50634;
  assign n50636 = ~n50625 & ~n50635;
  assign n50637 = n3374 & ~n50636;
  assign n50638 = n3374 & ~n50637;
  assign n50639 = n3655 & ~n50638;
  assign n50640 = ~n25499 & ~n34888;
  assign n50641 = controllable_nhgrant0 & ~n50640;
  assign n50642 = ~n4646 & ~n50641;
  assign n50643 = ~n3281 & ~n50642;
  assign n50644 = ~n3281 & ~n50643;
  assign n50645 = n3492 & ~n50644;
  assign n50646 = n3492 & ~n50645;
  assign n50647 = n3485 & ~n50646;
  assign n50648 = n3485 & ~n50647;
  assign n50649 = ~n3476 & ~n50648;
  assign n50650 = ~n25499 & ~n34914;
  assign n50651 = controllable_nhgrant0 & ~n50650;
  assign n50652 = ~n4646 & ~n50651;
  assign n50653 = ~n3281 & ~n50652;
  assign n50654 = ~n3281 & ~n50653;
  assign n50655 = n3492 & ~n50654;
  assign n50656 = ~n34669 & ~n50655;
  assign n50657 = n3485 & ~n50656;
  assign n50658 = ~n34668 & ~n50657;
  assign n50659 = n3476 & ~n50658;
  assign n50660 = ~n50649 & ~n50659;
  assign n50661 = n3374 & ~n50660;
  assign n50662 = n3374 & ~n50661;
  assign n50663 = ~n3655 & ~n50662;
  assign n50664 = ~n50639 & ~n50663;
  assign n50665 = ~n3652 & ~n50664;
  assign n50666 = ~n50615 & ~n50665;
  assign n50667 = n3368 & ~n50666;
  assign n50668 = ~n50565 & ~n50667;
  assign n50669 = ~n3362 & ~n50668;
  assign n50670 = ~n3362 & ~n50669;
  assign n50671 = ~n3359 & ~n50670;
  assign n50672 = ~n3359 & ~n50671;
  assign n50673 = n3356 & ~n50672;
  assign n50674 = ~n25649 & ~n34965;
  assign n50675 = controllable_nhgrant0 & ~n50674;
  assign n50676 = ~n5245 & ~n50675;
  assign n50677 = ~n3281 & ~n50676;
  assign n50678 = ~n3783 & ~n50677;
  assign n50679 = ~n3378 & ~n50678;
  assign n50680 = ~n34939 & ~n50679;
  assign n50681 = n3492 & ~n50680;
  assign n50682 = ~n3631 & ~n50681;
  assign n50683 = n3485 & ~n50682;
  assign n50684 = ~n3630 & ~n50683;
  assign n50685 = ~n3476 & ~n50684;
  assign n50686 = ~n34979 & ~n50681;
  assign n50687 = n3485 & ~n50686;
  assign n50688 = ~n34978 & ~n50687;
  assign n50689 = n3476 & ~n50688;
  assign n50690 = ~n50685 & ~n50689;
  assign n50691 = ~n3374 & ~n50690;
  assign n50692 = ~n25663 & ~n35031;
  assign n50693 = controllable_nhgrant0 & ~n50692;
  assign n50694 = ~n5363 & ~n50693;
  assign n50695 = ~n3281 & ~n50694;
  assign n50696 = ~n3950 & ~n50695;
  assign n50697 = n3378 & ~n50696;
  assign n50698 = ~n25684 & ~n35097;
  assign n50699 = controllable_nhgrant0 & ~n50698;
  assign n50700 = ~n5534 & ~n50699;
  assign n50701 = ~n3281 & ~n50700;
  assign n50702 = ~n3950 & ~n50701;
  assign n50703 = ~n3378 & ~n50702;
  assign n50704 = ~n50697 & ~n50703;
  assign n50705 = n3492 & ~n50704;
  assign n50706 = ~n3631 & ~n50705;
  assign n50707 = n3485 & ~n50706;
  assign n50708 = ~n3630 & ~n50707;
  assign n50709 = ~n3476 & ~n50708;
  assign n50710 = ~n25698 & ~n35189;
  assign n50711 = controllable_nhgrant0 & ~n50710;
  assign n50712 = ~n5809 & ~n50711;
  assign n50713 = ~n3281 & ~n50712;
  assign n50714 = ~n4089 & ~n50713;
  assign n50715 = n3378 & ~n50714;
  assign n50716 = ~n25726 & ~n35266;
  assign n50717 = controllable_nhgrant0 & ~n50716;
  assign n50718 = ~n6082 & ~n50717;
  assign n50719 = ~n3281 & ~n50718;
  assign n50720 = ~n4089 & ~n50719;
  assign n50721 = ~n3378 & ~n50720;
  assign n50722 = ~n50715 & ~n50721;
  assign n50723 = n3492 & ~n50722;
  assign n50724 = ~n34979 & ~n50723;
  assign n50725 = n3485 & ~n50724;
  assign n50726 = ~n34978 & ~n50725;
  assign n50727 = n3476 & ~n50726;
  assign n50728 = ~n50709 & ~n50727;
  assign n50729 = n3374 & ~n50728;
  assign n50730 = ~n50691 & ~n50729;
  assign n50731 = n3655 & ~n50730;
  assign n50732 = ~n25649 & ~n35307;
  assign n50733 = controllable_nhgrant0 & ~n50732;
  assign n50734 = ~n5245 & ~n50733;
  assign n50735 = ~n3281 & ~n50734;
  assign n50736 = ~n3783 & ~n50735;
  assign n50737 = ~n3378 & ~n50736;
  assign n50738 = ~n34939 & ~n50737;
  assign n50739 = n3492 & ~n50738;
  assign n50740 = ~n3631 & ~n50739;
  assign n50741 = n3485 & ~n50740;
  assign n50742 = ~n3630 & ~n50741;
  assign n50743 = ~n3476 & ~n50742;
  assign n50744 = ~n34979 & ~n50739;
  assign n50745 = n3485 & ~n50744;
  assign n50746 = ~n34978 & ~n50745;
  assign n50747 = n3476 & ~n50746;
  assign n50748 = ~n50743 & ~n50747;
  assign n50749 = ~n3374 & ~n50748;
  assign n50750 = ~n25663 & ~n35327;
  assign n50751 = controllable_nhgrant0 & ~n50750;
  assign n50752 = ~n5363 & ~n50751;
  assign n50753 = ~n3281 & ~n50752;
  assign n50754 = ~n3950 & ~n50753;
  assign n50755 = n3378 & ~n50754;
  assign n50756 = ~n25684 & ~n35406;
  assign n50757 = controllable_nhgrant0 & ~n50756;
  assign n50758 = ~n5534 & ~n50757;
  assign n50759 = ~n3281 & ~n50758;
  assign n50760 = ~n3950 & ~n50759;
  assign n50761 = ~n3378 & ~n50760;
  assign n50762 = ~n50755 & ~n50761;
  assign n50763 = n3492 & ~n50762;
  assign n50764 = ~n3631 & ~n50763;
  assign n50765 = n3485 & ~n50764;
  assign n50766 = ~n3630 & ~n50765;
  assign n50767 = ~n3476 & ~n50766;
  assign n50768 = ~n25698 & ~n35441;
  assign n50769 = controllable_nhgrant0 & ~n50768;
  assign n50770 = ~n5809 & ~n50769;
  assign n50771 = ~n3281 & ~n50770;
  assign n50772 = ~n4089 & ~n50771;
  assign n50773 = n3378 & ~n50772;
  assign n50774 = ~n25726 & ~n35530;
  assign n50775 = controllable_nhgrant0 & ~n50774;
  assign n50776 = ~n6082 & ~n50775;
  assign n50777 = ~n3281 & ~n50776;
  assign n50778 = ~n4089 & ~n50777;
  assign n50779 = ~n3378 & ~n50778;
  assign n50780 = ~n50773 & ~n50779;
  assign n50781 = n3492 & ~n50780;
  assign n50782 = ~n34979 & ~n50781;
  assign n50783 = n3485 & ~n50782;
  assign n50784 = ~n34978 & ~n50783;
  assign n50785 = n3476 & ~n50784;
  assign n50786 = ~n50767 & ~n50785;
  assign n50787 = n3374 & ~n50786;
  assign n50788 = ~n50749 & ~n50787;
  assign n50789 = ~n3655 & ~n50788;
  assign n50790 = ~n50731 & ~n50789;
  assign n50791 = n3652 & ~n50790;
  assign n50792 = ~n25649 & ~n35566;
  assign n50793 = controllable_nhgrant0 & ~n50792;
  assign n50794 = ~n5245 & ~n50793;
  assign n50795 = ~n3281 & ~n50794;
  assign n50796 = ~n3783 & ~n50795;
  assign n50797 = ~n3378 & ~n50796;
  assign n50798 = ~n34939 & ~n50797;
  assign n50799 = n3492 & ~n50798;
  assign n50800 = ~n3631 & ~n50799;
  assign n50801 = n3485 & ~n50800;
  assign n50802 = ~n3630 & ~n50801;
  assign n50803 = ~n3476 & ~n50802;
  assign n50804 = ~n34979 & ~n50799;
  assign n50805 = n3485 & ~n50804;
  assign n50806 = ~n34978 & ~n50805;
  assign n50807 = n3476 & ~n50806;
  assign n50808 = ~n50803 & ~n50807;
  assign n50809 = ~n3374 & ~n50808;
  assign n50810 = ~n25663 & ~n35586;
  assign n50811 = controllable_nhgrant0 & ~n50810;
  assign n50812 = ~n5363 & ~n50811;
  assign n50813 = ~n3281 & ~n50812;
  assign n50814 = ~n3950 & ~n50813;
  assign n50815 = n3378 & ~n50814;
  assign n50816 = ~n25684 & ~n35639;
  assign n50817 = controllable_nhgrant0 & ~n50816;
  assign n50818 = ~n5534 & ~n50817;
  assign n50819 = ~n3281 & ~n50818;
  assign n50820 = ~n3950 & ~n50819;
  assign n50821 = ~n3378 & ~n50820;
  assign n50822 = ~n50815 & ~n50821;
  assign n50823 = n3492 & ~n50822;
  assign n50824 = ~n3631 & ~n50823;
  assign n50825 = n3485 & ~n50824;
  assign n50826 = ~n3630 & ~n50825;
  assign n50827 = ~n3476 & ~n50826;
  assign n50828 = ~n25698 & ~n35667;
  assign n50829 = controllable_nhgrant0 & ~n50828;
  assign n50830 = ~n5809 & ~n50829;
  assign n50831 = ~n3281 & ~n50830;
  assign n50832 = ~n4089 & ~n50831;
  assign n50833 = n3378 & ~n50832;
  assign n50834 = ~n25726 & ~n35724;
  assign n50835 = controllable_nhgrant0 & ~n50834;
  assign n50836 = ~n6082 & ~n50835;
  assign n50837 = ~n3281 & ~n50836;
  assign n50838 = ~n4089 & ~n50837;
  assign n50839 = ~n3378 & ~n50838;
  assign n50840 = ~n50833 & ~n50839;
  assign n50841 = n3492 & ~n50840;
  assign n50842 = ~n34979 & ~n50841;
  assign n50843 = n3485 & ~n50842;
  assign n50844 = ~n34978 & ~n50843;
  assign n50845 = n3476 & ~n50844;
  assign n50846 = ~n50827 & ~n50845;
  assign n50847 = n3374 & ~n50846;
  assign n50848 = ~n50809 & ~n50847;
  assign n50849 = n3655 & ~n50848;
  assign n50850 = ~n25649 & ~n35758;
  assign n50851 = controllable_nhgrant0 & ~n50850;
  assign n50852 = ~n5245 & ~n50851;
  assign n50853 = ~n3281 & ~n50852;
  assign n50854 = ~n3783 & ~n50853;
  assign n50855 = ~n3378 & ~n50854;
  assign n50856 = ~n34939 & ~n50855;
  assign n50857 = n3492 & ~n50856;
  assign n50858 = ~n3631 & ~n50857;
  assign n50859 = n3485 & ~n50858;
  assign n50860 = ~n3630 & ~n50859;
  assign n50861 = ~n3476 & ~n50860;
  assign n50862 = ~n34979 & ~n50857;
  assign n50863 = n3485 & ~n50862;
  assign n50864 = ~n34978 & ~n50863;
  assign n50865 = n3476 & ~n50864;
  assign n50866 = ~n50861 & ~n50865;
  assign n50867 = ~n3374 & ~n50866;
  assign n50868 = ~n25663 & ~n35778;
  assign n50869 = controllable_nhgrant0 & ~n50868;
  assign n50870 = ~n5363 & ~n50869;
  assign n50871 = ~n3281 & ~n50870;
  assign n50872 = ~n3950 & ~n50871;
  assign n50873 = n3378 & ~n50872;
  assign n50874 = ~n25684 & ~n35831;
  assign n50875 = controllable_nhgrant0 & ~n50874;
  assign n50876 = ~n5534 & ~n50875;
  assign n50877 = ~n3281 & ~n50876;
  assign n50878 = ~n3950 & ~n50877;
  assign n50879 = ~n3378 & ~n50878;
  assign n50880 = ~n50873 & ~n50879;
  assign n50881 = n3492 & ~n50880;
  assign n50882 = ~n3631 & ~n50881;
  assign n50883 = n3485 & ~n50882;
  assign n50884 = ~n3630 & ~n50883;
  assign n50885 = ~n3476 & ~n50884;
  assign n50886 = ~n25698 & ~n35859;
  assign n50887 = controllable_nhgrant0 & ~n50886;
  assign n50888 = ~n5809 & ~n50887;
  assign n50889 = ~n3281 & ~n50888;
  assign n50890 = ~n4089 & ~n50889;
  assign n50891 = n3378 & ~n50890;
  assign n50892 = ~n25726 & ~n35916;
  assign n50893 = controllable_nhgrant0 & ~n50892;
  assign n50894 = ~n6082 & ~n50893;
  assign n50895 = ~n3281 & ~n50894;
  assign n50896 = ~n4089 & ~n50895;
  assign n50897 = ~n3378 & ~n50896;
  assign n50898 = ~n50891 & ~n50897;
  assign n50899 = n3492 & ~n50898;
  assign n50900 = ~n34979 & ~n50899;
  assign n50901 = n3485 & ~n50900;
  assign n50902 = ~n34978 & ~n50901;
  assign n50903 = n3476 & ~n50902;
  assign n50904 = ~n50885 & ~n50903;
  assign n50905 = n3374 & ~n50904;
  assign n50906 = ~n50867 & ~n50905;
  assign n50907 = ~n3655 & ~n50906;
  assign n50908 = ~n50849 & ~n50907;
  assign n50909 = ~n3652 & ~n50908;
  assign n50910 = ~n50791 & ~n50909;
  assign n50911 = ~n3368 & ~n50910;
  assign n50912 = ~n25905 & ~n35995;
  assign n50913 = controllable_nhgrant0 & ~n50912;
  assign n50914 = ~n7118 & ~n50913;
  assign n50915 = ~n3281 & ~n50914;
  assign n50916 = ~n3281 & ~n50915;
  assign n50917 = ~n3378 & ~n50916;
  assign n50918 = ~n35969 & ~n50917;
  assign n50919 = n3492 & ~n50918;
  assign n50920 = n3492 & ~n50919;
  assign n50921 = n3485 & ~n50920;
  assign n50922 = n3485 & ~n50921;
  assign n50923 = ~n3374 & ~n50922;
  assign n50924 = ~n25919 & ~n36061;
  assign n50925 = controllable_nhgrant0 & ~n50924;
  assign n50926 = ~n7166 & ~n50925;
  assign n50927 = ~n3281 & ~n50926;
  assign n50928 = ~n3281 & ~n50927;
  assign n50929 = n3378 & ~n50928;
  assign n50930 = ~n25927 & ~n36127;
  assign n50931 = controllable_nhgrant0 & ~n50930;
  assign n50932 = ~n7208 & ~n50931;
  assign n50933 = ~n3281 & ~n50932;
  assign n50934 = ~n3281 & ~n50933;
  assign n50935 = ~n3378 & ~n50934;
  assign n50936 = ~n50929 & ~n50935;
  assign n50937 = n3492 & ~n50936;
  assign n50938 = n3492 & ~n50937;
  assign n50939 = n3485 & ~n50938;
  assign n50940 = n3485 & ~n50939;
  assign n50941 = ~n3476 & ~n50940;
  assign n50942 = ~n25941 & ~n36228;
  assign n50943 = controllable_nhgrant0 & ~n50942;
  assign n50944 = ~n7432 & ~n50943;
  assign n50945 = ~n3281 & ~n50944;
  assign n50946 = ~n3281 & ~n50945;
  assign n50947 = n3378 & ~n50946;
  assign n50948 = ~n25949 & ~n36329;
  assign n50949 = controllable_nhgrant0 & ~n50948;
  assign n50950 = ~n7668 & ~n50949;
  assign n50951 = ~n3281 & ~n50950;
  assign n50952 = ~n3281 & ~n50951;
  assign n50953 = ~n3378 & ~n50952;
  assign n50954 = ~n50947 & ~n50953;
  assign n50955 = n3492 & ~n50954;
  assign n50956 = ~n34669 & ~n50955;
  assign n50957 = n3485 & ~n50956;
  assign n50958 = ~n34668 & ~n50957;
  assign n50959 = n3476 & ~n50958;
  assign n50960 = ~n50941 & ~n50959;
  assign n50961 = n3374 & ~n50960;
  assign n50962 = ~n50923 & ~n50961;
  assign n50963 = n3655 & ~n50962;
  assign n50964 = ~n25905 & ~n36370;
  assign n50965 = controllable_nhgrant0 & ~n50964;
  assign n50966 = ~n7118 & ~n50965;
  assign n50967 = ~n3281 & ~n50966;
  assign n50968 = ~n3281 & ~n50967;
  assign n50969 = ~n3378 & ~n50968;
  assign n50970 = ~n35969 & ~n50969;
  assign n50971 = n3492 & ~n50970;
  assign n50972 = n3492 & ~n50971;
  assign n50973 = n3485 & ~n50972;
  assign n50974 = n3485 & ~n50973;
  assign n50975 = ~n3374 & ~n50974;
  assign n50976 = ~n25919 & ~n36394;
  assign n50977 = controllable_nhgrant0 & ~n50976;
  assign n50978 = ~n7166 & ~n50977;
  assign n50979 = ~n3281 & ~n50978;
  assign n50980 = ~n3281 & ~n50979;
  assign n50981 = n3378 & ~n50980;
  assign n50982 = ~n25927 & ~n36459;
  assign n50983 = controllable_nhgrant0 & ~n50982;
  assign n50984 = ~n7208 & ~n50983;
  assign n50985 = ~n3281 & ~n50984;
  assign n50986 = ~n3281 & ~n50985;
  assign n50987 = ~n3378 & ~n50986;
  assign n50988 = ~n50981 & ~n50987;
  assign n50989 = n3492 & ~n50988;
  assign n50990 = n3492 & ~n50989;
  assign n50991 = n3485 & ~n50990;
  assign n50992 = n3485 & ~n50991;
  assign n50993 = ~n3476 & ~n50992;
  assign n50994 = ~n25941 & ~n36494;
  assign n50995 = controllable_nhgrant0 & ~n50994;
  assign n50996 = ~n7432 & ~n50995;
  assign n50997 = ~n3281 & ~n50996;
  assign n50998 = ~n3281 & ~n50997;
  assign n50999 = n3378 & ~n50998;
  assign n51000 = ~n25949 & ~n36583;
  assign n51001 = controllable_nhgrant0 & ~n51000;
  assign n51002 = ~n7668 & ~n51001;
  assign n51003 = ~n3281 & ~n51002;
  assign n51004 = ~n3281 & ~n51003;
  assign n51005 = ~n3378 & ~n51004;
  assign n51006 = ~n50999 & ~n51005;
  assign n51007 = n3492 & ~n51006;
  assign n51008 = ~n34669 & ~n51007;
  assign n51009 = n3485 & ~n51008;
  assign n51010 = ~n34668 & ~n51009;
  assign n51011 = n3476 & ~n51010;
  assign n51012 = ~n50993 & ~n51011;
  assign n51013 = n3374 & ~n51012;
  assign n51014 = ~n50975 & ~n51013;
  assign n51015 = ~n3655 & ~n51014;
  assign n51016 = ~n50963 & ~n51015;
  assign n51017 = n3652 & ~n51016;
  assign n51018 = ~n25905 & ~n36619;
  assign n51019 = controllable_nhgrant0 & ~n51018;
  assign n51020 = ~n7118 & ~n51019;
  assign n51021 = ~n3281 & ~n51020;
  assign n51022 = ~n3281 & ~n51021;
  assign n51023 = ~n3378 & ~n51022;
  assign n51024 = ~n35969 & ~n51023;
  assign n51025 = n3492 & ~n51024;
  assign n51026 = n3492 & ~n51025;
  assign n51027 = n3485 & ~n51026;
  assign n51028 = n3485 & ~n51027;
  assign n51029 = ~n3374 & ~n51028;
  assign n51030 = ~n25919 & ~n36643;
  assign n51031 = controllable_nhgrant0 & ~n51030;
  assign n51032 = ~n7166 & ~n51031;
  assign n51033 = ~n3281 & ~n51032;
  assign n51034 = ~n3281 & ~n51033;
  assign n51035 = n3378 & ~n51034;
  assign n51036 = ~n25927 & ~n36690;
  assign n51037 = controllable_nhgrant0 & ~n51036;
  assign n51038 = ~n7208 & ~n51037;
  assign n51039 = ~n3281 & ~n51038;
  assign n51040 = ~n3281 & ~n51039;
  assign n51041 = ~n3378 & ~n51040;
  assign n51042 = ~n51035 & ~n51041;
  assign n51043 = n3492 & ~n51042;
  assign n51044 = n3492 & ~n51043;
  assign n51045 = n3485 & ~n51044;
  assign n51046 = n3485 & ~n51045;
  assign n51047 = ~n3476 & ~n51046;
  assign n51048 = ~n25941 & ~n36718;
  assign n51049 = controllable_nhgrant0 & ~n51048;
  assign n51050 = ~n7432 & ~n51049;
  assign n51051 = ~n3281 & ~n51050;
  assign n51052 = ~n3281 & ~n51051;
  assign n51053 = n3378 & ~n51052;
  assign n51054 = ~n25949 & ~n36775;
  assign n51055 = controllable_nhgrant0 & ~n51054;
  assign n51056 = ~n7668 & ~n51055;
  assign n51057 = ~n3281 & ~n51056;
  assign n51058 = ~n3281 & ~n51057;
  assign n51059 = ~n3378 & ~n51058;
  assign n51060 = ~n51053 & ~n51059;
  assign n51061 = n3492 & ~n51060;
  assign n51062 = ~n34669 & ~n51061;
  assign n51063 = n3485 & ~n51062;
  assign n51064 = ~n34668 & ~n51063;
  assign n51065 = n3476 & ~n51064;
  assign n51066 = ~n51047 & ~n51065;
  assign n51067 = n3374 & ~n51066;
  assign n51068 = ~n51029 & ~n51067;
  assign n51069 = n3655 & ~n51068;
  assign n51070 = ~n25905 & ~n36809;
  assign n51071 = controllable_nhgrant0 & ~n51070;
  assign n51072 = ~n7118 & ~n51071;
  assign n51073 = ~n3281 & ~n51072;
  assign n51074 = ~n3281 & ~n51073;
  assign n51075 = ~n3378 & ~n51074;
  assign n51076 = ~n35969 & ~n51075;
  assign n51077 = n3492 & ~n51076;
  assign n51078 = n3492 & ~n51077;
  assign n51079 = n3485 & ~n51078;
  assign n51080 = n3485 & ~n51079;
  assign n51081 = ~n3374 & ~n51080;
  assign n51082 = ~n25919 & ~n36833;
  assign n51083 = controllable_nhgrant0 & ~n51082;
  assign n51084 = ~n7166 & ~n51083;
  assign n51085 = ~n3281 & ~n51084;
  assign n51086 = ~n3281 & ~n51085;
  assign n51087 = n3378 & ~n51086;
  assign n51088 = ~n25927 & ~n36880;
  assign n51089 = controllable_nhgrant0 & ~n51088;
  assign n51090 = ~n7208 & ~n51089;
  assign n51091 = ~n3281 & ~n51090;
  assign n51092 = ~n3281 & ~n51091;
  assign n51093 = ~n3378 & ~n51092;
  assign n51094 = ~n51087 & ~n51093;
  assign n51095 = n3492 & ~n51094;
  assign n51096 = n3492 & ~n51095;
  assign n51097 = n3485 & ~n51096;
  assign n51098 = n3485 & ~n51097;
  assign n51099 = ~n3476 & ~n51098;
  assign n51100 = ~n25941 & ~n36908;
  assign n51101 = controllable_nhgrant0 & ~n51100;
  assign n51102 = ~n7432 & ~n51101;
  assign n51103 = ~n3281 & ~n51102;
  assign n51104 = ~n3281 & ~n51103;
  assign n51105 = n3378 & ~n51104;
  assign n51106 = ~n25949 & ~n36965;
  assign n51107 = controllable_nhgrant0 & ~n51106;
  assign n51108 = ~n7668 & ~n51107;
  assign n51109 = ~n3281 & ~n51108;
  assign n51110 = ~n3281 & ~n51109;
  assign n51111 = ~n3378 & ~n51110;
  assign n51112 = ~n51105 & ~n51111;
  assign n51113 = n3492 & ~n51112;
  assign n51114 = ~n34669 & ~n51113;
  assign n51115 = n3485 & ~n51114;
  assign n51116 = ~n34668 & ~n51115;
  assign n51117 = n3476 & ~n51116;
  assign n51118 = ~n51099 & ~n51117;
  assign n51119 = n3374 & ~n51118;
  assign n51120 = ~n51081 & ~n51119;
  assign n51121 = ~n3655 & ~n51120;
  assign n51122 = ~n51069 & ~n51121;
  assign n51123 = ~n3652 & ~n51122;
  assign n51124 = ~n51017 & ~n51123;
  assign n51125 = n3368 & ~n51124;
  assign n51126 = ~n50911 & ~n51125;
  assign n51127 = n3362 & ~n51126;
  assign n51128 = n3492 & ~n50678;
  assign n51129 = ~n3631 & ~n51128;
  assign n51130 = n3485 & ~n51129;
  assign n51131 = ~n3630 & ~n51130;
  assign n51132 = ~n3476 & ~n51131;
  assign n51133 = ~n3793 & ~n26156;
  assign n51134 = controllable_hgrant3 & ~n51133;
  assign n51135 = ~n26172 & ~n34103;
  assign n51136 = ~controllable_hgrant3 & ~n51135;
  assign n51137 = ~n51134 & ~n51136;
  assign n51138 = controllable_nhgrant0 & ~n51137;
  assign n51139 = ~n3793 & ~n26172;
  assign n51140 = controllable_hgrant3 & ~n51139;
  assign n51141 = ~n3793 & ~n26192;
  assign n51142 = ~controllable_hgrant3 & ~n51141;
  assign n51143 = ~n51140 & ~n51142;
  assign n51144 = ~controllable_nhgrant0 & ~n51143;
  assign n51145 = ~n51138 & ~n51144;
  assign n51146 = ~n3281 & ~n51145;
  assign n51147 = ~n3783 & ~n51146;
  assign n51148 = ~n3492 & ~n51147;
  assign n51149 = ~n37007 & ~n51148;
  assign n51150 = ~n3485 & ~n51149;
  assign n51151 = ~n34979 & ~n51128;
  assign n51152 = n3485 & ~n51151;
  assign n51153 = ~n51150 & ~n51152;
  assign n51154 = n3476 & ~n51153;
  assign n51155 = ~n51132 & ~n51154;
  assign n51156 = ~n3374 & ~n51155;
  assign n51157 = n3492 & ~n50702;
  assign n51158 = ~n3631 & ~n51157;
  assign n51159 = n3485 & ~n51158;
  assign n51160 = ~n3630 & ~n51159;
  assign n51161 = ~n3476 & ~n51160;
  assign n51162 = n3492 & ~n50720;
  assign n51163 = ~n34979 & ~n51162;
  assign n51164 = n3485 & ~n51163;
  assign n51165 = ~n51150 & ~n51164;
  assign n51166 = n3476 & ~n51165;
  assign n51167 = ~n51161 & ~n51166;
  assign n51168 = n3374 & ~n51167;
  assign n51169 = ~n51156 & ~n51168;
  assign n51170 = n3655 & ~n51169;
  assign n51171 = n3492 & ~n50736;
  assign n51172 = ~n3631 & ~n51171;
  assign n51173 = n3485 & ~n51172;
  assign n51174 = ~n3630 & ~n51173;
  assign n51175 = ~n3476 & ~n51174;
  assign n51176 = ~n3793 & ~n26239;
  assign n51177 = controllable_hgrant3 & ~n51176;
  assign n51178 = ~n26255 & ~n34103;
  assign n51179 = ~controllable_hgrant3 & ~n51178;
  assign n51180 = ~n51177 & ~n51179;
  assign n51181 = controllable_nhgrant0 & ~n51180;
  assign n51182 = ~n3793 & ~n26273;
  assign n51183 = controllable_hgrant3 & ~n51182;
  assign n51184 = ~n3793 & ~n26289;
  assign n51185 = ~controllable_hgrant3 & ~n51184;
  assign n51186 = ~n51183 & ~n51185;
  assign n51187 = ~controllable_nhgrant0 & ~n51186;
  assign n51188 = ~n51181 & ~n51187;
  assign n51189 = ~n3281 & ~n51188;
  assign n51190 = ~n3783 & ~n51189;
  assign n51191 = ~n3492 & ~n51190;
  assign n51192 = ~n37007 & ~n51191;
  assign n51193 = ~n3485 & ~n51192;
  assign n51194 = ~n34979 & ~n51171;
  assign n51195 = n3485 & ~n51194;
  assign n51196 = ~n51193 & ~n51195;
  assign n51197 = n3476 & ~n51196;
  assign n51198 = ~n51175 & ~n51197;
  assign n51199 = ~n3374 & ~n51198;
  assign n51200 = n3492 & ~n50760;
  assign n51201 = ~n3631 & ~n51200;
  assign n51202 = n3485 & ~n51201;
  assign n51203 = ~n3630 & ~n51202;
  assign n51204 = ~n3476 & ~n51203;
  assign n51205 = n3492 & ~n50778;
  assign n51206 = ~n34979 & ~n51205;
  assign n51207 = n3485 & ~n51206;
  assign n51208 = ~n51193 & ~n51207;
  assign n51209 = n3476 & ~n51208;
  assign n51210 = ~n51204 & ~n51209;
  assign n51211 = n3374 & ~n51210;
  assign n51212 = ~n51199 & ~n51211;
  assign n51213 = ~n3655 & ~n51212;
  assign n51214 = ~n51170 & ~n51213;
  assign n51215 = n3652 & ~n51214;
  assign n51216 = n3492 & ~n50796;
  assign n51217 = ~n3631 & ~n51216;
  assign n51218 = n3485 & ~n51217;
  assign n51219 = ~n3630 & ~n51218;
  assign n51220 = ~n3476 & ~n51219;
  assign n51221 = ~n3793 & ~n26338;
  assign n51222 = controllable_hgrant3 & ~n51221;
  assign n51223 = ~n26354 & ~n34103;
  assign n51224 = ~controllable_hgrant3 & ~n51223;
  assign n51225 = ~n51222 & ~n51224;
  assign n51226 = controllable_nhgrant0 & ~n51225;
  assign n51227 = ~n3793 & ~n26372;
  assign n51228 = controllable_hgrant3 & ~n51227;
  assign n51229 = ~n3793 & ~n26388;
  assign n51230 = ~controllable_hgrant3 & ~n51229;
  assign n51231 = ~n51228 & ~n51230;
  assign n51232 = ~controllable_nhgrant0 & ~n51231;
  assign n51233 = ~n51226 & ~n51232;
  assign n51234 = ~n3281 & ~n51233;
  assign n51235 = ~n3783 & ~n51234;
  assign n51236 = ~n3492 & ~n51235;
  assign n51237 = ~n37007 & ~n51236;
  assign n51238 = ~n3485 & ~n51237;
  assign n51239 = ~n34979 & ~n51216;
  assign n51240 = n3485 & ~n51239;
  assign n51241 = ~n51238 & ~n51240;
  assign n51242 = n3476 & ~n51241;
  assign n51243 = ~n51220 & ~n51242;
  assign n51244 = ~n3374 & ~n51243;
  assign n51245 = n3492 & ~n50820;
  assign n51246 = ~n3631 & ~n51245;
  assign n51247 = n3485 & ~n51246;
  assign n51248 = ~n3630 & ~n51247;
  assign n51249 = ~n3476 & ~n51248;
  assign n51250 = n3492 & ~n50838;
  assign n51251 = ~n34979 & ~n51250;
  assign n51252 = n3485 & ~n51251;
  assign n51253 = ~n51238 & ~n51252;
  assign n51254 = n3476 & ~n51253;
  assign n51255 = ~n51249 & ~n51254;
  assign n51256 = n3374 & ~n51255;
  assign n51257 = ~n51244 & ~n51256;
  assign n51258 = n3655 & ~n51257;
  assign n51259 = n3492 & ~n50854;
  assign n51260 = ~n3631 & ~n51259;
  assign n51261 = n3485 & ~n51260;
  assign n51262 = ~n3630 & ~n51261;
  assign n51263 = ~n3476 & ~n51262;
  assign n51264 = ~n3793 & ~n25647;
  assign n51265 = controllable_hgrant3 & ~n51264;
  assign n51266 = ~n6887 & ~n34103;
  assign n51267 = ~controllable_hgrant3 & ~n51266;
  assign n51268 = ~n51265 & ~n51267;
  assign n51269 = controllable_nhgrant0 & ~n51268;
  assign n51270 = ~n3793 & ~n5187;
  assign n51271 = controllable_hgrant3 & ~n51270;
  assign n51272 = ~n3793 & ~n5241;
  assign n51273 = ~controllable_hgrant3 & ~n51272;
  assign n51274 = ~n51271 & ~n51273;
  assign n51275 = ~controllable_nhgrant0 & ~n51274;
  assign n51276 = ~n51269 & ~n51275;
  assign n51277 = ~n3281 & ~n51276;
  assign n51278 = ~n3783 & ~n51277;
  assign n51279 = ~n3492 & ~n51278;
  assign n51280 = ~n37007 & ~n51279;
  assign n51281 = ~n3485 & ~n51280;
  assign n51282 = ~n34979 & ~n51259;
  assign n51283 = n3485 & ~n51282;
  assign n51284 = ~n51281 & ~n51283;
  assign n51285 = n3476 & ~n51284;
  assign n51286 = ~n51263 & ~n51285;
  assign n51287 = ~n3374 & ~n51286;
  assign n51288 = n3492 & ~n50878;
  assign n51289 = ~n3631 & ~n51288;
  assign n51290 = n3485 & ~n51289;
  assign n51291 = ~n3630 & ~n51290;
  assign n51292 = ~n3476 & ~n51291;
  assign n51293 = n3492 & ~n50896;
  assign n51294 = ~n34979 & ~n51293;
  assign n51295 = n3485 & ~n51294;
  assign n51296 = ~n51281 & ~n51295;
  assign n51297 = n3476 & ~n51296;
  assign n51298 = ~n51292 & ~n51297;
  assign n51299 = n3374 & ~n51298;
  assign n51300 = ~n51287 & ~n51299;
  assign n51301 = ~n3655 & ~n51300;
  assign n51302 = ~n51258 & ~n51301;
  assign n51303 = ~n3652 & ~n51302;
  assign n51304 = ~n51215 & ~n51303;
  assign n51305 = ~n3368 & ~n51304;
  assign n51306 = n3492 & ~n50916;
  assign n51307 = n3492 & ~n51306;
  assign n51308 = n3485 & ~n51307;
  assign n51309 = n3485 & ~n51308;
  assign n51310 = ~n3476 & ~n51309;
  assign n51311 = ~n8525 & ~n51308;
  assign n51312 = n3476 & ~n51311;
  assign n51313 = ~n51310 & ~n51312;
  assign n51314 = ~n3374 & ~n51313;
  assign n51315 = n3492 & ~n50934;
  assign n51316 = n3492 & ~n51315;
  assign n51317 = n3485 & ~n51316;
  assign n51318 = n3485 & ~n51317;
  assign n51319 = ~n3476 & ~n51318;
  assign n51320 = ~n3281 & ~n51146;
  assign n51321 = ~n3492 & ~n51320;
  assign n51322 = ~n37175 & ~n51321;
  assign n51323 = ~n3485 & ~n51322;
  assign n51324 = n3492 & ~n50952;
  assign n51325 = ~n34669 & ~n51324;
  assign n51326 = n3485 & ~n51325;
  assign n51327 = ~n51323 & ~n51326;
  assign n51328 = n3476 & ~n51327;
  assign n51329 = ~n51319 & ~n51328;
  assign n51330 = n3374 & ~n51329;
  assign n51331 = ~n51314 & ~n51330;
  assign n51332 = n3655 & ~n51331;
  assign n51333 = n3492 & ~n50968;
  assign n51334 = n3492 & ~n51333;
  assign n51335 = n3485 & ~n51334;
  assign n51336 = n3485 & ~n51335;
  assign n51337 = ~n3476 & ~n51336;
  assign n51338 = ~n8525 & ~n51335;
  assign n51339 = n3476 & ~n51338;
  assign n51340 = ~n51337 & ~n51339;
  assign n51341 = ~n3374 & ~n51340;
  assign n51342 = n3492 & ~n50986;
  assign n51343 = n3492 & ~n51342;
  assign n51344 = n3485 & ~n51343;
  assign n51345 = n3485 & ~n51344;
  assign n51346 = ~n3476 & ~n51345;
  assign n51347 = ~n3281 & ~n51189;
  assign n51348 = ~n3492 & ~n51347;
  assign n51349 = ~n37175 & ~n51348;
  assign n51350 = ~n3485 & ~n51349;
  assign n51351 = n3492 & ~n51004;
  assign n51352 = ~n34669 & ~n51351;
  assign n51353 = n3485 & ~n51352;
  assign n51354 = ~n51350 & ~n51353;
  assign n51355 = n3476 & ~n51354;
  assign n51356 = ~n51346 & ~n51355;
  assign n51357 = n3374 & ~n51356;
  assign n51358 = ~n51341 & ~n51357;
  assign n51359 = ~n3655 & ~n51358;
  assign n51360 = ~n51332 & ~n51359;
  assign n51361 = n3652 & ~n51360;
  assign n51362 = n3492 & ~n51022;
  assign n51363 = n3492 & ~n51362;
  assign n51364 = n3485 & ~n51363;
  assign n51365 = n3485 & ~n51364;
  assign n51366 = ~n3476 & ~n51365;
  assign n51367 = ~n8525 & ~n51364;
  assign n51368 = n3476 & ~n51367;
  assign n51369 = ~n51366 & ~n51368;
  assign n51370 = ~n3374 & ~n51369;
  assign n51371 = n3492 & ~n51040;
  assign n51372 = n3492 & ~n51371;
  assign n51373 = n3485 & ~n51372;
  assign n51374 = n3485 & ~n51373;
  assign n51375 = ~n3476 & ~n51374;
  assign n51376 = ~n3281 & ~n51234;
  assign n51377 = ~n3492 & ~n51376;
  assign n51378 = ~n37175 & ~n51377;
  assign n51379 = ~n3485 & ~n51378;
  assign n51380 = n3492 & ~n51058;
  assign n51381 = ~n34669 & ~n51380;
  assign n51382 = n3485 & ~n51381;
  assign n51383 = ~n51379 & ~n51382;
  assign n51384 = n3476 & ~n51383;
  assign n51385 = ~n51375 & ~n51384;
  assign n51386 = n3374 & ~n51385;
  assign n51387 = ~n51370 & ~n51386;
  assign n51388 = n3655 & ~n51387;
  assign n51389 = n3492 & ~n51074;
  assign n51390 = n3492 & ~n51389;
  assign n51391 = n3485 & ~n51390;
  assign n51392 = n3485 & ~n51391;
  assign n51393 = ~n3476 & ~n51392;
  assign n51394 = ~n8525 & ~n51391;
  assign n51395 = n3476 & ~n51394;
  assign n51396 = ~n51393 & ~n51395;
  assign n51397 = ~n3374 & ~n51396;
  assign n51398 = n3492 & ~n51092;
  assign n51399 = n3492 & ~n51398;
  assign n51400 = n3485 & ~n51399;
  assign n51401 = n3485 & ~n51400;
  assign n51402 = ~n3476 & ~n51401;
  assign n51403 = ~n3281 & ~n51277;
  assign n51404 = ~n3492 & ~n51403;
  assign n51405 = ~n37175 & ~n51404;
  assign n51406 = ~n3485 & ~n51405;
  assign n51407 = n3492 & ~n51110;
  assign n51408 = ~n34669 & ~n51407;
  assign n51409 = n3485 & ~n51408;
  assign n51410 = ~n51406 & ~n51409;
  assign n51411 = n3476 & ~n51410;
  assign n51412 = ~n51402 & ~n51411;
  assign n51413 = n3374 & ~n51412;
  assign n51414 = ~n51397 & ~n51413;
  assign n51415 = ~n3655 & ~n51414;
  assign n51416 = ~n51388 & ~n51415;
  assign n51417 = ~n3652 & ~n51416;
  assign n51418 = ~n51361 & ~n51417;
  assign n51419 = n3368 & ~n51418;
  assign n51420 = ~n51305 & ~n51419;
  assign n51421 = ~n3362 & ~n51420;
  assign n51422 = ~n51127 & ~n51421;
  assign n51423 = n3359 & ~n51422;
  assign n51424 = ~n3485 & ~n51147;
  assign n51425 = ~n51152 & ~n51424;
  assign n51426 = n3476 & ~n51425;
  assign n51427 = ~n51132 & ~n51426;
  assign n51428 = ~n3374 & ~n51427;
  assign n51429 = ~n51164 & ~n51424;
  assign n51430 = n3476 & ~n51429;
  assign n51431 = ~n51161 & ~n51430;
  assign n51432 = n3374 & ~n51431;
  assign n51433 = ~n51428 & ~n51432;
  assign n51434 = n3655 & ~n51433;
  assign n51435 = ~n3485 & ~n51190;
  assign n51436 = ~n51195 & ~n51435;
  assign n51437 = n3476 & ~n51436;
  assign n51438 = ~n51175 & ~n51437;
  assign n51439 = ~n3374 & ~n51438;
  assign n51440 = ~n51207 & ~n51435;
  assign n51441 = n3476 & ~n51440;
  assign n51442 = ~n51204 & ~n51441;
  assign n51443 = n3374 & ~n51442;
  assign n51444 = ~n51439 & ~n51443;
  assign n51445 = ~n3655 & ~n51444;
  assign n51446 = ~n51434 & ~n51445;
  assign n51447 = n3652 & ~n51446;
  assign n51448 = ~n3485 & ~n51235;
  assign n51449 = ~n51240 & ~n51448;
  assign n51450 = n3476 & ~n51449;
  assign n51451 = ~n51220 & ~n51450;
  assign n51452 = ~n3374 & ~n51451;
  assign n51453 = ~n51252 & ~n51448;
  assign n51454 = n3476 & ~n51453;
  assign n51455 = ~n51249 & ~n51454;
  assign n51456 = n3374 & ~n51455;
  assign n51457 = ~n51452 & ~n51456;
  assign n51458 = n3655 & ~n51457;
  assign n51459 = ~n3485 & ~n51278;
  assign n51460 = ~n51283 & ~n51459;
  assign n51461 = n3476 & ~n51460;
  assign n51462 = ~n51263 & ~n51461;
  assign n51463 = ~n3374 & ~n51462;
  assign n51464 = ~n51295 & ~n51459;
  assign n51465 = n3476 & ~n51464;
  assign n51466 = ~n51292 & ~n51465;
  assign n51467 = n3374 & ~n51466;
  assign n51468 = ~n51463 & ~n51467;
  assign n51469 = ~n3655 & ~n51468;
  assign n51470 = ~n51458 & ~n51469;
  assign n51471 = ~n3652 & ~n51470;
  assign n51472 = ~n51447 & ~n51471;
  assign n51473 = ~n3368 & ~n51472;
  assign n51474 = ~n8689 & ~n51308;
  assign n51475 = n3476 & ~n51474;
  assign n51476 = ~n51310 & ~n51475;
  assign n51477 = ~n3374 & ~n51476;
  assign n51478 = ~n3485 & ~n51320;
  assign n51479 = ~n51326 & ~n51478;
  assign n51480 = n3476 & ~n51479;
  assign n51481 = ~n51319 & ~n51480;
  assign n51482 = n3374 & ~n51481;
  assign n51483 = ~n51477 & ~n51482;
  assign n51484 = n3655 & ~n51483;
  assign n51485 = ~n8689 & ~n51335;
  assign n51486 = n3476 & ~n51485;
  assign n51487 = ~n51337 & ~n51486;
  assign n51488 = ~n3374 & ~n51487;
  assign n51489 = ~n3485 & ~n51347;
  assign n51490 = ~n51353 & ~n51489;
  assign n51491 = n3476 & ~n51490;
  assign n51492 = ~n51346 & ~n51491;
  assign n51493 = n3374 & ~n51492;
  assign n51494 = ~n51488 & ~n51493;
  assign n51495 = ~n3655 & ~n51494;
  assign n51496 = ~n51484 & ~n51495;
  assign n51497 = n3652 & ~n51496;
  assign n51498 = ~n8689 & ~n51364;
  assign n51499 = n3476 & ~n51498;
  assign n51500 = ~n51366 & ~n51499;
  assign n51501 = ~n3374 & ~n51500;
  assign n51502 = ~n3485 & ~n51376;
  assign n51503 = ~n51382 & ~n51502;
  assign n51504 = n3476 & ~n51503;
  assign n51505 = ~n51375 & ~n51504;
  assign n51506 = n3374 & ~n51505;
  assign n51507 = ~n51501 & ~n51506;
  assign n51508 = n3655 & ~n51507;
  assign n51509 = ~n8689 & ~n51391;
  assign n51510 = n3476 & ~n51509;
  assign n51511 = ~n51393 & ~n51510;
  assign n51512 = ~n3374 & ~n51511;
  assign n51513 = ~n3485 & ~n51403;
  assign n51514 = ~n51409 & ~n51513;
  assign n51515 = n3476 & ~n51514;
  assign n51516 = ~n51402 & ~n51515;
  assign n51517 = n3374 & ~n51516;
  assign n51518 = ~n51512 & ~n51517;
  assign n51519 = ~n3655 & ~n51518;
  assign n51520 = ~n51508 & ~n51519;
  assign n51521 = ~n3652 & ~n51520;
  assign n51522 = ~n51497 & ~n51521;
  assign n51523 = n3368 & ~n51522;
  assign n51524 = ~n51473 & ~n51523;
  assign n51525 = n3362 & ~n51524;
  assign n51526 = n3378 & ~n50678;
  assign n51527 = ~n26684 & ~n37392;
  assign n51528 = controllable_nhgrant0 & ~n51527;
  assign n51529 = ~n8785 & ~n51528;
  assign n51530 = ~n3281 & ~n51529;
  assign n51531 = ~n3783 & ~n51530;
  assign n51532 = ~n3378 & ~n51531;
  assign n51533 = ~n51526 & ~n51532;
  assign n51534 = n3492 & ~n51533;
  assign n51535 = ~n3631 & ~n51534;
  assign n51536 = n3485 & ~n51535;
  assign n51537 = ~n3630 & ~n51536;
  assign n51538 = ~n3476 & ~n51537;
  assign n51539 = ~n51148 & ~n51534;
  assign n51540 = n3485 & ~n51539;
  assign n51541 = ~n51424 & ~n51540;
  assign n51542 = n3476 & ~n51541;
  assign n51543 = ~n51538 & ~n51542;
  assign n51544 = ~n3374 & ~n51543;
  assign n51545 = n3378 & ~n50702;
  assign n51546 = ~n26705 & ~n37466;
  assign n51547 = controllable_nhgrant0 & ~n51546;
  assign n51548 = ~n8902 & ~n51547;
  assign n51549 = ~n3281 & ~n51548;
  assign n51550 = ~n3950 & ~n51549;
  assign n51551 = ~n3378 & ~n51550;
  assign n51552 = ~n51545 & ~n51551;
  assign n51553 = n3492 & ~n51552;
  assign n51554 = ~n3631 & ~n51553;
  assign n51555 = n3485 & ~n51554;
  assign n51556 = ~n3630 & ~n51555;
  assign n51557 = ~n3476 & ~n51556;
  assign n51558 = n3378 & ~n50720;
  assign n51559 = ~n26720 & ~n37548;
  assign n51560 = controllable_nhgrant0 & ~n51559;
  assign n51561 = ~n9096 & ~n51560;
  assign n51562 = ~n3281 & ~n51561;
  assign n51563 = ~n4089 & ~n51562;
  assign n51564 = ~n3378 & ~n51563;
  assign n51565 = ~n51558 & ~n51564;
  assign n51566 = n3492 & ~n51565;
  assign n51567 = ~n51148 & ~n51566;
  assign n51568 = n3485 & ~n51567;
  assign n51569 = ~n51424 & ~n51568;
  assign n51570 = n3476 & ~n51569;
  assign n51571 = ~n51557 & ~n51570;
  assign n51572 = n3374 & ~n51571;
  assign n51573 = ~n51544 & ~n51572;
  assign n51574 = n3655 & ~n51573;
  assign n51575 = n3378 & ~n50736;
  assign n51576 = ~n26684 & ~n37582;
  assign n51577 = controllable_nhgrant0 & ~n51576;
  assign n51578 = ~n8785 & ~n51577;
  assign n51579 = ~n3281 & ~n51578;
  assign n51580 = ~n3783 & ~n51579;
  assign n51581 = ~n3378 & ~n51580;
  assign n51582 = ~n51575 & ~n51581;
  assign n51583 = n3492 & ~n51582;
  assign n51584 = ~n3631 & ~n51583;
  assign n51585 = n3485 & ~n51584;
  assign n51586 = ~n3630 & ~n51585;
  assign n51587 = ~n3476 & ~n51586;
  assign n51588 = ~n51191 & ~n51583;
  assign n51589 = n3485 & ~n51588;
  assign n51590 = ~n51435 & ~n51589;
  assign n51591 = n3476 & ~n51590;
  assign n51592 = ~n51587 & ~n51591;
  assign n51593 = ~n3374 & ~n51592;
  assign n51594 = n3378 & ~n50760;
  assign n51595 = ~n26705 & ~n37660;
  assign n51596 = controllable_nhgrant0 & ~n51595;
  assign n51597 = ~n8902 & ~n51596;
  assign n51598 = ~n3281 & ~n51597;
  assign n51599 = ~n3950 & ~n51598;
  assign n51600 = ~n3378 & ~n51599;
  assign n51601 = ~n51594 & ~n51600;
  assign n51602 = n3492 & ~n51601;
  assign n51603 = ~n3631 & ~n51602;
  assign n51604 = n3485 & ~n51603;
  assign n51605 = ~n3630 & ~n51604;
  assign n51606 = ~n3476 & ~n51605;
  assign n51607 = n3378 & ~n50778;
  assign n51608 = ~n26720 & ~n37751;
  assign n51609 = controllable_nhgrant0 & ~n51608;
  assign n51610 = ~n9096 & ~n51609;
  assign n51611 = ~n3281 & ~n51610;
  assign n51612 = ~n4089 & ~n51611;
  assign n51613 = ~n3378 & ~n51612;
  assign n51614 = ~n51607 & ~n51613;
  assign n51615 = n3492 & ~n51614;
  assign n51616 = ~n51191 & ~n51615;
  assign n51617 = n3485 & ~n51616;
  assign n51618 = ~n51435 & ~n51617;
  assign n51619 = n3476 & ~n51618;
  assign n51620 = ~n51606 & ~n51619;
  assign n51621 = n3374 & ~n51620;
  assign n51622 = ~n51593 & ~n51621;
  assign n51623 = ~n3655 & ~n51622;
  assign n51624 = ~n51574 & ~n51623;
  assign n51625 = n3652 & ~n51624;
  assign n51626 = n3378 & ~n50796;
  assign n51627 = ~n26684 & ~n37785;
  assign n51628 = controllable_nhgrant0 & ~n51627;
  assign n51629 = ~n8785 & ~n51628;
  assign n51630 = ~n3281 & ~n51629;
  assign n51631 = ~n3783 & ~n51630;
  assign n51632 = ~n3378 & ~n51631;
  assign n51633 = ~n51626 & ~n51632;
  assign n51634 = n3492 & ~n51633;
  assign n51635 = ~n3631 & ~n51634;
  assign n51636 = n3485 & ~n51635;
  assign n51637 = ~n3630 & ~n51636;
  assign n51638 = ~n3476 & ~n51637;
  assign n51639 = ~n51236 & ~n51634;
  assign n51640 = n3485 & ~n51639;
  assign n51641 = ~n51448 & ~n51640;
  assign n51642 = n3476 & ~n51641;
  assign n51643 = ~n51638 & ~n51642;
  assign n51644 = ~n3374 & ~n51643;
  assign n51645 = n3378 & ~n50820;
  assign n51646 = ~n26705 & ~n37845;
  assign n51647 = controllable_nhgrant0 & ~n51646;
  assign n51648 = ~n8902 & ~n51647;
  assign n51649 = ~n3281 & ~n51648;
  assign n51650 = ~n3950 & ~n51649;
  assign n51651 = ~n3378 & ~n51650;
  assign n51652 = ~n51645 & ~n51651;
  assign n51653 = n3492 & ~n51652;
  assign n51654 = ~n3631 & ~n51653;
  assign n51655 = n3485 & ~n51654;
  assign n51656 = ~n3630 & ~n51655;
  assign n51657 = ~n3476 & ~n51656;
  assign n51658 = n3378 & ~n50838;
  assign n51659 = ~n26720 & ~n37907;
  assign n51660 = controllable_nhgrant0 & ~n51659;
  assign n51661 = ~n9096 & ~n51660;
  assign n51662 = ~n3281 & ~n51661;
  assign n51663 = ~n4089 & ~n51662;
  assign n51664 = ~n3378 & ~n51663;
  assign n51665 = ~n51658 & ~n51664;
  assign n51666 = n3492 & ~n51665;
  assign n51667 = ~n51236 & ~n51666;
  assign n51668 = n3485 & ~n51667;
  assign n51669 = ~n51448 & ~n51668;
  assign n51670 = n3476 & ~n51669;
  assign n51671 = ~n51657 & ~n51670;
  assign n51672 = n3374 & ~n51671;
  assign n51673 = ~n51644 & ~n51672;
  assign n51674 = n3655 & ~n51673;
  assign n51675 = n3378 & ~n50854;
  assign n51676 = ~n26684 & ~n37939;
  assign n51677 = controllable_nhgrant0 & ~n51676;
  assign n51678 = ~n8785 & ~n51677;
  assign n51679 = ~n3281 & ~n51678;
  assign n51680 = ~n3783 & ~n51679;
  assign n51681 = ~n3378 & ~n51680;
  assign n51682 = ~n51675 & ~n51681;
  assign n51683 = n3492 & ~n51682;
  assign n51684 = ~n3631 & ~n51683;
  assign n51685 = n3485 & ~n51684;
  assign n51686 = ~n3630 & ~n51685;
  assign n51687 = ~n3476 & ~n51686;
  assign n51688 = ~n51279 & ~n51683;
  assign n51689 = n3485 & ~n51688;
  assign n51690 = ~n51459 & ~n51689;
  assign n51691 = n3476 & ~n51690;
  assign n51692 = ~n51687 & ~n51691;
  assign n51693 = ~n3374 & ~n51692;
  assign n51694 = n3378 & ~n50878;
  assign n51695 = ~n26705 & ~n37999;
  assign n51696 = controllable_nhgrant0 & ~n51695;
  assign n51697 = ~n8902 & ~n51696;
  assign n51698 = ~n3281 & ~n51697;
  assign n51699 = ~n3950 & ~n51698;
  assign n51700 = ~n3378 & ~n51699;
  assign n51701 = ~n51694 & ~n51700;
  assign n51702 = n3492 & ~n51701;
  assign n51703 = ~n3631 & ~n51702;
  assign n51704 = n3485 & ~n51703;
  assign n51705 = ~n3630 & ~n51704;
  assign n51706 = ~n3476 & ~n51705;
  assign n51707 = n3378 & ~n50896;
  assign n51708 = ~n26720 & ~n38061;
  assign n51709 = controllable_nhgrant0 & ~n51708;
  assign n51710 = ~n9096 & ~n51709;
  assign n51711 = ~n3281 & ~n51710;
  assign n51712 = ~n4089 & ~n51711;
  assign n51713 = ~n3378 & ~n51712;
  assign n51714 = ~n51707 & ~n51713;
  assign n51715 = n3492 & ~n51714;
  assign n51716 = ~n51279 & ~n51715;
  assign n51717 = n3485 & ~n51716;
  assign n51718 = ~n51459 & ~n51717;
  assign n51719 = n3476 & ~n51718;
  assign n51720 = ~n51706 & ~n51719;
  assign n51721 = n3374 & ~n51720;
  assign n51722 = ~n51693 & ~n51721;
  assign n51723 = ~n3655 & ~n51722;
  assign n51724 = ~n51674 & ~n51723;
  assign n51725 = ~n3652 & ~n51724;
  assign n51726 = ~n51625 & ~n51725;
  assign n51727 = ~n3368 & ~n51726;
  assign n51728 = n3378 & ~n50916;
  assign n51729 = ~n26891 & ~n38108;
  assign n51730 = controllable_nhgrant0 & ~n51729;
  assign n51731 = ~n9753 & ~n51730;
  assign n51732 = ~n3281 & ~n51731;
  assign n51733 = ~n3281 & ~n51732;
  assign n51734 = ~n3378 & ~n51733;
  assign n51735 = ~n51728 & ~n51734;
  assign n51736 = n3492 & ~n51735;
  assign n51737 = n3492 & ~n51736;
  assign n51738 = n3485 & ~n51737;
  assign n51739 = n3485 & ~n51738;
  assign n51740 = ~n3476 & ~n51739;
  assign n51741 = ~n8523 & ~n51736;
  assign n51742 = n3485 & ~n51741;
  assign n51743 = ~n8689 & ~n51742;
  assign n51744 = n3476 & ~n51743;
  assign n51745 = ~n51740 & ~n51744;
  assign n51746 = ~n3374 & ~n51745;
  assign n51747 = n3378 & ~n50934;
  assign n51748 = ~n26925 & ~n38180;
  assign n51749 = controllable_nhgrant0 & ~n51748;
  assign n51750 = ~n9861 & ~n51749;
  assign n51751 = ~n3281 & ~n51750;
  assign n51752 = ~n3281 & ~n51751;
  assign n51753 = ~n3378 & ~n51752;
  assign n51754 = ~n51747 & ~n51753;
  assign n51755 = n3492 & ~n51754;
  assign n51756 = n3492 & ~n51755;
  assign n51757 = n3485 & ~n51756;
  assign n51758 = n3485 & ~n51757;
  assign n51759 = ~n3476 & ~n51758;
  assign n51760 = ~n27061 & ~n38275;
  assign n51761 = controllable_nhgrant0 & ~n51760;
  assign n51762 = ~n10071 & ~n51761;
  assign n51763 = ~n3281 & ~n51762;
  assign n51764 = ~n3281 & ~n51763;
  assign n51765 = n3378 & ~n51764;
  assign n51766 = ~n27138 & ~n38365;
  assign n51767 = controllable_nhgrant0 & ~n51766;
  assign n51768 = ~n10240 & ~n51767;
  assign n51769 = ~n3281 & ~n51768;
  assign n51770 = ~n3281 & ~n51769;
  assign n51771 = ~n3378 & ~n51770;
  assign n51772 = ~n51765 & ~n51771;
  assign n51773 = n3492 & ~n51772;
  assign n51774 = ~n51321 & ~n51773;
  assign n51775 = n3485 & ~n51774;
  assign n51776 = ~n51478 & ~n51775;
  assign n51777 = n3476 & ~n51776;
  assign n51778 = ~n51759 & ~n51777;
  assign n51779 = n3374 & ~n51778;
  assign n51780 = ~n51746 & ~n51779;
  assign n51781 = n3655 & ~n51780;
  assign n51782 = n3378 & ~n50968;
  assign n51783 = ~n26891 & ~n38407;
  assign n51784 = controllable_nhgrant0 & ~n51783;
  assign n51785 = ~n9753 & ~n51784;
  assign n51786 = ~n3281 & ~n51785;
  assign n51787 = ~n3281 & ~n51786;
  assign n51788 = ~n3378 & ~n51787;
  assign n51789 = ~n51782 & ~n51788;
  assign n51790 = n3492 & ~n51789;
  assign n51791 = n3492 & ~n51790;
  assign n51792 = n3485 & ~n51791;
  assign n51793 = n3485 & ~n51792;
  assign n51794 = ~n3476 & ~n51793;
  assign n51795 = ~n8523 & ~n51790;
  assign n51796 = n3485 & ~n51795;
  assign n51797 = ~n8689 & ~n51796;
  assign n51798 = n3476 & ~n51797;
  assign n51799 = ~n51794 & ~n51798;
  assign n51800 = ~n3374 & ~n51799;
  assign n51801 = n3378 & ~n50986;
  assign n51802 = ~n26925 & ~n38479;
  assign n51803 = controllable_nhgrant0 & ~n51802;
  assign n51804 = ~n9861 & ~n51803;
  assign n51805 = ~n3281 & ~n51804;
  assign n51806 = ~n3281 & ~n51805;
  assign n51807 = ~n3378 & ~n51806;
  assign n51808 = ~n51801 & ~n51807;
  assign n51809 = n3492 & ~n51808;
  assign n51810 = n3492 & ~n51809;
  assign n51811 = n3485 & ~n51810;
  assign n51812 = n3485 & ~n51811;
  assign n51813 = ~n3476 & ~n51812;
  assign n51814 = ~n27061 & ~n38574;
  assign n51815 = controllable_nhgrant0 & ~n51814;
  assign n51816 = ~n10071 & ~n51815;
  assign n51817 = ~n3281 & ~n51816;
  assign n51818 = ~n3281 & ~n51817;
  assign n51819 = n3378 & ~n51818;
  assign n51820 = ~n27138 & ~n38653;
  assign n51821 = controllable_nhgrant0 & ~n51820;
  assign n51822 = ~n10240 & ~n51821;
  assign n51823 = ~n3281 & ~n51822;
  assign n51824 = ~n3281 & ~n51823;
  assign n51825 = ~n3378 & ~n51824;
  assign n51826 = ~n51819 & ~n51825;
  assign n51827 = n3492 & ~n51826;
  assign n51828 = ~n51348 & ~n51827;
  assign n51829 = n3485 & ~n51828;
  assign n51830 = ~n51489 & ~n51829;
  assign n51831 = n3476 & ~n51830;
  assign n51832 = ~n51813 & ~n51831;
  assign n51833 = n3374 & ~n51832;
  assign n51834 = ~n51800 & ~n51833;
  assign n51835 = ~n3655 & ~n51834;
  assign n51836 = ~n51781 & ~n51835;
  assign n51837 = n3652 & ~n51836;
  assign n51838 = n3378 & ~n51022;
  assign n51839 = ~n26891 & ~n38690;
  assign n51840 = controllable_nhgrant0 & ~n51839;
  assign n51841 = ~n9753 & ~n51840;
  assign n51842 = ~n3281 & ~n51841;
  assign n51843 = ~n3281 & ~n51842;
  assign n51844 = ~n3378 & ~n51843;
  assign n51845 = ~n51838 & ~n51844;
  assign n51846 = n3492 & ~n51845;
  assign n51847 = n3492 & ~n51846;
  assign n51848 = n3485 & ~n51847;
  assign n51849 = n3485 & ~n51848;
  assign n51850 = ~n3476 & ~n51849;
  assign n51851 = ~n8523 & ~n51846;
  assign n51852 = n3485 & ~n51851;
  assign n51853 = ~n8689 & ~n51852;
  assign n51854 = n3476 & ~n51853;
  assign n51855 = ~n51850 & ~n51854;
  assign n51856 = ~n3374 & ~n51855;
  assign n51857 = n3378 & ~n51040;
  assign n51858 = ~n26925 & ~n38748;
  assign n51859 = controllable_nhgrant0 & ~n51858;
  assign n51860 = ~n9861 & ~n51859;
  assign n51861 = ~n3281 & ~n51860;
  assign n51862 = ~n3281 & ~n51861;
  assign n51863 = ~n3378 & ~n51862;
  assign n51864 = ~n51857 & ~n51863;
  assign n51865 = n3492 & ~n51864;
  assign n51866 = n3492 & ~n51865;
  assign n51867 = n3485 & ~n51866;
  assign n51868 = n3485 & ~n51867;
  assign n51869 = ~n3476 & ~n51868;
  assign n51870 = ~n27061 & ~n38811;
  assign n51871 = controllable_nhgrant0 & ~n51870;
  assign n51872 = ~n10071 & ~n51871;
  assign n51873 = ~n3281 & ~n51872;
  assign n51874 = ~n3281 & ~n51873;
  assign n51875 = n3378 & ~n51874;
  assign n51876 = ~n27138 & ~n38864;
  assign n51877 = controllable_nhgrant0 & ~n51876;
  assign n51878 = ~n10240 & ~n51877;
  assign n51879 = ~n3281 & ~n51878;
  assign n51880 = ~n3281 & ~n51879;
  assign n51881 = ~n3378 & ~n51880;
  assign n51882 = ~n51875 & ~n51881;
  assign n51883 = n3492 & ~n51882;
  assign n51884 = ~n51377 & ~n51883;
  assign n51885 = n3485 & ~n51884;
  assign n51886 = ~n51502 & ~n51885;
  assign n51887 = n3476 & ~n51886;
  assign n51888 = ~n51869 & ~n51887;
  assign n51889 = n3374 & ~n51888;
  assign n51890 = ~n51856 & ~n51889;
  assign n51891 = n3655 & ~n51890;
  assign n51892 = n3378 & ~n51074;
  assign n51893 = ~n26891 & ~n38899;
  assign n51894 = controllable_nhgrant0 & ~n51893;
  assign n51895 = ~n9753 & ~n51894;
  assign n51896 = ~n3281 & ~n51895;
  assign n51897 = ~n3281 & ~n51896;
  assign n51898 = ~n3378 & ~n51897;
  assign n51899 = ~n51892 & ~n51898;
  assign n51900 = n3492 & ~n51899;
  assign n51901 = n3492 & ~n51900;
  assign n51902 = n3485 & ~n51901;
  assign n51903 = n3485 & ~n51902;
  assign n51904 = ~n3476 & ~n51903;
  assign n51905 = ~n8523 & ~n51900;
  assign n51906 = n3485 & ~n51905;
  assign n51907 = ~n8689 & ~n51906;
  assign n51908 = n3476 & ~n51907;
  assign n51909 = ~n51904 & ~n51908;
  assign n51910 = ~n3374 & ~n51909;
  assign n51911 = n3378 & ~n51092;
  assign n51912 = ~n26925 & ~n38957;
  assign n51913 = controllable_nhgrant0 & ~n51912;
  assign n51914 = ~n9861 & ~n51913;
  assign n51915 = ~n3281 & ~n51914;
  assign n51916 = ~n3281 & ~n51915;
  assign n51917 = ~n3378 & ~n51916;
  assign n51918 = ~n51911 & ~n51917;
  assign n51919 = n3492 & ~n51918;
  assign n51920 = n3492 & ~n51919;
  assign n51921 = n3485 & ~n51920;
  assign n51922 = n3485 & ~n51921;
  assign n51923 = ~n3476 & ~n51922;
  assign n51924 = ~n27061 & ~n39020;
  assign n51925 = controllable_nhgrant0 & ~n51924;
  assign n51926 = ~n10071 & ~n51925;
  assign n51927 = ~n3281 & ~n51926;
  assign n51928 = ~n3281 & ~n51927;
  assign n51929 = n3378 & ~n51928;
  assign n51930 = ~n27138 & ~n39073;
  assign n51931 = controllable_nhgrant0 & ~n51930;
  assign n51932 = ~n10240 & ~n51931;
  assign n51933 = ~n3281 & ~n51932;
  assign n51934 = ~n3281 & ~n51933;
  assign n51935 = ~n3378 & ~n51934;
  assign n51936 = ~n51929 & ~n51935;
  assign n51937 = n3492 & ~n51936;
  assign n51938 = ~n51404 & ~n51937;
  assign n51939 = n3485 & ~n51938;
  assign n51940 = ~n51513 & ~n51939;
  assign n51941 = n3476 & ~n51940;
  assign n51942 = ~n51923 & ~n51941;
  assign n51943 = n3374 & ~n51942;
  assign n51944 = ~n51910 & ~n51943;
  assign n51945 = ~n3655 & ~n51944;
  assign n51946 = ~n51891 & ~n51945;
  assign n51947 = ~n3652 & ~n51946;
  assign n51948 = ~n51837 & ~n51947;
  assign n51949 = n3368 & ~n51948;
  assign n51950 = ~n51727 & ~n51949;
  assign n51951 = ~n3362 & ~n51950;
  assign n51952 = ~n51525 & ~n51951;
  assign n51953 = ~n3359 & ~n51952;
  assign n51954 = ~n51423 & ~n51953;
  assign n51955 = ~n3356 & ~n51954;
  assign n51956 = ~n50673 & ~n51955;
  assign n51957 = n3345 & ~n51956;
  assign n51958 = ~n3649 & ~n51957;
  assign n51959 = ~n3341 & ~n51958;
  assign n51960 = ~n27406 & ~n39115;
  assign n51961 = controllable_nhgrant0 & ~n51960;
  assign n51962 = ~n11496 & ~n51961;
  assign n51963 = ~n3281 & ~n51962;
  assign n51964 = ~n3281 & ~n51963;
  assign n51965 = n3378 & ~n51964;
  assign n51966 = ~n27414 & ~n39123;
  assign n51967 = controllable_nhgrant0 & ~n51966;
  assign n51968 = ~n11512 & ~n51967;
  assign n51969 = ~n3281 & ~n51968;
  assign n51970 = ~n3950 & ~n51969;
  assign n51971 = ~n3378 & ~n51970;
  assign n51972 = ~n51965 & ~n51971;
  assign n51973 = n3492 & ~n51972;
  assign n51974 = ~n3493 & ~n51973;
  assign n51975 = n3485 & ~n51974;
  assign n51976 = ~n3486 & ~n51975;
  assign n51977 = ~n3476 & ~n51976;
  assign n51978 = ~n27440 & ~n39115;
  assign n51979 = controllable_nhgrant0 & ~n51978;
  assign n51980 = ~n11496 & ~n51979;
  assign n51981 = ~n3281 & ~n51980;
  assign n51982 = ~n3281 & ~n51981;
  assign n51983 = n3378 & ~n51982;
  assign n51984 = ~n27458 & ~n39164;
  assign n51985 = controllable_nhgrant0 & ~n51984;
  assign n51986 = ~n11512 & ~n51985;
  assign n51987 = ~n3281 & ~n51986;
  assign n51988 = ~n4089 & ~n51987;
  assign n51989 = ~n3378 & ~n51988;
  assign n51990 = ~n51983 & ~n51989;
  assign n51991 = n3492 & ~n51990;
  assign n51992 = ~n27390 & ~n51991;
  assign n51993 = n3485 & ~n51992;
  assign n51994 = ~n27389 & ~n51993;
  assign n51995 = n3476 & ~n51994;
  assign n51996 = ~n51977 & ~n51995;
  assign n51997 = n3374 & ~n51996;
  assign n51998 = ~n27396 & ~n51997;
  assign n51999 = n3655 & ~n51998;
  assign n52000 = ~n27406 & ~n39192;
  assign n52001 = controllable_nhgrant0 & ~n52000;
  assign n52002 = ~n11496 & ~n52001;
  assign n52003 = ~n3281 & ~n52002;
  assign n52004 = ~n3281 & ~n52003;
  assign n52005 = n3378 & ~n52004;
  assign n52006 = ~n27414 & ~n39200;
  assign n52007 = controllable_nhgrant0 & ~n52006;
  assign n52008 = ~n11512 & ~n52007;
  assign n52009 = ~n3281 & ~n52008;
  assign n52010 = ~n3950 & ~n52009;
  assign n52011 = ~n3378 & ~n52010;
  assign n52012 = ~n52005 & ~n52011;
  assign n52013 = n3492 & ~n52012;
  assign n52014 = ~n3493 & ~n52013;
  assign n52015 = n3485 & ~n52014;
  assign n52016 = ~n3486 & ~n52015;
  assign n52017 = ~n3476 & ~n52016;
  assign n52018 = ~n27440 & ~n39192;
  assign n52019 = controllable_nhgrant0 & ~n52018;
  assign n52020 = ~n11496 & ~n52019;
  assign n52021 = ~n3281 & ~n52020;
  assign n52022 = ~n3281 & ~n52021;
  assign n52023 = n3378 & ~n52022;
  assign n52024 = ~n27458 & ~n39241;
  assign n52025 = controllable_nhgrant0 & ~n52024;
  assign n52026 = ~n11512 & ~n52025;
  assign n52027 = ~n3281 & ~n52026;
  assign n52028 = ~n4089 & ~n52027;
  assign n52029 = ~n3378 & ~n52028;
  assign n52030 = ~n52023 & ~n52029;
  assign n52031 = n3492 & ~n52030;
  assign n52032 = ~n27390 & ~n52031;
  assign n52033 = n3485 & ~n52032;
  assign n52034 = ~n27389 & ~n52033;
  assign n52035 = n3476 & ~n52034;
  assign n52036 = ~n52017 & ~n52035;
  assign n52037 = n3374 & ~n52036;
  assign n52038 = ~n27396 & ~n52037;
  assign n52039 = ~n3655 & ~n52038;
  assign n52040 = ~n51999 & ~n52039;
  assign n52041 = n3652 & ~n52040;
  assign n52042 = ~n27406 & ~n39271;
  assign n52043 = controllable_nhgrant0 & ~n52042;
  assign n52044 = ~n11496 & ~n52043;
  assign n52045 = ~n3281 & ~n52044;
  assign n52046 = ~n3281 & ~n52045;
  assign n52047 = n3378 & ~n52046;
  assign n52048 = ~n27414 & ~n39279;
  assign n52049 = controllable_nhgrant0 & ~n52048;
  assign n52050 = ~n11512 & ~n52049;
  assign n52051 = ~n3281 & ~n52050;
  assign n52052 = ~n3950 & ~n52051;
  assign n52053 = ~n3378 & ~n52052;
  assign n52054 = ~n52047 & ~n52053;
  assign n52055 = n3492 & ~n52054;
  assign n52056 = ~n3493 & ~n52055;
  assign n52057 = n3485 & ~n52056;
  assign n52058 = ~n3486 & ~n52057;
  assign n52059 = ~n3476 & ~n52058;
  assign n52060 = ~n27440 & ~n39271;
  assign n52061 = controllable_nhgrant0 & ~n52060;
  assign n52062 = ~n11496 & ~n52061;
  assign n52063 = ~n3281 & ~n52062;
  assign n52064 = ~n3281 & ~n52063;
  assign n52065 = n3378 & ~n52064;
  assign n52066 = ~n27458 & ~n39313;
  assign n52067 = controllable_nhgrant0 & ~n52066;
  assign n52068 = ~n11512 & ~n52067;
  assign n52069 = ~n3281 & ~n52068;
  assign n52070 = ~n4089 & ~n52069;
  assign n52071 = ~n3378 & ~n52070;
  assign n52072 = ~n52065 & ~n52071;
  assign n52073 = n3492 & ~n52072;
  assign n52074 = ~n27390 & ~n52073;
  assign n52075 = n3485 & ~n52074;
  assign n52076 = ~n27389 & ~n52075;
  assign n52077 = n3476 & ~n52076;
  assign n52078 = ~n52059 & ~n52077;
  assign n52079 = n3374 & ~n52078;
  assign n52080 = ~n27396 & ~n52079;
  assign n52081 = n3655 & ~n52080;
  assign n52082 = ~n27406 & ~n39341;
  assign n52083 = controllable_nhgrant0 & ~n52082;
  assign n52084 = ~n11496 & ~n52083;
  assign n52085 = ~n3281 & ~n52084;
  assign n52086 = ~n3281 & ~n52085;
  assign n52087 = n3378 & ~n52086;
  assign n52088 = ~n27414 & ~n39349;
  assign n52089 = controllable_nhgrant0 & ~n52088;
  assign n52090 = ~n11512 & ~n52089;
  assign n52091 = ~n3281 & ~n52090;
  assign n52092 = ~n3950 & ~n52091;
  assign n52093 = ~n3378 & ~n52092;
  assign n52094 = ~n52087 & ~n52093;
  assign n52095 = n3492 & ~n52094;
  assign n52096 = ~n3493 & ~n52095;
  assign n52097 = n3485 & ~n52096;
  assign n52098 = ~n3486 & ~n52097;
  assign n52099 = ~n3476 & ~n52098;
  assign n52100 = ~n27440 & ~n39341;
  assign n52101 = controllable_nhgrant0 & ~n52100;
  assign n52102 = ~n11496 & ~n52101;
  assign n52103 = ~n3281 & ~n52102;
  assign n52104 = ~n3281 & ~n52103;
  assign n52105 = n3378 & ~n52104;
  assign n52106 = ~n27458 & ~n39383;
  assign n52107 = controllable_nhgrant0 & ~n52106;
  assign n52108 = ~n11512 & ~n52107;
  assign n52109 = ~n3281 & ~n52108;
  assign n52110 = ~n4089 & ~n52109;
  assign n52111 = ~n3378 & ~n52110;
  assign n52112 = ~n52105 & ~n52111;
  assign n52113 = n3492 & ~n52112;
  assign n52114 = ~n27390 & ~n52113;
  assign n52115 = n3485 & ~n52114;
  assign n52116 = ~n27389 & ~n52115;
  assign n52117 = n3476 & ~n52116;
  assign n52118 = ~n52099 & ~n52117;
  assign n52119 = n3374 & ~n52118;
  assign n52120 = ~n27396 & ~n52119;
  assign n52121 = ~n3655 & ~n52120;
  assign n52122 = ~n52081 & ~n52121;
  assign n52123 = ~n3652 & ~n52122;
  assign n52124 = ~n52041 & ~n52123;
  assign n52125 = ~n3368 & ~n52124;
  assign n52126 = ~n27610 & ~n39415;
  assign n52127 = controllable_nhgrant0 & ~n52126;
  assign n52128 = ~n11874 & ~n52127;
  assign n52129 = ~n3281 & ~n52128;
  assign n52130 = ~n3281 & ~n52129;
  assign n52131 = n3492 & ~n52130;
  assign n52132 = n3492 & ~n52131;
  assign n52133 = n3485 & ~n52132;
  assign n52134 = n3485 & ~n52133;
  assign n52135 = ~n3476 & ~n52134;
  assign n52136 = ~n27657 & ~n39415;
  assign n52137 = controllable_nhgrant0 & ~n52136;
  assign n52138 = ~n11874 & ~n52137;
  assign n52139 = ~n3281 & ~n52138;
  assign n52140 = ~n3281 & ~n52139;
  assign n52141 = n3492 & ~n52140;
  assign n52142 = ~n27622 & ~n52141;
  assign n52143 = n3485 & ~n52142;
  assign n52144 = ~n27621 & ~n52143;
  assign n52145 = n3476 & ~n52144;
  assign n52146 = ~n52135 & ~n52145;
  assign n52147 = n3374 & ~n52146;
  assign n52148 = n3374 & ~n52147;
  assign n52149 = n3655 & ~n52148;
  assign n52150 = ~n27610 & ~n39451;
  assign n52151 = controllable_nhgrant0 & ~n52150;
  assign n52152 = ~n11874 & ~n52151;
  assign n52153 = ~n3281 & ~n52152;
  assign n52154 = ~n3281 & ~n52153;
  assign n52155 = n3492 & ~n52154;
  assign n52156 = n3492 & ~n52155;
  assign n52157 = n3485 & ~n52156;
  assign n52158 = n3485 & ~n52157;
  assign n52159 = ~n3476 & ~n52158;
  assign n52160 = ~n27657 & ~n39451;
  assign n52161 = controllable_nhgrant0 & ~n52160;
  assign n52162 = ~n11874 & ~n52161;
  assign n52163 = ~n3281 & ~n52162;
  assign n52164 = ~n3281 & ~n52163;
  assign n52165 = n3492 & ~n52164;
  assign n52166 = ~n27622 & ~n52165;
  assign n52167 = n3485 & ~n52166;
  assign n52168 = ~n27621 & ~n52167;
  assign n52169 = n3476 & ~n52168;
  assign n52170 = ~n52159 & ~n52169;
  assign n52171 = n3374 & ~n52170;
  assign n52172 = n3374 & ~n52171;
  assign n52173 = ~n3655 & ~n52172;
  assign n52174 = ~n52149 & ~n52173;
  assign n52175 = n3652 & ~n52174;
  assign n52176 = ~n27610 & ~n39489;
  assign n52177 = controllable_nhgrant0 & ~n52176;
  assign n52178 = ~n11874 & ~n52177;
  assign n52179 = ~n3281 & ~n52178;
  assign n52180 = ~n3281 & ~n52179;
  assign n52181 = n3492 & ~n52180;
  assign n52182 = n3492 & ~n52181;
  assign n52183 = n3485 & ~n52182;
  assign n52184 = n3485 & ~n52183;
  assign n52185 = ~n3476 & ~n52184;
  assign n52186 = ~n27657 & ~n39489;
  assign n52187 = controllable_nhgrant0 & ~n52186;
  assign n52188 = ~n11874 & ~n52187;
  assign n52189 = ~n3281 & ~n52188;
  assign n52190 = ~n3281 & ~n52189;
  assign n52191 = n3492 & ~n52190;
  assign n52192 = ~n27622 & ~n52191;
  assign n52193 = n3485 & ~n52192;
  assign n52194 = ~n27621 & ~n52193;
  assign n52195 = n3476 & ~n52194;
  assign n52196 = ~n52185 & ~n52195;
  assign n52197 = n3374 & ~n52196;
  assign n52198 = n3374 & ~n52197;
  assign n52199 = n3655 & ~n52198;
  assign n52200 = ~n27610 & ~n39525;
  assign n52201 = controllable_nhgrant0 & ~n52200;
  assign n52202 = ~n11874 & ~n52201;
  assign n52203 = ~n3281 & ~n52202;
  assign n52204 = ~n3281 & ~n52203;
  assign n52205 = n3492 & ~n52204;
  assign n52206 = n3492 & ~n52205;
  assign n52207 = n3485 & ~n52206;
  assign n52208 = n3485 & ~n52207;
  assign n52209 = ~n3476 & ~n52208;
  assign n52210 = ~n27657 & ~n39525;
  assign n52211 = controllable_nhgrant0 & ~n52210;
  assign n52212 = ~n11874 & ~n52211;
  assign n52213 = ~n3281 & ~n52212;
  assign n52214 = ~n3281 & ~n52213;
  assign n52215 = n3492 & ~n52214;
  assign n52216 = ~n27622 & ~n52215;
  assign n52217 = n3485 & ~n52216;
  assign n52218 = ~n27621 & ~n52217;
  assign n52219 = n3476 & ~n52218;
  assign n52220 = ~n52209 & ~n52219;
  assign n52221 = n3374 & ~n52220;
  assign n52222 = n3374 & ~n52221;
  assign n52223 = ~n3655 & ~n52222;
  assign n52224 = ~n52199 & ~n52223;
  assign n52225 = ~n3652 & ~n52224;
  assign n52226 = ~n52175 & ~n52225;
  assign n52227 = n3368 & ~n52226;
  assign n52228 = ~n52125 & ~n52227;
  assign n52229 = ~n3362 & ~n52228;
  assign n52230 = ~n3362 & ~n52229;
  assign n52231 = ~n3359 & ~n52230;
  assign n52232 = ~n3359 & ~n52231;
  assign n52233 = n3356 & ~n52232;
  assign n52234 = ~n27765 & ~n39584;
  assign n52235 = controllable_nhgrant0 & ~n52234;
  assign n52236 = ~n5245 & ~n52235;
  assign n52237 = ~n3281 & ~n52236;
  assign n52238 = ~n3783 & ~n52237;
  assign n52239 = ~n3378 & ~n52238;
  assign n52240 = ~n27756 & ~n52239;
  assign n52241 = n3492 & ~n52240;
  assign n52242 = ~n3631 & ~n52241;
  assign n52243 = n3485 & ~n52242;
  assign n52244 = ~n3630 & ~n52243;
  assign n52245 = ~n3476 & ~n52244;
  assign n52246 = ~n27779 & ~n52241;
  assign n52247 = n3485 & ~n52246;
  assign n52248 = ~n27778 & ~n52247;
  assign n52249 = n3476 & ~n52248;
  assign n52250 = ~n52245 & ~n52249;
  assign n52251 = ~n3374 & ~n52250;
  assign n52252 = ~n27803 & ~n39608;
  assign n52253 = controllable_nhgrant0 & ~n52252;
  assign n52254 = ~n12101 & ~n52253;
  assign n52255 = ~n3281 & ~n52254;
  assign n52256 = ~n3950 & ~n52255;
  assign n52257 = n3378 & ~n52256;
  assign n52258 = ~n27817 & ~n39660;
  assign n52259 = controllable_nhgrant0 & ~n52258;
  assign n52260 = ~n5534 & ~n52259;
  assign n52261 = ~n3281 & ~n52260;
  assign n52262 = ~n3950 & ~n52261;
  assign n52263 = ~n3378 & ~n52262;
  assign n52264 = ~n52257 & ~n52263;
  assign n52265 = n3492 & ~n52264;
  assign n52266 = ~n3631 & ~n52265;
  assign n52267 = n3485 & ~n52266;
  assign n52268 = ~n3630 & ~n52267;
  assign n52269 = ~n3476 & ~n52268;
  assign n52270 = ~n27847 & ~n39697;
  assign n52271 = controllable_nhgrant0 & ~n52270;
  assign n52272 = ~n12249 & ~n52271;
  assign n52273 = ~n3281 & ~n52272;
  assign n52274 = ~n4089 & ~n52273;
  assign n52275 = n3378 & ~n52274;
  assign n52276 = ~n27865 & ~n39750;
  assign n52277 = controllable_nhgrant0 & ~n52276;
  assign n52278 = ~n6082 & ~n52277;
  assign n52279 = ~n3281 & ~n52278;
  assign n52280 = ~n4089 & ~n52279;
  assign n52281 = ~n3378 & ~n52280;
  assign n52282 = ~n52275 & ~n52281;
  assign n52283 = n3492 & ~n52282;
  assign n52284 = ~n27779 & ~n52283;
  assign n52285 = n3485 & ~n52284;
  assign n52286 = ~n27778 & ~n52285;
  assign n52287 = n3476 & ~n52286;
  assign n52288 = ~n52269 & ~n52287;
  assign n52289 = n3374 & ~n52288;
  assign n52290 = ~n52251 & ~n52289;
  assign n52291 = n3655 & ~n52290;
  assign n52292 = ~n27765 & ~n39791;
  assign n52293 = controllable_nhgrant0 & ~n52292;
  assign n52294 = ~n5245 & ~n52293;
  assign n52295 = ~n3281 & ~n52294;
  assign n52296 = ~n3783 & ~n52295;
  assign n52297 = ~n3378 & ~n52296;
  assign n52298 = ~n27756 & ~n52297;
  assign n52299 = n3492 & ~n52298;
  assign n52300 = ~n3631 & ~n52299;
  assign n52301 = n3485 & ~n52300;
  assign n52302 = ~n3630 & ~n52301;
  assign n52303 = ~n3476 & ~n52302;
  assign n52304 = ~n27779 & ~n52299;
  assign n52305 = n3485 & ~n52304;
  assign n52306 = ~n27778 & ~n52305;
  assign n52307 = n3476 & ~n52306;
  assign n52308 = ~n52303 & ~n52307;
  assign n52309 = ~n3374 & ~n52308;
  assign n52310 = ~n27803 & ~n39815;
  assign n52311 = controllable_nhgrant0 & ~n52310;
  assign n52312 = ~n12101 & ~n52311;
  assign n52313 = ~n3281 & ~n52312;
  assign n52314 = ~n3950 & ~n52313;
  assign n52315 = n3378 & ~n52314;
  assign n52316 = ~n27817 & ~n39867;
  assign n52317 = controllable_nhgrant0 & ~n52316;
  assign n52318 = ~n5534 & ~n52317;
  assign n52319 = ~n3281 & ~n52318;
  assign n52320 = ~n3950 & ~n52319;
  assign n52321 = ~n3378 & ~n52320;
  assign n52322 = ~n52315 & ~n52321;
  assign n52323 = n3492 & ~n52322;
  assign n52324 = ~n3631 & ~n52323;
  assign n52325 = n3485 & ~n52324;
  assign n52326 = ~n3630 & ~n52325;
  assign n52327 = ~n3476 & ~n52326;
  assign n52328 = ~n27847 & ~n39902;
  assign n52329 = controllable_nhgrant0 & ~n52328;
  assign n52330 = ~n12249 & ~n52329;
  assign n52331 = ~n3281 & ~n52330;
  assign n52332 = ~n4089 & ~n52331;
  assign n52333 = n3378 & ~n52332;
  assign n52334 = ~n27865 & ~n39955;
  assign n52335 = controllable_nhgrant0 & ~n52334;
  assign n52336 = ~n6082 & ~n52335;
  assign n52337 = ~n3281 & ~n52336;
  assign n52338 = ~n4089 & ~n52337;
  assign n52339 = ~n3378 & ~n52338;
  assign n52340 = ~n52333 & ~n52339;
  assign n52341 = n3492 & ~n52340;
  assign n52342 = ~n27779 & ~n52341;
  assign n52343 = n3485 & ~n52342;
  assign n52344 = ~n27778 & ~n52343;
  assign n52345 = n3476 & ~n52344;
  assign n52346 = ~n52327 & ~n52345;
  assign n52347 = n3374 & ~n52346;
  assign n52348 = ~n52309 & ~n52347;
  assign n52349 = ~n3655 & ~n52348;
  assign n52350 = ~n52291 & ~n52349;
  assign n52351 = n3652 & ~n52350;
  assign n52352 = ~n27765 & ~n39991;
  assign n52353 = controllable_nhgrant0 & ~n52352;
  assign n52354 = ~n5245 & ~n52353;
  assign n52355 = ~n3281 & ~n52354;
  assign n52356 = ~n3783 & ~n52355;
  assign n52357 = ~n3378 & ~n52356;
  assign n52358 = ~n27756 & ~n52357;
  assign n52359 = n3492 & ~n52358;
  assign n52360 = ~n3631 & ~n52359;
  assign n52361 = n3485 & ~n52360;
  assign n52362 = ~n3630 & ~n52361;
  assign n52363 = ~n3476 & ~n52362;
  assign n52364 = ~n27779 & ~n52359;
  assign n52365 = n3485 & ~n52364;
  assign n52366 = ~n27778 & ~n52365;
  assign n52367 = n3476 & ~n52366;
  assign n52368 = ~n52363 & ~n52367;
  assign n52369 = ~n3374 & ~n52368;
  assign n52370 = ~n27803 & ~n40015;
  assign n52371 = controllable_nhgrant0 & ~n52370;
  assign n52372 = ~n12101 & ~n52371;
  assign n52373 = ~n3281 & ~n52372;
  assign n52374 = ~n3950 & ~n52373;
  assign n52375 = n3378 & ~n52374;
  assign n52376 = ~n27817 & ~n40053;
  assign n52377 = controllable_nhgrant0 & ~n52376;
  assign n52378 = ~n5534 & ~n52377;
  assign n52379 = ~n3281 & ~n52378;
  assign n52380 = ~n3950 & ~n52379;
  assign n52381 = ~n3378 & ~n52380;
  assign n52382 = ~n52375 & ~n52381;
  assign n52383 = n3492 & ~n52382;
  assign n52384 = ~n3631 & ~n52383;
  assign n52385 = n3485 & ~n52384;
  assign n52386 = ~n3630 & ~n52385;
  assign n52387 = ~n3476 & ~n52386;
  assign n52388 = ~n27847 & ~n40081;
  assign n52389 = controllable_nhgrant0 & ~n52388;
  assign n52390 = ~n12249 & ~n52389;
  assign n52391 = ~n3281 & ~n52390;
  assign n52392 = ~n4089 & ~n52391;
  assign n52393 = n3378 & ~n52392;
  assign n52394 = ~n27865 & ~n40119;
  assign n52395 = controllable_nhgrant0 & ~n52394;
  assign n52396 = ~n6082 & ~n52395;
  assign n52397 = ~n3281 & ~n52396;
  assign n52398 = ~n4089 & ~n52397;
  assign n52399 = ~n3378 & ~n52398;
  assign n52400 = ~n52393 & ~n52399;
  assign n52401 = n3492 & ~n52400;
  assign n52402 = ~n27779 & ~n52401;
  assign n52403 = n3485 & ~n52402;
  assign n52404 = ~n27778 & ~n52403;
  assign n52405 = n3476 & ~n52404;
  assign n52406 = ~n52387 & ~n52405;
  assign n52407 = n3374 & ~n52406;
  assign n52408 = ~n52369 & ~n52407;
  assign n52409 = n3655 & ~n52408;
  assign n52410 = ~n27765 & ~n40153;
  assign n52411 = controllable_nhgrant0 & ~n52410;
  assign n52412 = ~n5245 & ~n52411;
  assign n52413 = ~n3281 & ~n52412;
  assign n52414 = ~n3783 & ~n52413;
  assign n52415 = ~n3378 & ~n52414;
  assign n52416 = ~n27756 & ~n52415;
  assign n52417 = n3492 & ~n52416;
  assign n52418 = ~n3631 & ~n52417;
  assign n52419 = n3485 & ~n52418;
  assign n52420 = ~n3630 & ~n52419;
  assign n52421 = ~n3476 & ~n52420;
  assign n52422 = ~n27779 & ~n52417;
  assign n52423 = n3485 & ~n52422;
  assign n52424 = ~n27778 & ~n52423;
  assign n52425 = n3476 & ~n52424;
  assign n52426 = ~n52421 & ~n52425;
  assign n52427 = ~n3374 & ~n52426;
  assign n52428 = ~n27803 & ~n40177;
  assign n52429 = controllable_nhgrant0 & ~n52428;
  assign n52430 = ~n12101 & ~n52429;
  assign n52431 = ~n3281 & ~n52430;
  assign n52432 = ~n3950 & ~n52431;
  assign n52433 = n3378 & ~n52432;
  assign n52434 = ~n27817 & ~n40215;
  assign n52435 = controllable_nhgrant0 & ~n52434;
  assign n52436 = ~n5534 & ~n52435;
  assign n52437 = ~n3281 & ~n52436;
  assign n52438 = ~n3950 & ~n52437;
  assign n52439 = ~n3378 & ~n52438;
  assign n52440 = ~n52433 & ~n52439;
  assign n52441 = n3492 & ~n52440;
  assign n52442 = ~n3631 & ~n52441;
  assign n52443 = n3485 & ~n52442;
  assign n52444 = ~n3630 & ~n52443;
  assign n52445 = ~n3476 & ~n52444;
  assign n52446 = ~n27847 & ~n40243;
  assign n52447 = controllable_nhgrant0 & ~n52446;
  assign n52448 = ~n12249 & ~n52447;
  assign n52449 = ~n3281 & ~n52448;
  assign n52450 = ~n4089 & ~n52449;
  assign n52451 = n3378 & ~n52450;
  assign n52452 = ~n27865 & ~n40281;
  assign n52453 = controllable_nhgrant0 & ~n52452;
  assign n52454 = ~n6082 & ~n52453;
  assign n52455 = ~n3281 & ~n52454;
  assign n52456 = ~n4089 & ~n52455;
  assign n52457 = ~n3378 & ~n52456;
  assign n52458 = ~n52451 & ~n52457;
  assign n52459 = n3492 & ~n52458;
  assign n52460 = ~n27779 & ~n52459;
  assign n52461 = n3485 & ~n52460;
  assign n52462 = ~n27778 & ~n52461;
  assign n52463 = n3476 & ~n52462;
  assign n52464 = ~n52445 & ~n52463;
  assign n52465 = n3374 & ~n52464;
  assign n52466 = ~n52427 & ~n52465;
  assign n52467 = ~n3655 & ~n52466;
  assign n52468 = ~n52409 & ~n52467;
  assign n52469 = ~n3652 & ~n52468;
  assign n52470 = ~n52351 & ~n52469;
  assign n52471 = ~n3368 & ~n52470;
  assign n52472 = ~n28091 & ~n40313;
  assign n52473 = controllable_nhgrant0 & ~n52472;
  assign n52474 = ~n7118 & ~n52473;
  assign n52475 = ~n3281 & ~n52474;
  assign n52476 = ~n3281 & ~n52475;
  assign n52477 = ~n3378 & ~n52476;
  assign n52478 = ~n28079 & ~n52477;
  assign n52479 = n3492 & ~n52478;
  assign n52480 = n3492 & ~n52479;
  assign n52481 = n3485 & ~n52480;
  assign n52482 = n3485 & ~n52481;
  assign n52483 = ~n3374 & ~n52482;
  assign n52484 = ~n28116 & ~n40337;
  assign n52485 = controllable_nhgrant0 & ~n52484;
  assign n52486 = ~n12773 & ~n52485;
  assign n52487 = ~n3281 & ~n52486;
  assign n52488 = ~n3281 & ~n52487;
  assign n52489 = n3378 & ~n52488;
  assign n52490 = ~n28139 & ~n40365;
  assign n52491 = controllable_nhgrant0 & ~n52490;
  assign n52492 = ~n12827 & ~n52491;
  assign n52493 = ~n3281 & ~n52492;
  assign n52494 = ~n3281 & ~n52493;
  assign n52495 = ~n3378 & ~n52494;
  assign n52496 = ~n52489 & ~n52495;
  assign n52497 = n3492 & ~n52496;
  assign n52498 = n3492 & ~n52497;
  assign n52499 = n3485 & ~n52498;
  assign n52500 = n3485 & ~n52499;
  assign n52501 = ~n3476 & ~n52500;
  assign n52502 = ~n28183 & ~n40402;
  assign n52503 = controllable_nhgrant0 & ~n52502;
  assign n52504 = ~n12942 & ~n52503;
  assign n52505 = ~n3281 & ~n52504;
  assign n52506 = ~n3281 & ~n52505;
  assign n52507 = n3378 & ~n52506;
  assign n52508 = ~n28235 & ~n40501;
  assign n52509 = controllable_nhgrant0 & ~n52508;
  assign n52510 = ~n13064 & ~n52509;
  assign n52511 = ~n3281 & ~n52510;
  assign n52512 = ~n3281 & ~n52511;
  assign n52513 = ~n3378 & ~n52512;
  assign n52514 = ~n52507 & ~n52513;
  assign n52515 = n3492 & ~n52514;
  assign n52516 = ~n27622 & ~n52515;
  assign n52517 = n3485 & ~n52516;
  assign n52518 = ~n27621 & ~n52517;
  assign n52519 = n3476 & ~n52518;
  assign n52520 = ~n52501 & ~n52519;
  assign n52521 = n3374 & ~n52520;
  assign n52522 = ~n52483 & ~n52521;
  assign n52523 = n3655 & ~n52522;
  assign n52524 = ~n28091 & ~n40529;
  assign n52525 = controllable_nhgrant0 & ~n52524;
  assign n52526 = ~n7118 & ~n52525;
  assign n52527 = ~n3281 & ~n52526;
  assign n52528 = ~n3281 & ~n52527;
  assign n52529 = ~n3378 & ~n52528;
  assign n52530 = ~n28079 & ~n52529;
  assign n52531 = n3492 & ~n52530;
  assign n52532 = n3492 & ~n52531;
  assign n52533 = n3485 & ~n52532;
  assign n52534 = n3485 & ~n52533;
  assign n52535 = ~n3374 & ~n52534;
  assign n52536 = ~n28116 & ~n40553;
  assign n52537 = controllable_nhgrant0 & ~n52536;
  assign n52538 = ~n12773 & ~n52537;
  assign n52539 = ~n3281 & ~n52538;
  assign n52540 = ~n3281 & ~n52539;
  assign n52541 = n3378 & ~n52540;
  assign n52542 = ~n28139 & ~n40581;
  assign n52543 = controllable_nhgrant0 & ~n52542;
  assign n52544 = ~n12827 & ~n52543;
  assign n52545 = ~n3281 & ~n52544;
  assign n52546 = ~n3281 & ~n52545;
  assign n52547 = ~n3378 & ~n52546;
  assign n52548 = ~n52541 & ~n52547;
  assign n52549 = n3492 & ~n52548;
  assign n52550 = n3492 & ~n52549;
  assign n52551 = n3485 & ~n52550;
  assign n52552 = n3485 & ~n52551;
  assign n52553 = ~n3476 & ~n52552;
  assign n52554 = ~n28183 & ~n40616;
  assign n52555 = controllable_nhgrant0 & ~n52554;
  assign n52556 = ~n12942 & ~n52555;
  assign n52557 = ~n3281 & ~n52556;
  assign n52558 = ~n3281 & ~n52557;
  assign n52559 = n3378 & ~n52558;
  assign n52560 = ~n28235 & ~n40713;
  assign n52561 = controllable_nhgrant0 & ~n52560;
  assign n52562 = ~n13064 & ~n52561;
  assign n52563 = ~n3281 & ~n52562;
  assign n52564 = ~n3281 & ~n52563;
  assign n52565 = ~n3378 & ~n52564;
  assign n52566 = ~n52559 & ~n52565;
  assign n52567 = n3492 & ~n52566;
  assign n52568 = ~n27622 & ~n52567;
  assign n52569 = n3485 & ~n52568;
  assign n52570 = ~n27621 & ~n52569;
  assign n52571 = n3476 & ~n52570;
  assign n52572 = ~n52553 & ~n52571;
  assign n52573 = n3374 & ~n52572;
  assign n52574 = ~n52535 & ~n52573;
  assign n52575 = ~n3655 & ~n52574;
  assign n52576 = ~n52523 & ~n52575;
  assign n52577 = n3652 & ~n52576;
  assign n52578 = ~n28091 & ~n40743;
  assign n52579 = controllable_nhgrant0 & ~n52578;
  assign n52580 = ~n7118 & ~n52579;
  assign n52581 = ~n3281 & ~n52580;
  assign n52582 = ~n3281 & ~n52581;
  assign n52583 = ~n3378 & ~n52582;
  assign n52584 = ~n28079 & ~n52583;
  assign n52585 = n3492 & ~n52584;
  assign n52586 = n3492 & ~n52585;
  assign n52587 = n3485 & ~n52586;
  assign n52588 = n3485 & ~n52587;
  assign n52589 = ~n3374 & ~n52588;
  assign n52590 = ~n28116 & ~n40767;
  assign n52591 = controllable_nhgrant0 & ~n52590;
  assign n52592 = ~n12773 & ~n52591;
  assign n52593 = ~n3281 & ~n52592;
  assign n52594 = ~n3281 & ~n52593;
  assign n52595 = n3378 & ~n52594;
  assign n52596 = ~n28139 & ~n40795;
  assign n52597 = controllable_nhgrant0 & ~n52596;
  assign n52598 = ~n12827 & ~n52597;
  assign n52599 = ~n3281 & ~n52598;
  assign n52600 = ~n3281 & ~n52599;
  assign n52601 = ~n3378 & ~n52600;
  assign n52602 = ~n52595 & ~n52601;
  assign n52603 = n3492 & ~n52602;
  assign n52604 = n3492 & ~n52603;
  assign n52605 = n3485 & ~n52604;
  assign n52606 = n3485 & ~n52605;
  assign n52607 = ~n3476 & ~n52606;
  assign n52608 = ~n28183 & ~n40823;
  assign n52609 = controllable_nhgrant0 & ~n52608;
  assign n52610 = ~n12942 & ~n52609;
  assign n52611 = ~n3281 & ~n52610;
  assign n52612 = ~n3281 & ~n52611;
  assign n52613 = n3378 & ~n52612;
  assign n52614 = ~n28235 & ~n40881;
  assign n52615 = controllable_nhgrant0 & ~n52614;
  assign n52616 = ~n13064 & ~n52615;
  assign n52617 = ~n3281 & ~n52616;
  assign n52618 = ~n3281 & ~n52617;
  assign n52619 = ~n3378 & ~n52618;
  assign n52620 = ~n52613 & ~n52619;
  assign n52621 = n3492 & ~n52620;
  assign n52622 = ~n27622 & ~n52621;
  assign n52623 = n3485 & ~n52622;
  assign n52624 = ~n27621 & ~n52623;
  assign n52625 = n3476 & ~n52624;
  assign n52626 = ~n52607 & ~n52625;
  assign n52627 = n3374 & ~n52626;
  assign n52628 = ~n52589 & ~n52627;
  assign n52629 = n3655 & ~n52628;
  assign n52630 = ~n28091 & ~n40909;
  assign n52631 = controllable_nhgrant0 & ~n52630;
  assign n52632 = ~n7118 & ~n52631;
  assign n52633 = ~n3281 & ~n52632;
  assign n52634 = ~n3281 & ~n52633;
  assign n52635 = ~n3378 & ~n52634;
  assign n52636 = ~n28079 & ~n52635;
  assign n52637 = n3492 & ~n52636;
  assign n52638 = n3492 & ~n52637;
  assign n52639 = n3485 & ~n52638;
  assign n52640 = n3485 & ~n52639;
  assign n52641 = ~n3374 & ~n52640;
  assign n52642 = ~n28116 & ~n40933;
  assign n52643 = controllable_nhgrant0 & ~n52642;
  assign n52644 = ~n12773 & ~n52643;
  assign n52645 = ~n3281 & ~n52644;
  assign n52646 = ~n3281 & ~n52645;
  assign n52647 = n3378 & ~n52646;
  assign n52648 = ~n28139 & ~n40961;
  assign n52649 = controllable_nhgrant0 & ~n52648;
  assign n52650 = ~n12827 & ~n52649;
  assign n52651 = ~n3281 & ~n52650;
  assign n52652 = ~n3281 & ~n52651;
  assign n52653 = ~n3378 & ~n52652;
  assign n52654 = ~n52647 & ~n52653;
  assign n52655 = n3492 & ~n52654;
  assign n52656 = n3492 & ~n52655;
  assign n52657 = n3485 & ~n52656;
  assign n52658 = n3485 & ~n52657;
  assign n52659 = ~n3476 & ~n52658;
  assign n52660 = ~n28183 & ~n40989;
  assign n52661 = controllable_nhgrant0 & ~n52660;
  assign n52662 = ~n12942 & ~n52661;
  assign n52663 = ~n3281 & ~n52662;
  assign n52664 = ~n3281 & ~n52663;
  assign n52665 = n3378 & ~n52664;
  assign n52666 = ~n28235 & ~n41047;
  assign n52667 = controllable_nhgrant0 & ~n52666;
  assign n52668 = ~n13064 & ~n52667;
  assign n52669 = ~n3281 & ~n52668;
  assign n52670 = ~n3281 & ~n52669;
  assign n52671 = ~n3378 & ~n52670;
  assign n52672 = ~n52665 & ~n52671;
  assign n52673 = n3492 & ~n52672;
  assign n52674 = ~n27622 & ~n52673;
  assign n52675 = n3485 & ~n52674;
  assign n52676 = ~n27621 & ~n52675;
  assign n52677 = n3476 & ~n52676;
  assign n52678 = ~n52659 & ~n52677;
  assign n52679 = n3374 & ~n52678;
  assign n52680 = ~n52641 & ~n52679;
  assign n52681 = ~n3655 & ~n52680;
  assign n52682 = ~n52629 & ~n52681;
  assign n52683 = ~n3652 & ~n52682;
  assign n52684 = ~n52577 & ~n52683;
  assign n52685 = n3368 & ~n52684;
  assign n52686 = ~n52471 & ~n52685;
  assign n52687 = n3362 & ~n52686;
  assign n52688 = n3492 & ~n52238;
  assign n52689 = ~n3631 & ~n52688;
  assign n52690 = n3485 & ~n52689;
  assign n52691 = ~n3630 & ~n52690;
  assign n52692 = ~n3476 & ~n52691;
  assign n52693 = ~n28421 & ~n51148;
  assign n52694 = ~n3485 & ~n52693;
  assign n52695 = ~n27779 & ~n52688;
  assign n52696 = n3485 & ~n52695;
  assign n52697 = ~n52694 & ~n52696;
  assign n52698 = n3476 & ~n52697;
  assign n52699 = ~n52692 & ~n52698;
  assign n52700 = ~n3374 & ~n52699;
  assign n52701 = n3492 & ~n52262;
  assign n52702 = ~n3631 & ~n52701;
  assign n52703 = n3485 & ~n52702;
  assign n52704 = ~n3630 & ~n52703;
  assign n52705 = ~n3476 & ~n52704;
  assign n52706 = n3492 & ~n52280;
  assign n52707 = ~n27779 & ~n52706;
  assign n52708 = n3485 & ~n52707;
  assign n52709 = ~n52694 & ~n52708;
  assign n52710 = n3476 & ~n52709;
  assign n52711 = ~n52705 & ~n52710;
  assign n52712 = n3374 & ~n52711;
  assign n52713 = ~n52700 & ~n52712;
  assign n52714 = n3655 & ~n52713;
  assign n52715 = n3492 & ~n52296;
  assign n52716 = ~n3631 & ~n52715;
  assign n52717 = n3485 & ~n52716;
  assign n52718 = ~n3630 & ~n52717;
  assign n52719 = ~n3476 & ~n52718;
  assign n52720 = ~n28421 & ~n51191;
  assign n52721 = ~n3485 & ~n52720;
  assign n52722 = ~n27779 & ~n52715;
  assign n52723 = n3485 & ~n52722;
  assign n52724 = ~n52721 & ~n52723;
  assign n52725 = n3476 & ~n52724;
  assign n52726 = ~n52719 & ~n52725;
  assign n52727 = ~n3374 & ~n52726;
  assign n52728 = n3492 & ~n52320;
  assign n52729 = ~n3631 & ~n52728;
  assign n52730 = n3485 & ~n52729;
  assign n52731 = ~n3630 & ~n52730;
  assign n52732 = ~n3476 & ~n52731;
  assign n52733 = n3492 & ~n52338;
  assign n52734 = ~n27779 & ~n52733;
  assign n52735 = n3485 & ~n52734;
  assign n52736 = ~n52721 & ~n52735;
  assign n52737 = n3476 & ~n52736;
  assign n52738 = ~n52732 & ~n52737;
  assign n52739 = n3374 & ~n52738;
  assign n52740 = ~n52727 & ~n52739;
  assign n52741 = ~n3655 & ~n52740;
  assign n52742 = ~n52714 & ~n52741;
  assign n52743 = n3652 & ~n52742;
  assign n52744 = n3492 & ~n52356;
  assign n52745 = ~n3631 & ~n52744;
  assign n52746 = n3485 & ~n52745;
  assign n52747 = ~n3630 & ~n52746;
  assign n52748 = ~n3476 & ~n52747;
  assign n52749 = ~n28421 & ~n51236;
  assign n52750 = ~n3485 & ~n52749;
  assign n52751 = ~n27779 & ~n52744;
  assign n52752 = n3485 & ~n52751;
  assign n52753 = ~n52750 & ~n52752;
  assign n52754 = n3476 & ~n52753;
  assign n52755 = ~n52748 & ~n52754;
  assign n52756 = ~n3374 & ~n52755;
  assign n52757 = n3492 & ~n52380;
  assign n52758 = ~n3631 & ~n52757;
  assign n52759 = n3485 & ~n52758;
  assign n52760 = ~n3630 & ~n52759;
  assign n52761 = ~n3476 & ~n52760;
  assign n52762 = n3492 & ~n52398;
  assign n52763 = ~n27779 & ~n52762;
  assign n52764 = n3485 & ~n52763;
  assign n52765 = ~n52750 & ~n52764;
  assign n52766 = n3476 & ~n52765;
  assign n52767 = ~n52761 & ~n52766;
  assign n52768 = n3374 & ~n52767;
  assign n52769 = ~n52756 & ~n52768;
  assign n52770 = n3655 & ~n52769;
  assign n52771 = n3492 & ~n52414;
  assign n52772 = ~n3631 & ~n52771;
  assign n52773 = n3485 & ~n52772;
  assign n52774 = ~n3630 & ~n52773;
  assign n52775 = ~n3476 & ~n52774;
  assign n52776 = ~n28421 & ~n51279;
  assign n52777 = ~n3485 & ~n52776;
  assign n52778 = ~n27779 & ~n52771;
  assign n52779 = n3485 & ~n52778;
  assign n52780 = ~n52777 & ~n52779;
  assign n52781 = n3476 & ~n52780;
  assign n52782 = ~n52775 & ~n52781;
  assign n52783 = ~n3374 & ~n52782;
  assign n52784 = n3492 & ~n52438;
  assign n52785 = ~n3631 & ~n52784;
  assign n52786 = n3485 & ~n52785;
  assign n52787 = ~n3630 & ~n52786;
  assign n52788 = ~n3476 & ~n52787;
  assign n52789 = n3492 & ~n52456;
  assign n52790 = ~n27779 & ~n52789;
  assign n52791 = n3485 & ~n52790;
  assign n52792 = ~n52777 & ~n52791;
  assign n52793 = n3476 & ~n52792;
  assign n52794 = ~n52788 & ~n52793;
  assign n52795 = n3374 & ~n52794;
  assign n52796 = ~n52783 & ~n52795;
  assign n52797 = ~n3655 & ~n52796;
  assign n52798 = ~n52770 & ~n52797;
  assign n52799 = ~n3652 & ~n52798;
  assign n52800 = ~n52743 & ~n52799;
  assign n52801 = ~n3368 & ~n52800;
  assign n52802 = n3492 & ~n52476;
  assign n52803 = n3492 & ~n52802;
  assign n52804 = n3485 & ~n52803;
  assign n52805 = n3485 & ~n52804;
  assign n52806 = ~n3476 & ~n52805;
  assign n52807 = ~n8525 & ~n52804;
  assign n52808 = n3476 & ~n52807;
  assign n52809 = ~n52806 & ~n52808;
  assign n52810 = ~n3374 & ~n52809;
  assign n52811 = n3492 & ~n52494;
  assign n52812 = n3492 & ~n52811;
  assign n52813 = n3485 & ~n52812;
  assign n52814 = n3485 & ~n52813;
  assign n52815 = ~n3476 & ~n52814;
  assign n52816 = ~n28545 & ~n51321;
  assign n52817 = ~n3485 & ~n52816;
  assign n52818 = n3492 & ~n52512;
  assign n52819 = ~n27622 & ~n52818;
  assign n52820 = n3485 & ~n52819;
  assign n52821 = ~n52817 & ~n52820;
  assign n52822 = n3476 & ~n52821;
  assign n52823 = ~n52815 & ~n52822;
  assign n52824 = n3374 & ~n52823;
  assign n52825 = ~n52810 & ~n52824;
  assign n52826 = n3655 & ~n52825;
  assign n52827 = n3492 & ~n52528;
  assign n52828 = n3492 & ~n52827;
  assign n52829 = n3485 & ~n52828;
  assign n52830 = n3485 & ~n52829;
  assign n52831 = ~n3476 & ~n52830;
  assign n52832 = ~n8525 & ~n52829;
  assign n52833 = n3476 & ~n52832;
  assign n52834 = ~n52831 & ~n52833;
  assign n52835 = ~n3374 & ~n52834;
  assign n52836 = n3492 & ~n52546;
  assign n52837 = n3492 & ~n52836;
  assign n52838 = n3485 & ~n52837;
  assign n52839 = n3485 & ~n52838;
  assign n52840 = ~n3476 & ~n52839;
  assign n52841 = ~n28545 & ~n51348;
  assign n52842 = ~n3485 & ~n52841;
  assign n52843 = n3492 & ~n52564;
  assign n52844 = ~n27622 & ~n52843;
  assign n52845 = n3485 & ~n52844;
  assign n52846 = ~n52842 & ~n52845;
  assign n52847 = n3476 & ~n52846;
  assign n52848 = ~n52840 & ~n52847;
  assign n52849 = n3374 & ~n52848;
  assign n52850 = ~n52835 & ~n52849;
  assign n52851 = ~n3655 & ~n52850;
  assign n52852 = ~n52826 & ~n52851;
  assign n52853 = n3652 & ~n52852;
  assign n52854 = n3492 & ~n52582;
  assign n52855 = n3492 & ~n52854;
  assign n52856 = n3485 & ~n52855;
  assign n52857 = n3485 & ~n52856;
  assign n52858 = ~n3476 & ~n52857;
  assign n52859 = ~n8525 & ~n52856;
  assign n52860 = n3476 & ~n52859;
  assign n52861 = ~n52858 & ~n52860;
  assign n52862 = ~n3374 & ~n52861;
  assign n52863 = n3492 & ~n52600;
  assign n52864 = n3492 & ~n52863;
  assign n52865 = n3485 & ~n52864;
  assign n52866 = n3485 & ~n52865;
  assign n52867 = ~n3476 & ~n52866;
  assign n52868 = ~n28545 & ~n51377;
  assign n52869 = ~n3485 & ~n52868;
  assign n52870 = n3492 & ~n52618;
  assign n52871 = ~n27622 & ~n52870;
  assign n52872 = n3485 & ~n52871;
  assign n52873 = ~n52869 & ~n52872;
  assign n52874 = n3476 & ~n52873;
  assign n52875 = ~n52867 & ~n52874;
  assign n52876 = n3374 & ~n52875;
  assign n52877 = ~n52862 & ~n52876;
  assign n52878 = n3655 & ~n52877;
  assign n52879 = n3492 & ~n52634;
  assign n52880 = n3492 & ~n52879;
  assign n52881 = n3485 & ~n52880;
  assign n52882 = n3485 & ~n52881;
  assign n52883 = ~n3476 & ~n52882;
  assign n52884 = ~n8525 & ~n52881;
  assign n52885 = n3476 & ~n52884;
  assign n52886 = ~n52883 & ~n52885;
  assign n52887 = ~n3374 & ~n52886;
  assign n52888 = n3492 & ~n52652;
  assign n52889 = n3492 & ~n52888;
  assign n52890 = n3485 & ~n52889;
  assign n52891 = n3485 & ~n52890;
  assign n52892 = ~n3476 & ~n52891;
  assign n52893 = ~n28545 & ~n51404;
  assign n52894 = ~n3485 & ~n52893;
  assign n52895 = n3492 & ~n52670;
  assign n52896 = ~n27622 & ~n52895;
  assign n52897 = n3485 & ~n52896;
  assign n52898 = ~n52894 & ~n52897;
  assign n52899 = n3476 & ~n52898;
  assign n52900 = ~n52892 & ~n52899;
  assign n52901 = n3374 & ~n52900;
  assign n52902 = ~n52887 & ~n52901;
  assign n52903 = ~n3655 & ~n52902;
  assign n52904 = ~n52878 & ~n52903;
  assign n52905 = ~n3652 & ~n52904;
  assign n52906 = ~n52853 & ~n52905;
  assign n52907 = n3368 & ~n52906;
  assign n52908 = ~n52801 & ~n52907;
  assign n52909 = ~n3362 & ~n52908;
  assign n52910 = ~n52687 & ~n52909;
  assign n52911 = n3359 & ~n52910;
  assign n52912 = ~n51424 & ~n52696;
  assign n52913 = n3476 & ~n52912;
  assign n52914 = ~n52692 & ~n52913;
  assign n52915 = ~n3374 & ~n52914;
  assign n52916 = ~n51424 & ~n52708;
  assign n52917 = n3476 & ~n52916;
  assign n52918 = ~n52705 & ~n52917;
  assign n52919 = n3374 & ~n52918;
  assign n52920 = ~n52915 & ~n52919;
  assign n52921 = n3655 & ~n52920;
  assign n52922 = ~n51435 & ~n52723;
  assign n52923 = n3476 & ~n52922;
  assign n52924 = ~n52719 & ~n52923;
  assign n52925 = ~n3374 & ~n52924;
  assign n52926 = ~n51435 & ~n52735;
  assign n52927 = n3476 & ~n52926;
  assign n52928 = ~n52732 & ~n52927;
  assign n52929 = n3374 & ~n52928;
  assign n52930 = ~n52925 & ~n52929;
  assign n52931 = ~n3655 & ~n52930;
  assign n52932 = ~n52921 & ~n52931;
  assign n52933 = n3652 & ~n52932;
  assign n52934 = ~n51448 & ~n52752;
  assign n52935 = n3476 & ~n52934;
  assign n52936 = ~n52748 & ~n52935;
  assign n52937 = ~n3374 & ~n52936;
  assign n52938 = ~n51448 & ~n52764;
  assign n52939 = n3476 & ~n52938;
  assign n52940 = ~n52761 & ~n52939;
  assign n52941 = n3374 & ~n52940;
  assign n52942 = ~n52937 & ~n52941;
  assign n52943 = n3655 & ~n52942;
  assign n52944 = ~n51459 & ~n52779;
  assign n52945 = n3476 & ~n52944;
  assign n52946 = ~n52775 & ~n52945;
  assign n52947 = ~n3374 & ~n52946;
  assign n52948 = ~n51459 & ~n52791;
  assign n52949 = n3476 & ~n52948;
  assign n52950 = ~n52788 & ~n52949;
  assign n52951 = n3374 & ~n52950;
  assign n52952 = ~n52947 & ~n52951;
  assign n52953 = ~n3655 & ~n52952;
  assign n52954 = ~n52943 & ~n52953;
  assign n52955 = ~n3652 & ~n52954;
  assign n52956 = ~n52933 & ~n52955;
  assign n52957 = ~n3368 & ~n52956;
  assign n52958 = ~n8689 & ~n52804;
  assign n52959 = n3476 & ~n52958;
  assign n52960 = ~n52806 & ~n52959;
  assign n52961 = ~n3374 & ~n52960;
  assign n52962 = ~n51478 & ~n52820;
  assign n52963 = n3476 & ~n52962;
  assign n52964 = ~n52815 & ~n52963;
  assign n52965 = n3374 & ~n52964;
  assign n52966 = ~n52961 & ~n52965;
  assign n52967 = n3655 & ~n52966;
  assign n52968 = ~n8689 & ~n52829;
  assign n52969 = n3476 & ~n52968;
  assign n52970 = ~n52831 & ~n52969;
  assign n52971 = ~n3374 & ~n52970;
  assign n52972 = ~n51489 & ~n52845;
  assign n52973 = n3476 & ~n52972;
  assign n52974 = ~n52840 & ~n52973;
  assign n52975 = n3374 & ~n52974;
  assign n52976 = ~n52971 & ~n52975;
  assign n52977 = ~n3655 & ~n52976;
  assign n52978 = ~n52967 & ~n52977;
  assign n52979 = n3652 & ~n52978;
  assign n52980 = ~n8689 & ~n52856;
  assign n52981 = n3476 & ~n52980;
  assign n52982 = ~n52858 & ~n52981;
  assign n52983 = ~n3374 & ~n52982;
  assign n52984 = ~n51502 & ~n52872;
  assign n52985 = n3476 & ~n52984;
  assign n52986 = ~n52867 & ~n52985;
  assign n52987 = n3374 & ~n52986;
  assign n52988 = ~n52983 & ~n52987;
  assign n52989 = n3655 & ~n52988;
  assign n52990 = ~n8689 & ~n52881;
  assign n52991 = n3476 & ~n52990;
  assign n52992 = ~n52883 & ~n52991;
  assign n52993 = ~n3374 & ~n52992;
  assign n52994 = ~n51513 & ~n52897;
  assign n52995 = n3476 & ~n52994;
  assign n52996 = ~n52892 & ~n52995;
  assign n52997 = n3374 & ~n52996;
  assign n52998 = ~n52993 & ~n52997;
  assign n52999 = ~n3655 & ~n52998;
  assign n53000 = ~n52989 & ~n52999;
  assign n53001 = ~n3652 & ~n53000;
  assign n53002 = ~n52979 & ~n53001;
  assign n53003 = n3368 & ~n53002;
  assign n53004 = ~n52957 & ~n53003;
  assign n53005 = n3362 & ~n53004;
  assign n53006 = n3378 & ~n52238;
  assign n53007 = ~n51532 & ~n53006;
  assign n53008 = n3492 & ~n53007;
  assign n53009 = ~n3631 & ~n53008;
  assign n53010 = n3485 & ~n53009;
  assign n53011 = ~n3630 & ~n53010;
  assign n53012 = ~n3476 & ~n53011;
  assign n53013 = ~n51148 & ~n53008;
  assign n53014 = n3485 & ~n53013;
  assign n53015 = ~n51424 & ~n53014;
  assign n53016 = n3476 & ~n53015;
  assign n53017 = ~n53012 & ~n53016;
  assign n53018 = ~n3374 & ~n53017;
  assign n53019 = n3378 & ~n52262;
  assign n53020 = ~n51551 & ~n53019;
  assign n53021 = n3492 & ~n53020;
  assign n53022 = ~n3631 & ~n53021;
  assign n53023 = n3485 & ~n53022;
  assign n53024 = ~n3630 & ~n53023;
  assign n53025 = ~n3476 & ~n53024;
  assign n53026 = n3378 & ~n52280;
  assign n53027 = ~n51564 & ~n53026;
  assign n53028 = n3492 & ~n53027;
  assign n53029 = ~n51148 & ~n53028;
  assign n53030 = n3485 & ~n53029;
  assign n53031 = ~n51424 & ~n53030;
  assign n53032 = n3476 & ~n53031;
  assign n53033 = ~n53025 & ~n53032;
  assign n53034 = n3374 & ~n53033;
  assign n53035 = ~n53018 & ~n53034;
  assign n53036 = n3655 & ~n53035;
  assign n53037 = n3378 & ~n52296;
  assign n53038 = ~n51581 & ~n53037;
  assign n53039 = n3492 & ~n53038;
  assign n53040 = ~n3631 & ~n53039;
  assign n53041 = n3485 & ~n53040;
  assign n53042 = ~n3630 & ~n53041;
  assign n53043 = ~n3476 & ~n53042;
  assign n53044 = ~n51191 & ~n53039;
  assign n53045 = n3485 & ~n53044;
  assign n53046 = ~n51435 & ~n53045;
  assign n53047 = n3476 & ~n53046;
  assign n53048 = ~n53043 & ~n53047;
  assign n53049 = ~n3374 & ~n53048;
  assign n53050 = n3378 & ~n52320;
  assign n53051 = ~n51600 & ~n53050;
  assign n53052 = n3492 & ~n53051;
  assign n53053 = ~n3631 & ~n53052;
  assign n53054 = n3485 & ~n53053;
  assign n53055 = ~n3630 & ~n53054;
  assign n53056 = ~n3476 & ~n53055;
  assign n53057 = n3378 & ~n52338;
  assign n53058 = ~n51613 & ~n53057;
  assign n53059 = n3492 & ~n53058;
  assign n53060 = ~n51191 & ~n53059;
  assign n53061 = n3485 & ~n53060;
  assign n53062 = ~n51435 & ~n53061;
  assign n53063 = n3476 & ~n53062;
  assign n53064 = ~n53056 & ~n53063;
  assign n53065 = n3374 & ~n53064;
  assign n53066 = ~n53049 & ~n53065;
  assign n53067 = ~n3655 & ~n53066;
  assign n53068 = ~n53036 & ~n53067;
  assign n53069 = n3652 & ~n53068;
  assign n53070 = n3378 & ~n52356;
  assign n53071 = ~n51632 & ~n53070;
  assign n53072 = n3492 & ~n53071;
  assign n53073 = ~n3631 & ~n53072;
  assign n53074 = n3485 & ~n53073;
  assign n53075 = ~n3630 & ~n53074;
  assign n53076 = ~n3476 & ~n53075;
  assign n53077 = ~n51236 & ~n53072;
  assign n53078 = n3485 & ~n53077;
  assign n53079 = ~n51448 & ~n53078;
  assign n53080 = n3476 & ~n53079;
  assign n53081 = ~n53076 & ~n53080;
  assign n53082 = ~n3374 & ~n53081;
  assign n53083 = n3378 & ~n52380;
  assign n53084 = ~n51651 & ~n53083;
  assign n53085 = n3492 & ~n53084;
  assign n53086 = ~n3631 & ~n53085;
  assign n53087 = n3485 & ~n53086;
  assign n53088 = ~n3630 & ~n53087;
  assign n53089 = ~n3476 & ~n53088;
  assign n53090 = n3378 & ~n52398;
  assign n53091 = ~n51664 & ~n53090;
  assign n53092 = n3492 & ~n53091;
  assign n53093 = ~n51236 & ~n53092;
  assign n53094 = n3485 & ~n53093;
  assign n53095 = ~n51448 & ~n53094;
  assign n53096 = n3476 & ~n53095;
  assign n53097 = ~n53089 & ~n53096;
  assign n53098 = n3374 & ~n53097;
  assign n53099 = ~n53082 & ~n53098;
  assign n53100 = n3655 & ~n53099;
  assign n53101 = n3378 & ~n52414;
  assign n53102 = ~n51681 & ~n53101;
  assign n53103 = n3492 & ~n53102;
  assign n53104 = ~n3631 & ~n53103;
  assign n53105 = n3485 & ~n53104;
  assign n53106 = ~n3630 & ~n53105;
  assign n53107 = ~n3476 & ~n53106;
  assign n53108 = ~n51279 & ~n53103;
  assign n53109 = n3485 & ~n53108;
  assign n53110 = ~n51459 & ~n53109;
  assign n53111 = n3476 & ~n53110;
  assign n53112 = ~n53107 & ~n53111;
  assign n53113 = ~n3374 & ~n53112;
  assign n53114 = n3378 & ~n52438;
  assign n53115 = ~n51700 & ~n53114;
  assign n53116 = n3492 & ~n53115;
  assign n53117 = ~n3631 & ~n53116;
  assign n53118 = n3485 & ~n53117;
  assign n53119 = ~n3630 & ~n53118;
  assign n53120 = ~n3476 & ~n53119;
  assign n53121 = n3378 & ~n52456;
  assign n53122 = ~n51713 & ~n53121;
  assign n53123 = n3492 & ~n53122;
  assign n53124 = ~n51279 & ~n53123;
  assign n53125 = n3485 & ~n53124;
  assign n53126 = ~n51459 & ~n53125;
  assign n53127 = n3476 & ~n53126;
  assign n53128 = ~n53120 & ~n53127;
  assign n53129 = n3374 & ~n53128;
  assign n53130 = ~n53113 & ~n53129;
  assign n53131 = ~n3655 & ~n53130;
  assign n53132 = ~n53100 & ~n53131;
  assign n53133 = ~n3652 & ~n53132;
  assign n53134 = ~n53069 & ~n53133;
  assign n53135 = ~n3368 & ~n53134;
  assign n53136 = n3378 & ~n52476;
  assign n53137 = ~n51734 & ~n53136;
  assign n53138 = n3492 & ~n53137;
  assign n53139 = n3492 & ~n53138;
  assign n53140 = n3485 & ~n53139;
  assign n53141 = n3485 & ~n53140;
  assign n53142 = ~n3476 & ~n53141;
  assign n53143 = ~n8523 & ~n53138;
  assign n53144 = n3485 & ~n53143;
  assign n53145 = ~n8689 & ~n53144;
  assign n53146 = n3476 & ~n53145;
  assign n53147 = ~n53142 & ~n53146;
  assign n53148 = ~n3374 & ~n53147;
  assign n53149 = n3378 & ~n52494;
  assign n53150 = ~n51753 & ~n53149;
  assign n53151 = n3492 & ~n53150;
  assign n53152 = n3492 & ~n53151;
  assign n53153 = n3485 & ~n53152;
  assign n53154 = n3485 & ~n53153;
  assign n53155 = ~n3476 & ~n53154;
  assign n53156 = ~n28235 & ~n41649;
  assign n53157 = controllable_nhgrant0 & ~n53156;
  assign n53158 = ~n13845 & ~n53157;
  assign n53159 = ~n3281 & ~n53158;
  assign n53160 = ~n3281 & ~n53159;
  assign n53161 = n3378 & ~n53160;
  assign n53162 = ~n51771 & ~n53161;
  assign n53163 = n3492 & ~n53162;
  assign n53164 = ~n51321 & ~n53163;
  assign n53165 = n3485 & ~n53164;
  assign n53166 = ~n51478 & ~n53165;
  assign n53167 = n3476 & ~n53166;
  assign n53168 = ~n53155 & ~n53167;
  assign n53169 = n3374 & ~n53168;
  assign n53170 = ~n53148 & ~n53169;
  assign n53171 = n3655 & ~n53170;
  assign n53172 = n3378 & ~n52528;
  assign n53173 = ~n51788 & ~n53172;
  assign n53174 = n3492 & ~n53173;
  assign n53175 = n3492 & ~n53174;
  assign n53176 = n3485 & ~n53175;
  assign n53177 = n3485 & ~n53176;
  assign n53178 = ~n3476 & ~n53177;
  assign n53179 = ~n8523 & ~n53174;
  assign n53180 = n3485 & ~n53179;
  assign n53181 = ~n8689 & ~n53180;
  assign n53182 = n3476 & ~n53181;
  assign n53183 = ~n53178 & ~n53182;
  assign n53184 = ~n3374 & ~n53183;
  assign n53185 = n3378 & ~n52546;
  assign n53186 = ~n51807 & ~n53185;
  assign n53187 = n3492 & ~n53186;
  assign n53188 = n3492 & ~n53187;
  assign n53189 = n3485 & ~n53188;
  assign n53190 = n3485 & ~n53189;
  assign n53191 = ~n3476 & ~n53190;
  assign n53192 = ~n28235 & ~n41771;
  assign n53193 = controllable_nhgrant0 & ~n53192;
  assign n53194 = ~n13845 & ~n53193;
  assign n53195 = ~n3281 & ~n53194;
  assign n53196 = ~n3281 & ~n53195;
  assign n53197 = n3378 & ~n53196;
  assign n53198 = ~n51825 & ~n53197;
  assign n53199 = n3492 & ~n53198;
  assign n53200 = ~n51348 & ~n53199;
  assign n53201 = n3485 & ~n53200;
  assign n53202 = ~n51489 & ~n53201;
  assign n53203 = n3476 & ~n53202;
  assign n53204 = ~n53191 & ~n53203;
  assign n53205 = n3374 & ~n53204;
  assign n53206 = ~n53184 & ~n53205;
  assign n53207 = ~n3655 & ~n53206;
  assign n53208 = ~n53171 & ~n53207;
  assign n53209 = n3652 & ~n53208;
  assign n53210 = n3378 & ~n52582;
  assign n53211 = ~n51844 & ~n53210;
  assign n53212 = n3492 & ~n53211;
  assign n53213 = n3492 & ~n53212;
  assign n53214 = n3485 & ~n53213;
  assign n53215 = n3485 & ~n53214;
  assign n53216 = ~n3476 & ~n53215;
  assign n53217 = ~n8523 & ~n53212;
  assign n53218 = n3485 & ~n53217;
  assign n53219 = ~n8689 & ~n53218;
  assign n53220 = n3476 & ~n53219;
  assign n53221 = ~n53216 & ~n53220;
  assign n53222 = ~n3374 & ~n53221;
  assign n53223 = n3378 & ~n52600;
  assign n53224 = ~n51863 & ~n53223;
  assign n53225 = n3492 & ~n53224;
  assign n53226 = n3492 & ~n53225;
  assign n53227 = n3485 & ~n53226;
  assign n53228 = n3485 & ~n53227;
  assign n53229 = ~n3476 & ~n53228;
  assign n53230 = ~n28235 & ~n41859;
  assign n53231 = controllable_nhgrant0 & ~n53230;
  assign n53232 = ~n13845 & ~n53231;
  assign n53233 = ~n3281 & ~n53232;
  assign n53234 = ~n3281 & ~n53233;
  assign n53235 = n3378 & ~n53234;
  assign n53236 = ~n51881 & ~n53235;
  assign n53237 = n3492 & ~n53236;
  assign n53238 = ~n51377 & ~n53237;
  assign n53239 = n3485 & ~n53238;
  assign n53240 = ~n51502 & ~n53239;
  assign n53241 = n3476 & ~n53240;
  assign n53242 = ~n53229 & ~n53241;
  assign n53243 = n3374 & ~n53242;
  assign n53244 = ~n53222 & ~n53243;
  assign n53245 = n3655 & ~n53244;
  assign n53246 = n3378 & ~n52634;
  assign n53247 = ~n51898 & ~n53246;
  assign n53248 = n3492 & ~n53247;
  assign n53249 = n3492 & ~n53248;
  assign n53250 = n3485 & ~n53249;
  assign n53251 = n3485 & ~n53250;
  assign n53252 = ~n3476 & ~n53251;
  assign n53253 = ~n8523 & ~n53248;
  assign n53254 = n3485 & ~n53253;
  assign n53255 = ~n8689 & ~n53254;
  assign n53256 = n3476 & ~n53255;
  assign n53257 = ~n53252 & ~n53256;
  assign n53258 = ~n3374 & ~n53257;
  assign n53259 = n3378 & ~n52652;
  assign n53260 = ~n51917 & ~n53259;
  assign n53261 = n3492 & ~n53260;
  assign n53262 = n3492 & ~n53261;
  assign n53263 = n3485 & ~n53262;
  assign n53264 = n3485 & ~n53263;
  assign n53265 = ~n3476 & ~n53264;
  assign n53266 = ~n28235 & ~n41945;
  assign n53267 = controllable_nhgrant0 & ~n53266;
  assign n53268 = ~n13845 & ~n53267;
  assign n53269 = ~n3281 & ~n53268;
  assign n53270 = ~n3281 & ~n53269;
  assign n53271 = n3378 & ~n53270;
  assign n53272 = ~n51935 & ~n53271;
  assign n53273 = n3492 & ~n53272;
  assign n53274 = ~n51404 & ~n53273;
  assign n53275 = n3485 & ~n53274;
  assign n53276 = ~n51513 & ~n53275;
  assign n53277 = n3476 & ~n53276;
  assign n53278 = ~n53265 & ~n53277;
  assign n53279 = n3374 & ~n53278;
  assign n53280 = ~n53258 & ~n53279;
  assign n53281 = ~n3655 & ~n53280;
  assign n53282 = ~n53245 & ~n53281;
  assign n53283 = ~n3652 & ~n53282;
  assign n53284 = ~n53209 & ~n53283;
  assign n53285 = n3368 & ~n53284;
  assign n53286 = ~n53135 & ~n53285;
  assign n53287 = ~n3362 & ~n53286;
  assign n53288 = ~n53005 & ~n53287;
  assign n53289 = ~n3359 & ~n53288;
  assign n53290 = ~n52911 & ~n53289;
  assign n53291 = ~n3356 & ~n53290;
  assign n53292 = ~n52233 & ~n53291;
  assign n53293 = ~n3345 & ~n53292;
  assign n53294 = ~n29024 & ~n41985;
  assign n53295 = controllable_nhgrant0 & ~n53294;
  assign n53296 = ~n14166 & ~n53295;
  assign n53297 = ~n3281 & ~n53296;
  assign n53298 = ~n3281 & ~n53297;
  assign n53299 = n3378 & ~n53298;
  assign n53300 = ~n29031 & ~n41993;
  assign n53301 = controllable_nhgrant0 & ~n53300;
  assign n53302 = ~n14180 & ~n53301;
  assign n53303 = ~n3281 & ~n53302;
  assign n53304 = ~n3950 & ~n53303;
  assign n53305 = ~n3378 & ~n53304;
  assign n53306 = ~n53299 & ~n53305;
  assign n53307 = n3492 & ~n53306;
  assign n53308 = ~n3493 & ~n53307;
  assign n53309 = n3485 & ~n53308;
  assign n53310 = ~n3486 & ~n53309;
  assign n53311 = ~n3476 & ~n53310;
  assign n53312 = ~n29024 & ~n42021;
  assign n53313 = controllable_nhgrant0 & ~n53312;
  assign n53314 = ~n14166 & ~n53313;
  assign n53315 = ~n3281 & ~n53314;
  assign n53316 = ~n3281 & ~n53315;
  assign n53317 = n3378 & ~n53316;
  assign n53318 = ~n29031 & ~n42043;
  assign n53319 = controllable_nhgrant0 & ~n53318;
  assign n53320 = ~n14180 & ~n53319;
  assign n53321 = ~n3281 & ~n53320;
  assign n53322 = ~n4089 & ~n53321;
  assign n53323 = ~n3378 & ~n53322;
  assign n53324 = ~n53317 & ~n53323;
  assign n53325 = n3492 & ~n53324;
  assign n53326 = ~n3493 & ~n53325;
  assign n53327 = n3485 & ~n53326;
  assign n53328 = ~n3486 & ~n53327;
  assign n53329 = n3476 & ~n53328;
  assign n53330 = ~n53311 & ~n53329;
  assign n53331 = n3374 & ~n53330;
  assign n53332 = ~n14130 & ~n53331;
  assign n53333 = n3655 & ~n53332;
  assign n53334 = ~n29024 & ~n42071;
  assign n53335 = controllable_nhgrant0 & ~n53334;
  assign n53336 = ~n14166 & ~n53335;
  assign n53337 = ~n3281 & ~n53336;
  assign n53338 = ~n3281 & ~n53337;
  assign n53339 = n3378 & ~n53338;
  assign n53340 = ~n29031 & ~n42079;
  assign n53341 = controllable_nhgrant0 & ~n53340;
  assign n53342 = ~n14180 & ~n53341;
  assign n53343 = ~n3281 & ~n53342;
  assign n53344 = ~n3950 & ~n53343;
  assign n53345 = ~n3378 & ~n53344;
  assign n53346 = ~n53339 & ~n53345;
  assign n53347 = n3492 & ~n53346;
  assign n53348 = ~n3493 & ~n53347;
  assign n53349 = n3485 & ~n53348;
  assign n53350 = ~n3486 & ~n53349;
  assign n53351 = ~n3476 & ~n53350;
  assign n53352 = ~n29024 & ~n42107;
  assign n53353 = controllable_nhgrant0 & ~n53352;
  assign n53354 = ~n14166 & ~n53353;
  assign n53355 = ~n3281 & ~n53354;
  assign n53356 = ~n3281 & ~n53355;
  assign n53357 = n3378 & ~n53356;
  assign n53358 = ~n29031 & ~n42129;
  assign n53359 = controllable_nhgrant0 & ~n53358;
  assign n53360 = ~n14180 & ~n53359;
  assign n53361 = ~n3281 & ~n53360;
  assign n53362 = ~n4089 & ~n53361;
  assign n53363 = ~n3378 & ~n53362;
  assign n53364 = ~n53357 & ~n53363;
  assign n53365 = n3492 & ~n53364;
  assign n53366 = ~n3493 & ~n53365;
  assign n53367 = n3485 & ~n53366;
  assign n53368 = ~n3486 & ~n53367;
  assign n53369 = n3476 & ~n53368;
  assign n53370 = ~n53351 & ~n53369;
  assign n53371 = n3374 & ~n53370;
  assign n53372 = ~n14130 & ~n53371;
  assign n53373 = ~n3655 & ~n53372;
  assign n53374 = ~n53333 & ~n53373;
  assign n53375 = n3652 & ~n53374;
  assign n53376 = ~n29024 & ~n42159;
  assign n53377 = controllable_nhgrant0 & ~n53376;
  assign n53378 = ~n14166 & ~n53377;
  assign n53379 = ~n3281 & ~n53378;
  assign n53380 = ~n3281 & ~n53379;
  assign n53381 = n3378 & ~n53380;
  assign n53382 = ~n29031 & ~n42167;
  assign n53383 = controllable_nhgrant0 & ~n53382;
  assign n53384 = ~n14180 & ~n53383;
  assign n53385 = ~n3281 & ~n53384;
  assign n53386 = ~n3950 & ~n53385;
  assign n53387 = ~n3378 & ~n53386;
  assign n53388 = ~n53381 & ~n53387;
  assign n53389 = n3492 & ~n53388;
  assign n53390 = ~n3493 & ~n53389;
  assign n53391 = n3485 & ~n53390;
  assign n53392 = ~n3486 & ~n53391;
  assign n53393 = ~n3476 & ~n53392;
  assign n53394 = ~n29024 & ~n42195;
  assign n53395 = controllable_nhgrant0 & ~n53394;
  assign n53396 = ~n14166 & ~n53395;
  assign n53397 = ~n3281 & ~n53396;
  assign n53398 = ~n3281 & ~n53397;
  assign n53399 = n3378 & ~n53398;
  assign n53400 = ~n29031 & ~n42217;
  assign n53401 = controllable_nhgrant0 & ~n53400;
  assign n53402 = ~n14180 & ~n53401;
  assign n53403 = ~n3281 & ~n53402;
  assign n53404 = ~n4089 & ~n53403;
  assign n53405 = ~n3378 & ~n53404;
  assign n53406 = ~n53399 & ~n53405;
  assign n53407 = n3492 & ~n53406;
  assign n53408 = ~n14433 & ~n53407;
  assign n53409 = n3485 & ~n53408;
  assign n53410 = ~n14432 & ~n53409;
  assign n53411 = n3476 & ~n53410;
  assign n53412 = ~n53393 & ~n53411;
  assign n53413 = n3374 & ~n53412;
  assign n53414 = ~n14439 & ~n53413;
  assign n53415 = n3655 & ~n53414;
  assign n53416 = ~n29024 & ~n42245;
  assign n53417 = controllable_nhgrant0 & ~n53416;
  assign n53418 = ~n14166 & ~n53417;
  assign n53419 = ~n3281 & ~n53418;
  assign n53420 = ~n3281 & ~n53419;
  assign n53421 = n3378 & ~n53420;
  assign n53422 = ~n29031 & ~n42253;
  assign n53423 = controllable_nhgrant0 & ~n53422;
  assign n53424 = ~n14180 & ~n53423;
  assign n53425 = ~n3281 & ~n53424;
  assign n53426 = ~n3950 & ~n53425;
  assign n53427 = ~n3378 & ~n53426;
  assign n53428 = ~n53421 & ~n53427;
  assign n53429 = n3492 & ~n53428;
  assign n53430 = ~n3493 & ~n53429;
  assign n53431 = n3485 & ~n53430;
  assign n53432 = ~n3486 & ~n53431;
  assign n53433 = ~n3476 & ~n53432;
  assign n53434 = ~n29024 & ~n42281;
  assign n53435 = controllable_nhgrant0 & ~n53434;
  assign n53436 = ~n14166 & ~n53435;
  assign n53437 = ~n3281 & ~n53436;
  assign n53438 = ~n3281 & ~n53437;
  assign n53439 = n3378 & ~n53438;
  assign n53440 = ~n29031 & ~n42303;
  assign n53441 = controllable_nhgrant0 & ~n53440;
  assign n53442 = ~n14180 & ~n53441;
  assign n53443 = ~n3281 & ~n53442;
  assign n53444 = ~n4089 & ~n53443;
  assign n53445 = ~n3378 & ~n53444;
  assign n53446 = ~n53439 & ~n53445;
  assign n53447 = n3492 & ~n53446;
  assign n53448 = ~n14433 & ~n53447;
  assign n53449 = n3485 & ~n53448;
  assign n53450 = ~n14432 & ~n53449;
  assign n53451 = n3476 & ~n53450;
  assign n53452 = ~n53433 & ~n53451;
  assign n53453 = n3374 & ~n53452;
  assign n53454 = ~n14439 & ~n53453;
  assign n53455 = ~n3655 & ~n53454;
  assign n53456 = ~n53415 & ~n53455;
  assign n53457 = ~n3652 & ~n53456;
  assign n53458 = ~n53375 & ~n53457;
  assign n53459 = ~n3368 & ~n53458;
  assign n53460 = ~n29192 & ~n42335;
  assign n53461 = controllable_nhgrant0 & ~n53460;
  assign n53462 = ~n14725 & ~n53461;
  assign n53463 = ~n3281 & ~n53462;
  assign n53464 = ~n3281 & ~n53463;
  assign n53465 = n3492 & ~n53464;
  assign n53466 = n3492 & ~n53465;
  assign n53467 = n3485 & ~n53466;
  assign n53468 = n3485 & ~n53467;
  assign n53469 = ~n3476 & ~n53468;
  assign n53470 = ~n29192 & ~n42361;
  assign n53471 = controllable_nhgrant0 & ~n53470;
  assign n53472 = ~n14725 & ~n53471;
  assign n53473 = ~n3281 & ~n53472;
  assign n53474 = ~n3281 & ~n53473;
  assign n53475 = n3492 & ~n53474;
  assign n53476 = n3492 & ~n53475;
  assign n53477 = n3485 & ~n53476;
  assign n53478 = n3485 & ~n53477;
  assign n53479 = n3476 & ~n53478;
  assign n53480 = ~n53469 & ~n53479;
  assign n53481 = n3374 & ~n53480;
  assign n53482 = n3374 & ~n53481;
  assign n53483 = n3655 & ~n53482;
  assign n53484 = ~n29192 & ~n42387;
  assign n53485 = controllable_nhgrant0 & ~n53484;
  assign n53486 = ~n14725 & ~n53485;
  assign n53487 = ~n3281 & ~n53486;
  assign n53488 = ~n3281 & ~n53487;
  assign n53489 = n3492 & ~n53488;
  assign n53490 = n3492 & ~n53489;
  assign n53491 = n3485 & ~n53490;
  assign n53492 = n3485 & ~n53491;
  assign n53493 = ~n3476 & ~n53492;
  assign n53494 = ~n29192 & ~n42413;
  assign n53495 = controllable_nhgrant0 & ~n53494;
  assign n53496 = ~n14725 & ~n53495;
  assign n53497 = ~n3281 & ~n53496;
  assign n53498 = ~n3281 & ~n53497;
  assign n53499 = n3492 & ~n53498;
  assign n53500 = n3492 & ~n53499;
  assign n53501 = n3485 & ~n53500;
  assign n53502 = n3485 & ~n53501;
  assign n53503 = n3476 & ~n53502;
  assign n53504 = ~n53493 & ~n53503;
  assign n53505 = n3374 & ~n53504;
  assign n53506 = n3374 & ~n53505;
  assign n53507 = ~n3655 & ~n53506;
  assign n53508 = ~n53483 & ~n53507;
  assign n53509 = n3652 & ~n53508;
  assign n53510 = ~n29192 & ~n42441;
  assign n53511 = controllable_nhgrant0 & ~n53510;
  assign n53512 = ~n14725 & ~n53511;
  assign n53513 = ~n3281 & ~n53512;
  assign n53514 = ~n3281 & ~n53513;
  assign n53515 = n3492 & ~n53514;
  assign n53516 = n3492 & ~n53515;
  assign n53517 = n3485 & ~n53516;
  assign n53518 = n3485 & ~n53517;
  assign n53519 = ~n3476 & ~n53518;
  assign n53520 = ~n29192 & ~n42467;
  assign n53521 = controllable_nhgrant0 & ~n53520;
  assign n53522 = ~n14725 & ~n53521;
  assign n53523 = ~n3281 & ~n53522;
  assign n53524 = ~n3281 & ~n53523;
  assign n53525 = n3492 & ~n53524;
  assign n53526 = ~n14836 & ~n53525;
  assign n53527 = n3485 & ~n53526;
  assign n53528 = ~n14835 & ~n53527;
  assign n53529 = n3476 & ~n53528;
  assign n53530 = ~n53519 & ~n53529;
  assign n53531 = n3374 & ~n53530;
  assign n53532 = n3374 & ~n53531;
  assign n53533 = n3655 & ~n53532;
  assign n53534 = ~n29192 & ~n42493;
  assign n53535 = controllable_nhgrant0 & ~n53534;
  assign n53536 = ~n14725 & ~n53535;
  assign n53537 = ~n3281 & ~n53536;
  assign n53538 = ~n3281 & ~n53537;
  assign n53539 = n3492 & ~n53538;
  assign n53540 = n3492 & ~n53539;
  assign n53541 = n3485 & ~n53540;
  assign n53542 = n3485 & ~n53541;
  assign n53543 = ~n3476 & ~n53542;
  assign n53544 = ~n29192 & ~n42519;
  assign n53545 = controllable_nhgrant0 & ~n53544;
  assign n53546 = ~n14725 & ~n53545;
  assign n53547 = ~n3281 & ~n53546;
  assign n53548 = ~n3281 & ~n53547;
  assign n53549 = n3492 & ~n53548;
  assign n53550 = ~n14836 & ~n53549;
  assign n53551 = n3485 & ~n53550;
  assign n53552 = ~n14835 & ~n53551;
  assign n53553 = n3476 & ~n53552;
  assign n53554 = ~n53543 & ~n53553;
  assign n53555 = n3374 & ~n53554;
  assign n53556 = n3374 & ~n53555;
  assign n53557 = ~n3655 & ~n53556;
  assign n53558 = ~n53533 & ~n53557;
  assign n53559 = ~n3652 & ~n53558;
  assign n53560 = ~n53509 & ~n53559;
  assign n53561 = n3368 & ~n53560;
  assign n53562 = ~n53459 & ~n53561;
  assign n53563 = ~n3362 & ~n53562;
  assign n53564 = ~n3362 & ~n53563;
  assign n53565 = ~n3359 & ~n53564;
  assign n53566 = ~n3359 & ~n53565;
  assign n53567 = n3356 & ~n53566;
  assign n53568 = ~n25649 & ~n39584;
  assign n53569 = controllable_nhgrant0 & ~n53568;
  assign n53570 = ~n5245 & ~n53569;
  assign n53571 = ~n3281 & ~n53570;
  assign n53572 = ~n3783 & ~n53571;
  assign n53573 = ~n3378 & ~n53572;
  assign n53574 = ~n14959 & ~n53573;
  assign n53575 = n3492 & ~n53574;
  assign n53576 = ~n3631 & ~n53575;
  assign n53577 = n3485 & ~n53576;
  assign n53578 = ~n3630 & ~n53577;
  assign n53579 = ~n3374 & ~n53578;
  assign n53580 = ~n29318 & ~n42561;
  assign n53581 = controllable_nhgrant0 & ~n53580;
  assign n53582 = ~n15006 & ~n53581;
  assign n53583 = ~n3281 & ~n53582;
  assign n53584 = ~n3950 & ~n53583;
  assign n53585 = n3378 & ~n53584;
  assign n53586 = ~n25684 & ~n42579;
  assign n53587 = controllable_nhgrant0 & ~n53586;
  assign n53588 = ~n5534 & ~n53587;
  assign n53589 = ~n3281 & ~n53588;
  assign n53590 = ~n3950 & ~n53589;
  assign n53591 = ~n3378 & ~n53590;
  assign n53592 = ~n53585 & ~n53591;
  assign n53593 = n3492 & ~n53592;
  assign n53594 = ~n3631 & ~n53593;
  assign n53595 = n3485 & ~n53594;
  assign n53596 = ~n3630 & ~n53595;
  assign n53597 = ~n3476 & ~n53596;
  assign n53598 = ~n29348 & ~n42607;
  assign n53599 = controllable_nhgrant0 & ~n53598;
  assign n53600 = ~n15088 & ~n53599;
  assign n53601 = ~n3281 & ~n53600;
  assign n53602 = ~n4089 & ~n53601;
  assign n53603 = n3378 & ~n53602;
  assign n53604 = ~n25726 & ~n42627;
  assign n53605 = controllable_nhgrant0 & ~n53604;
  assign n53606 = ~n6082 & ~n53605;
  assign n53607 = ~n3281 & ~n53606;
  assign n53608 = ~n4089 & ~n53607;
  assign n53609 = ~n3378 & ~n53608;
  assign n53610 = ~n53603 & ~n53609;
  assign n53611 = n3492 & ~n53610;
  assign n53612 = ~n3631 & ~n53611;
  assign n53613 = n3485 & ~n53612;
  assign n53614 = ~n3630 & ~n53613;
  assign n53615 = n3476 & ~n53614;
  assign n53616 = ~n53597 & ~n53615;
  assign n53617 = n3374 & ~n53616;
  assign n53618 = ~n53579 & ~n53617;
  assign n53619 = n3655 & ~n53618;
  assign n53620 = ~n25649 & ~n39791;
  assign n53621 = controllable_nhgrant0 & ~n53620;
  assign n53622 = ~n5245 & ~n53621;
  assign n53623 = ~n3281 & ~n53622;
  assign n53624 = ~n3783 & ~n53623;
  assign n53625 = ~n3378 & ~n53624;
  assign n53626 = ~n14959 & ~n53625;
  assign n53627 = n3492 & ~n53626;
  assign n53628 = ~n3631 & ~n53627;
  assign n53629 = n3485 & ~n53628;
  assign n53630 = ~n3630 & ~n53629;
  assign n53631 = ~n3374 & ~n53630;
  assign n53632 = ~n29318 & ~n42661;
  assign n53633 = controllable_nhgrant0 & ~n53632;
  assign n53634 = ~n15006 & ~n53633;
  assign n53635 = ~n3281 & ~n53634;
  assign n53636 = ~n3950 & ~n53635;
  assign n53637 = n3378 & ~n53636;
  assign n53638 = ~n25684 & ~n42679;
  assign n53639 = controllable_nhgrant0 & ~n53638;
  assign n53640 = ~n5534 & ~n53639;
  assign n53641 = ~n3281 & ~n53640;
  assign n53642 = ~n3950 & ~n53641;
  assign n53643 = ~n3378 & ~n53642;
  assign n53644 = ~n53637 & ~n53643;
  assign n53645 = n3492 & ~n53644;
  assign n53646 = ~n3631 & ~n53645;
  assign n53647 = n3485 & ~n53646;
  assign n53648 = ~n3630 & ~n53647;
  assign n53649 = ~n3476 & ~n53648;
  assign n53650 = ~n29348 & ~n42707;
  assign n53651 = controllable_nhgrant0 & ~n53650;
  assign n53652 = ~n15088 & ~n53651;
  assign n53653 = ~n3281 & ~n53652;
  assign n53654 = ~n4089 & ~n53653;
  assign n53655 = n3378 & ~n53654;
  assign n53656 = ~n25726 & ~n42727;
  assign n53657 = controllable_nhgrant0 & ~n53656;
  assign n53658 = ~n6082 & ~n53657;
  assign n53659 = ~n3281 & ~n53658;
  assign n53660 = ~n4089 & ~n53659;
  assign n53661 = ~n3378 & ~n53660;
  assign n53662 = ~n53655 & ~n53661;
  assign n53663 = n3492 & ~n53662;
  assign n53664 = ~n3631 & ~n53663;
  assign n53665 = n3485 & ~n53664;
  assign n53666 = ~n3630 & ~n53665;
  assign n53667 = n3476 & ~n53666;
  assign n53668 = ~n53649 & ~n53667;
  assign n53669 = n3374 & ~n53668;
  assign n53670 = ~n53631 & ~n53669;
  assign n53671 = ~n3655 & ~n53670;
  assign n53672 = ~n53619 & ~n53671;
  assign n53673 = n3652 & ~n53672;
  assign n53674 = ~n25649 & ~n42763;
  assign n53675 = controllable_nhgrant0 & ~n53674;
  assign n53676 = ~n5245 & ~n53675;
  assign n53677 = ~n3281 & ~n53676;
  assign n53678 = ~n3783 & ~n53677;
  assign n53679 = ~n3378 & ~n53678;
  assign n53680 = ~n15225 & ~n53679;
  assign n53681 = n3492 & ~n53680;
  assign n53682 = ~n3631 & ~n53681;
  assign n53683 = n3485 & ~n53682;
  assign n53684 = ~n3630 & ~n53683;
  assign n53685 = ~n3476 & ~n53684;
  assign n53686 = ~n15258 & ~n53681;
  assign n53687 = n3485 & ~n53686;
  assign n53688 = ~n15257 & ~n53687;
  assign n53689 = n3476 & ~n53688;
  assign n53690 = ~n53685 & ~n53689;
  assign n53691 = ~n3374 & ~n53690;
  assign n53692 = ~n29318 & ~n42793;
  assign n53693 = controllable_nhgrant0 & ~n53692;
  assign n53694 = ~n15006 & ~n53693;
  assign n53695 = ~n3281 & ~n53694;
  assign n53696 = ~n3950 & ~n53695;
  assign n53697 = n3378 & ~n53696;
  assign n53698 = ~n25684 & ~n42827;
  assign n53699 = controllable_nhgrant0 & ~n53698;
  assign n53700 = ~n5534 & ~n53699;
  assign n53701 = ~n3281 & ~n53700;
  assign n53702 = ~n3950 & ~n53701;
  assign n53703 = ~n3378 & ~n53702;
  assign n53704 = ~n53697 & ~n53703;
  assign n53705 = n3492 & ~n53704;
  assign n53706 = ~n3631 & ~n53705;
  assign n53707 = n3485 & ~n53706;
  assign n53708 = ~n3630 & ~n53707;
  assign n53709 = ~n3476 & ~n53708;
  assign n53710 = ~n29348 & ~n42855;
  assign n53711 = controllable_nhgrant0 & ~n53710;
  assign n53712 = ~n15088 & ~n53711;
  assign n53713 = ~n3281 & ~n53712;
  assign n53714 = ~n4089 & ~n53713;
  assign n53715 = n3378 & ~n53714;
  assign n53716 = ~n25726 & ~n42891;
  assign n53717 = controllable_nhgrant0 & ~n53716;
  assign n53718 = ~n6082 & ~n53717;
  assign n53719 = ~n3281 & ~n53718;
  assign n53720 = ~n4089 & ~n53719;
  assign n53721 = ~n3378 & ~n53720;
  assign n53722 = ~n53715 & ~n53721;
  assign n53723 = n3492 & ~n53722;
  assign n53724 = ~n15258 & ~n53723;
  assign n53725 = n3485 & ~n53724;
  assign n53726 = ~n15257 & ~n53725;
  assign n53727 = n3476 & ~n53726;
  assign n53728 = ~n53709 & ~n53727;
  assign n53729 = n3374 & ~n53728;
  assign n53730 = ~n53691 & ~n53729;
  assign n53731 = n3655 & ~n53730;
  assign n53732 = ~n25649 & ~n42925;
  assign n53733 = controllable_nhgrant0 & ~n53732;
  assign n53734 = ~n5245 & ~n53733;
  assign n53735 = ~n3281 & ~n53734;
  assign n53736 = ~n3783 & ~n53735;
  assign n53737 = ~n3378 & ~n53736;
  assign n53738 = ~n15225 & ~n53737;
  assign n53739 = n3492 & ~n53738;
  assign n53740 = ~n3631 & ~n53739;
  assign n53741 = n3485 & ~n53740;
  assign n53742 = ~n3630 & ~n53741;
  assign n53743 = ~n3476 & ~n53742;
  assign n53744 = ~n15258 & ~n53739;
  assign n53745 = n3485 & ~n53744;
  assign n53746 = ~n15257 & ~n53745;
  assign n53747 = n3476 & ~n53746;
  assign n53748 = ~n53743 & ~n53747;
  assign n53749 = ~n3374 & ~n53748;
  assign n53750 = ~n29318 & ~n42955;
  assign n53751 = controllable_nhgrant0 & ~n53750;
  assign n53752 = ~n15006 & ~n53751;
  assign n53753 = ~n3281 & ~n53752;
  assign n53754 = ~n3950 & ~n53753;
  assign n53755 = n3378 & ~n53754;
  assign n53756 = ~n25684 & ~n42989;
  assign n53757 = controllable_nhgrant0 & ~n53756;
  assign n53758 = ~n5534 & ~n53757;
  assign n53759 = ~n3281 & ~n53758;
  assign n53760 = ~n3950 & ~n53759;
  assign n53761 = ~n3378 & ~n53760;
  assign n53762 = ~n53755 & ~n53761;
  assign n53763 = n3492 & ~n53762;
  assign n53764 = ~n3631 & ~n53763;
  assign n53765 = n3485 & ~n53764;
  assign n53766 = ~n3630 & ~n53765;
  assign n53767 = ~n3476 & ~n53766;
  assign n53768 = ~n29348 & ~n43017;
  assign n53769 = controllable_nhgrant0 & ~n53768;
  assign n53770 = ~n15088 & ~n53769;
  assign n53771 = ~n3281 & ~n53770;
  assign n53772 = ~n4089 & ~n53771;
  assign n53773 = n3378 & ~n53772;
  assign n53774 = ~n25726 & ~n43053;
  assign n53775 = controllable_nhgrant0 & ~n53774;
  assign n53776 = ~n6082 & ~n53775;
  assign n53777 = ~n3281 & ~n53776;
  assign n53778 = ~n4089 & ~n53777;
  assign n53779 = ~n3378 & ~n53778;
  assign n53780 = ~n53773 & ~n53779;
  assign n53781 = n3492 & ~n53780;
  assign n53782 = ~n15258 & ~n53781;
  assign n53783 = n3485 & ~n53782;
  assign n53784 = ~n15257 & ~n53783;
  assign n53785 = n3476 & ~n53784;
  assign n53786 = ~n53767 & ~n53785;
  assign n53787 = n3374 & ~n53786;
  assign n53788 = ~n53749 & ~n53787;
  assign n53789 = ~n3655 & ~n53788;
  assign n53790 = ~n53731 & ~n53789;
  assign n53791 = ~n3652 & ~n53790;
  assign n53792 = ~n53673 & ~n53791;
  assign n53793 = ~n3368 & ~n53792;
  assign n53794 = ~n25905 & ~n40313;
  assign n53795 = controllable_nhgrant0 & ~n53794;
  assign n53796 = ~n7118 & ~n53795;
  assign n53797 = ~n3281 & ~n53796;
  assign n53798 = ~n3281 & ~n53797;
  assign n53799 = ~n3378 & ~n53798;
  assign n53800 = ~n7082 & ~n53799;
  assign n53801 = n3492 & ~n53800;
  assign n53802 = n3492 & ~n53801;
  assign n53803 = n3485 & ~n53802;
  assign n53804 = n3485 & ~n53803;
  assign n53805 = ~n3374 & ~n53804;
  assign n53806 = ~n29550 & ~n43085;
  assign n53807 = controllable_nhgrant0 & ~n53806;
  assign n53808 = ~n15675 & ~n53807;
  assign n53809 = ~n3281 & ~n53808;
  assign n53810 = ~n3281 & ~n53809;
  assign n53811 = n3378 & ~n53810;
  assign n53812 = ~n29568 & ~n43103;
  assign n53813 = controllable_nhgrant0 & ~n53812;
  assign n53814 = ~n15716 & ~n53813;
  assign n53815 = ~n3281 & ~n53814;
  assign n53816 = ~n3281 & ~n53815;
  assign n53817 = ~n3378 & ~n53816;
  assign n53818 = ~n53811 & ~n53817;
  assign n53819 = n3492 & ~n53818;
  assign n53820 = n3492 & ~n53819;
  assign n53821 = n3485 & ~n53820;
  assign n53822 = n3485 & ~n53821;
  assign n53823 = ~n3476 & ~n53822;
  assign n53824 = ~n29592 & ~n43131;
  assign n53825 = controllable_nhgrant0 & ~n53824;
  assign n53826 = ~n15783 & ~n53825;
  assign n53827 = ~n3281 & ~n53826;
  assign n53828 = ~n3281 & ~n53827;
  assign n53829 = n3378 & ~n53828;
  assign n53830 = ~n29610 & ~n43173;
  assign n53831 = controllable_nhgrant0 & ~n53830;
  assign n53832 = ~n15846 & ~n53831;
  assign n53833 = ~n3281 & ~n53832;
  assign n53834 = ~n3281 & ~n53833;
  assign n53835 = ~n3378 & ~n53834;
  assign n53836 = ~n53829 & ~n53835;
  assign n53837 = n3492 & ~n53836;
  assign n53838 = n3492 & ~n53837;
  assign n53839 = n3485 & ~n53838;
  assign n53840 = n3485 & ~n53839;
  assign n53841 = n3476 & ~n53840;
  assign n53842 = ~n53823 & ~n53841;
  assign n53843 = n3374 & ~n53842;
  assign n53844 = ~n53805 & ~n53843;
  assign n53845 = n3655 & ~n53844;
  assign n53846 = ~n25905 & ~n40529;
  assign n53847 = controllable_nhgrant0 & ~n53846;
  assign n53848 = ~n7118 & ~n53847;
  assign n53849 = ~n3281 & ~n53848;
  assign n53850 = ~n3281 & ~n53849;
  assign n53851 = ~n3378 & ~n53850;
  assign n53852 = ~n7082 & ~n53851;
  assign n53853 = n3492 & ~n53852;
  assign n53854 = n3492 & ~n53853;
  assign n53855 = n3485 & ~n53854;
  assign n53856 = n3485 & ~n53855;
  assign n53857 = ~n3374 & ~n53856;
  assign n53858 = ~n29550 & ~n43201;
  assign n53859 = controllable_nhgrant0 & ~n53858;
  assign n53860 = ~n15675 & ~n53859;
  assign n53861 = ~n3281 & ~n53860;
  assign n53862 = ~n3281 & ~n53861;
  assign n53863 = n3378 & ~n53862;
  assign n53864 = ~n29568 & ~n43219;
  assign n53865 = controllable_nhgrant0 & ~n53864;
  assign n53866 = ~n15716 & ~n53865;
  assign n53867 = ~n3281 & ~n53866;
  assign n53868 = ~n3281 & ~n53867;
  assign n53869 = ~n3378 & ~n53868;
  assign n53870 = ~n53863 & ~n53869;
  assign n53871 = n3492 & ~n53870;
  assign n53872 = n3492 & ~n53871;
  assign n53873 = n3485 & ~n53872;
  assign n53874 = n3485 & ~n53873;
  assign n53875 = ~n3476 & ~n53874;
  assign n53876 = ~n29592 & ~n43247;
  assign n53877 = controllable_nhgrant0 & ~n53876;
  assign n53878 = ~n15783 & ~n53877;
  assign n53879 = ~n3281 & ~n53878;
  assign n53880 = ~n3281 & ~n53879;
  assign n53881 = n3378 & ~n53880;
  assign n53882 = ~n29610 & ~n43289;
  assign n53883 = controllable_nhgrant0 & ~n53882;
  assign n53884 = ~n15846 & ~n53883;
  assign n53885 = ~n3281 & ~n53884;
  assign n53886 = ~n3281 & ~n53885;
  assign n53887 = ~n3378 & ~n53886;
  assign n53888 = ~n53881 & ~n53887;
  assign n53889 = n3492 & ~n53888;
  assign n53890 = n3492 & ~n53889;
  assign n53891 = n3485 & ~n53890;
  assign n53892 = n3485 & ~n53891;
  assign n53893 = n3476 & ~n53892;
  assign n53894 = ~n53875 & ~n53893;
  assign n53895 = n3374 & ~n53894;
  assign n53896 = ~n53857 & ~n53895;
  assign n53897 = ~n3655 & ~n53896;
  assign n53898 = ~n53845 & ~n53897;
  assign n53899 = n3652 & ~n53898;
  assign n53900 = ~n25905 & ~n43325;
  assign n53901 = controllable_nhgrant0 & ~n53900;
  assign n53902 = ~n7118 & ~n53901;
  assign n53903 = ~n3281 & ~n53902;
  assign n53904 = ~n3281 & ~n53903;
  assign n53905 = ~n3378 & ~n53904;
  assign n53906 = ~n16013 & ~n53905;
  assign n53907 = n3492 & ~n53906;
  assign n53908 = n3492 & ~n53907;
  assign n53909 = n3485 & ~n53908;
  assign n53910 = n3485 & ~n53909;
  assign n53911 = ~n3374 & ~n53910;
  assign n53912 = ~n29550 & ~n43349;
  assign n53913 = controllable_nhgrant0 & ~n53912;
  assign n53914 = ~n15675 & ~n53913;
  assign n53915 = ~n3281 & ~n53914;
  assign n53916 = ~n3281 & ~n53915;
  assign n53917 = n3378 & ~n53916;
  assign n53918 = ~n29568 & ~n43396;
  assign n53919 = controllable_nhgrant0 & ~n53918;
  assign n53920 = ~n15716 & ~n53919;
  assign n53921 = ~n3281 & ~n53920;
  assign n53922 = ~n3281 & ~n53921;
  assign n53923 = ~n3378 & ~n53922;
  assign n53924 = ~n53917 & ~n53923;
  assign n53925 = n3492 & ~n53924;
  assign n53926 = n3492 & ~n53925;
  assign n53927 = n3485 & ~n53926;
  assign n53928 = n3485 & ~n53927;
  assign n53929 = ~n3476 & ~n53928;
  assign n53930 = ~n29592 & ~n43424;
  assign n53931 = controllable_nhgrant0 & ~n53930;
  assign n53932 = ~n15783 & ~n53931;
  assign n53933 = ~n3281 & ~n53932;
  assign n53934 = ~n3281 & ~n53933;
  assign n53935 = n3378 & ~n53934;
  assign n53936 = ~n29610 & ~n43481;
  assign n53937 = controllable_nhgrant0 & ~n53936;
  assign n53938 = ~n15846 & ~n53937;
  assign n53939 = ~n3281 & ~n53938;
  assign n53940 = ~n3281 & ~n53939;
  assign n53941 = ~n3378 & ~n53940;
  assign n53942 = ~n53935 & ~n53941;
  assign n53943 = n3492 & ~n53942;
  assign n53944 = ~n14836 & ~n53943;
  assign n53945 = n3485 & ~n53944;
  assign n53946 = ~n14835 & ~n53945;
  assign n53947 = n3476 & ~n53946;
  assign n53948 = ~n53929 & ~n53947;
  assign n53949 = n3374 & ~n53948;
  assign n53950 = ~n53911 & ~n53949;
  assign n53951 = n3655 & ~n53950;
  assign n53952 = ~n25905 & ~n43515;
  assign n53953 = controllable_nhgrant0 & ~n53952;
  assign n53954 = ~n7118 & ~n53953;
  assign n53955 = ~n3281 & ~n53954;
  assign n53956 = ~n3281 & ~n53955;
  assign n53957 = ~n3378 & ~n53956;
  assign n53958 = ~n16013 & ~n53957;
  assign n53959 = n3492 & ~n53958;
  assign n53960 = n3492 & ~n53959;
  assign n53961 = n3485 & ~n53960;
  assign n53962 = n3485 & ~n53961;
  assign n53963 = ~n3374 & ~n53962;
  assign n53964 = ~n29550 & ~n43539;
  assign n53965 = controllable_nhgrant0 & ~n53964;
  assign n53966 = ~n15675 & ~n53965;
  assign n53967 = ~n3281 & ~n53966;
  assign n53968 = ~n3281 & ~n53967;
  assign n53969 = n3378 & ~n53968;
  assign n53970 = ~n29568 & ~n43586;
  assign n53971 = controllable_nhgrant0 & ~n53970;
  assign n53972 = ~n15716 & ~n53971;
  assign n53973 = ~n3281 & ~n53972;
  assign n53974 = ~n3281 & ~n53973;
  assign n53975 = ~n3378 & ~n53974;
  assign n53976 = ~n53969 & ~n53975;
  assign n53977 = n3492 & ~n53976;
  assign n53978 = n3492 & ~n53977;
  assign n53979 = n3485 & ~n53978;
  assign n53980 = n3485 & ~n53979;
  assign n53981 = ~n3476 & ~n53980;
  assign n53982 = ~n29592 & ~n43614;
  assign n53983 = controllable_nhgrant0 & ~n53982;
  assign n53984 = ~n15783 & ~n53983;
  assign n53985 = ~n3281 & ~n53984;
  assign n53986 = ~n3281 & ~n53985;
  assign n53987 = n3378 & ~n53986;
  assign n53988 = ~n29610 & ~n43671;
  assign n53989 = controllable_nhgrant0 & ~n53988;
  assign n53990 = ~n15846 & ~n53989;
  assign n53991 = ~n3281 & ~n53990;
  assign n53992 = ~n3281 & ~n53991;
  assign n53993 = ~n3378 & ~n53992;
  assign n53994 = ~n53987 & ~n53993;
  assign n53995 = n3492 & ~n53994;
  assign n53996 = ~n14836 & ~n53995;
  assign n53997 = n3485 & ~n53996;
  assign n53998 = ~n14835 & ~n53997;
  assign n53999 = n3476 & ~n53998;
  assign n54000 = ~n53981 & ~n53999;
  assign n54001 = n3374 & ~n54000;
  assign n54002 = ~n53963 & ~n54001;
  assign n54003 = ~n3655 & ~n54002;
  assign n54004 = ~n53951 & ~n54003;
  assign n54005 = ~n3652 & ~n54004;
  assign n54006 = ~n53899 & ~n54005;
  assign n54007 = n3368 & ~n54006;
  assign n54008 = ~n53793 & ~n54007;
  assign n54009 = n3362 & ~n54008;
  assign n54010 = n3492 & ~n53572;
  assign n54011 = ~n3631 & ~n54010;
  assign n54012 = n3485 & ~n54011;
  assign n54013 = ~n3630 & ~n54012;
  assign n54014 = ~n3476 & ~n54013;
  assign n54015 = ~n8310 & ~n51148;
  assign n54016 = ~n3485 & ~n54015;
  assign n54017 = ~n54012 & ~n54016;
  assign n54018 = n3476 & ~n54017;
  assign n54019 = ~n54014 & ~n54018;
  assign n54020 = ~n3374 & ~n54019;
  assign n54021 = n3492 & ~n53590;
  assign n54022 = ~n3631 & ~n54021;
  assign n54023 = n3485 & ~n54022;
  assign n54024 = ~n3630 & ~n54023;
  assign n54025 = ~n3476 & ~n54024;
  assign n54026 = n3492 & ~n53608;
  assign n54027 = ~n3631 & ~n54026;
  assign n54028 = n3485 & ~n54027;
  assign n54029 = ~n54016 & ~n54028;
  assign n54030 = n3476 & ~n54029;
  assign n54031 = ~n54025 & ~n54030;
  assign n54032 = n3374 & ~n54031;
  assign n54033 = ~n54020 & ~n54032;
  assign n54034 = n3655 & ~n54033;
  assign n54035 = n3492 & ~n53624;
  assign n54036 = ~n3631 & ~n54035;
  assign n54037 = n3485 & ~n54036;
  assign n54038 = ~n3630 & ~n54037;
  assign n54039 = ~n3476 & ~n54038;
  assign n54040 = ~n8310 & ~n51191;
  assign n54041 = ~n3485 & ~n54040;
  assign n54042 = ~n54037 & ~n54041;
  assign n54043 = n3476 & ~n54042;
  assign n54044 = ~n54039 & ~n54043;
  assign n54045 = ~n3374 & ~n54044;
  assign n54046 = n3492 & ~n53642;
  assign n54047 = ~n3631 & ~n54046;
  assign n54048 = n3485 & ~n54047;
  assign n54049 = ~n3630 & ~n54048;
  assign n54050 = ~n3476 & ~n54049;
  assign n54051 = n3492 & ~n53660;
  assign n54052 = ~n3631 & ~n54051;
  assign n54053 = n3485 & ~n54052;
  assign n54054 = ~n54041 & ~n54053;
  assign n54055 = n3476 & ~n54054;
  assign n54056 = ~n54050 & ~n54055;
  assign n54057 = n3374 & ~n54056;
  assign n54058 = ~n54045 & ~n54057;
  assign n54059 = ~n3655 & ~n54058;
  assign n54060 = ~n54034 & ~n54059;
  assign n54061 = n3652 & ~n54060;
  assign n54062 = n3492 & ~n53678;
  assign n54063 = ~n3631 & ~n54062;
  assign n54064 = n3485 & ~n54063;
  assign n54065 = ~n3630 & ~n54064;
  assign n54066 = ~n3476 & ~n54065;
  assign n54067 = ~n16588 & ~n51236;
  assign n54068 = ~n3485 & ~n54067;
  assign n54069 = ~n15258 & ~n54062;
  assign n54070 = n3485 & ~n54069;
  assign n54071 = ~n54068 & ~n54070;
  assign n54072 = n3476 & ~n54071;
  assign n54073 = ~n54066 & ~n54072;
  assign n54074 = ~n3374 & ~n54073;
  assign n54075 = n3492 & ~n53702;
  assign n54076 = ~n3631 & ~n54075;
  assign n54077 = n3485 & ~n54076;
  assign n54078 = ~n3630 & ~n54077;
  assign n54079 = ~n3476 & ~n54078;
  assign n54080 = n3492 & ~n53720;
  assign n54081 = ~n15258 & ~n54080;
  assign n54082 = n3485 & ~n54081;
  assign n54083 = ~n54068 & ~n54082;
  assign n54084 = n3476 & ~n54083;
  assign n54085 = ~n54079 & ~n54084;
  assign n54086 = n3374 & ~n54085;
  assign n54087 = ~n54074 & ~n54086;
  assign n54088 = n3655 & ~n54087;
  assign n54089 = n3492 & ~n53736;
  assign n54090 = ~n3631 & ~n54089;
  assign n54091 = n3485 & ~n54090;
  assign n54092 = ~n3630 & ~n54091;
  assign n54093 = ~n3476 & ~n54092;
  assign n54094 = ~n16588 & ~n51279;
  assign n54095 = ~n3485 & ~n54094;
  assign n54096 = ~n15258 & ~n54089;
  assign n54097 = n3485 & ~n54096;
  assign n54098 = ~n54095 & ~n54097;
  assign n54099 = n3476 & ~n54098;
  assign n54100 = ~n54093 & ~n54099;
  assign n54101 = ~n3374 & ~n54100;
  assign n54102 = n3492 & ~n53760;
  assign n54103 = ~n3631 & ~n54102;
  assign n54104 = n3485 & ~n54103;
  assign n54105 = ~n3630 & ~n54104;
  assign n54106 = ~n3476 & ~n54105;
  assign n54107 = n3492 & ~n53778;
  assign n54108 = ~n15258 & ~n54107;
  assign n54109 = n3485 & ~n54108;
  assign n54110 = ~n54095 & ~n54109;
  assign n54111 = n3476 & ~n54110;
  assign n54112 = ~n54106 & ~n54111;
  assign n54113 = n3374 & ~n54112;
  assign n54114 = ~n54101 & ~n54113;
  assign n54115 = ~n3655 & ~n54114;
  assign n54116 = ~n54088 & ~n54115;
  assign n54117 = ~n3652 & ~n54116;
  assign n54118 = ~n54061 & ~n54117;
  assign n54119 = ~n3368 & ~n54118;
  assign n54120 = n3492 & ~n53798;
  assign n54121 = n3492 & ~n54120;
  assign n54122 = n3485 & ~n54121;
  assign n54123 = n3485 & ~n54122;
  assign n54124 = ~n3476 & ~n54123;
  assign n54125 = ~n8525 & ~n54122;
  assign n54126 = n3476 & ~n54125;
  assign n54127 = ~n54124 & ~n54126;
  assign n54128 = ~n3374 & ~n54127;
  assign n54129 = n3492 & ~n53816;
  assign n54130 = n3492 & ~n54129;
  assign n54131 = n3485 & ~n54130;
  assign n54132 = n3485 & ~n54131;
  assign n54133 = ~n3476 & ~n54132;
  assign n54134 = ~n3492 & ~n51321;
  assign n54135 = ~n3485 & ~n54134;
  assign n54136 = n3492 & ~n53834;
  assign n54137 = n3492 & ~n54136;
  assign n54138 = n3485 & ~n54137;
  assign n54139 = ~n54135 & ~n54138;
  assign n54140 = n3476 & ~n54139;
  assign n54141 = ~n54133 & ~n54140;
  assign n54142 = n3374 & ~n54141;
  assign n54143 = ~n54128 & ~n54142;
  assign n54144 = n3655 & ~n54143;
  assign n54145 = n3492 & ~n53850;
  assign n54146 = n3492 & ~n54145;
  assign n54147 = n3485 & ~n54146;
  assign n54148 = n3485 & ~n54147;
  assign n54149 = ~n3476 & ~n54148;
  assign n54150 = ~n8525 & ~n54147;
  assign n54151 = n3476 & ~n54150;
  assign n54152 = ~n54149 & ~n54151;
  assign n54153 = ~n3374 & ~n54152;
  assign n54154 = n3492 & ~n53868;
  assign n54155 = n3492 & ~n54154;
  assign n54156 = n3485 & ~n54155;
  assign n54157 = n3485 & ~n54156;
  assign n54158 = ~n3476 & ~n54157;
  assign n54159 = ~n3492 & ~n51348;
  assign n54160 = ~n3485 & ~n54159;
  assign n54161 = n3492 & ~n53886;
  assign n54162 = n3492 & ~n54161;
  assign n54163 = n3485 & ~n54162;
  assign n54164 = ~n54160 & ~n54163;
  assign n54165 = n3476 & ~n54164;
  assign n54166 = ~n54158 & ~n54165;
  assign n54167 = n3374 & ~n54166;
  assign n54168 = ~n54153 & ~n54167;
  assign n54169 = ~n3655 & ~n54168;
  assign n54170 = ~n54144 & ~n54169;
  assign n54171 = n3652 & ~n54170;
  assign n54172 = n3492 & ~n53904;
  assign n54173 = n3492 & ~n54172;
  assign n54174 = n3485 & ~n54173;
  assign n54175 = n3485 & ~n54174;
  assign n54176 = ~n3476 & ~n54175;
  assign n54177 = ~n8525 & ~n54174;
  assign n54178 = n3476 & ~n54177;
  assign n54179 = ~n54176 & ~n54178;
  assign n54180 = ~n3374 & ~n54179;
  assign n54181 = n3492 & ~n53922;
  assign n54182 = n3492 & ~n54181;
  assign n54183 = n3485 & ~n54182;
  assign n54184 = n3485 & ~n54183;
  assign n54185 = ~n3476 & ~n54184;
  assign n54186 = ~n16686 & ~n51377;
  assign n54187 = ~n3485 & ~n54186;
  assign n54188 = n3492 & ~n53940;
  assign n54189 = ~n14836 & ~n54188;
  assign n54190 = n3485 & ~n54189;
  assign n54191 = ~n54187 & ~n54190;
  assign n54192 = n3476 & ~n54191;
  assign n54193 = ~n54185 & ~n54192;
  assign n54194 = n3374 & ~n54193;
  assign n54195 = ~n54180 & ~n54194;
  assign n54196 = n3655 & ~n54195;
  assign n54197 = n3492 & ~n53956;
  assign n54198 = n3492 & ~n54197;
  assign n54199 = n3485 & ~n54198;
  assign n54200 = n3485 & ~n54199;
  assign n54201 = ~n3476 & ~n54200;
  assign n54202 = ~n8525 & ~n54199;
  assign n54203 = n3476 & ~n54202;
  assign n54204 = ~n54201 & ~n54203;
  assign n54205 = ~n3374 & ~n54204;
  assign n54206 = n3492 & ~n53974;
  assign n54207 = n3492 & ~n54206;
  assign n54208 = n3485 & ~n54207;
  assign n54209 = n3485 & ~n54208;
  assign n54210 = ~n3476 & ~n54209;
  assign n54211 = ~n16686 & ~n51404;
  assign n54212 = ~n3485 & ~n54211;
  assign n54213 = n3492 & ~n53992;
  assign n54214 = ~n14836 & ~n54213;
  assign n54215 = n3485 & ~n54214;
  assign n54216 = ~n54212 & ~n54215;
  assign n54217 = n3476 & ~n54216;
  assign n54218 = ~n54210 & ~n54217;
  assign n54219 = n3374 & ~n54218;
  assign n54220 = ~n54205 & ~n54219;
  assign n54221 = ~n3655 & ~n54220;
  assign n54222 = ~n54196 & ~n54221;
  assign n54223 = ~n3652 & ~n54222;
  assign n54224 = ~n54171 & ~n54223;
  assign n54225 = n3368 & ~n54224;
  assign n54226 = ~n54119 & ~n54225;
  assign n54227 = ~n3362 & ~n54226;
  assign n54228 = ~n54009 & ~n54227;
  assign n54229 = n3359 & ~n54228;
  assign n54230 = ~n51424 & ~n54012;
  assign n54231 = n3476 & ~n54230;
  assign n54232 = ~n54014 & ~n54231;
  assign n54233 = ~n3374 & ~n54232;
  assign n54234 = ~n51424 & ~n54028;
  assign n54235 = n3476 & ~n54234;
  assign n54236 = ~n54025 & ~n54235;
  assign n54237 = n3374 & ~n54236;
  assign n54238 = ~n54233 & ~n54237;
  assign n54239 = n3655 & ~n54238;
  assign n54240 = ~n51435 & ~n54037;
  assign n54241 = n3476 & ~n54240;
  assign n54242 = ~n54039 & ~n54241;
  assign n54243 = ~n3374 & ~n54242;
  assign n54244 = ~n51435 & ~n54053;
  assign n54245 = n3476 & ~n54244;
  assign n54246 = ~n54050 & ~n54245;
  assign n54247 = n3374 & ~n54246;
  assign n54248 = ~n54243 & ~n54247;
  assign n54249 = ~n3655 & ~n54248;
  assign n54250 = ~n54239 & ~n54249;
  assign n54251 = n3652 & ~n54250;
  assign n54252 = ~n51448 & ~n54070;
  assign n54253 = n3476 & ~n54252;
  assign n54254 = ~n54066 & ~n54253;
  assign n54255 = ~n3374 & ~n54254;
  assign n54256 = ~n51448 & ~n54082;
  assign n54257 = n3476 & ~n54256;
  assign n54258 = ~n54079 & ~n54257;
  assign n54259 = n3374 & ~n54258;
  assign n54260 = ~n54255 & ~n54259;
  assign n54261 = n3655 & ~n54260;
  assign n54262 = ~n51459 & ~n54097;
  assign n54263 = n3476 & ~n54262;
  assign n54264 = ~n54093 & ~n54263;
  assign n54265 = ~n3374 & ~n54264;
  assign n54266 = ~n51459 & ~n54109;
  assign n54267 = n3476 & ~n54266;
  assign n54268 = ~n54106 & ~n54267;
  assign n54269 = n3374 & ~n54268;
  assign n54270 = ~n54265 & ~n54269;
  assign n54271 = ~n3655 & ~n54270;
  assign n54272 = ~n54261 & ~n54271;
  assign n54273 = ~n3652 & ~n54272;
  assign n54274 = ~n54251 & ~n54273;
  assign n54275 = ~n3368 & ~n54274;
  assign n54276 = ~n8689 & ~n54122;
  assign n54277 = n3476 & ~n54276;
  assign n54278 = ~n54124 & ~n54277;
  assign n54279 = ~n3374 & ~n54278;
  assign n54280 = ~n51478 & ~n54138;
  assign n54281 = n3476 & ~n54280;
  assign n54282 = ~n54133 & ~n54281;
  assign n54283 = n3374 & ~n54282;
  assign n54284 = ~n54279 & ~n54283;
  assign n54285 = n3655 & ~n54284;
  assign n54286 = ~n8689 & ~n54147;
  assign n54287 = n3476 & ~n54286;
  assign n54288 = ~n54149 & ~n54287;
  assign n54289 = ~n3374 & ~n54288;
  assign n54290 = ~n51489 & ~n54163;
  assign n54291 = n3476 & ~n54290;
  assign n54292 = ~n54158 & ~n54291;
  assign n54293 = n3374 & ~n54292;
  assign n54294 = ~n54289 & ~n54293;
  assign n54295 = ~n3655 & ~n54294;
  assign n54296 = ~n54285 & ~n54295;
  assign n54297 = n3652 & ~n54296;
  assign n54298 = ~n8689 & ~n54174;
  assign n54299 = n3476 & ~n54298;
  assign n54300 = ~n54176 & ~n54299;
  assign n54301 = ~n3374 & ~n54300;
  assign n54302 = ~n51502 & ~n54190;
  assign n54303 = n3476 & ~n54302;
  assign n54304 = ~n54185 & ~n54303;
  assign n54305 = n3374 & ~n54304;
  assign n54306 = ~n54301 & ~n54305;
  assign n54307 = n3655 & ~n54306;
  assign n54308 = ~n8689 & ~n54199;
  assign n54309 = n3476 & ~n54308;
  assign n54310 = ~n54201 & ~n54309;
  assign n54311 = ~n3374 & ~n54310;
  assign n54312 = ~n51513 & ~n54215;
  assign n54313 = n3476 & ~n54312;
  assign n54314 = ~n54210 & ~n54313;
  assign n54315 = n3374 & ~n54314;
  assign n54316 = ~n54311 & ~n54315;
  assign n54317 = ~n3655 & ~n54316;
  assign n54318 = ~n54307 & ~n54317;
  assign n54319 = ~n3652 & ~n54318;
  assign n54320 = ~n54297 & ~n54319;
  assign n54321 = n3368 & ~n54320;
  assign n54322 = ~n54275 & ~n54321;
  assign n54323 = n3362 & ~n54322;
  assign n54324 = n3378 & ~n53572;
  assign n54325 = ~n51532 & ~n54324;
  assign n54326 = n3492 & ~n54325;
  assign n54327 = ~n3631 & ~n54326;
  assign n54328 = n3485 & ~n54327;
  assign n54329 = ~n3630 & ~n54328;
  assign n54330 = ~n3476 & ~n54329;
  assign n54331 = ~n51148 & ~n54326;
  assign n54332 = n3485 & ~n54331;
  assign n54333 = ~n51424 & ~n54332;
  assign n54334 = n3476 & ~n54333;
  assign n54335 = ~n54330 & ~n54334;
  assign n54336 = ~n3374 & ~n54335;
  assign n54337 = n3378 & ~n53590;
  assign n54338 = ~n51551 & ~n54337;
  assign n54339 = n3492 & ~n54338;
  assign n54340 = ~n3631 & ~n54339;
  assign n54341 = n3485 & ~n54340;
  assign n54342 = ~n3630 & ~n54341;
  assign n54343 = ~n3476 & ~n54342;
  assign n54344 = n3378 & ~n53608;
  assign n54345 = ~n51564 & ~n54344;
  assign n54346 = n3492 & ~n54345;
  assign n54347 = ~n51148 & ~n54346;
  assign n54348 = n3485 & ~n54347;
  assign n54349 = ~n51424 & ~n54348;
  assign n54350 = n3476 & ~n54349;
  assign n54351 = ~n54343 & ~n54350;
  assign n54352 = n3374 & ~n54351;
  assign n54353 = ~n54336 & ~n54352;
  assign n54354 = n3655 & ~n54353;
  assign n54355 = n3378 & ~n53624;
  assign n54356 = ~n51581 & ~n54355;
  assign n54357 = n3492 & ~n54356;
  assign n54358 = ~n3631 & ~n54357;
  assign n54359 = n3485 & ~n54358;
  assign n54360 = ~n3630 & ~n54359;
  assign n54361 = ~n3476 & ~n54360;
  assign n54362 = ~n51191 & ~n54357;
  assign n54363 = n3485 & ~n54362;
  assign n54364 = ~n51435 & ~n54363;
  assign n54365 = n3476 & ~n54364;
  assign n54366 = ~n54361 & ~n54365;
  assign n54367 = ~n3374 & ~n54366;
  assign n54368 = n3378 & ~n53642;
  assign n54369 = ~n51600 & ~n54368;
  assign n54370 = n3492 & ~n54369;
  assign n54371 = ~n3631 & ~n54370;
  assign n54372 = n3485 & ~n54371;
  assign n54373 = ~n3630 & ~n54372;
  assign n54374 = ~n3476 & ~n54373;
  assign n54375 = n3378 & ~n53660;
  assign n54376 = ~n51613 & ~n54375;
  assign n54377 = n3492 & ~n54376;
  assign n54378 = ~n51191 & ~n54377;
  assign n54379 = n3485 & ~n54378;
  assign n54380 = ~n51435 & ~n54379;
  assign n54381 = n3476 & ~n54380;
  assign n54382 = ~n54374 & ~n54381;
  assign n54383 = n3374 & ~n54382;
  assign n54384 = ~n54367 & ~n54383;
  assign n54385 = ~n3655 & ~n54384;
  assign n54386 = ~n54354 & ~n54385;
  assign n54387 = n3652 & ~n54386;
  assign n54388 = n3378 & ~n53678;
  assign n54389 = ~n51632 & ~n54388;
  assign n54390 = n3492 & ~n54389;
  assign n54391 = ~n3631 & ~n54390;
  assign n54392 = n3485 & ~n54391;
  assign n54393 = ~n3630 & ~n54392;
  assign n54394 = ~n3476 & ~n54393;
  assign n54395 = ~n51236 & ~n54390;
  assign n54396 = n3485 & ~n54395;
  assign n54397 = ~n51448 & ~n54396;
  assign n54398 = n3476 & ~n54397;
  assign n54399 = ~n54394 & ~n54398;
  assign n54400 = ~n3374 & ~n54399;
  assign n54401 = n3378 & ~n53702;
  assign n54402 = ~n51651 & ~n54401;
  assign n54403 = n3492 & ~n54402;
  assign n54404 = ~n3631 & ~n54403;
  assign n54405 = n3485 & ~n54404;
  assign n54406 = ~n3630 & ~n54405;
  assign n54407 = ~n3476 & ~n54406;
  assign n54408 = n3378 & ~n53720;
  assign n54409 = ~n51664 & ~n54408;
  assign n54410 = n3492 & ~n54409;
  assign n54411 = ~n51236 & ~n54410;
  assign n54412 = n3485 & ~n54411;
  assign n54413 = ~n51448 & ~n54412;
  assign n54414 = n3476 & ~n54413;
  assign n54415 = ~n54407 & ~n54414;
  assign n54416 = n3374 & ~n54415;
  assign n54417 = ~n54400 & ~n54416;
  assign n54418 = n3655 & ~n54417;
  assign n54419 = n3378 & ~n53736;
  assign n54420 = ~n51681 & ~n54419;
  assign n54421 = n3492 & ~n54420;
  assign n54422 = ~n3631 & ~n54421;
  assign n54423 = n3485 & ~n54422;
  assign n54424 = ~n3630 & ~n54423;
  assign n54425 = ~n3476 & ~n54424;
  assign n54426 = ~n51279 & ~n54421;
  assign n54427 = n3485 & ~n54426;
  assign n54428 = ~n51459 & ~n54427;
  assign n54429 = n3476 & ~n54428;
  assign n54430 = ~n54425 & ~n54429;
  assign n54431 = ~n3374 & ~n54430;
  assign n54432 = n3378 & ~n53760;
  assign n54433 = ~n51700 & ~n54432;
  assign n54434 = n3492 & ~n54433;
  assign n54435 = ~n3631 & ~n54434;
  assign n54436 = n3485 & ~n54435;
  assign n54437 = ~n3630 & ~n54436;
  assign n54438 = ~n3476 & ~n54437;
  assign n54439 = n3378 & ~n53778;
  assign n54440 = ~n51713 & ~n54439;
  assign n54441 = n3492 & ~n54440;
  assign n54442 = ~n51279 & ~n54441;
  assign n54443 = n3485 & ~n54442;
  assign n54444 = ~n51459 & ~n54443;
  assign n54445 = n3476 & ~n54444;
  assign n54446 = ~n54438 & ~n54445;
  assign n54447 = n3374 & ~n54446;
  assign n54448 = ~n54431 & ~n54447;
  assign n54449 = ~n3655 & ~n54448;
  assign n54450 = ~n54418 & ~n54449;
  assign n54451 = ~n3652 & ~n54450;
  assign n54452 = ~n54387 & ~n54451;
  assign n54453 = ~n3368 & ~n54452;
  assign n54454 = n3378 & ~n53798;
  assign n54455 = ~n51734 & ~n54454;
  assign n54456 = n3492 & ~n54455;
  assign n54457 = n3492 & ~n54456;
  assign n54458 = n3485 & ~n54457;
  assign n54459 = n3485 & ~n54458;
  assign n54460 = ~n3476 & ~n54459;
  assign n54461 = ~n8523 & ~n54456;
  assign n54462 = n3485 & ~n54461;
  assign n54463 = ~n8689 & ~n54462;
  assign n54464 = n3476 & ~n54463;
  assign n54465 = ~n54460 & ~n54464;
  assign n54466 = ~n3374 & ~n54465;
  assign n54467 = n3378 & ~n53816;
  assign n54468 = ~n51753 & ~n54467;
  assign n54469 = n3492 & ~n54468;
  assign n54470 = n3492 & ~n54469;
  assign n54471 = n3485 & ~n54470;
  assign n54472 = n3485 & ~n54471;
  assign n54473 = ~n3476 & ~n54472;
  assign n54474 = ~n30177 & ~n44092;
  assign n54475 = controllable_nhgrant0 & ~n54474;
  assign n54476 = ~n16962 & ~n54475;
  assign n54477 = ~n3281 & ~n54476;
  assign n54478 = ~n3281 & ~n54477;
  assign n54479 = n3378 & ~n54478;
  assign n54480 = ~n51771 & ~n54479;
  assign n54481 = n3492 & ~n54480;
  assign n54482 = ~n51321 & ~n54481;
  assign n54483 = n3485 & ~n54482;
  assign n54484 = ~n51478 & ~n54483;
  assign n54485 = n3476 & ~n54484;
  assign n54486 = ~n54473 & ~n54485;
  assign n54487 = n3374 & ~n54486;
  assign n54488 = ~n54466 & ~n54487;
  assign n54489 = n3655 & ~n54488;
  assign n54490 = n3378 & ~n53850;
  assign n54491 = ~n51788 & ~n54490;
  assign n54492 = n3492 & ~n54491;
  assign n54493 = n3492 & ~n54492;
  assign n54494 = n3485 & ~n54493;
  assign n54495 = n3485 & ~n54494;
  assign n54496 = ~n3476 & ~n54495;
  assign n54497 = ~n8523 & ~n54492;
  assign n54498 = n3485 & ~n54497;
  assign n54499 = ~n8689 & ~n54498;
  assign n54500 = n3476 & ~n54499;
  assign n54501 = ~n54496 & ~n54500;
  assign n54502 = ~n3374 & ~n54501;
  assign n54503 = n3378 & ~n53868;
  assign n54504 = ~n51807 & ~n54503;
  assign n54505 = n3492 & ~n54504;
  assign n54506 = n3492 & ~n54505;
  assign n54507 = n3485 & ~n54506;
  assign n54508 = n3485 & ~n54507;
  assign n54509 = ~n3476 & ~n54508;
  assign n54510 = ~n30177 & ~n44149;
  assign n54511 = controllable_nhgrant0 & ~n54510;
  assign n54512 = ~n16962 & ~n54511;
  assign n54513 = ~n3281 & ~n54512;
  assign n54514 = ~n3281 & ~n54513;
  assign n54515 = n3378 & ~n54514;
  assign n54516 = ~n51825 & ~n54515;
  assign n54517 = n3492 & ~n54516;
  assign n54518 = ~n51348 & ~n54517;
  assign n54519 = n3485 & ~n54518;
  assign n54520 = ~n51489 & ~n54519;
  assign n54521 = n3476 & ~n54520;
  assign n54522 = ~n54509 & ~n54521;
  assign n54523 = n3374 & ~n54522;
  assign n54524 = ~n54502 & ~n54523;
  assign n54525 = ~n3655 & ~n54524;
  assign n54526 = ~n54489 & ~n54525;
  assign n54527 = n3652 & ~n54526;
  assign n54528 = n3378 & ~n53904;
  assign n54529 = ~n51844 & ~n54528;
  assign n54530 = n3492 & ~n54529;
  assign n54531 = n3492 & ~n54530;
  assign n54532 = n3485 & ~n54531;
  assign n54533 = n3485 & ~n54532;
  assign n54534 = ~n3476 & ~n54533;
  assign n54535 = ~n8523 & ~n54530;
  assign n54536 = n3485 & ~n54535;
  assign n54537 = ~n8689 & ~n54536;
  assign n54538 = n3476 & ~n54537;
  assign n54539 = ~n54534 & ~n54538;
  assign n54540 = ~n3374 & ~n54539;
  assign n54541 = n3378 & ~n53922;
  assign n54542 = ~n51863 & ~n54541;
  assign n54543 = n3492 & ~n54542;
  assign n54544 = n3492 & ~n54543;
  assign n54545 = n3485 & ~n54544;
  assign n54546 = n3485 & ~n54545;
  assign n54547 = ~n3476 & ~n54546;
  assign n54548 = ~n30177 & ~n44236;
  assign n54549 = controllable_nhgrant0 & ~n54548;
  assign n54550 = ~n16962 & ~n54549;
  assign n54551 = ~n3281 & ~n54550;
  assign n54552 = ~n3281 & ~n54551;
  assign n54553 = n3378 & ~n54552;
  assign n54554 = ~n51881 & ~n54553;
  assign n54555 = n3492 & ~n54554;
  assign n54556 = ~n51377 & ~n54555;
  assign n54557 = n3485 & ~n54556;
  assign n54558 = ~n51502 & ~n54557;
  assign n54559 = n3476 & ~n54558;
  assign n54560 = ~n54547 & ~n54559;
  assign n54561 = n3374 & ~n54560;
  assign n54562 = ~n54540 & ~n54561;
  assign n54563 = n3655 & ~n54562;
  assign n54564 = n3378 & ~n53956;
  assign n54565 = ~n51898 & ~n54564;
  assign n54566 = n3492 & ~n54565;
  assign n54567 = n3492 & ~n54566;
  assign n54568 = n3485 & ~n54567;
  assign n54569 = n3485 & ~n54568;
  assign n54570 = ~n3476 & ~n54569;
  assign n54571 = ~n8523 & ~n54566;
  assign n54572 = n3485 & ~n54571;
  assign n54573 = ~n8689 & ~n54572;
  assign n54574 = n3476 & ~n54573;
  assign n54575 = ~n54570 & ~n54574;
  assign n54576 = ~n3374 & ~n54575;
  assign n54577 = n3378 & ~n53974;
  assign n54578 = ~n51917 & ~n54577;
  assign n54579 = n3492 & ~n54578;
  assign n54580 = n3492 & ~n54579;
  assign n54581 = n3485 & ~n54580;
  assign n54582 = n3485 & ~n54581;
  assign n54583 = ~n3476 & ~n54582;
  assign n54584 = ~n30177 & ~n44321;
  assign n54585 = controllable_nhgrant0 & ~n54584;
  assign n54586 = ~n16962 & ~n54585;
  assign n54587 = ~n3281 & ~n54586;
  assign n54588 = ~n3281 & ~n54587;
  assign n54589 = n3378 & ~n54588;
  assign n54590 = ~n51935 & ~n54589;
  assign n54591 = n3492 & ~n54590;
  assign n54592 = ~n51404 & ~n54591;
  assign n54593 = n3485 & ~n54592;
  assign n54594 = ~n51513 & ~n54593;
  assign n54595 = n3476 & ~n54594;
  assign n54596 = ~n54583 & ~n54595;
  assign n54597 = n3374 & ~n54596;
  assign n54598 = ~n54576 & ~n54597;
  assign n54599 = ~n3655 & ~n54598;
  assign n54600 = ~n54563 & ~n54599;
  assign n54601 = ~n3652 & ~n54600;
  assign n54602 = ~n54527 & ~n54601;
  assign n54603 = n3368 & ~n54602;
  assign n54604 = ~n54453 & ~n54603;
  assign n54605 = ~n3362 & ~n54604;
  assign n54606 = ~n54323 & ~n54605;
  assign n54607 = ~n3359 & ~n54606;
  assign n54608 = ~n54229 & ~n54607;
  assign n54609 = ~n3356 & ~n54608;
  assign n54610 = ~n53567 & ~n54609;
  assign n54611 = n3345 & ~n54610;
  assign n54612 = ~n53293 & ~n54611;
  assign n54613 = n3341 & ~n54612;
  assign n54614 = ~n51959 & ~n54613;
  assign n54615 = ~n3337 & ~n54614;
  assign n54616 = ~n30307 & ~n44365;
  assign n54617 = controllable_nhgrant0 & ~n54616;
  assign n54618 = ~n17300 & ~n54617;
  assign n54619 = ~n3281 & ~n54618;
  assign n54620 = ~n3281 & ~n54619;
  assign n54621 = n3378 & ~n54620;
  assign n54622 = ~n30314 & ~n44373;
  assign n54623 = controllable_nhgrant0 & ~n54622;
  assign n54624 = ~n17314 & ~n54623;
  assign n54625 = ~n3281 & ~n54624;
  assign n54626 = ~n3950 & ~n54625;
  assign n54627 = ~n3378 & ~n54626;
  assign n54628 = ~n54621 & ~n54627;
  assign n54629 = n3492 & ~n54628;
  assign n54630 = ~n3493 & ~n54629;
  assign n54631 = n3485 & ~n54630;
  assign n54632 = ~n3486 & ~n54631;
  assign n54633 = ~n3476 & ~n54632;
  assign n54634 = ~n30307 & ~n44408;
  assign n54635 = controllable_nhgrant0 & ~n54634;
  assign n54636 = ~n17300 & ~n54635;
  assign n54637 = ~n3281 & ~n54636;
  assign n54638 = ~n3281 & ~n54637;
  assign n54639 = n3378 & ~n54638;
  assign n54640 = ~n30314 & ~n44437;
  assign n54641 = controllable_nhgrant0 & ~n54640;
  assign n54642 = ~n17314 & ~n54641;
  assign n54643 = ~n3281 & ~n54642;
  assign n54644 = ~n4089 & ~n54643;
  assign n54645 = ~n3378 & ~n54644;
  assign n54646 = ~n54639 & ~n54645;
  assign n54647 = n3492 & ~n54646;
  assign n54648 = ~n3493 & ~n54647;
  assign n54649 = n3485 & ~n54648;
  assign n54650 = ~n3486 & ~n54649;
  assign n54651 = n3476 & ~n54650;
  assign n54652 = ~n54633 & ~n54651;
  assign n54653 = n3374 & ~n54652;
  assign n54654 = ~n17268 & ~n54653;
  assign n54655 = n3655 & ~n54654;
  assign n54656 = ~n30307 & ~n44465;
  assign n54657 = controllable_nhgrant0 & ~n54656;
  assign n54658 = ~n17300 & ~n54657;
  assign n54659 = ~n3281 & ~n54658;
  assign n54660 = ~n3281 & ~n54659;
  assign n54661 = n3378 & ~n54660;
  assign n54662 = ~n30314 & ~n44473;
  assign n54663 = controllable_nhgrant0 & ~n54662;
  assign n54664 = ~n17314 & ~n54663;
  assign n54665 = ~n3281 & ~n54664;
  assign n54666 = ~n3950 & ~n54665;
  assign n54667 = ~n3378 & ~n54666;
  assign n54668 = ~n54661 & ~n54667;
  assign n54669 = n3492 & ~n54668;
  assign n54670 = ~n3493 & ~n54669;
  assign n54671 = n3485 & ~n54670;
  assign n54672 = ~n3486 & ~n54671;
  assign n54673 = ~n3476 & ~n54672;
  assign n54674 = ~n30307 & ~n44508;
  assign n54675 = controllable_nhgrant0 & ~n54674;
  assign n54676 = ~n17300 & ~n54675;
  assign n54677 = ~n3281 & ~n54676;
  assign n54678 = ~n3281 & ~n54677;
  assign n54679 = n3378 & ~n54678;
  assign n54680 = ~n30314 & ~n44537;
  assign n54681 = controllable_nhgrant0 & ~n54680;
  assign n54682 = ~n17314 & ~n54681;
  assign n54683 = ~n3281 & ~n54682;
  assign n54684 = ~n4089 & ~n54683;
  assign n54685 = ~n3378 & ~n54684;
  assign n54686 = ~n54679 & ~n54685;
  assign n54687 = n3492 & ~n54686;
  assign n54688 = ~n17612 & ~n54687;
  assign n54689 = n3485 & ~n54688;
  assign n54690 = ~n17611 & ~n54689;
  assign n54691 = n3476 & ~n54690;
  assign n54692 = ~n54673 & ~n54691;
  assign n54693 = n3374 & ~n54692;
  assign n54694 = ~n17618 & ~n54693;
  assign n54695 = ~n3655 & ~n54694;
  assign n54696 = ~n54655 & ~n54695;
  assign n54697 = n3652 & ~n54696;
  assign n54698 = ~n30307 & ~n44567;
  assign n54699 = controllable_nhgrant0 & ~n54698;
  assign n54700 = ~n17300 & ~n54699;
  assign n54701 = ~n3281 & ~n54700;
  assign n54702 = ~n3281 & ~n54701;
  assign n54703 = n3378 & ~n54702;
  assign n54704 = ~n30314 & ~n44575;
  assign n54705 = controllable_nhgrant0 & ~n54704;
  assign n54706 = ~n17314 & ~n54705;
  assign n54707 = ~n3281 & ~n54706;
  assign n54708 = ~n3950 & ~n54707;
  assign n54709 = ~n3378 & ~n54708;
  assign n54710 = ~n54703 & ~n54709;
  assign n54711 = n3492 & ~n54710;
  assign n54712 = ~n3493 & ~n54711;
  assign n54713 = n3485 & ~n54712;
  assign n54714 = ~n3486 & ~n54713;
  assign n54715 = ~n3476 & ~n54714;
  assign n54716 = ~n30307 & ~n44603;
  assign n54717 = controllable_nhgrant0 & ~n54716;
  assign n54718 = ~n17300 & ~n54717;
  assign n54719 = ~n3281 & ~n54718;
  assign n54720 = ~n3281 & ~n54719;
  assign n54721 = n3378 & ~n54720;
  assign n54722 = ~n30314 & ~n44625;
  assign n54723 = controllable_nhgrant0 & ~n54722;
  assign n54724 = ~n17314 & ~n54723;
  assign n54725 = ~n3281 & ~n54724;
  assign n54726 = ~n4089 & ~n54725;
  assign n54727 = ~n3378 & ~n54726;
  assign n54728 = ~n54721 & ~n54727;
  assign n54729 = n3492 & ~n54728;
  assign n54730 = ~n3493 & ~n54729;
  assign n54731 = n3485 & ~n54730;
  assign n54732 = ~n3486 & ~n54731;
  assign n54733 = n3476 & ~n54732;
  assign n54734 = ~n54715 & ~n54733;
  assign n54735 = n3374 & ~n54734;
  assign n54736 = ~n17268 & ~n54735;
  assign n54737 = n3655 & ~n54736;
  assign n54738 = ~n30307 & ~n44653;
  assign n54739 = controllable_nhgrant0 & ~n54738;
  assign n54740 = ~n17300 & ~n54739;
  assign n54741 = ~n3281 & ~n54740;
  assign n54742 = ~n3281 & ~n54741;
  assign n54743 = n3378 & ~n54742;
  assign n54744 = ~n30314 & ~n44661;
  assign n54745 = controllable_nhgrant0 & ~n54744;
  assign n54746 = ~n17314 & ~n54745;
  assign n54747 = ~n3281 & ~n54746;
  assign n54748 = ~n3950 & ~n54747;
  assign n54749 = ~n3378 & ~n54748;
  assign n54750 = ~n54743 & ~n54749;
  assign n54751 = n3492 & ~n54750;
  assign n54752 = ~n3493 & ~n54751;
  assign n54753 = n3485 & ~n54752;
  assign n54754 = ~n3486 & ~n54753;
  assign n54755 = ~n3476 & ~n54754;
  assign n54756 = ~n30307 & ~n44689;
  assign n54757 = controllable_nhgrant0 & ~n54756;
  assign n54758 = ~n17300 & ~n54757;
  assign n54759 = ~n3281 & ~n54758;
  assign n54760 = ~n3281 & ~n54759;
  assign n54761 = n3378 & ~n54760;
  assign n54762 = ~n30314 & ~n44711;
  assign n54763 = controllable_nhgrant0 & ~n54762;
  assign n54764 = ~n17314 & ~n54763;
  assign n54765 = ~n3281 & ~n54764;
  assign n54766 = ~n4089 & ~n54765;
  assign n54767 = ~n3378 & ~n54766;
  assign n54768 = ~n54761 & ~n54767;
  assign n54769 = n3492 & ~n54768;
  assign n54770 = ~n17612 & ~n54769;
  assign n54771 = n3485 & ~n54770;
  assign n54772 = ~n17611 & ~n54771;
  assign n54773 = n3476 & ~n54772;
  assign n54774 = ~n54755 & ~n54773;
  assign n54775 = n3374 & ~n54774;
  assign n54776 = ~n17618 & ~n54775;
  assign n54777 = ~n3655 & ~n54776;
  assign n54778 = ~n54737 & ~n54777;
  assign n54779 = ~n3652 & ~n54778;
  assign n54780 = ~n54697 & ~n54779;
  assign n54781 = ~n3368 & ~n54780;
  assign n54782 = ~n30475 & ~n44743;
  assign n54783 = controllable_nhgrant0 & ~n54782;
  assign n54784 = ~n18077 & ~n54783;
  assign n54785 = ~n3281 & ~n54784;
  assign n54786 = ~n3281 & ~n54785;
  assign n54787 = n3492 & ~n54786;
  assign n54788 = n3492 & ~n54787;
  assign n54789 = n3485 & ~n54788;
  assign n54790 = n3485 & ~n54789;
  assign n54791 = ~n3476 & ~n54790;
  assign n54792 = ~n30475 & ~n44776;
  assign n54793 = controllable_nhgrant0 & ~n54792;
  assign n54794 = ~n18077 & ~n54793;
  assign n54795 = ~n3281 & ~n54794;
  assign n54796 = ~n3281 & ~n54795;
  assign n54797 = n3492 & ~n54796;
  assign n54798 = n3492 & ~n54797;
  assign n54799 = n3485 & ~n54798;
  assign n54800 = n3485 & ~n54799;
  assign n54801 = n3476 & ~n54800;
  assign n54802 = ~n54791 & ~n54801;
  assign n54803 = n3374 & ~n54802;
  assign n54804 = n3374 & ~n54803;
  assign n54805 = n3655 & ~n54804;
  assign n54806 = ~n30475 & ~n44802;
  assign n54807 = controllable_nhgrant0 & ~n54806;
  assign n54808 = ~n18077 & ~n54807;
  assign n54809 = ~n3281 & ~n54808;
  assign n54810 = ~n3281 & ~n54809;
  assign n54811 = n3492 & ~n54810;
  assign n54812 = n3492 & ~n54811;
  assign n54813 = n3485 & ~n54812;
  assign n54814 = n3485 & ~n54813;
  assign n54815 = ~n3476 & ~n54814;
  assign n54816 = ~n30475 & ~n44835;
  assign n54817 = controllable_nhgrant0 & ~n54816;
  assign n54818 = ~n18077 & ~n54817;
  assign n54819 = ~n3281 & ~n54818;
  assign n54820 = ~n3281 & ~n54819;
  assign n54821 = n3492 & ~n54820;
  assign n54822 = ~n18151 & ~n54821;
  assign n54823 = n3485 & ~n54822;
  assign n54824 = ~n18150 & ~n54823;
  assign n54825 = n3476 & ~n54824;
  assign n54826 = ~n54815 & ~n54825;
  assign n54827 = n3374 & ~n54826;
  assign n54828 = n3374 & ~n54827;
  assign n54829 = ~n3655 & ~n54828;
  assign n54830 = ~n54805 & ~n54829;
  assign n54831 = n3652 & ~n54830;
  assign n54832 = ~n30475 & ~n44863;
  assign n54833 = controllable_nhgrant0 & ~n54832;
  assign n54834 = ~n18077 & ~n54833;
  assign n54835 = ~n3281 & ~n54834;
  assign n54836 = ~n3281 & ~n54835;
  assign n54837 = n3492 & ~n54836;
  assign n54838 = n3492 & ~n54837;
  assign n54839 = n3485 & ~n54838;
  assign n54840 = n3485 & ~n54839;
  assign n54841 = ~n3476 & ~n54840;
  assign n54842 = ~n30475 & ~n44889;
  assign n54843 = controllable_nhgrant0 & ~n54842;
  assign n54844 = ~n18077 & ~n54843;
  assign n54845 = ~n3281 & ~n54844;
  assign n54846 = ~n3281 & ~n54845;
  assign n54847 = n3492 & ~n54846;
  assign n54848 = n3492 & ~n54847;
  assign n54849 = n3485 & ~n54848;
  assign n54850 = n3485 & ~n54849;
  assign n54851 = n3476 & ~n54850;
  assign n54852 = ~n54841 & ~n54851;
  assign n54853 = n3374 & ~n54852;
  assign n54854 = n3374 & ~n54853;
  assign n54855 = n3655 & ~n54854;
  assign n54856 = ~n30475 & ~n44915;
  assign n54857 = controllable_nhgrant0 & ~n54856;
  assign n54858 = ~n18077 & ~n54857;
  assign n54859 = ~n3281 & ~n54858;
  assign n54860 = ~n3281 & ~n54859;
  assign n54861 = n3492 & ~n54860;
  assign n54862 = n3492 & ~n54861;
  assign n54863 = n3485 & ~n54862;
  assign n54864 = n3485 & ~n54863;
  assign n54865 = ~n3476 & ~n54864;
  assign n54866 = ~n30475 & ~n44941;
  assign n54867 = controllable_nhgrant0 & ~n54866;
  assign n54868 = ~n18077 & ~n54867;
  assign n54869 = ~n3281 & ~n54868;
  assign n54870 = ~n3281 & ~n54869;
  assign n54871 = n3492 & ~n54870;
  assign n54872 = ~n18151 & ~n54871;
  assign n54873 = n3485 & ~n54872;
  assign n54874 = ~n18150 & ~n54873;
  assign n54875 = n3476 & ~n54874;
  assign n54876 = ~n54865 & ~n54875;
  assign n54877 = n3374 & ~n54876;
  assign n54878 = n3374 & ~n54877;
  assign n54879 = ~n3655 & ~n54878;
  assign n54880 = ~n54855 & ~n54879;
  assign n54881 = ~n3652 & ~n54880;
  assign n54882 = ~n54831 & ~n54881;
  assign n54883 = n3368 & ~n54882;
  assign n54884 = ~n54781 & ~n54883;
  assign n54885 = ~n3362 & ~n54884;
  assign n54886 = ~n3362 & ~n54885;
  assign n54887 = ~n3359 & ~n54886;
  assign n54888 = ~n3359 & ~n54887;
  assign n54889 = n3356 & ~n54888;
  assign n54890 = ~n18369 & ~n53573;
  assign n54891 = n3492 & ~n54890;
  assign n54892 = ~n3631 & ~n54891;
  assign n54893 = n3485 & ~n54892;
  assign n54894 = ~n3630 & ~n54893;
  assign n54895 = ~n3374 & ~n54894;
  assign n54896 = ~n30599 & ~n44983;
  assign n54897 = controllable_nhgrant0 & ~n54896;
  assign n54898 = ~n18416 & ~n54897;
  assign n54899 = ~n3281 & ~n54898;
  assign n54900 = ~n3950 & ~n54899;
  assign n54901 = n3378 & ~n54900;
  assign n54902 = ~n25684 & ~n45001;
  assign n54903 = controllable_nhgrant0 & ~n54902;
  assign n54904 = ~n5534 & ~n54903;
  assign n54905 = ~n3281 & ~n54904;
  assign n54906 = ~n3950 & ~n54905;
  assign n54907 = ~n3378 & ~n54906;
  assign n54908 = ~n54901 & ~n54907;
  assign n54909 = n3492 & ~n54908;
  assign n54910 = ~n3631 & ~n54909;
  assign n54911 = n3485 & ~n54910;
  assign n54912 = ~n3630 & ~n54911;
  assign n54913 = ~n3476 & ~n54912;
  assign n54914 = ~n30627 & ~n45036;
  assign n54915 = controllable_nhgrant0 & ~n54914;
  assign n54916 = ~n18526 & ~n54915;
  assign n54917 = ~n3281 & ~n54916;
  assign n54918 = ~n4089 & ~n54917;
  assign n54919 = n3378 & ~n54918;
  assign n54920 = ~n25726 & ~n45060;
  assign n54921 = controllable_nhgrant0 & ~n54920;
  assign n54922 = ~n6082 & ~n54921;
  assign n54923 = ~n3281 & ~n54922;
  assign n54924 = ~n4089 & ~n54923;
  assign n54925 = ~n3378 & ~n54924;
  assign n54926 = ~n54919 & ~n54925;
  assign n54927 = n3492 & ~n54926;
  assign n54928 = ~n3631 & ~n54927;
  assign n54929 = n3485 & ~n54928;
  assign n54930 = ~n3630 & ~n54929;
  assign n54931 = n3476 & ~n54930;
  assign n54932 = ~n54913 & ~n54931;
  assign n54933 = n3374 & ~n54932;
  assign n54934 = ~n54895 & ~n54933;
  assign n54935 = n3655 & ~n54934;
  assign n54936 = ~n25649 & ~n45101;
  assign n54937 = controllable_nhgrant0 & ~n54936;
  assign n54938 = ~n5245 & ~n54937;
  assign n54939 = ~n3281 & ~n54938;
  assign n54940 = ~n3783 & ~n54939;
  assign n54941 = ~n3378 & ~n54940;
  assign n54942 = ~n18571 & ~n54941;
  assign n54943 = n3492 & ~n54942;
  assign n54944 = ~n3631 & ~n54943;
  assign n54945 = n3485 & ~n54944;
  assign n54946 = ~n3630 & ~n54945;
  assign n54947 = ~n3476 & ~n54946;
  assign n54948 = ~n18630 & ~n54943;
  assign n54949 = n3485 & ~n54948;
  assign n54950 = ~n18629 & ~n54949;
  assign n54951 = n3476 & ~n54950;
  assign n54952 = ~n54947 & ~n54951;
  assign n54953 = ~n3374 & ~n54952;
  assign n54954 = ~n30599 & ~n45131;
  assign n54955 = controllable_nhgrant0 & ~n54954;
  assign n54956 = ~n18416 & ~n54955;
  assign n54957 = ~n3281 & ~n54956;
  assign n54958 = ~n3950 & ~n54957;
  assign n54959 = n3378 & ~n54958;
  assign n54960 = ~n25684 & ~n45172;
  assign n54961 = controllable_nhgrant0 & ~n54960;
  assign n54962 = ~n5534 & ~n54961;
  assign n54963 = ~n3281 & ~n54962;
  assign n54964 = ~n3950 & ~n54963;
  assign n54965 = ~n3378 & ~n54964;
  assign n54966 = ~n54959 & ~n54965;
  assign n54967 = n3492 & ~n54966;
  assign n54968 = ~n3631 & ~n54967;
  assign n54969 = n3485 & ~n54968;
  assign n54970 = ~n3630 & ~n54969;
  assign n54971 = ~n3476 & ~n54970;
  assign n54972 = ~n30627 & ~n45207;
  assign n54973 = controllable_nhgrant0 & ~n54972;
  assign n54974 = ~n18526 & ~n54973;
  assign n54975 = ~n3281 & ~n54974;
  assign n54976 = ~n4089 & ~n54975;
  assign n54977 = n3378 & ~n54976;
  assign n54978 = ~n25726 & ~n45254;
  assign n54979 = controllable_nhgrant0 & ~n54978;
  assign n54980 = ~n6082 & ~n54979;
  assign n54981 = ~n3281 & ~n54980;
  assign n54982 = ~n4089 & ~n54981;
  assign n54983 = ~n3378 & ~n54982;
  assign n54984 = ~n54977 & ~n54983;
  assign n54985 = n3492 & ~n54984;
  assign n54986 = ~n18630 & ~n54985;
  assign n54987 = n3485 & ~n54986;
  assign n54988 = ~n18629 & ~n54987;
  assign n54989 = n3476 & ~n54988;
  assign n54990 = ~n54971 & ~n54989;
  assign n54991 = n3374 & ~n54990;
  assign n54992 = ~n54953 & ~n54991;
  assign n54993 = ~n3655 & ~n54992;
  assign n54994 = ~n54935 & ~n54993;
  assign n54995 = n3652 & ~n54994;
  assign n54996 = ~n25649 & ~n39991;
  assign n54997 = controllable_nhgrant0 & ~n54996;
  assign n54998 = ~n5245 & ~n54997;
  assign n54999 = ~n3281 & ~n54998;
  assign n55000 = ~n3783 & ~n54999;
  assign n55001 = ~n3378 & ~n55000;
  assign n55002 = ~n18369 & ~n55001;
  assign n55003 = n3492 & ~n55002;
  assign n55004 = ~n3631 & ~n55003;
  assign n55005 = n3485 & ~n55004;
  assign n55006 = ~n3630 & ~n55005;
  assign n55007 = ~n3374 & ~n55006;
  assign n55008 = ~n30599 & ~n45290;
  assign n55009 = controllable_nhgrant0 & ~n55008;
  assign n55010 = ~n18416 & ~n55009;
  assign n55011 = ~n3281 & ~n55010;
  assign n55012 = ~n3950 & ~n55011;
  assign n55013 = n3378 & ~n55012;
  assign n55014 = ~n25684 & ~n45308;
  assign n55015 = controllable_nhgrant0 & ~n55014;
  assign n55016 = ~n5534 & ~n55015;
  assign n55017 = ~n3281 & ~n55016;
  assign n55018 = ~n3950 & ~n55017;
  assign n55019 = ~n3378 & ~n55018;
  assign n55020 = ~n55013 & ~n55019;
  assign n55021 = n3492 & ~n55020;
  assign n55022 = ~n3631 & ~n55021;
  assign n55023 = n3485 & ~n55022;
  assign n55024 = ~n3630 & ~n55023;
  assign n55025 = ~n3476 & ~n55024;
  assign n55026 = ~n30627 & ~n45336;
  assign n55027 = controllable_nhgrant0 & ~n55026;
  assign n55028 = ~n18526 & ~n55027;
  assign n55029 = ~n3281 & ~n55028;
  assign n55030 = ~n4089 & ~n55029;
  assign n55031 = n3378 & ~n55030;
  assign n55032 = ~n25726 & ~n45356;
  assign n55033 = controllable_nhgrant0 & ~n55032;
  assign n55034 = ~n6082 & ~n55033;
  assign n55035 = ~n3281 & ~n55034;
  assign n55036 = ~n4089 & ~n55035;
  assign n55037 = ~n3378 & ~n55036;
  assign n55038 = ~n55031 & ~n55037;
  assign n55039 = n3492 & ~n55038;
  assign n55040 = ~n3631 & ~n55039;
  assign n55041 = n3485 & ~n55040;
  assign n55042 = ~n3630 & ~n55041;
  assign n55043 = n3476 & ~n55042;
  assign n55044 = ~n55025 & ~n55043;
  assign n55045 = n3374 & ~n55044;
  assign n55046 = ~n55007 & ~n55045;
  assign n55047 = n3655 & ~n55046;
  assign n55048 = ~n25649 & ~n45390;
  assign n55049 = controllable_nhgrant0 & ~n55048;
  assign n55050 = ~n5245 & ~n55049;
  assign n55051 = ~n3281 & ~n55050;
  assign n55052 = ~n3783 & ~n55051;
  assign n55053 = ~n3378 & ~n55052;
  assign n55054 = ~n18571 & ~n55053;
  assign n55055 = n3492 & ~n55054;
  assign n55056 = ~n3631 & ~n55055;
  assign n55057 = n3485 & ~n55056;
  assign n55058 = ~n3630 & ~n55057;
  assign n55059 = ~n3476 & ~n55058;
  assign n55060 = ~n18630 & ~n55055;
  assign n55061 = n3485 & ~n55060;
  assign n55062 = ~n18629 & ~n55061;
  assign n55063 = n3476 & ~n55062;
  assign n55064 = ~n55059 & ~n55063;
  assign n55065 = ~n3374 & ~n55064;
  assign n55066 = ~n30599 & ~n45420;
  assign n55067 = controllable_nhgrant0 & ~n55066;
  assign n55068 = ~n18416 & ~n55067;
  assign n55069 = ~n3281 & ~n55068;
  assign n55070 = ~n3950 & ~n55069;
  assign n55071 = n3378 & ~n55070;
  assign n55072 = ~n25684 & ~n45454;
  assign n55073 = controllable_nhgrant0 & ~n55072;
  assign n55074 = ~n5534 & ~n55073;
  assign n55075 = ~n3281 & ~n55074;
  assign n55076 = ~n3950 & ~n55075;
  assign n55077 = ~n3378 & ~n55076;
  assign n55078 = ~n55071 & ~n55077;
  assign n55079 = n3492 & ~n55078;
  assign n55080 = ~n3631 & ~n55079;
  assign n55081 = n3485 & ~n55080;
  assign n55082 = ~n3630 & ~n55081;
  assign n55083 = ~n3476 & ~n55082;
  assign n55084 = ~n30627 & ~n45482;
  assign n55085 = controllable_nhgrant0 & ~n55084;
  assign n55086 = ~n18526 & ~n55085;
  assign n55087 = ~n3281 & ~n55086;
  assign n55088 = ~n4089 & ~n55087;
  assign n55089 = n3378 & ~n55088;
  assign n55090 = ~n25726 & ~n45518;
  assign n55091 = controllable_nhgrant0 & ~n55090;
  assign n55092 = ~n6082 & ~n55091;
  assign n55093 = ~n3281 & ~n55092;
  assign n55094 = ~n4089 & ~n55093;
  assign n55095 = ~n3378 & ~n55094;
  assign n55096 = ~n55089 & ~n55095;
  assign n55097 = n3492 & ~n55096;
  assign n55098 = ~n18630 & ~n55097;
  assign n55099 = n3485 & ~n55098;
  assign n55100 = ~n18629 & ~n55099;
  assign n55101 = n3476 & ~n55100;
  assign n55102 = ~n55083 & ~n55101;
  assign n55103 = n3374 & ~n55102;
  assign n55104 = ~n55065 & ~n55103;
  assign n55105 = ~n3655 & ~n55104;
  assign n55106 = ~n55047 & ~n55105;
  assign n55107 = ~n3652 & ~n55106;
  assign n55108 = ~n54995 & ~n55107;
  assign n55109 = ~n3368 & ~n55108;
  assign n55110 = ~n30827 & ~n45550;
  assign n55111 = controllable_nhgrant0 & ~n55110;
  assign n55112 = ~n19213 & ~n55111;
  assign n55113 = ~n3281 & ~n55112;
  assign n55114 = ~n3281 & ~n55113;
  assign n55115 = n3378 & ~n55114;
  assign n55116 = ~n30844 & ~n45568;
  assign n55117 = controllable_nhgrant0 & ~n55116;
  assign n55118 = ~n19255 & ~n55117;
  assign n55119 = ~n3281 & ~n55118;
  assign n55120 = ~n3281 & ~n55119;
  assign n55121 = ~n3378 & ~n55120;
  assign n55122 = ~n55115 & ~n55121;
  assign n55123 = n3492 & ~n55122;
  assign n55124 = n3492 & ~n55123;
  assign n55125 = n3485 & ~n55124;
  assign n55126 = n3485 & ~n55125;
  assign n55127 = ~n3476 & ~n55126;
  assign n55128 = ~n30866 & ~n45603;
  assign n55129 = controllable_nhgrant0 & ~n55128;
  assign n55130 = ~n19385 & ~n55129;
  assign n55131 = ~n3281 & ~n55130;
  assign n55132 = ~n3281 & ~n55131;
  assign n55133 = n3378 & ~n55132;
  assign n55134 = ~n30883 & ~n45669;
  assign n55135 = controllable_nhgrant0 & ~n55134;
  assign n55136 = ~n19515 & ~n55135;
  assign n55137 = ~n3281 & ~n55136;
  assign n55138 = ~n3281 & ~n55137;
  assign n55139 = ~n3378 & ~n55138;
  assign n55140 = ~n55133 & ~n55139;
  assign n55141 = n3492 & ~n55140;
  assign n55142 = n3492 & ~n55141;
  assign n55143 = n3485 & ~n55142;
  assign n55144 = n3485 & ~n55143;
  assign n55145 = n3476 & ~n55144;
  assign n55146 = ~n55127 & ~n55145;
  assign n55147 = n3374 & ~n55146;
  assign n55148 = ~n53805 & ~n55147;
  assign n55149 = n3655 & ~n55148;
  assign n55150 = ~n25905 & ~n45710;
  assign n55151 = controllable_nhgrant0 & ~n55150;
  assign n55152 = ~n7118 & ~n55151;
  assign n55153 = ~n3281 & ~n55152;
  assign n55154 = ~n3281 & ~n55153;
  assign n55155 = ~n3378 & ~n55154;
  assign n55156 = ~n19575 & ~n55155;
  assign n55157 = n3492 & ~n55156;
  assign n55158 = n3492 & ~n55157;
  assign n55159 = n3485 & ~n55158;
  assign n55160 = n3485 & ~n55159;
  assign n55161 = ~n3374 & ~n55160;
  assign n55162 = ~n30827 & ~n45734;
  assign n55163 = controllable_nhgrant0 & ~n55162;
  assign n55164 = ~n19213 & ~n55163;
  assign n55165 = ~n3281 & ~n55164;
  assign n55166 = ~n3281 & ~n55165;
  assign n55167 = n3378 & ~n55166;
  assign n55168 = ~n30844 & ~n45799;
  assign n55169 = controllable_nhgrant0 & ~n55168;
  assign n55170 = ~n19255 & ~n55169;
  assign n55171 = ~n3281 & ~n55170;
  assign n55172 = ~n3281 & ~n55171;
  assign n55173 = ~n3378 & ~n55172;
  assign n55174 = ~n55167 & ~n55173;
  assign n55175 = n3492 & ~n55174;
  assign n55176 = n3492 & ~n55175;
  assign n55177 = n3485 & ~n55176;
  assign n55178 = n3485 & ~n55177;
  assign n55179 = ~n3476 & ~n55178;
  assign n55180 = ~n30866 & ~n45834;
  assign n55181 = controllable_nhgrant0 & ~n55180;
  assign n55182 = ~n19385 & ~n55181;
  assign n55183 = ~n3281 & ~n55182;
  assign n55184 = ~n3281 & ~n55183;
  assign n55185 = n3378 & ~n55184;
  assign n55186 = ~n30883 & ~n45923;
  assign n55187 = controllable_nhgrant0 & ~n55186;
  assign n55188 = ~n19515 & ~n55187;
  assign n55189 = ~n3281 & ~n55188;
  assign n55190 = ~n3281 & ~n55189;
  assign n55191 = ~n3378 & ~n55190;
  assign n55192 = ~n55185 & ~n55191;
  assign n55193 = n3492 & ~n55192;
  assign n55194 = ~n18151 & ~n55193;
  assign n55195 = n3485 & ~n55194;
  assign n55196 = ~n18150 & ~n55195;
  assign n55197 = n3476 & ~n55196;
  assign n55198 = ~n55179 & ~n55197;
  assign n55199 = n3374 & ~n55198;
  assign n55200 = ~n55161 & ~n55199;
  assign n55201 = ~n3655 & ~n55200;
  assign n55202 = ~n55149 & ~n55201;
  assign n55203 = n3652 & ~n55202;
  assign n55204 = ~n25905 & ~n40743;
  assign n55205 = controllable_nhgrant0 & ~n55204;
  assign n55206 = ~n7118 & ~n55205;
  assign n55207 = ~n3281 & ~n55206;
  assign n55208 = ~n3281 & ~n55207;
  assign n55209 = ~n3378 & ~n55208;
  assign n55210 = ~n7082 & ~n55209;
  assign n55211 = n3492 & ~n55210;
  assign n55212 = n3492 & ~n55211;
  assign n55213 = n3485 & ~n55212;
  assign n55214 = n3485 & ~n55213;
  assign n55215 = ~n3374 & ~n55214;
  assign n55216 = ~n30827 & ~n45953;
  assign n55217 = controllable_nhgrant0 & ~n55216;
  assign n55218 = ~n19213 & ~n55217;
  assign n55219 = ~n3281 & ~n55218;
  assign n55220 = ~n3281 & ~n55219;
  assign n55221 = n3378 & ~n55220;
  assign n55222 = ~n30844 & ~n45971;
  assign n55223 = controllable_nhgrant0 & ~n55222;
  assign n55224 = ~n19255 & ~n55223;
  assign n55225 = ~n3281 & ~n55224;
  assign n55226 = ~n3281 & ~n55225;
  assign n55227 = ~n3378 & ~n55226;
  assign n55228 = ~n55221 & ~n55227;
  assign n55229 = n3492 & ~n55228;
  assign n55230 = n3492 & ~n55229;
  assign n55231 = n3485 & ~n55230;
  assign n55232 = n3485 & ~n55231;
  assign n55233 = ~n3476 & ~n55232;
  assign n55234 = ~n30866 & ~n45999;
  assign n55235 = controllable_nhgrant0 & ~n55234;
  assign n55236 = ~n19385 & ~n55235;
  assign n55237 = ~n3281 & ~n55236;
  assign n55238 = ~n3281 & ~n55237;
  assign n55239 = n3378 & ~n55238;
  assign n55240 = ~n30883 & ~n46043;
  assign n55241 = controllable_nhgrant0 & ~n55240;
  assign n55242 = ~n19515 & ~n55241;
  assign n55243 = ~n3281 & ~n55242;
  assign n55244 = ~n3281 & ~n55243;
  assign n55245 = ~n3378 & ~n55244;
  assign n55246 = ~n55239 & ~n55245;
  assign n55247 = n3492 & ~n55246;
  assign n55248 = n3492 & ~n55247;
  assign n55249 = n3485 & ~n55248;
  assign n55250 = n3485 & ~n55249;
  assign n55251 = n3476 & ~n55250;
  assign n55252 = ~n55233 & ~n55251;
  assign n55253 = n3374 & ~n55252;
  assign n55254 = ~n55215 & ~n55253;
  assign n55255 = n3655 & ~n55254;
  assign n55256 = ~n25905 & ~n46077;
  assign n55257 = controllable_nhgrant0 & ~n55256;
  assign n55258 = ~n7118 & ~n55257;
  assign n55259 = ~n3281 & ~n55258;
  assign n55260 = ~n3281 & ~n55259;
  assign n55261 = ~n3378 & ~n55260;
  assign n55262 = ~n19575 & ~n55261;
  assign n55263 = n3492 & ~n55262;
  assign n55264 = n3492 & ~n55263;
  assign n55265 = n3485 & ~n55264;
  assign n55266 = n3485 & ~n55265;
  assign n55267 = ~n3374 & ~n55266;
  assign n55268 = ~n30827 & ~n46101;
  assign n55269 = controllable_nhgrant0 & ~n55268;
  assign n55270 = ~n19213 & ~n55269;
  assign n55271 = ~n3281 & ~n55270;
  assign n55272 = ~n3281 & ~n55271;
  assign n55273 = n3378 & ~n55272;
  assign n55274 = ~n30844 & ~n46148;
  assign n55275 = controllable_nhgrant0 & ~n55274;
  assign n55276 = ~n19255 & ~n55275;
  assign n55277 = ~n3281 & ~n55276;
  assign n55278 = ~n3281 & ~n55277;
  assign n55279 = ~n3378 & ~n55278;
  assign n55280 = ~n55273 & ~n55279;
  assign n55281 = n3492 & ~n55280;
  assign n55282 = n3492 & ~n55281;
  assign n55283 = n3485 & ~n55282;
  assign n55284 = n3485 & ~n55283;
  assign n55285 = ~n3476 & ~n55284;
  assign n55286 = ~n30866 & ~n46176;
  assign n55287 = controllable_nhgrant0 & ~n55286;
  assign n55288 = ~n19385 & ~n55287;
  assign n55289 = ~n3281 & ~n55288;
  assign n55290 = ~n3281 & ~n55289;
  assign n55291 = n3378 & ~n55290;
  assign n55292 = ~n30883 & ~n46233;
  assign n55293 = controllable_nhgrant0 & ~n55292;
  assign n55294 = ~n19515 & ~n55293;
  assign n55295 = ~n3281 & ~n55294;
  assign n55296 = ~n3281 & ~n55295;
  assign n55297 = ~n3378 & ~n55296;
  assign n55298 = ~n55291 & ~n55297;
  assign n55299 = n3492 & ~n55298;
  assign n55300 = ~n18151 & ~n55299;
  assign n55301 = n3485 & ~n55300;
  assign n55302 = ~n18150 & ~n55301;
  assign n55303 = n3476 & ~n55302;
  assign n55304 = ~n55285 & ~n55303;
  assign n55305 = n3374 & ~n55304;
  assign n55306 = ~n55267 & ~n55305;
  assign n55307 = ~n3655 & ~n55306;
  assign n55308 = ~n55255 & ~n55307;
  assign n55309 = ~n3652 & ~n55308;
  assign n55310 = ~n55203 & ~n55309;
  assign n55311 = n3368 & ~n55310;
  assign n55312 = ~n55109 & ~n55311;
  assign n55313 = n3362 & ~n55312;
  assign n55314 = n3492 & ~n54906;
  assign n55315 = ~n3631 & ~n55314;
  assign n55316 = n3485 & ~n55315;
  assign n55317 = ~n3630 & ~n55316;
  assign n55318 = ~n3476 & ~n55317;
  assign n55319 = n3492 & ~n54924;
  assign n55320 = ~n3631 & ~n55319;
  assign n55321 = n3485 & ~n55320;
  assign n55322 = ~n54016 & ~n55321;
  assign n55323 = n3476 & ~n55322;
  assign n55324 = ~n55318 & ~n55323;
  assign n55325 = n3374 & ~n55324;
  assign n55326 = ~n54020 & ~n55325;
  assign n55327 = n3655 & ~n55326;
  assign n55328 = n3492 & ~n54940;
  assign n55329 = ~n3631 & ~n55328;
  assign n55330 = n3485 & ~n55329;
  assign n55331 = ~n3630 & ~n55330;
  assign n55332 = ~n3476 & ~n55331;
  assign n55333 = ~n20467 & ~n51191;
  assign n55334 = ~n3485 & ~n55333;
  assign n55335 = ~n18630 & ~n55328;
  assign n55336 = n3485 & ~n55335;
  assign n55337 = ~n55334 & ~n55336;
  assign n55338 = n3476 & ~n55337;
  assign n55339 = ~n55332 & ~n55338;
  assign n55340 = ~n3374 & ~n55339;
  assign n55341 = n3492 & ~n54964;
  assign n55342 = ~n3631 & ~n55341;
  assign n55343 = n3485 & ~n55342;
  assign n55344 = ~n3630 & ~n55343;
  assign n55345 = ~n3476 & ~n55344;
  assign n55346 = n3492 & ~n54982;
  assign n55347 = ~n18630 & ~n55346;
  assign n55348 = n3485 & ~n55347;
  assign n55349 = ~n55334 & ~n55348;
  assign n55350 = n3476 & ~n55349;
  assign n55351 = ~n55345 & ~n55350;
  assign n55352 = n3374 & ~n55351;
  assign n55353 = ~n55340 & ~n55352;
  assign n55354 = ~n3655 & ~n55353;
  assign n55355 = ~n55327 & ~n55354;
  assign n55356 = n3652 & ~n55355;
  assign n55357 = n3492 & ~n55000;
  assign n55358 = ~n3631 & ~n55357;
  assign n55359 = n3485 & ~n55358;
  assign n55360 = ~n3630 & ~n55359;
  assign n55361 = ~n3476 & ~n55360;
  assign n55362 = ~n8310 & ~n51236;
  assign n55363 = ~n3485 & ~n55362;
  assign n55364 = ~n55359 & ~n55363;
  assign n55365 = n3476 & ~n55364;
  assign n55366 = ~n55361 & ~n55365;
  assign n55367 = ~n3374 & ~n55366;
  assign n55368 = n3492 & ~n55018;
  assign n55369 = ~n3631 & ~n55368;
  assign n55370 = n3485 & ~n55369;
  assign n55371 = ~n3630 & ~n55370;
  assign n55372 = ~n3476 & ~n55371;
  assign n55373 = n3492 & ~n55036;
  assign n55374 = ~n3631 & ~n55373;
  assign n55375 = n3485 & ~n55374;
  assign n55376 = ~n55363 & ~n55375;
  assign n55377 = n3476 & ~n55376;
  assign n55378 = ~n55372 & ~n55377;
  assign n55379 = n3374 & ~n55378;
  assign n55380 = ~n55367 & ~n55379;
  assign n55381 = n3655 & ~n55380;
  assign n55382 = n3492 & ~n55052;
  assign n55383 = ~n3631 & ~n55382;
  assign n55384 = n3485 & ~n55383;
  assign n55385 = ~n3630 & ~n55384;
  assign n55386 = ~n3476 & ~n55385;
  assign n55387 = ~n20467 & ~n51279;
  assign n55388 = ~n3485 & ~n55387;
  assign n55389 = ~n18630 & ~n55382;
  assign n55390 = n3485 & ~n55389;
  assign n55391 = ~n55388 & ~n55390;
  assign n55392 = n3476 & ~n55391;
  assign n55393 = ~n55386 & ~n55392;
  assign n55394 = ~n3374 & ~n55393;
  assign n55395 = n3492 & ~n55076;
  assign n55396 = ~n3631 & ~n55395;
  assign n55397 = n3485 & ~n55396;
  assign n55398 = ~n3630 & ~n55397;
  assign n55399 = ~n3476 & ~n55398;
  assign n55400 = n3492 & ~n55094;
  assign n55401 = ~n18630 & ~n55400;
  assign n55402 = n3485 & ~n55401;
  assign n55403 = ~n55388 & ~n55402;
  assign n55404 = n3476 & ~n55403;
  assign n55405 = ~n55399 & ~n55404;
  assign n55406 = n3374 & ~n55405;
  assign n55407 = ~n55394 & ~n55406;
  assign n55408 = ~n3655 & ~n55407;
  assign n55409 = ~n55381 & ~n55408;
  assign n55410 = ~n3652 & ~n55409;
  assign n55411 = ~n55356 & ~n55410;
  assign n55412 = ~n3368 & ~n55411;
  assign n55413 = n3492 & ~n55120;
  assign n55414 = n3492 & ~n55413;
  assign n55415 = n3485 & ~n55414;
  assign n55416 = n3485 & ~n55415;
  assign n55417 = ~n3476 & ~n55416;
  assign n55418 = n3492 & ~n55138;
  assign n55419 = n3492 & ~n55418;
  assign n55420 = n3485 & ~n55419;
  assign n55421 = ~n54135 & ~n55420;
  assign n55422 = n3476 & ~n55421;
  assign n55423 = ~n55417 & ~n55422;
  assign n55424 = n3374 & ~n55423;
  assign n55425 = ~n54128 & ~n55424;
  assign n55426 = n3655 & ~n55425;
  assign n55427 = n3492 & ~n55154;
  assign n55428 = n3492 & ~n55427;
  assign n55429 = n3485 & ~n55428;
  assign n55430 = n3485 & ~n55429;
  assign n55431 = ~n3476 & ~n55430;
  assign n55432 = ~n8525 & ~n55429;
  assign n55433 = n3476 & ~n55432;
  assign n55434 = ~n55431 & ~n55433;
  assign n55435 = ~n3374 & ~n55434;
  assign n55436 = n3492 & ~n55172;
  assign n55437 = n3492 & ~n55436;
  assign n55438 = n3485 & ~n55437;
  assign n55439 = n3485 & ~n55438;
  assign n55440 = ~n3476 & ~n55439;
  assign n55441 = ~n20565 & ~n51348;
  assign n55442 = ~n3485 & ~n55441;
  assign n55443 = n3492 & ~n55190;
  assign n55444 = ~n18151 & ~n55443;
  assign n55445 = n3485 & ~n55444;
  assign n55446 = ~n55442 & ~n55445;
  assign n55447 = n3476 & ~n55446;
  assign n55448 = ~n55440 & ~n55447;
  assign n55449 = n3374 & ~n55448;
  assign n55450 = ~n55435 & ~n55449;
  assign n55451 = ~n3655 & ~n55450;
  assign n55452 = ~n55426 & ~n55451;
  assign n55453 = n3652 & ~n55452;
  assign n55454 = n3492 & ~n55208;
  assign n55455 = n3492 & ~n55454;
  assign n55456 = n3485 & ~n55455;
  assign n55457 = n3485 & ~n55456;
  assign n55458 = ~n3476 & ~n55457;
  assign n55459 = ~n8525 & ~n55456;
  assign n55460 = n3476 & ~n55459;
  assign n55461 = ~n55458 & ~n55460;
  assign n55462 = ~n3374 & ~n55461;
  assign n55463 = n3492 & ~n55226;
  assign n55464 = n3492 & ~n55463;
  assign n55465 = n3485 & ~n55464;
  assign n55466 = n3485 & ~n55465;
  assign n55467 = ~n3476 & ~n55466;
  assign n55468 = ~n3492 & ~n51377;
  assign n55469 = ~n3485 & ~n55468;
  assign n55470 = n3492 & ~n55244;
  assign n55471 = n3492 & ~n55470;
  assign n55472 = n3485 & ~n55471;
  assign n55473 = ~n55469 & ~n55472;
  assign n55474 = n3476 & ~n55473;
  assign n55475 = ~n55467 & ~n55474;
  assign n55476 = n3374 & ~n55475;
  assign n55477 = ~n55462 & ~n55476;
  assign n55478 = n3655 & ~n55477;
  assign n55479 = n3492 & ~n55260;
  assign n55480 = n3492 & ~n55479;
  assign n55481 = n3485 & ~n55480;
  assign n55482 = n3485 & ~n55481;
  assign n55483 = ~n3476 & ~n55482;
  assign n55484 = ~n8525 & ~n55481;
  assign n55485 = n3476 & ~n55484;
  assign n55486 = ~n55483 & ~n55485;
  assign n55487 = ~n3374 & ~n55486;
  assign n55488 = n3492 & ~n55278;
  assign n55489 = n3492 & ~n55488;
  assign n55490 = n3485 & ~n55489;
  assign n55491 = n3485 & ~n55490;
  assign n55492 = ~n3476 & ~n55491;
  assign n55493 = ~n20565 & ~n51404;
  assign n55494 = ~n3485 & ~n55493;
  assign n55495 = n3492 & ~n55296;
  assign n55496 = ~n18151 & ~n55495;
  assign n55497 = n3485 & ~n55496;
  assign n55498 = ~n55494 & ~n55497;
  assign n55499 = n3476 & ~n55498;
  assign n55500 = ~n55492 & ~n55499;
  assign n55501 = n3374 & ~n55500;
  assign n55502 = ~n55487 & ~n55501;
  assign n55503 = ~n3655 & ~n55502;
  assign n55504 = ~n55478 & ~n55503;
  assign n55505 = ~n3652 & ~n55504;
  assign n55506 = ~n55453 & ~n55505;
  assign n55507 = n3368 & ~n55506;
  assign n55508 = ~n55412 & ~n55507;
  assign n55509 = ~n3362 & ~n55508;
  assign n55510 = ~n55313 & ~n55509;
  assign n55511 = n3359 & ~n55510;
  assign n55512 = ~n51424 & ~n55321;
  assign n55513 = n3476 & ~n55512;
  assign n55514 = ~n55318 & ~n55513;
  assign n55515 = n3374 & ~n55514;
  assign n55516 = ~n54233 & ~n55515;
  assign n55517 = n3655 & ~n55516;
  assign n55518 = ~n51435 & ~n55336;
  assign n55519 = n3476 & ~n55518;
  assign n55520 = ~n55332 & ~n55519;
  assign n55521 = ~n3374 & ~n55520;
  assign n55522 = ~n51435 & ~n55348;
  assign n55523 = n3476 & ~n55522;
  assign n55524 = ~n55345 & ~n55523;
  assign n55525 = n3374 & ~n55524;
  assign n55526 = ~n55521 & ~n55525;
  assign n55527 = ~n3655 & ~n55526;
  assign n55528 = ~n55517 & ~n55527;
  assign n55529 = n3652 & ~n55528;
  assign n55530 = ~n51448 & ~n55359;
  assign n55531 = n3476 & ~n55530;
  assign n55532 = ~n55361 & ~n55531;
  assign n55533 = ~n3374 & ~n55532;
  assign n55534 = ~n51448 & ~n55375;
  assign n55535 = n3476 & ~n55534;
  assign n55536 = ~n55372 & ~n55535;
  assign n55537 = n3374 & ~n55536;
  assign n55538 = ~n55533 & ~n55537;
  assign n55539 = n3655 & ~n55538;
  assign n55540 = ~n51459 & ~n55390;
  assign n55541 = n3476 & ~n55540;
  assign n55542 = ~n55386 & ~n55541;
  assign n55543 = ~n3374 & ~n55542;
  assign n55544 = ~n51459 & ~n55402;
  assign n55545 = n3476 & ~n55544;
  assign n55546 = ~n55399 & ~n55545;
  assign n55547 = n3374 & ~n55546;
  assign n55548 = ~n55543 & ~n55547;
  assign n55549 = ~n3655 & ~n55548;
  assign n55550 = ~n55539 & ~n55549;
  assign n55551 = ~n3652 & ~n55550;
  assign n55552 = ~n55529 & ~n55551;
  assign n55553 = ~n3368 & ~n55552;
  assign n55554 = ~n51478 & ~n55420;
  assign n55555 = n3476 & ~n55554;
  assign n55556 = ~n55417 & ~n55555;
  assign n55557 = n3374 & ~n55556;
  assign n55558 = ~n54279 & ~n55557;
  assign n55559 = n3655 & ~n55558;
  assign n55560 = ~n8689 & ~n55429;
  assign n55561 = n3476 & ~n55560;
  assign n55562 = ~n55431 & ~n55561;
  assign n55563 = ~n3374 & ~n55562;
  assign n55564 = ~n51489 & ~n55445;
  assign n55565 = n3476 & ~n55564;
  assign n55566 = ~n55440 & ~n55565;
  assign n55567 = n3374 & ~n55566;
  assign n55568 = ~n55563 & ~n55567;
  assign n55569 = ~n3655 & ~n55568;
  assign n55570 = ~n55559 & ~n55569;
  assign n55571 = n3652 & ~n55570;
  assign n55572 = ~n8689 & ~n55456;
  assign n55573 = n3476 & ~n55572;
  assign n55574 = ~n55458 & ~n55573;
  assign n55575 = ~n3374 & ~n55574;
  assign n55576 = ~n51502 & ~n55472;
  assign n55577 = n3476 & ~n55576;
  assign n55578 = ~n55467 & ~n55577;
  assign n55579 = n3374 & ~n55578;
  assign n55580 = ~n55575 & ~n55579;
  assign n55581 = n3655 & ~n55580;
  assign n55582 = ~n8689 & ~n55481;
  assign n55583 = n3476 & ~n55582;
  assign n55584 = ~n55483 & ~n55583;
  assign n55585 = ~n3374 & ~n55584;
  assign n55586 = ~n51513 & ~n55497;
  assign n55587 = n3476 & ~n55586;
  assign n55588 = ~n55492 & ~n55587;
  assign n55589 = n3374 & ~n55588;
  assign n55590 = ~n55585 & ~n55589;
  assign n55591 = ~n3655 & ~n55590;
  assign n55592 = ~n55581 & ~n55591;
  assign n55593 = ~n3652 & ~n55592;
  assign n55594 = ~n55571 & ~n55593;
  assign n55595 = n3368 & ~n55594;
  assign n55596 = ~n55553 & ~n55595;
  assign n55597 = n3362 & ~n55596;
  assign n55598 = n3378 & ~n54906;
  assign n55599 = ~n51551 & ~n55598;
  assign n55600 = n3492 & ~n55599;
  assign n55601 = ~n3631 & ~n55600;
  assign n55602 = n3485 & ~n55601;
  assign n55603 = ~n3630 & ~n55602;
  assign n55604 = ~n3476 & ~n55603;
  assign n55605 = n3378 & ~n54924;
  assign n55606 = ~n51564 & ~n55605;
  assign n55607 = n3492 & ~n55606;
  assign n55608 = ~n51148 & ~n55607;
  assign n55609 = n3485 & ~n55608;
  assign n55610 = ~n51424 & ~n55609;
  assign n55611 = n3476 & ~n55610;
  assign n55612 = ~n55604 & ~n55611;
  assign n55613 = n3374 & ~n55612;
  assign n55614 = ~n54336 & ~n55613;
  assign n55615 = n3655 & ~n55614;
  assign n55616 = n3378 & ~n54940;
  assign n55617 = ~n51581 & ~n55616;
  assign n55618 = n3492 & ~n55617;
  assign n55619 = ~n3631 & ~n55618;
  assign n55620 = n3485 & ~n55619;
  assign n55621 = ~n3630 & ~n55620;
  assign n55622 = ~n3476 & ~n55621;
  assign n55623 = ~n51191 & ~n55618;
  assign n55624 = n3485 & ~n55623;
  assign n55625 = ~n51435 & ~n55624;
  assign n55626 = n3476 & ~n55625;
  assign n55627 = ~n55622 & ~n55626;
  assign n55628 = ~n3374 & ~n55627;
  assign n55629 = n3378 & ~n54964;
  assign n55630 = ~n51600 & ~n55629;
  assign n55631 = n3492 & ~n55630;
  assign n55632 = ~n3631 & ~n55631;
  assign n55633 = n3485 & ~n55632;
  assign n55634 = ~n3630 & ~n55633;
  assign n55635 = ~n3476 & ~n55634;
  assign n55636 = n3378 & ~n54982;
  assign n55637 = ~n51613 & ~n55636;
  assign n55638 = n3492 & ~n55637;
  assign n55639 = ~n51191 & ~n55638;
  assign n55640 = n3485 & ~n55639;
  assign n55641 = ~n51435 & ~n55640;
  assign n55642 = n3476 & ~n55641;
  assign n55643 = ~n55635 & ~n55642;
  assign n55644 = n3374 & ~n55643;
  assign n55645 = ~n55628 & ~n55644;
  assign n55646 = ~n3655 & ~n55645;
  assign n55647 = ~n55615 & ~n55646;
  assign n55648 = n3652 & ~n55647;
  assign n55649 = n3378 & ~n55000;
  assign n55650 = ~n51632 & ~n55649;
  assign n55651 = n3492 & ~n55650;
  assign n55652 = ~n3631 & ~n55651;
  assign n55653 = n3485 & ~n55652;
  assign n55654 = ~n3630 & ~n55653;
  assign n55655 = ~n3476 & ~n55654;
  assign n55656 = ~n51236 & ~n55651;
  assign n55657 = n3485 & ~n55656;
  assign n55658 = ~n51448 & ~n55657;
  assign n55659 = n3476 & ~n55658;
  assign n55660 = ~n55655 & ~n55659;
  assign n55661 = ~n3374 & ~n55660;
  assign n55662 = n3378 & ~n55018;
  assign n55663 = ~n51651 & ~n55662;
  assign n55664 = n3492 & ~n55663;
  assign n55665 = ~n3631 & ~n55664;
  assign n55666 = n3485 & ~n55665;
  assign n55667 = ~n3630 & ~n55666;
  assign n55668 = ~n3476 & ~n55667;
  assign n55669 = n3378 & ~n55036;
  assign n55670 = ~n51664 & ~n55669;
  assign n55671 = n3492 & ~n55670;
  assign n55672 = ~n51236 & ~n55671;
  assign n55673 = n3485 & ~n55672;
  assign n55674 = ~n51448 & ~n55673;
  assign n55675 = n3476 & ~n55674;
  assign n55676 = ~n55668 & ~n55675;
  assign n55677 = n3374 & ~n55676;
  assign n55678 = ~n55661 & ~n55677;
  assign n55679 = n3655 & ~n55678;
  assign n55680 = n3378 & ~n55052;
  assign n55681 = ~n51681 & ~n55680;
  assign n55682 = n3492 & ~n55681;
  assign n55683 = ~n3631 & ~n55682;
  assign n55684 = n3485 & ~n55683;
  assign n55685 = ~n3630 & ~n55684;
  assign n55686 = ~n3476 & ~n55685;
  assign n55687 = ~n51279 & ~n55682;
  assign n55688 = n3485 & ~n55687;
  assign n55689 = ~n51459 & ~n55688;
  assign n55690 = n3476 & ~n55689;
  assign n55691 = ~n55686 & ~n55690;
  assign n55692 = ~n3374 & ~n55691;
  assign n55693 = n3378 & ~n55076;
  assign n55694 = ~n51700 & ~n55693;
  assign n55695 = n3492 & ~n55694;
  assign n55696 = ~n3631 & ~n55695;
  assign n55697 = n3485 & ~n55696;
  assign n55698 = ~n3630 & ~n55697;
  assign n55699 = ~n3476 & ~n55698;
  assign n55700 = n3378 & ~n55094;
  assign n55701 = ~n51713 & ~n55700;
  assign n55702 = n3492 & ~n55701;
  assign n55703 = ~n51279 & ~n55702;
  assign n55704 = n3485 & ~n55703;
  assign n55705 = ~n51459 & ~n55704;
  assign n55706 = n3476 & ~n55705;
  assign n55707 = ~n55699 & ~n55706;
  assign n55708 = n3374 & ~n55707;
  assign n55709 = ~n55692 & ~n55708;
  assign n55710 = ~n3655 & ~n55709;
  assign n55711 = ~n55679 & ~n55710;
  assign n55712 = ~n3652 & ~n55711;
  assign n55713 = ~n55648 & ~n55712;
  assign n55714 = ~n3368 & ~n55713;
  assign n55715 = n3378 & ~n55120;
  assign n55716 = ~n51753 & ~n55715;
  assign n55717 = n3492 & ~n55716;
  assign n55718 = n3492 & ~n55717;
  assign n55719 = n3485 & ~n55718;
  assign n55720 = n3485 & ~n55719;
  assign n55721 = ~n3476 & ~n55720;
  assign n55722 = ~n31444 & ~n46675;
  assign n55723 = controllable_nhgrant0 & ~n55722;
  assign n55724 = ~n20915 & ~n55723;
  assign n55725 = ~n3281 & ~n55724;
  assign n55726 = ~n3281 & ~n55725;
  assign n55727 = n3378 & ~n55726;
  assign n55728 = ~n51771 & ~n55727;
  assign n55729 = n3492 & ~n55728;
  assign n55730 = ~n51321 & ~n55729;
  assign n55731 = n3485 & ~n55730;
  assign n55732 = ~n51478 & ~n55731;
  assign n55733 = n3476 & ~n55732;
  assign n55734 = ~n55721 & ~n55733;
  assign n55735 = n3374 & ~n55734;
  assign n55736 = ~n54466 & ~n55735;
  assign n55737 = n3655 & ~n55736;
  assign n55738 = n3378 & ~n55154;
  assign n55739 = ~n51788 & ~n55738;
  assign n55740 = n3492 & ~n55739;
  assign n55741 = n3492 & ~n55740;
  assign n55742 = n3485 & ~n55741;
  assign n55743 = n3485 & ~n55742;
  assign n55744 = ~n3476 & ~n55743;
  assign n55745 = ~n8523 & ~n55740;
  assign n55746 = n3485 & ~n55745;
  assign n55747 = ~n8689 & ~n55746;
  assign n55748 = n3476 & ~n55747;
  assign n55749 = ~n55744 & ~n55748;
  assign n55750 = ~n3374 & ~n55749;
  assign n55751 = n3378 & ~n55172;
  assign n55752 = ~n51807 & ~n55751;
  assign n55753 = n3492 & ~n55752;
  assign n55754 = n3492 & ~n55753;
  assign n55755 = n3485 & ~n55754;
  assign n55756 = n3485 & ~n55755;
  assign n55757 = ~n3476 & ~n55756;
  assign n55758 = ~n31444 & ~n46789;
  assign n55759 = controllable_nhgrant0 & ~n55758;
  assign n55760 = ~n20915 & ~n55759;
  assign n55761 = ~n3281 & ~n55760;
  assign n55762 = ~n3281 & ~n55761;
  assign n55763 = n3378 & ~n55762;
  assign n55764 = ~n51825 & ~n55763;
  assign n55765 = n3492 & ~n55764;
  assign n55766 = ~n51348 & ~n55765;
  assign n55767 = n3485 & ~n55766;
  assign n55768 = ~n51489 & ~n55767;
  assign n55769 = n3476 & ~n55768;
  assign n55770 = ~n55757 & ~n55769;
  assign n55771 = n3374 & ~n55770;
  assign n55772 = ~n55750 & ~n55771;
  assign n55773 = ~n3655 & ~n55772;
  assign n55774 = ~n55737 & ~n55773;
  assign n55775 = n3652 & ~n55774;
  assign n55776 = n3378 & ~n55208;
  assign n55777 = ~n51844 & ~n55776;
  assign n55778 = n3492 & ~n55777;
  assign n55779 = n3492 & ~n55778;
  assign n55780 = n3485 & ~n55779;
  assign n55781 = n3485 & ~n55780;
  assign n55782 = ~n3476 & ~n55781;
  assign n55783 = ~n8523 & ~n55778;
  assign n55784 = n3485 & ~n55783;
  assign n55785 = ~n8689 & ~n55784;
  assign n55786 = n3476 & ~n55785;
  assign n55787 = ~n55782 & ~n55786;
  assign n55788 = ~n3374 & ~n55787;
  assign n55789 = n3378 & ~n55226;
  assign n55790 = ~n51863 & ~n55789;
  assign n55791 = n3492 & ~n55790;
  assign n55792 = n3492 & ~n55791;
  assign n55793 = n3485 & ~n55792;
  assign n55794 = n3485 & ~n55793;
  assign n55795 = ~n3476 & ~n55794;
  assign n55796 = ~n31444 & ~n46850;
  assign n55797 = controllable_nhgrant0 & ~n55796;
  assign n55798 = ~n20915 & ~n55797;
  assign n55799 = ~n3281 & ~n55798;
  assign n55800 = ~n3281 & ~n55799;
  assign n55801 = n3378 & ~n55800;
  assign n55802 = ~n51881 & ~n55801;
  assign n55803 = n3492 & ~n55802;
  assign n55804 = ~n51377 & ~n55803;
  assign n55805 = n3485 & ~n55804;
  assign n55806 = ~n51502 & ~n55805;
  assign n55807 = n3476 & ~n55806;
  assign n55808 = ~n55795 & ~n55807;
  assign n55809 = n3374 & ~n55808;
  assign n55810 = ~n55788 & ~n55809;
  assign n55811 = n3655 & ~n55810;
  assign n55812 = n3378 & ~n55260;
  assign n55813 = ~n51898 & ~n55812;
  assign n55814 = n3492 & ~n55813;
  assign n55815 = n3492 & ~n55814;
  assign n55816 = n3485 & ~n55815;
  assign n55817 = n3485 & ~n55816;
  assign n55818 = ~n3476 & ~n55817;
  assign n55819 = ~n8523 & ~n55814;
  assign n55820 = n3485 & ~n55819;
  assign n55821 = ~n8689 & ~n55820;
  assign n55822 = n3476 & ~n55821;
  assign n55823 = ~n55818 & ~n55822;
  assign n55824 = ~n3374 & ~n55823;
  assign n55825 = n3378 & ~n55278;
  assign n55826 = ~n51917 & ~n55825;
  assign n55827 = n3492 & ~n55826;
  assign n55828 = n3492 & ~n55827;
  assign n55829 = n3485 & ~n55828;
  assign n55830 = n3485 & ~n55829;
  assign n55831 = ~n3476 & ~n55830;
  assign n55832 = ~n31444 & ~n46935;
  assign n55833 = controllable_nhgrant0 & ~n55832;
  assign n55834 = ~n20915 & ~n55833;
  assign n55835 = ~n3281 & ~n55834;
  assign n55836 = ~n3281 & ~n55835;
  assign n55837 = n3378 & ~n55836;
  assign n55838 = ~n51935 & ~n55837;
  assign n55839 = n3492 & ~n55838;
  assign n55840 = ~n51404 & ~n55839;
  assign n55841 = n3485 & ~n55840;
  assign n55842 = ~n51513 & ~n55841;
  assign n55843 = n3476 & ~n55842;
  assign n55844 = ~n55831 & ~n55843;
  assign n55845 = n3374 & ~n55844;
  assign n55846 = ~n55824 & ~n55845;
  assign n55847 = ~n3655 & ~n55846;
  assign n55848 = ~n55811 & ~n55847;
  assign n55849 = ~n3652 & ~n55848;
  assign n55850 = ~n55775 & ~n55849;
  assign n55851 = n3368 & ~n55850;
  assign n55852 = ~n55714 & ~n55851;
  assign n55853 = ~n3362 & ~n55852;
  assign n55854 = ~n55597 & ~n55853;
  assign n55855 = ~n3359 & ~n55854;
  assign n55856 = ~n55511 & ~n55855;
  assign n55857 = ~n3356 & ~n55856;
  assign n55858 = ~n54889 & ~n55857;
  assign n55859 = ~n3345 & ~n55858;
  assign n55860 = ~n31577 & ~n46975;
  assign n55861 = controllable_nhgrant0 & ~n55860;
  assign n55862 = ~n21332 & ~n55861;
  assign n55863 = ~n3281 & ~n55862;
  assign n55864 = ~n3281 & ~n55863;
  assign n55865 = n3378 & ~n55864;
  assign n55866 = ~n31585 & ~n46983;
  assign n55867 = controllable_nhgrant0 & ~n55866;
  assign n55868 = ~n21347 & ~n55867;
  assign n55869 = ~n3281 & ~n55868;
  assign n55870 = ~n3950 & ~n55869;
  assign n55871 = ~n3378 & ~n55870;
  assign n55872 = ~n55865 & ~n55871;
  assign n55873 = n3492 & ~n55872;
  assign n55874 = ~n3493 & ~n55873;
  assign n55875 = n3485 & ~n55874;
  assign n55876 = ~n3486 & ~n55875;
  assign n55877 = ~n3476 & ~n55876;
  assign n55878 = ~n21383 & ~n55861;
  assign n55879 = ~n3281 & ~n55878;
  assign n55880 = ~n3281 & ~n55879;
  assign n55881 = n3378 & ~n55880;
  assign n55882 = ~n31585 & ~n47018;
  assign n55883 = controllable_nhgrant0 & ~n55882;
  assign n55884 = ~n21461 & ~n55883;
  assign n55885 = ~n3281 & ~n55884;
  assign n55886 = ~n4089 & ~n55885;
  assign n55887 = ~n3378 & ~n55886;
  assign n55888 = ~n55881 & ~n55887;
  assign n55889 = n3492 & ~n55888;
  assign n55890 = ~n21290 & ~n55889;
  assign n55891 = n3485 & ~n55890;
  assign n55892 = ~n21289 & ~n55891;
  assign n55893 = n3476 & ~n55892;
  assign n55894 = ~n55877 & ~n55893;
  assign n55895 = n3374 & ~n55894;
  assign n55896 = ~n21296 & ~n55895;
  assign n55897 = n3655 & ~n55896;
  assign n55898 = ~n31577 & ~n47046;
  assign n55899 = controllable_nhgrant0 & ~n55898;
  assign n55900 = ~n21332 & ~n55899;
  assign n55901 = ~n3281 & ~n55900;
  assign n55902 = ~n3281 & ~n55901;
  assign n55903 = n3378 & ~n55902;
  assign n55904 = ~n31585 & ~n47054;
  assign n55905 = controllable_nhgrant0 & ~n55904;
  assign n55906 = ~n21347 & ~n55905;
  assign n55907 = ~n3281 & ~n55906;
  assign n55908 = ~n3950 & ~n55907;
  assign n55909 = ~n3378 & ~n55908;
  assign n55910 = ~n55903 & ~n55909;
  assign n55911 = n3492 & ~n55910;
  assign n55912 = ~n3493 & ~n55911;
  assign n55913 = n3485 & ~n55912;
  assign n55914 = ~n3486 & ~n55913;
  assign n55915 = ~n3476 & ~n55914;
  assign n55916 = ~n21383 & ~n55899;
  assign n55917 = ~n3281 & ~n55916;
  assign n55918 = ~n3281 & ~n55917;
  assign n55919 = n3378 & ~n55918;
  assign n55920 = ~n31585 & ~n47089;
  assign n55921 = controllable_nhgrant0 & ~n55920;
  assign n55922 = ~n21461 & ~n55921;
  assign n55923 = ~n3281 & ~n55922;
  assign n55924 = ~n4089 & ~n55923;
  assign n55925 = ~n3378 & ~n55924;
  assign n55926 = ~n55919 & ~n55925;
  assign n55927 = n3492 & ~n55926;
  assign n55928 = ~n21290 & ~n55927;
  assign n55929 = n3485 & ~n55928;
  assign n55930 = ~n21289 & ~n55929;
  assign n55931 = n3476 & ~n55930;
  assign n55932 = ~n55915 & ~n55931;
  assign n55933 = n3374 & ~n55932;
  assign n55934 = ~n21296 & ~n55933;
  assign n55935 = ~n3655 & ~n55934;
  assign n55936 = ~n55897 & ~n55935;
  assign n55937 = n3652 & ~n55936;
  assign n55938 = ~n31577 & ~n47119;
  assign n55939 = controllable_nhgrant0 & ~n55938;
  assign n55940 = ~n21332 & ~n55939;
  assign n55941 = ~n3281 & ~n55940;
  assign n55942 = ~n3281 & ~n55941;
  assign n55943 = n3378 & ~n55942;
  assign n55944 = ~n31585 & ~n47127;
  assign n55945 = controllable_nhgrant0 & ~n55944;
  assign n55946 = ~n21347 & ~n55945;
  assign n55947 = ~n3281 & ~n55946;
  assign n55948 = ~n3950 & ~n55947;
  assign n55949 = ~n3378 & ~n55948;
  assign n55950 = ~n55943 & ~n55949;
  assign n55951 = n3492 & ~n55950;
  assign n55952 = ~n3493 & ~n55951;
  assign n55953 = n3485 & ~n55952;
  assign n55954 = ~n3486 & ~n55953;
  assign n55955 = ~n3476 & ~n55954;
  assign n55956 = ~n21383 & ~n55939;
  assign n55957 = ~n3281 & ~n55956;
  assign n55958 = ~n3281 & ~n55957;
  assign n55959 = n3378 & ~n55958;
  assign n55960 = ~n31585 & ~n47158;
  assign n55961 = controllable_nhgrant0 & ~n55960;
  assign n55962 = ~n21461 & ~n55961;
  assign n55963 = ~n3281 & ~n55962;
  assign n55964 = ~n4089 & ~n55963;
  assign n55965 = ~n3378 & ~n55964;
  assign n55966 = ~n55959 & ~n55965;
  assign n55967 = n3492 & ~n55966;
  assign n55968 = ~n21290 & ~n55967;
  assign n55969 = n3485 & ~n55968;
  assign n55970 = ~n21289 & ~n55969;
  assign n55971 = n3476 & ~n55970;
  assign n55972 = ~n55955 & ~n55971;
  assign n55973 = n3374 & ~n55972;
  assign n55974 = ~n21296 & ~n55973;
  assign n55975 = n3655 & ~n55974;
  assign n55976 = ~n31577 & ~n47186;
  assign n55977 = controllable_nhgrant0 & ~n55976;
  assign n55978 = ~n21332 & ~n55977;
  assign n55979 = ~n3281 & ~n55978;
  assign n55980 = ~n3281 & ~n55979;
  assign n55981 = n3378 & ~n55980;
  assign n55982 = ~n31585 & ~n47194;
  assign n55983 = controllable_nhgrant0 & ~n55982;
  assign n55984 = ~n21347 & ~n55983;
  assign n55985 = ~n3281 & ~n55984;
  assign n55986 = ~n3950 & ~n55985;
  assign n55987 = ~n3378 & ~n55986;
  assign n55988 = ~n55981 & ~n55987;
  assign n55989 = n3492 & ~n55988;
  assign n55990 = ~n3493 & ~n55989;
  assign n55991 = n3485 & ~n55990;
  assign n55992 = ~n3486 & ~n55991;
  assign n55993 = ~n3476 & ~n55992;
  assign n55994 = ~n21383 & ~n55977;
  assign n55995 = ~n3281 & ~n55994;
  assign n55996 = ~n3281 & ~n55995;
  assign n55997 = n3378 & ~n55996;
  assign n55998 = ~n31585 & ~n47225;
  assign n55999 = controllable_nhgrant0 & ~n55998;
  assign n56000 = ~n21461 & ~n55999;
  assign n56001 = ~n3281 & ~n56000;
  assign n56002 = ~n4089 & ~n56001;
  assign n56003 = ~n3378 & ~n56002;
  assign n56004 = ~n55997 & ~n56003;
  assign n56005 = n3492 & ~n56004;
  assign n56006 = ~n21290 & ~n56005;
  assign n56007 = n3485 & ~n56006;
  assign n56008 = ~n21289 & ~n56007;
  assign n56009 = n3476 & ~n56008;
  assign n56010 = ~n55993 & ~n56009;
  assign n56011 = n3374 & ~n56010;
  assign n56012 = ~n21296 & ~n56011;
  assign n56013 = ~n3655 & ~n56012;
  assign n56014 = ~n55975 & ~n56013;
  assign n56015 = ~n3652 & ~n56014;
  assign n56016 = ~n55937 & ~n56015;
  assign n56017 = ~n3368 & ~n56016;
  assign n56018 = ~n31740 & ~n47251;
  assign n56019 = controllable_nhgrant0 & ~n56018;
  assign n56020 = ~n21712 & ~n56019;
  assign n56021 = ~n3281 & ~n56020;
  assign n56022 = ~n3281 & ~n56021;
  assign n56023 = n3492 & ~n56022;
  assign n56024 = n3492 & ~n56023;
  assign n56025 = n3485 & ~n56024;
  assign n56026 = n3485 & ~n56025;
  assign n56027 = ~n3476 & ~n56026;
  assign n56028 = ~n21740 & ~n56019;
  assign n56029 = ~n3281 & ~n56028;
  assign n56030 = ~n3281 & ~n56029;
  assign n56031 = n3492 & ~n56030;
  assign n56032 = ~n21722 & ~n56031;
  assign n56033 = n3485 & ~n56032;
  assign n56034 = ~n21721 & ~n56033;
  assign n56035 = n3476 & ~n56034;
  assign n56036 = ~n56027 & ~n56035;
  assign n56037 = n3374 & ~n56036;
  assign n56038 = n3374 & ~n56037;
  assign n56039 = n3655 & ~n56038;
  assign n56040 = ~n31740 & ~n47279;
  assign n56041 = controllable_nhgrant0 & ~n56040;
  assign n56042 = ~n21712 & ~n56041;
  assign n56043 = ~n3281 & ~n56042;
  assign n56044 = ~n3281 & ~n56043;
  assign n56045 = n3492 & ~n56044;
  assign n56046 = n3492 & ~n56045;
  assign n56047 = n3485 & ~n56046;
  assign n56048 = n3485 & ~n56047;
  assign n56049 = ~n3476 & ~n56048;
  assign n56050 = ~n21740 & ~n56041;
  assign n56051 = ~n3281 & ~n56050;
  assign n56052 = ~n3281 & ~n56051;
  assign n56053 = n3492 & ~n56052;
  assign n56054 = ~n21722 & ~n56053;
  assign n56055 = n3485 & ~n56054;
  assign n56056 = ~n21721 & ~n56055;
  assign n56057 = n3476 & ~n56056;
  assign n56058 = ~n56049 & ~n56057;
  assign n56059 = n3374 & ~n56058;
  assign n56060 = n3374 & ~n56059;
  assign n56061 = ~n3655 & ~n56060;
  assign n56062 = ~n56039 & ~n56061;
  assign n56063 = n3652 & ~n56062;
  assign n56064 = ~n31740 & ~n47309;
  assign n56065 = controllable_nhgrant0 & ~n56064;
  assign n56066 = ~n21712 & ~n56065;
  assign n56067 = ~n3281 & ~n56066;
  assign n56068 = ~n3281 & ~n56067;
  assign n56069 = n3492 & ~n56068;
  assign n56070 = n3492 & ~n56069;
  assign n56071 = n3485 & ~n56070;
  assign n56072 = n3485 & ~n56071;
  assign n56073 = ~n3476 & ~n56072;
  assign n56074 = ~n21740 & ~n56065;
  assign n56075 = ~n3281 & ~n56074;
  assign n56076 = ~n3281 & ~n56075;
  assign n56077 = n3492 & ~n56076;
  assign n56078 = ~n21722 & ~n56077;
  assign n56079 = n3485 & ~n56078;
  assign n56080 = ~n21721 & ~n56079;
  assign n56081 = n3476 & ~n56080;
  assign n56082 = ~n56073 & ~n56081;
  assign n56083 = n3374 & ~n56082;
  assign n56084 = n3374 & ~n56083;
  assign n56085 = n3655 & ~n56084;
  assign n56086 = ~n31740 & ~n47337;
  assign n56087 = controllable_nhgrant0 & ~n56086;
  assign n56088 = ~n21712 & ~n56087;
  assign n56089 = ~n3281 & ~n56088;
  assign n56090 = ~n3281 & ~n56089;
  assign n56091 = n3492 & ~n56090;
  assign n56092 = n3492 & ~n56091;
  assign n56093 = n3485 & ~n56092;
  assign n56094 = n3485 & ~n56093;
  assign n56095 = ~n3476 & ~n56094;
  assign n56096 = ~n21740 & ~n56087;
  assign n56097 = ~n3281 & ~n56096;
  assign n56098 = ~n3281 & ~n56097;
  assign n56099 = n3492 & ~n56098;
  assign n56100 = ~n21722 & ~n56099;
  assign n56101 = n3485 & ~n56100;
  assign n56102 = ~n21721 & ~n56101;
  assign n56103 = n3476 & ~n56102;
  assign n56104 = ~n56095 & ~n56103;
  assign n56105 = n3374 & ~n56104;
  assign n56106 = n3374 & ~n56105;
  assign n56107 = ~n3655 & ~n56106;
  assign n56108 = ~n56085 & ~n56107;
  assign n56109 = ~n3652 & ~n56108;
  assign n56110 = ~n56063 & ~n56109;
  assign n56111 = n3368 & ~n56110;
  assign n56112 = ~n56017 & ~n56111;
  assign n56113 = ~n3362 & ~n56112;
  assign n56114 = ~n3362 & ~n56113;
  assign n56115 = ~n3359 & ~n56114;
  assign n56116 = ~n3359 & ~n56115;
  assign n56117 = n3356 & ~n56116;
  assign n56118 = ~n31848 & ~n47377;
  assign n56119 = controllable_nhgrant0 & ~n56118;
  assign n56120 = ~n8785 & ~n56119;
  assign n56121 = ~n3281 & ~n56120;
  assign n56122 = ~n3783 & ~n56121;
  assign n56123 = ~n3378 & ~n56122;
  assign n56124 = ~n21849 & ~n56123;
  assign n56125 = n3492 & ~n56124;
  assign n56126 = ~n3631 & ~n56125;
  assign n56127 = n3485 & ~n56126;
  assign n56128 = ~n3630 & ~n56127;
  assign n56129 = ~n3476 & ~n56128;
  assign n56130 = ~n8309 & ~n56125;
  assign n56131 = n3485 & ~n56130;
  assign n56132 = ~n8639 & ~n56131;
  assign n56133 = n3476 & ~n56132;
  assign n56134 = ~n56129 & ~n56133;
  assign n56135 = ~n3374 & ~n56134;
  assign n56136 = ~n31876 & ~n47407;
  assign n56137 = controllable_nhgrant0 & ~n56136;
  assign n56138 = ~n8902 & ~n56137;
  assign n56139 = ~n3281 & ~n56138;
  assign n56140 = ~n3950 & ~n56139;
  assign n56141 = n3378 & ~n56140;
  assign n56142 = ~n31890 & ~n47431;
  assign n56143 = controllable_nhgrant0 & ~n56142;
  assign n56144 = ~n8902 & ~n56143;
  assign n56145 = ~n3281 & ~n56144;
  assign n56146 = ~n3950 & ~n56145;
  assign n56147 = ~n3378 & ~n56146;
  assign n56148 = ~n56141 & ~n56147;
  assign n56149 = n3492 & ~n56148;
  assign n56150 = ~n3631 & ~n56149;
  assign n56151 = n3485 & ~n56150;
  assign n56152 = ~n3630 & ~n56151;
  assign n56153 = ~n3476 & ~n56152;
  assign n56154 = ~n31915 & ~n47463;
  assign n56155 = controllable_nhgrant0 & ~n56154;
  assign n56156 = ~n9096 & ~n56155;
  assign n56157 = ~n3281 & ~n56156;
  assign n56158 = ~n4089 & ~n56157;
  assign n56159 = n3378 & ~n56158;
  assign n56160 = ~n31933 & ~n47517;
  assign n56161 = controllable_nhgrant0 & ~n56160;
  assign n56162 = ~n9096 & ~n56161;
  assign n56163 = ~n3281 & ~n56162;
  assign n56164 = ~n4089 & ~n56163;
  assign n56165 = ~n3378 & ~n56164;
  assign n56166 = ~n56159 & ~n56165;
  assign n56167 = n3492 & ~n56166;
  assign n56168 = ~n8309 & ~n56167;
  assign n56169 = n3485 & ~n56168;
  assign n56170 = ~n8639 & ~n56169;
  assign n56171 = n3476 & ~n56170;
  assign n56172 = ~n56153 & ~n56171;
  assign n56173 = n3374 & ~n56172;
  assign n56174 = ~n56135 & ~n56173;
  assign n56175 = n3655 & ~n56174;
  assign n56176 = ~n31848 & ~n47541;
  assign n56177 = controllable_nhgrant0 & ~n56176;
  assign n56178 = ~n8785 & ~n56177;
  assign n56179 = ~n3281 & ~n56178;
  assign n56180 = ~n3783 & ~n56179;
  assign n56181 = ~n3378 & ~n56180;
  assign n56182 = ~n21849 & ~n56181;
  assign n56183 = n3492 & ~n56182;
  assign n56184 = ~n3631 & ~n56183;
  assign n56185 = n3485 & ~n56184;
  assign n56186 = ~n3630 & ~n56185;
  assign n56187 = ~n3476 & ~n56186;
  assign n56188 = ~n8309 & ~n56183;
  assign n56189 = n3485 & ~n56188;
  assign n56190 = ~n8639 & ~n56189;
  assign n56191 = n3476 & ~n56190;
  assign n56192 = ~n56187 & ~n56191;
  assign n56193 = ~n3374 & ~n56192;
  assign n56194 = ~n31876 & ~n47571;
  assign n56195 = controllable_nhgrant0 & ~n56194;
  assign n56196 = ~n8902 & ~n56195;
  assign n56197 = ~n3281 & ~n56196;
  assign n56198 = ~n3950 & ~n56197;
  assign n56199 = n3378 & ~n56198;
  assign n56200 = ~n31890 & ~n47595;
  assign n56201 = controllable_nhgrant0 & ~n56200;
  assign n56202 = ~n8902 & ~n56201;
  assign n56203 = ~n3281 & ~n56202;
  assign n56204 = ~n3950 & ~n56203;
  assign n56205 = ~n3378 & ~n56204;
  assign n56206 = ~n56199 & ~n56205;
  assign n56207 = n3492 & ~n56206;
  assign n56208 = ~n3631 & ~n56207;
  assign n56209 = n3485 & ~n56208;
  assign n56210 = ~n3630 & ~n56209;
  assign n56211 = ~n3476 & ~n56210;
  assign n56212 = ~n31915 & ~n47626;
  assign n56213 = controllable_nhgrant0 & ~n56212;
  assign n56214 = ~n9096 & ~n56213;
  assign n56215 = ~n3281 & ~n56214;
  assign n56216 = ~n4089 & ~n56215;
  assign n56217 = n3378 & ~n56216;
  assign n56218 = ~n31933 & ~n47679;
  assign n56219 = controllable_nhgrant0 & ~n56218;
  assign n56220 = ~n9096 & ~n56219;
  assign n56221 = ~n3281 & ~n56220;
  assign n56222 = ~n4089 & ~n56221;
  assign n56223 = ~n3378 & ~n56222;
  assign n56224 = ~n56217 & ~n56223;
  assign n56225 = n3492 & ~n56224;
  assign n56226 = ~n8309 & ~n56225;
  assign n56227 = n3485 & ~n56226;
  assign n56228 = ~n8639 & ~n56227;
  assign n56229 = n3476 & ~n56228;
  assign n56230 = ~n56211 & ~n56229;
  assign n56231 = n3374 & ~n56230;
  assign n56232 = ~n56193 & ~n56231;
  assign n56233 = ~n3655 & ~n56232;
  assign n56234 = ~n56175 & ~n56233;
  assign n56235 = n3652 & ~n56234;
  assign n56236 = ~n31848 & ~n47705;
  assign n56237 = controllable_nhgrant0 & ~n56236;
  assign n56238 = ~n8785 & ~n56237;
  assign n56239 = ~n3281 & ~n56238;
  assign n56240 = ~n3783 & ~n56239;
  assign n56241 = ~n3378 & ~n56240;
  assign n56242 = ~n21849 & ~n56241;
  assign n56243 = n3492 & ~n56242;
  assign n56244 = ~n3631 & ~n56243;
  assign n56245 = n3485 & ~n56244;
  assign n56246 = ~n3630 & ~n56245;
  assign n56247 = ~n3476 & ~n56246;
  assign n56248 = ~n8309 & ~n56243;
  assign n56249 = n3485 & ~n56248;
  assign n56250 = ~n8639 & ~n56249;
  assign n56251 = n3476 & ~n56250;
  assign n56252 = ~n56247 & ~n56251;
  assign n56253 = ~n3374 & ~n56252;
  assign n56254 = ~n31876 & ~n47735;
  assign n56255 = controllable_nhgrant0 & ~n56254;
  assign n56256 = ~n8902 & ~n56255;
  assign n56257 = ~n3281 & ~n56256;
  assign n56258 = ~n3950 & ~n56257;
  assign n56259 = n3378 & ~n56258;
  assign n56260 = ~n31890 & ~n47759;
  assign n56261 = controllable_nhgrant0 & ~n56260;
  assign n56262 = ~n8902 & ~n56261;
  assign n56263 = ~n3281 & ~n56262;
  assign n56264 = ~n3950 & ~n56263;
  assign n56265 = ~n3378 & ~n56264;
  assign n56266 = ~n56259 & ~n56265;
  assign n56267 = n3492 & ~n56266;
  assign n56268 = ~n3631 & ~n56267;
  assign n56269 = n3485 & ~n56268;
  assign n56270 = ~n3630 & ~n56269;
  assign n56271 = ~n3476 & ~n56270;
  assign n56272 = ~n31915 & ~n47786;
  assign n56273 = controllable_nhgrant0 & ~n56272;
  assign n56274 = ~n9096 & ~n56273;
  assign n56275 = ~n3281 & ~n56274;
  assign n56276 = ~n4089 & ~n56275;
  assign n56277 = n3378 & ~n56276;
  assign n56278 = ~n31933 & ~n47823;
  assign n56279 = controllable_nhgrant0 & ~n56278;
  assign n56280 = ~n9096 & ~n56279;
  assign n56281 = ~n3281 & ~n56280;
  assign n56282 = ~n4089 & ~n56281;
  assign n56283 = ~n3378 & ~n56282;
  assign n56284 = ~n56277 & ~n56283;
  assign n56285 = n3492 & ~n56284;
  assign n56286 = ~n8309 & ~n56285;
  assign n56287 = n3485 & ~n56286;
  assign n56288 = ~n8639 & ~n56287;
  assign n56289 = n3476 & ~n56288;
  assign n56290 = ~n56271 & ~n56289;
  assign n56291 = n3374 & ~n56290;
  assign n56292 = ~n56253 & ~n56291;
  assign n56293 = n3655 & ~n56292;
  assign n56294 = ~n31848 & ~n47847;
  assign n56295 = controllable_nhgrant0 & ~n56294;
  assign n56296 = ~n8785 & ~n56295;
  assign n56297 = ~n3281 & ~n56296;
  assign n56298 = ~n3783 & ~n56297;
  assign n56299 = ~n3378 & ~n56298;
  assign n56300 = ~n21849 & ~n56299;
  assign n56301 = n3492 & ~n56300;
  assign n56302 = ~n3631 & ~n56301;
  assign n56303 = n3485 & ~n56302;
  assign n56304 = ~n3630 & ~n56303;
  assign n56305 = ~n3476 & ~n56304;
  assign n56306 = ~n8309 & ~n56301;
  assign n56307 = n3485 & ~n56306;
  assign n56308 = ~n8639 & ~n56307;
  assign n56309 = n3476 & ~n56308;
  assign n56310 = ~n56305 & ~n56309;
  assign n56311 = ~n3374 & ~n56310;
  assign n56312 = ~n31876 & ~n47877;
  assign n56313 = controllable_nhgrant0 & ~n56312;
  assign n56314 = ~n8902 & ~n56313;
  assign n56315 = ~n3281 & ~n56314;
  assign n56316 = ~n3950 & ~n56315;
  assign n56317 = n3378 & ~n56316;
  assign n56318 = ~n31890 & ~n47901;
  assign n56319 = controllable_nhgrant0 & ~n56318;
  assign n56320 = ~n8902 & ~n56319;
  assign n56321 = ~n3281 & ~n56320;
  assign n56322 = ~n3950 & ~n56321;
  assign n56323 = ~n3378 & ~n56322;
  assign n56324 = ~n56317 & ~n56323;
  assign n56325 = n3492 & ~n56324;
  assign n56326 = ~n3631 & ~n56325;
  assign n56327 = n3485 & ~n56326;
  assign n56328 = ~n3630 & ~n56327;
  assign n56329 = ~n3476 & ~n56328;
  assign n56330 = ~n31915 & ~n47928;
  assign n56331 = controllable_nhgrant0 & ~n56330;
  assign n56332 = ~n9096 & ~n56331;
  assign n56333 = ~n3281 & ~n56332;
  assign n56334 = ~n4089 & ~n56333;
  assign n56335 = n3378 & ~n56334;
  assign n56336 = ~n31933 & ~n47965;
  assign n56337 = controllable_nhgrant0 & ~n56336;
  assign n56338 = ~n9096 & ~n56337;
  assign n56339 = ~n3281 & ~n56338;
  assign n56340 = ~n4089 & ~n56339;
  assign n56341 = ~n3378 & ~n56340;
  assign n56342 = ~n56335 & ~n56341;
  assign n56343 = n3492 & ~n56342;
  assign n56344 = ~n8309 & ~n56343;
  assign n56345 = n3485 & ~n56344;
  assign n56346 = ~n8639 & ~n56345;
  assign n56347 = n3476 & ~n56346;
  assign n56348 = ~n56329 & ~n56347;
  assign n56349 = n3374 & ~n56348;
  assign n56350 = ~n56311 & ~n56349;
  assign n56351 = ~n3655 & ~n56350;
  assign n56352 = ~n56293 & ~n56351;
  assign n56353 = ~n3652 & ~n56352;
  assign n56354 = ~n56235 & ~n56353;
  assign n56355 = ~n3368 & ~n56354;
  assign n56356 = ~n32138 & ~n48001;
  assign n56357 = controllable_nhgrant0 & ~n56356;
  assign n56358 = ~n9753 & ~n56357;
  assign n56359 = ~n3281 & ~n56358;
  assign n56360 = ~n3281 & ~n56359;
  assign n56361 = ~n3378 & ~n56360;
  assign n56362 = ~n22618 & ~n56361;
  assign n56363 = n3492 & ~n56362;
  assign n56364 = n3492 & ~n56363;
  assign n56365 = n3485 & ~n56364;
  assign n56366 = n3485 & ~n56365;
  assign n56367 = ~n3374 & ~n56366;
  assign n56368 = ~n32160 & ~n48025;
  assign n56369 = controllable_nhgrant0 & ~n56368;
  assign n56370 = ~n9861 & ~n56369;
  assign n56371 = ~n3281 & ~n56370;
  assign n56372 = ~n3281 & ~n56371;
  assign n56373 = n3378 & ~n56372;
  assign n56374 = ~n32182 & ~n48071;
  assign n56375 = controllable_nhgrant0 & ~n56374;
  assign n56376 = ~n9861 & ~n56375;
  assign n56377 = ~n3281 & ~n56376;
  assign n56378 = ~n3281 & ~n56377;
  assign n56379 = ~n3378 & ~n56378;
  assign n56380 = ~n56373 & ~n56379;
  assign n56381 = n3492 & ~n56380;
  assign n56382 = n3492 & ~n56381;
  assign n56383 = n3485 & ~n56382;
  assign n56384 = n3485 & ~n56383;
  assign n56385 = ~n3476 & ~n56384;
  assign n56386 = ~n32204 & ~n48096;
  assign n56387 = controllable_nhgrant0 & ~n56386;
  assign n56388 = ~n10240 & ~n56387;
  assign n56389 = ~n3281 & ~n56388;
  assign n56390 = ~n3281 & ~n56389;
  assign n56391 = n3378 & ~n56390;
  assign n56392 = ~n32232 & ~n48152;
  assign n56393 = controllable_nhgrant0 & ~n56392;
  assign n56394 = ~n10240 & ~n56393;
  assign n56395 = ~n3281 & ~n56394;
  assign n56396 = ~n3281 & ~n56395;
  assign n56397 = ~n3378 & ~n56396;
  assign n56398 = ~n56391 & ~n56397;
  assign n56399 = n3492 & ~n56398;
  assign n56400 = ~n21722 & ~n56399;
  assign n56401 = n3485 & ~n56400;
  assign n56402 = ~n21721 & ~n56401;
  assign n56403 = n3476 & ~n56402;
  assign n56404 = ~n56385 & ~n56403;
  assign n56405 = n3374 & ~n56404;
  assign n56406 = ~n56367 & ~n56405;
  assign n56407 = n3655 & ~n56406;
  assign n56408 = ~n32138 & ~n48183;
  assign n56409 = controllable_nhgrant0 & ~n56408;
  assign n56410 = ~n9753 & ~n56409;
  assign n56411 = ~n3281 & ~n56410;
  assign n56412 = ~n3281 & ~n56411;
  assign n56413 = ~n3378 & ~n56412;
  assign n56414 = ~n22618 & ~n56413;
  assign n56415 = n3492 & ~n56414;
  assign n56416 = n3492 & ~n56415;
  assign n56417 = n3485 & ~n56416;
  assign n56418 = n3485 & ~n56417;
  assign n56419 = ~n3374 & ~n56418;
  assign n56420 = ~n32160 & ~n48207;
  assign n56421 = controllable_nhgrant0 & ~n56420;
  assign n56422 = ~n9861 & ~n56421;
  assign n56423 = ~n3281 & ~n56422;
  assign n56424 = ~n3281 & ~n56423;
  assign n56425 = n3378 & ~n56424;
  assign n56426 = ~n32182 & ~n48253;
  assign n56427 = controllable_nhgrant0 & ~n56426;
  assign n56428 = ~n9861 & ~n56427;
  assign n56429 = ~n3281 & ~n56428;
  assign n56430 = ~n3281 & ~n56429;
  assign n56431 = ~n3378 & ~n56430;
  assign n56432 = ~n56425 & ~n56431;
  assign n56433 = n3492 & ~n56432;
  assign n56434 = n3492 & ~n56433;
  assign n56435 = n3485 & ~n56434;
  assign n56436 = n3485 & ~n56435;
  assign n56437 = ~n3476 & ~n56436;
  assign n56438 = ~n32204 & ~n48278;
  assign n56439 = controllable_nhgrant0 & ~n56438;
  assign n56440 = ~n10240 & ~n56439;
  assign n56441 = ~n3281 & ~n56440;
  assign n56442 = ~n3281 & ~n56441;
  assign n56443 = n3378 & ~n56442;
  assign n56444 = ~n32232 & ~n48334;
  assign n56445 = controllable_nhgrant0 & ~n56444;
  assign n56446 = ~n10240 & ~n56445;
  assign n56447 = ~n3281 & ~n56446;
  assign n56448 = ~n3281 & ~n56447;
  assign n56449 = ~n3378 & ~n56448;
  assign n56450 = ~n56443 & ~n56449;
  assign n56451 = n3492 & ~n56450;
  assign n56452 = ~n21722 & ~n56451;
  assign n56453 = n3485 & ~n56452;
  assign n56454 = ~n21721 & ~n56453;
  assign n56455 = n3476 & ~n56454;
  assign n56456 = ~n56437 & ~n56455;
  assign n56457 = n3374 & ~n56456;
  assign n56458 = ~n56419 & ~n56457;
  assign n56459 = ~n3655 & ~n56458;
  assign n56460 = ~n56407 & ~n56459;
  assign n56461 = n3652 & ~n56460;
  assign n56462 = ~n32138 & ~n48363;
  assign n56463 = controllable_nhgrant0 & ~n56462;
  assign n56464 = ~n9753 & ~n56463;
  assign n56465 = ~n3281 & ~n56464;
  assign n56466 = ~n3281 & ~n56465;
  assign n56467 = ~n3378 & ~n56466;
  assign n56468 = ~n22618 & ~n56467;
  assign n56469 = n3492 & ~n56468;
  assign n56470 = n3492 & ~n56469;
  assign n56471 = n3485 & ~n56470;
  assign n56472 = n3485 & ~n56471;
  assign n56473 = ~n3374 & ~n56472;
  assign n56474 = ~n32160 & ~n48387;
  assign n56475 = controllable_nhgrant0 & ~n56474;
  assign n56476 = ~n9861 & ~n56475;
  assign n56477 = ~n3281 & ~n56476;
  assign n56478 = ~n3281 & ~n56477;
  assign n56479 = n3378 & ~n56478;
  assign n56480 = ~n32182 & ~n48421;
  assign n56481 = controllable_nhgrant0 & ~n56480;
  assign n56482 = ~n9861 & ~n56481;
  assign n56483 = ~n3281 & ~n56482;
  assign n56484 = ~n3281 & ~n56483;
  assign n56485 = ~n3378 & ~n56484;
  assign n56486 = ~n56479 & ~n56485;
  assign n56487 = n3492 & ~n56486;
  assign n56488 = n3492 & ~n56487;
  assign n56489 = n3485 & ~n56488;
  assign n56490 = n3485 & ~n56489;
  assign n56491 = ~n3476 & ~n56490;
  assign n56492 = ~n32204 & ~n48446;
  assign n56493 = controllable_nhgrant0 & ~n56492;
  assign n56494 = ~n10240 & ~n56493;
  assign n56495 = ~n3281 & ~n56494;
  assign n56496 = ~n3281 & ~n56495;
  assign n56497 = n3378 & ~n56496;
  assign n56498 = ~n32232 & ~n48484;
  assign n56499 = controllable_nhgrant0 & ~n56498;
  assign n56500 = ~n10240 & ~n56499;
  assign n56501 = ~n3281 & ~n56500;
  assign n56502 = ~n3281 & ~n56501;
  assign n56503 = ~n3378 & ~n56502;
  assign n56504 = ~n56497 & ~n56503;
  assign n56505 = n3492 & ~n56504;
  assign n56506 = ~n21722 & ~n56505;
  assign n56507 = n3485 & ~n56506;
  assign n56508 = ~n21721 & ~n56507;
  assign n56509 = n3476 & ~n56508;
  assign n56510 = ~n56491 & ~n56509;
  assign n56511 = n3374 & ~n56510;
  assign n56512 = ~n56473 & ~n56511;
  assign n56513 = n3655 & ~n56512;
  assign n56514 = ~n32138 & ~n48511;
  assign n56515 = controllable_nhgrant0 & ~n56514;
  assign n56516 = ~n9753 & ~n56515;
  assign n56517 = ~n3281 & ~n56516;
  assign n56518 = ~n3281 & ~n56517;
  assign n56519 = ~n3378 & ~n56518;
  assign n56520 = ~n22618 & ~n56519;
  assign n56521 = n3492 & ~n56520;
  assign n56522 = n3492 & ~n56521;
  assign n56523 = n3485 & ~n56522;
  assign n56524 = n3485 & ~n56523;
  assign n56525 = ~n3374 & ~n56524;
  assign n56526 = ~n32160 & ~n48535;
  assign n56527 = controllable_nhgrant0 & ~n56526;
  assign n56528 = ~n9861 & ~n56527;
  assign n56529 = ~n3281 & ~n56528;
  assign n56530 = ~n3281 & ~n56529;
  assign n56531 = n3378 & ~n56530;
  assign n56532 = ~n32182 & ~n48569;
  assign n56533 = controllable_nhgrant0 & ~n56532;
  assign n56534 = ~n9861 & ~n56533;
  assign n56535 = ~n3281 & ~n56534;
  assign n56536 = ~n3281 & ~n56535;
  assign n56537 = ~n3378 & ~n56536;
  assign n56538 = ~n56531 & ~n56537;
  assign n56539 = n3492 & ~n56538;
  assign n56540 = n3492 & ~n56539;
  assign n56541 = n3485 & ~n56540;
  assign n56542 = n3485 & ~n56541;
  assign n56543 = ~n3476 & ~n56542;
  assign n56544 = ~n32204 & ~n48594;
  assign n56545 = controllable_nhgrant0 & ~n56544;
  assign n56546 = ~n10240 & ~n56545;
  assign n56547 = ~n3281 & ~n56546;
  assign n56548 = ~n3281 & ~n56547;
  assign n56549 = n3378 & ~n56548;
  assign n56550 = ~n32232 & ~n48635;
  assign n56551 = controllable_nhgrant0 & ~n56550;
  assign n56552 = ~n10240 & ~n56551;
  assign n56553 = ~n3281 & ~n56552;
  assign n56554 = ~n3281 & ~n56553;
  assign n56555 = ~n3378 & ~n56554;
  assign n56556 = ~n56549 & ~n56555;
  assign n56557 = n3492 & ~n56556;
  assign n56558 = ~n21722 & ~n56557;
  assign n56559 = n3485 & ~n56558;
  assign n56560 = ~n21721 & ~n56559;
  assign n56561 = n3476 & ~n56560;
  assign n56562 = ~n56543 & ~n56561;
  assign n56563 = n3374 & ~n56562;
  assign n56564 = ~n56525 & ~n56563;
  assign n56565 = ~n3655 & ~n56564;
  assign n56566 = ~n56513 & ~n56565;
  assign n56567 = ~n3652 & ~n56566;
  assign n56568 = ~n56461 & ~n56567;
  assign n56569 = n3368 & ~n56568;
  assign n56570 = ~n56355 & ~n56569;
  assign n56571 = n3362 & ~n56570;
  assign n56572 = n3492 & ~n56122;
  assign n56573 = ~n3631 & ~n56572;
  assign n56574 = n3485 & ~n56573;
  assign n56575 = ~n3630 & ~n56574;
  assign n56576 = ~n3476 & ~n56575;
  assign n56577 = ~n23549 & ~n51148;
  assign n56578 = ~n3485 & ~n56577;
  assign n56579 = ~n8309 & ~n56572;
  assign n56580 = n3485 & ~n56579;
  assign n56581 = ~n56578 & ~n56580;
  assign n56582 = n3476 & ~n56581;
  assign n56583 = ~n56576 & ~n56582;
  assign n56584 = ~n3374 & ~n56583;
  assign n56585 = n3492 & ~n56146;
  assign n56586 = ~n3631 & ~n56585;
  assign n56587 = n3485 & ~n56586;
  assign n56588 = ~n3630 & ~n56587;
  assign n56589 = ~n3476 & ~n56588;
  assign n56590 = n3492 & ~n56164;
  assign n56591 = ~n8309 & ~n56590;
  assign n56592 = n3485 & ~n56591;
  assign n56593 = ~n56578 & ~n56592;
  assign n56594 = n3476 & ~n56593;
  assign n56595 = ~n56589 & ~n56594;
  assign n56596 = n3374 & ~n56595;
  assign n56597 = ~n56584 & ~n56596;
  assign n56598 = n3655 & ~n56597;
  assign n56599 = n3492 & ~n56180;
  assign n56600 = ~n3631 & ~n56599;
  assign n56601 = n3485 & ~n56600;
  assign n56602 = ~n3630 & ~n56601;
  assign n56603 = ~n3476 & ~n56602;
  assign n56604 = ~n23549 & ~n51191;
  assign n56605 = ~n3485 & ~n56604;
  assign n56606 = ~n8309 & ~n56599;
  assign n56607 = n3485 & ~n56606;
  assign n56608 = ~n56605 & ~n56607;
  assign n56609 = n3476 & ~n56608;
  assign n56610 = ~n56603 & ~n56609;
  assign n56611 = ~n3374 & ~n56610;
  assign n56612 = n3492 & ~n56204;
  assign n56613 = ~n3631 & ~n56612;
  assign n56614 = n3485 & ~n56613;
  assign n56615 = ~n3630 & ~n56614;
  assign n56616 = ~n3476 & ~n56615;
  assign n56617 = n3492 & ~n56222;
  assign n56618 = ~n8309 & ~n56617;
  assign n56619 = n3485 & ~n56618;
  assign n56620 = ~n56605 & ~n56619;
  assign n56621 = n3476 & ~n56620;
  assign n56622 = ~n56616 & ~n56621;
  assign n56623 = n3374 & ~n56622;
  assign n56624 = ~n56611 & ~n56623;
  assign n56625 = ~n3655 & ~n56624;
  assign n56626 = ~n56598 & ~n56625;
  assign n56627 = n3652 & ~n56626;
  assign n56628 = n3492 & ~n56240;
  assign n56629 = ~n3631 & ~n56628;
  assign n56630 = n3485 & ~n56629;
  assign n56631 = ~n3630 & ~n56630;
  assign n56632 = ~n3476 & ~n56631;
  assign n56633 = ~n23549 & ~n51236;
  assign n56634 = ~n3485 & ~n56633;
  assign n56635 = ~n8309 & ~n56628;
  assign n56636 = n3485 & ~n56635;
  assign n56637 = ~n56634 & ~n56636;
  assign n56638 = n3476 & ~n56637;
  assign n56639 = ~n56632 & ~n56638;
  assign n56640 = ~n3374 & ~n56639;
  assign n56641 = n3492 & ~n56264;
  assign n56642 = ~n3631 & ~n56641;
  assign n56643 = n3485 & ~n56642;
  assign n56644 = ~n3630 & ~n56643;
  assign n56645 = ~n3476 & ~n56644;
  assign n56646 = n3492 & ~n56282;
  assign n56647 = ~n8309 & ~n56646;
  assign n56648 = n3485 & ~n56647;
  assign n56649 = ~n56634 & ~n56648;
  assign n56650 = n3476 & ~n56649;
  assign n56651 = ~n56645 & ~n56650;
  assign n56652 = n3374 & ~n56651;
  assign n56653 = ~n56640 & ~n56652;
  assign n56654 = n3655 & ~n56653;
  assign n56655 = n3492 & ~n56298;
  assign n56656 = ~n3631 & ~n56655;
  assign n56657 = n3485 & ~n56656;
  assign n56658 = ~n3630 & ~n56657;
  assign n56659 = ~n3476 & ~n56658;
  assign n56660 = ~n23549 & ~n51279;
  assign n56661 = ~n3485 & ~n56660;
  assign n56662 = ~n8309 & ~n56655;
  assign n56663 = n3485 & ~n56662;
  assign n56664 = ~n56661 & ~n56663;
  assign n56665 = n3476 & ~n56664;
  assign n56666 = ~n56659 & ~n56665;
  assign n56667 = ~n3374 & ~n56666;
  assign n56668 = n3492 & ~n56322;
  assign n56669 = ~n3631 & ~n56668;
  assign n56670 = n3485 & ~n56669;
  assign n56671 = ~n3630 & ~n56670;
  assign n56672 = ~n3476 & ~n56671;
  assign n56673 = n3492 & ~n56340;
  assign n56674 = ~n8309 & ~n56673;
  assign n56675 = n3485 & ~n56674;
  assign n56676 = ~n56661 & ~n56675;
  assign n56677 = n3476 & ~n56676;
  assign n56678 = ~n56672 & ~n56677;
  assign n56679 = n3374 & ~n56678;
  assign n56680 = ~n56667 & ~n56679;
  assign n56681 = ~n3655 & ~n56680;
  assign n56682 = ~n56654 & ~n56681;
  assign n56683 = ~n3652 & ~n56682;
  assign n56684 = ~n56627 & ~n56683;
  assign n56685 = ~n3368 & ~n56684;
  assign n56686 = n3492 & ~n56360;
  assign n56687 = n3492 & ~n56686;
  assign n56688 = n3485 & ~n56687;
  assign n56689 = n3485 & ~n56688;
  assign n56690 = ~n3476 & ~n56689;
  assign n56691 = ~n8525 & ~n56688;
  assign n56692 = n3476 & ~n56691;
  assign n56693 = ~n56690 & ~n56692;
  assign n56694 = ~n3374 & ~n56693;
  assign n56695 = n3492 & ~n56378;
  assign n56696 = n3492 & ~n56695;
  assign n56697 = n3485 & ~n56696;
  assign n56698 = n3485 & ~n56697;
  assign n56699 = ~n3476 & ~n56698;
  assign n56700 = ~n23646 & ~n51321;
  assign n56701 = ~n3485 & ~n56700;
  assign n56702 = n3492 & ~n56396;
  assign n56703 = ~n21722 & ~n56702;
  assign n56704 = n3485 & ~n56703;
  assign n56705 = ~n56701 & ~n56704;
  assign n56706 = n3476 & ~n56705;
  assign n56707 = ~n56699 & ~n56706;
  assign n56708 = n3374 & ~n56707;
  assign n56709 = ~n56694 & ~n56708;
  assign n56710 = n3655 & ~n56709;
  assign n56711 = n3492 & ~n56412;
  assign n56712 = n3492 & ~n56711;
  assign n56713 = n3485 & ~n56712;
  assign n56714 = n3485 & ~n56713;
  assign n56715 = ~n3476 & ~n56714;
  assign n56716 = ~n8525 & ~n56713;
  assign n56717 = n3476 & ~n56716;
  assign n56718 = ~n56715 & ~n56717;
  assign n56719 = ~n3374 & ~n56718;
  assign n56720 = n3492 & ~n56430;
  assign n56721 = n3492 & ~n56720;
  assign n56722 = n3485 & ~n56721;
  assign n56723 = n3485 & ~n56722;
  assign n56724 = ~n3476 & ~n56723;
  assign n56725 = ~n23646 & ~n51348;
  assign n56726 = ~n3485 & ~n56725;
  assign n56727 = n3492 & ~n56448;
  assign n56728 = ~n21722 & ~n56727;
  assign n56729 = n3485 & ~n56728;
  assign n56730 = ~n56726 & ~n56729;
  assign n56731 = n3476 & ~n56730;
  assign n56732 = ~n56724 & ~n56731;
  assign n56733 = n3374 & ~n56732;
  assign n56734 = ~n56719 & ~n56733;
  assign n56735 = ~n3655 & ~n56734;
  assign n56736 = ~n56710 & ~n56735;
  assign n56737 = n3652 & ~n56736;
  assign n56738 = n3492 & ~n56466;
  assign n56739 = n3492 & ~n56738;
  assign n56740 = n3485 & ~n56739;
  assign n56741 = n3485 & ~n56740;
  assign n56742 = ~n3476 & ~n56741;
  assign n56743 = ~n8525 & ~n56740;
  assign n56744 = n3476 & ~n56743;
  assign n56745 = ~n56742 & ~n56744;
  assign n56746 = ~n3374 & ~n56745;
  assign n56747 = n3492 & ~n56484;
  assign n56748 = n3492 & ~n56747;
  assign n56749 = n3485 & ~n56748;
  assign n56750 = n3485 & ~n56749;
  assign n56751 = ~n3476 & ~n56750;
  assign n56752 = ~n23646 & ~n51377;
  assign n56753 = ~n3485 & ~n56752;
  assign n56754 = n3492 & ~n56502;
  assign n56755 = ~n21722 & ~n56754;
  assign n56756 = n3485 & ~n56755;
  assign n56757 = ~n56753 & ~n56756;
  assign n56758 = n3476 & ~n56757;
  assign n56759 = ~n56751 & ~n56758;
  assign n56760 = n3374 & ~n56759;
  assign n56761 = ~n56746 & ~n56760;
  assign n56762 = n3655 & ~n56761;
  assign n56763 = n3492 & ~n56518;
  assign n56764 = n3492 & ~n56763;
  assign n56765 = n3485 & ~n56764;
  assign n56766 = n3485 & ~n56765;
  assign n56767 = ~n3476 & ~n56766;
  assign n56768 = ~n8525 & ~n56765;
  assign n56769 = n3476 & ~n56768;
  assign n56770 = ~n56767 & ~n56769;
  assign n56771 = ~n3374 & ~n56770;
  assign n56772 = n3492 & ~n56536;
  assign n56773 = n3492 & ~n56772;
  assign n56774 = n3485 & ~n56773;
  assign n56775 = n3485 & ~n56774;
  assign n56776 = ~n3476 & ~n56775;
  assign n56777 = ~n23646 & ~n51404;
  assign n56778 = ~n3485 & ~n56777;
  assign n56779 = n3492 & ~n56554;
  assign n56780 = ~n21722 & ~n56779;
  assign n56781 = n3485 & ~n56780;
  assign n56782 = ~n56778 & ~n56781;
  assign n56783 = n3476 & ~n56782;
  assign n56784 = ~n56776 & ~n56783;
  assign n56785 = n3374 & ~n56784;
  assign n56786 = ~n56771 & ~n56785;
  assign n56787 = ~n3655 & ~n56786;
  assign n56788 = ~n56762 & ~n56787;
  assign n56789 = ~n3652 & ~n56788;
  assign n56790 = ~n56737 & ~n56789;
  assign n56791 = n3368 & ~n56790;
  assign n56792 = ~n56685 & ~n56791;
  assign n56793 = ~n3362 & ~n56792;
  assign n56794 = ~n56571 & ~n56793;
  assign n56795 = n3359 & ~n56794;
  assign n56796 = ~n51424 & ~n56580;
  assign n56797 = n3476 & ~n56796;
  assign n56798 = ~n56576 & ~n56797;
  assign n56799 = ~n3374 & ~n56798;
  assign n56800 = ~n51424 & ~n56592;
  assign n56801 = n3476 & ~n56800;
  assign n56802 = ~n56589 & ~n56801;
  assign n56803 = n3374 & ~n56802;
  assign n56804 = ~n56799 & ~n56803;
  assign n56805 = n3655 & ~n56804;
  assign n56806 = ~n51435 & ~n56607;
  assign n56807 = n3476 & ~n56806;
  assign n56808 = ~n56603 & ~n56807;
  assign n56809 = ~n3374 & ~n56808;
  assign n56810 = ~n51435 & ~n56619;
  assign n56811 = n3476 & ~n56810;
  assign n56812 = ~n56616 & ~n56811;
  assign n56813 = n3374 & ~n56812;
  assign n56814 = ~n56809 & ~n56813;
  assign n56815 = ~n3655 & ~n56814;
  assign n56816 = ~n56805 & ~n56815;
  assign n56817 = n3652 & ~n56816;
  assign n56818 = ~n51448 & ~n56636;
  assign n56819 = n3476 & ~n56818;
  assign n56820 = ~n56632 & ~n56819;
  assign n56821 = ~n3374 & ~n56820;
  assign n56822 = ~n51448 & ~n56648;
  assign n56823 = n3476 & ~n56822;
  assign n56824 = ~n56645 & ~n56823;
  assign n56825 = n3374 & ~n56824;
  assign n56826 = ~n56821 & ~n56825;
  assign n56827 = n3655 & ~n56826;
  assign n56828 = ~n51459 & ~n56663;
  assign n56829 = n3476 & ~n56828;
  assign n56830 = ~n56659 & ~n56829;
  assign n56831 = ~n3374 & ~n56830;
  assign n56832 = ~n51459 & ~n56675;
  assign n56833 = n3476 & ~n56832;
  assign n56834 = ~n56672 & ~n56833;
  assign n56835 = n3374 & ~n56834;
  assign n56836 = ~n56831 & ~n56835;
  assign n56837 = ~n3655 & ~n56836;
  assign n56838 = ~n56827 & ~n56837;
  assign n56839 = ~n3652 & ~n56838;
  assign n56840 = ~n56817 & ~n56839;
  assign n56841 = ~n3368 & ~n56840;
  assign n56842 = ~n8689 & ~n56688;
  assign n56843 = n3476 & ~n56842;
  assign n56844 = ~n56690 & ~n56843;
  assign n56845 = ~n3374 & ~n56844;
  assign n56846 = ~n51478 & ~n56704;
  assign n56847 = n3476 & ~n56846;
  assign n56848 = ~n56699 & ~n56847;
  assign n56849 = n3374 & ~n56848;
  assign n56850 = ~n56845 & ~n56849;
  assign n56851 = n3655 & ~n56850;
  assign n56852 = ~n8689 & ~n56713;
  assign n56853 = n3476 & ~n56852;
  assign n56854 = ~n56715 & ~n56853;
  assign n56855 = ~n3374 & ~n56854;
  assign n56856 = ~n51489 & ~n56729;
  assign n56857 = n3476 & ~n56856;
  assign n56858 = ~n56724 & ~n56857;
  assign n56859 = n3374 & ~n56858;
  assign n56860 = ~n56855 & ~n56859;
  assign n56861 = ~n3655 & ~n56860;
  assign n56862 = ~n56851 & ~n56861;
  assign n56863 = n3652 & ~n56862;
  assign n56864 = ~n8689 & ~n56740;
  assign n56865 = n3476 & ~n56864;
  assign n56866 = ~n56742 & ~n56865;
  assign n56867 = ~n3374 & ~n56866;
  assign n56868 = ~n51502 & ~n56756;
  assign n56869 = n3476 & ~n56868;
  assign n56870 = ~n56751 & ~n56869;
  assign n56871 = n3374 & ~n56870;
  assign n56872 = ~n56867 & ~n56871;
  assign n56873 = n3655 & ~n56872;
  assign n56874 = ~n8689 & ~n56765;
  assign n56875 = n3476 & ~n56874;
  assign n56876 = ~n56767 & ~n56875;
  assign n56877 = ~n3374 & ~n56876;
  assign n56878 = ~n51513 & ~n56781;
  assign n56879 = n3476 & ~n56878;
  assign n56880 = ~n56776 & ~n56879;
  assign n56881 = n3374 & ~n56880;
  assign n56882 = ~n56877 & ~n56881;
  assign n56883 = ~n3655 & ~n56882;
  assign n56884 = ~n56873 & ~n56883;
  assign n56885 = ~n3652 & ~n56884;
  assign n56886 = ~n56863 & ~n56885;
  assign n56887 = n3368 & ~n56886;
  assign n56888 = ~n56841 & ~n56887;
  assign n56889 = n3362 & ~n56888;
  assign n56890 = n3378 & ~n56122;
  assign n56891 = ~n51532 & ~n56890;
  assign n56892 = n3492 & ~n56891;
  assign n56893 = ~n3631 & ~n56892;
  assign n56894 = n3485 & ~n56893;
  assign n56895 = ~n3630 & ~n56894;
  assign n56896 = ~n3476 & ~n56895;
  assign n56897 = ~n51148 & ~n56892;
  assign n56898 = n3485 & ~n56897;
  assign n56899 = ~n51424 & ~n56898;
  assign n56900 = n3476 & ~n56899;
  assign n56901 = ~n56896 & ~n56900;
  assign n56902 = ~n3374 & ~n56901;
  assign n56903 = n3378 & ~n56146;
  assign n56904 = ~n51551 & ~n56903;
  assign n56905 = n3492 & ~n56904;
  assign n56906 = ~n3631 & ~n56905;
  assign n56907 = n3485 & ~n56906;
  assign n56908 = ~n3630 & ~n56907;
  assign n56909 = ~n3476 & ~n56908;
  assign n56910 = n3378 & ~n56164;
  assign n56911 = ~n51564 & ~n56910;
  assign n56912 = n3492 & ~n56911;
  assign n56913 = ~n51148 & ~n56912;
  assign n56914 = n3485 & ~n56913;
  assign n56915 = ~n51424 & ~n56914;
  assign n56916 = n3476 & ~n56915;
  assign n56917 = ~n56909 & ~n56916;
  assign n56918 = n3374 & ~n56917;
  assign n56919 = ~n56902 & ~n56918;
  assign n56920 = n3655 & ~n56919;
  assign n56921 = n3378 & ~n56180;
  assign n56922 = ~n51581 & ~n56921;
  assign n56923 = n3492 & ~n56922;
  assign n56924 = ~n3631 & ~n56923;
  assign n56925 = n3485 & ~n56924;
  assign n56926 = ~n3630 & ~n56925;
  assign n56927 = ~n3476 & ~n56926;
  assign n56928 = ~n51191 & ~n56923;
  assign n56929 = n3485 & ~n56928;
  assign n56930 = ~n51435 & ~n56929;
  assign n56931 = n3476 & ~n56930;
  assign n56932 = ~n56927 & ~n56931;
  assign n56933 = ~n3374 & ~n56932;
  assign n56934 = n3378 & ~n56204;
  assign n56935 = ~n51600 & ~n56934;
  assign n56936 = n3492 & ~n56935;
  assign n56937 = ~n3631 & ~n56936;
  assign n56938 = n3485 & ~n56937;
  assign n56939 = ~n3630 & ~n56938;
  assign n56940 = ~n3476 & ~n56939;
  assign n56941 = n3378 & ~n56222;
  assign n56942 = ~n51613 & ~n56941;
  assign n56943 = n3492 & ~n56942;
  assign n56944 = ~n51191 & ~n56943;
  assign n56945 = n3485 & ~n56944;
  assign n56946 = ~n51435 & ~n56945;
  assign n56947 = n3476 & ~n56946;
  assign n56948 = ~n56940 & ~n56947;
  assign n56949 = n3374 & ~n56948;
  assign n56950 = ~n56933 & ~n56949;
  assign n56951 = ~n3655 & ~n56950;
  assign n56952 = ~n56920 & ~n56951;
  assign n56953 = n3652 & ~n56952;
  assign n56954 = n3378 & ~n56240;
  assign n56955 = ~n51632 & ~n56954;
  assign n56956 = n3492 & ~n56955;
  assign n56957 = ~n3631 & ~n56956;
  assign n56958 = n3485 & ~n56957;
  assign n56959 = ~n3630 & ~n56958;
  assign n56960 = ~n3476 & ~n56959;
  assign n56961 = ~n51236 & ~n56956;
  assign n56962 = n3485 & ~n56961;
  assign n56963 = ~n51448 & ~n56962;
  assign n56964 = n3476 & ~n56963;
  assign n56965 = ~n56960 & ~n56964;
  assign n56966 = ~n3374 & ~n56965;
  assign n56967 = n3378 & ~n56264;
  assign n56968 = ~n51651 & ~n56967;
  assign n56969 = n3492 & ~n56968;
  assign n56970 = ~n3631 & ~n56969;
  assign n56971 = n3485 & ~n56970;
  assign n56972 = ~n3630 & ~n56971;
  assign n56973 = ~n3476 & ~n56972;
  assign n56974 = n3378 & ~n56282;
  assign n56975 = ~n51664 & ~n56974;
  assign n56976 = n3492 & ~n56975;
  assign n56977 = ~n51236 & ~n56976;
  assign n56978 = n3485 & ~n56977;
  assign n56979 = ~n51448 & ~n56978;
  assign n56980 = n3476 & ~n56979;
  assign n56981 = ~n56973 & ~n56980;
  assign n56982 = n3374 & ~n56981;
  assign n56983 = ~n56966 & ~n56982;
  assign n56984 = n3655 & ~n56983;
  assign n56985 = n3378 & ~n56298;
  assign n56986 = ~n51681 & ~n56985;
  assign n56987 = n3492 & ~n56986;
  assign n56988 = ~n3631 & ~n56987;
  assign n56989 = n3485 & ~n56988;
  assign n56990 = ~n3630 & ~n56989;
  assign n56991 = ~n3476 & ~n56990;
  assign n56992 = ~n51279 & ~n56987;
  assign n56993 = n3485 & ~n56992;
  assign n56994 = ~n51459 & ~n56993;
  assign n56995 = n3476 & ~n56994;
  assign n56996 = ~n56991 & ~n56995;
  assign n56997 = ~n3374 & ~n56996;
  assign n56998 = n3378 & ~n56322;
  assign n56999 = ~n51700 & ~n56998;
  assign n57000 = n3492 & ~n56999;
  assign n57001 = ~n3631 & ~n57000;
  assign n57002 = n3485 & ~n57001;
  assign n57003 = ~n3630 & ~n57002;
  assign n57004 = ~n3476 & ~n57003;
  assign n57005 = n3378 & ~n56340;
  assign n57006 = ~n51713 & ~n57005;
  assign n57007 = n3492 & ~n57006;
  assign n57008 = ~n51279 & ~n57007;
  assign n57009 = n3485 & ~n57008;
  assign n57010 = ~n51459 & ~n57009;
  assign n57011 = n3476 & ~n57010;
  assign n57012 = ~n57004 & ~n57011;
  assign n57013 = n3374 & ~n57012;
  assign n57014 = ~n56997 & ~n57013;
  assign n57015 = ~n3655 & ~n57014;
  assign n57016 = ~n56984 & ~n57015;
  assign n57017 = ~n3652 & ~n57016;
  assign n57018 = ~n56953 & ~n57017;
  assign n57019 = ~n3368 & ~n57018;
  assign n57020 = n3378 & ~n56360;
  assign n57021 = ~n51734 & ~n57020;
  assign n57022 = n3492 & ~n57021;
  assign n57023 = n3492 & ~n57022;
  assign n57024 = n3485 & ~n57023;
  assign n57025 = n3485 & ~n57024;
  assign n57026 = ~n3476 & ~n57025;
  assign n57027 = ~n8523 & ~n57022;
  assign n57028 = n3485 & ~n57027;
  assign n57029 = ~n8689 & ~n57028;
  assign n57030 = n3476 & ~n57029;
  assign n57031 = ~n57026 & ~n57030;
  assign n57032 = ~n3374 & ~n57031;
  assign n57033 = n3378 & ~n56378;
  assign n57034 = ~n51753 & ~n57033;
  assign n57035 = n3492 & ~n57034;
  assign n57036 = n3492 & ~n57035;
  assign n57037 = n3485 & ~n57036;
  assign n57038 = n3485 & ~n57037;
  assign n57039 = ~n3476 & ~n57038;
  assign n57040 = ~n32932 & ~n49184;
  assign n57041 = controllable_nhgrant0 & ~n57040;
  assign n57042 = ~n10240 & ~n57041;
  assign n57043 = ~n3281 & ~n57042;
  assign n57044 = ~n3281 & ~n57043;
  assign n57045 = n3378 & ~n57044;
  assign n57046 = ~n51771 & ~n57045;
  assign n57047 = n3492 & ~n57046;
  assign n57048 = ~n51321 & ~n57047;
  assign n57049 = n3485 & ~n57048;
  assign n57050 = ~n51478 & ~n57049;
  assign n57051 = n3476 & ~n57050;
  assign n57052 = ~n57039 & ~n57051;
  assign n57053 = n3374 & ~n57052;
  assign n57054 = ~n57032 & ~n57053;
  assign n57055 = n3655 & ~n57054;
  assign n57056 = n3378 & ~n56412;
  assign n57057 = ~n51788 & ~n57056;
  assign n57058 = n3492 & ~n57057;
  assign n57059 = n3492 & ~n57058;
  assign n57060 = n3485 & ~n57059;
  assign n57061 = n3485 & ~n57060;
  assign n57062 = ~n3476 & ~n57061;
  assign n57063 = ~n8523 & ~n57058;
  assign n57064 = n3485 & ~n57063;
  assign n57065 = ~n8689 & ~n57064;
  assign n57066 = n3476 & ~n57065;
  assign n57067 = ~n57062 & ~n57066;
  assign n57068 = ~n3374 & ~n57067;
  assign n57069 = n3378 & ~n56430;
  assign n57070 = ~n51807 & ~n57069;
  assign n57071 = n3492 & ~n57070;
  assign n57072 = n3492 & ~n57071;
  assign n57073 = n3485 & ~n57072;
  assign n57074 = n3485 & ~n57073;
  assign n57075 = ~n3476 & ~n57074;
  assign n57076 = ~n32932 & ~n49269;
  assign n57077 = controllable_nhgrant0 & ~n57076;
  assign n57078 = ~n10240 & ~n57077;
  assign n57079 = ~n3281 & ~n57078;
  assign n57080 = ~n3281 & ~n57079;
  assign n57081 = n3378 & ~n57080;
  assign n57082 = ~n51825 & ~n57081;
  assign n57083 = n3492 & ~n57082;
  assign n57084 = ~n51348 & ~n57083;
  assign n57085 = n3485 & ~n57084;
  assign n57086 = ~n51489 & ~n57085;
  assign n57087 = n3476 & ~n57086;
  assign n57088 = ~n57075 & ~n57087;
  assign n57089 = n3374 & ~n57088;
  assign n57090 = ~n57068 & ~n57089;
  assign n57091 = ~n3655 & ~n57090;
  assign n57092 = ~n57055 & ~n57091;
  assign n57093 = n3652 & ~n57092;
  assign n57094 = n3378 & ~n56466;
  assign n57095 = ~n51844 & ~n57094;
  assign n57096 = n3492 & ~n57095;
  assign n57097 = n3492 & ~n57096;
  assign n57098 = n3485 & ~n57097;
  assign n57099 = n3485 & ~n57098;
  assign n57100 = ~n3476 & ~n57099;
  assign n57101 = ~n8523 & ~n57096;
  assign n57102 = n3485 & ~n57101;
  assign n57103 = ~n8689 & ~n57102;
  assign n57104 = n3476 & ~n57103;
  assign n57105 = ~n57100 & ~n57104;
  assign n57106 = ~n3374 & ~n57105;
  assign n57107 = n3378 & ~n56484;
  assign n57108 = ~n51863 & ~n57107;
  assign n57109 = n3492 & ~n57108;
  assign n57110 = n3492 & ~n57109;
  assign n57111 = n3485 & ~n57110;
  assign n57112 = n3485 & ~n57111;
  assign n57113 = ~n3476 & ~n57112;
  assign n57114 = ~n32932 & ~n49338;
  assign n57115 = controllable_nhgrant0 & ~n57114;
  assign n57116 = ~n10240 & ~n57115;
  assign n57117 = ~n3281 & ~n57116;
  assign n57118 = ~n3281 & ~n57117;
  assign n57119 = n3378 & ~n57118;
  assign n57120 = ~n51881 & ~n57119;
  assign n57121 = n3492 & ~n57120;
  assign n57122 = ~n51377 & ~n57121;
  assign n57123 = n3485 & ~n57122;
  assign n57124 = ~n51502 & ~n57123;
  assign n57125 = n3476 & ~n57124;
  assign n57126 = ~n57113 & ~n57125;
  assign n57127 = n3374 & ~n57126;
  assign n57128 = ~n57106 & ~n57127;
  assign n57129 = n3655 & ~n57128;
  assign n57130 = n3378 & ~n56518;
  assign n57131 = ~n51898 & ~n57130;
  assign n57132 = n3492 & ~n57131;
  assign n57133 = n3492 & ~n57132;
  assign n57134 = n3485 & ~n57133;
  assign n57135 = n3485 & ~n57134;
  assign n57136 = ~n3476 & ~n57135;
  assign n57137 = ~n8523 & ~n57132;
  assign n57138 = n3485 & ~n57137;
  assign n57139 = ~n8689 & ~n57138;
  assign n57140 = n3476 & ~n57139;
  assign n57141 = ~n57136 & ~n57140;
  assign n57142 = ~n3374 & ~n57141;
  assign n57143 = n3378 & ~n56536;
  assign n57144 = ~n51917 & ~n57143;
  assign n57145 = n3492 & ~n57144;
  assign n57146 = n3492 & ~n57145;
  assign n57147 = n3485 & ~n57146;
  assign n57148 = n3485 & ~n57147;
  assign n57149 = ~n3476 & ~n57148;
  assign n57150 = ~n32932 & ~n49408;
  assign n57151 = controllable_nhgrant0 & ~n57150;
  assign n57152 = ~n10240 & ~n57151;
  assign n57153 = ~n3281 & ~n57152;
  assign n57154 = ~n3281 & ~n57153;
  assign n57155 = n3378 & ~n57154;
  assign n57156 = ~n51935 & ~n57155;
  assign n57157 = n3492 & ~n57156;
  assign n57158 = ~n51404 & ~n57157;
  assign n57159 = n3485 & ~n57158;
  assign n57160 = ~n51513 & ~n57159;
  assign n57161 = n3476 & ~n57160;
  assign n57162 = ~n57149 & ~n57161;
  assign n57163 = n3374 & ~n57162;
  assign n57164 = ~n57142 & ~n57163;
  assign n57165 = ~n3655 & ~n57164;
  assign n57166 = ~n57129 & ~n57165;
  assign n57167 = ~n3652 & ~n57166;
  assign n57168 = ~n57093 & ~n57167;
  assign n57169 = n3368 & ~n57168;
  assign n57170 = ~n57019 & ~n57169;
  assign n57171 = ~n3362 & ~n57170;
  assign n57172 = ~n56889 & ~n57171;
  assign n57173 = ~n3359 & ~n57172;
  assign n57174 = ~n56795 & ~n57173;
  assign n57175 = ~n3356 & ~n57174;
  assign n57176 = ~n56117 & ~n57175;
  assign n57177 = n3345 & ~n57176;
  assign n57178 = ~n55859 & ~n57177;
  assign n57179 = ~n3341 & ~n57178;
  assign n57180 = ~n33073 & ~n49444;
  assign n57181 = controllable_nhgrant0 & ~n57180;
  assign n57182 = ~n24376 & ~n57181;
  assign n57183 = ~n3281 & ~n57182;
  assign n57184 = ~n3783 & ~n57183;
  assign n57185 = ~n3378 & ~n57184;
  assign n57186 = ~n3378 & ~n57185;
  assign n57187 = n3492 & ~n57186;
  assign n57188 = ~n3493 & ~n57187;
  assign n57189 = n3485 & ~n57188;
  assign n57190 = ~n3486 & ~n57189;
  assign n57191 = ~n3476 & ~n57190;
  assign n57192 = ~n3281 & ~n51530;
  assign n57193 = n3378 & ~n57192;
  assign n57194 = ~n51532 & ~n57193;
  assign n57195 = n3492 & ~n57194;
  assign n57196 = ~n3493 & ~n57195;
  assign n57197 = n3485 & ~n57196;
  assign n57198 = ~n3486 & ~n57197;
  assign n57199 = n3476 & ~n57198;
  assign n57200 = ~n57191 & ~n57199;
  assign n57201 = ~n3374 & ~n57200;
  assign n57202 = ~n3950 & ~n57183;
  assign n57203 = ~n3378 & ~n57202;
  assign n57204 = ~n3378 & ~n57203;
  assign n57205 = n3492 & ~n57204;
  assign n57206 = ~n3493 & ~n57205;
  assign n57207 = n3485 & ~n57206;
  assign n57208 = ~n3486 & ~n57207;
  assign n57209 = ~n3476 & ~n57208;
  assign n57210 = ~n3281 & ~n51562;
  assign n57211 = n3378 & ~n57210;
  assign n57212 = ~n51564 & ~n57211;
  assign n57213 = n3492 & ~n57212;
  assign n57214 = ~n3493 & ~n57213;
  assign n57215 = n3485 & ~n57214;
  assign n57216 = ~n3486 & ~n57215;
  assign n57217 = n3476 & ~n57216;
  assign n57218 = ~n57209 & ~n57217;
  assign n57219 = n3374 & ~n57218;
  assign n57220 = ~n57201 & ~n57219;
  assign n57221 = n3655 & ~n57220;
  assign n57222 = ~n33073 & ~n49492;
  assign n57223 = controllable_nhgrant0 & ~n57222;
  assign n57224 = ~n24376 & ~n57223;
  assign n57225 = ~n3281 & ~n57224;
  assign n57226 = ~n3783 & ~n57225;
  assign n57227 = ~n3378 & ~n57226;
  assign n57228 = ~n3378 & ~n57227;
  assign n57229 = n3492 & ~n57228;
  assign n57230 = ~n3493 & ~n57229;
  assign n57231 = n3485 & ~n57230;
  assign n57232 = ~n3486 & ~n57231;
  assign n57233 = ~n3476 & ~n57232;
  assign n57234 = ~n3281 & ~n51579;
  assign n57235 = n3378 & ~n57234;
  assign n57236 = ~n51581 & ~n57235;
  assign n57237 = n3492 & ~n57236;
  assign n57238 = ~n3493 & ~n57237;
  assign n57239 = n3485 & ~n57238;
  assign n57240 = ~n3486 & ~n57239;
  assign n57241 = n3476 & ~n57240;
  assign n57242 = ~n57233 & ~n57241;
  assign n57243 = ~n3374 & ~n57242;
  assign n57244 = ~n3950 & ~n57225;
  assign n57245 = ~n3378 & ~n57244;
  assign n57246 = ~n3378 & ~n57245;
  assign n57247 = n3492 & ~n57246;
  assign n57248 = ~n3493 & ~n57247;
  assign n57249 = n3485 & ~n57248;
  assign n57250 = ~n3486 & ~n57249;
  assign n57251 = ~n3476 & ~n57250;
  assign n57252 = ~n3281 & ~n51611;
  assign n57253 = n3378 & ~n57252;
  assign n57254 = ~n51613 & ~n57253;
  assign n57255 = n3492 & ~n57254;
  assign n57256 = ~n3493 & ~n57255;
  assign n57257 = n3485 & ~n57256;
  assign n57258 = ~n3486 & ~n57257;
  assign n57259 = n3476 & ~n57258;
  assign n57260 = ~n57251 & ~n57259;
  assign n57261 = n3374 & ~n57260;
  assign n57262 = ~n57243 & ~n57261;
  assign n57263 = ~n3655 & ~n57262;
  assign n57264 = ~n57221 & ~n57263;
  assign n57265 = n3652 & ~n57264;
  assign n57266 = ~n33073 & ~n49542;
  assign n57267 = controllable_nhgrant0 & ~n57266;
  assign n57268 = ~n24376 & ~n57267;
  assign n57269 = ~n3281 & ~n57268;
  assign n57270 = ~n3783 & ~n57269;
  assign n57271 = ~n3378 & ~n57270;
  assign n57272 = ~n3378 & ~n57271;
  assign n57273 = n3492 & ~n57272;
  assign n57274 = ~n3493 & ~n57273;
  assign n57275 = n3485 & ~n57274;
  assign n57276 = ~n3486 & ~n57275;
  assign n57277 = ~n3476 & ~n57276;
  assign n57278 = ~n3281 & ~n51630;
  assign n57279 = n3378 & ~n57278;
  assign n57280 = ~n51632 & ~n57279;
  assign n57281 = n3492 & ~n57280;
  assign n57282 = ~n3493 & ~n57281;
  assign n57283 = n3485 & ~n57282;
  assign n57284 = ~n3486 & ~n57283;
  assign n57285 = n3476 & ~n57284;
  assign n57286 = ~n57277 & ~n57285;
  assign n57287 = ~n3374 & ~n57286;
  assign n57288 = ~n3950 & ~n57269;
  assign n57289 = ~n3378 & ~n57288;
  assign n57290 = ~n3378 & ~n57289;
  assign n57291 = n3492 & ~n57290;
  assign n57292 = ~n3493 & ~n57291;
  assign n57293 = n3485 & ~n57292;
  assign n57294 = ~n3486 & ~n57293;
  assign n57295 = ~n3476 & ~n57294;
  assign n57296 = ~n3281 & ~n51662;
  assign n57297 = n3378 & ~n57296;
  assign n57298 = ~n51664 & ~n57297;
  assign n57299 = n3492 & ~n57298;
  assign n57300 = ~n3493 & ~n57299;
  assign n57301 = n3485 & ~n57300;
  assign n57302 = ~n3486 & ~n57301;
  assign n57303 = n3476 & ~n57302;
  assign n57304 = ~n57295 & ~n57303;
  assign n57305 = n3374 & ~n57304;
  assign n57306 = ~n57287 & ~n57305;
  assign n57307 = n3655 & ~n57306;
  assign n57308 = ~n33073 & ~n49590;
  assign n57309 = controllable_nhgrant0 & ~n57308;
  assign n57310 = ~n24376 & ~n57309;
  assign n57311 = ~n3281 & ~n57310;
  assign n57312 = ~n3783 & ~n57311;
  assign n57313 = ~n3378 & ~n57312;
  assign n57314 = ~n3378 & ~n57313;
  assign n57315 = n3492 & ~n57314;
  assign n57316 = ~n3493 & ~n57315;
  assign n57317 = n3485 & ~n57316;
  assign n57318 = ~n3486 & ~n57317;
  assign n57319 = ~n3476 & ~n57318;
  assign n57320 = ~n3281 & ~n51679;
  assign n57321 = n3378 & ~n57320;
  assign n57322 = ~n51681 & ~n57321;
  assign n57323 = n3492 & ~n57322;
  assign n57324 = ~n3493 & ~n57323;
  assign n57325 = n3485 & ~n57324;
  assign n57326 = ~n3486 & ~n57325;
  assign n57327 = n3476 & ~n57326;
  assign n57328 = ~n57319 & ~n57327;
  assign n57329 = ~n3374 & ~n57328;
  assign n57330 = ~n3950 & ~n57311;
  assign n57331 = ~n3378 & ~n57330;
  assign n57332 = ~n3378 & ~n57331;
  assign n57333 = n3492 & ~n57332;
  assign n57334 = ~n3493 & ~n57333;
  assign n57335 = n3485 & ~n57334;
  assign n57336 = ~n3486 & ~n57335;
  assign n57337 = ~n3476 & ~n57336;
  assign n57338 = ~n3281 & ~n51711;
  assign n57339 = n3378 & ~n57338;
  assign n57340 = ~n51713 & ~n57339;
  assign n57341 = n3492 & ~n57340;
  assign n57342 = ~n3493 & ~n57341;
  assign n57343 = n3485 & ~n57342;
  assign n57344 = ~n3486 & ~n57343;
  assign n57345 = n3476 & ~n57344;
  assign n57346 = ~n57337 & ~n57345;
  assign n57347 = n3374 & ~n57346;
  assign n57348 = ~n57329 & ~n57347;
  assign n57349 = ~n3655 & ~n57348;
  assign n57350 = ~n57307 & ~n57349;
  assign n57351 = ~n3652 & ~n57350;
  assign n57352 = ~n57265 & ~n57351;
  assign n57353 = ~n3368 & ~n57352;
  assign n57354 = n3492 & ~n51733;
  assign n57355 = n3492 & ~n57354;
  assign n57356 = n3485 & ~n57355;
  assign n57357 = n3485 & ~n57356;
  assign n57358 = n3476 & ~n57357;
  assign n57359 = n3476 & ~n57358;
  assign n57360 = ~n3374 & ~n57359;
  assign n57361 = n3492 & ~n51770;
  assign n57362 = n3492 & ~n57361;
  assign n57363 = n3485 & ~n57362;
  assign n57364 = n3485 & ~n57363;
  assign n57365 = n3476 & ~n57364;
  assign n57366 = n3476 & ~n57365;
  assign n57367 = n3374 & ~n57366;
  assign n57368 = ~n57360 & ~n57367;
  assign n57369 = n3655 & ~n57368;
  assign n57370 = n3492 & ~n51787;
  assign n57371 = n3492 & ~n57370;
  assign n57372 = n3485 & ~n57371;
  assign n57373 = n3485 & ~n57372;
  assign n57374 = n3476 & ~n57373;
  assign n57375 = n3476 & ~n57374;
  assign n57376 = ~n3374 & ~n57375;
  assign n57377 = n3492 & ~n51824;
  assign n57378 = n3492 & ~n57377;
  assign n57379 = n3485 & ~n57378;
  assign n57380 = n3485 & ~n57379;
  assign n57381 = n3476 & ~n57380;
  assign n57382 = n3476 & ~n57381;
  assign n57383 = n3374 & ~n57382;
  assign n57384 = ~n57376 & ~n57383;
  assign n57385 = ~n3655 & ~n57384;
  assign n57386 = ~n57369 & ~n57385;
  assign n57387 = n3652 & ~n57386;
  assign n57388 = n3492 & ~n51843;
  assign n57389 = n3492 & ~n57388;
  assign n57390 = n3485 & ~n57389;
  assign n57391 = n3485 & ~n57390;
  assign n57392 = n3476 & ~n57391;
  assign n57393 = n3476 & ~n57392;
  assign n57394 = ~n3374 & ~n57393;
  assign n57395 = n3492 & ~n51880;
  assign n57396 = n3492 & ~n57395;
  assign n57397 = n3485 & ~n57396;
  assign n57398 = n3485 & ~n57397;
  assign n57399 = n3476 & ~n57398;
  assign n57400 = n3476 & ~n57399;
  assign n57401 = n3374 & ~n57400;
  assign n57402 = ~n57394 & ~n57401;
  assign n57403 = n3655 & ~n57402;
  assign n57404 = n3492 & ~n51897;
  assign n57405 = n3492 & ~n57404;
  assign n57406 = n3485 & ~n57405;
  assign n57407 = n3485 & ~n57406;
  assign n57408 = n3476 & ~n57407;
  assign n57409 = n3476 & ~n57408;
  assign n57410 = ~n3374 & ~n57409;
  assign n57411 = n3492 & ~n51934;
  assign n57412 = n3492 & ~n57411;
  assign n57413 = n3485 & ~n57412;
  assign n57414 = n3485 & ~n57413;
  assign n57415 = n3476 & ~n57414;
  assign n57416 = n3476 & ~n57415;
  assign n57417 = n3374 & ~n57416;
  assign n57418 = ~n57410 & ~n57417;
  assign n57419 = ~n3655 & ~n57418;
  assign n57420 = ~n57403 & ~n57419;
  assign n57421 = ~n3652 & ~n57420;
  assign n57422 = ~n57387 & ~n57421;
  assign n57423 = n3368 & ~n57422;
  assign n57424 = ~n57353 & ~n57423;
  assign n57425 = ~n3362 & ~n57424;
  assign n57426 = ~n3362 & ~n57425;
  assign n57427 = ~n3359 & ~n57426;
  assign n57428 = ~n3359 & ~n57427;
  assign n57429 = n3356 & ~n57428;
  assign n57430 = n3492 & ~n51531;
  assign n57431 = ~n3631 & ~n57430;
  assign n57432 = n3485 & ~n57431;
  assign n57433 = ~n3630 & ~n57432;
  assign n57434 = ~n3374 & ~n57433;
  assign n57435 = n3492 & ~n51550;
  assign n57436 = ~n3631 & ~n57435;
  assign n57437 = n3485 & ~n57436;
  assign n57438 = ~n3630 & ~n57437;
  assign n57439 = ~n3476 & ~n57438;
  assign n57440 = n3492 & ~n51563;
  assign n57441 = ~n3631 & ~n57440;
  assign n57442 = n3485 & ~n57441;
  assign n57443 = ~n3630 & ~n57442;
  assign n57444 = n3476 & ~n57443;
  assign n57445 = ~n57439 & ~n57444;
  assign n57446 = n3374 & ~n57445;
  assign n57447 = ~n57434 & ~n57446;
  assign n57448 = n3655 & ~n57447;
  assign n57449 = n3492 & ~n51580;
  assign n57450 = ~n3631 & ~n57449;
  assign n57451 = n3485 & ~n57450;
  assign n57452 = ~n3630 & ~n57451;
  assign n57453 = ~n3374 & ~n57452;
  assign n57454 = n3492 & ~n51599;
  assign n57455 = ~n3631 & ~n57454;
  assign n57456 = n3485 & ~n57455;
  assign n57457 = ~n3630 & ~n57456;
  assign n57458 = ~n3476 & ~n57457;
  assign n57459 = n3492 & ~n51612;
  assign n57460 = ~n3631 & ~n57459;
  assign n57461 = n3485 & ~n57460;
  assign n57462 = ~n3630 & ~n57461;
  assign n57463 = n3476 & ~n57462;
  assign n57464 = ~n57458 & ~n57463;
  assign n57465 = n3374 & ~n57464;
  assign n57466 = ~n57453 & ~n57465;
  assign n57467 = ~n3655 & ~n57466;
  assign n57468 = ~n57448 & ~n57467;
  assign n57469 = n3652 & ~n57468;
  assign n57470 = n3492 & ~n51631;
  assign n57471 = ~n3631 & ~n57470;
  assign n57472 = n3485 & ~n57471;
  assign n57473 = ~n3630 & ~n57472;
  assign n57474 = ~n3374 & ~n57473;
  assign n57475 = n3492 & ~n51650;
  assign n57476 = ~n3631 & ~n57475;
  assign n57477 = n3485 & ~n57476;
  assign n57478 = ~n3630 & ~n57477;
  assign n57479 = ~n3476 & ~n57478;
  assign n57480 = n3492 & ~n51663;
  assign n57481 = ~n3631 & ~n57480;
  assign n57482 = n3485 & ~n57481;
  assign n57483 = ~n3630 & ~n57482;
  assign n57484 = n3476 & ~n57483;
  assign n57485 = ~n57479 & ~n57484;
  assign n57486 = n3374 & ~n57485;
  assign n57487 = ~n57474 & ~n57486;
  assign n57488 = n3655 & ~n57487;
  assign n57489 = n3492 & ~n51680;
  assign n57490 = ~n3631 & ~n57489;
  assign n57491 = n3485 & ~n57490;
  assign n57492 = ~n3630 & ~n57491;
  assign n57493 = ~n3374 & ~n57492;
  assign n57494 = n3492 & ~n51699;
  assign n57495 = ~n3631 & ~n57494;
  assign n57496 = n3485 & ~n57495;
  assign n57497 = ~n3630 & ~n57496;
  assign n57498 = ~n3476 & ~n57497;
  assign n57499 = n3492 & ~n51712;
  assign n57500 = ~n3631 & ~n57499;
  assign n57501 = n3485 & ~n57500;
  assign n57502 = ~n3630 & ~n57501;
  assign n57503 = n3476 & ~n57502;
  assign n57504 = ~n57498 & ~n57503;
  assign n57505 = n3374 & ~n57504;
  assign n57506 = ~n57493 & ~n57505;
  assign n57507 = ~n3655 & ~n57506;
  assign n57508 = ~n57488 & ~n57507;
  assign n57509 = ~n3652 & ~n57508;
  assign n57510 = ~n57469 & ~n57509;
  assign n57511 = ~n3368 & ~n57510;
  assign n57512 = ~n3374 & ~n57357;
  assign n57513 = n3492 & ~n51752;
  assign n57514 = n3492 & ~n57513;
  assign n57515 = n3485 & ~n57514;
  assign n57516 = n3485 & ~n57515;
  assign n57517 = ~n3476 & ~n57516;
  assign n57518 = ~n57365 & ~n57517;
  assign n57519 = n3374 & ~n57518;
  assign n57520 = ~n57512 & ~n57519;
  assign n57521 = n3655 & ~n57520;
  assign n57522 = ~n3374 & ~n57373;
  assign n57523 = n3492 & ~n51806;
  assign n57524 = n3492 & ~n57523;
  assign n57525 = n3485 & ~n57524;
  assign n57526 = n3485 & ~n57525;
  assign n57527 = ~n3476 & ~n57526;
  assign n57528 = ~n57381 & ~n57527;
  assign n57529 = n3374 & ~n57528;
  assign n57530 = ~n57522 & ~n57529;
  assign n57531 = ~n3655 & ~n57530;
  assign n57532 = ~n57521 & ~n57531;
  assign n57533 = n3652 & ~n57532;
  assign n57534 = ~n3374 & ~n57391;
  assign n57535 = n3492 & ~n51862;
  assign n57536 = n3492 & ~n57535;
  assign n57537 = n3485 & ~n57536;
  assign n57538 = n3485 & ~n57537;
  assign n57539 = ~n3476 & ~n57538;
  assign n57540 = ~n57399 & ~n57539;
  assign n57541 = n3374 & ~n57540;
  assign n57542 = ~n57534 & ~n57541;
  assign n57543 = n3655 & ~n57542;
  assign n57544 = ~n3374 & ~n57407;
  assign n57545 = n3492 & ~n51916;
  assign n57546 = n3492 & ~n57545;
  assign n57547 = n3485 & ~n57546;
  assign n57548 = n3485 & ~n57547;
  assign n57549 = ~n3476 & ~n57548;
  assign n57550 = ~n57415 & ~n57549;
  assign n57551 = n3374 & ~n57550;
  assign n57552 = ~n57544 & ~n57551;
  assign n57553 = ~n3655 & ~n57552;
  assign n57554 = ~n57543 & ~n57553;
  assign n57555 = ~n3652 & ~n57554;
  assign n57556 = ~n57533 & ~n57555;
  assign n57557 = n3368 & ~n57556;
  assign n57558 = ~n57511 & ~n57557;
  assign n57559 = n3362 & ~n57558;
  assign n57560 = ~n3476 & ~n57433;
  assign n57561 = ~n54016 & ~n57432;
  assign n57562 = n3476 & ~n57561;
  assign n57563 = ~n57560 & ~n57562;
  assign n57564 = ~n3374 & ~n57563;
  assign n57565 = ~n54016 & ~n57442;
  assign n57566 = n3476 & ~n57565;
  assign n57567 = ~n57439 & ~n57566;
  assign n57568 = n3374 & ~n57567;
  assign n57569 = ~n57564 & ~n57568;
  assign n57570 = n3655 & ~n57569;
  assign n57571 = ~n3476 & ~n57452;
  assign n57572 = ~n54041 & ~n57451;
  assign n57573 = n3476 & ~n57572;
  assign n57574 = ~n57571 & ~n57573;
  assign n57575 = ~n3374 & ~n57574;
  assign n57576 = ~n54041 & ~n57461;
  assign n57577 = n3476 & ~n57576;
  assign n57578 = ~n57458 & ~n57577;
  assign n57579 = n3374 & ~n57578;
  assign n57580 = ~n57575 & ~n57579;
  assign n57581 = ~n3655 & ~n57580;
  assign n57582 = ~n57570 & ~n57581;
  assign n57583 = n3652 & ~n57582;
  assign n57584 = ~n3476 & ~n57473;
  assign n57585 = ~n55363 & ~n57472;
  assign n57586 = n3476 & ~n57585;
  assign n57587 = ~n57584 & ~n57586;
  assign n57588 = ~n3374 & ~n57587;
  assign n57589 = ~n55363 & ~n57482;
  assign n57590 = n3476 & ~n57589;
  assign n57591 = ~n57479 & ~n57590;
  assign n57592 = n3374 & ~n57591;
  assign n57593 = ~n57588 & ~n57592;
  assign n57594 = n3655 & ~n57593;
  assign n57595 = ~n3476 & ~n57492;
  assign n57596 = ~n8310 & ~n51279;
  assign n57597 = ~n3485 & ~n57596;
  assign n57598 = ~n57491 & ~n57597;
  assign n57599 = n3476 & ~n57598;
  assign n57600 = ~n57595 & ~n57599;
  assign n57601 = ~n3374 & ~n57600;
  assign n57602 = ~n57501 & ~n57597;
  assign n57603 = n3476 & ~n57602;
  assign n57604 = ~n57498 & ~n57603;
  assign n57605 = n3374 & ~n57604;
  assign n57606 = ~n57601 & ~n57605;
  assign n57607 = ~n3655 & ~n57606;
  assign n57608 = ~n57594 & ~n57607;
  assign n57609 = ~n3652 & ~n57608;
  assign n57610 = ~n57583 & ~n57609;
  assign n57611 = ~n3368 & ~n57610;
  assign n57612 = ~n3476 & ~n57357;
  assign n57613 = ~n8525 & ~n57356;
  assign n57614 = n3476 & ~n57613;
  assign n57615 = ~n57612 & ~n57614;
  assign n57616 = ~n3374 & ~n57615;
  assign n57617 = ~n54135 & ~n57363;
  assign n57618 = n3476 & ~n57617;
  assign n57619 = ~n57517 & ~n57618;
  assign n57620 = n3374 & ~n57619;
  assign n57621 = ~n57616 & ~n57620;
  assign n57622 = n3655 & ~n57621;
  assign n57623 = ~n3476 & ~n57373;
  assign n57624 = ~n8525 & ~n57372;
  assign n57625 = n3476 & ~n57624;
  assign n57626 = ~n57623 & ~n57625;
  assign n57627 = ~n3374 & ~n57626;
  assign n57628 = ~n54160 & ~n57379;
  assign n57629 = n3476 & ~n57628;
  assign n57630 = ~n57527 & ~n57629;
  assign n57631 = n3374 & ~n57630;
  assign n57632 = ~n57627 & ~n57631;
  assign n57633 = ~n3655 & ~n57632;
  assign n57634 = ~n57622 & ~n57633;
  assign n57635 = n3652 & ~n57634;
  assign n57636 = ~n3476 & ~n57391;
  assign n57637 = ~n8525 & ~n57390;
  assign n57638 = n3476 & ~n57637;
  assign n57639 = ~n57636 & ~n57638;
  assign n57640 = ~n3374 & ~n57639;
  assign n57641 = ~n55469 & ~n57397;
  assign n57642 = n3476 & ~n57641;
  assign n57643 = ~n57539 & ~n57642;
  assign n57644 = n3374 & ~n57643;
  assign n57645 = ~n57640 & ~n57644;
  assign n57646 = n3655 & ~n57645;
  assign n57647 = ~n3476 & ~n57407;
  assign n57648 = ~n8525 & ~n57406;
  assign n57649 = n3476 & ~n57648;
  assign n57650 = ~n57647 & ~n57649;
  assign n57651 = ~n3374 & ~n57650;
  assign n57652 = ~n3492 & ~n51404;
  assign n57653 = ~n3485 & ~n57652;
  assign n57654 = ~n57413 & ~n57653;
  assign n57655 = n3476 & ~n57654;
  assign n57656 = ~n57549 & ~n57655;
  assign n57657 = n3374 & ~n57656;
  assign n57658 = ~n57651 & ~n57657;
  assign n57659 = ~n3655 & ~n57658;
  assign n57660 = ~n57646 & ~n57659;
  assign n57661 = ~n3652 & ~n57660;
  assign n57662 = ~n57635 & ~n57661;
  assign n57663 = n3368 & ~n57662;
  assign n57664 = ~n57611 & ~n57663;
  assign n57665 = ~n3362 & ~n57664;
  assign n57666 = ~n57559 & ~n57665;
  assign n57667 = n3359 & ~n57666;
  assign n57668 = ~n51424 & ~n57432;
  assign n57669 = n3476 & ~n57668;
  assign n57670 = ~n57560 & ~n57669;
  assign n57671 = ~n3374 & ~n57670;
  assign n57672 = ~n51424 & ~n57442;
  assign n57673 = n3476 & ~n57672;
  assign n57674 = ~n57439 & ~n57673;
  assign n57675 = n3374 & ~n57674;
  assign n57676 = ~n57671 & ~n57675;
  assign n57677 = n3655 & ~n57676;
  assign n57678 = ~n51435 & ~n57451;
  assign n57679 = n3476 & ~n57678;
  assign n57680 = ~n57571 & ~n57679;
  assign n57681 = ~n3374 & ~n57680;
  assign n57682 = ~n51435 & ~n57461;
  assign n57683 = n3476 & ~n57682;
  assign n57684 = ~n57458 & ~n57683;
  assign n57685 = n3374 & ~n57684;
  assign n57686 = ~n57681 & ~n57685;
  assign n57687 = ~n3655 & ~n57686;
  assign n57688 = ~n57677 & ~n57687;
  assign n57689 = n3652 & ~n57688;
  assign n57690 = ~n51448 & ~n57472;
  assign n57691 = n3476 & ~n57690;
  assign n57692 = ~n57584 & ~n57691;
  assign n57693 = ~n3374 & ~n57692;
  assign n57694 = ~n51448 & ~n57482;
  assign n57695 = n3476 & ~n57694;
  assign n57696 = ~n57479 & ~n57695;
  assign n57697 = n3374 & ~n57696;
  assign n57698 = ~n57693 & ~n57697;
  assign n57699 = n3655 & ~n57698;
  assign n57700 = ~n51459 & ~n57491;
  assign n57701 = n3476 & ~n57700;
  assign n57702 = ~n57595 & ~n57701;
  assign n57703 = ~n3374 & ~n57702;
  assign n57704 = ~n51459 & ~n57501;
  assign n57705 = n3476 & ~n57704;
  assign n57706 = ~n57498 & ~n57705;
  assign n57707 = n3374 & ~n57706;
  assign n57708 = ~n57703 & ~n57707;
  assign n57709 = ~n3655 & ~n57708;
  assign n57710 = ~n57699 & ~n57709;
  assign n57711 = ~n3652 & ~n57710;
  assign n57712 = ~n57689 & ~n57711;
  assign n57713 = ~n3368 & ~n57712;
  assign n57714 = ~n8689 & ~n57356;
  assign n57715 = n3476 & ~n57714;
  assign n57716 = ~n57612 & ~n57715;
  assign n57717 = ~n3374 & ~n57716;
  assign n57718 = ~n51478 & ~n57363;
  assign n57719 = n3476 & ~n57718;
  assign n57720 = ~n57517 & ~n57719;
  assign n57721 = n3374 & ~n57720;
  assign n57722 = ~n57717 & ~n57721;
  assign n57723 = n3655 & ~n57722;
  assign n57724 = ~n8689 & ~n57372;
  assign n57725 = n3476 & ~n57724;
  assign n57726 = ~n57623 & ~n57725;
  assign n57727 = ~n3374 & ~n57726;
  assign n57728 = ~n51489 & ~n57379;
  assign n57729 = n3476 & ~n57728;
  assign n57730 = ~n57527 & ~n57729;
  assign n57731 = n3374 & ~n57730;
  assign n57732 = ~n57727 & ~n57731;
  assign n57733 = ~n3655 & ~n57732;
  assign n57734 = ~n57723 & ~n57733;
  assign n57735 = n3652 & ~n57734;
  assign n57736 = ~n8689 & ~n57390;
  assign n57737 = n3476 & ~n57736;
  assign n57738 = ~n57636 & ~n57737;
  assign n57739 = ~n3374 & ~n57738;
  assign n57740 = ~n51502 & ~n57397;
  assign n57741 = n3476 & ~n57740;
  assign n57742 = ~n57539 & ~n57741;
  assign n57743 = n3374 & ~n57742;
  assign n57744 = ~n57739 & ~n57743;
  assign n57745 = n3655 & ~n57744;
  assign n57746 = ~n8689 & ~n57406;
  assign n57747 = n3476 & ~n57746;
  assign n57748 = ~n57647 & ~n57747;
  assign n57749 = ~n3374 & ~n57748;
  assign n57750 = ~n51513 & ~n57413;
  assign n57751 = n3476 & ~n57750;
  assign n57752 = ~n57549 & ~n57751;
  assign n57753 = n3374 & ~n57752;
  assign n57754 = ~n57749 & ~n57753;
  assign n57755 = ~n3655 & ~n57754;
  assign n57756 = ~n57745 & ~n57755;
  assign n57757 = ~n3652 & ~n57756;
  assign n57758 = ~n57735 & ~n57757;
  assign n57759 = n3368 & ~n57758;
  assign n57760 = ~n57713 & ~n57759;
  assign n57761 = n3362 & ~n57760;
  assign n57762 = ~n51148 & ~n57430;
  assign n57763 = n3485 & ~n57762;
  assign n57764 = ~n51424 & ~n57763;
  assign n57765 = n3476 & ~n57764;
  assign n57766 = ~n57560 & ~n57765;
  assign n57767 = ~n3374 & ~n57766;
  assign n57768 = ~n51148 & ~n57440;
  assign n57769 = n3485 & ~n57768;
  assign n57770 = ~n51424 & ~n57769;
  assign n57771 = n3476 & ~n57770;
  assign n57772 = ~n57439 & ~n57771;
  assign n57773 = n3374 & ~n57772;
  assign n57774 = ~n57767 & ~n57773;
  assign n57775 = n3655 & ~n57774;
  assign n57776 = ~n51191 & ~n57449;
  assign n57777 = n3485 & ~n57776;
  assign n57778 = ~n51435 & ~n57777;
  assign n57779 = n3476 & ~n57778;
  assign n57780 = ~n57571 & ~n57779;
  assign n57781 = ~n3374 & ~n57780;
  assign n57782 = ~n51191 & ~n57459;
  assign n57783 = n3485 & ~n57782;
  assign n57784 = ~n51435 & ~n57783;
  assign n57785 = n3476 & ~n57784;
  assign n57786 = ~n57458 & ~n57785;
  assign n57787 = n3374 & ~n57786;
  assign n57788 = ~n57781 & ~n57787;
  assign n57789 = ~n3655 & ~n57788;
  assign n57790 = ~n57775 & ~n57789;
  assign n57791 = n3652 & ~n57790;
  assign n57792 = ~n51236 & ~n57470;
  assign n57793 = n3485 & ~n57792;
  assign n57794 = ~n51448 & ~n57793;
  assign n57795 = n3476 & ~n57794;
  assign n57796 = ~n57584 & ~n57795;
  assign n57797 = ~n3374 & ~n57796;
  assign n57798 = ~n51236 & ~n57480;
  assign n57799 = n3485 & ~n57798;
  assign n57800 = ~n51448 & ~n57799;
  assign n57801 = n3476 & ~n57800;
  assign n57802 = ~n57479 & ~n57801;
  assign n57803 = n3374 & ~n57802;
  assign n57804 = ~n57797 & ~n57803;
  assign n57805 = n3655 & ~n57804;
  assign n57806 = ~n51279 & ~n57489;
  assign n57807 = n3485 & ~n57806;
  assign n57808 = ~n51459 & ~n57807;
  assign n57809 = n3476 & ~n57808;
  assign n57810 = ~n57595 & ~n57809;
  assign n57811 = ~n3374 & ~n57810;
  assign n57812 = ~n51279 & ~n57499;
  assign n57813 = n3485 & ~n57812;
  assign n57814 = ~n51459 & ~n57813;
  assign n57815 = n3476 & ~n57814;
  assign n57816 = ~n57498 & ~n57815;
  assign n57817 = n3374 & ~n57816;
  assign n57818 = ~n57811 & ~n57817;
  assign n57819 = ~n3655 & ~n57818;
  assign n57820 = ~n57805 & ~n57819;
  assign n57821 = ~n3652 & ~n57820;
  assign n57822 = ~n57791 & ~n57821;
  assign n57823 = ~n3368 & ~n57822;
  assign n57824 = ~n8523 & ~n57354;
  assign n57825 = n3485 & ~n57824;
  assign n57826 = ~n8689 & ~n57825;
  assign n57827 = n3476 & ~n57826;
  assign n57828 = ~n57612 & ~n57827;
  assign n57829 = ~n3374 & ~n57828;
  assign n57830 = ~n51321 & ~n57361;
  assign n57831 = n3485 & ~n57830;
  assign n57832 = ~n51478 & ~n57831;
  assign n57833 = n3476 & ~n57832;
  assign n57834 = ~n57517 & ~n57833;
  assign n57835 = n3374 & ~n57834;
  assign n57836 = ~n57829 & ~n57835;
  assign n57837 = n3655 & ~n57836;
  assign n57838 = ~n8523 & ~n57370;
  assign n57839 = n3485 & ~n57838;
  assign n57840 = ~n8689 & ~n57839;
  assign n57841 = n3476 & ~n57840;
  assign n57842 = ~n57623 & ~n57841;
  assign n57843 = ~n3374 & ~n57842;
  assign n57844 = ~n51348 & ~n57377;
  assign n57845 = n3485 & ~n57844;
  assign n57846 = ~n51489 & ~n57845;
  assign n57847 = n3476 & ~n57846;
  assign n57848 = ~n57527 & ~n57847;
  assign n57849 = n3374 & ~n57848;
  assign n57850 = ~n57843 & ~n57849;
  assign n57851 = ~n3655 & ~n57850;
  assign n57852 = ~n57837 & ~n57851;
  assign n57853 = n3652 & ~n57852;
  assign n57854 = ~n8523 & ~n57388;
  assign n57855 = n3485 & ~n57854;
  assign n57856 = ~n8689 & ~n57855;
  assign n57857 = n3476 & ~n57856;
  assign n57858 = ~n57636 & ~n57857;
  assign n57859 = ~n3374 & ~n57858;
  assign n57860 = ~n51377 & ~n57395;
  assign n57861 = n3485 & ~n57860;
  assign n57862 = ~n51502 & ~n57861;
  assign n57863 = n3476 & ~n57862;
  assign n57864 = ~n57539 & ~n57863;
  assign n57865 = n3374 & ~n57864;
  assign n57866 = ~n57859 & ~n57865;
  assign n57867 = n3655 & ~n57866;
  assign n57868 = ~n8523 & ~n57404;
  assign n57869 = n3485 & ~n57868;
  assign n57870 = ~n8689 & ~n57869;
  assign n57871 = n3476 & ~n57870;
  assign n57872 = ~n57647 & ~n57871;
  assign n57873 = ~n3374 & ~n57872;
  assign n57874 = ~n51404 & ~n57411;
  assign n57875 = n3485 & ~n57874;
  assign n57876 = ~n51513 & ~n57875;
  assign n57877 = n3476 & ~n57876;
  assign n57878 = ~n57549 & ~n57877;
  assign n57879 = n3374 & ~n57878;
  assign n57880 = ~n57873 & ~n57879;
  assign n57881 = ~n3655 & ~n57880;
  assign n57882 = ~n57867 & ~n57881;
  assign n57883 = ~n3652 & ~n57882;
  assign n57884 = ~n57853 & ~n57883;
  assign n57885 = n3368 & ~n57884;
  assign n57886 = ~n57823 & ~n57885;
  assign n57887 = ~n3362 & ~n57886;
  assign n57888 = ~n57761 & ~n57887;
  assign n57889 = ~n3359 & ~n57888;
  assign n57890 = ~n57667 & ~n57889;
  assign n57891 = ~n3356 & ~n57890;
  assign n57892 = ~n57429 & ~n57891;
  assign n57893 = ~n3345 & ~n57892;
  assign n57894 = ~n3378 & ~n51532;
  assign n57895 = n3492 & ~n57894;
  assign n57896 = ~n3493 & ~n57895;
  assign n57897 = n3485 & ~n57896;
  assign n57898 = ~n3486 & ~n57897;
  assign n57899 = ~n3476 & ~n57898;
  assign n57900 = ~n3378 & ~n51147;
  assign n57901 = ~n3378 & ~n57900;
  assign n57902 = ~n3485 & ~n57901;
  assign n57903 = ~n3492 & ~n57901;
  assign n57904 = ~n57895 & ~n57903;
  assign n57905 = n3485 & ~n57904;
  assign n57906 = ~n57902 & ~n57905;
  assign n57907 = n3476 & ~n57906;
  assign n57908 = ~n57899 & ~n57907;
  assign n57909 = ~n3374 & ~n57908;
  assign n57910 = ~n3281 & ~n51549;
  assign n57911 = n3378 & ~n57910;
  assign n57912 = ~n51551 & ~n57911;
  assign n57913 = n3492 & ~n57912;
  assign n57914 = ~n25115 & ~n57913;
  assign n57915 = n3485 & ~n57914;
  assign n57916 = ~n25114 & ~n57915;
  assign n57917 = ~n3476 & ~n57916;
  assign n57918 = n3378 & ~n51320;
  assign n57919 = ~n57900 & ~n57918;
  assign n57920 = ~n3485 & ~n57919;
  assign n57921 = ~n3492 & ~n57919;
  assign n57922 = ~n57213 & ~n57921;
  assign n57923 = n3485 & ~n57922;
  assign n57924 = ~n57920 & ~n57923;
  assign n57925 = n3476 & ~n57924;
  assign n57926 = ~n57917 & ~n57925;
  assign n57927 = n3374 & ~n57926;
  assign n57928 = ~n57909 & ~n57927;
  assign n57929 = n3655 & ~n57928;
  assign n57930 = ~n3378 & ~n51581;
  assign n57931 = n3492 & ~n57930;
  assign n57932 = ~n3493 & ~n57931;
  assign n57933 = n3485 & ~n57932;
  assign n57934 = ~n3486 & ~n57933;
  assign n57935 = ~n3476 & ~n57934;
  assign n57936 = ~n3378 & ~n51190;
  assign n57937 = ~n3378 & ~n57936;
  assign n57938 = ~n3485 & ~n57937;
  assign n57939 = ~n3492 & ~n57937;
  assign n57940 = ~n57931 & ~n57939;
  assign n57941 = n3485 & ~n57940;
  assign n57942 = ~n57938 & ~n57941;
  assign n57943 = n3476 & ~n57942;
  assign n57944 = ~n57935 & ~n57943;
  assign n57945 = ~n3374 & ~n57944;
  assign n57946 = ~n3281 & ~n51598;
  assign n57947 = n3378 & ~n57946;
  assign n57948 = ~n51600 & ~n57947;
  assign n57949 = n3492 & ~n57948;
  assign n57950 = ~n25115 & ~n57949;
  assign n57951 = n3485 & ~n57950;
  assign n57952 = ~n25114 & ~n57951;
  assign n57953 = ~n3476 & ~n57952;
  assign n57954 = n3378 & ~n51347;
  assign n57955 = ~n57936 & ~n57954;
  assign n57956 = ~n3485 & ~n57955;
  assign n57957 = ~n3492 & ~n57955;
  assign n57958 = ~n57255 & ~n57957;
  assign n57959 = n3485 & ~n57958;
  assign n57960 = ~n57956 & ~n57959;
  assign n57961 = n3476 & ~n57960;
  assign n57962 = ~n57953 & ~n57961;
  assign n57963 = n3374 & ~n57962;
  assign n57964 = ~n57945 & ~n57963;
  assign n57965 = ~n3655 & ~n57964;
  assign n57966 = ~n57929 & ~n57965;
  assign n57967 = n3652 & ~n57966;
  assign n57968 = ~n3378 & ~n51632;
  assign n57969 = n3492 & ~n57968;
  assign n57970 = ~n3493 & ~n57969;
  assign n57971 = n3485 & ~n57970;
  assign n57972 = ~n3486 & ~n57971;
  assign n57973 = ~n3476 & ~n57972;
  assign n57974 = ~n3378 & ~n51235;
  assign n57975 = ~n3378 & ~n57974;
  assign n57976 = ~n3485 & ~n57975;
  assign n57977 = ~n3492 & ~n57975;
  assign n57978 = ~n57969 & ~n57977;
  assign n57979 = n3485 & ~n57978;
  assign n57980 = ~n57976 & ~n57979;
  assign n57981 = n3476 & ~n57980;
  assign n57982 = ~n57973 & ~n57981;
  assign n57983 = ~n3374 & ~n57982;
  assign n57984 = ~n3281 & ~n51649;
  assign n57985 = n3378 & ~n57984;
  assign n57986 = ~n51651 & ~n57985;
  assign n57987 = n3492 & ~n57986;
  assign n57988 = ~n25115 & ~n57987;
  assign n57989 = n3485 & ~n57988;
  assign n57990 = ~n25114 & ~n57989;
  assign n57991 = ~n3476 & ~n57990;
  assign n57992 = n3378 & ~n51376;
  assign n57993 = ~n57974 & ~n57992;
  assign n57994 = ~n3485 & ~n57993;
  assign n57995 = ~n3492 & ~n57993;
  assign n57996 = ~n57299 & ~n57995;
  assign n57997 = n3485 & ~n57996;
  assign n57998 = ~n57994 & ~n57997;
  assign n57999 = n3476 & ~n57998;
  assign n58000 = ~n57991 & ~n57999;
  assign n58001 = n3374 & ~n58000;
  assign n58002 = ~n57983 & ~n58001;
  assign n58003 = n3655 & ~n58002;
  assign n58004 = ~n3378 & ~n51681;
  assign n58005 = n3492 & ~n58004;
  assign n58006 = ~n3493 & ~n58005;
  assign n58007 = n3485 & ~n58006;
  assign n58008 = ~n3486 & ~n58007;
  assign n58009 = ~n3476 & ~n58008;
  assign n58010 = ~n3378 & ~n51278;
  assign n58011 = ~n3378 & ~n58010;
  assign n58012 = ~n3485 & ~n58011;
  assign n58013 = ~n3492 & ~n58011;
  assign n58014 = ~n58005 & ~n58013;
  assign n58015 = n3485 & ~n58014;
  assign n58016 = ~n58012 & ~n58015;
  assign n58017 = n3476 & ~n58016;
  assign n58018 = ~n58009 & ~n58017;
  assign n58019 = ~n3374 & ~n58018;
  assign n58020 = ~n3281 & ~n51698;
  assign n58021 = n3378 & ~n58020;
  assign n58022 = ~n51700 & ~n58021;
  assign n58023 = n3492 & ~n58022;
  assign n58024 = ~n25115 & ~n58023;
  assign n58025 = n3485 & ~n58024;
  assign n58026 = ~n25114 & ~n58025;
  assign n58027 = ~n3476 & ~n58026;
  assign n58028 = n3378 & ~n51403;
  assign n58029 = ~n58010 & ~n58028;
  assign n58030 = ~n3485 & ~n58029;
  assign n58031 = ~n3492 & ~n58029;
  assign n58032 = ~n57341 & ~n58031;
  assign n58033 = n3485 & ~n58032;
  assign n58034 = ~n58030 & ~n58033;
  assign n58035 = n3476 & ~n58034;
  assign n58036 = ~n58027 & ~n58035;
  assign n58037 = n3374 & ~n58036;
  assign n58038 = ~n58019 & ~n58037;
  assign n58039 = ~n3655 & ~n58038;
  assign n58040 = ~n58003 & ~n58039;
  assign n58041 = ~n3652 & ~n58040;
  assign n58042 = ~n57967 & ~n58041;
  assign n58043 = ~n3368 & ~n58042;
  assign n58044 = ~n3378 & ~n51734;
  assign n58045 = n3492 & ~n58044;
  assign n58046 = n3492 & ~n58045;
  assign n58047 = n3485 & ~n58046;
  assign n58048 = n3485 & ~n58047;
  assign n58049 = ~n3476 & ~n58048;
  assign n58050 = ~n25259 & ~n58045;
  assign n58051 = n3485 & ~n58050;
  assign n58052 = ~n25258 & ~n58051;
  assign n58053 = n3476 & ~n58052;
  assign n58054 = ~n58049 & ~n58053;
  assign n58055 = ~n3374 & ~n58054;
  assign n58056 = ~n57835 & ~n58055;
  assign n58057 = n3655 & ~n58056;
  assign n58058 = ~n3378 & ~n51788;
  assign n58059 = n3492 & ~n58058;
  assign n58060 = n3492 & ~n58059;
  assign n58061 = n3485 & ~n58060;
  assign n58062 = n3485 & ~n58061;
  assign n58063 = ~n3476 & ~n58062;
  assign n58064 = ~n25259 & ~n58059;
  assign n58065 = n3485 & ~n58064;
  assign n58066 = ~n25258 & ~n58065;
  assign n58067 = n3476 & ~n58066;
  assign n58068 = ~n58063 & ~n58067;
  assign n58069 = ~n3374 & ~n58068;
  assign n58070 = ~n57849 & ~n58069;
  assign n58071 = ~n3655 & ~n58070;
  assign n58072 = ~n58057 & ~n58071;
  assign n58073 = n3652 & ~n58072;
  assign n58074 = ~n3378 & ~n51844;
  assign n58075 = n3492 & ~n58074;
  assign n58076 = n3492 & ~n58075;
  assign n58077 = n3485 & ~n58076;
  assign n58078 = n3485 & ~n58077;
  assign n58079 = ~n3476 & ~n58078;
  assign n58080 = ~n25259 & ~n58075;
  assign n58081 = n3485 & ~n58080;
  assign n58082 = ~n25258 & ~n58081;
  assign n58083 = n3476 & ~n58082;
  assign n58084 = ~n58079 & ~n58083;
  assign n58085 = ~n3374 & ~n58084;
  assign n58086 = ~n57865 & ~n58085;
  assign n58087 = n3655 & ~n58086;
  assign n58088 = ~n3378 & ~n51898;
  assign n58089 = n3492 & ~n58088;
  assign n58090 = n3492 & ~n58089;
  assign n58091 = n3485 & ~n58090;
  assign n58092 = n3485 & ~n58091;
  assign n58093 = ~n3476 & ~n58092;
  assign n58094 = ~n25259 & ~n58089;
  assign n58095 = n3485 & ~n58094;
  assign n58096 = ~n25258 & ~n58095;
  assign n58097 = n3476 & ~n58096;
  assign n58098 = ~n58093 & ~n58097;
  assign n58099 = ~n3374 & ~n58098;
  assign n58100 = ~n57879 & ~n58099;
  assign n58101 = ~n3655 & ~n58100;
  assign n58102 = ~n58087 & ~n58101;
  assign n58103 = ~n3652 & ~n58102;
  assign n58104 = ~n58073 & ~n58103;
  assign n58105 = n3368 & ~n58104;
  assign n58106 = ~n58043 & ~n58105;
  assign n58107 = ~n3362 & ~n58106;
  assign n58108 = ~n3362 & ~n58107;
  assign n58109 = ~n3359 & ~n58108;
  assign n58110 = ~n3359 & ~n58109;
  assign n58111 = n3356 & ~n58110;
  assign n58112 = ~n3356 & ~n57886;
  assign n58113 = ~n58111 & ~n58112;
  assign n58114 = n3345 & ~n58113;
  assign n58115 = ~n57893 & ~n58114;
  assign n58116 = n3341 & ~n58115;
  assign n58117 = ~n57179 & ~n58116;
  assign n58118 = n3337 & ~n58117;
  assign n58119 = ~n54615 & ~n58118;
  assign n58120 = ~n3280 & ~n58119;
  assign n58121 = ~n50399 & ~n58120;
  assign n58122 = n3277 & n58121;
  assign n58123 = n3277 & ~n58122;
  assign n58124 = ~n3266 & ~n58123;
  assign n58125 = ~n34014 & ~n58124;
  assign inductivity_check  = ~n3263 & n58125;
endmodule


