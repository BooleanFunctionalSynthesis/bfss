// Benchmark "amba2c7y_cert" written by ABC on Sat Jul 29 15:45:24 2017

module amba2c7y_cert ( 
    n33, next_env_fair_out, reg_stateG3_0_out, reg_controllable_locked_out,
    reg_stateG3_1_out, reg_controllable_ndecide_out, reg_stateG3_2_out,
    reg_i_hbusreq0_out, reg_controllable_busreq_out,
    reg_controllable_nstart_out, reg_i_hbusreq1_out, reg_stateG2_out,
    reg_stateG10_1_out, reg_controllable_nhgrant0_out, reg_stateA1_out,
    reg_controllable_hmastlock_out, next_sys_fair<0>_out ,
    next_sys_fair<1>_out , next_sys_fair<2>_out , reg_i_hlock1_out,
    fair_cnt<0>_out , fair_cnt<1>_out , fair_cnt<2>_out ,
    env_safe_err_happened_out, reg_i_hlock0_out, reg_i_hready_out,
    reg_controllable_hgrant1_out, reg_controllable_hmaster0_out,
    i_hbusreq0, i_hbusreq1, i_hburst1, i_hburst0, i_hlock0, i_hlock1,
    i_hready, controllable_hmastlock, controllable_nstart,
    controllable_locked, controllable_hmaster0, controllable_hgrant1,
    controllable_busreq, controllable_ndecide, controllable_nhgrant0,
    inductivity_check   );
  input  n33, next_env_fair_out, reg_stateG3_0_out,
    reg_controllable_locked_out, reg_stateG3_1_out,
    reg_controllable_ndecide_out, reg_stateG3_2_out, reg_i_hbusreq0_out,
    reg_controllable_busreq_out, reg_controllable_nstart_out,
    reg_i_hbusreq1_out, reg_stateG2_out, reg_stateG10_1_out,
    reg_controllable_nhgrant0_out, reg_stateA1_out,
    reg_controllable_hmastlock_out, next_sys_fair<0>_out ,
    next_sys_fair<1>_out , next_sys_fair<2>_out , reg_i_hlock1_out,
    fair_cnt<0>_out , fair_cnt<1>_out , fair_cnt<2>_out ,
    env_safe_err_happened_out, reg_i_hlock0_out, reg_i_hready_out,
    reg_controllable_hgrant1_out, reg_controllable_hmaster0_out,
    i_hbusreq0, i_hbusreq1, i_hburst1, i_hburst0, i_hlock0, i_hlock1,
    i_hready, controllable_hmastlock, controllable_nstart,
    controllable_locked, controllable_hmaster0, controllable_hgrant1,
    controllable_busreq, controllable_ndecide, controllable_nhgrant0;
  output inductivity_check ;
  wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
    n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
    n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
    n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335;
  assign n45 = ~reg_stateG3_0_out & reg_stateG3_1_out;
  assign n46 = ~reg_stateG3_0_out & ~n45;
  assign n47 = ~reg_stateG3_2_out & ~n46;
  assign n48 = ~reg_stateG3_2_out & ~n47;
  assign n49 = ~fair_cnt<0>_out  & ~n48;
  assign n50 = ~fair_cnt<0>_out  & ~n49;
  assign n51 = ~fair_cnt<1>_out  & ~n50;
  assign n52 = ~fair_cnt<1>_out  & ~n51;
  assign n53 = ~fair_cnt<2>_out  & ~n52;
  assign n54 = ~fair_cnt<2>_out  & ~n53;
  assign n55 = ~reg_stateA1_out & ~n54;
  assign n56 = ~reg_stateA1_out & ~n55;
  assign n57 = reg_i_hready_out & ~n56;
  assign n58 = reg_i_hready_out & ~n57;
  assign n59 = next_sys_fair<1>_out  & ~n58;
  assign n60 = fair_cnt<1>_out  & ~n50;
  assign n61 = ~fair_cnt<1>_out  & ~n48;
  assign n62 = ~n60 & ~n61;
  assign n63 = fair_cnt<2>_out  & ~n62;
  assign n64 = ~fair_cnt<2>_out  & ~n48;
  assign n65 = ~n63 & ~n64;
  assign n66 = ~reg_stateA1_out & ~n65;
  assign n67 = ~reg_stateA1_out & ~n66;
  assign n68 = reg_i_hready_out & ~n67;
  assign n69 = reg_i_hready_out & ~n68;
  assign n70 = ~next_sys_fair<1>_out  & ~n69;
  assign n71 = ~n59 & ~n70;
  assign n72 = reg_controllable_locked_out & ~n71;
  assign n73 = next_env_fair_out & ~n52;
  assign n74 = ~fair_cnt<1>_out  & ~n61;
  assign n75 = ~next_env_fair_out & ~n74;
  assign n76 = ~n73 & ~n75;
  assign n77 = fair_cnt<2>_out  & ~n76;
  assign n78 = ~n64 & ~n77;
  assign n79 = reg_i_hready_out & ~n78;
  assign n80 = ~fair_cnt<0>_out  & ~n46;
  assign n81 = ~fair_cnt<0>_out  & ~n80;
  assign n82 = fair_cnt<1>_out  & ~n81;
  assign n83 = ~fair_cnt<1>_out  & ~n46;
  assign n84 = ~n82 & ~n83;
  assign n85 = fair_cnt<2>_out  & ~n84;
  assign n86 = ~fair_cnt<2>_out  & ~n46;
  assign n87 = ~n85 & ~n86;
  assign n88 = ~reg_i_hready_out & ~n87;
  assign n89 = ~n79 & ~n88;
  assign n90 = next_sys_fair<1>_out  & ~n89;
  assign n91 = reg_i_hready_out & ~n65;
  assign n92 = ~n60 & ~n83;
  assign n93 = fair_cnt<2>_out  & ~n92;
  assign n94 = ~n86 & ~n93;
  assign n95 = ~reg_i_hready_out & ~n94;
  assign n96 = ~n91 & ~n95;
  assign n97 = ~next_sys_fair<1>_out  & ~n96;
  assign n98 = ~n90 & ~n97;
  assign n99 = ~reg_controllable_locked_out & ~n98;
  assign n100 = ~n72 & ~n99;
  assign n101 = next_sys_fair<0>_out  & ~n100;
  assign n102 = reg_controllable_locked_out & ~n69;
  assign n103 = ~fair_cnt<1>_out  & ~n83;
  assign n104 = fair_cnt<2>_out  & ~n103;
  assign n105 = ~n86 & ~n104;
  assign n106 = ~reg_i_hready_out & ~n105;
  assign n107 = ~n91 & ~n106;
  assign n108 = next_sys_fair<1>_out  & ~n107;
  assign n109 = ~n88 & ~n91;
  assign n110 = ~next_sys_fair<1>_out  & ~n109;
  assign n111 = ~n108 & ~n110;
  assign n112 = ~reg_controllable_locked_out & ~n111;
  assign n113 = ~n102 & ~n112;
  assign n114 = ~next_sys_fair<0>_out  & ~n113;
  assign n115 = ~n101 & ~n114;
  assign n116 = ~reg_controllable_nhgrant0_out & ~n115;
  assign n117 = ~reg_controllable_nhgrant0_out & ~n116;
  assign n118 = ~reg_controllable_hgrant1_out & ~n117;
  assign n119 = ~reg_controllable_hgrant1_out & ~n118;
  assign n120 = reg_controllable_hmastlock_out & ~n119;
  assign n121 = ~reg_stateA1_out & ~n87;
  assign n122 = ~reg_stateA1_out & ~n121;
  assign n123 = ~reg_i_hready_out & ~n122;
  assign n124 = ~n57 & ~n123;
  assign n125 = next_sys_fair<1>_out  & ~n124;
  assign n126 = ~reg_stateA1_out & ~n94;
  assign n127 = ~reg_stateA1_out & ~n126;
  assign n128 = ~reg_i_hready_out & ~n127;
  assign n129 = ~n68 & ~n128;
  assign n130 = ~next_sys_fair<1>_out  & ~n129;
  assign n131 = ~n125 & ~n130;
  assign n132 = reg_controllable_locked_out & ~n131;
  assign n133 = ~n99 & ~n132;
  assign n134 = next_sys_fair<0>_out  & ~n133;
  assign n135 = ~reg_stateA1_out & ~n105;
  assign n136 = ~reg_stateA1_out & ~n135;
  assign n137 = ~reg_i_hready_out & ~n136;
  assign n138 = ~n68 & ~n137;
  assign n139 = next_sys_fair<1>_out  & ~n138;
  assign n140 = ~n68 & ~n123;
  assign n141 = ~next_sys_fair<1>_out  & ~n140;
  assign n142 = ~n139 & ~n141;
  assign n143 = reg_controllable_locked_out & ~n142;
  assign n144 = ~n112 & ~n143;
  assign n145 = ~next_sys_fair<0>_out  & ~n144;
  assign n146 = ~n134 & ~n145;
  assign n147 = ~reg_controllable_nhgrant0_out & ~n146;
  assign n148 = ~reg_controllable_nhgrant0_out & ~n147;
  assign n149 = ~reg_controllable_hgrant1_out & ~n148;
  assign n150 = ~reg_controllable_hgrant1_out & ~n149;
  assign n151 = ~reg_controllable_hmastlock_out & ~n150;
  assign n152 = ~n120 & ~n151;
  assign n153 = ~reg_stateG2_out & ~n152;
  assign n154 = ~reg_stateG2_out & ~n153;
  assign n155 = reg_controllable_hmaster0_out & ~n154;
  assign n156 = ~fair_cnt<1>_out  & ~n81;
  assign n157 = ~fair_cnt<1>_out  & ~n156;
  assign n158 = ~next_env_fair_out & ~n157;
  assign n159 = ~next_env_fair_out & ~n158;
  assign n160 = fair_cnt<2>_out  & ~n159;
  assign n161 = fair_cnt<0>_out  & ~n46;
  assign n162 = reg_stateG3_2_out & ~n46;
  assign n163 = reg_stateG3_0_out & reg_stateG3_1_out;
  assign n164 = ~reg_stateG3_0_out & ~reg_stateG3_1_out;
  assign n165 = ~n163 & ~n164;
  assign n166 = ~reg_stateG3_2_out & n165;
  assign n167 = ~n162 & ~n166;
  assign n168 = ~fair_cnt<0>_out  & ~n167;
  assign n169 = ~n161 & ~n168;
  assign n170 = fair_cnt<1>_out  & ~n169;
  assign n171 = reg_stateG3_0_out & ~n163;
  assign n172 = ~reg_stateG3_2_out & n171;
  assign n173 = ~n162 & ~n172;
  assign n174 = fair_cnt<0>_out  & ~n173;
  assign n175 = ~fair_cnt<0>_out  & n162;
  assign n176 = ~n174 & ~n175;
  assign n177 = ~fair_cnt<1>_out  & ~n176;
  assign n178 = ~n170 & ~n177;
  assign n179 = ~fair_cnt<2>_out  & ~n178;
  assign n180 = ~n160 & ~n179;
  assign n181 = reg_stateA1_out & ~n180;
  assign n182 = reg_stateA1_out & ~n181;
  assign n183 = next_sys_fair<1>_out  & ~n182;
  assign n184 = ~fair_cnt<1>_out  & ~n169;
  assign n185 = ~n60 & ~n184;
  assign n186 = fair_cnt<2>_out  & ~n185;
  assign n187 = fair_cnt<1>_out  & ~n176;
  assign n188 = ~fair_cnt<1>_out  & n162;
  assign n189 = ~n187 & ~n188;
  assign n190 = ~fair_cnt<2>_out  & ~n189;
  assign n191 = ~n186 & ~n190;
  assign n192 = reg_stateA1_out & ~n191;
  assign n193 = reg_stateA1_out & ~n192;
  assign n194 = ~next_sys_fair<1>_out  & ~n193;
  assign n195 = ~n183 & ~n194;
  assign n196 = reg_controllable_locked_out & ~n195;
  assign n197 = reg_controllable_locked_out & ~n196;
  assign n198 = next_sys_fair<0>_out  & ~n197;
  assign n199 = ~fair_cnt<0>_out  & ~n175;
  assign n200 = fair_cnt<1>_out  & ~n199;
  assign n201 = ~n188 & ~n200;
  assign n202 = fair_cnt<2>_out  & ~n201;
  assign n203 = ~fair_cnt<2>_out  & n162;
  assign n204 = ~n202 & ~n203;
  assign n205 = reg_stateA1_out & ~n204;
  assign n206 = reg_stateA1_out & ~n205;
  assign n207 = next_sys_fair<1>_out  & ~n206;
  assign n208 = ~fair_cnt<1>_out  & ~n188;
  assign n209 = next_env_fair_out & ~n208;
  assign n210 = ~next_env_fair_out & ~n201;
  assign n211 = ~n209 & ~n210;
  assign n212 = fair_cnt<2>_out  & ~n211;
  assign n213 = ~n203 & ~n212;
  assign n214 = reg_stateA1_out & ~n213;
  assign n215 = reg_stateA1_out & ~n214;
  assign n216 = ~next_sys_fair<1>_out  & ~n215;
  assign n217 = ~n207 & ~n216;
  assign n218 = reg_controllable_locked_out & ~n217;
  assign n219 = reg_controllable_locked_out & ~n218;
  assign n220 = ~next_sys_fair<0>_out  & ~n219;
  assign n221 = ~n198 & ~n220;
  assign n222 = ~reg_controllable_nhgrant0_out & ~n221;
  assign n223 = ~reg_controllable_nhgrant0_out & ~n222;
  assign n224 = ~reg_controllable_hgrant1_out & ~n223;
  assign n225 = ~reg_controllable_hgrant1_out & ~n224;
  assign n226 = reg_controllable_hmastlock_out & ~n225;
  assign n227 = ~fair_cnt<0>_out  & ~n168;
  assign n228 = ~fair_cnt<1>_out  & ~n227;
  assign n229 = ~fair_cnt<1>_out  & ~n228;
  assign n230 = next_env_fair_out & ~n229;
  assign n231 = ~fair_cnt<1>_out  & ~n184;
  assign n232 = ~next_env_fair_out & ~n231;
  assign n233 = ~n230 & ~n232;
  assign n234 = fair_cnt<2>_out  & ~n233;
  assign n235 = ~n190 & ~n234;
  assign n236 = reg_stateA1_out & ~n235;
  assign n237 = reg_stateA1_out & ~n236;
  assign n238 = next_sys_fair<1>_out  & ~n237;
  assign n239 = ~n194 & ~n238;
  assign n240 = ~reg_controllable_locked_out & ~n239;
  assign n241 = ~reg_controllable_locked_out & ~n240;
  assign n242 = next_sys_fair<0>_out  & ~n241;
  assign n243 = ~reg_controllable_locked_out & ~n217;
  assign n244 = ~reg_controllable_locked_out & ~n243;
  assign n245 = ~next_sys_fair<0>_out  & ~n244;
  assign n246 = ~n242 & ~n245;
  assign n247 = ~reg_controllable_nhgrant0_out & ~n246;
  assign n248 = ~reg_controllable_nhgrant0_out & ~n247;
  assign n249 = ~reg_controllable_hgrant1_out & ~n248;
  assign n250 = ~reg_controllable_hgrant1_out & ~n249;
  assign n251 = ~reg_controllable_hmastlock_out & ~n250;
  assign n252 = ~n226 & ~n251;
  assign n253 = reg_stateG2_out & ~n252;
  assign n254 = fair_cnt<1>_out  & ~n227;
  assign n255 = ~n177 & ~n254;
  assign n256 = next_env_fair_out & ~n255;
  assign n257 = ~next_env_fair_out & ~n178;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~fair_cnt<2>_out  & ~n258;
  assign n260 = ~fair_cnt<2>_out  & ~n259;
  assign n261 = ~reg_stateA1_out & ~n260;
  assign n262 = ~n181 & ~n261;
  assign n263 = next_sys_fair<1>_out  & ~n262;
  assign n264 = ~next_sys_fair<1>_out  & ~n191;
  assign n265 = ~n263 & ~n264;
  assign n266 = reg_controllable_locked_out & ~n265;
  assign n267 = fair_cnt<2>_out  & ~n157;
  assign n268 = ~n86 & ~n267;
  assign n269 = ~reg_i_hready_out & ~n268;
  assign n270 = ~n79 & ~n269;
  assign n271 = next_sys_fair<1>_out  & ~n270;
  assign n272 = ~n97 & ~n271;
  assign n273 = ~reg_controllable_locked_out & ~n272;
  assign n274 = ~n266 & ~n273;
  assign n275 = next_sys_fair<0>_out  & ~n274;
  assign n276 = reg_controllable_locked_out & ~n204;
  assign n277 = ~reg_controllable_locked_out & ~n109;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~next_sys_fair<0>_out  & ~n278;
  assign n280 = ~n275 & ~n279;
  assign n281 = ~reg_controllable_nhgrant0_out & ~n280;
  assign n282 = ~reg_controllable_nhgrant0_out & ~n281;
  assign n283 = ~reg_controllable_hgrant1_out & ~n282;
  assign n284 = ~reg_controllable_hgrant1_out & ~n283;
  assign n285 = reg_controllable_hmastlock_out & ~n284;
  assign n286 = ~fair_cnt<2>_out  & ~n159;
  assign n287 = ~fair_cnt<2>_out  & ~n286;
  assign n288 = ~reg_stateA1_out & ~n287;
  assign n289 = ~reg_stateA1_out & ~n288;
  assign n290 = ~reg_i_hready_out & ~n289;
  assign n291 = ~n57 & ~n290;
  assign n292 = next_sys_fair<1>_out  & ~n291;
  assign n293 = ~n130 & ~n292;
  assign n294 = reg_controllable_locked_out & ~n293;
  assign n295 = next_sys_fair<1>_out  & ~n235;
  assign n296 = ~n264 & ~n295;
  assign n297 = ~reg_controllable_locked_out & ~n296;
  assign n298 = ~n294 & ~n297;
  assign n299 = next_sys_fair<0>_out  & ~n298;
  assign n300 = reg_controllable_locked_out & ~n140;
  assign n301 = ~reg_controllable_locked_out & ~n204;
  assign n302 = ~n300 & ~n301;
  assign n303 = ~next_sys_fair<0>_out  & ~n302;
  assign n304 = ~n299 & ~n303;
  assign n305 = ~reg_controllable_nhgrant0_out & ~n304;
  assign n306 = ~reg_controllable_nhgrant0_out & ~n305;
  assign n307 = ~reg_controllable_hgrant1_out & ~n306;
  assign n308 = ~reg_controllable_hgrant1_out & ~n307;
  assign n309 = ~reg_controllable_hmastlock_out & ~n308;
  assign n310 = ~n285 & ~n309;
  assign n311 = ~reg_stateG2_out & ~n310;
  assign n312 = ~n253 & ~n311;
  assign n313 = ~reg_controllable_hmaster0_out & ~n312;
  assign n314 = ~n155 & ~n313;
  assign n315 = reg_controllable_ndecide_out & ~n314;
  assign n316 = reg_stateA1_out & ~n87;
  assign n317 = reg_stateA1_out & ~n316;
  assign n318 = next_sys_fair<1>_out  & ~n317;
  assign n319 = reg_stateA1_out & ~n94;
  assign n320 = reg_stateA1_out & ~n319;
  assign n321 = ~next_sys_fair<1>_out  & ~n320;
  assign n322 = ~n318 & ~n321;
  assign n323 = reg_controllable_locked_out & ~n322;
  assign n324 = ~reg_i_hready_out & ~n317;
  assign n325 = ~reg_i_hready_out & ~n324;
  assign n326 = next_sys_fair<1>_out  & ~n325;
  assign n327 = ~reg_i_hready_out & ~n320;
  assign n328 = ~reg_i_hready_out & ~n327;
  assign n329 = ~next_sys_fair<1>_out  & ~n328;
  assign n330 = ~n326 & ~n329;
  assign n331 = ~reg_controllable_locked_out & ~n330;
  assign n332 = ~n323 & ~n331;
  assign n333 = next_sys_fair<0>_out  & ~n332;
  assign n334 = ~n86 & ~n160;
  assign n335 = reg_stateA1_out & ~n334;
  assign n336 = reg_stateA1_out & ~n335;
  assign n337 = next_sys_fair<1>_out  & ~n336;
  assign n338 = next_env_fair_out & ~n103;
  assign n339 = ~next_env_fair_out & ~n84;
  assign n340 = ~n338 & ~n339;
  assign n341 = fair_cnt<2>_out  & ~n340;
  assign n342 = ~n86 & ~n341;
  assign n343 = reg_stateA1_out & ~n342;
  assign n344 = reg_stateA1_out & ~n343;
  assign n345 = ~next_sys_fair<1>_out  & ~n344;
  assign n346 = ~n337 & ~n345;
  assign n347 = reg_controllable_locked_out & ~n346;
  assign n348 = ~reg_i_hready_out & ~n336;
  assign n349 = ~reg_i_hready_out & ~n348;
  assign n350 = next_sys_fair<1>_out  & ~n349;
  assign n351 = ~reg_i_hready_out & ~n344;
  assign n352 = ~reg_i_hready_out & ~n351;
  assign n353 = ~next_sys_fair<1>_out  & ~n352;
  assign n354 = ~n350 & ~n353;
  assign n355 = ~reg_controllable_locked_out & ~n354;
  assign n356 = ~n347 & ~n355;
  assign n357 = ~next_sys_fair<0>_out  & ~n356;
  assign n358 = ~n333 & ~n357;
  assign n359 = reg_i_hbusreq0_out & ~n358;
  assign n360 = reg_i_hbusreq1_out & ~n358;
  assign n361 = reg_i_hbusreq1_out & ~n360;
  assign n362 = ~reg_i_hbusreq0_out & ~n361;
  assign n363 = ~n359 & ~n362;
  assign n364 = reg_controllable_nhgrant0_out & ~n363;
  assign n365 = next_sys_fair<0>_out  & ~n330;
  assign n366 = ~next_sys_fair<0>_out  & ~n354;
  assign n367 = ~n365 & ~n366;
  assign n368 = reg_i_hbusreq0_out & ~n367;
  assign n369 = reg_i_hbusreq1_out & ~n367;
  assign n370 = reg_i_hbusreq1_out & ~n369;
  assign n371 = ~reg_i_hbusreq0_out & ~n370;
  assign n372 = ~n368 & ~n371;
  assign n373 = ~reg_controllable_nhgrant0_out & ~n372;
  assign n374 = ~n364 & ~n373;
  assign n375 = reg_controllable_hgrant1_out & ~n374;
  assign n376 = ~reg_controllable_hgrant1_out & ~n372;
  assign n377 = ~n375 & ~n376;
  assign n378 = reg_controllable_hmastlock_out & ~n377;
  assign n379 = reg_controllable_hmastlock_out & ~n378;
  assign n380 = ~reg_i_hlock0_out & ~n379;
  assign n381 = ~reg_i_hlock0_out & ~n380;
  assign n382 = reg_stateG2_out & ~n381;
  assign n383 = ~reg_controllable_locked_out & ~n69;
  assign n384 = ~reg_controllable_locked_out & ~n383;
  assign n385 = next_sys_fair<0>_out  & ~n384;
  assign n386 = fair_cnt<2>_out  & ~n74;
  assign n387 = ~n64 & ~n386;
  assign n388 = ~reg_stateA1_out & ~n387;
  assign n389 = ~reg_stateA1_out & ~n388;
  assign n390 = reg_i_hready_out & ~n389;
  assign n391 = reg_i_hready_out & ~n390;
  assign n392 = next_sys_fair<1>_out  & ~n391;
  assign n393 = ~n70 & ~n392;
  assign n394 = ~reg_controllable_locked_out & ~n393;
  assign n395 = ~reg_controllable_locked_out & ~n394;
  assign n396 = ~next_sys_fair<0>_out  & ~n395;
  assign n397 = ~n385 & ~n396;
  assign n398 = reg_controllable_nhgrant0_out & ~n397;
  assign n399 = reg_controllable_nhgrant0_out & ~n398;
  assign n400 = reg_controllable_hgrant1_out & ~n399;
  assign n401 = ~n72 & ~n394;
  assign n402 = next_sys_fair<0>_out  & ~n401;
  assign n403 = ~next_sys_fair<0>_out  & ~n69;
  assign n404 = ~n402 & ~n403;
  assign n405 = reg_i_hbusreq0_out & ~n404;
  assign n406 = reg_i_hbusreq1_out & ~n404;
  assign n407 = ~next_env_fair_out & ~n52;
  assign n408 = ~next_env_fair_out & ~n407;
  assign n409 = ~fair_cnt<2>_out  & ~n408;
  assign n410 = ~fair_cnt<2>_out  & ~n409;
  assign n411 = ~reg_stateA1_out & ~n410;
  assign n412 = ~reg_stateA1_out & ~n411;
  assign n413 = reg_i_hready_out & ~n412;
  assign n414 = reg_i_hready_out & ~n413;
  assign n415 = next_sys_fair<1>_out  & ~n414;
  assign n416 = ~n70 & ~n415;
  assign n417 = ~reg_controllable_locked_out & ~n416;
  assign n418 = ~n72 & ~n417;
  assign n419 = next_sys_fair<0>_out  & ~n418;
  assign n420 = ~n403 & ~n419;
  assign n421 = ~reg_i_hbusreq1_out & ~n420;
  assign n422 = ~n406 & ~n421;
  assign n423 = ~reg_i_hbusreq0_out & ~n422;
  assign n424 = ~n405 & ~n423;
  assign n425 = ~reg_controllable_nhgrant0_out & ~n424;
  assign n426 = ~reg_controllable_nhgrant0_out & ~n425;
  assign n427 = ~reg_controllable_hgrant1_out & ~n426;
  assign n428 = ~n400 & ~n427;
  assign n429 = reg_controllable_hmastlock_out & ~n428;
  assign n430 = ~reg_i_hready_out & ~n123;
  assign n431 = next_sys_fair<1>_out  & ~n430;
  assign n432 = ~reg_i_hready_out & ~n128;
  assign n433 = ~next_sys_fair<1>_out  & ~n432;
  assign n434 = ~n431 & ~n433;
  assign n435 = reg_controllable_locked_out & ~n434;
  assign n436 = next_sys_fair<1>_out  & ~n122;
  assign n437 = ~next_sys_fair<1>_out  & ~n127;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~reg_controllable_locked_out & ~n438;
  assign n440 = ~n435 & ~n439;
  assign n441 = next_sys_fair<0>_out  & ~n440;
  assign n442 = ~reg_i_hready_out & ~n137;
  assign n443 = next_sys_fair<1>_out  & ~n442;
  assign n444 = ~next_sys_fair<1>_out  & ~n430;
  assign n445 = ~n443 & ~n444;
  assign n446 = reg_controllable_locked_out & ~n445;
  assign n447 = next_sys_fair<1>_out  & ~n136;
  assign n448 = ~next_sys_fair<1>_out  & ~n122;
  assign n449 = ~n447 & ~n448;
  assign n450 = ~reg_controllable_locked_out & ~n449;
  assign n451 = ~n446 & ~n450;
  assign n452 = ~next_sys_fair<0>_out  & ~n451;
  assign n453 = ~n441 & ~n452;
  assign n454 = reg_controllable_nhgrant0_out & ~n453;
  assign n455 = next_sys_fair<0>_out  & ~n434;
  assign n456 = ~next_sys_fair<0>_out  & ~n445;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~reg_controllable_nhgrant0_out & ~n457;
  assign n459 = ~n454 & ~n458;
  assign n460 = reg_controllable_hgrant1_out & ~n459;
  assign n461 = reg_controllable_nhgrant0_out & ~n457;
  assign n462 = ~n123 & ~n390;
  assign n463 = next_sys_fair<1>_out  & ~n462;
  assign n464 = ~n130 & ~n463;
  assign n465 = ~reg_controllable_locked_out & ~n464;
  assign n466 = ~n132 & ~n465;
  assign n467 = next_sys_fair<0>_out  & ~n466;
  assign n468 = ~next_sys_fair<0>_out  & ~n142;
  assign n469 = ~n467 & ~n468;
  assign n470 = reg_i_hbusreq0_out & ~n469;
  assign n471 = reg_i_hbusreq1_out & ~n469;
  assign n472 = ~n123 & ~n413;
  assign n473 = next_sys_fair<1>_out  & ~n472;
  assign n474 = ~n130 & ~n473;
  assign n475 = ~reg_controllable_locked_out & ~n474;
  assign n476 = ~n132 & ~n475;
  assign n477 = next_sys_fair<0>_out  & ~n476;
  assign n478 = ~n468 & ~n477;
  assign n479 = ~reg_i_hbusreq1_out & ~n478;
  assign n480 = ~n471 & ~n479;
  assign n481 = ~reg_i_hbusreq0_out & ~n480;
  assign n482 = ~n470 & ~n481;
  assign n483 = ~reg_controllable_nhgrant0_out & ~n482;
  assign n484 = ~n461 & ~n483;
  assign n485 = ~reg_controllable_hgrant1_out & ~n484;
  assign n486 = ~n460 & ~n485;
  assign n487 = ~reg_controllable_hmastlock_out & ~n486;
  assign n488 = ~n429 & ~n487;
  assign n489 = reg_i_hlock0_out & ~n488;
  assign n490 = next_sys_fair<1>_out  & ~n87;
  assign n491 = ~next_sys_fair<1>_out  & ~n94;
  assign n492 = ~n490 & ~n491;
  assign n493 = reg_controllable_locked_out & ~n492;
  assign n494 = next_sys_fair<1>_out  & ~n109;
  assign n495 = ~n97 & ~n494;
  assign n496 = ~reg_controllable_locked_out & ~n495;
  assign n497 = ~n493 & ~n496;
  assign n498 = next_sys_fair<0>_out  & ~n497;
  assign n499 = next_sys_fair<1>_out  & ~n105;
  assign n500 = ~next_sys_fair<1>_out  & ~n87;
  assign n501 = ~n499 & ~n500;
  assign n502 = reg_controllable_locked_out & ~n501;
  assign n503 = reg_i_hready_out & ~n387;
  assign n504 = ~n106 & ~n503;
  assign n505 = next_sys_fair<1>_out  & ~n504;
  assign n506 = ~n110 & ~n505;
  assign n507 = ~reg_controllable_locked_out & ~n506;
  assign n508 = ~n502 & ~n507;
  assign n509 = ~next_sys_fair<0>_out  & ~n508;
  assign n510 = ~n498 & ~n509;
  assign n511 = reg_controllable_nhgrant0_out & ~n510;
  assign n512 = ~reg_i_hready_out & ~n88;
  assign n513 = next_sys_fair<1>_out  & ~n512;
  assign n514 = ~reg_i_hready_out & ~n95;
  assign n515 = ~next_sys_fair<1>_out  & ~n514;
  assign n516 = ~n513 & ~n515;
  assign n517 = next_sys_fair<0>_out  & ~n516;
  assign n518 = ~reg_i_hready_out & ~n106;
  assign n519 = next_sys_fair<1>_out  & ~n518;
  assign n520 = ~next_sys_fair<1>_out  & ~n512;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~next_sys_fair<0>_out  & ~n521;
  assign n523 = ~n517 & ~n522;
  assign n524 = ~reg_controllable_nhgrant0_out & ~n523;
  assign n525 = ~n511 & ~n524;
  assign n526 = reg_controllable_hgrant1_out & ~n525;
  assign n527 = reg_controllable_nhgrant0_out & ~n523;
  assign n528 = reg_controllable_locked_out & ~n516;
  assign n529 = reg_stateA1_out & ~n78;
  assign n530 = ~n388 & ~n529;
  assign n531 = reg_i_hready_out & ~n530;
  assign n532 = ~n88 & ~n531;
  assign n533 = next_sys_fair<1>_out  & ~n532;
  assign n534 = ~n97 & ~n533;
  assign n535 = ~reg_controllable_locked_out & ~n534;
  assign n536 = ~n528 & ~n535;
  assign n537 = next_sys_fair<0>_out  & ~n536;
  assign n538 = reg_controllable_locked_out & ~n521;
  assign n539 = ~n112 & ~n538;
  assign n540 = ~next_sys_fair<0>_out  & ~n539;
  assign n541 = ~n537 & ~n540;
  assign n542 = reg_i_hbusreq0_out & ~n541;
  assign n543 = reg_i_hbusreq1_out & ~n541;
  assign n544 = ~n99 & ~n528;
  assign n545 = next_sys_fair<0>_out  & ~n544;
  assign n546 = ~n540 & ~n545;
  assign n547 = ~reg_i_hbusreq1_out & ~n546;
  assign n548 = ~n543 & ~n547;
  assign n549 = ~reg_i_hbusreq0_out & ~n548;
  assign n550 = ~n542 & ~n549;
  assign n551 = ~reg_controllable_nhgrant0_out & ~n550;
  assign n552 = ~n527 & ~n551;
  assign n553 = ~reg_controllable_hgrant1_out & ~n552;
  assign n554 = ~n526 & ~n553;
  assign n555 = reg_controllable_hmastlock_out & ~n554;
  assign n556 = ~reg_controllable_locked_out & ~n492;
  assign n557 = ~n528 & ~n556;
  assign n558 = next_sys_fair<0>_out  & ~n557;
  assign n559 = ~reg_controllable_locked_out & ~n501;
  assign n560 = ~n538 & ~n559;
  assign n561 = ~next_sys_fair<0>_out  & ~n560;
  assign n562 = ~n558 & ~n561;
  assign n563 = reg_controllable_nhgrant0_out & ~n562;
  assign n564 = ~n524 & ~n563;
  assign n565 = reg_controllable_hgrant1_out & ~n564;
  assign n566 = ~n553 & ~n565;
  assign n567 = ~reg_controllable_hmastlock_out & ~n566;
  assign n568 = ~n555 & ~n567;
  assign n569 = ~reg_i_hlock0_out & ~n568;
  assign n570 = ~n489 & ~n569;
  assign n571 = ~reg_stateG2_out & ~n570;
  assign n572 = ~n382 & ~n571;
  assign n573 = reg_controllable_hmaster0_out & ~n572;
  assign n574 = ~reg_i_hready_out & ~n182;
  assign n575 = ~reg_i_hready_out & ~n574;
  assign n576 = next_sys_fair<1>_out  & ~n575;
  assign n577 = ~reg_i_hready_out & ~n193;
  assign n578 = ~reg_i_hready_out & ~n577;
  assign n579 = ~next_sys_fair<1>_out  & ~n578;
  assign n580 = ~n576 & ~n579;
  assign n581 = next_sys_fair<0>_out  & ~n580;
  assign n582 = ~reg_i_hready_out & ~n206;
  assign n583 = ~reg_i_hready_out & ~n582;
  assign n584 = next_sys_fair<1>_out  & ~n583;
  assign n585 = ~reg_i_hready_out & ~n215;
  assign n586 = ~reg_i_hready_out & ~n585;
  assign n587 = ~next_sys_fair<1>_out  & ~n586;
  assign n588 = ~n584 & ~n587;
  assign n589 = ~next_sys_fair<0>_out  & ~n588;
  assign n590 = ~n581 & ~n589;
  assign n591 = reg_controllable_hgrant1_out & ~n590;
  assign n592 = reg_controllable_nhgrant0_out & ~n590;
  assign n593 = ~reg_controllable_locked_out & ~n580;
  assign n594 = ~n196 & ~n593;
  assign n595 = next_sys_fair<0>_out  & ~n594;
  assign n596 = ~reg_controllable_locked_out & ~n588;
  assign n597 = ~n218 & ~n596;
  assign n598 = ~next_sys_fair<0>_out  & ~n597;
  assign n599 = ~n595 & ~n598;
  assign n600 = ~reg_controllable_nhgrant0_out & ~n599;
  assign n601 = ~n592 & ~n600;
  assign n602 = ~reg_controllable_hgrant1_out & ~n601;
  assign n603 = ~n591 & ~n602;
  assign n604 = reg_controllable_hmastlock_out & ~n603;
  assign n605 = reg_controllable_hmastlock_out & ~n604;
  assign n606 = reg_i_hlock0_out & ~n605;
  assign n607 = ~reg_i_hready_out & ~n237;
  assign n608 = ~reg_i_hready_out & ~n607;
  assign n609 = next_sys_fair<1>_out  & ~n608;
  assign n610 = ~n579 & ~n609;
  assign n611 = next_sys_fair<0>_out  & ~n610;
  assign n612 = ~n589 & ~n611;
  assign n613 = reg_controllable_hgrant1_out & ~n612;
  assign n614 = reg_controllable_nhgrant0_out & ~n612;
  assign n615 = reg_controllable_locked_out & ~n610;
  assign n616 = ~n240 & ~n615;
  assign n617 = next_sys_fair<0>_out  & ~n616;
  assign n618 = reg_controllable_locked_out & ~n588;
  assign n619 = ~n243 & ~n618;
  assign n620 = ~next_sys_fair<0>_out  & ~n619;
  assign n621 = ~n617 & ~n620;
  assign n622 = ~reg_controllable_nhgrant0_out & ~n621;
  assign n623 = ~n614 & ~n622;
  assign n624 = ~reg_controllable_hgrant1_out & ~n623;
  assign n625 = ~n613 & ~n624;
  assign n626 = ~reg_controllable_hmastlock_out & ~n625;
  assign n627 = ~reg_controllable_hmastlock_out & ~n626;
  assign n628 = ~reg_i_hlock0_out & ~n627;
  assign n629 = ~n606 & ~n628;
  assign n630 = reg_stateG2_out & ~n629;
  assign n631 = ~fair_cnt<2>_out  & ~n179;
  assign n632 = ~reg_stateA1_out & ~n631;
  assign n633 = ~n181 & ~n632;
  assign n634 = ~reg_i_hready_out & ~n633;
  assign n635 = ~reg_i_hready_out & ~n634;
  assign n636 = next_sys_fair<1>_out  & ~n635;
  assign n637 = ~reg_i_hready_out & ~n191;
  assign n638 = ~reg_i_hready_out & ~n637;
  assign n639 = ~next_sys_fair<1>_out  & ~n638;
  assign n640 = ~n636 & ~n639;
  assign n641 = reg_controllable_locked_out & ~n640;
  assign n642 = ~n68 & ~n634;
  assign n643 = next_sys_fair<1>_out  & ~n642;
  assign n644 = ~n68 & ~n637;
  assign n645 = ~next_sys_fair<1>_out  & ~n644;
  assign n646 = ~n643 & ~n645;
  assign n647 = ~reg_controllable_locked_out & ~n646;
  assign n648 = ~n641 & ~n647;
  assign n649 = next_sys_fair<0>_out  & ~n648;
  assign n650 = ~reg_i_hready_out & ~n204;
  assign n651 = ~reg_i_hready_out & ~n650;
  assign n652 = reg_controllable_locked_out & ~n651;
  assign n653 = ~n390 & ~n650;
  assign n654 = next_sys_fair<1>_out  & ~n653;
  assign n655 = ~n68 & ~n650;
  assign n656 = ~next_sys_fair<1>_out  & ~n655;
  assign n657 = ~n654 & ~n656;
  assign n658 = ~reg_controllable_locked_out & ~n657;
  assign n659 = ~n652 & ~n658;
  assign n660 = ~next_sys_fair<0>_out  & ~n659;
  assign n661 = ~n649 & ~n660;
  assign n662 = reg_i_hbusreq0_out & ~n661;
  assign n663 = reg_i_hbusreq1_out & ~n661;
  assign n664 = ~reg_i_hready_out & ~n262;
  assign n665 = ~reg_i_hready_out & ~n664;
  assign n666 = next_sys_fair<1>_out  & ~n665;
  assign n667 = ~n639 & ~n666;
  assign n668 = reg_controllable_locked_out & ~n667;
  assign n669 = ~n68 & ~n664;
  assign n670 = next_sys_fair<1>_out  & ~n669;
  assign n671 = ~n645 & ~n670;
  assign n672 = ~reg_controllable_locked_out & ~n671;
  assign n673 = ~n668 & ~n672;
  assign n674 = next_sys_fair<0>_out  & ~n673;
  assign n675 = ~n660 & ~n674;
  assign n676 = ~reg_i_hbusreq1_out & ~n675;
  assign n677 = ~n663 & ~n676;
  assign n678 = ~reg_i_hbusreq0_out & ~n677;
  assign n679 = ~n662 & ~n678;
  assign n680 = reg_controllable_nhgrant0_out & ~n679;
  assign n681 = next_sys_fair<0>_out  & ~n640;
  assign n682 = ~next_sys_fair<0>_out  & ~n651;
  assign n683 = ~n681 & ~n682;
  assign n684 = reg_i_hbusreq0_out & ~n683;
  assign n685 = reg_i_hbusreq1_out & ~n683;
  assign n686 = next_sys_fair<0>_out  & ~n667;
  assign n687 = ~n682 & ~n686;
  assign n688 = ~reg_i_hbusreq1_out & ~n687;
  assign n689 = ~n685 & ~n688;
  assign n690 = ~reg_i_hbusreq0_out & ~n689;
  assign n691 = ~n684 & ~n690;
  assign n692 = ~reg_controllable_nhgrant0_out & ~n691;
  assign n693 = ~n680 & ~n692;
  assign n694 = reg_controllable_hgrant1_out & ~n693;
  assign n695 = reg_controllable_nhgrant0_out & ~n691;
  assign n696 = next_sys_fair<1>_out  & ~n633;
  assign n697 = ~n264 & ~n696;
  assign n698 = reg_controllable_locked_out & ~n697;
  assign n699 = ~n390 & ~n634;
  assign n700 = next_sys_fair<1>_out  & ~n699;
  assign n701 = ~n645 & ~n700;
  assign n702 = ~reg_controllable_locked_out & ~n701;
  assign n703 = ~n698 & ~n702;
  assign n704 = next_sys_fair<0>_out  & ~n703;
  assign n705 = ~reg_controllable_locked_out & ~n655;
  assign n706 = ~n276 & ~n705;
  assign n707 = ~next_sys_fair<0>_out  & ~n706;
  assign n708 = ~n704 & ~n707;
  assign n709 = reg_i_hbusreq0_out & ~n708;
  assign n710 = reg_i_hbusreq1_out & ~n708;
  assign n711 = ~n413 & ~n664;
  assign n712 = next_sys_fair<1>_out  & ~n711;
  assign n713 = ~n645 & ~n712;
  assign n714 = ~reg_controllable_locked_out & ~n713;
  assign n715 = ~n266 & ~n714;
  assign n716 = next_sys_fair<0>_out  & ~n715;
  assign n717 = ~n707 & ~n716;
  assign n718 = ~reg_i_hbusreq1_out & ~n717;
  assign n719 = ~n710 & ~n718;
  assign n720 = ~reg_i_hbusreq0_out & ~n719;
  assign n721 = ~n709 & ~n720;
  assign n722 = ~reg_controllable_nhgrant0_out & ~n721;
  assign n723 = ~n695 & ~n722;
  assign n724 = ~reg_controllable_hgrant1_out & ~n723;
  assign n725 = ~n694 & ~n724;
  assign n726 = reg_controllable_hmastlock_out & ~n725;
  assign n727 = ~n433 & ~n443;
  assign n728 = reg_controllable_locked_out & ~n727;
  assign n729 = ~n130 & ~n139;
  assign n730 = ~reg_controllable_locked_out & ~n729;
  assign n731 = ~n728 & ~n730;
  assign n732 = next_sys_fair<0>_out  & ~n731;
  assign n733 = reg_controllable_locked_out & ~n430;
  assign n734 = ~n141 & ~n463;
  assign n735 = ~reg_controllable_locked_out & ~n734;
  assign n736 = ~n733 & ~n735;
  assign n737 = ~next_sys_fair<0>_out  & ~n736;
  assign n738 = ~n732 & ~n737;
  assign n739 = reg_i_hbusreq0_out & ~n738;
  assign n740 = reg_i_hbusreq1_out & ~n738;
  assign n741 = ~reg_i_hready_out & ~n290;
  assign n742 = next_sys_fair<1>_out  & ~n741;
  assign n743 = ~n433 & ~n742;
  assign n744 = reg_controllable_locked_out & ~n743;
  assign n745 = ~n68 & ~n290;
  assign n746 = next_sys_fair<1>_out  & ~n745;
  assign n747 = ~n130 & ~n746;
  assign n748 = ~reg_controllable_locked_out & ~n747;
  assign n749 = ~n744 & ~n748;
  assign n750 = next_sys_fair<0>_out  & ~n749;
  assign n751 = ~n737 & ~n750;
  assign n752 = ~reg_i_hbusreq1_out & ~n751;
  assign n753 = ~n740 & ~n752;
  assign n754 = ~reg_i_hbusreq0_out & ~n753;
  assign n755 = ~n739 & ~n754;
  assign n756 = reg_controllable_nhgrant0_out & ~n755;
  assign n757 = next_sys_fair<0>_out  & ~n727;
  assign n758 = ~next_sys_fair<0>_out  & ~n430;
  assign n759 = ~n757 & ~n758;
  assign n760 = reg_i_hbusreq0_out & ~n759;
  assign n761 = reg_i_hbusreq1_out & ~n759;
  assign n762 = next_sys_fair<0>_out  & ~n743;
  assign n763 = ~n758 & ~n762;
  assign n764 = ~reg_i_hbusreq1_out & ~n763;
  assign n765 = ~n761 & ~n764;
  assign n766 = ~reg_i_hbusreq0_out & ~n765;
  assign n767 = ~n760 & ~n766;
  assign n768 = ~reg_controllable_nhgrant0_out & ~n767;
  assign n769 = ~n756 & ~n768;
  assign n770 = reg_controllable_hgrant1_out & ~n769;
  assign n771 = reg_controllable_nhgrant0_out & ~n767;
  assign n772 = ~n57 & ~n137;
  assign n773 = next_sys_fair<1>_out  & ~n772;
  assign n774 = ~n130 & ~n773;
  assign n775 = reg_controllable_locked_out & ~n774;
  assign n776 = ~n437 & ~n447;
  assign n777 = ~reg_controllable_locked_out & ~n776;
  assign n778 = ~n775 & ~n777;
  assign n779 = next_sys_fair<0>_out  & ~n778;
  assign n780 = ~reg_controllable_locked_out & ~n122;
  assign n781 = ~n300 & ~n780;
  assign n782 = ~next_sys_fair<0>_out  & ~n781;
  assign n783 = ~n779 & ~n782;
  assign n784 = reg_i_hbusreq0_out & ~n783;
  assign n785 = reg_i_hbusreq1_out & ~n783;
  assign n786 = next_sys_fair<1>_out  & ~n289;
  assign n787 = ~n437 & ~n786;
  assign n788 = ~reg_controllable_locked_out & ~n787;
  assign n789 = ~n294 & ~n788;
  assign n790 = next_sys_fair<0>_out  & ~n789;
  assign n791 = ~n782 & ~n790;
  assign n792 = ~reg_i_hbusreq1_out & ~n791;
  assign n793 = ~n785 & ~n792;
  assign n794 = ~reg_i_hbusreq0_out & ~n793;
  assign n795 = ~n784 & ~n794;
  assign n796 = ~reg_controllable_nhgrant0_out & ~n795;
  assign n797 = ~n771 & ~n796;
  assign n798 = ~reg_controllable_hgrant1_out & ~n797;
  assign n799 = ~n770 & ~n798;
  assign n800 = ~reg_controllable_hmastlock_out & ~n799;
  assign n801 = ~n726 & ~n800;
  assign n802 = reg_i_hlock0_out & ~n801;
  assign n803 = ~reg_i_hready_out & ~n269;
  assign n804 = next_sys_fair<1>_out  & ~n803;
  assign n805 = ~n515 & ~n804;
  assign n806 = reg_controllable_locked_out & ~n805;
  assign n807 = ~n91 & ~n269;
  assign n808 = next_sys_fair<1>_out  & ~n807;
  assign n809 = ~n97 & ~n808;
  assign n810 = ~reg_controllable_locked_out & ~n809;
  assign n811 = ~n806 & ~n810;
  assign n812 = next_sys_fair<0>_out  & ~n811;
  assign n813 = reg_controllable_locked_out & ~n512;
  assign n814 = ~n88 & ~n503;
  assign n815 = next_sys_fair<1>_out  & ~n814;
  assign n816 = ~n110 & ~n815;
  assign n817 = ~reg_controllable_locked_out & ~n816;
  assign n818 = ~n813 & ~n817;
  assign n819 = ~next_sys_fair<0>_out  & ~n818;
  assign n820 = ~n812 & ~n819;
  assign n821 = reg_controllable_nhgrant0_out & ~n820;
  assign n822 = next_sys_fair<0>_out  & ~n805;
  assign n823 = ~next_sys_fair<0>_out  & ~n512;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~reg_controllable_nhgrant0_out & ~n824;
  assign n826 = ~n821 & ~n825;
  assign n827 = reg_controllable_hgrant1_out & ~n826;
  assign n828 = reg_controllable_nhgrant0_out & ~n824;
  assign n829 = next_sys_fair<1>_out  & ~n268;
  assign n830 = ~n491 & ~n829;
  assign n831 = reg_controllable_locked_out & ~n830;
  assign n832 = ~n269 & ~n531;
  assign n833 = next_sys_fair<1>_out  & ~n832;
  assign n834 = ~n97 & ~n833;
  assign n835 = ~reg_controllable_locked_out & ~n834;
  assign n836 = ~n831 & ~n835;
  assign n837 = next_sys_fair<0>_out  & ~n836;
  assign n838 = reg_controllable_locked_out & ~n87;
  assign n839 = ~n277 & ~n838;
  assign n840 = ~next_sys_fair<0>_out  & ~n839;
  assign n841 = ~n837 & ~n840;
  assign n842 = reg_i_hbusreq0_out & ~n841;
  assign n843 = reg_i_hbusreq1_out & ~n841;
  assign n844 = ~n273 & ~n831;
  assign n845 = next_sys_fair<0>_out  & ~n844;
  assign n846 = ~n840 & ~n845;
  assign n847 = ~reg_i_hbusreq1_out & ~n846;
  assign n848 = ~n843 & ~n847;
  assign n849 = ~reg_i_hbusreq0_out & ~n848;
  assign n850 = ~n842 & ~n849;
  assign n851 = ~reg_controllable_nhgrant0_out & ~n850;
  assign n852 = ~n828 & ~n851;
  assign n853 = ~reg_controllable_hgrant1_out & ~n852;
  assign n854 = ~n827 & ~n853;
  assign n855 = reg_controllable_hmastlock_out & ~n854;
  assign n856 = fair_cnt<2>_out  & ~n231;
  assign n857 = ~n190 & ~n856;
  assign n858 = ~reg_stateA1_out & ~n857;
  assign n859 = ~n236 & ~n858;
  assign n860 = ~reg_i_hready_out & ~n859;
  assign n861 = ~reg_i_hready_out & ~n860;
  assign n862 = next_sys_fair<1>_out  & ~n861;
  assign n863 = ~n639 & ~n862;
  assign n864 = reg_controllable_locked_out & ~n863;
  assign n865 = ~n91 & ~n860;
  assign n866 = next_sys_fair<1>_out  & ~n865;
  assign n867 = ~n91 & ~n637;
  assign n868 = ~next_sys_fair<1>_out  & ~n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = ~reg_controllable_locked_out & ~n869;
  assign n871 = ~n864 & ~n870;
  assign n872 = next_sys_fair<0>_out  & ~n871;
  assign n873 = ~n503 & ~n650;
  assign n874 = next_sys_fair<1>_out  & ~n873;
  assign n875 = ~n91 & ~n650;
  assign n876 = ~next_sys_fair<1>_out  & ~n875;
  assign n877 = ~n874 & ~n876;
  assign n878 = ~reg_controllable_locked_out & ~n877;
  assign n879 = ~n652 & ~n878;
  assign n880 = ~next_sys_fair<0>_out  & ~n879;
  assign n881 = ~n872 & ~n880;
  assign n882 = reg_i_hbusreq0_out & ~n881;
  assign n883 = reg_i_hbusreq1_out & ~n881;
  assign n884 = ~reg_i_hready_out & ~n235;
  assign n885 = ~reg_i_hready_out & ~n884;
  assign n886 = next_sys_fair<1>_out  & ~n885;
  assign n887 = ~n639 & ~n886;
  assign n888 = reg_controllable_locked_out & ~n887;
  assign n889 = ~n91 & ~n884;
  assign n890 = next_sys_fair<1>_out  & ~n889;
  assign n891 = ~n868 & ~n890;
  assign n892 = ~reg_controllable_locked_out & ~n891;
  assign n893 = ~n888 & ~n892;
  assign n894 = next_sys_fair<0>_out  & ~n893;
  assign n895 = ~n880 & ~n894;
  assign n896 = ~reg_i_hbusreq1_out & ~n895;
  assign n897 = ~n883 & ~n896;
  assign n898 = ~reg_i_hbusreq0_out & ~n897;
  assign n899 = ~n882 & ~n898;
  assign n900 = reg_controllable_nhgrant0_out & ~n899;
  assign n901 = next_sys_fair<0>_out  & ~n863;
  assign n902 = ~n682 & ~n901;
  assign n903 = reg_i_hbusreq0_out & ~n902;
  assign n904 = reg_i_hbusreq1_out & ~n902;
  assign n905 = next_sys_fair<0>_out  & ~n887;
  assign n906 = ~n682 & ~n905;
  assign n907 = ~reg_i_hbusreq1_out & ~n906;
  assign n908 = ~n904 & ~n907;
  assign n909 = ~reg_i_hbusreq0_out & ~n908;
  assign n910 = ~n903 & ~n909;
  assign n911 = ~reg_controllable_nhgrant0_out & ~n910;
  assign n912 = ~n900 & ~n911;
  assign n913 = reg_controllable_hgrant1_out & ~n912;
  assign n914 = reg_controllable_nhgrant0_out & ~n910;
  assign n915 = next_sys_fair<1>_out  & ~n859;
  assign n916 = ~n264 & ~n915;
  assign n917 = ~reg_controllable_locked_out & ~n916;
  assign n918 = ~n864 & ~n917;
  assign n919 = next_sys_fair<0>_out  & ~n918;
  assign n920 = ~n301 & ~n652;
  assign n921 = ~next_sys_fair<0>_out  & ~n920;
  assign n922 = ~n919 & ~n921;
  assign n923 = reg_i_hbusreq0_out & ~n922;
  assign n924 = reg_i_hbusreq1_out & ~n922;
  assign n925 = ~n297 & ~n888;
  assign n926 = next_sys_fair<0>_out  & ~n925;
  assign n927 = ~n921 & ~n926;
  assign n928 = ~reg_i_hbusreq1_out & ~n927;
  assign n929 = ~n924 & ~n928;
  assign n930 = ~reg_i_hbusreq0_out & ~n929;
  assign n931 = ~n923 & ~n930;
  assign n932 = ~reg_controllable_nhgrant0_out & ~n931;
  assign n933 = ~n914 & ~n932;
  assign n934 = ~reg_controllable_hgrant1_out & ~n933;
  assign n935 = ~n913 & ~n934;
  assign n936 = ~reg_controllable_hmastlock_out & ~n935;
  assign n937 = ~n855 & ~n936;
  assign n938 = ~reg_i_hlock0_out & ~n937;
  assign n939 = ~n802 & ~n938;
  assign n940 = ~reg_stateG2_out & ~n939;
  assign n941 = ~n630 & ~n940;
  assign n942 = ~reg_controllable_hmaster0_out & ~n941;
  assign n943 = ~n573 & ~n942;
  assign n944 = reg_i_hlock1_out & ~n943;
  assign n945 = reg_controllable_locked_out & ~n330;
  assign n946 = ~reg_controllable_locked_out & ~n322;
  assign n947 = ~n945 & ~n946;
  assign n948 = next_sys_fair<0>_out  & ~n947;
  assign n949 = next_env_fair_out & ~n157;
  assign n950 = ~next_env_fair_out & ~n103;
  assign n951 = ~n949 & ~n950;
  assign n952 = fair_cnt<2>_out  & ~n951;
  assign n953 = ~n86 & ~n952;
  assign n954 = reg_stateA1_out & ~n953;
  assign n955 = reg_stateA1_out & ~n954;
  assign n956 = ~reg_i_hready_out & ~n955;
  assign n957 = ~reg_i_hready_out & ~n956;
  assign n958 = next_sys_fair<1>_out  & ~n957;
  assign n959 = ~n353 & ~n958;
  assign n960 = reg_controllable_locked_out & ~n959;
  assign n961 = next_sys_fair<1>_out  & ~n955;
  assign n962 = ~n345 & ~n961;
  assign n963 = ~reg_controllable_locked_out & ~n962;
  assign n964 = ~n960 & ~n963;
  assign n965 = ~next_sys_fair<0>_out  & ~n964;
  assign n966 = ~n948 & ~n965;
  assign n967 = reg_i_hbusreq0_out & ~n966;
  assign n968 = reg_i_hbusreq1_out & ~n966;
  assign n969 = reg_i_hbusreq1_out & ~n968;
  assign n970 = ~reg_i_hbusreq0_out & ~n969;
  assign n971 = ~n967 & ~n970;
  assign n972 = reg_controllable_nhgrant0_out & ~n971;
  assign n973 = ~next_sys_fair<0>_out  & ~n959;
  assign n974 = ~n365 & ~n973;
  assign n975 = reg_i_hbusreq0_out & ~n974;
  assign n976 = reg_i_hbusreq1_out & ~n974;
  assign n977 = reg_i_hbusreq1_out & ~n976;
  assign n978 = ~reg_i_hbusreq0_out & ~n977;
  assign n979 = ~n975 & ~n978;
  assign n980 = ~reg_controllable_nhgrant0_out & ~n979;
  assign n981 = ~n972 & ~n980;
  assign n982 = reg_controllable_hgrant1_out & ~n981;
  assign n983 = ~reg_controllable_hgrant1_out & ~n979;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~reg_controllable_hmastlock_out & ~n984;
  assign n986 = ~reg_controllable_hmastlock_out & ~n985;
  assign n987 = reg_stateG2_out & ~n986;
  assign n988 = reg_i_hready_out & ~n91;
  assign n989 = ~reg_controllable_locked_out & ~n988;
  assign n990 = ~reg_controllable_locked_out & ~n989;
  assign n991 = next_sys_fair<0>_out  & ~n990;
  assign n992 = reg_i_hready_out & ~n531;
  assign n993 = next_sys_fair<1>_out  & ~n992;
  assign n994 = ~next_sys_fair<1>_out  & ~n988;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~reg_controllable_locked_out & ~n995;
  assign n997 = ~reg_controllable_locked_out & ~n996;
  assign n998 = ~next_sys_fair<0>_out  & ~n997;
  assign n999 = ~n991 & ~n998;
  assign n1000 = reg_i_hbusreq0_out & ~n999;
  assign n1001 = reg_i_hbusreq1_out & ~n999;
  assign n1002 = ~reg_i_hbusreq1_out & ~n397;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~reg_i_hbusreq0_out & ~n1003;
  assign n1005 = ~n1000 & ~n1004;
  assign n1006 = reg_controllable_nhgrant0_out & ~n1005;
  assign n1007 = reg_controllable_nhgrant0_out & ~n1006;
  assign n1008 = reg_controllable_hgrant1_out & ~n1007;
  assign n1009 = ~n427 & ~n1008;
  assign n1010 = reg_controllable_hmastlock_out & ~n1009;
  assign n1011 = ~n135 & ~n954;
  assign n1012 = ~reg_i_hready_out & ~n1011;
  assign n1013 = ~reg_i_hready_out & ~n1012;
  assign n1014 = next_sys_fair<1>_out  & ~n1013;
  assign n1015 = ~n520 & ~n1014;
  assign n1016 = reg_controllable_locked_out & ~n1015;
  assign n1017 = next_sys_fair<1>_out  & ~n1011;
  assign n1018 = ~n500 & ~n1017;
  assign n1019 = ~reg_controllable_locked_out & ~n1018;
  assign n1020 = ~n1016 & ~n1019;
  assign n1021 = ~next_sys_fair<0>_out  & ~n1020;
  assign n1022 = ~n558 & ~n1021;
  assign n1023 = reg_i_hbusreq0_out & ~n1022;
  assign n1024 = reg_i_hbusreq1_out & ~n1022;
  assign n1025 = ~reg_i_hbusreq1_out & ~n453;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~reg_i_hbusreq0_out & ~n1026;
  assign n1028 = ~n1023 & ~n1027;
  assign n1029 = reg_controllable_nhgrant0_out & ~n1028;
  assign n1030 = ~next_sys_fair<0>_out  & ~n1015;
  assign n1031 = ~n517 & ~n1030;
  assign n1032 = reg_i_hbusreq0_out & ~n1031;
  assign n1033 = reg_i_hbusreq1_out & ~n1031;
  assign n1034 = ~reg_i_hbusreq1_out & ~n457;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = ~reg_i_hbusreq0_out & ~n1035;
  assign n1037 = ~n1032 & ~n1036;
  assign n1038 = ~reg_controllable_nhgrant0_out & ~n1037;
  assign n1039 = ~n1029 & ~n1038;
  assign n1040 = reg_controllable_hgrant1_out & ~n1039;
  assign n1041 = reg_controllable_nhgrant0_out & ~n1037;
  assign n1042 = ~n57 & ~n88;
  assign n1043 = next_sys_fair<1>_out  & ~n1042;
  assign n1044 = ~n68 & ~n95;
  assign n1045 = ~next_sys_fair<1>_out  & ~n1044;
  assign n1046 = ~n1043 & ~n1045;
  assign n1047 = reg_controllable_locked_out & ~n1046;
  assign n1048 = ~n88 & ~n390;
  assign n1049 = next_sys_fair<1>_out  & ~n1048;
  assign n1050 = ~n1045 & ~n1049;
  assign n1051 = ~reg_controllable_locked_out & ~n1050;
  assign n1052 = ~n1047 & ~n1051;
  assign n1053 = next_sys_fair<0>_out  & ~n1052;
  assign n1054 = ~n68 & ~n1012;
  assign n1055 = next_sys_fair<1>_out  & ~n1054;
  assign n1056 = ~n68 & ~n88;
  assign n1057 = ~next_sys_fair<1>_out  & ~n1056;
  assign n1058 = ~n1055 & ~n1057;
  assign n1059 = ~next_sys_fair<0>_out  & ~n1058;
  assign n1060 = ~n1053 & ~n1059;
  assign n1061 = reg_i_hbusreq0_out & ~n1060;
  assign n1062 = reg_i_hbusreq1_out & ~n1060;
  assign n1063 = ~n479 & ~n1062;
  assign n1064 = ~reg_i_hbusreq0_out & ~n1063;
  assign n1065 = ~n1061 & ~n1064;
  assign n1066 = ~reg_controllable_nhgrant0_out & ~n1065;
  assign n1067 = ~n1041 & ~n1066;
  assign n1068 = ~reg_controllable_hgrant1_out & ~n1067;
  assign n1069 = ~n1040 & ~n1068;
  assign n1070 = ~reg_controllable_hmastlock_out & ~n1069;
  assign n1071 = ~n1010 & ~n1070;
  assign n1072 = reg_i_hlock0_out & ~n1071;
  assign n1073 = ~n97 & ~n815;
  assign n1074 = ~reg_controllable_locked_out & ~n1073;
  assign n1075 = ~n528 & ~n1074;
  assign n1076 = next_sys_fair<0>_out  & ~n1075;
  assign n1077 = ~n540 & ~n1076;
  assign n1078 = reg_i_hbusreq0_out & ~n1077;
  assign n1079 = reg_i_hbusreq1_out & ~n1077;
  assign n1080 = ~n547 & ~n1079;
  assign n1081 = ~reg_i_hbusreq0_out & ~n1080;
  assign n1082 = ~n1078 & ~n1081;
  assign n1083 = ~reg_controllable_nhgrant0_out & ~n1082;
  assign n1084 = ~n527 & ~n1083;
  assign n1085 = ~reg_controllable_hgrant1_out & ~n1084;
  assign n1086 = ~n526 & ~n1085;
  assign n1087 = reg_controllable_hmastlock_out & ~n1086;
  assign n1088 = ~n565 & ~n1085;
  assign n1089 = ~reg_controllable_hmastlock_out & ~n1088;
  assign n1090 = ~n1087 & ~n1089;
  assign n1091 = ~reg_i_hlock0_out & ~n1090;
  assign n1092 = ~n1072 & ~n1091;
  assign n1093 = ~reg_stateG2_out & ~n1092;
  assign n1094 = ~n987 & ~n1093;
  assign n1095 = reg_controllable_hmaster0_out & ~n1094;
  assign n1096 = ~n104 & ~n179;
  assign n1097 = ~reg_i_hready_out & ~n1096;
  assign n1098 = ~reg_i_hready_out & ~n1097;
  assign n1099 = next_sys_fair<1>_out  & ~n1098;
  assign n1100 = ~n639 & ~n1099;
  assign n1101 = reg_controllable_locked_out & ~n1100;
  assign n1102 = ~n91 & ~n1097;
  assign n1103 = next_sys_fair<1>_out  & ~n1102;
  assign n1104 = ~n868 & ~n1103;
  assign n1105 = ~reg_controllable_locked_out & ~n1104;
  assign n1106 = ~n1101 & ~n1105;
  assign n1107 = next_sys_fair<0>_out  & ~n1106;
  assign n1108 = ~n531 & ~n650;
  assign n1109 = next_sys_fair<1>_out  & ~n1108;
  assign n1110 = ~n876 & ~n1109;
  assign n1111 = ~reg_controllable_locked_out & ~n1110;
  assign n1112 = ~n652 & ~n1111;
  assign n1113 = ~next_sys_fair<0>_out  & ~n1112;
  assign n1114 = ~n1107 & ~n1113;
  assign n1115 = reg_i_hbusreq0_out & ~n1114;
  assign n1116 = reg_i_hbusreq1_out & ~n1114;
  assign n1117 = ~n676 & ~n1116;
  assign n1118 = ~reg_i_hbusreq0_out & ~n1117;
  assign n1119 = ~n1115 & ~n1118;
  assign n1120 = reg_controllable_nhgrant0_out & ~n1119;
  assign n1121 = next_sys_fair<0>_out  & ~n1100;
  assign n1122 = ~n682 & ~n1121;
  assign n1123 = reg_i_hbusreq0_out & ~n1122;
  assign n1124 = reg_i_hbusreq1_out & ~n1122;
  assign n1125 = ~n688 & ~n1124;
  assign n1126 = ~reg_i_hbusreq0_out & ~n1125;
  assign n1127 = ~n1123 & ~n1126;
  assign n1128 = ~reg_controllable_nhgrant0_out & ~n1127;
  assign n1129 = ~n1120 & ~n1128;
  assign n1130 = reg_controllable_hgrant1_out & ~n1129;
  assign n1131 = reg_controllable_nhgrant0_out & ~n1127;
  assign n1132 = next_sys_fair<1>_out  & ~n1096;
  assign n1133 = ~n264 & ~n1132;
  assign n1134 = reg_controllable_locked_out & ~n1133;
  assign n1135 = ~n390 & ~n1097;
  assign n1136 = next_sys_fair<1>_out  & ~n1135;
  assign n1137 = ~n645 & ~n1136;
  assign n1138 = ~reg_controllable_locked_out & ~n1137;
  assign n1139 = ~n1134 & ~n1138;
  assign n1140 = next_sys_fair<0>_out  & ~n1139;
  assign n1141 = ~n707 & ~n1140;
  assign n1142 = reg_i_hbusreq0_out & ~n1141;
  assign n1143 = reg_i_hbusreq1_out & ~n1141;
  assign n1144 = ~n718 & ~n1143;
  assign n1145 = ~reg_i_hbusreq0_out & ~n1144;
  assign n1146 = ~n1142 & ~n1145;
  assign n1147 = ~reg_controllable_nhgrant0_out & ~n1146;
  assign n1148 = ~n1131 & ~n1147;
  assign n1149 = ~reg_controllable_hgrant1_out & ~n1148;
  assign n1150 = ~n1130 & ~n1149;
  assign n1151 = reg_controllable_hmastlock_out & ~n1150;
  assign n1152 = ~n91 & ~n137;
  assign n1153 = next_sys_fair<1>_out  & ~n1152;
  assign n1154 = ~n91 & ~n128;
  assign n1155 = ~next_sys_fair<1>_out  & ~n1154;
  assign n1156 = ~n1153 & ~n1155;
  assign n1157 = ~reg_controllable_locked_out & ~n1156;
  assign n1158 = ~n728 & ~n1157;
  assign n1159 = next_sys_fair<0>_out  & ~n1158;
  assign n1160 = ~n123 & ~n531;
  assign n1161 = next_sys_fair<1>_out  & ~n1160;
  assign n1162 = ~n91 & ~n123;
  assign n1163 = ~next_sys_fair<1>_out  & ~n1162;
  assign n1164 = ~n1161 & ~n1163;
  assign n1165 = ~reg_controllable_locked_out & ~n1164;
  assign n1166 = ~n733 & ~n1165;
  assign n1167 = ~next_sys_fair<0>_out  & ~n1166;
  assign n1168 = ~n1159 & ~n1167;
  assign n1169 = reg_i_hbusreq0_out & ~n1168;
  assign n1170 = reg_i_hbusreq1_out & ~n1168;
  assign n1171 = ~n752 & ~n1170;
  assign n1172 = ~reg_i_hbusreq0_out & ~n1171;
  assign n1173 = ~n1169 & ~n1172;
  assign n1174 = reg_controllable_nhgrant0_out & ~n1173;
  assign n1175 = ~n768 & ~n1174;
  assign n1176 = reg_controllable_hgrant1_out & ~n1175;
  assign n1177 = ~n798 & ~n1176;
  assign n1178 = ~reg_controllable_hmastlock_out & ~n1177;
  assign n1179 = ~n1151 & ~n1178;
  assign n1180 = reg_i_hlock0_out & ~n1179;
  assign n1181 = ~n515 & ~n519;
  assign n1182 = reg_controllable_locked_out & ~n1181;
  assign n1183 = ~n97 & ~n108;
  assign n1184 = ~reg_controllable_locked_out & ~n1183;
  assign n1185 = ~n1182 & ~n1184;
  assign n1186 = next_sys_fair<0>_out  & ~n1185;
  assign n1187 = ~n819 & ~n1186;
  assign n1188 = reg_i_hbusreq0_out & ~n1187;
  assign n1189 = reg_i_hbusreq1_out & ~n1187;
  assign n1190 = ~reg_i_hbusreq1_out & ~n820;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~reg_i_hbusreq0_out & ~n1191;
  assign n1193 = ~n1188 & ~n1192;
  assign n1194 = reg_controllable_nhgrant0_out & ~n1193;
  assign n1195 = next_sys_fair<0>_out  & ~n1181;
  assign n1196 = ~n823 & ~n1195;
  assign n1197 = reg_i_hbusreq0_out & ~n1196;
  assign n1198 = reg_i_hbusreq1_out & ~n1196;
  assign n1199 = ~reg_i_hbusreq1_out & ~n824;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~reg_i_hbusreq0_out & ~n1200;
  assign n1202 = ~n1197 & ~n1201;
  assign n1203 = ~reg_controllable_nhgrant0_out & ~n1202;
  assign n1204 = ~n1194 & ~n1203;
  assign n1205 = reg_controllable_hgrant1_out & ~n1204;
  assign n1206 = reg_controllable_nhgrant0_out & ~n1202;
  assign n1207 = ~n491 & ~n499;
  assign n1208 = reg_controllable_locked_out & ~n1207;
  assign n1209 = ~n97 & ~n505;
  assign n1210 = ~reg_controllable_locked_out & ~n1209;
  assign n1211 = ~n1208 & ~n1210;
  assign n1212 = next_sys_fair<0>_out  & ~n1211;
  assign n1213 = ~n840 & ~n1212;
  assign n1214 = reg_i_hbusreq0_out & ~n1213;
  assign n1215 = reg_i_hbusreq1_out & ~n1213;
  assign n1216 = ~n847 & ~n1215;
  assign n1217 = ~reg_i_hbusreq0_out & ~n1216;
  assign n1218 = ~n1214 & ~n1217;
  assign n1219 = ~reg_controllable_nhgrant0_out & ~n1218;
  assign n1220 = ~n1206 & ~n1219;
  assign n1221 = ~reg_controllable_hgrant1_out & ~n1220;
  assign n1222 = ~n1205 & ~n1221;
  assign n1223 = reg_controllable_hmastlock_out & ~n1222;
  assign n1224 = ~reg_i_hready_out & ~n857;
  assign n1225 = ~reg_i_hready_out & ~n1224;
  assign n1226 = next_sys_fair<1>_out  & ~n1225;
  assign n1227 = ~n639 & ~n1226;
  assign n1228 = reg_controllable_locked_out & ~n1227;
  assign n1229 = ~n91 & ~n1224;
  assign n1230 = next_sys_fair<1>_out  & ~n1229;
  assign n1231 = ~n868 & ~n1230;
  assign n1232 = ~reg_controllable_locked_out & ~n1231;
  assign n1233 = ~n1228 & ~n1232;
  assign n1234 = next_sys_fair<0>_out  & ~n1233;
  assign n1235 = ~n880 & ~n1234;
  assign n1236 = reg_i_hbusreq0_out & ~n1235;
  assign n1237 = reg_i_hbusreq1_out & ~n1235;
  assign n1238 = ~n896 & ~n1237;
  assign n1239 = ~reg_i_hbusreq0_out & ~n1238;
  assign n1240 = ~n1236 & ~n1239;
  assign n1241 = reg_controllable_nhgrant0_out & ~n1240;
  assign n1242 = next_sys_fair<0>_out  & ~n1227;
  assign n1243 = ~n682 & ~n1242;
  assign n1244 = reg_i_hbusreq0_out & ~n1243;
  assign n1245 = reg_i_hbusreq1_out & ~n1243;
  assign n1246 = ~n907 & ~n1245;
  assign n1247 = ~reg_i_hbusreq0_out & ~n1246;
  assign n1248 = ~n1244 & ~n1247;
  assign n1249 = ~reg_controllable_nhgrant0_out & ~n1248;
  assign n1250 = ~n1241 & ~n1249;
  assign n1251 = reg_controllable_hgrant1_out & ~n1250;
  assign n1252 = reg_controllable_nhgrant0_out & ~n1248;
  assign n1253 = next_sys_fair<1>_out  & ~n857;
  assign n1254 = ~n264 & ~n1253;
  assign n1255 = ~reg_controllable_locked_out & ~n1254;
  assign n1256 = ~n1228 & ~n1255;
  assign n1257 = next_sys_fair<0>_out  & ~n1256;
  assign n1258 = ~n921 & ~n1257;
  assign n1259 = reg_i_hbusreq0_out & ~n1258;
  assign n1260 = reg_i_hbusreq1_out & ~n1258;
  assign n1261 = ~n928 & ~n1260;
  assign n1262 = ~reg_i_hbusreq0_out & ~n1261;
  assign n1263 = ~n1259 & ~n1262;
  assign n1264 = ~reg_controllable_nhgrant0_out & ~n1263;
  assign n1265 = ~n1252 & ~n1264;
  assign n1266 = ~reg_controllable_hgrant1_out & ~n1265;
  assign n1267 = ~n1251 & ~n1266;
  assign n1268 = ~reg_controllable_hmastlock_out & ~n1267;
  assign n1269 = ~n1223 & ~n1268;
  assign n1270 = ~reg_i_hlock0_out & ~n1269;
  assign n1271 = ~n1180 & ~n1270;
  assign n1272 = ~reg_stateG2_out & ~n1271;
  assign n1273 = ~n630 & ~n1272;
  assign n1274 = ~reg_controllable_hmaster0_out & ~n1273;
  assign n1275 = ~n1095 & ~n1274;
  assign n1276 = ~reg_i_hlock1_out & ~n1275;
  assign n1277 = ~n944 & ~n1276;
  assign n1278 = ~reg_controllable_ndecide_out & ~n1277;
  assign n1279 = ~n315 & ~n1278;
  assign n1280 = reg_stateG10_1_out & ~n1279;
  assign n1281 = ~n194 & ~n207;
  assign n1282 = reg_controllable_locked_out & ~n1281;
  assign n1283 = reg_controllable_locked_out & ~n1282;
  assign n1284 = next_sys_fair<0>_out  & ~n1283;
  assign n1285 = ~n183 & ~n216;
  assign n1286 = reg_controllable_locked_out & ~n1285;
  assign n1287 = reg_controllable_locked_out & ~n1286;
  assign n1288 = ~next_sys_fair<0>_out  & ~n1287;
  assign n1289 = ~n1284 & ~n1288;
  assign n1290 = reg_controllable_nhgrant0_out & ~n1289;
  assign n1291 = reg_controllable_nhgrant0_out & ~n1290;
  assign n1292 = reg_controllable_hgrant1_out & ~n1291;
  assign n1293 = reg_controllable_hgrant1_out & ~n1292;
  assign n1294 = reg_controllable_hmastlock_out & ~n1293;
  assign n1295 = ~reg_controllable_locked_out & ~n1281;
  assign n1296 = ~reg_controllable_locked_out & ~n1295;
  assign n1297 = next_sys_fair<0>_out  & ~n1296;
  assign n1298 = ~n216 & ~n238;
  assign n1299 = ~reg_controllable_locked_out & ~n1298;
  assign n1300 = ~reg_controllable_locked_out & ~n1299;
  assign n1301 = ~next_sys_fair<0>_out  & ~n1300;
  assign n1302 = ~n1297 & ~n1301;
  assign n1303 = reg_controllable_nhgrant0_out & ~n1302;
  assign n1304 = reg_controllable_nhgrant0_out & ~n1303;
  assign n1305 = reg_controllable_hgrant1_out & ~n1304;
  assign n1306 = reg_controllable_hgrant1_out & ~n1305;
  assign n1307 = ~reg_controllable_hmastlock_out & ~n1306;
  assign n1308 = ~n1294 & ~n1307;
  assign n1309 = reg_stateG2_out & ~n1308;
  assign n1310 = next_sys_fair<1>_out  & ~n204;
  assign n1311 = ~n264 & ~n1310;
  assign n1312 = reg_controllable_locked_out & ~n1311;
  assign n1313 = ~n496 & ~n1312;
  assign n1314 = next_sys_fair<0>_out  & ~n1313;
  assign n1315 = ~next_sys_fair<1>_out  & ~n204;
  assign n1316 = ~n263 & ~n1315;
  assign n1317 = reg_controllable_locked_out & ~n1316;
  assign n1318 = ~n110 & ~n271;
  assign n1319 = ~reg_controllable_locked_out & ~n1318;
  assign n1320 = ~n1317 & ~n1319;
  assign n1321 = ~next_sys_fair<0>_out  & ~n1320;
  assign n1322 = ~n1314 & ~n1321;
  assign n1323 = reg_controllable_nhgrant0_out & ~n1322;
  assign n1324 = reg_controllable_nhgrant0_out & ~n1323;
  assign n1325 = reg_controllable_hgrant1_out & ~n1324;
  assign n1326 = ~n118 & ~n1325;
  assign n1327 = reg_controllable_hmastlock_out & ~n1326;
  assign n1328 = next_sys_fair<1>_out  & ~n140;
  assign n1329 = ~n130 & ~n1328;
  assign n1330 = reg_controllable_locked_out & ~n1329;
  assign n1331 = ~reg_controllable_locked_out & ~n1311;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = next_sys_fair<0>_out  & ~n1332;
  assign n1334 = ~n141 & ~n292;
  assign n1335 = reg_controllable_locked_out & ~n1334;
  assign n1336 = ~n295 & ~n1315;
  assign n1337 = ~reg_controllable_locked_out & ~n1336;
  assign n1338 = ~n1335 & ~n1337;
  assign n1339 = ~next_sys_fair<0>_out  & ~n1338;
  assign n1340 = ~n1333 & ~n1339;
  assign n1341 = reg_controllable_nhgrant0_out & ~n1340;
  assign n1342 = reg_controllable_nhgrant0_out & ~n1341;
  assign n1343 = reg_controllable_hgrant1_out & ~n1342;
  assign n1344 = ~n149 & ~n1343;
  assign n1345 = ~reg_controllable_hmastlock_out & ~n1344;
  assign n1346 = ~n1327 & ~n1345;
  assign n1347 = ~reg_stateG2_out & ~n1346;
  assign n1348 = ~n1309 & ~n1347;
  assign n1349 = reg_controllable_hmaster0_out & ~n1348;
  assign n1350 = ~n102 & ~n1184;
  assign n1351 = next_sys_fair<0>_out  & ~n1350;
  assign n1352 = ~n90 & ~n110;
  assign n1353 = ~reg_controllable_locked_out & ~n1352;
  assign n1354 = ~n72 & ~n1353;
  assign n1355 = ~next_sys_fair<0>_out  & ~n1354;
  assign n1356 = ~n1351 & ~n1355;
  assign n1357 = reg_controllable_nhgrant0_out & ~n1356;
  assign n1358 = reg_controllable_nhgrant0_out & ~n1357;
  assign n1359 = reg_controllable_hgrant1_out & ~n1358;
  assign n1360 = ~n283 & ~n1359;
  assign n1361 = reg_controllable_hmastlock_out & ~n1360;
  assign n1362 = reg_controllable_locked_out & ~n729;
  assign n1363 = ~n1184 & ~n1362;
  assign n1364 = next_sys_fair<0>_out  & ~n1363;
  assign n1365 = ~n125 & ~n141;
  assign n1366 = reg_controllable_locked_out & ~n1365;
  assign n1367 = ~n1353 & ~n1366;
  assign n1368 = ~next_sys_fair<0>_out  & ~n1367;
  assign n1369 = ~n1364 & ~n1368;
  assign n1370 = reg_controllable_nhgrant0_out & ~n1369;
  assign n1371 = reg_controllable_nhgrant0_out & ~n1370;
  assign n1372 = reg_controllable_hgrant1_out & ~n1371;
  assign n1373 = ~n307 & ~n1372;
  assign n1374 = ~reg_controllable_hmastlock_out & ~n1373;
  assign n1375 = ~n1361 & ~n1374;
  assign n1376 = ~reg_stateG2_out & ~n1375;
  assign n1377 = ~n253 & ~n1376;
  assign n1378 = ~reg_controllable_hmaster0_out & ~n1377;
  assign n1379 = ~n1349 & ~n1378;
  assign n1380 = reg_controllable_ndecide_out & ~n1379;
  assign n1381 = ~n579 & ~n584;
  assign n1382 = ~reg_controllable_locked_out & ~n1381;
  assign n1383 = ~n1282 & ~n1382;
  assign n1384 = next_sys_fair<0>_out  & ~n1383;
  assign n1385 = ~n576 & ~n587;
  assign n1386 = ~reg_controllable_locked_out & ~n1385;
  assign n1387 = ~n1286 & ~n1386;
  assign n1388 = ~next_sys_fair<0>_out  & ~n1387;
  assign n1389 = ~n1384 & ~n1388;
  assign n1390 = reg_i_hbusreq0_out & ~n1389;
  assign n1391 = reg_i_hbusreq1_out & ~n1389;
  assign n1392 = reg_i_hbusreq1_out & ~n1391;
  assign n1393 = ~reg_i_hbusreq0_out & ~n1392;
  assign n1394 = ~n1390 & ~n1393;
  assign n1395 = reg_controllable_nhgrant0_out & ~n1394;
  assign n1396 = next_sys_fair<0>_out  & ~n1381;
  assign n1397 = ~next_sys_fair<0>_out  & ~n1385;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = reg_i_hbusreq0_out & ~n1398;
  assign n1400 = reg_i_hbusreq1_out & ~n1398;
  assign n1401 = reg_i_hbusreq1_out & ~n1400;
  assign n1402 = ~reg_i_hbusreq0_out & ~n1401;
  assign n1403 = ~n1399 & ~n1402;
  assign n1404 = ~reg_controllable_nhgrant0_out & ~n1403;
  assign n1405 = ~n1395 & ~n1404;
  assign n1406 = reg_controllable_hgrant1_out & ~n1405;
  assign n1407 = ~reg_controllable_hgrant1_out & ~n1403;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = reg_controllable_hmastlock_out & ~n1408;
  assign n1410 = reg_controllable_hmastlock_out & ~n1409;
  assign n1411 = reg_stateG2_out & ~n1410;
  assign n1412 = next_sys_fair<1>_out  & ~n655;
  assign n1413 = ~n645 & ~n1412;
  assign n1414 = ~reg_controllable_locked_out & ~n1413;
  assign n1415 = ~n1312 & ~n1414;
  assign n1416 = next_sys_fair<0>_out  & ~n1415;
  assign n1417 = ~n696 & ~n1315;
  assign n1418 = reg_controllable_locked_out & ~n1417;
  assign n1419 = ~n656 & ~n700;
  assign n1420 = ~reg_controllable_locked_out & ~n1419;
  assign n1421 = ~n1418 & ~n1420;
  assign n1422 = ~next_sys_fair<0>_out  & ~n1421;
  assign n1423 = ~n1416 & ~n1422;
  assign n1424 = reg_i_hbusreq0_out & ~n1423;
  assign n1425 = reg_i_hbusreq1_out & ~n1423;
  assign n1426 = ~n1002 & ~n1425;
  assign n1427 = ~reg_i_hbusreq0_out & ~n1426;
  assign n1428 = ~n1424 & ~n1427;
  assign n1429 = reg_controllable_nhgrant0_out & ~n1428;
  assign n1430 = next_sys_fair<1>_out  & ~n651;
  assign n1431 = ~n639 & ~n1430;
  assign n1432 = next_sys_fair<0>_out  & ~n1431;
  assign n1433 = ~next_sys_fair<1>_out  & ~n651;
  assign n1434 = ~n636 & ~n1433;
  assign n1435 = ~next_sys_fair<0>_out  & ~n1434;
  assign n1436 = ~n1432 & ~n1435;
  assign n1437 = reg_i_hbusreq0_out & ~n1436;
  assign n1438 = reg_i_hbusreq1_out & ~n1436;
  assign n1439 = reg_i_hbusreq1_out & ~n1438;
  assign n1440 = ~reg_i_hbusreq0_out & ~n1439;
  assign n1441 = ~n1437 & ~n1440;
  assign n1442 = ~reg_controllable_nhgrant0_out & ~n1441;
  assign n1443 = ~n1429 & ~n1442;
  assign n1444 = reg_controllable_hgrant1_out & ~n1443;
  assign n1445 = reg_controllable_nhgrant0_out & ~n1441;
  assign n1446 = ~n57 & ~n650;
  assign n1447 = next_sys_fair<1>_out  & ~n1446;
  assign n1448 = ~n645 & ~n1447;
  assign n1449 = reg_controllable_locked_out & ~n1448;
  assign n1450 = ~n645 & ~n654;
  assign n1451 = ~reg_controllable_locked_out & ~n1450;
  assign n1452 = ~n1449 & ~n1451;
  assign n1453 = next_sys_fair<0>_out  & ~n1452;
  assign n1454 = ~n643 & ~n656;
  assign n1455 = ~next_sys_fair<0>_out  & ~n1454;
  assign n1456 = ~n1453 & ~n1455;
  assign n1457 = reg_i_hbusreq0_out & ~n1456;
  assign n1458 = reg_i_hbusreq1_out & ~n1456;
  assign n1459 = ~n421 & ~n1458;
  assign n1460 = ~reg_i_hbusreq0_out & ~n1459;
  assign n1461 = ~n1457 & ~n1460;
  assign n1462 = ~reg_controllable_nhgrant0_out & ~n1461;
  assign n1463 = ~n1445 & ~n1462;
  assign n1464 = ~reg_controllable_hgrant1_out & ~n1463;
  assign n1465 = ~n1444 & ~n1464;
  assign n1466 = reg_controllable_hmastlock_out & ~n1465;
  assign n1467 = ~n439 & ~n1330;
  assign n1468 = next_sys_fair<0>_out  & ~n1467;
  assign n1469 = ~n141 & ~n773;
  assign n1470 = reg_controllable_locked_out & ~n1469;
  assign n1471 = ~n450 & ~n1470;
  assign n1472 = ~next_sys_fair<0>_out  & ~n1471;
  assign n1473 = ~n1468 & ~n1472;
  assign n1474 = reg_i_hbusreq0_out & ~n1473;
  assign n1475 = reg_i_hbusreq1_out & ~n1473;
  assign n1476 = ~n1025 & ~n1475;
  assign n1477 = ~reg_i_hbusreq0_out & ~n1476;
  assign n1478 = ~n1474 & ~n1477;
  assign n1479 = reg_controllable_nhgrant0_out & ~n1478;
  assign n1480 = ~n458 & ~n1479;
  assign n1481 = reg_controllable_hgrant1_out & ~n1480;
  assign n1482 = ~n485 & ~n1481;
  assign n1483 = ~reg_controllable_hmastlock_out & ~n1482;
  assign n1484 = ~n1466 & ~n1483;
  assign n1485 = reg_i_hlock0_out & ~n1484;
  assign n1486 = next_sys_fair<1>_out  & ~n875;
  assign n1487 = ~n868 & ~n1486;
  assign n1488 = ~reg_controllable_locked_out & ~n1487;
  assign n1489 = ~n1312 & ~n1488;
  assign n1490 = next_sys_fair<0>_out  & ~n1489;
  assign n1491 = ~n1132 & ~n1315;
  assign n1492 = reg_controllable_locked_out & ~n1491;
  assign n1493 = ~n503 & ~n1097;
  assign n1494 = next_sys_fair<1>_out  & ~n1493;
  assign n1495 = ~n876 & ~n1494;
  assign n1496 = ~reg_controllable_locked_out & ~n1495;
  assign n1497 = ~n1492 & ~n1496;
  assign n1498 = ~next_sys_fair<0>_out  & ~n1497;
  assign n1499 = ~n1490 & ~n1498;
  assign n1500 = reg_i_hbusreq0_out & ~n1499;
  assign n1501 = reg_i_hbusreq1_out & ~n1499;
  assign n1502 = ~reg_i_hbusreq1_out & ~n510;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~reg_i_hbusreq0_out & ~n1503;
  assign n1505 = ~n1500 & ~n1504;
  assign n1506 = reg_controllable_nhgrant0_out & ~n1505;
  assign n1507 = ~n1099 & ~n1433;
  assign n1508 = ~next_sys_fair<0>_out  & ~n1507;
  assign n1509 = ~n1432 & ~n1508;
  assign n1510 = reg_i_hbusreq0_out & ~n1509;
  assign n1511 = reg_i_hbusreq1_out & ~n1509;
  assign n1512 = ~reg_i_hbusreq1_out & ~n523;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = ~reg_i_hbusreq0_out & ~n1513;
  assign n1515 = ~n1510 & ~n1514;
  assign n1516 = ~reg_controllable_nhgrant0_out & ~n1515;
  assign n1517 = ~n1506 & ~n1516;
  assign n1518 = reg_controllable_hgrant1_out & ~n1517;
  assign n1519 = reg_controllable_nhgrant0_out & ~n1515;
  assign n1520 = reg_controllable_locked_out & ~n1431;
  assign n1521 = ~n868 & ~n1109;
  assign n1522 = ~reg_controllable_locked_out & ~n1521;
  assign n1523 = ~n1520 & ~n1522;
  assign n1524 = next_sys_fair<0>_out  & ~n1523;
  assign n1525 = reg_controllable_locked_out & ~n1507;
  assign n1526 = ~n876 & ~n1103;
  assign n1527 = ~reg_controllable_locked_out & ~n1526;
  assign n1528 = ~n1525 & ~n1527;
  assign n1529 = ~next_sys_fair<0>_out  & ~n1528;
  assign n1530 = ~n1524 & ~n1529;
  assign n1531 = reg_i_hbusreq0_out & ~n1530;
  assign n1532 = reg_i_hbusreq1_out & ~n1530;
  assign n1533 = ~n547 & ~n1532;
  assign n1534 = ~reg_i_hbusreq0_out & ~n1533;
  assign n1535 = ~n1531 & ~n1534;
  assign n1536 = ~reg_controllable_nhgrant0_out & ~n1535;
  assign n1537 = ~n1519 & ~n1536;
  assign n1538 = ~reg_controllable_hgrant1_out & ~n1537;
  assign n1539 = ~n1518 & ~n1538;
  assign n1540 = reg_controllable_hmastlock_out & ~n1539;
  assign n1541 = next_sys_fair<1>_out  & ~n1056;
  assign n1542 = ~n1045 & ~n1541;
  assign n1543 = reg_controllable_locked_out & ~n1542;
  assign n1544 = ~n556 & ~n1543;
  assign n1545 = next_sys_fair<0>_out  & ~n1544;
  assign n1546 = ~n57 & ~n106;
  assign n1547 = next_sys_fair<1>_out  & ~n1546;
  assign n1548 = ~n1057 & ~n1547;
  assign n1549 = reg_controllable_locked_out & ~n1548;
  assign n1550 = ~n559 & ~n1549;
  assign n1551 = ~next_sys_fair<0>_out  & ~n1550;
  assign n1552 = ~n1545 & ~n1551;
  assign n1553 = reg_i_hbusreq0_out & ~n1552;
  assign n1554 = reg_i_hbusreq1_out & ~n1552;
  assign n1555 = ~reg_i_hbusreq1_out & ~n562;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~reg_i_hbusreq0_out & ~n1556;
  assign n1558 = ~n1553 & ~n1557;
  assign n1559 = reg_controllable_nhgrant0_out & ~n1558;
  assign n1560 = ~n524 & ~n1559;
  assign n1561 = reg_controllable_hgrant1_out & ~n1560;
  assign n1562 = ~n553 & ~n1561;
  assign n1563 = ~reg_controllable_hmastlock_out & ~n1562;
  assign n1564 = ~n1540 & ~n1563;
  assign n1565 = ~reg_i_hlock0_out & ~n1564;
  assign n1566 = ~n1485 & ~n1565;
  assign n1567 = ~reg_stateG2_out & ~n1566;
  assign n1568 = ~n1411 & ~n1567;
  assign n1569 = reg_controllable_hmaster0_out & ~n1568;
  assign n1570 = next_sys_fair<0>_out  & ~n646;
  assign n1571 = ~n656 & ~n1447;
  assign n1572 = reg_controllable_locked_out & ~n1571;
  assign n1573 = ~n658 & ~n1572;
  assign n1574 = ~next_sys_fair<0>_out  & ~n1573;
  assign n1575 = ~n1570 & ~n1574;
  assign n1576 = reg_i_hbusreq0_out & ~n1575;
  assign n1577 = reg_i_hbusreq1_out & ~n1575;
  assign n1578 = ~n676 & ~n1577;
  assign n1579 = ~reg_i_hbusreq0_out & ~n1578;
  assign n1580 = ~n1576 & ~n1579;
  assign n1581 = reg_controllable_nhgrant0_out & ~n1580;
  assign n1582 = ~n692 & ~n1581;
  assign n1583 = reg_controllable_hgrant1_out & ~n1582;
  assign n1584 = ~n724 & ~n1583;
  assign n1585 = reg_controllable_hmastlock_out & ~n1584;
  assign n1586 = next_sys_fair<0>_out  & ~n729;
  assign n1587 = ~n735 & ~n1366;
  assign n1588 = ~next_sys_fair<0>_out  & ~n1587;
  assign n1589 = ~n1586 & ~n1588;
  assign n1590 = reg_i_hbusreq0_out & ~n1589;
  assign n1591 = reg_i_hbusreq1_out & ~n1589;
  assign n1592 = ~n752 & ~n1591;
  assign n1593 = ~reg_i_hbusreq0_out & ~n1592;
  assign n1594 = ~n1590 & ~n1593;
  assign n1595 = reg_controllable_nhgrant0_out & ~n1594;
  assign n1596 = ~n768 & ~n1595;
  assign n1597 = reg_controllable_hgrant1_out & ~n1596;
  assign n1598 = ~n798 & ~n1597;
  assign n1599 = ~reg_controllable_hmastlock_out & ~n1598;
  assign n1600 = ~n1585 & ~n1599;
  assign n1601 = reg_i_hlock0_out & ~n1600;
  assign n1602 = ~n68 & ~n269;
  assign n1603 = next_sys_fair<1>_out  & ~n1602;
  assign n1604 = ~n1045 & ~n1603;
  assign n1605 = reg_controllable_locked_out & ~n1604;
  assign n1606 = ~n810 & ~n1605;
  assign n1607 = next_sys_fair<0>_out  & ~n1606;
  assign n1608 = ~n1043 & ~n1057;
  assign n1609 = reg_controllable_locked_out & ~n1608;
  assign n1610 = ~n817 & ~n1609;
  assign n1611 = ~next_sys_fair<0>_out  & ~n1610;
  assign n1612 = ~n1607 & ~n1611;
  assign n1613 = reg_i_hbusreq0_out & ~n1612;
  assign n1614 = reg_i_hbusreq1_out & ~n1612;
  assign n1615 = ~n1190 & ~n1614;
  assign n1616 = ~reg_i_hbusreq0_out & ~n1615;
  assign n1617 = ~n1613 & ~n1616;
  assign n1618 = reg_controllable_nhgrant0_out & ~n1617;
  assign n1619 = ~n825 & ~n1618;
  assign n1620 = reg_controllable_hgrant1_out & ~n1619;
  assign n1621 = ~n853 & ~n1620;
  assign n1622 = reg_controllable_hmastlock_out & ~n1621;
  assign n1623 = ~n68 & ~n860;
  assign n1624 = next_sys_fair<1>_out  & ~n1623;
  assign n1625 = ~n645 & ~n1624;
  assign n1626 = reg_controllable_locked_out & ~n1625;
  assign n1627 = ~n870 & ~n1626;
  assign n1628 = next_sys_fair<0>_out  & ~n1627;
  assign n1629 = ~n878 & ~n1572;
  assign n1630 = ~next_sys_fair<0>_out  & ~n1629;
  assign n1631 = ~n1628 & ~n1630;
  assign n1632 = reg_i_hbusreq0_out & ~n1631;
  assign n1633 = reg_i_hbusreq1_out & ~n1631;
  assign n1634 = ~n896 & ~n1633;
  assign n1635 = ~reg_i_hbusreq0_out & ~n1634;
  assign n1636 = ~n1632 & ~n1635;
  assign n1637 = reg_controllable_nhgrant0_out & ~n1636;
  assign n1638 = ~n911 & ~n1637;
  assign n1639 = reg_controllable_hgrant1_out & ~n1638;
  assign n1640 = ~n934 & ~n1639;
  assign n1641 = ~reg_controllable_hmastlock_out & ~n1640;
  assign n1642 = ~n1622 & ~n1641;
  assign n1643 = ~reg_i_hlock0_out & ~n1642;
  assign n1644 = ~n1601 & ~n1643;
  assign n1645 = ~reg_stateG2_out & ~n1644;
  assign n1646 = ~n630 & ~n1645;
  assign n1647 = ~reg_controllable_hmaster0_out & ~n1646;
  assign n1648 = ~n1569 & ~n1647;
  assign n1649 = reg_i_hlock1_out & ~n1648;
  assign n1650 = reg_controllable_locked_out & ~n1381;
  assign n1651 = ~n1295 & ~n1650;
  assign n1652 = next_sys_fair<0>_out  & ~n1651;
  assign n1653 = ~n587 & ~n609;
  assign n1654 = reg_controllable_locked_out & ~n1653;
  assign n1655 = ~n1299 & ~n1654;
  assign n1656 = ~next_sys_fair<0>_out  & ~n1655;
  assign n1657 = ~n1652 & ~n1656;
  assign n1658 = reg_i_hbusreq0_out & ~n1657;
  assign n1659 = reg_i_hbusreq1_out & ~n1657;
  assign n1660 = reg_i_hbusreq1_out & ~n1659;
  assign n1661 = ~reg_i_hbusreq0_out & ~n1660;
  assign n1662 = ~n1658 & ~n1661;
  assign n1663 = reg_controllable_nhgrant0_out & ~n1662;
  assign n1664 = ~next_sys_fair<0>_out  & ~n1653;
  assign n1665 = ~n1396 & ~n1664;
  assign n1666 = reg_i_hbusreq0_out & ~n1665;
  assign n1667 = reg_i_hbusreq1_out & ~n1665;
  assign n1668 = reg_i_hbusreq1_out & ~n1667;
  assign n1669 = ~reg_i_hbusreq0_out & ~n1668;
  assign n1670 = ~n1666 & ~n1669;
  assign n1671 = ~reg_controllable_nhgrant0_out & ~n1670;
  assign n1672 = ~n1663 & ~n1671;
  assign n1673 = reg_controllable_hgrant1_out & ~n1672;
  assign n1674 = ~reg_controllable_hgrant1_out & ~n1670;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~reg_controllable_hmastlock_out & ~n1675;
  assign n1677 = ~reg_controllable_hmastlock_out & ~n1676;
  assign n1678 = reg_stateG2_out & ~n1677;
  assign n1679 = ~n500 & ~n829;
  assign n1680 = reg_controllable_locked_out & ~n1679;
  assign n1681 = ~n110 & ~n833;
  assign n1682 = ~reg_controllable_locked_out & ~n1681;
  assign n1683 = ~n1680 & ~n1682;
  assign n1684 = ~next_sys_fair<0>_out  & ~n1683;
  assign n1685 = ~n498 & ~n1684;
  assign n1686 = reg_i_hbusreq0_out & ~n1685;
  assign n1687 = reg_i_hbusreq1_out & ~n1685;
  assign n1688 = ~n1002 & ~n1687;
  assign n1689 = ~reg_i_hbusreq0_out & ~n1688;
  assign n1690 = ~n1686 & ~n1689;
  assign n1691 = reg_controllable_nhgrant0_out & ~n1690;
  assign n1692 = ~n520 & ~n804;
  assign n1693 = ~next_sys_fair<0>_out  & ~n1692;
  assign n1694 = ~n517 & ~n1693;
  assign n1695 = reg_i_hbusreq0_out & ~n1694;
  assign n1696 = reg_i_hbusreq1_out & ~n1694;
  assign n1697 = reg_i_hbusreq1_out & ~n1696;
  assign n1698 = ~reg_i_hbusreq0_out & ~n1697;
  assign n1699 = ~n1695 & ~n1698;
  assign n1700 = ~reg_controllable_nhgrant0_out & ~n1699;
  assign n1701 = ~n1691 & ~n1700;
  assign n1702 = reg_controllable_hgrant1_out & ~n1701;
  assign n1703 = reg_controllable_nhgrant0_out & ~n1699;
  assign n1704 = ~n1047 & ~n1074;
  assign n1705 = next_sys_fair<0>_out  & ~n1704;
  assign n1706 = ~n1057 & ~n1603;
  assign n1707 = reg_controllable_locked_out & ~n1706;
  assign n1708 = ~n110 & ~n808;
  assign n1709 = ~reg_controllable_locked_out & ~n1708;
  assign n1710 = ~n1707 & ~n1709;
  assign n1711 = ~next_sys_fair<0>_out  & ~n1710;
  assign n1712 = ~n1705 & ~n1711;
  assign n1713 = reg_i_hbusreq0_out & ~n1712;
  assign n1714 = reg_i_hbusreq1_out & ~n1712;
  assign n1715 = ~n421 & ~n1714;
  assign n1716 = ~reg_i_hbusreq0_out & ~n1715;
  assign n1717 = ~n1713 & ~n1716;
  assign n1718 = ~reg_controllable_nhgrant0_out & ~n1717;
  assign n1719 = ~n1703 & ~n1718;
  assign n1720 = ~reg_controllable_hgrant1_out & ~n1719;
  assign n1721 = ~n1702 & ~n1720;
  assign n1722 = reg_controllable_hmastlock_out & ~n1721;
  assign n1723 = ~n1331 & ~n1520;
  assign n1724 = next_sys_fair<0>_out  & ~n1723;
  assign n1725 = ~n862 & ~n1433;
  assign n1726 = reg_controllable_locked_out & ~n1725;
  assign n1727 = ~n915 & ~n1315;
  assign n1728 = ~reg_controllable_locked_out & ~n1727;
  assign n1729 = ~n1726 & ~n1728;
  assign n1730 = ~next_sys_fair<0>_out  & ~n1729;
  assign n1731 = ~n1724 & ~n1730;
  assign n1732 = reg_i_hbusreq0_out & ~n1731;
  assign n1733 = reg_i_hbusreq1_out & ~n1731;
  assign n1734 = ~n1025 & ~n1733;
  assign n1735 = ~reg_i_hbusreq0_out & ~n1734;
  assign n1736 = ~n1732 & ~n1735;
  assign n1737 = reg_controllable_nhgrant0_out & ~n1736;
  assign n1738 = ~next_sys_fair<0>_out  & ~n1725;
  assign n1739 = ~n1432 & ~n1738;
  assign n1740 = reg_i_hbusreq0_out & ~n1739;
  assign n1741 = reg_i_hbusreq1_out & ~n1739;
  assign n1742 = ~n1034 & ~n1741;
  assign n1743 = ~reg_i_hbusreq0_out & ~n1742;
  assign n1744 = ~n1740 & ~n1743;
  assign n1745 = ~reg_controllable_nhgrant0_out & ~n1744;
  assign n1746 = ~n1737 & ~n1745;
  assign n1747 = reg_controllable_hgrant1_out & ~n1746;
  assign n1748 = reg_controllable_nhgrant0_out & ~n1744;
  assign n1749 = ~n868 & ~n874;
  assign n1750 = ~reg_controllable_locked_out & ~n1749;
  assign n1751 = ~n1449 & ~n1750;
  assign n1752 = next_sys_fair<0>_out  & ~n1751;
  assign n1753 = ~n656 & ~n1624;
  assign n1754 = reg_controllable_locked_out & ~n1753;
  assign n1755 = ~n866 & ~n876;
  assign n1756 = ~reg_controllable_locked_out & ~n1755;
  assign n1757 = ~n1754 & ~n1756;
  assign n1758 = ~next_sys_fair<0>_out  & ~n1757;
  assign n1759 = ~n1752 & ~n1758;
  assign n1760 = reg_i_hbusreq0_out & ~n1759;
  assign n1761 = reg_i_hbusreq1_out & ~n1759;
  assign n1762 = ~n479 & ~n1761;
  assign n1763 = ~reg_i_hbusreq0_out & ~n1762;
  assign n1764 = ~n1760 & ~n1763;
  assign n1765 = ~reg_controllable_nhgrant0_out & ~n1764;
  assign n1766 = ~n1748 & ~n1765;
  assign n1767 = ~reg_controllable_hgrant1_out & ~n1766;
  assign n1768 = ~n1747 & ~n1767;
  assign n1769 = ~reg_controllable_hmastlock_out & ~n1768;
  assign n1770 = ~n1722 & ~n1769;
  assign n1771 = reg_i_hlock0_out & ~n1770;
  assign n1772 = ~n1226 & ~n1433;
  assign n1773 = reg_controllable_locked_out & ~n1772;
  assign n1774 = ~n1253 & ~n1315;
  assign n1775 = ~reg_controllable_locked_out & ~n1774;
  assign n1776 = ~n1773 & ~n1775;
  assign n1777 = ~next_sys_fair<0>_out  & ~n1776;
  assign n1778 = ~n1724 & ~n1777;
  assign n1779 = reg_i_hbusreq0_out & ~n1778;
  assign n1780 = reg_i_hbusreq1_out & ~n1778;
  assign n1781 = ~n1555 & ~n1780;
  assign n1782 = ~reg_i_hbusreq0_out & ~n1781;
  assign n1783 = ~n1779 & ~n1782;
  assign n1784 = reg_controllable_nhgrant0_out & ~n1783;
  assign n1785 = ~next_sys_fair<0>_out  & ~n1772;
  assign n1786 = ~n1432 & ~n1785;
  assign n1787 = reg_i_hbusreq0_out & ~n1786;
  assign n1788 = reg_i_hbusreq1_out & ~n1786;
  assign n1789 = ~n1512 & ~n1788;
  assign n1790 = ~reg_i_hbusreq0_out & ~n1789;
  assign n1791 = ~n1787 & ~n1790;
  assign n1792 = ~reg_controllable_nhgrant0_out & ~n1791;
  assign n1793 = ~n1784 & ~n1792;
  assign n1794 = reg_controllable_hgrant1_out & ~n1793;
  assign n1795 = reg_controllable_nhgrant0_out & ~n1791;
  assign n1796 = ~n1520 & ~n1750;
  assign n1797 = next_sys_fair<0>_out  & ~n1796;
  assign n1798 = ~n876 & ~n1230;
  assign n1799 = ~reg_controllable_locked_out & ~n1798;
  assign n1800 = ~n1773 & ~n1799;
  assign n1801 = ~next_sys_fair<0>_out  & ~n1800;
  assign n1802 = ~n1797 & ~n1801;
  assign n1803 = reg_i_hbusreq0_out & ~n1802;
  assign n1804 = reg_i_hbusreq1_out & ~n1802;
  assign n1805 = ~n547 & ~n1804;
  assign n1806 = ~reg_i_hbusreq0_out & ~n1805;
  assign n1807 = ~n1803 & ~n1806;
  assign n1808 = ~reg_controllable_nhgrant0_out & ~n1807;
  assign n1809 = ~n1795 & ~n1808;
  assign n1810 = ~reg_controllable_hgrant1_out & ~n1809;
  assign n1811 = ~n1794 & ~n1810;
  assign n1812 = ~reg_controllable_hmastlock_out & ~n1811;
  assign n1813 = ~n1087 & ~n1812;
  assign n1814 = ~reg_i_hlock0_out & ~n1813;
  assign n1815 = ~n1771 & ~n1814;
  assign n1816 = ~reg_stateG2_out & ~n1815;
  assign n1817 = ~n1678 & ~n1816;
  assign n1818 = reg_controllable_hmaster0_out & ~n1817;
  assign n1819 = ~n868 & ~n1494;
  assign n1820 = ~reg_controllable_locked_out & ~n1819;
  assign n1821 = ~n1134 & ~n1820;
  assign n1822 = next_sys_fair<0>_out  & ~n1821;
  assign n1823 = ~reg_controllable_locked_out & ~n875;
  assign n1824 = ~n276 & ~n1823;
  assign n1825 = ~next_sys_fair<0>_out  & ~n1824;
  assign n1826 = ~n1822 & ~n1825;
  assign n1827 = reg_i_hbusreq0_out & ~n1826;
  assign n1828 = reg_i_hbusreq1_out & ~n1826;
  assign n1829 = ~n718 & ~n1828;
  assign n1830 = ~reg_i_hbusreq0_out & ~n1829;
  assign n1831 = ~n1827 & ~n1830;
  assign n1832 = ~reg_controllable_nhgrant0_out & ~n1831;
  assign n1833 = ~n1131 & ~n1832;
  assign n1834 = ~reg_controllable_hgrant1_out & ~n1833;
  assign n1835 = ~n1130 & ~n1834;
  assign n1836 = reg_controllable_hmastlock_out & ~n1835;
  assign n1837 = ~n110 & ~n533;
  assign n1838 = ~reg_controllable_locked_out & ~n1837;
  assign n1839 = ~n813 & ~n1838;
  assign n1840 = ~next_sys_fair<0>_out  & ~n1839;
  assign n1841 = ~n1186 & ~n1840;
  assign n1842 = reg_i_hbusreq0_out & ~n1841;
  assign n1843 = reg_i_hbusreq1_out & ~n1841;
  assign n1844 = ~n752 & ~n1843;
  assign n1845 = ~reg_i_hbusreq0_out & ~n1844;
  assign n1846 = ~n1842 & ~n1845;
  assign n1847 = reg_controllable_nhgrant0_out & ~n1846;
  assign n1848 = ~n764 & ~n1198;
  assign n1849 = ~reg_i_hbusreq0_out & ~n1848;
  assign n1850 = ~n1197 & ~n1849;
  assign n1851 = ~reg_controllable_nhgrant0_out & ~n1850;
  assign n1852 = ~n1847 & ~n1851;
  assign n1853 = reg_controllable_hgrant1_out & ~n1852;
  assign n1854 = reg_controllable_nhgrant0_out & ~n1850;
  assign n1855 = ~n1045 & ~n1547;
  assign n1856 = reg_controllable_locked_out & ~n1855;
  assign n1857 = ~reg_controllable_locked_out & ~n1207;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = next_sys_fair<0>_out  & ~n1858;
  assign n1860 = reg_controllable_locked_out & ~n1056;
  assign n1861 = ~reg_controllable_locked_out & ~n87;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = ~next_sys_fair<0>_out  & ~n1862;
  assign n1864 = ~n1859 & ~n1863;
  assign n1865 = reg_i_hbusreq0_out & ~n1864;
  assign n1866 = reg_i_hbusreq1_out & ~n1864;
  assign n1867 = ~n792 & ~n1866;
  assign n1868 = ~reg_i_hbusreq0_out & ~n1867;
  assign n1869 = ~n1865 & ~n1868;
  assign n1870 = ~reg_controllable_nhgrant0_out & ~n1869;
  assign n1871 = ~n1854 & ~n1870;
  assign n1872 = ~reg_controllable_hgrant1_out & ~n1871;
  assign n1873 = ~n1853 & ~n1872;
  assign n1874 = ~reg_controllable_hmastlock_out & ~n1873;
  assign n1875 = ~n1836 & ~n1874;
  assign n1876 = reg_i_hlock0_out & ~n1875;
  assign n1877 = ~n1270 & ~n1876;
  assign n1878 = ~reg_stateG2_out & ~n1877;
  assign n1879 = ~n630 & ~n1878;
  assign n1880 = ~reg_controllable_hmaster0_out & ~n1879;
  assign n1881 = ~n1818 & ~n1880;
  assign n1882 = ~reg_i_hlock1_out & ~n1881;
  assign n1883 = ~n1649 & ~n1882;
  assign n1884 = ~reg_controllable_ndecide_out & ~n1883;
  assign n1885 = ~n1380 & ~n1884;
  assign n1886 = ~reg_stateG10_1_out & ~n1885;
  assign n1887 = ~n1280 & ~n1886;
  assign n1888 = ~next_sys_fair<2>_out  & ~n1887;
  assign n1889 = ~next_sys_fair<2>_out  & ~n1888;
  assign n1890 = ~env_safe_err_happened_out & n1889;
  assign n1891 = ~env_safe_err_happened_out & ~n1890;
  assign n1892 = n33 & ~n1891;
  assign n1893 = n33 & ~n1892;
  assign n1894 = ~i_hbusreq0 & i_hlock0;
  assign n1895 = ~i_hbusreq1 & i_hlock1;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = n33 & env_safe_err_happened_out;
  assign n1898 = n1896 & ~n1897;
  assign n1899 = n33 & next_sys_fair<2>_out ;
  assign n1900 = n33 & next_sys_fair<0>_out ;
  assign n1901 = n33 & next_sys_fair<1>_out ;
  assign n1902 = n1900 & n1901;
  assign n1903 = ~n1899 & n1902;
  assign n1904 = i_hbusreq1 & ~controllable_hmaster0;
  assign n1905 = n1903 & ~n1904;
  assign n1906 = n33 & reg_stateG2_out;
  assign n1907 = ~n1900 & ~n1901;
  assign n1908 = ~n1899 & n1907;
  assign n1909 = ~n1906 & n1908;
  assign n1910 = ~n1900 & n1901;
  assign n1911 = ~n1899 & n1910;
  assign n1912 = i_hbusreq0 & controllable_hmaster0;
  assign n1913 = n1911 & ~n1912;
  assign n1914 = n33 & reg_stateG3_0_out;
  assign n1915 = n33 & reg_stateG3_1_out;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n33 & reg_stateG3_2_out;
  assign n1918 = n1916 & ~n1917;
  assign n1919 = n1900 & ~n1901;
  assign n1920 = ~n1899 & n1919;
  assign n1921 = n1918 & n1920;
  assign n1922 = ~n1913 & ~n1921;
  assign n1923 = ~n1909 & n1922;
  assign n1924 = ~n1905 & n1923;
  assign n1925 = n33 & next_env_fair_out;
  assign n1926 = i_hready & n1925;
  assign n1927 = n33 & fair_cnt<0>_out ;
  assign n1928 = n33 & fair_cnt<1>_out ;
  assign n1929 = n1927 & n1928;
  assign n1930 = n1926 & n1929;
  assign n1931 = n33 & fair_cnt<2>_out ;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = n1930 & n1931;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1924 & n1934;
  assign n1936 = n1926 & n1927;
  assign n1937 = ~n1928 & ~n1936;
  assign n1938 = ~n1930 & ~n1937;
  assign n1939 = n1924 & n1938;
  assign n1940 = ~n1926 & ~n1927;
  assign n1941 = ~n1936 & ~n1940;
  assign n1942 = n1924 & n1941;
  assign n1943 = n1901 & n1924;
  assign n1944 = n1922 & ~n1943;
  assign n1945 = n1900 & n1924;
  assign n1946 = ~n1909 & ~n1913;
  assign n1947 = ~n1945 & n1946;
  assign n1948 = n33 & reg_stateA1_out;
  assign n1949 = controllable_hmastlock & ~n1948;
  assign n1950 = ~i_hburst1 & ~i_hburst0;
  assign n1951 = n1949 & n1950;
  assign n1952 = controllable_busreq & n1948;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = n33 & reg_stateG10_1_out;
  assign n1955 = controllable_hgrant1 & ~n1954;
  assign n1956 = ~i_hbusreq1 & ~n1955;
  assign n1957 = controllable_busreq & n1906;
  assign n1958 = controllable_hmastlock & ~controllable_nstart;
  assign n1959 = ~i_hburst0 & n1958;
  assign n1960 = ~i_hburst1 & ~n1906;
  assign n1961 = n1959 & n1960;
  assign n1962 = ~n1957 & ~n1961;
  assign n1963 = n1918 & n1959;
  assign n1964 = i_hburst1 & n1963;
  assign n1965 = i_hready & n1964;
  assign n1966 = n1914 & n1915;
  assign n1967 = ~n1917 & n1966;
  assign n1968 = i_hready & n1967;
  assign n1969 = n1915 & ~n1968;
  assign n1970 = i_hready & ~n1917;
  assign n1971 = n1914 & ~n1915;
  assign n1972 = n1970 & n1971;
  assign n1973 = ~n1969 & ~n1972;
  assign n1974 = ~n1965 & n1973;
  assign n1975 = ~i_hready & n1964;
  assign n1976 = ~n1914 & ~n1970;
  assign n1977 = n1914 & n1970;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1916 & n1978;
  assign n1980 = ~n1975 & ~n1979;
  assign n1981 = i_hready & ~controllable_hmastlock;
  assign n1982 = ~controllable_hmastlock & ~n1981;
  assign n1983 = controllable_locked & ~n1982;
  assign n1984 = controllable_hmastlock & ~controllable_locked;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = controllable_nhgrant0 & ~n1985;
  assign n1987 = ~controllable_nhgrant0 & ~n1982;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = controllable_hgrant1 & ~n1988;
  assign n1990 = ~controllable_hgrant1 & ~n1982;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = ~i_hlock1 & ~n1991;
  assign n1993 = ~i_hlock1 & ~n1992;
  assign n1994 = ~controllable_ndecide & ~n1993;
  assign n1995 = ~controllable_ndecide & ~n1994;
  assign n1996 = controllable_hmaster0 & ~n1995;
  assign n1997 = controllable_hmaster0 & ~n1996;
  assign n1998 = i_hlock0 & ~n1997;
  assign n1999 = controllable_hmastlock & controllable_locked;
  assign n2000 = i_hready & controllable_hmastlock;
  assign n2001 = controllable_hmastlock & ~n2000;
  assign n2002 = ~controllable_locked & n2001;
  assign n2003 = ~n1999 & ~n2002;
  assign n2004 = controllable_nhgrant0 & ~n2003;
  assign n2005 = ~controllable_nhgrant0 & n2001;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = controllable_hgrant1 & ~n2006;
  assign n2008 = ~controllable_hgrant1 & n2001;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = i_hlock1 & ~n2009;
  assign n2011 = ~i_hlock1 & n1991;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~controllable_ndecide & n2012;
  assign n2014 = ~controllable_ndecide & ~n2013;
  assign n2015 = controllable_hmaster0 & ~n2014;
  assign n2016 = controllable_hmaster0 & ~n2015;
  assign n2017 = ~i_hlock0 & ~n2016;
  assign n2018 = ~n1998 & ~n2017;
  assign n2019 = i_hbusreq0 & ~n2018;
  assign n2020 = i_hbusreq1 & ~n1995;
  assign n2021 = i_hbusreq1 & ~n2020;
  assign n2022 = controllable_hmaster0 & ~n2021;
  assign n2023 = controllable_hmaster0 & ~n2022;
  assign n2024 = i_hlock0 & ~n2023;
  assign n2025 = i_hbusreq1 & ~n2014;
  assign n2026 = i_hbusreq1 & ~n2025;
  assign n2027 = controllable_hmaster0 & ~n2026;
  assign n2028 = controllable_hmaster0 & ~n2027;
  assign n2029 = ~i_hlock0 & ~n2028;
  assign n2030 = ~n2024 & ~n2029;
  assign n2031 = ~i_hbusreq0 & ~n2030;
  assign n2032 = ~n2019 & ~n2031;
  assign n2033 = ~n1899 & ~n2032;
  assign n2034 = ~n1899 & ~n2033;
  assign n2035 = n1980 & ~n2034;
  assign n2036 = n1980 & ~n2035;
  assign n2037 = n1974 & ~n2036;
  assign n2038 = n1974 & ~n2037;
  assign n2039 = ~n1962 & ~n2038;
  assign n2040 = i_hready & n1916;
  assign n2041 = n1917 & ~n2040;
  assign n2042 = ~n1968 & ~n2041;
  assign n2043 = i_hready & ~controllable_locked;
  assign n2044 = ~controllable_locked & ~n2043;
  assign n2045 = ~controllable_nhgrant0 & ~n2044;
  assign n2046 = ~controllable_nhgrant0 & ~n2045;
  assign n2047 = ~controllable_hgrant1 & ~n2046;
  assign n2048 = ~controllable_hgrant1 & ~n2047;
  assign n2049 = controllable_ndecide & ~n2048;
  assign n2050 = ~n1994 & ~n2049;
  assign n2051 = controllable_hmaster0 & ~n2050;
  assign n2052 = controllable_hmaster0 & ~n2051;
  assign n2053 = i_hlock0 & ~n2052;
  assign n2054 = ~i_hready & ~controllable_hmastlock;
  assign n2055 = ~controllable_hmastlock & ~n2054;
  assign n2056 = controllable_locked & ~n2055;
  assign n2057 = ~controllable_locked & ~n2000;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = controllable_nhgrant0 & ~n2058;
  assign n2060 = ~i_hready & ~controllable_nhgrant0;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = controllable_hgrant1 & ~n2061;
  assign n2063 = ~i_hready & ~controllable_hgrant1;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~controllable_ndecide & n2064;
  assign n2066 = ~n2049 & ~n2065;
  assign n2067 = controllable_hmaster0 & ~n2066;
  assign n2068 = controllable_hmaster0 & ~n2067;
  assign n2069 = ~i_hlock0 & ~n2068;
  assign n2070 = ~n2053 & ~n2069;
  assign n2071 = i_hbusreq0 & ~n2070;
  assign n2072 = i_hbusreq1 & ~n2050;
  assign n2073 = controllable_ndecide & ~n2049;
  assign n2074 = ~i_hbusreq1 & ~n2073;
  assign n2075 = ~n2072 & ~n2074;
  assign n2076 = controllable_hmaster0 & ~n2075;
  assign n2077 = controllable_hmaster0 & ~n2076;
  assign n2078 = i_hlock0 & ~n2077;
  assign n2079 = ~n2069 & ~n2078;
  assign n2080 = ~i_hbusreq0 & ~n2079;
  assign n2081 = ~n2071 & ~n2080;
  assign n2082 = ~n1899 & ~n2081;
  assign n2083 = ~n1899 & ~n2082;
  assign n2084 = n1980 & ~n2083;
  assign n2085 = n1980 & ~n2084;
  assign n2086 = n1974 & ~n2085;
  assign n2087 = n1974 & ~n2086;
  assign n2088 = ~n2042 & ~n2087;
  assign n2089 = ~n1983 & ~n2002;
  assign n2090 = controllable_nhgrant0 & ~n2089;
  assign n2091 = ~n1987 & ~n2090;
  assign n2092 = controllable_hgrant1 & ~n2091;
  assign n2093 = ~n1990 & ~n2092;
  assign n2094 = ~i_hlock1 & ~n2093;
  assign n2095 = ~i_hlock1 & ~n2094;
  assign n2096 = ~controllable_ndecide & ~n2095;
  assign n2097 = ~n2049 & ~n2096;
  assign n2098 = controllable_hmaster0 & ~n2097;
  assign n2099 = ~i_hready & ~controllable_locked;
  assign n2100 = ~controllable_locked & ~n2099;
  assign n2101 = controllable_nhgrant0 & ~n2100;
  assign n2102 = controllable_nhgrant0 & ~n2101;
  assign n2103 = controllable_hgrant1 & ~n2102;
  assign n2104 = controllable_hgrant1 & ~n2103;
  assign n2105 = ~i_hlock1 & ~n2104;
  assign n2106 = ~i_hlock1 & ~n2105;
  assign n2107 = ~controllable_ndecide & ~n2106;
  assign n2108 = ~controllable_ndecide & ~n2107;
  assign n2109 = ~controllable_hmaster0 & ~n2108;
  assign n2110 = ~n2098 & ~n2109;
  assign n2111 = i_hlock0 & ~n2110;
  assign n2112 = controllable_locked & ~n2056;
  assign n2113 = controllable_nhgrant0 & ~n2112;
  assign n2114 = ~n2060 & ~n2113;
  assign n2115 = controllable_hgrant1 & ~n2114;
  assign n2116 = ~n2063 & ~n2115;
  assign n2117 = ~controllable_ndecide & n2116;
  assign n2118 = ~n2049 & ~n2117;
  assign n2119 = controllable_hmaster0 & ~n2118;
  assign n2120 = ~controllable_ndecide & ~n2104;
  assign n2121 = ~controllable_ndecide & ~n2120;
  assign n2122 = ~controllable_hmaster0 & ~n2121;
  assign n2123 = ~n2119 & ~n2122;
  assign n2124 = ~i_hlock0 & ~n2123;
  assign n2125 = ~n2111 & ~n2124;
  assign n2126 = i_hbusreq0 & ~n2125;
  assign n2127 = i_hbusreq1 & ~n2097;
  assign n2128 = ~n2074 & ~n2127;
  assign n2129 = controllable_hmaster0 & ~n2128;
  assign n2130 = i_hbusreq1 & ~n2108;
  assign n2131 = i_hbusreq1 & ~n2130;
  assign n2132 = ~controllable_hmaster0 & ~n2131;
  assign n2133 = ~n2129 & ~n2132;
  assign n2134 = i_hlock0 & ~n2133;
  assign n2135 = ~n2124 & ~n2134;
  assign n2136 = ~i_hbusreq0 & ~n2135;
  assign n2137 = ~n2126 & ~n2136;
  assign n2138 = ~n1899 & ~n2137;
  assign n2139 = ~n1899 & ~n2138;
  assign n2140 = n1980 & ~n2139;
  assign n2141 = n1980 & ~n2140;
  assign n2142 = n1974 & ~n2141;
  assign n2143 = n1974 & ~n2142;
  assign n2144 = n2042 & ~n2143;
  assign n2145 = ~n2088 & ~n2144;
  assign n2146 = n1962 & ~n2145;
  assign n2147 = ~n2039 & ~n2146;
  assign n2148 = n1956 & ~n2147;
  assign n2149 = ~controllable_hmastlock & ~controllable_locked;
  assign n2150 = ~n1999 & ~n2149;
  assign n2151 = controllable_nhgrant0 & ~n2150;
  assign n2152 = controllable_hgrant1 & n2151;
  assign n2153 = controllable_ndecide & n2152;
  assign n2154 = ~controllable_ndecide & ~n2012;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = controllable_hmaster0 & ~n2155;
  assign n2157 = i_hbusreq0 & n2156;
  assign n2158 = i_hbusreq1 & ~n2155;
  assign n2159 = ~i_hbusreq1 & n2153;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = controllable_hmaster0 & ~n2160;
  assign n2162 = ~i_hbusreq0 & n2161;
  assign n2163 = ~n2157 & ~n2162;
  assign n2164 = ~n1899 & n2163;
  assign n2165 = ~n1899 & ~n2164;
  assign n2166 = n1980 & ~n2165;
  assign n2167 = n1980 & ~n2166;
  assign n2168 = n1974 & ~n2167;
  assign n2169 = n1974 & ~n2168;
  assign n2170 = ~n2042 & ~n2169;
  assign n2171 = n2042 & ~n2165;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n1962 & ~n2172;
  assign n2174 = ~n1999 & ~n2057;
  assign n2175 = controllable_nhgrant0 & ~n2174;
  assign n2176 = controllable_hgrant1 & n2175;
  assign n2177 = ~controllable_hgrant1 & n2046;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = controllable_ndecide & ~n2178;
  assign n2180 = ~i_hlock1 & ~n2064;
  assign n2181 = ~n2010 & ~n2180;
  assign n2182 = ~controllable_ndecide & ~n2181;
  assign n2183 = ~n2179 & ~n2182;
  assign n2184 = controllable_hmaster0 & ~n2183;
  assign n2185 = i_hlock0 & n2184;
  assign n2186 = ~controllable_ndecide & ~n2064;
  assign n2187 = ~n2179 & ~n2186;
  assign n2188 = controllable_hmaster0 & ~n2187;
  assign n2189 = ~i_hlock0 & n2188;
  assign n2190 = ~n2185 & ~n2189;
  assign n2191 = i_hbusreq0 & ~n2190;
  assign n2192 = i_hbusreq1 & ~n2183;
  assign n2193 = ~i_hbusreq1 & n2179;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = controllable_hmaster0 & ~n2194;
  assign n2196 = i_hlock0 & n2195;
  assign n2197 = ~n2189 & ~n2196;
  assign n2198 = ~i_hbusreq0 & ~n2197;
  assign n2199 = ~n2191 & ~n2198;
  assign n2200 = ~n1899 & n2199;
  assign n2201 = ~n1899 & ~n2200;
  assign n2202 = n1980 & ~n2201;
  assign n2203 = n1980 & ~n2202;
  assign n2204 = n1974 & ~n2203;
  assign n2205 = n1974 & ~n2204;
  assign n2206 = ~n2042 & ~n2205;
  assign n2207 = ~n1974 & ~n2165;
  assign n2208 = ~n1980 & ~n2165;
  assign n2209 = controllable_locked & ~n1999;
  assign n2210 = controllable_nhgrant0 & ~n2209;
  assign n2211 = controllable_hgrant1 & n2210;
  assign n2212 = ~n2177 & ~n2211;
  assign n2213 = controllable_ndecide & ~n2212;
  assign n2214 = ~i_hlock1 & ~n2116;
  assign n2215 = ~n2010 & ~n2214;
  assign n2216 = ~controllable_ndecide & ~n2215;
  assign n2217 = ~n2213 & ~n2216;
  assign n2218 = controllable_hmaster0 & ~n2217;
  assign n2219 = controllable_ndecide & ~n2104;
  assign n2220 = ~n2107 & ~n2219;
  assign n2221 = ~controllable_hmaster0 & n2220;
  assign n2222 = ~n2218 & ~n2221;
  assign n2223 = i_hlock0 & ~n2222;
  assign n2224 = ~controllable_ndecide & ~n2116;
  assign n2225 = ~n2213 & ~n2224;
  assign n2226 = controllable_hmaster0 & ~n2225;
  assign n2227 = ~controllable_hmaster0 & n2104;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = ~i_hlock0 & ~n2228;
  assign n2230 = ~n2223 & ~n2229;
  assign n2231 = i_hbusreq0 & ~n2230;
  assign n2232 = i_hbusreq1 & ~n2217;
  assign n2233 = ~i_hbusreq1 & n2213;
  assign n2234 = ~n2232 & ~n2233;
  assign n2235 = controllable_hmaster0 & ~n2234;
  assign n2236 = i_hbusreq1 & ~n2220;
  assign n2237 = controllable_ndecide & ~n2219;
  assign n2238 = ~i_hbusreq1 & ~n2237;
  assign n2239 = ~n2236 & ~n2238;
  assign n2240 = ~controllable_hmaster0 & n2239;
  assign n2241 = ~n2235 & ~n2240;
  assign n2242 = i_hlock0 & ~n2241;
  assign n2243 = ~n2229 & ~n2242;
  assign n2244 = ~i_hbusreq0 & ~n2243;
  assign n2245 = ~n2231 & ~n2244;
  assign n2246 = ~n1899 & n2245;
  assign n2247 = ~n1899 & ~n2246;
  assign n2248 = n1980 & ~n2247;
  assign n2249 = ~n2208 & ~n2248;
  assign n2250 = n1974 & ~n2249;
  assign n2251 = ~n2207 & ~n2250;
  assign n2252 = n2042 & ~n2251;
  assign n2253 = ~n2206 & ~n2252;
  assign n2254 = n1962 & ~n2253;
  assign n2255 = ~n2173 & ~n2254;
  assign n2256 = ~n1956 & ~n2255;
  assign n2257 = ~n2148 & ~n2256;
  assign n2258 = ~n1953 & ~n2257;
  assign n2259 = ~n1983 & ~n2043;
  assign n2260 = ~controllable_nhgrant0 & ~n2259;
  assign n2261 = ~controllable_nhgrant0 & ~n2260;
  assign n2262 = ~controllable_hgrant1 & ~n2261;
  assign n2263 = ~controllable_hgrant1 & ~n2262;
  assign n2264 = controllable_ndecide & ~n2263;
  assign n2265 = ~controllable_ndecide & ~n1991;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = controllable_hmaster0 & ~n2266;
  assign n2268 = controllable_hmaster0 & ~n2267;
  assign n2269 = i_hlock0 & ~n2268;
  assign n2270 = ~n2065 & ~n2264;
  assign n2271 = controllable_hmaster0 & ~n2270;
  assign n2272 = controllable_hmaster0 & ~n2271;
  assign n2273 = ~i_hlock0 & ~n2272;
  assign n2274 = ~n2269 & ~n2273;
  assign n2275 = ~n1899 & ~n2274;
  assign n2276 = ~n1899 & ~n2275;
  assign n2277 = n1980 & ~n2276;
  assign n2278 = n1980 & ~n2277;
  assign n2279 = n1974 & ~n2278;
  assign n2280 = n1974 & ~n2279;
  assign n2281 = ~n2042 & ~n2280;
  assign n2282 = ~controllable_ndecide & ~n2093;
  assign n2283 = ~n2264 & ~n2282;
  assign n2284 = controllable_hmaster0 & ~n2283;
  assign n2285 = ~n2122 & ~n2284;
  assign n2286 = i_hlock0 & ~n2285;
  assign n2287 = ~n2117 & ~n2264;
  assign n2288 = controllable_hmaster0 & ~n2287;
  assign n2289 = ~n2122 & ~n2288;
  assign n2290 = ~i_hlock0 & ~n2289;
  assign n2291 = ~n2286 & ~n2290;
  assign n2292 = ~n1899 & ~n2291;
  assign n2293 = ~n1899 & ~n2292;
  assign n2294 = n1980 & ~n2293;
  assign n2295 = n1980 & ~n2294;
  assign n2296 = n1974 & ~n2295;
  assign n2297 = n1974 & ~n2296;
  assign n2298 = n2042 & ~n2297;
  assign n2299 = ~n2281 & ~n2298;
  assign n2300 = n1962 & ~n2299;
  assign n2301 = n1962 & ~n2300;
  assign n2302 = n1956 & ~n2301;
  assign n2303 = controllable_hgrant1 & n2059;
  assign n2304 = ~controllable_hgrant1 & n2261;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = controllable_ndecide & ~n2305;
  assign n2307 = ~n2186 & ~n2306;
  assign n2308 = controllable_hmaster0 & ~n2307;
  assign n2309 = i_hbusreq0 & n2308;
  assign n2310 = i_hbusreq1 & ~n2307;
  assign n2311 = ~controllable_ndecide & n1991;
  assign n2312 = ~n2306 & ~n2311;
  assign n2313 = ~i_hbusreq1 & ~n2312;
  assign n2314 = ~n2310 & ~n2313;
  assign n2315 = controllable_hmaster0 & ~n2314;
  assign n2316 = i_hlock0 & n2315;
  assign n2317 = ~i_hlock0 & n2308;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = ~i_hbusreq0 & ~n2318;
  assign n2320 = ~n2309 & ~n2319;
  assign n2321 = ~n1899 & n2320;
  assign n2322 = ~n1899 & ~n2321;
  assign n2323 = n1980 & ~n2322;
  assign n2324 = n1980 & ~n2323;
  assign n2325 = n1974 & ~n2324;
  assign n2326 = n1974 & ~n2325;
  assign n2327 = ~n2042 & ~n2326;
  assign n2328 = controllable_hgrant1 & controllable_nhgrant0;
  assign n2329 = ~n2304 & ~n2328;
  assign n2330 = controllable_ndecide & ~n2329;
  assign n2331 = ~controllable_nhgrant0 & ~n2060;
  assign n2332 = controllable_hgrant1 & ~n2331;
  assign n2333 = ~n2063 & ~n2332;
  assign n2334 = i_hlock1 & ~n2333;
  assign n2335 = ~n2214 & ~n2334;
  assign n2336 = ~controllable_ndecide & ~n2335;
  assign n2337 = ~n2330 & ~n2336;
  assign n2338 = controllable_hmaster0 & ~n2337;
  assign n2339 = i_hready & controllable_nhgrant0;
  assign n2340 = controllable_hgrant1 & n2339;
  assign n2341 = controllable_ndecide & n2340;
  assign n2342 = i_hlock1 & n2340;
  assign n2343 = ~i_hlock1 & n2104;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~controllable_ndecide & ~n2344;
  assign n2346 = ~n2341 & ~n2345;
  assign n2347 = ~controllable_hmaster0 & ~n2346;
  assign n2348 = ~n2338 & ~n2347;
  assign n2349 = i_hbusreq0 & ~n2348;
  assign n2350 = i_hbusreq1 & ~n2337;
  assign n2351 = ~controllable_ndecide & n2093;
  assign n2352 = ~n2330 & ~n2351;
  assign n2353 = ~i_hbusreq1 & ~n2352;
  assign n2354 = ~n2350 & ~n2353;
  assign n2355 = controllable_hmaster0 & ~n2354;
  assign n2356 = i_hbusreq1 & ~n2346;
  assign n2357 = ~controllable_ndecide & n2104;
  assign n2358 = ~n2341 & ~n2357;
  assign n2359 = ~i_hbusreq1 & ~n2358;
  assign n2360 = ~n2356 & ~n2359;
  assign n2361 = ~controllable_hmaster0 & ~n2360;
  assign n2362 = ~n2355 & ~n2361;
  assign n2363 = i_hlock0 & ~n2362;
  assign n2364 = ~n2224 & ~n2330;
  assign n2365 = ~i_hbusreq1 & ~n2364;
  assign n2366 = ~n2350 & ~n2365;
  assign n2367 = controllable_hmaster0 & ~n2366;
  assign n2368 = ~n2361 & ~n2367;
  assign n2369 = ~i_hlock0 & ~n2368;
  assign n2370 = ~n2363 & ~n2369;
  assign n2371 = ~i_hbusreq0 & ~n2370;
  assign n2372 = ~n2349 & ~n2371;
  assign n2373 = ~n1899 & n2372;
  assign n2374 = ~n1899 & ~n2373;
  assign n2375 = n1980 & ~n2374;
  assign n2376 = ~n2208 & ~n2375;
  assign n2377 = n1974 & ~n2376;
  assign n2378 = ~n2207 & ~n2377;
  assign n2379 = n2042 & ~n2378;
  assign n2380 = ~n2327 & ~n2379;
  assign n2381 = n1962 & ~n2380;
  assign n2382 = n1962 & ~n2381;
  assign n2383 = ~n1956 & ~n2382;
  assign n2384 = ~n2302 & ~n2383;
  assign n2385 = n1953 & ~n2384;
  assign n2386 = ~n2258 & ~n2385;
  assign n2387 = ~n1947 & ~n2386;
  assign n2388 = ~controllable_nhgrant0 & n2150;
  assign n2389 = ~controllable_nhgrant0 & ~n2388;
  assign n2390 = ~controllable_hgrant1 & ~n2389;
  assign n2391 = ~controllable_hgrant1 & ~n2390;
  assign n2392 = controllable_ndecide & ~n2391;
  assign n2393 = controllable_hgrant1 & ~n2001;
  assign n2394 = controllable_nhgrant0 & ~n2001;
  assign n2395 = ~controllable_nhgrant0 & n2003;
  assign n2396 = ~n2394 & ~n2395;
  assign n2397 = ~controllable_hgrant1 & ~n2396;
  assign n2398 = ~n2393 & ~n2397;
  assign n2399 = ~controllable_ndecide & ~n2398;
  assign n2400 = ~n2392 & ~n2399;
  assign n2401 = ~controllable_hmaster0 & ~n2400;
  assign n2402 = ~controllable_hmaster0 & ~n2401;
  assign n2403 = i_hlock0 & ~n2402;
  assign n2404 = controllable_hgrant1 & ~n1982;
  assign n2405 = controllable_nhgrant0 & ~n1982;
  assign n2406 = ~controllable_nhgrant0 & ~n1985;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = ~controllable_hgrant1 & ~n2407;
  assign n2409 = ~n2404 & ~n2408;
  assign n2410 = ~controllable_ndecide & ~n2409;
  assign n2411 = ~n2392 & ~n2410;
  assign n2412 = ~controllable_hmaster0 & ~n2411;
  assign n2413 = ~controllable_hmaster0 & ~n2412;
  assign n2414 = ~i_hlock0 & ~n2413;
  assign n2415 = ~n2403 & ~n2414;
  assign n2416 = ~n1899 & ~n2415;
  assign n2417 = ~n1899 & ~n2416;
  assign n2418 = n1980 & ~n2417;
  assign n2419 = n1980 & ~n2418;
  assign n2420 = n1974 & ~n2419;
  assign n2421 = n1974 & ~n2420;
  assign n2422 = ~n2042 & ~n2421;
  assign n2423 = n2042 & ~n2417;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n1962 & ~n2424;
  assign n2426 = ~controllable_nhgrant0 & n2174;
  assign n2427 = ~controllable_nhgrant0 & ~n2426;
  assign n2428 = ~controllable_hgrant1 & ~n2427;
  assign n2429 = ~controllable_hgrant1 & ~n2428;
  assign n2430 = controllable_ndecide & ~n2429;
  assign n2431 = ~n2399 & ~n2430;
  assign n2432 = ~controllable_hmaster0 & ~n2431;
  assign n2433 = ~controllable_hmaster0 & ~n2432;
  assign n2434 = i_hlock0 & ~n2433;
  assign n2435 = i_hready & controllable_hgrant1;
  assign n2436 = ~controllable_nhgrant0 & n2058;
  assign n2437 = ~n2339 & ~n2436;
  assign n2438 = ~controllable_hgrant1 & ~n2437;
  assign n2439 = ~n2435 & ~n2438;
  assign n2440 = ~controllable_ndecide & ~n2439;
  assign n2441 = ~n2430 & ~n2440;
  assign n2442 = ~controllable_hmaster0 & ~n2441;
  assign n2443 = ~controllable_hmaster0 & ~n2442;
  assign n2444 = ~i_hlock0 & ~n2443;
  assign n2445 = ~n2434 & ~n2444;
  assign n2446 = ~n1899 & ~n2445;
  assign n2447 = ~n1899 & ~n2446;
  assign n2448 = n1980 & ~n2447;
  assign n2449 = n1980 & ~n2448;
  assign n2450 = n1974 & ~n2449;
  assign n2451 = n1974 & ~n2450;
  assign n2452 = ~n2042 & ~n2451;
  assign n2453 = ~n1974 & ~n2417;
  assign n2454 = ~n1980 & ~n2417;
  assign n2455 = ~controllable_nhgrant0 & ~n2100;
  assign n2456 = ~controllable_nhgrant0 & ~n2455;
  assign n2457 = ~controllable_hgrant1 & ~n2456;
  assign n2458 = ~controllable_hgrant1 & ~n2457;
  assign n2459 = controllable_ndecide & ~n2458;
  assign n2460 = controllable_ndecide & ~n2459;
  assign n2461 = controllable_hmaster0 & ~n2460;
  assign n2462 = ~controllable_nhgrant0 & n2209;
  assign n2463 = ~controllable_nhgrant0 & ~n2462;
  assign n2464 = ~controllable_hgrant1 & ~n2463;
  assign n2465 = ~controllable_hgrant1 & ~n2464;
  assign n2466 = controllable_ndecide & ~n2465;
  assign n2467 = ~n2399 & ~n2466;
  assign n2468 = ~controllable_hmaster0 & ~n2467;
  assign n2469 = ~n2461 & ~n2468;
  assign n2470 = i_hlock0 & ~n2469;
  assign n2471 = controllable_hmaster0 & ~n2458;
  assign n2472 = ~controllable_nhgrant0 & n2112;
  assign n2473 = ~n2339 & ~n2472;
  assign n2474 = ~controllable_hgrant1 & ~n2473;
  assign n2475 = ~n2435 & ~n2474;
  assign n2476 = ~controllable_ndecide & ~n2475;
  assign n2477 = ~n2466 & ~n2476;
  assign n2478 = ~controllable_hmaster0 & ~n2477;
  assign n2479 = ~n2471 & ~n2478;
  assign n2480 = ~i_hlock0 & ~n2479;
  assign n2481 = ~n2470 & ~n2480;
  assign n2482 = ~n1899 & ~n2481;
  assign n2483 = ~n1899 & ~n2482;
  assign n2484 = n1980 & ~n2483;
  assign n2485 = ~n2454 & ~n2484;
  assign n2486 = n1974 & ~n2485;
  assign n2487 = ~n2453 & ~n2486;
  assign n2488 = n2042 & ~n2487;
  assign n2489 = ~n2452 & ~n2488;
  assign n2490 = n1962 & ~n2489;
  assign n2491 = ~n2425 & ~n2490;
  assign n2492 = n1956 & ~n2491;
  assign n2493 = controllable_nhgrant0 & ~n2044;
  assign n2494 = controllable_nhgrant0 & ~n2493;
  assign n2495 = controllable_hgrant1 & ~n2494;
  assign n2496 = ~n2428 & ~n2495;
  assign n2497 = controllable_ndecide & ~n2496;
  assign n2498 = i_hlock1 & ~n2398;
  assign n2499 = ~i_hlock1 & ~n2439;
  assign n2500 = ~n2498 & ~n2499;
  assign n2501 = ~controllable_ndecide & ~n2500;
  assign n2502 = ~n2497 & ~n2501;
  assign n2503 = ~controllable_hmaster0 & ~n2502;
  assign n2504 = ~controllable_hmaster0 & ~n2503;
  assign n2505 = i_hlock0 & ~n2504;
  assign n2506 = ~n2440 & ~n2497;
  assign n2507 = ~controllable_hmaster0 & ~n2506;
  assign n2508 = ~controllable_hmaster0 & ~n2507;
  assign n2509 = ~i_hlock0 & ~n2508;
  assign n2510 = ~n2505 & ~n2509;
  assign n2511 = i_hbusreq0 & ~n2510;
  assign n2512 = i_hbusreq1 & ~n2502;
  assign n2513 = ~n2399 & ~n2497;
  assign n2514 = ~i_hbusreq1 & ~n2513;
  assign n2515 = ~n2512 & ~n2514;
  assign n2516 = ~controllable_hmaster0 & ~n2515;
  assign n2517 = ~controllable_hmaster0 & ~n2516;
  assign n2518 = i_hlock0 & ~n2517;
  assign n2519 = ~n2509 & ~n2518;
  assign n2520 = ~i_hbusreq0 & ~n2519;
  assign n2521 = ~n2511 & ~n2520;
  assign n2522 = ~n1899 & ~n2521;
  assign n2523 = ~n1899 & ~n2522;
  assign n2524 = n1980 & ~n2523;
  assign n2525 = n1980 & ~n2524;
  assign n2526 = n1974 & ~n2525;
  assign n2527 = n1974 & ~n2526;
  assign n2528 = ~n2042 & ~n2527;
  assign n2529 = ~i_hlock1 & ~n2458;
  assign n2530 = ~i_hlock1 & ~n2529;
  assign n2531 = ~controllable_ndecide & ~n2530;
  assign n2532 = ~n2459 & ~n2531;
  assign n2533 = controllable_hmaster0 & ~n2532;
  assign n2534 = ~n2464 & ~n2495;
  assign n2535 = controllable_ndecide & ~n2534;
  assign n2536 = ~i_hlock1 & ~n2475;
  assign n2537 = ~n2498 & ~n2536;
  assign n2538 = ~controllable_ndecide & ~n2537;
  assign n2539 = ~n2535 & ~n2538;
  assign n2540 = ~controllable_hmaster0 & ~n2539;
  assign n2541 = ~n2533 & ~n2540;
  assign n2542 = i_hlock0 & ~n2541;
  assign n2543 = ~n2476 & ~n2535;
  assign n2544 = ~controllable_hmaster0 & ~n2543;
  assign n2545 = ~n2471 & ~n2544;
  assign n2546 = ~i_hlock0 & ~n2545;
  assign n2547 = ~n2542 & ~n2546;
  assign n2548 = i_hbusreq0 & ~n2547;
  assign n2549 = i_hbusreq1 & ~n2532;
  assign n2550 = ~i_hbusreq1 & ~n2460;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = controllable_hmaster0 & ~n2551;
  assign n2553 = i_hbusreq1 & ~n2539;
  assign n2554 = ~n2399 & ~n2535;
  assign n2555 = ~i_hbusreq1 & ~n2554;
  assign n2556 = ~n2553 & ~n2555;
  assign n2557 = ~controllable_hmaster0 & ~n2556;
  assign n2558 = ~n2552 & ~n2557;
  assign n2559 = i_hlock0 & ~n2558;
  assign n2560 = ~n2546 & ~n2559;
  assign n2561 = ~i_hbusreq0 & ~n2560;
  assign n2562 = ~n2548 & ~n2561;
  assign n2563 = ~n1899 & ~n2562;
  assign n2564 = ~n1899 & ~n2563;
  assign n2565 = n1980 & ~n2564;
  assign n2566 = ~n2454 & ~n2565;
  assign n2567 = n1974 & ~n2566;
  assign n2568 = ~n2453 & ~n2567;
  assign n2569 = n2042 & ~n2568;
  assign n2570 = ~n2528 & ~n2569;
  assign n2571 = n1962 & ~n2570;
  assign n2572 = ~n2425 & ~n2571;
  assign n2573 = ~n1956 & ~n2572;
  assign n2574 = ~n2492 & ~n2573;
  assign n2575 = ~n1953 & ~n2574;
  assign n2576 = ~controllable_nhgrant0 & ~n2436;
  assign n2577 = ~controllable_hgrant1 & ~n2576;
  assign n2578 = ~controllable_hgrant1 & ~n2577;
  assign n2579 = controllable_ndecide & ~n2578;
  assign n2580 = ~n2440 & ~n2579;
  assign n2581 = ~controllable_hmaster0 & ~n2580;
  assign n2582 = ~controllable_hmaster0 & ~n2581;
  assign n2583 = ~n1899 & ~n2582;
  assign n2584 = ~n1899 & ~n2583;
  assign n2585 = n1980 & ~n2584;
  assign n2586 = n1980 & ~n2585;
  assign n2587 = n1974 & ~n2586;
  assign n2588 = n1974 & ~n2587;
  assign n2589 = ~n2042 & ~n2588;
  assign n2590 = ~controllable_hgrant1 & ~n2331;
  assign n2591 = ~controllable_hgrant1 & ~n2590;
  assign n2592 = controllable_hmaster0 & ~n2591;
  assign n2593 = ~controllable_hgrant1 & controllable_nhgrant0;
  assign n2594 = ~controllable_hgrant1 & ~n2593;
  assign n2595 = controllable_ndecide & ~n2594;
  assign n2596 = ~controllable_hgrant1 & n2339;
  assign n2597 = ~n2435 & ~n2596;
  assign n2598 = ~controllable_ndecide & ~n2597;
  assign n2599 = ~n2595 & ~n2598;
  assign n2600 = ~controllable_hmaster0 & ~n2599;
  assign n2601 = ~n2592 & ~n2600;
  assign n2602 = i_hlock0 & ~n2601;
  assign n2603 = controllable_ndecide & ~n2591;
  assign n2604 = ~controllable_ndecide & ~n2458;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = controllable_hmaster0 & ~n2605;
  assign n2607 = ~n2476 & ~n2595;
  assign n2608 = ~controllable_hmaster0 & ~n2607;
  assign n2609 = ~n2606 & ~n2608;
  assign n2610 = ~i_hlock0 & ~n2609;
  assign n2611 = ~n2602 & ~n2610;
  assign n2612 = ~n1899 & ~n2611;
  assign n2613 = ~n1899 & ~n2612;
  assign n2614 = n1980 & ~n2613;
  assign n2615 = ~n2454 & ~n2614;
  assign n2616 = n1974 & ~n2615;
  assign n2617 = ~n2453 & ~n2616;
  assign n2618 = n2042 & ~n2617;
  assign n2619 = ~n2589 & ~n2618;
  assign n2620 = n1962 & ~n2619;
  assign n2621 = n1962 & ~n2620;
  assign n2622 = n1956 & ~n2621;
  assign n2623 = controllable_nhgrant0 & ~n2259;
  assign n2624 = controllable_nhgrant0 & ~n2623;
  assign n2625 = controllable_hgrant1 & ~n2624;
  assign n2626 = ~n2577 & ~n2625;
  assign n2627 = controllable_ndecide & ~n2626;
  assign n2628 = ~n2440 & ~n2627;
  assign n2629 = ~controllable_hmaster0 & ~n2628;
  assign n2630 = ~controllable_hmaster0 & ~n2629;
  assign n2631 = ~n1899 & ~n2630;
  assign n2632 = ~n1899 & ~n2631;
  assign n2633 = n1980 & ~n2632;
  assign n2634 = n1980 & ~n2633;
  assign n2635 = n1974 & ~n2634;
  assign n2636 = n1974 & ~n2635;
  assign n2637 = ~n2042 & ~n2636;
  assign n2638 = ~n2593 & ~n2625;
  assign n2639 = controllable_ndecide & ~n2638;
  assign n2640 = ~n2598 & ~n2639;
  assign n2641 = ~controllable_hmaster0 & ~n2640;
  assign n2642 = ~n2592 & ~n2641;
  assign n2643 = i_hlock0 & ~n2642;
  assign n2644 = ~n2476 & ~n2639;
  assign n2645 = ~controllable_hmaster0 & ~n2644;
  assign n2646 = ~n2606 & ~n2645;
  assign n2647 = ~i_hlock0 & ~n2646;
  assign n2648 = ~n2643 & ~n2647;
  assign n2649 = ~n1899 & ~n2648;
  assign n2650 = ~n1899 & ~n2649;
  assign n2651 = n1980 & ~n2650;
  assign n2652 = ~n2454 & ~n2651;
  assign n2653 = n1974 & ~n2652;
  assign n2654 = ~n2453 & ~n2653;
  assign n2655 = n2042 & ~n2654;
  assign n2656 = ~n2637 & ~n2655;
  assign n2657 = n1962 & ~n2656;
  assign n2658 = n1962 & ~n2657;
  assign n2659 = ~n1956 & ~n2658;
  assign n2660 = ~n2622 & ~n2659;
  assign n2661 = n1953 & ~n2660;
  assign n2662 = ~n2575 & ~n2661;
  assign n2663 = n1947 & ~n2662;
  assign n2664 = ~n2387 & ~n2663;
  assign n2665 = ~n1944 & ~n2664;
  assign n2666 = ~n1996 & ~n2401;
  assign n2667 = i_hlock0 & ~n2666;
  assign n2668 = ~n2015 & ~n2412;
  assign n2669 = ~i_hlock0 & ~n2668;
  assign n2670 = ~n2667 & ~n2669;
  assign n2671 = i_hbusreq0 & ~n2670;
  assign n2672 = ~n2022 & ~n2401;
  assign n2673 = i_hlock0 & ~n2672;
  assign n2674 = ~n2027 & ~n2412;
  assign n2675 = ~i_hlock0 & ~n2674;
  assign n2676 = ~n2673 & ~n2675;
  assign n2677 = ~i_hbusreq0 & ~n2676;
  assign n2678 = ~n2671 & ~n2677;
  assign n2679 = ~n1899 & ~n2678;
  assign n2680 = ~n1899 & ~n2679;
  assign n2681 = n1980 & ~n2680;
  assign n2682 = n1980 & ~n2681;
  assign n2683 = n1974 & ~n2682;
  assign n2684 = n1974 & ~n2683;
  assign n2685 = n2042 & ~n2684;
  assign n2686 = n2042 & ~n2685;
  assign n2687 = ~n1962 & ~n2686;
  assign n2688 = controllable_locked & ~controllable_nhgrant0;
  assign n2689 = ~controllable_nhgrant0 & ~n2688;
  assign n2690 = ~controllable_hgrant1 & ~n2689;
  assign n2691 = ~controllable_hgrant1 & ~n2690;
  assign n2692 = controllable_ndecide & ~n2691;
  assign n2693 = ~n2096 & ~n2692;
  assign n2694 = controllable_hmaster0 & ~n2693;
  assign n2695 = controllable_locked & ~n2001;
  assign n2696 = ~controllable_locked & n1982;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = controllable_nhgrant0 & ~n2697;
  assign n2699 = ~controllable_nhgrant0 & ~n2001;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = controllable_hgrant1 & ~n2700;
  assign n2702 = ~n2397 & ~n2701;
  assign n2703 = ~i_hlock1 & ~n2702;
  assign n2704 = ~n2498 & ~n2703;
  assign n2705 = ~controllable_ndecide & ~n2704;
  assign n2706 = ~n2466 & ~n2705;
  assign n2707 = ~controllable_hmaster0 & ~n2706;
  assign n2708 = ~n2694 & ~n2707;
  assign n2709 = i_hlock0 & ~n2708;
  assign n2710 = i_hready & controllable_locked;
  assign n2711 = ~controllable_nhgrant0 & n2710;
  assign n2712 = ~n2339 & ~n2711;
  assign n2713 = ~controllable_hgrant1 & n2712;
  assign n2714 = ~n2115 & ~n2713;
  assign n2715 = ~controllable_ndecide & n2714;
  assign n2716 = ~n2692 & ~n2715;
  assign n2717 = controllable_hmaster0 & ~n2716;
  assign n2718 = controllable_nhgrant0 & n2710;
  assign n2719 = i_hready & ~controllable_nhgrant0;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = controllable_hgrant1 & ~n2720;
  assign n2722 = ~n2474 & ~n2721;
  assign n2723 = ~controllable_ndecide & ~n2722;
  assign n2724 = ~n2466 & ~n2723;
  assign n2725 = ~controllable_hmaster0 & ~n2724;
  assign n2726 = ~n2717 & ~n2725;
  assign n2727 = ~i_hlock0 & ~n2726;
  assign n2728 = ~n2709 & ~n2727;
  assign n2729 = i_hbusreq0 & ~n2728;
  assign n2730 = i_hbusreq1 & ~n2693;
  assign n2731 = controllable_ndecide & ~n2692;
  assign n2732 = ~i_hbusreq1 & ~n2731;
  assign n2733 = ~n2730 & ~n2732;
  assign n2734 = controllable_hmaster0 & ~n2733;
  assign n2735 = i_hbusreq1 & ~n2706;
  assign n2736 = ~i_hbusreq1 & ~n2467;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = ~controllable_hmaster0 & ~n2737;
  assign n2739 = ~n2734 & ~n2738;
  assign n2740 = i_hlock0 & ~n2739;
  assign n2741 = ~n2727 & ~n2740;
  assign n2742 = ~i_hbusreq0 & ~n2741;
  assign n2743 = ~n2729 & ~n2742;
  assign n2744 = ~n1899 & ~n2743;
  assign n2745 = ~n1899 & ~n2744;
  assign n2746 = n1980 & ~n2745;
  assign n2747 = n1980 & ~n2746;
  assign n2748 = n1974 & ~n2747;
  assign n2749 = n1974 & ~n2748;
  assign n2750 = n2042 & ~n2749;
  assign n2751 = n2042 & ~n2750;
  assign n2752 = n1962 & ~n2751;
  assign n2753 = ~n2687 & ~n2752;
  assign n2754 = n1956 & ~n2753;
  assign n2755 = ~controllable_hmaster0 & n2400;
  assign n2756 = ~n2156 & ~n2755;
  assign n2757 = i_hlock0 & ~n2756;
  assign n2758 = ~controllable_hmaster0 & n2411;
  assign n2759 = ~n2156 & ~n2758;
  assign n2760 = ~i_hlock0 & ~n2759;
  assign n2761 = ~n2757 & ~n2760;
  assign n2762 = i_hbusreq0 & ~n2761;
  assign n2763 = ~n2161 & ~n2755;
  assign n2764 = i_hlock0 & ~n2763;
  assign n2765 = ~n2161 & ~n2758;
  assign n2766 = ~i_hlock0 & ~n2765;
  assign n2767 = ~n2764 & ~n2766;
  assign n2768 = ~i_hbusreq0 & ~n2767;
  assign n2769 = ~n2762 & ~n2768;
  assign n2770 = ~n1899 & n2769;
  assign n2771 = ~n1899 & ~n2770;
  assign n2772 = n1980 & ~n2771;
  assign n2773 = n1980 & ~n2772;
  assign n2774 = n1974 & ~n2773;
  assign n2775 = n1974 & ~n2774;
  assign n2776 = n2042 & ~n2775;
  assign n2777 = n2042 & ~n2776;
  assign n2778 = ~n1962 & ~n2777;
  assign n2779 = ~controllable_hgrant1 & n2689;
  assign n2780 = ~n2211 & ~n2779;
  assign n2781 = controllable_ndecide & ~n2780;
  assign n2782 = ~i_hlock1 & ~n2714;
  assign n2783 = ~n2010 & ~n2782;
  assign n2784 = ~controllable_ndecide & ~n2783;
  assign n2785 = ~n2781 & ~n2784;
  assign n2786 = controllable_hmaster0 & ~n2785;
  assign n2787 = controllable_locked & controllable_nhgrant0;
  assign n2788 = controllable_nhgrant0 & ~n2787;
  assign n2789 = controllable_hgrant1 & ~n2788;
  assign n2790 = ~n2464 & ~n2789;
  assign n2791 = controllable_ndecide & ~n2790;
  assign n2792 = ~i_hlock1 & ~n2722;
  assign n2793 = ~n2498 & ~n2792;
  assign n2794 = ~controllable_ndecide & ~n2793;
  assign n2795 = ~n2791 & ~n2794;
  assign n2796 = ~controllable_hmaster0 & n2795;
  assign n2797 = ~n2786 & ~n2796;
  assign n2798 = i_hlock0 & ~n2797;
  assign n2799 = ~controllable_ndecide & ~n2714;
  assign n2800 = ~n2781 & ~n2799;
  assign n2801 = controllable_hmaster0 & ~n2800;
  assign n2802 = ~n2723 & ~n2791;
  assign n2803 = ~controllable_hmaster0 & n2802;
  assign n2804 = ~n2801 & ~n2803;
  assign n2805 = ~i_hlock0 & ~n2804;
  assign n2806 = ~n2798 & ~n2805;
  assign n2807 = i_hbusreq0 & ~n2806;
  assign n2808 = i_hbusreq1 & ~n2785;
  assign n2809 = ~i_hbusreq1 & n2781;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = controllable_hmaster0 & ~n2810;
  assign n2812 = i_hbusreq1 & ~n2795;
  assign n2813 = ~n2399 & ~n2791;
  assign n2814 = ~i_hbusreq1 & ~n2813;
  assign n2815 = ~n2812 & ~n2814;
  assign n2816 = ~controllable_hmaster0 & n2815;
  assign n2817 = ~n2811 & ~n2816;
  assign n2818 = i_hlock0 & ~n2817;
  assign n2819 = ~n2805 & ~n2818;
  assign n2820 = ~i_hbusreq0 & ~n2819;
  assign n2821 = ~n2807 & ~n2820;
  assign n2822 = ~n1899 & n2821;
  assign n2823 = ~n1899 & ~n2822;
  assign n2824 = n1980 & ~n2823;
  assign n2825 = n1980 & ~n2824;
  assign n2826 = n1974 & ~n2825;
  assign n2827 = n1974 & ~n2826;
  assign n2828 = n2042 & ~n2827;
  assign n2829 = n2042 & ~n2828;
  assign n2830 = n1962 & ~n2829;
  assign n2831 = ~n2778 & ~n2830;
  assign n2832 = ~n1956 & ~n2831;
  assign n2833 = ~n2754 & ~n2832;
  assign n2834 = ~n1953 & ~n2833;
  assign n2835 = controllable_locked & ~n2695;
  assign n2836 = ~controllable_nhgrant0 & n2835;
  assign n2837 = ~controllable_nhgrant0 & ~n2836;
  assign n2838 = ~controllable_hgrant1 & ~n2837;
  assign n2839 = ~controllable_hgrant1 & ~n2838;
  assign n2840 = controllable_ndecide & ~n2839;
  assign n2841 = ~n2005 & ~n2405;
  assign n2842 = ~controllable_hgrant1 & ~n2841;
  assign n2843 = ~n2092 & ~n2842;
  assign n2844 = ~controllable_ndecide & ~n2843;
  assign n2845 = ~n2840 & ~n2844;
  assign n2846 = controllable_hmaster0 & ~n2845;
  assign n2847 = ~n2596 & ~n2721;
  assign n2848 = ~controllable_ndecide & ~n2847;
  assign n2849 = ~n2595 & ~n2848;
  assign n2850 = ~controllable_hmaster0 & ~n2849;
  assign n2851 = ~n2846 & ~n2850;
  assign n2852 = i_hlock0 & ~n2851;
  assign n2853 = ~n2715 & ~n2840;
  assign n2854 = controllable_hmaster0 & ~n2853;
  assign n2855 = ~n2595 & ~n2723;
  assign n2856 = ~controllable_hmaster0 & ~n2855;
  assign n2857 = ~n2854 & ~n2856;
  assign n2858 = ~i_hlock0 & ~n2857;
  assign n2859 = ~n2852 & ~n2858;
  assign n2860 = ~n1899 & ~n2859;
  assign n2861 = ~n1899 & ~n2860;
  assign n2862 = n1980 & ~n2861;
  assign n2863 = n1980 & ~n2862;
  assign n2864 = n1974 & ~n2863;
  assign n2865 = n1974 & ~n2864;
  assign n2866 = n2042 & ~n2865;
  assign n2867 = n2042 & ~n2866;
  assign n2868 = n1962 & ~n2867;
  assign n2869 = n1962 & ~n2868;
  assign n2870 = n1956 & ~n2869;
  assign n2871 = ~controllable_hgrant1 & n2837;
  assign n2872 = ~n2328 & ~n2871;
  assign n2873 = controllable_ndecide & ~n2872;
  assign n2874 = ~controllable_hgrant1 & ~n2339;
  assign n2875 = ~n2332 & ~n2874;
  assign n2876 = i_hlock1 & ~n2875;
  assign n2877 = ~n2115 & ~n2874;
  assign n2878 = ~i_hlock1 & ~n2877;
  assign n2879 = ~n2876 & ~n2878;
  assign n2880 = ~controllable_ndecide & ~n2879;
  assign n2881 = ~n2873 & ~n2880;
  assign n2882 = controllable_hmaster0 & ~n2881;
  assign n2883 = controllable_nhgrant0 & ~n2835;
  assign n2884 = controllable_hgrant1 & n2883;
  assign n2885 = ~controllable_hgrant1 & ~controllable_nhgrant0;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = controllable_ndecide & ~n2886;
  assign n2888 = ~i_hlock1 & n2847;
  assign n2889 = ~n2876 & ~n2888;
  assign n2890 = ~controllable_ndecide & ~n2889;
  assign n2891 = ~n2887 & ~n2890;
  assign n2892 = ~controllable_hmaster0 & ~n2891;
  assign n2893 = ~n2882 & ~n2892;
  assign n2894 = i_hlock0 & ~n2893;
  assign n2895 = ~n2332 & ~n2713;
  assign n2896 = i_hlock1 & ~n2895;
  assign n2897 = ~n2782 & ~n2896;
  assign n2898 = ~controllable_ndecide & ~n2897;
  assign n2899 = ~n2873 & ~n2898;
  assign n2900 = controllable_hmaster0 & ~n2899;
  assign n2901 = ~controllable_hgrant1 & n2473;
  assign n2902 = ~n2332 & ~n2901;
  assign n2903 = i_hlock1 & ~n2902;
  assign n2904 = ~i_hlock1 & n2722;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = ~controllable_ndecide & ~n2905;
  assign n2907 = ~n2887 & ~n2906;
  assign n2908 = ~controllable_hmaster0 & ~n2907;
  assign n2909 = ~n2900 & ~n2908;
  assign n2910 = ~i_hlock0 & ~n2909;
  assign n2911 = ~n2894 & ~n2910;
  assign n2912 = i_hbusreq0 & ~n2911;
  assign n2913 = i_hbusreq1 & ~n2881;
  assign n2914 = ~controllable_ndecide & n2843;
  assign n2915 = ~n2873 & ~n2914;
  assign n2916 = ~i_hbusreq1 & ~n2915;
  assign n2917 = ~n2913 & ~n2916;
  assign n2918 = controllable_hmaster0 & ~n2917;
  assign n2919 = i_hbusreq1 & ~n2891;
  assign n2920 = ~controllable_ndecide & n2847;
  assign n2921 = ~n2887 & ~n2920;
  assign n2922 = ~i_hbusreq1 & ~n2921;
  assign n2923 = ~n2919 & ~n2922;
  assign n2924 = ~controllable_hmaster0 & ~n2923;
  assign n2925 = ~n2918 & ~n2924;
  assign n2926 = i_hlock0 & ~n2925;
  assign n2927 = i_hbusreq1 & ~n2899;
  assign n2928 = ~n2799 & ~n2873;
  assign n2929 = ~i_hbusreq1 & ~n2928;
  assign n2930 = ~n2927 & ~n2929;
  assign n2931 = controllable_hmaster0 & ~n2930;
  assign n2932 = i_hbusreq1 & ~n2907;
  assign n2933 = ~controllable_ndecide & n2722;
  assign n2934 = ~n2887 & ~n2933;
  assign n2935 = ~i_hbusreq1 & ~n2934;
  assign n2936 = ~n2932 & ~n2935;
  assign n2937 = ~controllable_hmaster0 & ~n2936;
  assign n2938 = ~n2931 & ~n2937;
  assign n2939 = ~i_hlock0 & ~n2938;
  assign n2940 = ~n2926 & ~n2939;
  assign n2941 = ~i_hbusreq0 & ~n2940;
  assign n2942 = ~n2912 & ~n2941;
  assign n2943 = ~n1899 & n2942;
  assign n2944 = ~n1899 & ~n2943;
  assign n2945 = n1980 & ~n2944;
  assign n2946 = n1980 & ~n2945;
  assign n2947 = n1974 & ~n2946;
  assign n2948 = n1974 & ~n2947;
  assign n2949 = n2042 & ~n2948;
  assign n2950 = n2042 & ~n2949;
  assign n2951 = n1962 & ~n2950;
  assign n2952 = n1962 & ~n2951;
  assign n2953 = ~n1956 & ~n2952;
  assign n2954 = ~n2870 & ~n2953;
  assign n2955 = n1953 & ~n2954;
  assign n2956 = ~n2834 & ~n2955;
  assign n2957 = ~n1947 & ~n2956;
  assign n2958 = ~n1925 & n1948;
  assign n2959 = ~n1926 & ~n2958;
  assign n2960 = n1924 & n2959;
  assign n2961 = ~n2680 & ~n2960;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = n1980 & ~n2962;
  assign n2964 = n1980 & ~n2963;
  assign n2965 = n1974 & ~n2964;
  assign n2966 = n1974 & ~n2965;
  assign n2967 = ~n2042 & ~n2966;
  assign n2968 = ~n2417 & ~n2960;
  assign n2969 = ~n2960 & ~n2968;
  assign n2970 = ~n1974 & ~n2969;
  assign n2971 = ~n1980 & ~n2969;
  assign n2972 = ~n2963 & ~n2971;
  assign n2973 = n1974 & ~n2972;
  assign n2974 = ~n2970 & ~n2973;
  assign n2975 = n2042 & ~n2974;
  assign n2976 = ~n2967 & ~n2975;
  assign n2977 = ~n1962 & ~n2976;
  assign n2978 = ~n2051 & ~n2432;
  assign n2979 = i_hlock0 & ~n2978;
  assign n2980 = ~n2067 & ~n2442;
  assign n2981 = ~i_hlock0 & ~n2980;
  assign n2982 = ~n2979 & ~n2981;
  assign n2983 = i_hbusreq0 & ~n2982;
  assign n2984 = ~n2076 & ~n2432;
  assign n2985 = i_hlock0 & ~n2984;
  assign n2986 = ~n2981 & ~n2985;
  assign n2987 = ~i_hbusreq0 & ~n2986;
  assign n2988 = ~n2983 & ~n2987;
  assign n2989 = ~n1899 & ~n2988;
  assign n2990 = ~n1899 & ~n2989;
  assign n2991 = n1980 & ~n2990;
  assign n2992 = n1980 & ~n2991;
  assign n2993 = n1974 & ~n2992;
  assign n2994 = n1974 & ~n2993;
  assign n2995 = ~n2042 & ~n2994;
  assign n2996 = ~n2454 & ~n2746;
  assign n2997 = n1974 & ~n2996;
  assign n2998 = ~n2453 & ~n2997;
  assign n2999 = n2042 & ~n2998;
  assign n3000 = ~n2995 & ~n2999;
  assign n3001 = n1962 & ~n3000;
  assign n3002 = ~n2977 & ~n3001;
  assign n3003 = n1956 & ~n3002;
  assign n3004 = ~n2771 & ~n2960;
  assign n3005 = ~n2960 & ~n3004;
  assign n3006 = n1980 & ~n3005;
  assign n3007 = n1980 & ~n3006;
  assign n3008 = n1974 & ~n3007;
  assign n3009 = n1974 & ~n3008;
  assign n3010 = ~n2042 & ~n3009;
  assign n3011 = n2042 & ~n3005;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n1962 & ~n3012;
  assign n3014 = ~controllable_hmaster0 & n2502;
  assign n3015 = ~n2184 & ~n3014;
  assign n3016 = i_hlock0 & ~n3015;
  assign n3017 = ~controllable_hmaster0 & n2506;
  assign n3018 = ~n2188 & ~n3017;
  assign n3019 = ~i_hlock0 & ~n3018;
  assign n3020 = ~n3016 & ~n3019;
  assign n3021 = i_hbusreq0 & ~n3020;
  assign n3022 = ~controllable_hmaster0 & n2515;
  assign n3023 = ~n2195 & ~n3022;
  assign n3024 = i_hlock0 & ~n3023;
  assign n3025 = ~n3019 & ~n3024;
  assign n3026 = ~i_hbusreq0 & ~n3025;
  assign n3027 = ~n3021 & ~n3026;
  assign n3028 = ~n1899 & n3027;
  assign n3029 = ~n1899 & ~n3028;
  assign n3030 = n1980 & ~n3029;
  assign n3031 = n1980 & ~n3030;
  assign n3032 = n1974 & ~n3031;
  assign n3033 = n1974 & ~n3032;
  assign n3034 = ~n2042 & ~n3033;
  assign n3035 = ~n1974 & ~n2771;
  assign n3036 = ~n1980 & ~n2771;
  assign n3037 = ~n2824 & ~n3036;
  assign n3038 = n1974 & ~n3037;
  assign n3039 = ~n3035 & ~n3038;
  assign n3040 = n2042 & ~n3039;
  assign n3041 = ~n3034 & ~n3040;
  assign n3042 = n1962 & ~n3041;
  assign n3043 = ~n3013 & ~n3042;
  assign n3044 = ~n1956 & ~n3043;
  assign n3045 = ~n3003 & ~n3044;
  assign n3046 = ~n1953 & ~n3045;
  assign n3047 = ~n2267 & ~n2581;
  assign n3048 = i_hlock0 & ~n3047;
  assign n3049 = ~n2271 & ~n2581;
  assign n3050 = ~i_hlock0 & ~n3049;
  assign n3051 = ~n3048 & ~n3050;
  assign n3052 = ~n1899 & ~n3051;
  assign n3053 = ~n1899 & ~n3052;
  assign n3054 = n1980 & ~n3053;
  assign n3055 = n1980 & ~n3054;
  assign n3056 = n1974 & ~n3055;
  assign n3057 = n1974 & ~n3056;
  assign n3058 = ~n2042 & ~n3057;
  assign n3059 = ~n2454 & ~n2862;
  assign n3060 = n1974 & ~n3059;
  assign n3061 = ~n2453 & ~n3060;
  assign n3062 = n2042 & ~n3061;
  assign n3063 = ~n3058 & ~n3062;
  assign n3064 = n1962 & ~n3063;
  assign n3065 = n1962 & ~n3064;
  assign n3066 = n1956 & ~n3065;
  assign n3067 = ~controllable_hmaster0 & n2628;
  assign n3068 = ~n2308 & ~n3067;
  assign n3069 = i_hbusreq0 & ~n3068;
  assign n3070 = ~n2315 & ~n3067;
  assign n3071 = i_hlock0 & ~n3070;
  assign n3072 = ~i_hlock0 & ~n3068;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~i_hbusreq0 & ~n3073;
  assign n3075 = ~n3069 & ~n3074;
  assign n3076 = ~n1899 & n3075;
  assign n3077 = ~n1899 & ~n3076;
  assign n3078 = n1980 & ~n3077;
  assign n3079 = n1980 & ~n3078;
  assign n3080 = n1974 & ~n3079;
  assign n3081 = n1974 & ~n3080;
  assign n3082 = ~n2042 & ~n3081;
  assign n3083 = ~n2945 & ~n3036;
  assign n3084 = n1974 & ~n3083;
  assign n3085 = ~n3035 & ~n3084;
  assign n3086 = n2042 & ~n3085;
  assign n3087 = ~n3082 & ~n3086;
  assign n3088 = n1962 & ~n3087;
  assign n3089 = n1962 & ~n3088;
  assign n3090 = ~n1956 & ~n3089;
  assign n3091 = ~n3066 & ~n3090;
  assign n3092 = n1953 & ~n3091;
  assign n3093 = ~n3046 & ~n3092;
  assign n3094 = n1947 & ~n3093;
  assign n3095 = ~n2957 & ~n3094;
  assign n3096 = n1944 & ~n3095;
  assign n3097 = ~n2665 & ~n3096;
  assign n3098 = ~n1942 & ~n3097;
  assign n3099 = ~n1942 & ~n3098;
  assign n3100 = n1939 & ~n3099;
  assign n3101 = ~n2034 & n2960;
  assign n3102 = ~controllable_locked & ~n1984;
  assign n3103 = ~controllable_nhgrant0 & ~n3102;
  assign n3104 = ~controllable_nhgrant0 & ~n3103;
  assign n3105 = ~controllable_hgrant1 & ~n3104;
  assign n3106 = ~controllable_hgrant1 & ~n3105;
  assign n3107 = controllable_ndecide & ~n3106;
  assign n3108 = controllable_ndecide & ~n3107;
  assign n3109 = ~controllable_hmaster0 & ~n3108;
  assign n3110 = ~n1996 & ~n3109;
  assign n3111 = i_hlock0 & ~n3110;
  assign n3112 = ~n2410 & ~n3107;
  assign n3113 = ~controllable_hmaster0 & ~n3112;
  assign n3114 = ~n2015 & ~n3113;
  assign n3115 = ~i_hlock0 & ~n3114;
  assign n3116 = ~n3111 & ~n3115;
  assign n3117 = i_hbusreq0 & ~n3116;
  assign n3118 = ~n2022 & ~n3109;
  assign n3119 = i_hlock0 & ~n3118;
  assign n3120 = ~n2027 & ~n3113;
  assign n3121 = ~i_hlock0 & ~n3120;
  assign n3122 = ~n3119 & ~n3121;
  assign n3123 = ~i_hbusreq0 & ~n3122;
  assign n3124 = ~n3117 & ~n3123;
  assign n3125 = ~n1899 & ~n3124;
  assign n3126 = ~n1899 & ~n3125;
  assign n3127 = ~n2960 & ~n3126;
  assign n3128 = ~n3101 & ~n3127;
  assign n3129 = n1980 & ~n3128;
  assign n3130 = n1980 & ~n3129;
  assign n3131 = n1974 & ~n3130;
  assign n3132 = n1974 & ~n3131;
  assign n3133 = ~n1962 & ~n3132;
  assign n3134 = ~i_hlock1 & ~n2398;
  assign n3135 = ~i_hlock1 & ~n3134;
  assign n3136 = ~controllable_ndecide & ~n3135;
  assign n3137 = ~controllable_ndecide & ~n3136;
  assign n3138 = ~controllable_hmaster0 & ~n3137;
  assign n3139 = ~n2051 & ~n3138;
  assign n3140 = i_hlock0 & ~n3139;
  assign n3141 = ~i_hlock1 & ~n2499;
  assign n3142 = ~controllable_ndecide & ~n3141;
  assign n3143 = ~controllable_ndecide & ~n3142;
  assign n3144 = ~controllable_hmaster0 & ~n3143;
  assign n3145 = ~n2067 & ~n3144;
  assign n3146 = ~i_hlock0 & ~n3145;
  assign n3147 = ~n3140 & ~n3146;
  assign n3148 = i_hbusreq0 & ~n3147;
  assign n3149 = i_hbusreq1 & ~n3137;
  assign n3150 = i_hbusreq1 & ~n3149;
  assign n3151 = ~controllable_hmaster0 & ~n3150;
  assign n3152 = ~n2076 & ~n3151;
  assign n3153 = i_hlock0 & ~n3152;
  assign n3154 = i_hbusreq1 & ~n3143;
  assign n3155 = i_hbusreq1 & ~n3154;
  assign n3156 = ~controllable_hmaster0 & ~n3155;
  assign n3157 = ~n2067 & ~n3156;
  assign n3158 = ~i_hlock0 & ~n3157;
  assign n3159 = ~n3153 & ~n3158;
  assign n3160 = ~i_hbusreq0 & ~n3159;
  assign n3161 = ~n3148 & ~n3160;
  assign n3162 = ~n1899 & ~n3161;
  assign n3163 = ~n1899 & ~n3162;
  assign n3164 = n2960 & ~n3163;
  assign n3165 = ~n3107 & ~n3136;
  assign n3166 = ~controllable_hmaster0 & ~n3165;
  assign n3167 = ~n2051 & ~n3166;
  assign n3168 = i_hlock0 & ~n3167;
  assign n3169 = i_hlock1 & ~n2409;
  assign n3170 = ~n2499 & ~n3169;
  assign n3171 = ~controllable_ndecide & ~n3170;
  assign n3172 = ~n3107 & ~n3171;
  assign n3173 = ~controllable_hmaster0 & ~n3172;
  assign n3174 = ~n2067 & ~n3173;
  assign n3175 = ~i_hlock0 & ~n3174;
  assign n3176 = ~n3168 & ~n3175;
  assign n3177 = i_hbusreq0 & ~n3176;
  assign n3178 = i_hbusreq1 & ~n3165;
  assign n3179 = ~i_hbusreq1 & ~n3108;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~controllable_hmaster0 & ~n3180;
  assign n3182 = ~n2076 & ~n3181;
  assign n3183 = i_hlock0 & ~n3182;
  assign n3184 = i_hbusreq1 & ~n3172;
  assign n3185 = ~i_hbusreq1 & ~n3112;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~controllable_hmaster0 & ~n3186;
  assign n3188 = ~n2067 & ~n3187;
  assign n3189 = ~i_hlock0 & ~n3188;
  assign n3190 = ~n3183 & ~n3189;
  assign n3191 = ~i_hbusreq0 & ~n3190;
  assign n3192 = ~n3177 & ~n3191;
  assign n3193 = ~n1899 & ~n3192;
  assign n3194 = ~n1899 & ~n3193;
  assign n3195 = ~n2960 & ~n3194;
  assign n3196 = ~n3164 & ~n3195;
  assign n3197 = n1980 & ~n3196;
  assign n3198 = n1980 & ~n3197;
  assign n3199 = n1974 & ~n3198;
  assign n3200 = n1974 & ~n3199;
  assign n3201 = ~n2042 & ~n3200;
  assign n3202 = ~i_hlock1 & ~n2703;
  assign n3203 = ~controllable_ndecide & ~n3202;
  assign n3204 = ~controllable_ndecide & ~n3203;
  assign n3205 = ~controllable_hmaster0 & ~n3204;
  assign n3206 = ~n2098 & ~n3205;
  assign n3207 = i_hlock0 & ~n3206;
  assign n3208 = i_hlock1 & ~n2116;
  assign n3209 = ~n2782 & ~n3208;
  assign n3210 = ~controllable_ndecide & n3209;
  assign n3211 = ~n2049 & ~n3210;
  assign n3212 = controllable_hmaster0 & ~n3211;
  assign n3213 = i_hlock1 & ~n2104;
  assign n3214 = ~n2792 & ~n3213;
  assign n3215 = ~controllable_ndecide & ~n3214;
  assign n3216 = ~controllable_ndecide & ~n3215;
  assign n3217 = ~controllable_hmaster0 & ~n3216;
  assign n3218 = ~n3212 & ~n3217;
  assign n3219 = ~i_hlock0 & ~n3218;
  assign n3220 = ~n3207 & ~n3219;
  assign n3221 = i_hbusreq0 & ~n3220;
  assign n3222 = i_hbusreq1 & ~n3204;
  assign n3223 = i_hbusreq1 & ~n3222;
  assign n3224 = ~controllable_hmaster0 & ~n3223;
  assign n3225 = ~n2129 & ~n3224;
  assign n3226 = i_hlock0 & ~n3225;
  assign n3227 = i_hbusreq1 & ~n3211;
  assign n3228 = ~i_hbusreq1 & ~n2118;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = controllable_hmaster0 & ~n3229;
  assign n3231 = i_hbusreq1 & ~n3216;
  assign n3232 = ~i_hbusreq1 & ~n2121;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = ~controllable_hmaster0 & ~n3233;
  assign n3235 = ~n3230 & ~n3234;
  assign n3236 = ~i_hlock0 & ~n3235;
  assign n3237 = ~n3226 & ~n3236;
  assign n3238 = ~i_hbusreq0 & ~n3237;
  assign n3239 = ~n3221 & ~n3238;
  assign n3240 = ~n1899 & ~n3239;
  assign n3241 = ~n1899 & ~n3240;
  assign n3242 = n2960 & ~n3241;
  assign n3243 = ~controllable_locked & ~n2002;
  assign n3244 = ~controllable_nhgrant0 & ~n3243;
  assign n3245 = ~controllable_nhgrant0 & ~n3244;
  assign n3246 = ~controllable_hgrant1 & ~n3245;
  assign n3247 = ~controllable_hgrant1 & ~n3246;
  assign n3248 = controllable_ndecide & ~n3247;
  assign n3249 = ~n3203 & ~n3248;
  assign n3250 = ~controllable_hmaster0 & ~n3249;
  assign n3251 = ~n2694 & ~n3250;
  assign n3252 = i_hlock0 & ~n3251;
  assign n3253 = ~controllable_nhgrant0 & ~n2089;
  assign n3254 = ~n2405 & ~n3253;
  assign n3255 = ~controllable_hgrant1 & ~n3254;
  assign n3256 = ~n2092 & ~n3255;
  assign n3257 = i_hlock1 & ~n3256;
  assign n3258 = ~n2792 & ~n3257;
  assign n3259 = ~controllable_ndecide & ~n3258;
  assign n3260 = ~n3248 & ~n3259;
  assign n3261 = ~controllable_hmaster0 & ~n3260;
  assign n3262 = ~n2717 & ~n3261;
  assign n3263 = ~i_hlock0 & ~n3262;
  assign n3264 = ~n3252 & ~n3263;
  assign n3265 = i_hbusreq0 & ~n3264;
  assign n3266 = i_hbusreq1 & ~n3249;
  assign n3267 = controllable_ndecide & ~n3248;
  assign n3268 = ~i_hbusreq1 & ~n3267;
  assign n3269 = ~n3266 & ~n3268;
  assign n3270 = ~controllable_hmaster0 & ~n3269;
  assign n3271 = ~n2734 & ~n3270;
  assign n3272 = i_hlock0 & ~n3271;
  assign n3273 = i_hbusreq1 & ~n3260;
  assign n3274 = ~controllable_ndecide & ~n3256;
  assign n3275 = ~n3248 & ~n3274;
  assign n3276 = ~i_hbusreq1 & ~n3275;
  assign n3277 = ~n3273 & ~n3276;
  assign n3278 = ~controllable_hmaster0 & ~n3277;
  assign n3279 = ~n2717 & ~n3278;
  assign n3280 = ~i_hlock0 & ~n3279;
  assign n3281 = ~n3272 & ~n3280;
  assign n3282 = ~i_hbusreq0 & ~n3281;
  assign n3283 = ~n3265 & ~n3282;
  assign n3284 = ~n1899 & ~n3283;
  assign n3285 = ~n1899 & ~n3284;
  assign n3286 = ~n2960 & ~n3285;
  assign n3287 = ~n3242 & ~n3286;
  assign n3288 = n1980 & ~n3287;
  assign n3289 = n1980 & ~n3288;
  assign n3290 = n1974 & ~n3289;
  assign n3291 = n1974 & ~n3290;
  assign n3292 = n2042 & ~n3291;
  assign n3293 = ~n3201 & ~n3292;
  assign n3294 = n1962 & ~n3293;
  assign n3295 = ~n3133 & ~n3294;
  assign n3296 = n1956 & ~n3295;
  assign n3297 = ~n2165 & n2960;
  assign n3298 = ~controllable_hmaster0 & n3108;
  assign n3299 = ~n2156 & ~n3298;
  assign n3300 = i_hlock0 & ~n3299;
  assign n3301 = ~controllable_hmaster0 & n3112;
  assign n3302 = ~n2156 & ~n3301;
  assign n3303 = ~i_hlock0 & ~n3302;
  assign n3304 = ~n3300 & ~n3303;
  assign n3305 = i_hbusreq0 & ~n3304;
  assign n3306 = ~n2161 & ~n3298;
  assign n3307 = i_hlock0 & ~n3306;
  assign n3308 = ~n2161 & ~n3301;
  assign n3309 = ~i_hlock0 & ~n3308;
  assign n3310 = ~n3307 & ~n3309;
  assign n3311 = ~i_hbusreq0 & ~n3310;
  assign n3312 = ~n3305 & ~n3311;
  assign n3313 = ~n1899 & n3312;
  assign n3314 = ~n1899 & ~n3313;
  assign n3315 = ~n2960 & ~n3314;
  assign n3316 = ~n3297 & ~n3315;
  assign n3317 = n1980 & ~n3316;
  assign n3318 = n1980 & ~n3317;
  assign n3319 = n1974 & ~n3318;
  assign n3320 = n1974 & ~n3319;
  assign n3321 = ~n2042 & ~n3320;
  assign n3322 = ~n2208 & ~n3317;
  assign n3323 = n1974 & ~n3322;
  assign n3324 = ~n2207 & ~n3323;
  assign n3325 = n2042 & ~n3324;
  assign n3326 = ~n3321 & ~n3325;
  assign n3327 = ~n1962 & ~n3326;
  assign n3328 = controllable_hgrant1 & ~n2495;
  assign n3329 = controllable_ndecide & ~n3328;
  assign n3330 = ~n3142 & ~n3329;
  assign n3331 = ~controllable_hmaster0 & n3330;
  assign n3332 = ~n2184 & ~n3331;
  assign n3333 = i_hlock0 & ~n3332;
  assign n3334 = ~n2188 & ~n3331;
  assign n3335 = ~i_hlock0 & ~n3334;
  assign n3336 = ~n3333 & ~n3335;
  assign n3337 = i_hbusreq0 & ~n3336;
  assign n3338 = i_hbusreq1 & ~n3330;
  assign n3339 = controllable_ndecide & ~n3329;
  assign n3340 = ~i_hbusreq1 & ~n3339;
  assign n3341 = ~n3338 & ~n3340;
  assign n3342 = ~controllable_hmaster0 & n3341;
  assign n3343 = ~n2195 & ~n3342;
  assign n3344 = i_hlock0 & ~n3343;
  assign n3345 = ~n2188 & ~n3342;
  assign n3346 = ~i_hlock0 & ~n3345;
  assign n3347 = ~n3344 & ~n3346;
  assign n3348 = ~i_hbusreq0 & ~n3347;
  assign n3349 = ~n3337 & ~n3348;
  assign n3350 = ~n1899 & n3349;
  assign n3351 = ~n1899 & ~n3350;
  assign n3352 = n2960 & ~n3351;
  assign n3353 = ~n2495 & ~n3105;
  assign n3354 = controllable_ndecide & ~n3353;
  assign n3355 = ~n3142 & ~n3354;
  assign n3356 = ~controllable_hmaster0 & n3355;
  assign n3357 = ~n2184 & ~n3356;
  assign n3358 = i_hlock0 & ~n3357;
  assign n3359 = ~n3171 & ~n3354;
  assign n3360 = ~controllable_hmaster0 & n3359;
  assign n3361 = ~n2188 & ~n3360;
  assign n3362 = ~i_hlock0 & ~n3361;
  assign n3363 = ~n3358 & ~n3362;
  assign n3364 = i_hbusreq0 & ~n3363;
  assign n3365 = i_hbusreq1 & ~n3355;
  assign n3366 = controllable_ndecide & ~n3354;
  assign n3367 = ~i_hbusreq1 & ~n3366;
  assign n3368 = ~n3365 & ~n3367;
  assign n3369 = ~controllable_hmaster0 & n3368;
  assign n3370 = ~n2195 & ~n3369;
  assign n3371 = i_hlock0 & ~n3370;
  assign n3372 = i_hbusreq1 & ~n3359;
  assign n3373 = ~n2410 & ~n3354;
  assign n3374 = ~i_hbusreq1 & ~n3373;
  assign n3375 = ~n3372 & ~n3374;
  assign n3376 = ~controllable_hmaster0 & n3375;
  assign n3377 = ~n2188 & ~n3376;
  assign n3378 = ~i_hlock0 & ~n3377;
  assign n3379 = ~n3371 & ~n3378;
  assign n3380 = ~i_hbusreq0 & ~n3379;
  assign n3381 = ~n3364 & ~n3380;
  assign n3382 = ~n1899 & n3381;
  assign n3383 = ~n1899 & ~n3382;
  assign n3384 = ~n2960 & ~n3383;
  assign n3385 = ~n3352 & ~n3384;
  assign n3386 = n1980 & ~n3385;
  assign n3387 = n1980 & ~n3386;
  assign n3388 = n1974 & ~n3387;
  assign n3389 = n1974 & ~n3388;
  assign n3390 = ~n2042 & ~n3389;
  assign n3391 = ~n2213 & ~n2784;
  assign n3392 = controllable_hmaster0 & ~n3391;
  assign n3393 = controllable_hgrant1 & ~n2789;
  assign n3394 = controllable_ndecide & ~n3393;
  assign n3395 = ~i_hlock1 & ~n2792;
  assign n3396 = ~controllable_ndecide & ~n3395;
  assign n3397 = ~n3394 & ~n3396;
  assign n3398 = ~controllable_hmaster0 & n3397;
  assign n3399 = ~n3392 & ~n3398;
  assign n3400 = i_hlock0 & ~n3399;
  assign n3401 = ~controllable_ndecide & ~n3209;
  assign n3402 = ~n2213 & ~n3401;
  assign n3403 = controllable_hmaster0 & ~n3402;
  assign n3404 = ~n3215 & ~n3394;
  assign n3405 = ~controllable_hmaster0 & n3404;
  assign n3406 = ~n3403 & ~n3405;
  assign n3407 = ~i_hlock0 & ~n3406;
  assign n3408 = ~n3400 & ~n3407;
  assign n3409 = i_hbusreq0 & ~n3408;
  assign n3410 = i_hbusreq1 & ~n3391;
  assign n3411 = ~n2233 & ~n3410;
  assign n3412 = controllable_hmaster0 & ~n3411;
  assign n3413 = i_hbusreq1 & ~n3397;
  assign n3414 = controllable_ndecide & ~n3394;
  assign n3415 = ~i_hbusreq1 & ~n3414;
  assign n3416 = ~n3413 & ~n3415;
  assign n3417 = ~controllable_hmaster0 & n3416;
  assign n3418 = ~n3412 & ~n3417;
  assign n3419 = i_hlock0 & ~n3418;
  assign n3420 = i_hbusreq1 & ~n3402;
  assign n3421 = ~i_hbusreq1 & ~n2225;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = controllable_hmaster0 & ~n3422;
  assign n3424 = i_hbusreq1 & ~n3404;
  assign n3425 = ~n2120 & ~n3394;
  assign n3426 = ~i_hbusreq1 & ~n3425;
  assign n3427 = ~n3424 & ~n3426;
  assign n3428 = ~controllable_hmaster0 & n3427;
  assign n3429 = ~n3423 & ~n3428;
  assign n3430 = ~i_hlock0 & ~n3429;
  assign n3431 = ~n3419 & ~n3430;
  assign n3432 = ~i_hbusreq0 & ~n3431;
  assign n3433 = ~n3409 & ~n3432;
  assign n3434 = ~n1899 & n3433;
  assign n3435 = ~n1899 & ~n3434;
  assign n3436 = n2960 & ~n3435;
  assign n3437 = ~n2789 & ~n3246;
  assign n3438 = controllable_ndecide & ~n3437;
  assign n3439 = ~n3396 & ~n3438;
  assign n3440 = ~controllable_hmaster0 & n3439;
  assign n3441 = ~n2786 & ~n3440;
  assign n3442 = i_hlock0 & ~n3441;
  assign n3443 = ~n3259 & ~n3438;
  assign n3444 = ~controllable_hmaster0 & n3443;
  assign n3445 = ~n2801 & ~n3444;
  assign n3446 = ~i_hlock0 & ~n3445;
  assign n3447 = ~n3442 & ~n3446;
  assign n3448 = i_hbusreq0 & ~n3447;
  assign n3449 = i_hbusreq1 & ~n3439;
  assign n3450 = controllable_ndecide & ~n3438;
  assign n3451 = ~i_hbusreq1 & ~n3450;
  assign n3452 = ~n3449 & ~n3451;
  assign n3453 = ~controllable_hmaster0 & n3452;
  assign n3454 = ~n2811 & ~n3453;
  assign n3455 = i_hlock0 & ~n3454;
  assign n3456 = i_hbusreq1 & ~n3443;
  assign n3457 = ~n3274 & ~n3438;
  assign n3458 = ~i_hbusreq1 & ~n3457;
  assign n3459 = ~n3456 & ~n3458;
  assign n3460 = ~controllable_hmaster0 & n3459;
  assign n3461 = ~n2801 & ~n3460;
  assign n3462 = ~i_hlock0 & ~n3461;
  assign n3463 = ~n3455 & ~n3462;
  assign n3464 = ~i_hbusreq0 & ~n3463;
  assign n3465 = ~n3448 & ~n3464;
  assign n3466 = ~n1899 & n3465;
  assign n3467 = ~n1899 & ~n3466;
  assign n3468 = ~n2960 & ~n3467;
  assign n3469 = ~n3436 & ~n3468;
  assign n3470 = n1980 & ~n3469;
  assign n3471 = ~n2208 & ~n3470;
  assign n3472 = n1974 & ~n3471;
  assign n3473 = ~n2207 & ~n3472;
  assign n3474 = n2042 & ~n3473;
  assign n3475 = ~n3390 & ~n3474;
  assign n3476 = n1962 & ~n3475;
  assign n3477 = ~n3327 & ~n3476;
  assign n3478 = ~n1956 & ~n3477;
  assign n3479 = ~n3296 & ~n3478;
  assign n3480 = ~n1953 & ~n3479;
  assign n3481 = ~controllable_ndecide & ~n3171;
  assign n3482 = ~controllable_hmaster0 & ~n3481;
  assign n3483 = ~n2267 & ~n3482;
  assign n3484 = i_hlock0 & ~n3483;
  assign n3485 = ~n2271 & ~n3482;
  assign n3486 = ~i_hlock0 & ~n3485;
  assign n3487 = ~n3484 & ~n3486;
  assign n3488 = i_hbusreq0 & ~n3487;
  assign n3489 = i_hbusreq1 & ~n3481;
  assign n3490 = i_hbusreq1 & ~n3489;
  assign n3491 = ~controllable_hmaster0 & ~n3490;
  assign n3492 = ~n2267 & ~n3491;
  assign n3493 = i_hlock0 & ~n3492;
  assign n3494 = ~n2271 & ~n3491;
  assign n3495 = ~i_hlock0 & ~n3494;
  assign n3496 = ~n3493 & ~n3495;
  assign n3497 = ~i_hbusreq0 & ~n3496;
  assign n3498 = ~n3488 & ~n3497;
  assign n3499 = ~n1899 & ~n3498;
  assign n3500 = ~n1899 & ~n3499;
  assign n3501 = n2960 & ~n3500;
  assign n3502 = ~n2267 & ~n3173;
  assign n3503 = i_hlock0 & ~n3502;
  assign n3504 = ~n2271 & ~n3173;
  assign n3505 = ~i_hlock0 & ~n3504;
  assign n3506 = ~n3503 & ~n3505;
  assign n3507 = i_hbusreq0 & ~n3506;
  assign n3508 = ~n3179 & ~n3184;
  assign n3509 = ~controllable_hmaster0 & ~n3508;
  assign n3510 = ~n2267 & ~n3509;
  assign n3511 = i_hlock0 & ~n3510;
  assign n3512 = ~n2271 & ~n3187;
  assign n3513 = ~i_hlock0 & ~n3512;
  assign n3514 = ~n3511 & ~n3513;
  assign n3515 = ~i_hbusreq0 & ~n3514;
  assign n3516 = ~n3507 & ~n3515;
  assign n3517 = ~n1899 & ~n3516;
  assign n3518 = ~n1899 & ~n3517;
  assign n3519 = ~n2960 & ~n3518;
  assign n3520 = ~n3501 & ~n3519;
  assign n3521 = n1980 & ~n3520;
  assign n3522 = n1980 & ~n3521;
  assign n3523 = n1974 & ~n3522;
  assign n3524 = n1974 & ~n3523;
  assign n3525 = ~n2042 & ~n3524;
  assign n3526 = ~n2264 & ~n3274;
  assign n3527 = controllable_hmaster0 & ~n3526;
  assign n3528 = ~controllable_ndecide & ~n3259;
  assign n3529 = ~controllable_hmaster0 & ~n3528;
  assign n3530 = ~n3527 & ~n3529;
  assign n3531 = i_hlock0 & ~n3530;
  assign n3532 = ~n2264 & ~n2715;
  assign n3533 = controllable_hmaster0 & ~n3532;
  assign n3534 = ~n3529 & ~n3533;
  assign n3535 = ~i_hlock0 & ~n3534;
  assign n3536 = ~n3531 & ~n3535;
  assign n3537 = i_hbusreq0 & ~n3536;
  assign n3538 = i_hbusreq1 & ~n3526;
  assign n3539 = ~i_hbusreq1 & ~n2283;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = controllable_hmaster0 & ~n3540;
  assign n3542 = i_hbusreq1 & ~n3528;
  assign n3543 = ~n3232 & ~n3542;
  assign n3544 = ~controllable_hmaster0 & ~n3543;
  assign n3545 = ~n3541 & ~n3544;
  assign n3546 = i_hlock0 & ~n3545;
  assign n3547 = i_hbusreq1 & ~n3532;
  assign n3548 = ~i_hbusreq1 & ~n2287;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = controllable_hmaster0 & ~n3549;
  assign n3551 = ~n3544 & ~n3550;
  assign n3552 = ~i_hlock0 & ~n3551;
  assign n3553 = ~n3546 & ~n3552;
  assign n3554 = ~i_hbusreq0 & ~n3553;
  assign n3555 = ~n3537 & ~n3554;
  assign n3556 = ~n1899 & ~n3555;
  assign n3557 = ~n1899 & ~n3556;
  assign n3558 = n2960 & ~n3557;
  assign n3559 = ~controllable_nhgrant0 & n1983;
  assign n3560 = ~controllable_nhgrant0 & ~n3559;
  assign n3561 = ~controllable_hgrant1 & ~n3560;
  assign n3562 = ~controllable_hgrant1 & ~n3561;
  assign n3563 = controllable_ndecide & ~n3562;
  assign n3564 = ~n3274 & ~n3563;
  assign n3565 = controllable_hmaster0 & ~n3564;
  assign n3566 = ~n3261 & ~n3565;
  assign n3567 = i_hlock0 & ~n3566;
  assign n3568 = ~n2715 & ~n3563;
  assign n3569 = controllable_hmaster0 & ~n3568;
  assign n3570 = ~n3261 & ~n3569;
  assign n3571 = ~i_hlock0 & ~n3570;
  assign n3572 = ~n3567 & ~n3571;
  assign n3573 = i_hbusreq0 & ~n3572;
  assign n3574 = i_hbusreq1 & ~n3564;
  assign n3575 = ~n2282 & ~n3563;
  assign n3576 = ~i_hbusreq1 & ~n3575;
  assign n3577 = ~n3574 & ~n3576;
  assign n3578 = controllable_hmaster0 & ~n3577;
  assign n3579 = ~n2120 & ~n3248;
  assign n3580 = ~i_hbusreq1 & ~n3579;
  assign n3581 = ~n3273 & ~n3580;
  assign n3582 = ~controllable_hmaster0 & ~n3581;
  assign n3583 = ~n3578 & ~n3582;
  assign n3584 = i_hlock0 & ~n3583;
  assign n3585 = ~n3278 & ~n3569;
  assign n3586 = ~i_hlock0 & ~n3585;
  assign n3587 = ~n3584 & ~n3586;
  assign n3588 = ~i_hbusreq0 & ~n3587;
  assign n3589 = ~n3573 & ~n3588;
  assign n3590 = ~n1899 & ~n3589;
  assign n3591 = ~n1899 & ~n3590;
  assign n3592 = ~n2960 & ~n3591;
  assign n3593 = ~n3558 & ~n3592;
  assign n3594 = n1980 & ~n3593;
  assign n3595 = n1980 & ~n3594;
  assign n3596 = n1974 & ~n3595;
  assign n3597 = n1974 & ~n3596;
  assign n3598 = n2042 & ~n3597;
  assign n3599 = ~n3525 & ~n3598;
  assign n3600 = n1962 & ~n3599;
  assign n3601 = n1962 & ~n3600;
  assign n3602 = n1956 & ~n3601;
  assign n3603 = controllable_hgrant1 & ~n2625;
  assign n3604 = controllable_ndecide & ~n3603;
  assign n3605 = ~n3171 & ~n3604;
  assign n3606 = ~controllable_hmaster0 & n3605;
  assign n3607 = ~n2308 & ~n3606;
  assign n3608 = i_hbusreq0 & ~n3607;
  assign n3609 = i_hbusreq1 & ~n3605;
  assign n3610 = controllable_ndecide & ~n3604;
  assign n3611 = ~i_hbusreq1 & ~n3610;
  assign n3612 = ~n3609 & ~n3611;
  assign n3613 = ~controllable_hmaster0 & n3612;
  assign n3614 = ~n2315 & ~n3613;
  assign n3615 = i_hlock0 & ~n3614;
  assign n3616 = ~n2308 & ~n3613;
  assign n3617 = ~i_hlock0 & ~n3616;
  assign n3618 = ~n3615 & ~n3617;
  assign n3619 = ~i_hbusreq0 & ~n3618;
  assign n3620 = ~n3608 & ~n3619;
  assign n3621 = ~n1899 & n3620;
  assign n3622 = ~n1899 & ~n3621;
  assign n3623 = n2960 & ~n3622;
  assign n3624 = ~n2625 & ~n3105;
  assign n3625 = controllable_ndecide & ~n3624;
  assign n3626 = ~n3171 & ~n3625;
  assign n3627 = ~controllable_hmaster0 & n3626;
  assign n3628 = ~n2308 & ~n3627;
  assign n3629 = i_hbusreq0 & ~n3628;
  assign n3630 = i_hbusreq1 & ~n3626;
  assign n3631 = controllable_ndecide & ~n3625;
  assign n3632 = ~i_hbusreq1 & ~n3631;
  assign n3633 = ~n3630 & ~n3632;
  assign n3634 = ~controllable_hmaster0 & n3633;
  assign n3635 = ~n2315 & ~n3634;
  assign n3636 = i_hlock0 & ~n3635;
  assign n3637 = ~n2410 & ~n3625;
  assign n3638 = ~i_hbusreq1 & ~n3637;
  assign n3639 = ~n3630 & ~n3638;
  assign n3640 = ~controllable_hmaster0 & n3639;
  assign n3641 = ~n2308 & ~n3640;
  assign n3642 = ~i_hlock0 & ~n3641;
  assign n3643 = ~n3636 & ~n3642;
  assign n3644 = ~i_hbusreq0 & ~n3643;
  assign n3645 = ~n3629 & ~n3644;
  assign n3646 = ~n1899 & n3645;
  assign n3647 = ~n1899 & ~n3646;
  assign n3648 = ~n2960 & ~n3647;
  assign n3649 = ~n3623 & ~n3648;
  assign n3650 = n1980 & ~n3649;
  assign n3651 = n1980 & ~n3650;
  assign n3652 = n1974 & ~n3651;
  assign n3653 = n1974 & ~n3652;
  assign n3654 = ~n2042 & ~n3653;
  assign n3655 = ~n2330 & ~n2898;
  assign n3656 = controllable_hmaster0 & ~n3655;
  assign n3657 = controllable_ndecide & n2884;
  assign n3658 = ~controllable_nhgrant0 & n1982;
  assign n3659 = ~n2394 & ~n3658;
  assign n3660 = controllable_hgrant1 & ~n3659;
  assign n3661 = ~controllable_hgrant1 & n3254;
  assign n3662 = ~n3660 & ~n3661;
  assign n3663 = i_hlock1 & ~n3662;
  assign n3664 = ~n2904 & ~n3663;
  assign n3665 = ~controllable_ndecide & ~n3664;
  assign n3666 = ~n3657 & ~n3665;
  assign n3667 = ~controllable_hmaster0 & ~n3666;
  assign n3668 = ~n3656 & ~n3667;
  assign n3669 = i_hbusreq0 & ~n3668;
  assign n3670 = i_hbusreq1 & ~n3655;
  assign n3671 = ~n2353 & ~n3670;
  assign n3672 = controllable_hmaster0 & ~n3671;
  assign n3673 = i_hbusreq1 & ~n3666;
  assign n3674 = ~n2357 & ~n3657;
  assign n3675 = ~i_hbusreq1 & ~n3674;
  assign n3676 = ~n3673 & ~n3675;
  assign n3677 = ~controllable_hmaster0 & ~n3676;
  assign n3678 = ~n3672 & ~n3677;
  assign n3679 = i_hlock0 & ~n3678;
  assign n3680 = ~n2365 & ~n3670;
  assign n3681 = controllable_hmaster0 & ~n3680;
  assign n3682 = ~n3677 & ~n3681;
  assign n3683 = ~i_hlock0 & ~n3682;
  assign n3684 = ~n3679 & ~n3683;
  assign n3685 = ~i_hbusreq0 & ~n3684;
  assign n3686 = ~n3669 & ~n3685;
  assign n3687 = ~n1899 & n3686;
  assign n3688 = ~n1899 & ~n3687;
  assign n3689 = n2960 & ~n3688;
  assign n3690 = ~controllable_hgrant1 & n3560;
  assign n3691 = ~n2328 & ~n3690;
  assign n3692 = controllable_ndecide & ~n3691;
  assign n3693 = ~n2898 & ~n3692;
  assign n3694 = controllable_hmaster0 & ~n3693;
  assign n3695 = ~controllable_hgrant1 & n3245;
  assign n3696 = ~n2884 & ~n3695;
  assign n3697 = controllable_ndecide & ~n3696;
  assign n3698 = ~n3665 & ~n3697;
  assign n3699 = ~controllable_hmaster0 & ~n3698;
  assign n3700 = ~n3694 & ~n3699;
  assign n3701 = i_hbusreq0 & ~n3700;
  assign n3702 = i_hbusreq1 & ~n3693;
  assign n3703 = ~n2351 & ~n3692;
  assign n3704 = ~i_hbusreq1 & ~n3703;
  assign n3705 = ~n3702 & ~n3704;
  assign n3706 = controllable_hmaster0 & ~n3705;
  assign n3707 = i_hbusreq1 & ~n3698;
  assign n3708 = ~n2357 & ~n3697;
  assign n3709 = ~i_hbusreq1 & ~n3708;
  assign n3710 = ~n3707 & ~n3709;
  assign n3711 = ~controllable_hmaster0 & ~n3710;
  assign n3712 = ~n3706 & ~n3711;
  assign n3713 = i_hlock0 & ~n3712;
  assign n3714 = ~n2799 & ~n3692;
  assign n3715 = ~i_hbusreq1 & ~n3714;
  assign n3716 = ~n3702 & ~n3715;
  assign n3717 = controllable_hmaster0 & ~n3716;
  assign n3718 = ~controllable_ndecide & n3256;
  assign n3719 = ~n3697 & ~n3718;
  assign n3720 = ~i_hbusreq1 & ~n3719;
  assign n3721 = ~n3707 & ~n3720;
  assign n3722 = ~controllable_hmaster0 & ~n3721;
  assign n3723 = ~n3717 & ~n3722;
  assign n3724 = ~i_hlock0 & ~n3723;
  assign n3725 = ~n3713 & ~n3724;
  assign n3726 = ~i_hbusreq0 & ~n3725;
  assign n3727 = ~n3701 & ~n3726;
  assign n3728 = ~n1899 & n3727;
  assign n3729 = ~n1899 & ~n3728;
  assign n3730 = ~n2960 & ~n3729;
  assign n3731 = ~n3689 & ~n3730;
  assign n3732 = n1980 & ~n3731;
  assign n3733 = ~n2208 & ~n3732;
  assign n3734 = n1974 & ~n3733;
  assign n3735 = ~n2207 & ~n3734;
  assign n3736 = n2042 & ~n3735;
  assign n3737 = ~n3654 & ~n3736;
  assign n3738 = n1962 & ~n3737;
  assign n3739 = n1962 & ~n3738;
  assign n3740 = ~n1956 & ~n3739;
  assign n3741 = ~n3602 & ~n3740;
  assign n3742 = n1953 & ~n3741;
  assign n3743 = ~n3480 & ~n3742;
  assign n3744 = ~n1947 & ~n3743;
  assign n3745 = ~n2417 & n2960;
  assign n3746 = ~n1996 & ~n2412;
  assign n3747 = ~i_hlock0 & ~n3746;
  assign n3748 = ~n2667 & ~n3747;
  assign n3749 = i_hbusreq0 & ~n3748;
  assign n3750 = ~n2022 & ~n2412;
  assign n3751 = ~i_hlock0 & ~n3750;
  assign n3752 = ~n2673 & ~n3751;
  assign n3753 = ~i_hbusreq0 & ~n3752;
  assign n3754 = ~n3749 & ~n3753;
  assign n3755 = ~n1899 & ~n3754;
  assign n3756 = ~n1899 & ~n3755;
  assign n3757 = ~n2960 & ~n3756;
  assign n3758 = ~n3745 & ~n3757;
  assign n3759 = n1980 & ~n3758;
  assign n3760 = n1980 & ~n3759;
  assign n3761 = n1974 & ~n3760;
  assign n3762 = n1974 & ~n3761;
  assign n3763 = ~n2042 & ~n3762;
  assign n3764 = ~n2454 & ~n3759;
  assign n3765 = n1974 & ~n3764;
  assign n3766 = ~n2453 & ~n3765;
  assign n3767 = n2042 & ~n3766;
  assign n3768 = ~n3763 & ~n3767;
  assign n3769 = ~n1962 & ~n3768;
  assign n3770 = controllable_hmaster0 & ~n2073;
  assign n3771 = ~n2432 & ~n3770;
  assign n3772 = i_hlock0 & ~n3771;
  assign n3773 = ~n2981 & ~n3772;
  assign n3774 = ~n1899 & ~n3773;
  assign n3775 = ~n1899 & ~n3774;
  assign n3776 = n2960 & ~n3775;
  assign n3777 = ~n2960 & ~n2990;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = n1980 & ~n3778;
  assign n3780 = n1980 & ~n3779;
  assign n3781 = n1974 & ~n3780;
  assign n3782 = n1974 & ~n3781;
  assign n3783 = ~n2042 & ~n3782;
  assign n3784 = controllable_hmaster0 & ~n2731;
  assign n3785 = ~n2468 & ~n3784;
  assign n3786 = i_hlock0 & ~n3785;
  assign n3787 = ~n2727 & ~n3786;
  assign n3788 = ~n1899 & ~n3787;
  assign n3789 = ~n1899 & ~n3788;
  assign n3790 = n2960 & ~n3789;
  assign n3791 = ~n2745 & ~n2960;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = n1980 & ~n3792;
  assign n3794 = ~n2454 & ~n3793;
  assign n3795 = n1974 & ~n3794;
  assign n3796 = ~n2453 & ~n3795;
  assign n3797 = n2042 & ~n3796;
  assign n3798 = ~n3783 & ~n3797;
  assign n3799 = n1962 & ~n3798;
  assign n3800 = ~n3769 & ~n3799;
  assign n3801 = n1956 & ~n3800;
  assign n3802 = controllable_nhgrant0 & ~n3102;
  assign n3803 = controllable_nhgrant0 & ~n3802;
  assign n3804 = controllable_hgrant1 & ~n3803;
  assign n3805 = controllable_hgrant1 & ~n3804;
  assign n3806 = controllable_ndecide & ~n3805;
  assign n3807 = ~n1994 & ~n3806;
  assign n3808 = controllable_hmaster0 & ~n3807;
  assign n3809 = ~n2401 & ~n3808;
  assign n3810 = i_hlock0 & ~n3809;
  assign n3811 = ~n2412 & ~n3808;
  assign n3812 = ~i_hlock0 & ~n3811;
  assign n3813 = ~n3810 & ~n3812;
  assign n3814 = i_hbusreq0 & ~n3813;
  assign n3815 = i_hbusreq1 & ~n3807;
  assign n3816 = controllable_ndecide & ~n3806;
  assign n3817 = ~i_hbusreq1 & ~n3816;
  assign n3818 = ~n3815 & ~n3817;
  assign n3819 = controllable_hmaster0 & ~n3818;
  assign n3820 = ~n2401 & ~n3819;
  assign n3821 = i_hlock0 & ~n3820;
  assign n3822 = ~n2412 & ~n3819;
  assign n3823 = ~i_hlock0 & ~n3822;
  assign n3824 = ~n3821 & ~n3823;
  assign n3825 = ~i_hbusreq0 & ~n3824;
  assign n3826 = ~n3814 & ~n3825;
  assign n3827 = ~n1899 & ~n3826;
  assign n3828 = ~n1899 & ~n3827;
  assign n3829 = ~n2960 & ~n3828;
  assign n3830 = ~n3745 & ~n3829;
  assign n3831 = n1980 & ~n3830;
  assign n3832 = n1980 & ~n3831;
  assign n3833 = n1974 & ~n3832;
  assign n3834 = n1974 & ~n3833;
  assign n3835 = ~n2042 & ~n3834;
  assign n3836 = ~n2454 & ~n3831;
  assign n3837 = n1974 & ~n3836;
  assign n3838 = ~n2453 & ~n3837;
  assign n3839 = n2042 & ~n3838;
  assign n3840 = ~n3835 & ~n3839;
  assign n3841 = ~n1962 & ~n3840;
  assign n3842 = ~n2503 & ~n3770;
  assign n3843 = i_hlock0 & ~n3842;
  assign n3844 = ~n2067 & ~n2507;
  assign n3845 = ~i_hlock0 & ~n3844;
  assign n3846 = ~n3843 & ~n3845;
  assign n3847 = i_hbusreq0 & ~n3846;
  assign n3848 = ~n2516 & ~n3770;
  assign n3849 = i_hlock0 & ~n3848;
  assign n3850 = ~n3845 & ~n3849;
  assign n3851 = ~i_hbusreq0 & ~n3850;
  assign n3852 = ~n3847 & ~n3851;
  assign n3853 = ~n1899 & ~n3852;
  assign n3854 = ~n1899 & ~n3853;
  assign n3855 = n2960 & ~n3854;
  assign n3856 = ~n2047 & ~n3804;
  assign n3857 = controllable_ndecide & ~n3856;
  assign n3858 = ~n1994 & ~n3857;
  assign n3859 = controllable_hmaster0 & ~n3858;
  assign n3860 = ~n2503 & ~n3859;
  assign n3861 = i_hlock0 & ~n3860;
  assign n3862 = ~n2065 & ~n3857;
  assign n3863 = controllable_hmaster0 & ~n3862;
  assign n3864 = ~n2507 & ~n3863;
  assign n3865 = ~i_hlock0 & ~n3864;
  assign n3866 = ~n3861 & ~n3865;
  assign n3867 = i_hbusreq0 & ~n3866;
  assign n3868 = i_hbusreq1 & ~n3858;
  assign n3869 = controllable_ndecide & ~n3857;
  assign n3870 = ~i_hbusreq1 & ~n3869;
  assign n3871 = ~n3868 & ~n3870;
  assign n3872 = controllable_hmaster0 & ~n3871;
  assign n3873 = ~n2516 & ~n3872;
  assign n3874 = i_hlock0 & ~n3873;
  assign n3875 = ~n3865 & ~n3874;
  assign n3876 = ~i_hbusreq0 & ~n3875;
  assign n3877 = ~n3867 & ~n3876;
  assign n3878 = ~n1899 & ~n3877;
  assign n3879 = ~n1899 & ~n3878;
  assign n3880 = ~n2960 & ~n3879;
  assign n3881 = ~n3855 & ~n3880;
  assign n3882 = n1980 & ~n3881;
  assign n3883 = n1980 & ~n3882;
  assign n3884 = n1974 & ~n3883;
  assign n3885 = n1974 & ~n3884;
  assign n3886 = ~n2042 & ~n3885;
  assign n3887 = ~n2531 & ~n2692;
  assign n3888 = controllable_hmaster0 & ~n3887;
  assign n3889 = ~n2540 & ~n3888;
  assign n3890 = i_hlock0 & ~n3889;
  assign n3891 = ~n2535 & ~n2723;
  assign n3892 = ~controllable_hmaster0 & ~n3891;
  assign n3893 = ~n2717 & ~n3892;
  assign n3894 = ~i_hlock0 & ~n3893;
  assign n3895 = ~n3890 & ~n3894;
  assign n3896 = i_hbusreq0 & ~n3895;
  assign n3897 = i_hbusreq1 & ~n3887;
  assign n3898 = ~n2732 & ~n3897;
  assign n3899 = controllable_hmaster0 & ~n3898;
  assign n3900 = ~n2557 & ~n3899;
  assign n3901 = i_hlock0 & ~n3900;
  assign n3902 = ~n3894 & ~n3901;
  assign n3903 = ~i_hbusreq0 & ~n3902;
  assign n3904 = ~n3896 & ~n3903;
  assign n3905 = ~n1899 & ~n3904;
  assign n3906 = ~n1899 & ~n3905;
  assign n3907 = n2960 & ~n3906;
  assign n3908 = controllable_nhgrant0 & ~n3243;
  assign n3909 = controllable_nhgrant0 & ~n3908;
  assign n3910 = controllable_hgrant1 & ~n3909;
  assign n3911 = ~n2690 & ~n3910;
  assign n3912 = controllable_ndecide & ~n3911;
  assign n3913 = ~i_hlock1 & ~n3256;
  assign n3914 = ~i_hlock1 & ~n3913;
  assign n3915 = ~controllable_ndecide & ~n3914;
  assign n3916 = ~n3912 & ~n3915;
  assign n3917 = controllable_hmaster0 & ~n3916;
  assign n3918 = ~controllable_hmaster0 & ~n2795;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = i_hlock0 & ~n3919;
  assign n3921 = ~n2715 & ~n3912;
  assign n3922 = controllable_hmaster0 & ~n3921;
  assign n3923 = ~controllable_hmaster0 & ~n2802;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~i_hlock0 & ~n3924;
  assign n3926 = ~n3920 & ~n3925;
  assign n3927 = i_hbusreq0 & ~n3926;
  assign n3928 = i_hbusreq1 & ~n3916;
  assign n3929 = controllable_ndecide & ~n3912;
  assign n3930 = ~i_hbusreq1 & ~n3929;
  assign n3931 = ~n3928 & ~n3930;
  assign n3932 = controllable_hmaster0 & ~n3931;
  assign n3933 = ~controllable_hmaster0 & ~n2815;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = i_hlock0 & ~n3934;
  assign n3936 = ~n3925 & ~n3935;
  assign n3937 = ~i_hbusreq0 & ~n3936;
  assign n3938 = ~n3927 & ~n3937;
  assign n3939 = ~n1899 & ~n3938;
  assign n3940 = ~n1899 & ~n3939;
  assign n3941 = ~n2960 & ~n3940;
  assign n3942 = ~n3907 & ~n3941;
  assign n3943 = n1980 & ~n3942;
  assign n3944 = ~n2454 & ~n3943;
  assign n3945 = n1974 & ~n3944;
  assign n3946 = ~n2453 & ~n3945;
  assign n3947 = n2042 & ~n3946;
  assign n3948 = ~n3886 & ~n3947;
  assign n3949 = n1962 & ~n3948;
  assign n3950 = ~n3841 & ~n3949;
  assign n3951 = ~n1956 & ~n3950;
  assign n3952 = ~n3801 & ~n3951;
  assign n3953 = ~n1953 & ~n3952;
  assign n3954 = ~n2267 & ~n2629;
  assign n3955 = i_hlock0 & ~n3954;
  assign n3956 = ~n2271 & ~n2629;
  assign n3957 = ~i_hlock0 & ~n3956;
  assign n3958 = ~n3955 & ~n3957;
  assign n3959 = ~n1899 & ~n3958;
  assign n3960 = ~n1899 & ~n3959;
  assign n3961 = n2960 & ~n3960;
  assign n3962 = ~n2262 & ~n3804;
  assign n3963 = controllable_ndecide & ~n3962;
  assign n3964 = ~n2265 & ~n3963;
  assign n3965 = controllable_hmaster0 & ~n3964;
  assign n3966 = ~n2629 & ~n3965;
  assign n3967 = i_hlock0 & ~n3966;
  assign n3968 = ~n2065 & ~n3963;
  assign n3969 = controllable_hmaster0 & ~n3968;
  assign n3970 = ~n2629 & ~n3969;
  assign n3971 = ~i_hlock0 & ~n3970;
  assign n3972 = ~n3967 & ~n3971;
  assign n3973 = ~n1899 & ~n3972;
  assign n3974 = ~n1899 & ~n3973;
  assign n3975 = ~n2960 & ~n3974;
  assign n3976 = ~n3961 & ~n3975;
  assign n3977 = n1980 & ~n3976;
  assign n3978 = n1980 & ~n3977;
  assign n3979 = n1974 & ~n3978;
  assign n3980 = n1974 & ~n3979;
  assign n3981 = ~n2042 & ~n3980;
  assign n3982 = ~n2639 & ~n2848;
  assign n3983 = ~controllable_hmaster0 & ~n3982;
  assign n3984 = ~n2846 & ~n3983;
  assign n3985 = i_hlock0 & ~n3984;
  assign n3986 = ~n2639 & ~n2723;
  assign n3987 = ~controllable_hmaster0 & ~n3986;
  assign n3988 = ~n2854 & ~n3987;
  assign n3989 = ~i_hlock0 & ~n3988;
  assign n3990 = ~n3985 & ~n3989;
  assign n3991 = ~n1899 & ~n3990;
  assign n3992 = ~n1899 & ~n3991;
  assign n3993 = n2960 & ~n3992;
  assign n3994 = ~n2838 & ~n3910;
  assign n3995 = controllable_ndecide & ~n3994;
  assign n3996 = ~n2844 & ~n3995;
  assign n3997 = controllable_hmaster0 & ~n3996;
  assign n3998 = controllable_nhgrant0 & n1983;
  assign n3999 = controllable_nhgrant0 & ~n3998;
  assign n4000 = controllable_hgrant1 & ~n3999;
  assign n4001 = ~n2593 & ~n4000;
  assign n4002 = controllable_ndecide & ~n4001;
  assign n4003 = ~n2848 & ~n4002;
  assign n4004 = ~controllable_hmaster0 & ~n4003;
  assign n4005 = ~n3997 & ~n4004;
  assign n4006 = i_hlock0 & ~n4005;
  assign n4007 = ~n2715 & ~n3995;
  assign n4008 = controllable_hmaster0 & ~n4007;
  assign n4009 = ~n2723 & ~n4002;
  assign n4010 = ~controllable_hmaster0 & ~n4009;
  assign n4011 = ~n4008 & ~n4010;
  assign n4012 = ~i_hlock0 & ~n4011;
  assign n4013 = ~n4006 & ~n4012;
  assign n4014 = ~n1899 & ~n4013;
  assign n4015 = ~n1899 & ~n4014;
  assign n4016 = ~n2960 & ~n4015;
  assign n4017 = ~n3993 & ~n4016;
  assign n4018 = n1980 & ~n4017;
  assign n4019 = ~n2454 & ~n4018;
  assign n4020 = n1974 & ~n4019;
  assign n4021 = ~n2453 & ~n4020;
  assign n4022 = n2042 & ~n4021;
  assign n4023 = ~n3981 & ~n4022;
  assign n4024 = n1962 & ~n4023;
  assign n4025 = n1962 & ~n4024;
  assign n4026 = ~n1956 & ~n4025;
  assign n4027 = ~n3066 & ~n4026;
  assign n4028 = n1953 & ~n4027;
  assign n4029 = ~n3953 & ~n4028;
  assign n4030 = n1947 & ~n4029;
  assign n4031 = ~n3744 & ~n4030;
  assign n4032 = ~n1944 & ~n4031;
  assign n4033 = ~n1962 & ~n2684;
  assign n4034 = ~n2750 & ~n2995;
  assign n4035 = n1962 & ~n4034;
  assign n4036 = ~n4033 & ~n4035;
  assign n4037 = n1956 & ~n4036;
  assign n4038 = ~n1962 & ~n2775;
  assign n4039 = ~n2828 & ~n3034;
  assign n4040 = n1962 & ~n4039;
  assign n4041 = ~n4038 & ~n4040;
  assign n4042 = ~n1956 & ~n4041;
  assign n4043 = ~n4037 & ~n4042;
  assign n4044 = ~n1953 & ~n4043;
  assign n4045 = ~n2866 & ~n3058;
  assign n4046 = n1962 & ~n4045;
  assign n4047 = n1962 & ~n4046;
  assign n4048 = n1956 & ~n4047;
  assign n4049 = ~n2949 & ~n3082;
  assign n4050 = n1962 & ~n4049;
  assign n4051 = n1962 & ~n4050;
  assign n4052 = ~n1956 & ~n4051;
  assign n4053 = ~n4048 & ~n4052;
  assign n4054 = n1953 & ~n4053;
  assign n4055 = ~n4044 & ~n4054;
  assign n4056 = ~n1947 & ~n4055;
  assign n4057 = ~n2042 & ~n2684;
  assign n4058 = ~n2454 & ~n2681;
  assign n4059 = n1974 & ~n4058;
  assign n4060 = ~n2453 & ~n4059;
  assign n4061 = n2042 & ~n4060;
  assign n4062 = ~n4057 & ~n4061;
  assign n4063 = ~n1962 & ~n4062;
  assign n4064 = ~n3001 & ~n4063;
  assign n4065 = n1956 & ~n4064;
  assign n4066 = ~n2042 & ~n2775;
  assign n4067 = n2042 & ~n2771;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n1962 & ~n4068;
  assign n4070 = ~n3042 & ~n4069;
  assign n4071 = ~n1956 & ~n4070;
  assign n4072 = ~n4065 & ~n4071;
  assign n4073 = ~n1953 & ~n4072;
  assign n4074 = ~n3092 & ~n4073;
  assign n4075 = n1947 & ~n4074;
  assign n4076 = ~n4056 & ~n4075;
  assign n4077 = n1944 & ~n4076;
  assign n4078 = ~n4032 & ~n4077;
  assign n4079 = n1942 & ~n4078;
  assign n4080 = n2960 & ~n3126;
  assign n4081 = ~n2961 & ~n4080;
  assign n4082 = n1980 & ~n4081;
  assign n4083 = n1980 & ~n4082;
  assign n4084 = n1974 & ~n4083;
  assign n4085 = n1974 & ~n4084;
  assign n4086 = ~n2042 & ~n4085;
  assign n4087 = ~controllable_hmaster0 & ~n3109;
  assign n4088 = i_hlock0 & ~n4087;
  assign n4089 = ~controllable_hmaster0 & ~n3113;
  assign n4090 = ~i_hlock0 & ~n4089;
  assign n4091 = ~n4088 & ~n4090;
  assign n4092 = ~n1899 & ~n4091;
  assign n4093 = ~n1899 & ~n4092;
  assign n4094 = ~n1980 & ~n4093;
  assign n4095 = ~n1980 & ~n4094;
  assign n4096 = ~n1974 & ~n4095;
  assign n4097 = ~n4084 & ~n4096;
  assign n4098 = n2042 & ~n4097;
  assign n4099 = ~n4086 & ~n4098;
  assign n4100 = ~n1962 & ~n4099;
  assign n4101 = ~controllable_locked & n2000;
  assign n4102 = ~controllable_locked & ~n4101;
  assign n4103 = ~controllable_nhgrant0 & ~n4102;
  assign n4104 = ~controllable_nhgrant0 & ~n4103;
  assign n4105 = ~controllable_hgrant1 & ~n4104;
  assign n4106 = ~controllable_hgrant1 & ~n4105;
  assign n4107 = controllable_ndecide & ~n4106;
  assign n4108 = ~n3136 & ~n4107;
  assign n4109 = ~controllable_hmaster0 & ~n4108;
  assign n4110 = ~n2051 & ~n4109;
  assign n4111 = i_hlock0 & ~n4110;
  assign n4112 = ~n2440 & ~n4107;
  assign n4113 = ~controllable_hmaster0 & ~n4112;
  assign n4114 = ~n2067 & ~n4113;
  assign n4115 = ~i_hlock0 & ~n4114;
  assign n4116 = ~n4111 & ~n4115;
  assign n4117 = i_hbusreq0 & ~n4116;
  assign n4118 = i_hbusreq1 & ~n4108;
  assign n4119 = controllable_ndecide & ~n4107;
  assign n4120 = ~i_hbusreq1 & ~n4119;
  assign n4121 = ~n4118 & ~n4120;
  assign n4122 = ~controllable_hmaster0 & ~n4121;
  assign n4123 = ~n2076 & ~n4122;
  assign n4124 = i_hlock0 & ~n4123;
  assign n4125 = ~n4115 & ~n4124;
  assign n4126 = ~i_hbusreq0 & ~n4125;
  assign n4127 = ~n4117 & ~n4126;
  assign n4128 = ~n1899 & ~n4127;
  assign n4129 = ~n1899 & ~n4128;
  assign n4130 = n2960 & ~n4129;
  assign n4131 = ~n3777 & ~n4130;
  assign n4132 = n1980 & ~n4131;
  assign n4133 = n1980 & ~n4132;
  assign n4134 = n1974 & ~n4133;
  assign n4135 = n1974 & ~n4134;
  assign n4136 = ~n2042 & ~n4135;
  assign n4137 = ~n2692 & ~n3203;
  assign n4138 = ~controllable_hmaster0 & ~n4137;
  assign n4139 = ~n2694 & ~n4138;
  assign n4140 = i_hlock0 & ~n4139;
  assign n4141 = ~n2692 & ~n2723;
  assign n4142 = ~controllable_hmaster0 & ~n4141;
  assign n4143 = ~n2717 & ~n4142;
  assign n4144 = ~i_hlock0 & ~n4143;
  assign n4145 = ~n4140 & ~n4144;
  assign n4146 = i_hbusreq0 & ~n4145;
  assign n4147 = i_hbusreq1 & ~n4137;
  assign n4148 = ~n2732 & ~n4147;
  assign n4149 = ~controllable_hmaster0 & ~n4148;
  assign n4150 = ~n2734 & ~n4149;
  assign n4151 = i_hlock0 & ~n4150;
  assign n4152 = ~n4144 & ~n4151;
  assign n4153 = ~i_hbusreq0 & ~n4152;
  assign n4154 = ~n4146 & ~n4153;
  assign n4155 = ~n1899 & ~n4154;
  assign n4156 = ~n1899 & ~n4155;
  assign n4157 = n2960 & ~n4156;
  assign n4158 = ~n3791 & ~n4157;
  assign n4159 = n1980 & ~n4158;
  assign n4160 = n1980 & ~n4159;
  assign n4161 = n1974 & ~n4160;
  assign n4162 = ~n4096 & ~n4161;
  assign n4163 = n2042 & ~n4162;
  assign n4164 = ~n4136 & ~n4163;
  assign n4165 = n1962 & ~n4164;
  assign n4166 = ~n4100 & ~n4165;
  assign n4167 = n1956 & ~n4166;
  assign n4168 = n2960 & ~n3314;
  assign n4169 = ~n3004 & ~n4168;
  assign n4170 = n1980 & ~n4169;
  assign n4171 = n1980 & ~n4170;
  assign n4172 = n1974 & ~n4171;
  assign n4173 = n1974 & ~n4172;
  assign n4174 = ~n2042 & ~n4173;
  assign n4175 = ~n1980 & ~n3314;
  assign n4176 = ~n2166 & ~n4175;
  assign n4177 = ~n1974 & ~n4176;
  assign n4178 = ~n2208 & ~n4170;
  assign n4179 = n1974 & ~n4178;
  assign n4180 = ~n4177 & ~n4179;
  assign n4181 = n2042 & ~n4180;
  assign n4182 = ~n4174 & ~n4181;
  assign n4183 = ~n1962 & ~n4182;
  assign n4184 = ~n2495 & ~n4105;
  assign n4185 = controllable_ndecide & ~n4184;
  assign n4186 = ~n3142 & ~n4185;
  assign n4187 = ~controllable_hmaster0 & n4186;
  assign n4188 = ~n2184 & ~n4187;
  assign n4189 = i_hlock0 & ~n4188;
  assign n4190 = ~n2440 & ~n4185;
  assign n4191 = ~controllable_hmaster0 & n4190;
  assign n4192 = ~n2188 & ~n4191;
  assign n4193 = ~i_hlock0 & ~n4192;
  assign n4194 = ~n4189 & ~n4193;
  assign n4195 = i_hbusreq0 & ~n4194;
  assign n4196 = i_hbusreq1 & ~n4186;
  assign n4197 = controllable_ndecide & ~n4185;
  assign n4198 = ~i_hbusreq1 & ~n4197;
  assign n4199 = ~n4196 & ~n4198;
  assign n4200 = ~controllable_hmaster0 & n4199;
  assign n4201 = ~n2195 & ~n4200;
  assign n4202 = i_hlock0 & ~n4201;
  assign n4203 = ~n4193 & ~n4202;
  assign n4204 = ~i_hbusreq0 & ~n4203;
  assign n4205 = ~n4195 & ~n4204;
  assign n4206 = ~n1899 & n4205;
  assign n4207 = ~n1899 & ~n4206;
  assign n4208 = n2960 & ~n4207;
  assign n4209 = ~n2960 & ~n3029;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = n1980 & ~n4210;
  assign n4212 = n1980 & ~n4211;
  assign n4213 = n1974 & ~n4212;
  assign n4214 = n1974 & ~n4213;
  assign n4215 = ~n2042 & ~n4214;
  assign n4216 = ~n2690 & ~n2789;
  assign n4217 = controllable_ndecide & ~n4216;
  assign n4218 = ~n3396 & ~n4217;
  assign n4219 = ~controllable_hmaster0 & n4218;
  assign n4220 = ~n2786 & ~n4219;
  assign n4221 = i_hlock0 & ~n4220;
  assign n4222 = ~n2723 & ~n4217;
  assign n4223 = ~controllable_hmaster0 & n4222;
  assign n4224 = ~n2801 & ~n4223;
  assign n4225 = ~i_hlock0 & ~n4224;
  assign n4226 = ~n4221 & ~n4225;
  assign n4227 = i_hbusreq0 & ~n4226;
  assign n4228 = i_hbusreq1 & ~n4218;
  assign n4229 = controllable_ndecide & ~n4217;
  assign n4230 = ~i_hbusreq1 & ~n4229;
  assign n4231 = ~n4228 & ~n4230;
  assign n4232 = ~controllable_hmaster0 & n4231;
  assign n4233 = ~n2811 & ~n4232;
  assign n4234 = i_hlock0 & ~n4233;
  assign n4235 = ~n4225 & ~n4234;
  assign n4236 = ~i_hbusreq0 & ~n4235;
  assign n4237 = ~n4227 & ~n4236;
  assign n4238 = ~n1899 & n4237;
  assign n4239 = ~n1899 & ~n4238;
  assign n4240 = n2960 & ~n4239;
  assign n4241 = ~n2823 & ~n2960;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = n1980 & ~n4242;
  assign n4244 = ~n2208 & ~n4243;
  assign n4245 = n1974 & ~n4244;
  assign n4246 = ~n4177 & ~n4245;
  assign n4247 = n2042 & ~n4246;
  assign n4248 = ~n4215 & ~n4247;
  assign n4249 = n1962 & ~n4248;
  assign n4250 = ~n4183 & ~n4249;
  assign n4251 = ~n1956 & ~n4250;
  assign n4252 = ~n4167 & ~n4251;
  assign n4253 = ~n1953 & ~n4252;
  assign n4254 = ~n3171 & ~n4107;
  assign n4255 = ~controllable_hmaster0 & ~n4254;
  assign n4256 = ~n2267 & ~n4255;
  assign n4257 = i_hlock0 & ~n4256;
  assign n4258 = ~n2271 & ~n4113;
  assign n4259 = ~i_hlock0 & ~n4258;
  assign n4260 = ~n4257 & ~n4259;
  assign n4261 = i_hbusreq0 & ~n4260;
  assign n4262 = i_hbusreq1 & ~n4254;
  assign n4263 = ~n4120 & ~n4262;
  assign n4264 = ~controllable_hmaster0 & ~n4263;
  assign n4265 = ~n2267 & ~n4264;
  assign n4266 = i_hlock0 & ~n4265;
  assign n4267 = ~n4259 & ~n4266;
  assign n4268 = ~i_hbusreq0 & ~n4267;
  assign n4269 = ~n4261 & ~n4268;
  assign n4270 = ~n1899 & ~n4269;
  assign n4271 = ~n1899 & ~n4270;
  assign n4272 = n1980 & ~n4271;
  assign n4273 = n1980 & ~n4272;
  assign n4274 = n1974 & ~n4273;
  assign n4275 = n1974 & ~n4274;
  assign n4276 = ~n2042 & ~n4275;
  assign n4277 = ~n2692 & ~n3259;
  assign n4278 = ~controllable_hmaster0 & ~n4277;
  assign n4279 = ~n3565 & ~n4278;
  assign n4280 = i_hlock0 & ~n4279;
  assign n4281 = ~n3569 & ~n4142;
  assign n4282 = ~i_hlock0 & ~n4281;
  assign n4283 = ~n4280 & ~n4282;
  assign n4284 = i_hbusreq0 & ~n4283;
  assign n4285 = i_hbusreq1 & ~n4277;
  assign n4286 = ~n2120 & ~n2692;
  assign n4287 = ~i_hbusreq1 & ~n4286;
  assign n4288 = ~n4285 & ~n4287;
  assign n4289 = ~controllable_hmaster0 & ~n4288;
  assign n4290 = ~n3578 & ~n4289;
  assign n4291 = i_hlock0 & ~n4290;
  assign n4292 = ~n4282 & ~n4291;
  assign n4293 = ~i_hbusreq0 & ~n4292;
  assign n4294 = ~n4284 & ~n4293;
  assign n4295 = ~n1899 & ~n4294;
  assign n4296 = ~n1899 & ~n4295;
  assign n4297 = n1980 & ~n4296;
  assign n4298 = n1980 & ~n4297;
  assign n4299 = n1974 & ~n4298;
  assign n4300 = ~n4096 & ~n4299;
  assign n4301 = n2042 & ~n4300;
  assign n4302 = ~n4276 & ~n4301;
  assign n4303 = n1962 & ~n4302;
  assign n4304 = n1962 & ~n4303;
  assign n4305 = n1956 & ~n4304;
  assign n4306 = ~n2625 & ~n4105;
  assign n4307 = controllable_ndecide & ~n4306;
  assign n4308 = ~n3171 & ~n4307;
  assign n4309 = ~controllable_hmaster0 & n4308;
  assign n4310 = ~n2308 & ~n4309;
  assign n4311 = i_hlock0 & ~n4310;
  assign n4312 = ~n2440 & ~n4307;
  assign n4313 = ~controllable_hmaster0 & n4312;
  assign n4314 = ~n2308 & ~n4313;
  assign n4315 = ~i_hlock0 & ~n4314;
  assign n4316 = ~n4311 & ~n4315;
  assign n4317 = i_hbusreq0 & ~n4316;
  assign n4318 = i_hbusreq1 & ~n4308;
  assign n4319 = controllable_ndecide & ~n4307;
  assign n4320 = ~i_hbusreq1 & ~n4319;
  assign n4321 = ~n4318 & ~n4320;
  assign n4322 = ~controllable_hmaster0 & n4321;
  assign n4323 = ~n2315 & ~n4322;
  assign n4324 = i_hlock0 & ~n4323;
  assign n4325 = ~n4315 & ~n4324;
  assign n4326 = ~i_hbusreq0 & ~n4325;
  assign n4327 = ~n4317 & ~n4326;
  assign n4328 = ~n1899 & n4327;
  assign n4329 = ~n1899 & ~n4328;
  assign n4330 = n1980 & ~n4329;
  assign n4331 = n1980 & ~n4330;
  assign n4332 = n1974 & ~n4331;
  assign n4333 = n1974 & ~n4332;
  assign n4334 = ~n2042 & ~n4333;
  assign n4335 = ~n2779 & ~n2884;
  assign n4336 = controllable_ndecide & ~n4335;
  assign n4337 = ~n3665 & ~n4336;
  assign n4338 = ~controllable_hmaster0 & ~n4337;
  assign n4339 = ~n3694 & ~n4338;
  assign n4340 = i_hlock0 & ~n4339;
  assign n4341 = ~n2906 & ~n4336;
  assign n4342 = ~controllable_hmaster0 & ~n4341;
  assign n4343 = ~n3694 & ~n4342;
  assign n4344 = ~i_hlock0 & ~n4343;
  assign n4345 = ~n4340 & ~n4344;
  assign n4346 = i_hbusreq0 & ~n4345;
  assign n4347 = i_hbusreq1 & ~n4337;
  assign n4348 = ~n2357 & ~n4336;
  assign n4349 = ~i_hbusreq1 & ~n4348;
  assign n4350 = ~n4347 & ~n4349;
  assign n4351 = ~controllable_hmaster0 & ~n4350;
  assign n4352 = ~n3706 & ~n4351;
  assign n4353 = i_hlock0 & ~n4352;
  assign n4354 = i_hbusreq1 & ~n4341;
  assign n4355 = ~n2933 & ~n4336;
  assign n4356 = ~i_hbusreq1 & ~n4355;
  assign n4357 = ~n4354 & ~n4356;
  assign n4358 = ~controllable_hmaster0 & ~n4357;
  assign n4359 = ~n3717 & ~n4358;
  assign n4360 = ~i_hlock0 & ~n4359;
  assign n4361 = ~n4353 & ~n4360;
  assign n4362 = ~i_hbusreq0 & ~n4361;
  assign n4363 = ~n4346 & ~n4362;
  assign n4364 = ~n1899 & n4363;
  assign n4365 = ~n1899 & ~n4364;
  assign n4366 = n1980 & ~n4365;
  assign n4367 = ~n2208 & ~n4366;
  assign n4368 = n1974 & ~n4367;
  assign n4369 = ~n4177 & ~n4368;
  assign n4370 = n2042 & ~n4369;
  assign n4371 = ~n4334 & ~n4370;
  assign n4372 = n1962 & ~n4371;
  assign n4373 = n1962 & ~n4372;
  assign n4374 = ~n1956 & ~n4373;
  assign n4375 = ~n4305 & ~n4374;
  assign n4376 = n1953 & ~n4375;
  assign n4377 = ~n4253 & ~n4376;
  assign n4378 = ~n1947 & ~n4377;
  assign n4379 = n2960 & ~n3756;
  assign n4380 = ~n2961 & ~n4379;
  assign n4381 = n1980 & ~n4380;
  assign n4382 = n1980 & ~n4381;
  assign n4383 = n1974 & ~n4382;
  assign n4384 = n1974 & ~n4383;
  assign n4385 = ~n2042 & ~n4384;
  assign n4386 = ~n2454 & ~n4381;
  assign n4387 = n1974 & ~n4386;
  assign n4388 = ~n2453 & ~n4387;
  assign n4389 = n2042 & ~n4388;
  assign n4390 = ~n4385 & ~n4389;
  assign n4391 = ~n1962 & ~n4390;
  assign n4392 = ~n3001 & ~n4391;
  assign n4393 = n1956 & ~n4392;
  assign n4394 = n2960 & ~n3828;
  assign n4395 = ~n3004 & ~n4394;
  assign n4396 = n1980 & ~n4395;
  assign n4397 = n1980 & ~n4396;
  assign n4398 = n1974 & ~n4397;
  assign n4399 = n1974 & ~n4398;
  assign n4400 = ~n2042 & ~n4399;
  assign n4401 = ~n1980 & ~n3828;
  assign n4402 = ~n2418 & ~n4401;
  assign n4403 = ~n1974 & ~n4402;
  assign n4404 = ~n2454 & ~n4396;
  assign n4405 = n1974 & ~n4404;
  assign n4406 = ~n4403 & ~n4405;
  assign n4407 = n2042 & ~n4406;
  assign n4408 = ~n4400 & ~n4407;
  assign n4409 = ~n1962 & ~n4408;
  assign n4410 = controllable_nhgrant0 & ~n4102;
  assign n4411 = controllable_nhgrant0 & ~n4410;
  assign n4412 = controllable_hgrant1 & ~n4411;
  assign n4413 = ~n2047 & ~n4412;
  assign n4414 = controllable_ndecide & ~n4413;
  assign n4415 = ~i_hlock1 & n2064;
  assign n4416 = ~i_hlock1 & ~n4415;
  assign n4417 = ~controllable_ndecide & ~n4416;
  assign n4418 = ~n4414 & ~n4417;
  assign n4419 = controllable_hmaster0 & ~n4418;
  assign n4420 = ~n2503 & ~n4419;
  assign n4421 = i_hlock0 & ~n4420;
  assign n4422 = ~n2065 & ~n4414;
  assign n4423 = controllable_hmaster0 & ~n4422;
  assign n4424 = ~n2507 & ~n4423;
  assign n4425 = ~i_hlock0 & ~n4424;
  assign n4426 = ~n4421 & ~n4425;
  assign n4427 = i_hbusreq0 & ~n4426;
  assign n4428 = i_hbusreq1 & ~n4418;
  assign n4429 = controllable_ndecide & ~n4414;
  assign n4430 = ~i_hbusreq1 & ~n4429;
  assign n4431 = ~n4428 & ~n4430;
  assign n4432 = controllable_hmaster0 & ~n4431;
  assign n4433 = ~n2516 & ~n4432;
  assign n4434 = i_hlock0 & ~n4433;
  assign n4435 = ~n4425 & ~n4434;
  assign n4436 = ~i_hbusreq0 & ~n4435;
  assign n4437 = ~n4427 & ~n4436;
  assign n4438 = ~n1899 & ~n4437;
  assign n4439 = ~n1899 & ~n4438;
  assign n4440 = n2960 & ~n4439;
  assign n4441 = ~n4209 & ~n4440;
  assign n4442 = n1980 & ~n4441;
  assign n4443 = n1980 & ~n4442;
  assign n4444 = n1974 & ~n4443;
  assign n4445 = n1974 & ~n4444;
  assign n4446 = ~n2042 & ~n4445;
  assign n4447 = ~i_hlock1 & n2714;
  assign n4448 = ~i_hlock1 & ~n4447;
  assign n4449 = ~controllable_ndecide & ~n4448;
  assign n4450 = ~n4217 & ~n4449;
  assign n4451 = controllable_hmaster0 & ~n4450;
  assign n4452 = ~n3918 & ~n4451;
  assign n4453 = i_hlock0 & ~n4452;
  assign n4454 = ~n2715 & ~n4217;
  assign n4455 = controllable_hmaster0 & ~n4454;
  assign n4456 = ~n3923 & ~n4455;
  assign n4457 = ~i_hlock0 & ~n4456;
  assign n4458 = ~n4453 & ~n4457;
  assign n4459 = i_hbusreq0 & ~n4458;
  assign n4460 = i_hbusreq1 & ~n4450;
  assign n4461 = ~n4230 & ~n4460;
  assign n4462 = controllable_hmaster0 & ~n4461;
  assign n4463 = ~n3933 & ~n4462;
  assign n4464 = i_hlock0 & ~n4463;
  assign n4465 = ~n4457 & ~n4464;
  assign n4466 = ~i_hbusreq0 & ~n4465;
  assign n4467 = ~n4459 & ~n4466;
  assign n4468 = ~n1899 & ~n4467;
  assign n4469 = ~n1899 & ~n4468;
  assign n4470 = n2960 & ~n4469;
  assign n4471 = ~n4241 & ~n4470;
  assign n4472 = n1980 & ~n4471;
  assign n4473 = ~n2454 & ~n4472;
  assign n4474 = n1974 & ~n4473;
  assign n4475 = ~n4403 & ~n4474;
  assign n4476 = n2042 & ~n4475;
  assign n4477 = ~n4446 & ~n4476;
  assign n4478 = n1962 & ~n4477;
  assign n4479 = ~n4409 & ~n4478;
  assign n4480 = ~n1956 & ~n4479;
  assign n4481 = ~n4393 & ~n4480;
  assign n4482 = ~n1953 & ~n4481;
  assign n4483 = ~n2262 & ~n4412;
  assign n4484 = controllable_ndecide & ~n4483;
  assign n4485 = i_hlock1 & ~n1991;
  assign n4486 = ~n4415 & ~n4485;
  assign n4487 = ~controllable_ndecide & ~n4486;
  assign n4488 = ~n4484 & ~n4487;
  assign n4489 = controllable_hmaster0 & ~n4488;
  assign n4490 = ~n2629 & ~n4489;
  assign n4491 = i_hlock0 & ~n4490;
  assign n4492 = ~n2065 & ~n4484;
  assign n4493 = controllable_hmaster0 & ~n4492;
  assign n4494 = ~n2629 & ~n4493;
  assign n4495 = ~i_hlock0 & ~n4494;
  assign n4496 = ~n4491 & ~n4495;
  assign n4497 = i_hbusreq0 & ~n4496;
  assign n4498 = i_hbusreq1 & ~n4488;
  assign n4499 = ~n2265 & ~n4484;
  assign n4500 = ~i_hbusreq1 & ~n4499;
  assign n4501 = ~n4498 & ~n4500;
  assign n4502 = controllable_hmaster0 & ~n4501;
  assign n4503 = ~n2629 & ~n4502;
  assign n4504 = i_hlock0 & ~n4503;
  assign n4505 = ~n4495 & ~n4504;
  assign n4506 = ~i_hbusreq0 & ~n4505;
  assign n4507 = ~n4497 & ~n4506;
  assign n4508 = ~n1899 & ~n4507;
  assign n4509 = ~n1899 & ~n4508;
  assign n4510 = n1980 & ~n4509;
  assign n4511 = n1980 & ~n4510;
  assign n4512 = n1974 & ~n4511;
  assign n4513 = n1974 & ~n4512;
  assign n4514 = ~n2042 & ~n4513;
  assign n4515 = ~n2789 & ~n2838;
  assign n4516 = controllable_ndecide & ~n4515;
  assign n4517 = i_hlock1 & ~n2843;
  assign n4518 = ~i_hlock1 & n2877;
  assign n4519 = ~n4517 & ~n4518;
  assign n4520 = ~controllable_ndecide & ~n4519;
  assign n4521 = ~n4516 & ~n4520;
  assign n4522 = controllable_hmaster0 & ~n4521;
  assign n4523 = ~n4004 & ~n4522;
  assign n4524 = i_hlock0 & ~n4523;
  assign n4525 = ~n2715 & ~n4516;
  assign n4526 = controllable_hmaster0 & ~n4525;
  assign n4527 = ~n4010 & ~n4526;
  assign n4528 = ~i_hlock0 & ~n4527;
  assign n4529 = ~n4524 & ~n4528;
  assign n4530 = i_hbusreq0 & ~n4529;
  assign n4531 = i_hbusreq1 & ~n4521;
  assign n4532 = ~n2844 & ~n4516;
  assign n4533 = ~i_hbusreq1 & ~n4532;
  assign n4534 = ~n4531 & ~n4533;
  assign n4535 = controllable_hmaster0 & ~n4534;
  assign n4536 = ~n4004 & ~n4535;
  assign n4537 = i_hlock0 & ~n4536;
  assign n4538 = ~n4528 & ~n4537;
  assign n4539 = ~i_hbusreq0 & ~n4538;
  assign n4540 = ~n4530 & ~n4539;
  assign n4541 = ~n1899 & ~n4540;
  assign n4542 = ~n1899 & ~n4541;
  assign n4543 = n1980 & ~n4542;
  assign n4544 = ~n2454 & ~n4543;
  assign n4545 = n1974 & ~n4544;
  assign n4546 = ~n4403 & ~n4545;
  assign n4547 = n2042 & ~n4546;
  assign n4548 = ~n4514 & ~n4547;
  assign n4549 = n1962 & ~n4548;
  assign n4550 = n1962 & ~n4549;
  assign n4551 = ~n1956 & ~n4550;
  assign n4552 = ~n3066 & ~n4551;
  assign n4553 = n1953 & ~n4552;
  assign n4554 = ~n4482 & ~n4553;
  assign n4555 = n1947 & ~n4554;
  assign n4556 = ~n4378 & ~n4555;
  assign n4557 = ~n1944 & ~n4556;
  assign n4558 = ~n1980 & ~n2454;
  assign n4559 = ~n1974 & ~n4558;
  assign n4560 = ~n2683 & ~n4559;
  assign n4561 = n2042 & ~n4560;
  assign n4562 = ~n4057 & ~n4561;
  assign n4563 = ~n1962 & ~n4562;
  assign n4564 = ~n2748 & ~n4559;
  assign n4565 = n2042 & ~n4564;
  assign n4566 = ~n2995 & ~n4565;
  assign n4567 = n1962 & ~n4566;
  assign n4568 = ~n4563 & ~n4567;
  assign n4569 = n1956 & ~n4568;
  assign n4570 = ~n1980 & ~n3036;
  assign n4571 = ~n1974 & ~n4570;
  assign n4572 = ~n2774 & ~n4571;
  assign n4573 = n2042 & ~n4572;
  assign n4574 = ~n4066 & ~n4573;
  assign n4575 = ~n1962 & ~n4574;
  assign n4576 = ~n2826 & ~n4571;
  assign n4577 = n2042 & ~n4576;
  assign n4578 = ~n3034 & ~n4577;
  assign n4579 = n1962 & ~n4578;
  assign n4580 = ~n4575 & ~n4579;
  assign n4581 = ~n1956 & ~n4580;
  assign n4582 = ~n4569 & ~n4581;
  assign n4583 = ~n1953 & ~n4582;
  assign n4584 = ~n2864 & ~n4559;
  assign n4585 = n2042 & ~n4584;
  assign n4586 = ~n3058 & ~n4585;
  assign n4587 = n1962 & ~n4586;
  assign n4588 = n1962 & ~n4587;
  assign n4589 = n1956 & ~n4588;
  assign n4590 = ~n2947 & ~n4571;
  assign n4591 = n2042 & ~n4590;
  assign n4592 = ~n3082 & ~n4591;
  assign n4593 = n1962 & ~n4592;
  assign n4594 = n1962 & ~n4593;
  assign n4595 = ~n1956 & ~n4594;
  assign n4596 = ~n4589 & ~n4595;
  assign n4597 = n1953 & ~n4596;
  assign n4598 = ~n4583 & ~n4597;
  assign n4599 = ~n1947 & ~n4598;
  assign n4600 = ~n4075 & ~n4599;
  assign n4601 = n1944 & ~n4600;
  assign n4602 = ~n4557 & ~n4601;
  assign n4603 = ~n1942 & ~n4602;
  assign n4604 = ~n4079 & ~n4603;
  assign n4605 = ~n1939 & ~n4604;
  assign n4606 = ~n3100 & ~n4605;
  assign n4607 = n1935 & ~n4606;
  assign n4608 = ~n1974 & ~n4093;
  assign n4609 = ~n2683 & ~n4608;
  assign n4610 = n2042 & ~n4609;
  assign n4611 = ~n4057 & ~n4610;
  assign n4612 = ~n1962 & ~n4611;
  assign n4613 = ~n2748 & ~n4608;
  assign n4614 = n2042 & ~n4613;
  assign n4615 = ~n2995 & ~n4614;
  assign n4616 = n1962 & ~n4615;
  assign n4617 = ~n4612 & ~n4616;
  assign n4618 = n1956 & ~n4617;
  assign n4619 = ~n1974 & ~n3314;
  assign n4620 = ~n2208 & ~n2772;
  assign n4621 = n1974 & ~n4620;
  assign n4622 = ~n4619 & ~n4621;
  assign n4623 = n2042 & ~n4622;
  assign n4624 = ~n4066 & ~n4623;
  assign n4625 = ~n1962 & ~n4624;
  assign n4626 = ~n2208 & ~n2824;
  assign n4627 = n1974 & ~n4626;
  assign n4628 = ~n4619 & ~n4627;
  assign n4629 = n2042 & ~n4628;
  assign n4630 = ~n3034 & ~n4629;
  assign n4631 = n1962 & ~n4630;
  assign n4632 = ~n4625 & ~n4631;
  assign n4633 = ~n1956 & ~n4632;
  assign n4634 = ~n4618 & ~n4633;
  assign n4635 = ~n1953 & ~n4634;
  assign n4636 = ~n2267 & ~n4113;
  assign n4637 = i_hlock0 & ~n4636;
  assign n4638 = ~n4259 & ~n4637;
  assign n4639 = i_hbusreq0 & ~n4638;
  assign n4640 = i_hbusreq1 & ~n4112;
  assign n4641 = ~n4120 & ~n4640;
  assign n4642 = ~controllable_hmaster0 & ~n4641;
  assign n4643 = ~n2267 & ~n4642;
  assign n4644 = i_hlock0 & ~n4643;
  assign n4645 = ~n4259 & ~n4644;
  assign n4646 = ~i_hbusreq0 & ~n4645;
  assign n4647 = ~n4639 & ~n4646;
  assign n4648 = ~n1899 & ~n4647;
  assign n4649 = ~n1899 & ~n4648;
  assign n4650 = n2960 & ~n4649;
  assign n4651 = ~n2267 & ~n2442;
  assign n4652 = i_hlock0 & ~n4651;
  assign n4653 = ~n2271 & ~n2442;
  assign n4654 = ~i_hlock0 & ~n4653;
  assign n4655 = ~n4652 & ~n4654;
  assign n4656 = i_hbusreq0 & ~n4655;
  assign n4657 = i_hbusreq1 & ~n2441;
  assign n4658 = ~i_hbusreq1 & ~n2431;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~controllable_hmaster0 & ~n4659;
  assign n4661 = ~n2267 & ~n4660;
  assign n4662 = i_hlock0 & ~n4661;
  assign n4663 = ~n4654 & ~n4662;
  assign n4664 = ~i_hbusreq0 & ~n4663;
  assign n4665 = ~n4656 & ~n4664;
  assign n4666 = ~n1899 & ~n4665;
  assign n4667 = ~n1899 & ~n4666;
  assign n4668 = ~n2960 & ~n4667;
  assign n4669 = ~n4650 & ~n4668;
  assign n4670 = n1980 & ~n4669;
  assign n4671 = n1980 & ~n4670;
  assign n4672 = n1974 & ~n4671;
  assign n4673 = n1974 & ~n4672;
  assign n4674 = ~n2042 & ~n4673;
  assign n4675 = ~n3565 & ~n4142;
  assign n4676 = i_hlock0 & ~n4675;
  assign n4677 = ~n4282 & ~n4676;
  assign n4678 = i_hbusreq0 & ~n4677;
  assign n4679 = i_hbusreq1 & ~n4141;
  assign n4680 = ~n4287 & ~n4679;
  assign n4681 = ~controllable_hmaster0 & ~n4680;
  assign n4682 = ~n3578 & ~n4681;
  assign n4683 = i_hlock0 & ~n4682;
  assign n4684 = ~n4282 & ~n4683;
  assign n4685 = ~i_hbusreq0 & ~n4684;
  assign n4686 = ~n4678 & ~n4685;
  assign n4687 = ~n1899 & ~n4686;
  assign n4688 = ~n1899 & ~n4687;
  assign n4689 = n2960 & ~n4688;
  assign n4690 = ~n2725 & ~n3565;
  assign n4691 = i_hlock0 & ~n4690;
  assign n4692 = ~n2725 & ~n3569;
  assign n4693 = ~i_hlock0 & ~n4692;
  assign n4694 = ~n4691 & ~n4693;
  assign n4695 = i_hbusreq0 & ~n4694;
  assign n4696 = i_hbusreq1 & ~n2724;
  assign n4697 = ~controllable_ndecide & ~n2702;
  assign n4698 = ~n2466 & ~n4697;
  assign n4699 = ~i_hbusreq1 & ~n4698;
  assign n4700 = ~n4696 & ~n4699;
  assign n4701 = ~controllable_hmaster0 & ~n4700;
  assign n4702 = ~n3578 & ~n4701;
  assign n4703 = i_hlock0 & ~n4702;
  assign n4704 = ~n4693 & ~n4703;
  assign n4705 = ~i_hbusreq0 & ~n4704;
  assign n4706 = ~n4695 & ~n4705;
  assign n4707 = ~n1899 & ~n4706;
  assign n4708 = ~n1899 & ~n4707;
  assign n4709 = ~n2960 & ~n4708;
  assign n4710 = ~n4689 & ~n4709;
  assign n4711 = n1980 & ~n4710;
  assign n4712 = n1980 & ~n4711;
  assign n4713 = n1974 & ~n4712;
  assign n4714 = ~n4608 & ~n4713;
  assign n4715 = n2042 & ~n4714;
  assign n4716 = ~n4674 & ~n4715;
  assign n4717 = n1962 & ~n4716;
  assign n4718 = n1962 & ~n4717;
  assign n4719 = n1956 & ~n4718;
  assign n4720 = i_hbusreq0 & ~n4314;
  assign n4721 = i_hbusreq1 & ~n4312;
  assign n4722 = ~n4320 & ~n4721;
  assign n4723 = ~controllable_hmaster0 & n4722;
  assign n4724 = ~n2315 & ~n4723;
  assign n4725 = i_hlock0 & ~n4724;
  assign n4726 = ~n4315 & ~n4725;
  assign n4727 = ~i_hbusreq0 & ~n4726;
  assign n4728 = ~n4720 & ~n4727;
  assign n4729 = ~n1899 & n4728;
  assign n4730 = ~n1899 & ~n4729;
  assign n4731 = n2960 & ~n4730;
  assign n4732 = ~n2428 & ~n2625;
  assign n4733 = controllable_ndecide & ~n4732;
  assign n4734 = ~n2440 & ~n4733;
  assign n4735 = ~controllable_hmaster0 & n4734;
  assign n4736 = ~n2308 & ~n4735;
  assign n4737 = i_hbusreq0 & ~n4736;
  assign n4738 = i_hbusreq1 & ~n4734;
  assign n4739 = ~n2399 & ~n4733;
  assign n4740 = ~i_hbusreq1 & ~n4739;
  assign n4741 = ~n4738 & ~n4740;
  assign n4742 = ~controllable_hmaster0 & n4741;
  assign n4743 = ~n2315 & ~n4742;
  assign n4744 = i_hlock0 & ~n4743;
  assign n4745 = ~i_hlock0 & ~n4736;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~i_hbusreq0 & ~n4746;
  assign n4748 = ~n4737 & ~n4747;
  assign n4749 = ~n1899 & n4748;
  assign n4750 = ~n1899 & ~n4749;
  assign n4751 = ~n2960 & ~n4750;
  assign n4752 = ~n4731 & ~n4751;
  assign n4753 = n1980 & ~n4752;
  assign n4754 = n1980 & ~n4753;
  assign n4755 = n1974 & ~n4754;
  assign n4756 = n1974 & ~n4755;
  assign n4757 = ~n2042 & ~n4756;
  assign n4758 = i_hbusreq0 & ~n4343;
  assign n4759 = ~n4349 & ~n4354;
  assign n4760 = ~controllable_hmaster0 & ~n4759;
  assign n4761 = ~n3706 & ~n4760;
  assign n4762 = i_hlock0 & ~n4761;
  assign n4763 = ~n4360 & ~n4762;
  assign n4764 = ~i_hbusreq0 & ~n4763;
  assign n4765 = ~n4758 & ~n4764;
  assign n4766 = ~n1899 & n4765;
  assign n4767 = ~n1899 & ~n4766;
  assign n4768 = n2960 & ~n4767;
  assign n4769 = ~controllable_hgrant1 & n2463;
  assign n4770 = ~n2884 & ~n4769;
  assign n4771 = controllable_ndecide & ~n4770;
  assign n4772 = ~n2906 & ~n4771;
  assign n4773 = ~controllable_hmaster0 & ~n4772;
  assign n4774 = ~n3694 & ~n4773;
  assign n4775 = i_hbusreq0 & ~n4774;
  assign n4776 = i_hbusreq1 & ~n4772;
  assign n4777 = ~controllable_ndecide & n2702;
  assign n4778 = ~n4771 & ~n4777;
  assign n4779 = ~i_hbusreq1 & ~n4778;
  assign n4780 = ~n4776 & ~n4779;
  assign n4781 = ~controllable_hmaster0 & ~n4780;
  assign n4782 = ~n3706 & ~n4781;
  assign n4783 = i_hlock0 & ~n4782;
  assign n4784 = ~n2933 & ~n4771;
  assign n4785 = ~i_hbusreq1 & ~n4784;
  assign n4786 = ~n4776 & ~n4785;
  assign n4787 = ~controllable_hmaster0 & ~n4786;
  assign n4788 = ~n3717 & ~n4787;
  assign n4789 = ~i_hlock0 & ~n4788;
  assign n4790 = ~n4783 & ~n4789;
  assign n4791 = ~i_hbusreq0 & ~n4790;
  assign n4792 = ~n4775 & ~n4791;
  assign n4793 = ~n1899 & n4792;
  assign n4794 = ~n1899 & ~n4793;
  assign n4795 = ~n2960 & ~n4794;
  assign n4796 = ~n4768 & ~n4795;
  assign n4797 = n1980 & ~n4796;
  assign n4798 = ~n2208 & ~n4797;
  assign n4799 = n1974 & ~n4798;
  assign n4800 = ~n4619 & ~n4799;
  assign n4801 = n2042 & ~n4800;
  assign n4802 = ~n4757 & ~n4801;
  assign n4803 = n1962 & ~n4802;
  assign n4804 = n1962 & ~n4803;
  assign n4805 = ~n1956 & ~n4804;
  assign n4806 = ~n4719 & ~n4805;
  assign n4807 = n1953 & ~n4806;
  assign n4808 = ~n4635 & ~n4807;
  assign n4809 = ~n1947 & ~n4808;
  assign n4810 = ~n1974 & ~n3828;
  assign n4811 = ~n2454 & ~n2772;
  assign n4812 = n1974 & ~n4811;
  assign n4813 = ~n4810 & ~n4812;
  assign n4814 = n2042 & ~n4813;
  assign n4815 = ~n4066 & ~n4814;
  assign n4816 = ~n1962 & ~n4815;
  assign n4817 = ~n2454 & ~n2824;
  assign n4818 = n1974 & ~n4817;
  assign n4819 = ~n4810 & ~n4818;
  assign n4820 = n2042 & ~n4819;
  assign n4821 = ~n3034 & ~n4820;
  assign n4822 = n1962 & ~n4821;
  assign n4823 = ~n4816 & ~n4822;
  assign n4824 = ~n1956 & ~n4823;
  assign n4825 = ~n4065 & ~n4824;
  assign n4826 = ~n1953 & ~n4825;
  assign n4827 = i_hbusreq0 & ~n4494;
  assign n4828 = i_hbusreq1 & ~n4492;
  assign n4829 = ~n4500 & ~n4828;
  assign n4830 = controllable_hmaster0 & ~n4829;
  assign n4831 = ~n2629 & ~n4830;
  assign n4832 = i_hlock0 & ~n4831;
  assign n4833 = ~n4495 & ~n4832;
  assign n4834 = ~i_hbusreq0 & ~n4833;
  assign n4835 = ~n4827 & ~n4834;
  assign n4836 = ~n1899 & ~n4835;
  assign n4837 = ~n1899 & ~n4836;
  assign n4838 = n2960 & ~n4837;
  assign n4839 = ~n2176 & ~n2304;
  assign n4840 = controllable_ndecide & ~n4839;
  assign n4841 = ~n2186 & ~n4840;
  assign n4842 = controllable_hmaster0 & ~n4841;
  assign n4843 = ~n3067 & ~n4842;
  assign n4844 = i_hbusreq0 & ~n4843;
  assign n4845 = i_hbusreq1 & ~n4841;
  assign n4846 = ~n2311 & ~n4840;
  assign n4847 = ~i_hbusreq1 & ~n4846;
  assign n4848 = ~n4845 & ~n4847;
  assign n4849 = controllable_hmaster0 & ~n4848;
  assign n4850 = ~n3067 & ~n4849;
  assign n4851 = i_hlock0 & ~n4850;
  assign n4852 = ~i_hlock0 & ~n4843;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~i_hbusreq0 & ~n4853;
  assign n4855 = ~n4844 & ~n4854;
  assign n4856 = ~n1899 & n4855;
  assign n4857 = ~n1899 & ~n4856;
  assign n4858 = ~n2960 & ~n4857;
  assign n4859 = ~n4838 & ~n4858;
  assign n4860 = n1980 & ~n4859;
  assign n4861 = n1980 & ~n4860;
  assign n4862 = n1974 & ~n4861;
  assign n4863 = n1974 & ~n4862;
  assign n4864 = ~n2042 & ~n4863;
  assign n4865 = ~controllable_ndecide & n2877;
  assign n4866 = ~n4516 & ~n4865;
  assign n4867 = controllable_hmaster0 & ~n4866;
  assign n4868 = ~n4004 & ~n4867;
  assign n4869 = i_hlock0 & ~n4868;
  assign n4870 = ~n4528 & ~n4869;
  assign n4871 = i_hbusreq0 & ~n4870;
  assign n4872 = i_hbusreq1 & ~n4866;
  assign n4873 = ~n4533 & ~n4872;
  assign n4874 = controllable_hmaster0 & ~n4873;
  assign n4875 = ~n4004 & ~n4874;
  assign n4876 = i_hlock0 & ~n4875;
  assign n4877 = ~n4528 & ~n4876;
  assign n4878 = ~i_hbusreq0 & ~n4877;
  assign n4879 = ~n4871 & ~n4878;
  assign n4880 = ~n1899 & ~n4879;
  assign n4881 = ~n1899 & ~n4880;
  assign n4882 = n2960 & ~n4881;
  assign n4883 = ~n2211 & ~n2871;
  assign n4884 = controllable_ndecide & ~n4883;
  assign n4885 = ~controllable_ndecide & ~n2877;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = controllable_hmaster0 & ~n4886;
  assign n4888 = ~controllable_hmaster0 & n4003;
  assign n4889 = ~n4887 & ~n4888;
  assign n4890 = i_hlock0 & ~n4889;
  assign n4891 = ~n2799 & ~n4884;
  assign n4892 = controllable_hmaster0 & ~n4891;
  assign n4893 = ~controllable_hmaster0 & n4009;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = ~i_hlock0 & ~n4894;
  assign n4896 = ~n4890 & ~n4895;
  assign n4897 = i_hbusreq0 & ~n4896;
  assign n4898 = i_hbusreq1 & ~n4886;
  assign n4899 = ~n2914 & ~n4884;
  assign n4900 = ~i_hbusreq1 & ~n4899;
  assign n4901 = ~n4898 & ~n4900;
  assign n4902 = controllable_hmaster0 & ~n4901;
  assign n4903 = ~n4888 & ~n4902;
  assign n4904 = i_hlock0 & ~n4903;
  assign n4905 = ~n4895 & ~n4904;
  assign n4906 = ~i_hbusreq0 & ~n4905;
  assign n4907 = ~n4897 & ~n4906;
  assign n4908 = ~n1899 & n4907;
  assign n4909 = ~n1899 & ~n4908;
  assign n4910 = ~n2960 & ~n4909;
  assign n4911 = ~n4882 & ~n4910;
  assign n4912 = n1980 & ~n4911;
  assign n4913 = ~n2454 & ~n4912;
  assign n4914 = n1974 & ~n4913;
  assign n4915 = ~n4810 & ~n4914;
  assign n4916 = n2042 & ~n4915;
  assign n4917 = ~n4864 & ~n4916;
  assign n4918 = n1962 & ~n4917;
  assign n4919 = n1962 & ~n4918;
  assign n4920 = ~n1956 & ~n4919;
  assign n4921 = ~n3066 & ~n4920;
  assign n4922 = n1953 & ~n4921;
  assign n4923 = ~n4826 & ~n4922;
  assign n4924 = n1947 & ~n4923;
  assign n4925 = ~n4809 & ~n4924;
  assign n4926 = ~n1944 & ~n4925;
  assign n4927 = ~n2453 & ~n2683;
  assign n4928 = n2042 & ~n4927;
  assign n4929 = ~n4057 & ~n4928;
  assign n4930 = ~n1962 & ~n4929;
  assign n4931 = ~n2453 & ~n2748;
  assign n4932 = n2042 & ~n4931;
  assign n4933 = ~n2995 & ~n4932;
  assign n4934 = n1962 & ~n4933;
  assign n4935 = ~n4930 & ~n4934;
  assign n4936 = n1956 & ~n4935;
  assign n4937 = ~n2774 & ~n3035;
  assign n4938 = n2042 & ~n4937;
  assign n4939 = ~n4066 & ~n4938;
  assign n4940 = ~n1962 & ~n4939;
  assign n4941 = ~n2826 & ~n3035;
  assign n4942 = n2042 & ~n4941;
  assign n4943 = ~n3034 & ~n4942;
  assign n4944 = n1962 & ~n4943;
  assign n4945 = ~n4940 & ~n4944;
  assign n4946 = ~n1956 & ~n4945;
  assign n4947 = ~n4936 & ~n4946;
  assign n4948 = ~n1953 & ~n4947;
  assign n4949 = ~n2453 & ~n2864;
  assign n4950 = n2042 & ~n4949;
  assign n4951 = ~n3058 & ~n4950;
  assign n4952 = n1962 & ~n4951;
  assign n4953 = n1962 & ~n4952;
  assign n4954 = n1956 & ~n4953;
  assign n4955 = ~n2947 & ~n3035;
  assign n4956 = n2042 & ~n4955;
  assign n4957 = ~n3082 & ~n4956;
  assign n4958 = n1962 & ~n4957;
  assign n4959 = n1962 & ~n4958;
  assign n4960 = ~n1956 & ~n4959;
  assign n4961 = ~n4954 & ~n4960;
  assign n4962 = n1953 & ~n4961;
  assign n4963 = ~n4948 & ~n4962;
  assign n4964 = ~n1947 & ~n4963;
  assign n4965 = ~n4075 & ~n4964;
  assign n4966 = n1944 & ~n4965;
  assign n4967 = ~n4926 & ~n4966;
  assign n4968 = n1942 & ~n4967;
  assign n4969 = n1980 & ~n4093;
  assign n4970 = ~n2454 & ~n4969;
  assign n4971 = ~n1974 & ~n4970;
  assign n4972 = ~n2681 & ~n4094;
  assign n4973 = n1974 & ~n4972;
  assign n4974 = ~n4971 & ~n4973;
  assign n4975 = n2042 & ~n4974;
  assign n4976 = ~n4057 & ~n4975;
  assign n4977 = ~n1962 & ~n4976;
  assign n4978 = ~n2746 & ~n4094;
  assign n4979 = n1974 & ~n4978;
  assign n4980 = ~n4971 & ~n4979;
  assign n4981 = n2042 & ~n4980;
  assign n4982 = ~n2995 & ~n4981;
  assign n4983 = n1962 & ~n4982;
  assign n4984 = ~n4977 & ~n4983;
  assign n4985 = n1956 & ~n4984;
  assign n4986 = n1980 & ~n3314;
  assign n4987 = ~n3036 & ~n4986;
  assign n4988 = ~n1974 & ~n4987;
  assign n4989 = ~n2772 & ~n4175;
  assign n4990 = n1974 & ~n4989;
  assign n4991 = ~n4988 & ~n4990;
  assign n4992 = n2042 & ~n4991;
  assign n4993 = ~n4066 & ~n4992;
  assign n4994 = ~n1962 & ~n4993;
  assign n4995 = ~n2824 & ~n4175;
  assign n4996 = n1974 & ~n4995;
  assign n4997 = ~n4988 & ~n4996;
  assign n4998 = n2042 & ~n4997;
  assign n4999 = ~n3034 & ~n4998;
  assign n5000 = n1962 & ~n4999;
  assign n5001 = ~n4994 & ~n5000;
  assign n5002 = ~n1956 & ~n5001;
  assign n5003 = ~n4985 & ~n5002;
  assign n5004 = ~n1953 & ~n5003;
  assign n5005 = n1980 & ~n4667;
  assign n5006 = n1980 & ~n5005;
  assign n5007 = n1974 & ~n5006;
  assign n5008 = n1974 & ~n5007;
  assign n5009 = ~n2042 & ~n5008;
  assign n5010 = n1980 & ~n4708;
  assign n5011 = ~n4094 & ~n5010;
  assign n5012 = n1974 & ~n5011;
  assign n5013 = ~n4971 & ~n5012;
  assign n5014 = n2042 & ~n5013;
  assign n5015 = ~n5009 & ~n5014;
  assign n5016 = n1962 & ~n5015;
  assign n5017 = n1962 & ~n5016;
  assign n5018 = n1956 & ~n5017;
  assign n5019 = n1980 & ~n4750;
  assign n5020 = n1980 & ~n5019;
  assign n5021 = n1974 & ~n5020;
  assign n5022 = n1974 & ~n5021;
  assign n5023 = ~n2042 & ~n5022;
  assign n5024 = n1980 & ~n4794;
  assign n5025 = ~n4175 & ~n5024;
  assign n5026 = n1974 & ~n5025;
  assign n5027 = ~n4988 & ~n5026;
  assign n5028 = n2042 & ~n5027;
  assign n5029 = ~n5023 & ~n5028;
  assign n5030 = n1962 & ~n5029;
  assign n5031 = n1962 & ~n5030;
  assign n5032 = ~n1956 & ~n5031;
  assign n5033 = ~n5018 & ~n5032;
  assign n5034 = n1953 & ~n5033;
  assign n5035 = ~n5004 & ~n5034;
  assign n5036 = ~n1947 & ~n5035;
  assign n5037 = n1980 & ~n3828;
  assign n5038 = ~n3036 & ~n5037;
  assign n5039 = ~n1974 & ~n5038;
  assign n5040 = ~n2772 & ~n4401;
  assign n5041 = n1974 & ~n5040;
  assign n5042 = ~n5039 & ~n5041;
  assign n5043 = n2042 & ~n5042;
  assign n5044 = ~n4066 & ~n5043;
  assign n5045 = ~n1962 & ~n5044;
  assign n5046 = ~n2824 & ~n4401;
  assign n5047 = n1974 & ~n5046;
  assign n5048 = ~n5039 & ~n5047;
  assign n5049 = n2042 & ~n5048;
  assign n5050 = ~n3034 & ~n5049;
  assign n5051 = n1962 & ~n5050;
  assign n5052 = ~n5045 & ~n5051;
  assign n5053 = ~n1956 & ~n5052;
  assign n5054 = ~n4065 & ~n5053;
  assign n5055 = ~n1953 & ~n5054;
  assign n5056 = n1980 & ~n4857;
  assign n5057 = n1980 & ~n5056;
  assign n5058 = n1974 & ~n5057;
  assign n5059 = n1974 & ~n5058;
  assign n5060 = ~n2042 & ~n5059;
  assign n5061 = n1980 & ~n4909;
  assign n5062 = ~n4401 & ~n5061;
  assign n5063 = n1974 & ~n5062;
  assign n5064 = ~n5039 & ~n5063;
  assign n5065 = n2042 & ~n5064;
  assign n5066 = ~n5060 & ~n5065;
  assign n5067 = n1962 & ~n5066;
  assign n5068 = n1962 & ~n5067;
  assign n5069 = ~n1956 & ~n5068;
  assign n5070 = ~n3066 & ~n5069;
  assign n5071 = n1953 & ~n5070;
  assign n5072 = ~n5055 & ~n5071;
  assign n5073 = n1947 & ~n5072;
  assign n5074 = ~n5036 & ~n5073;
  assign n5075 = ~n1944 & ~n5074;
  assign n5076 = n1944 & ~n4074;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n1942 & ~n5077;
  assign n5079 = ~n4968 & ~n5078;
  assign n5080 = n1939 & ~n5079;
  assign n5081 = ~n2453 & ~n4973;
  assign n5082 = n2042 & ~n5081;
  assign n5083 = ~n4057 & ~n5082;
  assign n5084 = ~n1962 & ~n5083;
  assign n5085 = ~n2453 & ~n4979;
  assign n5086 = n2042 & ~n5085;
  assign n5087 = ~n2995 & ~n5086;
  assign n5088 = n1962 & ~n5087;
  assign n5089 = ~n5084 & ~n5088;
  assign n5090 = n1956 & ~n5089;
  assign n5091 = ~n3035 & ~n4990;
  assign n5092 = n2042 & ~n5091;
  assign n5093 = ~n4066 & ~n5092;
  assign n5094 = ~n1962 & ~n5093;
  assign n5095 = ~n3035 & ~n4996;
  assign n5096 = n2042 & ~n5095;
  assign n5097 = ~n3034 & ~n5096;
  assign n5098 = n1962 & ~n5097;
  assign n5099 = ~n5094 & ~n5098;
  assign n5100 = ~n1956 & ~n5099;
  assign n5101 = ~n5090 & ~n5100;
  assign n5102 = ~n1953 & ~n5101;
  assign n5103 = ~n2453 & ~n5012;
  assign n5104 = n2042 & ~n5103;
  assign n5105 = ~n5009 & ~n5104;
  assign n5106 = n1962 & ~n5105;
  assign n5107 = n1962 & ~n5106;
  assign n5108 = n1956 & ~n5107;
  assign n5109 = ~n3035 & ~n5026;
  assign n5110 = n2042 & ~n5109;
  assign n5111 = ~n5023 & ~n5110;
  assign n5112 = n1962 & ~n5111;
  assign n5113 = n1962 & ~n5112;
  assign n5114 = ~n1956 & ~n5113;
  assign n5115 = ~n5108 & ~n5114;
  assign n5116 = n1953 & ~n5115;
  assign n5117 = ~n5102 & ~n5116;
  assign n5118 = ~n1947 & ~n5117;
  assign n5119 = ~n3035 & ~n5041;
  assign n5120 = n2042 & ~n5119;
  assign n5121 = ~n4066 & ~n5120;
  assign n5122 = ~n1962 & ~n5121;
  assign n5123 = ~n3035 & ~n5047;
  assign n5124 = n2042 & ~n5123;
  assign n5125 = ~n3034 & ~n5124;
  assign n5126 = n1962 & ~n5125;
  assign n5127 = ~n5122 & ~n5126;
  assign n5128 = ~n1956 & ~n5127;
  assign n5129 = ~n4065 & ~n5128;
  assign n5130 = ~n1953 & ~n5129;
  assign n5131 = ~n3035 & ~n5063;
  assign n5132 = n2042 & ~n5131;
  assign n5133 = ~n5060 & ~n5132;
  assign n5134 = n1962 & ~n5133;
  assign n5135 = n1962 & ~n5134;
  assign n5136 = ~n1956 & ~n5135;
  assign n5137 = ~n3066 & ~n5136;
  assign n5138 = n1953 & ~n5137;
  assign n5139 = ~n5130 & ~n5138;
  assign n5140 = n1947 & ~n5139;
  assign n5141 = ~n5118 & ~n5140;
  assign n5142 = ~n1944 & ~n5141;
  assign n5143 = ~n5076 & ~n5142;
  assign n5144 = n1942 & ~n5143;
  assign n5145 = n2960 & ~n4667;
  assign n5146 = ~n2960 & ~n3053;
  assign n5147 = ~n5145 & ~n5146;
  assign n5148 = n1980 & ~n5147;
  assign n5149 = n1980 & ~n5148;
  assign n5150 = n1974 & ~n5149;
  assign n5151 = n1974 & ~n5150;
  assign n5152 = ~n2042 & ~n5151;
  assign n5153 = controllable_locked & ~n1983;
  assign n5154 = ~controllable_nhgrant0 & n5153;
  assign n5155 = ~controllable_nhgrant0 & ~n5154;
  assign n5156 = ~controllable_hgrant1 & ~n5155;
  assign n5157 = ~controllable_hgrant1 & ~n5156;
  assign n5158 = controllable_ndecide & ~n5157;
  assign n5159 = ~n2848 & ~n5158;
  assign n5160 = ~controllable_hmaster0 & ~n5159;
  assign n5161 = ~n2846 & ~n5160;
  assign n5162 = i_hlock0 & ~n5161;
  assign n5163 = ~n2723 & ~n5158;
  assign n5164 = ~controllable_hmaster0 & ~n5163;
  assign n5165 = ~n2854 & ~n5164;
  assign n5166 = ~i_hlock0 & ~n5165;
  assign n5167 = ~n5162 & ~n5166;
  assign n5168 = i_hbusreq0 & ~n5167;
  assign n5169 = i_hbusreq1 & ~n2845;
  assign n5170 = ~controllable_nhgrant0 & n2697;
  assign n5171 = ~n2405 & ~n5170;
  assign n5172 = ~controllable_hgrant1 & ~n5171;
  assign n5173 = ~n2092 & ~n5172;
  assign n5174 = ~controllable_ndecide & ~n5173;
  assign n5175 = ~n2840 & ~n5174;
  assign n5176 = ~i_hbusreq1 & ~n5175;
  assign n5177 = ~n5169 & ~n5176;
  assign n5178 = controllable_hmaster0 & ~n5177;
  assign n5179 = i_hbusreq1 & ~n5159;
  assign n5180 = ~controllable_nhgrant0 & n2089;
  assign n5181 = ~n2394 & ~n5180;
  assign n5182 = ~controllable_hgrant1 & ~n5181;
  assign n5183 = ~n2701 & ~n5182;
  assign n5184 = ~controllable_ndecide & ~n5183;
  assign n5185 = ~n5158 & ~n5184;
  assign n5186 = ~i_hbusreq1 & ~n5185;
  assign n5187 = ~n5179 & ~n5186;
  assign n5188 = ~controllable_hmaster0 & ~n5187;
  assign n5189 = ~n5178 & ~n5188;
  assign n5190 = i_hlock0 & ~n5189;
  assign n5191 = ~n5166 & ~n5190;
  assign n5192 = ~i_hbusreq0 & ~n5191;
  assign n5193 = ~n5168 & ~n5192;
  assign n5194 = ~n1899 & ~n5193;
  assign n5195 = ~n1899 & ~n5194;
  assign n5196 = n2960 & ~n5195;
  assign n5197 = ~n2861 & ~n2960;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = n1980 & ~n5198;
  assign n5200 = ~n2454 & ~n5199;
  assign n5201 = n1974 & ~n5200;
  assign n5202 = ~n2453 & ~n5201;
  assign n5203 = n2042 & ~n5202;
  assign n5204 = ~n5152 & ~n5203;
  assign n5205 = n1962 & ~n5204;
  assign n5206 = n1962 & ~n5205;
  assign n5207 = n1956 & ~n5206;
  assign n5208 = n2960 & ~n4750;
  assign n5209 = ~n2960 & ~n3077;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = n1980 & ~n5210;
  assign n5212 = n1980 & ~n5211;
  assign n5213 = n1974 & ~n5212;
  assign n5214 = n1974 & ~n5213;
  assign n5215 = ~n2042 & ~n5214;
  assign n5216 = ~controllable_hgrant1 & n5155;
  assign n5217 = ~n2884 & ~n5216;
  assign n5218 = controllable_ndecide & ~n5217;
  assign n5219 = ~n2890 & ~n5218;
  assign n5220 = ~controllable_hmaster0 & ~n5219;
  assign n5221 = ~n2882 & ~n5220;
  assign n5222 = i_hlock0 & ~n5221;
  assign n5223 = ~n2906 & ~n5218;
  assign n5224 = ~controllable_hmaster0 & ~n5223;
  assign n5225 = ~n2900 & ~n5224;
  assign n5226 = ~i_hlock0 & ~n5225;
  assign n5227 = ~n5222 & ~n5226;
  assign n5228 = i_hbusreq0 & ~n5227;
  assign n5229 = ~controllable_ndecide & n5173;
  assign n5230 = ~n2873 & ~n5229;
  assign n5231 = ~i_hbusreq1 & ~n5230;
  assign n5232 = ~n2913 & ~n5231;
  assign n5233 = controllable_hmaster0 & ~n5232;
  assign n5234 = i_hbusreq1 & ~n5219;
  assign n5235 = ~controllable_ndecide & n5183;
  assign n5236 = ~n5218 & ~n5235;
  assign n5237 = ~i_hbusreq1 & ~n5236;
  assign n5238 = ~n5234 & ~n5237;
  assign n5239 = ~controllable_hmaster0 & ~n5238;
  assign n5240 = ~n5233 & ~n5239;
  assign n5241 = i_hlock0 & ~n5240;
  assign n5242 = i_hbusreq1 & ~n5223;
  assign n5243 = ~n2933 & ~n5218;
  assign n5244 = ~i_hbusreq1 & ~n5243;
  assign n5245 = ~n5242 & ~n5244;
  assign n5246 = ~controllable_hmaster0 & ~n5245;
  assign n5247 = ~n2931 & ~n5246;
  assign n5248 = ~i_hlock0 & ~n5247;
  assign n5249 = ~n5241 & ~n5248;
  assign n5250 = ~i_hbusreq0 & ~n5249;
  assign n5251 = ~n5228 & ~n5250;
  assign n5252 = ~n1899 & n5251;
  assign n5253 = ~n1899 & ~n5252;
  assign n5254 = n2960 & ~n5253;
  assign n5255 = ~n2944 & ~n2960;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = n1980 & ~n5256;
  assign n5258 = ~n3036 & ~n5257;
  assign n5259 = n1974 & ~n5258;
  assign n5260 = ~n3035 & ~n5259;
  assign n5261 = n2042 & ~n5260;
  assign n5262 = ~n5215 & ~n5261;
  assign n5263 = n1962 & ~n5262;
  assign n5264 = n1962 & ~n5263;
  assign n5265 = ~n1956 & ~n5264;
  assign n5266 = ~n5207 & ~n5265;
  assign n5267 = n1953 & ~n5266;
  assign n5268 = ~n4073 & ~n5267;
  assign n5269 = ~n1947 & ~n5268;
  assign n5270 = n2960 & ~n4857;
  assign n5271 = ~n5209 & ~n5270;
  assign n5272 = n1980 & ~n5271;
  assign n5273 = n1980 & ~n5272;
  assign n5274 = n1974 & ~n5273;
  assign n5275 = n1974 & ~n5274;
  assign n5276 = ~n2042 & ~n5275;
  assign n5277 = controllable_nhgrant0 & ~n5153;
  assign n5278 = controllable_hgrant1 & n5277;
  assign n5279 = ~n2871 & ~n5278;
  assign n5280 = controllable_ndecide & ~n5279;
  assign n5281 = ~n2880 & ~n5280;
  assign n5282 = controllable_hmaster0 & ~n5281;
  assign n5283 = ~n2892 & ~n5282;
  assign n5284 = i_hlock0 & ~n5283;
  assign n5285 = ~n2898 & ~n5280;
  assign n5286 = controllable_hmaster0 & ~n5285;
  assign n5287 = ~n2908 & ~n5286;
  assign n5288 = ~i_hlock0 & ~n5287;
  assign n5289 = ~n5284 & ~n5288;
  assign n5290 = i_hbusreq0 & ~n5289;
  assign n5291 = i_hbusreq1 & ~n5281;
  assign n5292 = ~n2914 & ~n5280;
  assign n5293 = ~i_hbusreq1 & ~n5292;
  assign n5294 = ~n5291 & ~n5293;
  assign n5295 = controllable_hmaster0 & ~n5294;
  assign n5296 = ~n2924 & ~n5295;
  assign n5297 = i_hlock0 & ~n5296;
  assign n5298 = i_hbusreq1 & ~n5285;
  assign n5299 = ~n2799 & ~n5280;
  assign n5300 = ~i_hbusreq1 & ~n5299;
  assign n5301 = ~n5298 & ~n5300;
  assign n5302 = controllable_hmaster0 & ~n5301;
  assign n5303 = ~n2937 & ~n5302;
  assign n5304 = ~i_hlock0 & ~n5303;
  assign n5305 = ~n5297 & ~n5304;
  assign n5306 = ~i_hbusreq0 & ~n5305;
  assign n5307 = ~n5290 & ~n5306;
  assign n5308 = ~n1899 & n5307;
  assign n5309 = ~n1899 & ~n5308;
  assign n5310 = n2960 & ~n5309;
  assign n5311 = ~n5255 & ~n5310;
  assign n5312 = n1980 & ~n5311;
  assign n5313 = ~n3036 & ~n5312;
  assign n5314 = n1974 & ~n5313;
  assign n5315 = ~n3035 & ~n5314;
  assign n5316 = n2042 & ~n5315;
  assign n5317 = ~n5276 & ~n5316;
  assign n5318 = n1962 & ~n5317;
  assign n5319 = n1962 & ~n5318;
  assign n5320 = ~n1956 & ~n5319;
  assign n5321 = ~n3066 & ~n5320;
  assign n5322 = n1953 & ~n5321;
  assign n5323 = ~n4073 & ~n5322;
  assign n5324 = n1947 & ~n5323;
  assign n5325 = ~n5269 & ~n5324;
  assign n5326 = ~n1944 & ~n5325;
  assign n5327 = ~n5076 & ~n5326;
  assign n5328 = ~n1942 & ~n5327;
  assign n5329 = ~n5144 & ~n5328;
  assign n5330 = ~n1939 & ~n5329;
  assign n5331 = ~n5080 & ~n5330;
  assign n5332 = ~n1935 & ~n5331;
  assign n5333 = ~n4607 & ~n5332;
  assign n5334 = n1898 & n5333;
  assign n5335 = n1898 & ~n5334;
  assign inductivity_check  = ~n1893 & n5335;
endmodule


