// Generated using findDep.cpp 
module stmt44_554_604 (v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_15, v_20, v_22, v_24, v_25, v_26, v_29, v_31, v_33, v_34, v_36, v_38, v_40, v_41, v_43, v_45, v_47, v_49, v_51, v_53, v_55, v_58, v_59, v_66, v_68, v_72, v_76, v_78, v_80, v_84, v_91, v_96, v_101, v_107, v_108, v_112, v_115, v_116, v_125, v_130, v_133, v_134, v_141, v_142, v_146, v_150, v_151, v_154, v_158, v_162, v_164, v_166, v_168, v_170, v_171, v_175, v_179, v_181, v_185, v_189, v_194, v_196, v_200, v_202, v_203, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_460, v_465, v_467, v_469, v_470, v_471, v_474, v_476, v_478, v_479, v_481, v_483, v_485, v_486, v_488, v_490, v_492, v_494, v_496, v_498, v_500, v_503, v_504, v_511, v_513, v_517, v_521, v_523, v_525, v_529, v_536, v_541, v_546, v_552, v_553, v_557, v_560, v_561, v_570, v_575, v_578, v_579, v_586, v_587, v_591, v_595, v_596, v_599, v_603, v_607, v_609, v_611, v_613, v_615, v_616, v_620, v_624, v_626, v_630, v_634, v_639, v_641, v_645, o_1);
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_15;
input v_20;
input v_22;
input v_24;
input v_25;
input v_26;
input v_29;
input v_31;
input v_33;
input v_34;
input v_36;
input v_38;
input v_40;
input v_41;
input v_43;
input v_45;
input v_47;
input v_49;
input v_51;
input v_53;
input v_55;
input v_58;
input v_59;
input v_66;
input v_68;
input v_72;
input v_76;
input v_78;
input v_80;
input v_84;
input v_91;
input v_96;
input v_101;
input v_107;
input v_108;
input v_112;
input v_115;
input v_116;
input v_125;
input v_130;
input v_133;
input v_134;
input v_141;
input v_142;
input v_146;
input v_150;
input v_151;
input v_154;
input v_158;
input v_162;
input v_164;
input v_166;
input v_168;
input v_170;
input v_171;
input v_175;
input v_179;
input v_181;
input v_185;
input v_189;
input v_194;
input v_196;
input v_200;
input v_202;
input v_203;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_460;
input v_465;
input v_467;
input v_469;
input v_470;
input v_471;
input v_474;
input v_476;
input v_478;
input v_479;
input v_481;
input v_483;
input v_485;
input v_486;
input v_488;
input v_490;
input v_492;
input v_494;
input v_496;
input v_498;
input v_500;
input v_503;
input v_504;
input v_511;
input v_513;
input v_517;
input v_521;
input v_523;
input v_525;
input v_529;
input v_536;
input v_541;
input v_546;
input v_552;
input v_553;
input v_557;
input v_560;
input v_561;
input v_570;
input v_575;
input v_578;
input v_579;
input v_586;
input v_587;
input v_591;
input v_595;
input v_596;
input v_599;
input v_603;
input v_607;
input v_609;
input v_611;
input v_613;
input v_615;
input v_616;
input v_620;
input v_624;
input v_626;
input v_630;
input v_634;
input v_639;
input v_641;
input v_645;
output o_1;
wire v_1;
wire v_12;
wire v_13;
wire v_14;
wire v_16;
wire v_17;
wire v_18;
wire v_19;
wire v_21;
wire v_23;
wire v_27;
wire v_28;
wire v_30;
wire v_32;
wire v_35;
wire v_37;
wire v_39;
wire v_42;
wire v_44;
wire v_46;
wire v_48;
wire v_50;
wire v_52;
wire v_54;
wire v_56;
wire v_57;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_67;
wire v_69;
wire v_70;
wire v_71;
wire v_73;
wire v_74;
wire v_75;
wire v_77;
wire v_79;
wire v_81;
wire v_82;
wire v_83;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_109;
wire v_110;
wire v_111;
wire v_113;
wire v_114;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_131;
wire v_132;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_143;
wire v_144;
wire v_145;
wire v_147;
wire v_148;
wire v_149;
wire v_152;
wire v_153;
wire v_155;
wire v_156;
wire v_157;
wire v_159;
wire v_160;
wire v_161;
wire v_163;
wire v_165;
wire v_167;
wire v_169;
wire v_172;
wire v_173;
wire v_174;
wire v_176;
wire v_177;
wire v_178;
wire v_180;
wire v_182;
wire v_183;
wire v_184;
wire v_186;
wire v_187;
wire v_188;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_195;
wire v_197;
wire v_198;
wire v_199;
wire v_201;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_457;
wire v_458;
wire v_459;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_466;
wire v_468;
wire v_472;
wire v_473;
wire v_475;
wire v_477;
wire v_480;
wire v_482;
wire v_484;
wire v_487;
wire v_489;
wire v_491;
wire v_493;
wire v_495;
wire v_497;
wire v_499;
wire v_501;
wire v_502;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_512;
wire v_514;
wire v_515;
wire v_516;
wire v_518;
wire v_519;
wire v_520;
wire v_522;
wire v_524;
wire v_526;
wire v_527;
wire v_528;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_554;
wire v_555;
wire v_556;
wire v_558;
wire v_559;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_576;
wire v_577;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_588;
wire v_589;
wire v_590;
wire v_592;
wire v_593;
wire v_594;
wire v_597;
wire v_598;
wire v_600;
wire v_601;
wire v_602;
wire v_604;
wire v_605;
wire v_606;
wire v_608;
wire v_610;
wire v_612;
wire v_614;
wire v_617;
wire v_618;
wire v_619;
wire v_621;
wire v_622;
wire v_623;
wire v_625;
wire v_627;
wire v_628;
wire v_629;
wire v_631;
wire v_632;
wire v_633;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_640;
wire v_642;
wire v_643;
wire v_644;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire x_1;
assign v_1 = 1;
assign v_16 = 1;
assign v_21 = 1;
assign v_23 = 1;
assign v_30 = 1;
assign v_35 = 1;
assign v_54 = 1;
assign v_77 = 1;
assign v_81 = 1;
assign v_92 = 1;
assign v_97 = 1;
assign v_102 = 1;
assign v_113 = 1;
assign v_117 = 1;
assign v_126 = 1;
assign v_131 = 1;
assign v_135 = 1;
assign v_201 = 1;
assign v_204 = 1;
assign v_208 = 1;
assign v_329 = 1;
assign v_461 = 1;
assign v_466 = 1;
assign v_468 = 1;
assign v_475 = 1;
assign v_480 = 1;
assign v_499 = 1;
assign v_522 = 1;
assign v_526 = 1;
assign v_537 = 1;
assign v_542 = 1;
assign v_547 = 1;
assign v_558 = 1;
assign v_562 = 1;
assign v_571 = 1;
assign v_576 = 1;
assign v_580 = 1;
assign v_646 = 1;
assign v_648 = 1;
assign v_766 = 1;
assign v_12 = v_10 & v_11;
assign v_13 = v_10 & ~v_11;
assign v_17 = v_9 & v_14;
assign v_18 = ~v_9 & v_14;
assign v_27 = v_25 & ~v_26;
assign v_32 = v_31;
assign v_37 = ~v_36;
assign v_39 = v_36 & v_38;
assign v_42 = v_36 & ~v_38 & v_40 & v_41;
assign v_44 = v_36 & ~v_38 & v_40 & ~v_41 & ~v_43;
assign v_46 = v_36 & ~v_38 & ~v_40 & ~v_45;
assign v_48 = v_36 & ~v_38 & ~v_40 & v_45 & v_47;
assign v_50 = v_884 & v_885;
assign v_52 = v_886 & v_887;
assign v_56 = v_888 & v_889;
assign v_57 = v_890 & v_891;
assign v_60 = v_58 & v_59;
assign v_61 = v_58 & ~v_59;
assign v_63 = v_892 & v_893;
assign v_65 = ~v_31 & ~v_33 & v_64;
assign v_67 = ~v_31 & v_33 & ~v_66;
assign v_69 = ~v_31 & v_33 & v_66 & ~v_68;
assign v_70 = ~v_31 & v_33 & v_66 & v_68;
assign v_73 = v_71 & v_72;
assign v_74 = v_71 & ~v_72;
assign v_79 = v_24 & v_28 & v_75 & v_78;
assign v_82 = v_24 & v_28 & v_75 & ~v_78;
assign v_85 = v_83 & v_84;
assign v_86 = v_83 & ~v_84;
assign v_88 = v_8 & v_19 & v_87;
assign v_89 = ~v_8 & v_19;
assign v_93 = v_7 & v_90;
assign v_94 = ~v_7 & v_90;
assign v_98 = v_6 & v_95;
assign v_99 = ~v_6 & v_95;
assign v_103 = v_5 & v_100;
assign v_104 = ~v_5 & v_100;
assign v_106 = v_4 & v_105;
assign v_109 = v_108 & v_100;
assign v_110 = ~v_108 & v_100;
assign v_114 = v_107 & v_111;
assign v_118 = v_115 & v_111;
assign v_119 = ~v_115 & v_111;
assign v_121 = ~v_107 & v_120;
assign v_123 = ~v_4 & v_122;
assign v_127 = v_3 & v_124;
assign v_128 = ~v_3 & v_124;
assign v_132 = v_2 & v_129;
assign v_136 = v_133 & v_129;
assign v_137 = ~v_133 & v_129;
assign v_139 = ~v_2 & v_138;
assign v_143 = v_141 & v_142;
assign v_144 = v_141 & ~v_142;
assign v_147 = v_145 & v_146;
assign v_148 = v_145 & ~v_146;
assign v_152 = v_149 & ~v_150 & v_151;
assign v_153 = v_149 & ~v_150 & ~v_151;
assign v_155 = v_149 & v_150 & v_154;
assign v_156 = v_149 & v_150 & ~v_154;
assign v_159 = v_157 & v_158;
assign v_160 = v_157 & ~v_158;
assign v_163 = v_161 & v_162;
assign v_165 = v_161 & ~v_162 & v_164;
assign v_167 = v_161 & ~v_162 & ~v_164 & v_166;
assign v_169 = v_161 & ~v_162 & ~v_164 & ~v_166 & v_168;
assign v_172 = v_894 & v_895;
assign v_173 = v_896 & v_897;
assign v_176 = v_174 & v_175;
assign v_177 = v_174 & ~v_175;
assign v_180 = v_178 & v_179;
assign v_182 = v_898 & v_899;
assign v_183 = v_900 & v_901;
assign v_186 = v_184 & v_185;
assign v_187 = v_184 & ~v_185;
assign v_190 = v_188 & v_189;
assign v_191 = v_178 & ~v_179;
assign v_192 = v_188 & ~v_189;
assign v_195 = v_193 & ~v_194;
assign v_197 = v_193 & v_194 & v_196;
assign v_198 = v_193 & v_194 & ~v_196;
assign v_205 = v_202;
assign v_207 = v_140 & v_199 & v_206;
assign v_209 = v_9;
assign v_211 = v_210 & ~v_24;
assign v_212 = v_210 & v_31;
assign v_213 = v_210 & ~v_31 & v_33 & v_66 & ~v_68;
assign v_214 = v_210 & ~v_31 & v_33 & v_66 & v_68;
assign v_215 = v_210 & ~v_31 & v_33 & ~v_66;
assign v_216 = v_210 & v_34;
assign v_217 = v_210 & ~v_34;
assign v_220 = v_218 & v_219;
assign v_221 = v_902 & v_903;
assign v_223 = v_218 & v_222;
assign v_225 = v_224 & ~v_31 & ~v_33 & v_64;
assign v_227 = v_226 & v_71 & v_72;
assign v_228 = v_226 & v_71 & ~v_72;
assign v_230 = v_229 & v_24 & v_28 & v_75 & v_78;
assign v_231 = v_229 & v_24 & v_28 & v_75 & ~v_78;
assign v_234 = v_232 & v_233;
assign v_236 = v_8 & v_235;
assign v_237 = ~v_8 & v_210;
assign v_239 = v_238 & ~v_91;
assign v_240 = v_238 & v_91;
assign v_242 = v_7 & v_241;
assign v_243 = ~v_7 & v_238;
assign v_245 = v_244 & ~v_96;
assign v_246 = v_244 & v_96;
assign v_248 = v_6 & v_247;
assign v_249 = ~v_6 & v_244;
assign v_251 = v_250 & ~v_101;
assign v_252 = v_250 & v_101;
assign v_254 = v_5 & v_253;
assign v_255 = ~v_5 & v_250;
assign v_257 = v_4 & v_256;
assign v_258 = v_108 & v_253;
assign v_259 = ~v_108 & v_250;
assign v_261 = v_260 & ~v_112;
assign v_262 = v_260 & v_112;
assign v_264 = v_107 & v_263;
assign v_265 = v_260 & ~v_116;
assign v_266 = v_260 & v_116;
assign v_268 = v_115 & v_267;
assign v_269 = ~v_115 & v_260;
assign v_271 = ~v_107 & v_270;
assign v_273 = ~v_4 & v_272;
assign v_275 = v_274 & ~v_125;
assign v_276 = v_274 & v_125;
assign v_278 = v_3 & v_277;
assign v_279 = ~v_3 & v_274;
assign v_281 = v_280 & ~v_130;
assign v_282 = v_280 & v_130;
assign v_284 = v_2 & v_283;
assign v_285 = v_280 & ~v_134;
assign v_286 = v_280 & v_134;
assign v_288 = v_133 & v_287;
assign v_289 = ~v_133 & v_280;
assign v_291 = ~v_2 & v_290;
assign v_293 = v_292 & ~v_141;
assign v_294 = v_292 & v_141 & v_142;
assign v_295 = v_292 & v_141 & ~v_142;
assign v_297 = v_296 & v_145 & v_146;
assign v_298 = v_296 & v_145 & ~v_146;
assign v_300 = v_299 & v_157 & v_158;
assign v_301 = v_299 & v_157 & ~v_158;
assign v_304 = v_302 & v_303;
assign v_305 = v_904 & v_905;
assign v_306 = v_906 & v_907;
assign v_308 = v_307 & v_184 & v_185;
assign v_309 = v_307 & v_184 & ~v_185;
assign v_311 = v_310 & v_188 & v_189;
assign v_312 = v_310 & v_188 & ~v_189;
assign v_313 = v_908 & v_909;
assign v_314 = v_910 & v_911;
assign v_316 = v_315 & v_174 & v_175;
assign v_317 = v_315 & v_174 & ~v_175;
assign v_319 = v_318 & v_178 & v_179;
assign v_320 = v_318 & v_178 & ~v_179;
assign v_324 = v_321 & v_323;
assign v_326 = v_325 & v_202;
assign v_327 = v_325 & ~v_202;
assign v_330 = v_9;
assign v_332 = v_331 & ~v_24;
assign v_333 = v_331 & v_31;
assign v_334 = v_331 & ~v_31 & v_33 & v_66 & ~v_68;
assign v_335 = v_331 & ~v_31 & v_33 & v_66 & v_68;
assign v_336 = v_331 & ~v_31 & v_33 & ~v_66;
assign v_337 = v_331 & v_34;
assign v_338 = v_331 & ~v_34;
assign v_341 = v_339 & v_340;
assign v_342 = v_912 & v_913;
assign v_343 = v_339 & v_222;
assign v_345 = v_344 & ~v_31 & ~v_33 & v_64;
assign v_347 = v_346 & v_71 & v_72;
assign v_348 = v_346 & v_71 & ~v_72;
assign v_350 = v_349 & v_24 & v_28 & v_75 & v_78;
assign v_351 = v_349 & v_24 & v_28 & v_75 & ~v_78;
assign v_353 = v_352 & v_233;
assign v_355 = v_8 & v_354;
assign v_356 = ~v_8 & v_331;
assign v_358 = v_357 & ~v_91;
assign v_359 = v_357 & v_91;
assign v_361 = v_7 & v_360;
assign v_362 = ~v_7 & v_357;
assign v_364 = v_363 & ~v_96;
assign v_365 = v_363 & v_96;
assign v_367 = v_6 & v_366;
assign v_368 = ~v_6 & v_363;
assign v_370 = v_369 & ~v_101;
assign v_371 = v_369 & v_101;
assign v_373 = v_5 & v_372;
assign v_374 = ~v_5 & v_369;
assign v_376 = v_4 & v_375;
assign v_377 = v_108 & v_372;
assign v_378 = ~v_108 & v_369;
assign v_380 = v_379 & ~v_112;
assign v_381 = v_379 & v_112;
assign v_383 = v_107 & v_382;
assign v_384 = v_379 & ~v_116;
assign v_385 = v_379 & v_116;
assign v_387 = v_115 & v_386;
assign v_388 = ~v_115 & v_379;
assign v_390 = ~v_107 & v_389;
assign v_392 = ~v_4 & v_391;
assign v_394 = v_393 & ~v_125;
assign v_395 = v_393 & v_125;
assign v_397 = v_3 & v_396;
assign v_398 = ~v_3 & v_393;
assign v_400 = v_399 & ~v_130;
assign v_401 = v_399 & v_130;
assign v_403 = v_2 & v_402;
assign v_404 = v_399 & ~v_134;
assign v_405 = v_399 & v_134;
assign v_407 = v_133 & v_406;
assign v_408 = ~v_133 & v_399;
assign v_410 = ~v_2 & v_409;
assign v_412 = v_411 & ~v_141;
assign v_413 = v_411 & v_141 & v_142;
assign v_414 = v_411 & v_141 & ~v_142;
assign v_416 = v_415 & v_145 & v_146;
assign v_417 = v_415 & v_145 & ~v_146;
assign v_419 = v_418 & v_157 & v_158;
assign v_420 = v_418 & v_157 & ~v_158;
assign v_423 = v_421 & v_422;
assign v_424 = v_914 & v_915;
assign v_425 = v_916 & v_917;
assign v_427 = v_426 & v_184 & v_185;
assign v_428 = v_426 & v_184 & ~v_185;
assign v_430 = v_429 & v_188 & v_189;
assign v_431 = v_429 & v_188 & ~v_189;
assign v_432 = v_918 & v_919;
assign v_433 = v_920 & v_921;
assign v_435 = v_434 & v_174 & v_175;
assign v_436 = v_434 & v_174 & ~v_175;
assign v_438 = v_437 & v_178 & v_179;
assign v_439 = v_437 & v_178 & ~v_179;
assign v_442 = v_440 & v_441;
assign v_444 = v_443 & v_202;
assign v_445 = v_443 & ~v_202;
assign v_457 = v_455 & v_456;
assign v_458 = v_455 & ~v_456;
assign v_462 = v_454 & v_459;
assign v_463 = ~v_454 & v_459;
assign v_472 = v_470 & ~v_471;
assign v_477 = v_476;
assign v_482 = ~v_481;
assign v_484 = v_481 & v_483;
assign v_487 = v_481 & ~v_483 & v_485 & v_486;
assign v_489 = v_481 & ~v_483 & v_485 & ~v_486 & ~v_488;
assign v_491 = v_481 & ~v_483 & ~v_485 & ~v_490;
assign v_493 = v_481 & ~v_483 & ~v_485 & v_490 & v_492;
assign v_495 = v_922 & v_923;
assign v_497 = v_924 & v_925;
assign v_501 = v_926 & v_927;
assign v_502 = v_928 & v_929;
assign v_505 = v_503 & v_504;
assign v_506 = v_503 & ~v_504;
assign v_508 = v_930 & v_931;
assign v_510 = ~v_476 & ~v_478 & v_509;
assign v_512 = ~v_476 & v_478 & ~v_511;
assign v_514 = ~v_476 & v_478 & v_511 & ~v_513;
assign v_515 = ~v_476 & v_478 & v_511 & v_513;
assign v_518 = v_516 & v_517;
assign v_519 = v_516 & ~v_517;
assign v_524 = v_469 & v_473 & v_520 & v_523;
assign v_527 = v_469 & v_473 & v_520 & ~v_523;
assign v_530 = v_528 & v_529;
assign v_531 = v_528 & ~v_529;
assign v_533 = v_453 & v_464 & v_532;
assign v_534 = ~v_453 & v_464;
assign v_538 = v_452 & v_535;
assign v_539 = ~v_452 & v_535;
assign v_543 = v_451 & v_540;
assign v_544 = ~v_451 & v_540;
assign v_548 = v_450 & v_545;
assign v_549 = ~v_450 & v_545;
assign v_551 = v_449 & v_550;
assign v_554 = v_553 & v_545;
assign v_555 = ~v_553 & v_545;
assign v_559 = v_552 & v_556;
assign v_563 = v_560 & v_556;
assign v_564 = ~v_560 & v_556;
assign v_566 = ~v_552 & v_565;
assign v_568 = ~v_449 & v_567;
assign v_572 = v_448 & v_569;
assign v_573 = ~v_448 & v_569;
assign v_577 = v_447 & v_574;
assign v_581 = v_578 & v_574;
assign v_582 = ~v_578 & v_574;
assign v_584 = ~v_447 & v_583;
assign v_588 = v_586 & v_587;
assign v_589 = v_586 & ~v_587;
assign v_592 = v_590 & v_591;
assign v_593 = v_590 & ~v_591;
assign v_597 = v_594 & ~v_595 & v_596;
assign v_598 = v_594 & ~v_595 & ~v_596;
assign v_600 = v_594 & v_595 & v_599;
assign v_601 = v_594 & v_595 & ~v_599;
assign v_604 = v_602 & v_603;
assign v_605 = v_602 & ~v_603;
assign v_608 = v_606 & v_607;
assign v_610 = v_606 & ~v_607 & v_609;
assign v_612 = v_606 & ~v_607 & ~v_609 & v_611;
assign v_614 = v_606 & ~v_607 & ~v_609 & ~v_611 & v_613;
assign v_617 = v_932 & v_933;
assign v_618 = v_934 & v_935;
assign v_621 = v_619 & v_620;
assign v_622 = v_619 & ~v_620;
assign v_625 = v_623 & v_624;
assign v_627 = v_936 & v_937;
assign v_628 = v_938 & v_939;
assign v_631 = v_629 & v_630;
assign v_632 = v_629 & ~v_630;
assign v_635 = v_633 & v_634;
assign v_636 = v_623 & ~v_624;
assign v_637 = v_633 & ~v_634;
assign v_640 = v_638 & ~v_639;
assign v_642 = v_638 & v_639 & v_641;
assign v_643 = v_638 & v_639 & ~v_641;
assign v_647 = v_585 & v_644;
assign v_649 = v_454;
assign v_651 = v_650 & ~v_469;
assign v_652 = v_650 & v_476;
assign v_653 = v_650 & ~v_476 & v_478 & v_511 & ~v_513;
assign v_654 = v_650 & ~v_476 & v_478 & v_511 & v_513;
assign v_655 = v_650 & ~v_476 & v_478 & ~v_511;
assign v_656 = v_650 & v_479;
assign v_657 = v_650 & ~v_479;
assign v_660 = v_658 & v_659;
assign v_661 = v_940 & v_941;
assign v_663 = v_658 & v_662;
assign v_665 = v_664 & ~v_476 & ~v_478 & v_509;
assign v_667 = v_666 & v_516 & v_517;
assign v_668 = v_666 & v_516 & ~v_517;
assign v_670 = v_669 & v_469 & v_473 & v_520 & v_523;
assign v_671 = v_669 & v_469 & v_473 & v_520 & ~v_523;
assign v_674 = v_672 & v_673;
assign v_676 = v_453 & v_675;
assign v_677 = ~v_453 & v_650;
assign v_679 = v_678 & ~v_536;
assign v_680 = v_678 & v_536;
assign v_682 = v_452 & v_681;
assign v_683 = ~v_452 & v_678;
assign v_685 = v_684 & ~v_541;
assign v_686 = v_684 & v_541;
assign v_688 = v_451 & v_687;
assign v_689 = ~v_451 & v_684;
assign v_691 = v_690 & ~v_546;
assign v_692 = v_690 & v_546;
assign v_694 = v_450 & v_693;
assign v_695 = ~v_450 & v_690;
assign v_697 = v_449 & v_696;
assign v_698 = v_553 & v_693;
assign v_699 = ~v_553 & v_690;
assign v_701 = v_700 & ~v_557;
assign v_702 = v_700 & v_557;
assign v_704 = v_552 & v_703;
assign v_705 = v_700 & ~v_561;
assign v_706 = v_700 & v_561;
assign v_708 = v_560 & v_707;
assign v_709 = ~v_560 & v_700;
assign v_711 = ~v_552 & v_710;
assign v_713 = ~v_449 & v_712;
assign v_715 = v_714 & ~v_570;
assign v_716 = v_714 & v_570;
assign v_718 = v_448 & v_717;
assign v_719 = ~v_448 & v_714;
assign v_721 = v_720 & ~v_575;
assign v_722 = v_720 & v_575;
assign v_724 = v_447 & v_723;
assign v_725 = v_720 & ~v_579;
assign v_726 = v_720 & v_579;
assign v_728 = v_578 & v_727;
assign v_729 = ~v_578 & v_720;
assign v_731 = ~v_447 & v_730;
assign v_733 = v_732 & ~v_586;
assign v_734 = v_732 & v_586 & v_587;
assign v_735 = v_732 & v_586 & ~v_587;
assign v_737 = v_736 & v_590 & v_591;
assign v_738 = v_736 & v_590 & ~v_591;
assign v_740 = v_739 & v_602 & v_603;
assign v_741 = v_739 & v_602 & ~v_603;
assign v_744 = v_742 & v_743;
assign v_745 = v_942 & v_943;
assign v_746 = v_944 & v_945;
assign v_748 = v_747 & v_629 & v_630;
assign v_749 = v_747 & v_629 & ~v_630;
assign v_751 = v_750 & v_633 & v_634;
assign v_752 = v_750 & v_633 & ~v_634;
assign v_753 = v_946 & v_947;
assign v_754 = v_948 & v_949;
assign v_756 = v_755 & v_619 & v_620;
assign v_757 = v_755 & v_619 & ~v_620;
assign v_759 = v_758 & v_623 & v_624;
assign v_760 = v_758 & v_623 & ~v_624;
assign v_764 = v_761 & v_763;
assign v_767 = v_454;
assign v_769 = v_768 & ~v_469;
assign v_770 = v_768 & v_476;
assign v_771 = v_768 & ~v_476 & v_478 & v_511 & ~v_513;
assign v_772 = v_768 & ~v_476 & v_478 & v_511 & v_513;
assign v_773 = v_768 & ~v_476 & v_478 & ~v_511;
assign v_774 = v_768 & v_479;
assign v_775 = v_768 & ~v_479;
assign v_778 = v_776 & v_777;
assign v_779 = v_950 & v_951;
assign v_780 = v_776 & v_662;
assign v_782 = v_781 & ~v_476 & ~v_478 & v_509;
assign v_784 = v_783 & v_516 & v_517;
assign v_785 = v_783 & v_516 & ~v_517;
assign v_787 = v_786 & v_469 & v_473 & v_520 & v_523;
assign v_788 = v_786 & v_469 & v_473 & v_520 & ~v_523;
assign v_790 = v_789 & v_673;
assign v_792 = v_453 & v_791;
assign v_793 = ~v_453 & v_768;
assign v_795 = v_794 & ~v_536;
assign v_796 = v_794 & v_536;
assign v_798 = v_452 & v_797;
assign v_799 = ~v_452 & v_794;
assign v_801 = v_800 & ~v_541;
assign v_802 = v_800 & v_541;
assign v_804 = v_451 & v_803;
assign v_805 = ~v_451 & v_800;
assign v_807 = v_806 & ~v_546;
assign v_808 = v_806 & v_546;
assign v_810 = v_450 & v_809;
assign v_811 = ~v_450 & v_806;
assign v_813 = v_449 & v_812;
assign v_814 = v_553 & v_809;
assign v_815 = ~v_553 & v_806;
assign v_817 = v_816 & ~v_557;
assign v_818 = v_816 & v_557;
assign v_820 = v_552 & v_819;
assign v_821 = v_816 & ~v_561;
assign v_822 = v_816 & v_561;
assign v_824 = v_560 & v_823;
assign v_825 = ~v_560 & v_816;
assign v_827 = ~v_552 & v_826;
assign v_829 = ~v_449 & v_828;
assign v_831 = v_830 & ~v_570;
assign v_832 = v_830 & v_570;
assign v_834 = v_448 & v_833;
assign v_835 = ~v_448 & v_830;
assign v_837 = v_836 & ~v_575;
assign v_838 = v_836 & v_575;
assign v_840 = v_447 & v_839;
assign v_841 = v_836 & ~v_579;
assign v_842 = v_836 & v_579;
assign v_844 = v_578 & v_843;
assign v_845 = ~v_578 & v_836;
assign v_847 = ~v_447 & v_846;
assign v_849 = v_848 & ~v_586;
assign v_850 = v_848 & v_586 & v_587;
assign v_851 = v_848 & v_586 & ~v_587;
assign v_853 = v_852 & v_590 & v_591;
assign v_854 = v_852 & v_590 & ~v_591;
assign v_856 = v_855 & v_602 & v_603;
assign v_857 = v_855 & v_602 & ~v_603;
assign v_860 = v_858 & v_859;
assign v_861 = v_952 & v_953;
assign v_862 = v_954 & v_955;
assign v_864 = v_863 & v_629 & v_630;
assign v_865 = v_863 & v_629 & ~v_630;
assign v_867 = v_866 & v_633 & v_634;
assign v_868 = v_866 & v_633 & ~v_634;
assign v_869 = v_956 & v_957;
assign v_870 = v_958 & v_959;
assign v_872 = v_871 & v_619 & v_620;
assign v_873 = v_871 & v_619 & ~v_620;
assign v_875 = v_874 & v_623 & v_624;
assign v_876 = v_874 & v_623 & ~v_624;
assign v_879 = v_877 & v_878;
assign v_883 = ~v_881 & ~v_882 & v_647;
assign v_884 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_885 = v_49;
assign v_886 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_887 = ~v_49 & v_51;
assign v_888 = v_36 & ~v_38 & ~v_40 & v_45 & ~v_47;
assign v_889 = v_55;
assign v_890 = v_36 & ~v_38 & ~v_40 & v_45 & ~v_47;
assign v_891 = ~v_55;
assign v_892 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_893 = ~v_49 & ~v_51 & v_62;
assign v_894 = v_161 & ~v_162 & ~v_164 & ~v_166 & ~v_168;
assign v_895 = v_170 & v_171;
assign v_896 = v_161 & ~v_162 & ~v_164 & ~v_166 & ~v_168;
assign v_897 = v_170 & ~v_171;
assign v_898 = v_161 & ~v_162 & ~v_164 & ~v_166 & ~v_168;
assign v_899 = ~v_170 & v_181;
assign v_900 = v_161 & ~v_162 & ~v_164 & ~v_166 & ~v_168;
assign v_901 = ~v_170 & ~v_181;
assign v_902 = v_218 & v_36 & ~v_38 & v_40 & ~v_41;
assign v_903 = v_43 & ~v_49 & ~v_51 & v_62;
assign v_904 = v_302 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_905 = ~v_168 & ~v_170 & v_181;
assign v_906 = v_302 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_907 = ~v_168 & ~v_170 & ~v_181;
assign v_908 = v_302 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_909 = ~v_168 & v_170 & v_171;
assign v_910 = v_302 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_911 = ~v_168 & v_170 & ~v_171;
assign v_912 = v_339 & v_36 & ~v_38 & v_40 & ~v_41;
assign v_913 = v_43 & ~v_49 & ~v_51 & v_62;
assign v_914 = v_421 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_915 = ~v_168 & ~v_170 & v_181;
assign v_916 = v_421 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_917 = ~v_168 & ~v_170 & ~v_181;
assign v_918 = v_421 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_919 = ~v_168 & v_170 & v_171;
assign v_920 = v_421 & v_161 & ~v_162 & ~v_164 & ~v_166;
assign v_921 = ~v_168 & v_170 & ~v_171;
assign v_922 = v_481 & ~v_483 & v_485 & ~v_486 & v_488;
assign v_923 = v_494;
assign v_924 = v_481 & ~v_483 & v_485 & ~v_486 & v_488;
assign v_925 = ~v_494 & v_496;
assign v_926 = v_481 & ~v_483 & ~v_485 & v_490 & ~v_492;
assign v_927 = v_500;
assign v_928 = v_481 & ~v_483 & ~v_485 & v_490 & ~v_492;
assign v_929 = ~v_500;
assign v_930 = v_481 & ~v_483 & v_485 & ~v_486 & v_488;
assign v_931 = ~v_494 & ~v_496 & v_507;
assign v_932 = v_606 & ~v_607 & ~v_609 & ~v_611 & ~v_613;
assign v_933 = v_615 & v_616;
assign v_934 = v_606 & ~v_607 & ~v_609 & ~v_611 & ~v_613;
assign v_935 = v_615 & ~v_616;
assign v_936 = v_606 & ~v_607 & ~v_609 & ~v_611 & ~v_613;
assign v_937 = ~v_615 & v_626;
assign v_938 = v_606 & ~v_607 & ~v_609 & ~v_611 & ~v_613;
assign v_939 = ~v_615 & ~v_626;
assign v_940 = v_658 & v_481 & ~v_483 & v_485 & ~v_486;
assign v_941 = v_488 & ~v_494 & ~v_496 & v_507;
assign v_942 = v_742 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_943 = ~v_613 & ~v_615 & v_626;
assign v_944 = v_742 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_945 = ~v_613 & ~v_615 & ~v_626;
assign v_946 = v_742 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_947 = ~v_613 & v_615 & v_616;
assign v_948 = v_742 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_949 = ~v_613 & v_615 & ~v_616;
assign v_950 = v_776 & v_481 & ~v_483 & v_485 & ~v_486;
assign v_951 = v_488 & ~v_494 & ~v_496 & v_507;
assign v_952 = v_858 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_953 = ~v_613 & ~v_615 & v_626;
assign v_954 = v_858 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_955 = ~v_613 & ~v_615 & ~v_626;
assign v_956 = v_858 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_957 = ~v_613 & v_615 & v_616;
assign v_958 = v_858 & v_606 & ~v_607 & ~v_609 & ~v_611;
assign v_959 = ~v_613 & v_615 & ~v_616;
assign v_14 = ~v_10 | v_12 | v_13;
assign v_19 = v_17 | v_18;
assign v_28 = ~v_25 | v_27;
assign v_62 = ~v_58 | v_60 | v_61;
assign v_64 = v_960 | v_961 | v_962;
assign v_71 = v_65 | v_67 | v_69 | v_70;
assign v_75 = v_32 | v_73 | v_74;
assign v_83 = v_79 | v_82;
assign v_87 = ~v_24 | v_85 | v_86;
assign v_90 = v_88 | v_89;
assign v_95 = v_93 | v_94;
assign v_100 = v_98 | v_99;
assign v_105 = v_103 | v_104;
assign v_111 = v_109 | v_110;
assign v_120 = v_118 | v_119;
assign v_122 = v_114 | v_121;
assign v_124 = v_106 | v_123;
assign v_129 = v_127 | v_128;
assign v_138 = v_136 | v_137;
assign v_140 = v_132 | v_139;
assign v_145 = v_143 | v_144;
assign v_149 = v_147 | v_148;
assign v_157 = v_152 | v_153 | v_155 | v_156;
assign v_161 = v_159 | v_160;
assign v_174 = v_172 | v_173;
assign v_178 = v_176 | v_177;
assign v_184 = v_182 | v_183;
assign v_188 = v_186 | v_187;
assign v_193 = v_180 | v_190 | v_191 | v_192;
assign v_199 = v_963 | v_964;
assign v_206 = ~v_202 | v_205;
assign v_210 = v_209 | ~v_9;
assign v_218 = v_216 | v_217;
assign v_219 = v_965 | v_966;
assign v_222 = v_56 | v_57;
assign v_224 = v_220 | v_221 | v_223;
assign v_226 = v_213 | v_214 | v_215 | v_225;
assign v_229 = v_212 | v_227 | v_228;
assign v_232 = v_230 | v_231;
assign v_233 = v_85 | v_86;
assign v_235 = v_211 | v_234;
assign v_238 = v_236 | v_237;
assign v_241 = v_239 | v_240;
assign v_244 = v_242 | v_243;
assign v_247 = v_245 | v_246;
assign v_250 = v_248 | v_249;
assign v_253 = v_251 | v_252;
assign v_256 = v_254 | v_255;
assign v_260 = v_258 | v_259;
assign v_263 = v_261 | v_262;
assign v_267 = v_265 | v_266;
assign v_270 = v_268 | v_269;
assign v_272 = v_264 | v_271;
assign v_274 = v_257 | v_273;
assign v_277 = v_275 | v_276;
assign v_280 = v_278 | v_279;
assign v_283 = v_281 | v_282;
assign v_287 = v_285 | v_286;
assign v_290 = v_288 | v_289;
assign v_292 = v_284 | v_291;
assign v_296 = v_294 | v_295;
assign v_299 = v_297 | v_298;
assign v_302 = v_300 | v_301;
assign v_303 = v_163 | v_165 | v_167 | v_169;
assign v_307 = v_305 | v_306;
assign v_310 = v_308 | v_309;
assign v_315 = v_313 | v_314;
assign v_318 = v_316 | v_317;
assign v_321 = v_311 | v_312 | v_319 | v_320;
assign v_322 = v_197 | v_198;
assign v_323 = v_195 | v_322;
assign v_325 = v_293 | v_304 | v_324;
assign v_328 = v_326 | v_327;
assign v_331 = v_330 | ~v_9;
assign v_339 = v_337 | v_338;
assign v_340 = v_967 | v_968;
assign v_344 = v_341 | v_342 | v_343;
assign v_346 = v_334 | v_335 | v_336 | v_345;
assign v_349 = v_333 | v_347 | v_348;
assign v_352 = v_350 | v_351;
assign v_354 = v_332 | v_353;
assign v_357 = v_355 | v_356;
assign v_360 = v_358 | v_359;
assign v_363 = v_361 | v_362;
assign v_366 = v_364 | v_365;
assign v_369 = v_367 | v_368;
assign v_372 = v_370 | v_371;
assign v_375 = v_373 | v_374;
assign v_379 = v_377 | v_378;
assign v_382 = v_380 | v_381;
assign v_386 = v_384 | v_385;
assign v_389 = v_387 | v_388;
assign v_391 = v_383 | v_390;
assign v_393 = v_376 | v_392;
assign v_396 = v_394 | v_395;
assign v_399 = v_397 | v_398;
assign v_402 = v_400 | v_401;
assign v_406 = v_404 | v_405;
assign v_409 = v_407 | v_408;
assign v_411 = v_403 | v_410;
assign v_415 = v_413 | v_414;
assign v_418 = v_416 | v_417;
assign v_421 = v_419 | v_420;
assign v_422 = v_163 | v_165 | v_167 | v_169;
assign v_426 = v_424 | v_425;
assign v_429 = v_427 | v_428;
assign v_434 = v_432 | v_433;
assign v_437 = v_435 | v_436;
assign v_440 = v_430 | v_431 | v_438 | v_439;
assign v_441 = v_195 | v_322;
assign v_443 = v_412 | v_423 | v_442;
assign v_446 = v_444 | v_445;
assign v_459 = ~v_455 | v_457 | v_458;
assign v_464 = v_462 | v_463;
assign v_473 = ~v_470 | v_472;
assign v_507 = ~v_503 | v_505 | v_506;
assign v_509 = v_969 | v_970 | v_971;
assign v_516 = v_510 | v_512 | v_514 | v_515;
assign v_520 = v_477 | v_518 | v_519;
assign v_528 = v_524 | v_527;
assign v_532 = ~v_469 | v_530 | v_531;
assign v_535 = v_533 | v_534;
assign v_540 = v_538 | v_539;
assign v_545 = v_543 | v_544;
assign v_550 = v_548 | v_549;
assign v_556 = v_554 | v_555;
assign v_565 = v_563 | v_564;
assign v_567 = v_559 | v_566;
assign v_569 = v_551 | v_568;
assign v_574 = v_572 | v_573;
assign v_583 = v_581 | v_582;
assign v_585 = v_577 | v_584;
assign v_590 = v_588 | v_589;
assign v_594 = v_592 | v_593;
assign v_602 = v_597 | v_598 | v_600 | v_601;
assign v_606 = v_604 | v_605;
assign v_619 = v_617 | v_618;
assign v_623 = v_621 | v_622;
assign v_629 = v_627 | v_628;
assign v_633 = v_631 | v_632;
assign v_638 = v_625 | v_635 | v_636 | v_637;
assign v_644 = v_972 | v_973;
assign v_650 = v_649 | ~v_454;
assign v_658 = v_656 | v_657;
assign v_659 = v_974 | v_975;
assign v_662 = v_501 | v_502;
assign v_664 = v_660 | v_661 | v_663;
assign v_666 = v_653 | v_654 | v_655 | v_665;
assign v_669 = v_652 | v_667 | v_668;
assign v_672 = v_670 | v_671;
assign v_673 = v_530 | v_531;
assign v_675 = v_651 | v_674;
assign v_678 = v_676 | v_677;
assign v_681 = v_679 | v_680;
assign v_684 = v_682 | v_683;
assign v_687 = v_685 | v_686;
assign v_690 = v_688 | v_689;
assign v_693 = v_691 | v_692;
assign v_696 = v_694 | v_695;
assign v_700 = v_698 | v_699;
assign v_703 = v_701 | v_702;
assign v_707 = v_705 | v_706;
assign v_710 = v_708 | v_709;
assign v_712 = v_704 | v_711;
assign v_714 = v_697 | v_713;
assign v_717 = v_715 | v_716;
assign v_720 = v_718 | v_719;
assign v_723 = v_721 | v_722;
assign v_727 = v_725 | v_726;
assign v_730 = v_728 | v_729;
assign v_732 = v_724 | v_731;
assign v_736 = v_734 | v_735;
assign v_739 = v_737 | v_738;
assign v_742 = v_740 | v_741;
assign v_743 = v_608 | v_610 | v_612 | v_614;
assign v_747 = v_745 | v_746;
assign v_750 = v_748 | v_749;
assign v_755 = v_753 | v_754;
assign v_758 = v_756 | v_757;
assign v_761 = v_751 | v_752 | v_759 | v_760;
assign v_762 = v_642 | v_643;
assign v_763 = v_640 | v_762;
assign v_765 = v_733 | v_744 | v_764;
assign v_768 = v_767 | ~v_454;
assign v_776 = v_774 | v_775;
assign v_777 = v_976 | v_977;
assign v_781 = v_778 | v_779 | v_780;
assign v_783 = v_771 | v_772 | v_773 | v_782;
assign v_786 = v_770 | v_784 | v_785;
assign v_789 = v_787 | v_788;
assign v_791 = v_769 | v_790;
assign v_794 = v_792 | v_793;
assign v_797 = v_795 | v_796;
assign v_800 = v_798 | v_799;
assign v_803 = v_801 | v_802;
assign v_806 = v_804 | v_805;
assign v_809 = v_807 | v_808;
assign v_812 = v_810 | v_811;
assign v_816 = v_814 | v_815;
assign v_819 = v_817 | v_818;
assign v_823 = v_821 | v_822;
assign v_826 = v_824 | v_825;
assign v_828 = v_820 | v_827;
assign v_830 = v_813 | v_829;
assign v_833 = v_831 | v_832;
assign v_836 = v_834 | v_835;
assign v_839 = v_837 | v_838;
assign v_843 = v_841 | v_842;
assign v_846 = v_844 | v_845;
assign v_848 = v_840 | v_847;
assign v_852 = v_850 | v_851;
assign v_855 = v_853 | v_854;
assign v_858 = v_856 | v_857;
assign v_859 = v_608 | v_610 | v_612 | v_614;
assign v_863 = v_861 | v_862;
assign v_866 = v_864 | v_865;
assign v_871 = v_869 | v_870;
assign v_874 = v_872 | v_873;
assign v_877 = v_867 | v_868 | v_875 | v_876;
assign v_878 = v_640 | v_762;
assign v_880 = v_849 | v_860 | v_879;
assign v_960 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_961 = v_48 | v_50 | v_52 | v_56 | v_57;
assign v_962 = v_63;
assign v_963 = ~v_141 | v_163 | v_165 | v_167 | v_169;
assign v_964 = v_195 | v_197 | v_198;
assign v_965 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_966 = v_48 | v_50 | v_52;
assign v_967 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_968 = v_48 | v_50 | v_52;
assign v_969 = v_482 | v_484 | v_487 | v_489 | v_491;
assign v_970 = v_493 | v_495 | v_497 | v_501 | v_502;
assign v_971 = v_508;
assign v_972 = ~v_586 | v_608 | v_610 | v_612 | v_614;
assign v_973 = v_640 | v_642 | v_643;
assign v_974 = v_482 | v_484 | v_487 | v_489 | v_491;
assign v_975 = v_493 | v_495 | v_497;
assign v_976 = v_482 | v_484 | v_487 | v_489 | v_491;
assign v_977 = v_493 | v_495 | v_497;
assign v_881 = ~v_765 ^ ~v_328;
assign v_882 = ~v_880 ^ ~v_446;
assign x_1 = ~v_207 | v_883;
assign o_1 = x_1;
endmodule
