// Benchmark "genbuf15b4y_cert" written by ABC on Sun Jul 30 12:02:19 2017

module genbuf15b4y_cert ( 
    n87, reg_i_StoB_REQ4_out, reg_controllable_SLC1_out, sys_fair8done_out,
    reg_i_RtoB_ACK1_out, sys_fair14done_out, reg_i_StoB_REQ3_out,
    reg_controllable_SLC2_out, sys_fair7done_out, reg_i_StoB_REQ2_out,
    reg_controllable_SLC3_out, sys_fair9done_out,
    reg_controllable_BtoS_ACK10_out, env_fair1done_out,
    reg_i_StoB_REQ1_out, reg_controllable_BtoS_ACK11_out,
    sys_fair10done_out, reg_i_StoB_REQ0_out,
    reg_controllable_BtoS_ACK12_out, sys_fair6done_out, sys_fair11done_out,
    reg_controllable_BtoR_REQ0_out, reg_controllable_DEQ_out,
    reg_controllable_BtoS_ACK13_out, reg_controllable_BtoS_ACK14_out,
    sys_fair5done_out, reg_controllable_BtoR_REQ1_out,
    reg_controllable_ENQ_out, sys_fair12done_out, sys_fair4done_out,
    env_fair0done_out, reg_controllable_BtoS_ACK0_out, reg_nstateG7_1_out,
    reg_controllable_BtoS_ACK1_out, sys_fair13done_out,
    reg_controllable_BtoS_ACK2_out, sys_fair3done_out, reg_stateG7_0_out,
    reg_controllable_BtoS_ACK3_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , reg_controllable_BtoS_ACK4_out, sys_fair2done_out,
    reg_controllable_BtoS_ACK5_out, reg_controllable_BtoS_ACK6_out,
    sys_fair1done_out, reg_controllable_BtoS_ACK7_out, reg_i_nEMPTY_out,
    reg_controllable_BtoS_ACK8_out, reg_stateG12_out, sys_fair0done_out,
    reg_controllable_BtoS_ACK9_out, reg_i_StoB_REQ14_out, reg_i_FULL_out,
    reg_i_StoB_REQ13_out, reg_i_StoB_REQ9_out, env_safe_err_happened_out,
    reg_i_StoB_REQ8_out, reg_i_StoB_REQ12_out, reg_i_StoB_REQ7_out,
    reg_i_StoB_REQ11_out, reg_i_StoB_REQ6_out, reg_i_StoB_REQ10_out,
    sys_fair15done_out, reg_i_RtoB_ACK0_out, reg_i_StoB_REQ5_out,
    reg_controllable_SLC0_out, i_StoB_REQ0, i_StoB_REQ1, i_FULL,
    i_StoB_REQ2, i_StoB_REQ3, i_StoB_REQ4, i_StoB_REQ5, i_StoB_REQ6,
    i_StoB_REQ7, i_StoB_REQ8, i_StoB_REQ9, i_StoB_REQ10, i_StoB_REQ11,
    i_StoB_REQ12, i_StoB_REQ13, i_StoB_REQ14, i_nEMPTY, i_RtoB_ACK1,
    i_RtoB_ACK0, controllable_SLC2, controllable_SLC3, controllable_DEQ,
    controllable_BtoR_REQ0, controllable_BtoR_REQ1, controllable_BtoS_ACK0,
    controllable_BtoS_ACK1, controllable_BtoS_ACK2, controllable_BtoS_ACK3,
    controllable_BtoS_ACK4, controllable_BtoS_ACK5, controllable_BtoS_ACK6,
    controllable_BtoS_ACK7, controllable_BtoS_ACK8, controllable_BtoS_ACK9,
    controllable_BtoS_ACK10, controllable_ENQ, controllable_BtoS_ACK11,
    controllable_BtoS_ACK12, controllable_BtoS_ACK13,
    controllable_BtoS_ACK14, controllable_SLC0, controllable_SLC1,
    inductivity_check   );
  input  n87, reg_i_StoB_REQ4_out, reg_controllable_SLC1_out,
    sys_fair8done_out, reg_i_RtoB_ACK1_out, sys_fair14done_out,
    reg_i_StoB_REQ3_out, reg_controllable_SLC2_out, sys_fair7done_out,
    reg_i_StoB_REQ2_out, reg_controllable_SLC3_out, sys_fair9done_out,
    reg_controllable_BtoS_ACK10_out, env_fair1done_out,
    reg_i_StoB_REQ1_out, reg_controllable_BtoS_ACK11_out,
    sys_fair10done_out, reg_i_StoB_REQ0_out,
    reg_controllable_BtoS_ACK12_out, sys_fair6done_out, sys_fair11done_out,
    reg_controllable_BtoR_REQ0_out, reg_controllable_DEQ_out,
    reg_controllable_BtoS_ACK13_out, reg_controllable_BtoS_ACK14_out,
    sys_fair5done_out, reg_controllable_BtoR_REQ1_out,
    reg_controllable_ENQ_out, sys_fair12done_out, sys_fair4done_out,
    env_fair0done_out, reg_controllable_BtoS_ACK0_out, reg_nstateG7_1_out,
    reg_controllable_BtoS_ACK1_out, sys_fair13done_out,
    reg_controllable_BtoS_ACK2_out, sys_fair3done_out, reg_stateG7_0_out,
    reg_controllable_BtoS_ACK3_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , reg_controllable_BtoS_ACK4_out, sys_fair2done_out,
    reg_controllable_BtoS_ACK5_out, reg_controllable_BtoS_ACK6_out,
    sys_fair1done_out, reg_controllable_BtoS_ACK7_out, reg_i_nEMPTY_out,
    reg_controllable_BtoS_ACK8_out, reg_stateG12_out, sys_fair0done_out,
    reg_controllable_BtoS_ACK9_out, reg_i_StoB_REQ14_out, reg_i_FULL_out,
    reg_i_StoB_REQ13_out, reg_i_StoB_REQ9_out, env_safe_err_happened_out,
    reg_i_StoB_REQ8_out, reg_i_StoB_REQ12_out, reg_i_StoB_REQ7_out,
    reg_i_StoB_REQ11_out, reg_i_StoB_REQ6_out, reg_i_StoB_REQ10_out,
    sys_fair15done_out, reg_i_RtoB_ACK0_out, reg_i_StoB_REQ5_out,
    reg_controllable_SLC0_out, i_StoB_REQ0, i_StoB_REQ1, i_FULL,
    i_StoB_REQ2, i_StoB_REQ3, i_StoB_REQ4, i_StoB_REQ5, i_StoB_REQ6,
    i_StoB_REQ7, i_StoB_REQ8, i_StoB_REQ9, i_StoB_REQ10, i_StoB_REQ11,
    i_StoB_REQ12, i_StoB_REQ13, i_StoB_REQ14, i_nEMPTY, i_RtoB_ACK1,
    i_RtoB_ACK0, controllable_SLC2, controllable_SLC3, controllable_DEQ,
    controllable_BtoR_REQ0, controllable_BtoR_REQ1, controllable_BtoS_ACK0,
    controllable_BtoS_ACK1, controllable_BtoS_ACK2, controllable_BtoS_ACK3,
    controllable_BtoS_ACK4, controllable_BtoS_ACK5, controllable_BtoS_ACK6,
    controllable_BtoS_ACK7, controllable_BtoS_ACK8, controllable_BtoS_ACK9,
    controllable_BtoS_ACK10, controllable_ENQ, controllable_BtoS_ACK11,
    controllable_BtoS_ACK12, controllable_BtoS_ACK13,
    controllable_BtoS_ACK14, controllable_SLC0, controllable_SLC1;
  output inductivity_check ;
  wire n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
    n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
    n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
    n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
    n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
    n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
    n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
    n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
    n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
    n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
    n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
    n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
    n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
    n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
    n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
    n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
    n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
    n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
    n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
    n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
    n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
    n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
    n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
    n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
    n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
    n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
    n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
    n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
    n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
    n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
    n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
    n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
    n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
    n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
    n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
    n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
    n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
    n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
    n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
    n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
    n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
    n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
    n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
    n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
    n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
    n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
    n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
    n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
    n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
    n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
    n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
    n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
    n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
    n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
    n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
    n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
    n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
    n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
    n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
    n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
    n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
    n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
    n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
    n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
    n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
    n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
    n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
    n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
    n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
    n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
    n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
    n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
    n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
    n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
    n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
    n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
    n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
    n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
    n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
    n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
    n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
    n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
    n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
    n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
    n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
    n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
    n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
    n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
    n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
    n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
    n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
    n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
    n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
    n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
    n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
    n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
    n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
    n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
    n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
    n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
    n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
    n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
    n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
    n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
    n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
    n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
    n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
    n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
    n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
    n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
    n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
    n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
    n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
    n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
    n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
    n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
    n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
    n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
    n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
    n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
    n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
    n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
    n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
    n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
    n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
    n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
    n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
    n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
    n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
    n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
    n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
    n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
    n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
    n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
    n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
    n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
    n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
    n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
    n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
    n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
    n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
    n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
    n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
    n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
    n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
    n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
    n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
    n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
    n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
    n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
    n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
    n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
    n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
    n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
    n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
    n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
    n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
    n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
    n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
    n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
    n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
    n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
    n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
    n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
    n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
    n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
    n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
    n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
    n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
    n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
    n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
    n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
    n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
    n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
    n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
    n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
    n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
    n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
    n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
    n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
    n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
    n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
    n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
    n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
    n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
    n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
    n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
    n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
    n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
    n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
    n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
    n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
    n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
    n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
    n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
    n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
    n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
    n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
    n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
    n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
    n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
    n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
    n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
    n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
    n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
    n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
    n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
    n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
    n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
    n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
    n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
    n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
    n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
    n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
    n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
    n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
    n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
    n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
    n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
    n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
    n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
    n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
    n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
    n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
    n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
    n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
    n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
    n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
    n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
    n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
    n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
    n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
    n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
    n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
    n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
    n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
    n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
    n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
    n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
    n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
    n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
    n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
    n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
    n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
    n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
    n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
    n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
    n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
    n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
    n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
    n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
    n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
    n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
    n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
    n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
    n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
    n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
    n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
    n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
    n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
    n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
    n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
    n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
    n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
    n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
    n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
    n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
    n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
    n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
    n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
    n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
    n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
    n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
    n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
    n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
    n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
    n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
    n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
    n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
    n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
    n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
    n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
    n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
    n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
    n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
    n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
    n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
    n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
    n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
    n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
    n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
    n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
    n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
    n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
    n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
    n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
    n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
    n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
    n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
    n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
    n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
    n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
    n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
    n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
    n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
    n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
    n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
    n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
    n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
    n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
    n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
    n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
    n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
    n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
    n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
    n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
    n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
    n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
    n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
    n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
    n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
    n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
    n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
    n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
    n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
    n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
    n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
    n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
    n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
    n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
    n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
    n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
    n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
    n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
    n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
    n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
    n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
    n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
    n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
    n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
    n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
    n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
    n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
    n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
    n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
    n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
    n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
    n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
    n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
    n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
    n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
    n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
    n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
    n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
    n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
    n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
    n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
    n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
    n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
    n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
    n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
    n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
    n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
    n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
    n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
    n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
    n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
    n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
    n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
    n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
    n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
    n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
    n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
    n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
    n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
    n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
    n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
    n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
    n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
    n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
    n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
    n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
    n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
    n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
    n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
    n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
    n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
    n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
    n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
    n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
    n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
    n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
    n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
    n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
    n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
    n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
    n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
    n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
    n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
    n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
    n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
    n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
    n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
    n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
    n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
    n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
    n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
    n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
    n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
    n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
    n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
    n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
    n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
    n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
    n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
    n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
    n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
    n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
    n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758,
    n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
    n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
    n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
    n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
    n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
    n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
    n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
    n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
    n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
    n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
    n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
    n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
    n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
    n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
    n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
    n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
    n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
    n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
    n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
    n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
    n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
    n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
    n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
    n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046,
    n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
    n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
    n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
    n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
    n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
    n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
    n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
    n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
    n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
    n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
    n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
    n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
    n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
    n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
    n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
    n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
    n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
    n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
    n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
    n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
    n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
    n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
    n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
    n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
    n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
    n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
    n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
    n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
    n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
    n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
    n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
    n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
    n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
    n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
    n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
    n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
    n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
    n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
    n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
    n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
    n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
    n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
    n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
    n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
    n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
    n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
    n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
    n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
    n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
    n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
    n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
    n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
    n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
    n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
    n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
    n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
    n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
    n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
    n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
    n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
    n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
    n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
    n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
    n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
    n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
    n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
    n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
    n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
    n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
    n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
    n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
    n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
    n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
    n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
    n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
    n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
    n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
    n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
    n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
    n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
    n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
    n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
    n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
    n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
    n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
    n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
    n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
    n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
    n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
    n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
    n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
    n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
    n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
    n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
    n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
    n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
    n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
    n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
    n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
    n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
    n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
    n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
    n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
    n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
    n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
    n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
    n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
    n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
    n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
    n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
    n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
    n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
    n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
    n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
    n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
    n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
    n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
    n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
    n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
    n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
    n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
    n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
    n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
    n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
    n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
    n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
    n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
    n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
    n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
    n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422,
    n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
    n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
    n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
    n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
    n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485,
    n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494,
    n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
    n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
    n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
    n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
    n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
    n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
    n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566,
    n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
    n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
    n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
    n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
    n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
    n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
    n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
    n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638,
    n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
    n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
    n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
    n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
    n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
    n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
    n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
    n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710,
    n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
    n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
    n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
    n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
    n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
    n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
    n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
    n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
    n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
    n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
    n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
    n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
    n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
    n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
    n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
    n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
    n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
    n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
    n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
    n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
    n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
    n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
    n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
    n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998,
    n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
    n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016,
    n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
    n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
    n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
    n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
    n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
    n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
    n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
    n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088,
    n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
    n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
    n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
    n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
    n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133,
    n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142,
    n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
    n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160,
    n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
    n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
    n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
    n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
    n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
    n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
    n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
    n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
    n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
    n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
    n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
    n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
    n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
    n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
    n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
    n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
    n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
    n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
    n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
    n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
    n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
    n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
    n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
    n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
    n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
    n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
    n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
    n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
    n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
    n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
    n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
    n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
    n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
    n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
    n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
    n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
    n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
    n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
    n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
    n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
    n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
    n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
    n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
    n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
    n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
    n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
    n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925,
    n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
    n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
    n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
    n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
    n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997,
    n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006,
    n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
    n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
    n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
    n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
    n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
    n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
    n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069,
    n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
    n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
    n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
    n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
    n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
    n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
    n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
    n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
    n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
    n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
    n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
    n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
    n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204,
    n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213,
    n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
    n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
    n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
    n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
    n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
    n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
    n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
    n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
    n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357,
    n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
    n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
    n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
    n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
    n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
    n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
    n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
    n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501,
    n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
    n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
    n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
    n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573,
    n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
    n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
    n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
    n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645,
    n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
    n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
    n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
    n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
    n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
    n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708,
    n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
    n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
    n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
    n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
    n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
    n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
    n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
    n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
    n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
    n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
    n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852,
    n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861,
    n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
    n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
    n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
    n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
    n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
    n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
    n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924,
    n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933,
    n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
    n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
    n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
    n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996,
    n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005,
    n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
    n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
    n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
    n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
    n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
    n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
    n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068,
    n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077,
    n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
    n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
    n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
    n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
    n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
    n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
    n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
    n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
    n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
    n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
    n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
    n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212,
    n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221,
    n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
    n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
    n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
    n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
    n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
    n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
    n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284,
    n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
    n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
    n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
    n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
    n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
    n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
    n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
    n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356,
    n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365,
    n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
    n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
    n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
    n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428,
    n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
    n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
    n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
    n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
    n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
    n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
    n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500,
    n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509,
    n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
    n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
    n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
    n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
    n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572,
    n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581,
    n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
    n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
    n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
    n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
    n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
    n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
    n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644,
    n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653,
    n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662,
    n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
    n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
    n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
    n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
    n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
    n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716,
    n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734,
    n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
    n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
    n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
    n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
    n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
    n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
    n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860,
    n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869,
    n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878,
    n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
    n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
    n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
    n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
    n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
    n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950,
    n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
    n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
    n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
    n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
    n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
    n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013,
    n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022,
    n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
    n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
    n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
    n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
    n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
    n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
    n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085,
    n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
    n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
    n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
    n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
    n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
    n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
    n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
    n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157,
    n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166,
    n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
    n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
    n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
    n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
    n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
    n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
    n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229,
    n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
    n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
    n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
    n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
    n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
    n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
    n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301,
    n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
    n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
    n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
    n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
    n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
    n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
    n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
    n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373,
    n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
    n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
    n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
    n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
    n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
    n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
    n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445,
    n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454,
    n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
    n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
    n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
    n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517,
    n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
    n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
    n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
    n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
    n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589,
    n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
    n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
    n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
    n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661,
    n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670,
    n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
    n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
    n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
    n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
    n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
    n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733,
    n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
    n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
    n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
    n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
    n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805,
    n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814,
    n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
    n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
    n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
    n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
    n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
    n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
    n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877,
    n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886,
    n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
    n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
    n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
    n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
    n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
    n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949,
    n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958,
    n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
    n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
    n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
    n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
    n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
    n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
    n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021,
    n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
    n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039,
    n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
    n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
    n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
    n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
    n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
    n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
    n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
    n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
    n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
    n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
    n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
    n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165,
    n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
    n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
    n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
    n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237,
    n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
    n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264,
    n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
    n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
    n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
    n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
    n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309,
    n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318,
    n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
    n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336,
    n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
    n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
    n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
    n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
    n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381,
    n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
    n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
    n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
    n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453,
    n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471,
    n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
    n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
    n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
    n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
    n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
    n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525,
    n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534,
    n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
    n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
    n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
    n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
    n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
    n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
    n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597,
    n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606,
    n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615,
    n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
    n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
    n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
    n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
    n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
    n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669,
    n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
    n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
    n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
    n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
    n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
    n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
    n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
    n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
    n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
    n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
    n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
    n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
    n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
    n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813,
    n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
    n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
    n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
    n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
    n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
    n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
    n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885,
    n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
    n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
    n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
    n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
    n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
    n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
    n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957,
    n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
    n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
    n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
    n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
    n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
    n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
    n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
    n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029,
    n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
    n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
    n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
    n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
    n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
    n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
    n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101,
    n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
    n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
    n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
    n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
    n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
    n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
    n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173,
    n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
    n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
    n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
    n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245,
    n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
    n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263,
    n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
    n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
    n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
    n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
    n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
    n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317,
    n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
    n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
    n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
    n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
    n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
    n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
    n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
    n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389,
    n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
    n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407,
    n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
    n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
    n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
    n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
    n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
    n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
    n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
    n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
    n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
    n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
    n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
    n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
    n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
    n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
    n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
    n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
    n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
    n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
    n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
    n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
    n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605,
    n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
    n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623,
    n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
    n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
    n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
    n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
    n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
    n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677,
    n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
    n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695,
    n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
    n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
    n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
    n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
    n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
    n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749,
    n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
    n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767,
    n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
    n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
    n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
    n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
    n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
    n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821,
    n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
    n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839,
    n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
    n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
    n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
    n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
    n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
    n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893,
    n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
    n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
    n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
    n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
    n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965,
    n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
    n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
    n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
    n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
    n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037,
    n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
    n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
    n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
    n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
    n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
    n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
    n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109,
    n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
    n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
    n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
    n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
    n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
    n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
    n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
    n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181,
    n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
    n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
    n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
    n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
    n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
    n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
    n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
    n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253,
    n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
    n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
    n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
    n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
    n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
    n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
    n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
    n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325,
    n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
    n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
    n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
    n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
    n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
    n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
    n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
    n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397,
    n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
    n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
    n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
    n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
    n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
    n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
    n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
    n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469,
    n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
    n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
    n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
    n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
    n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
    n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
    n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
    n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541,
    n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
    n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
    n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
    n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
    n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
    n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
    n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
    n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613,
    n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
    n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
    n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
    n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
    n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
    n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
    n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685,
    n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
    n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
    n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
    n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
    n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
    n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
    n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757,
    n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
    n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
    n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
    n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
    n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
    n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
    n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
    n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829,
    n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
    n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
    n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856,
    n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
    n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
    n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
    n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892,
    n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901,
    n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
    n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
    n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928,
    n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
    n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
    n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
    n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964,
    n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973,
    n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
    n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
    n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000,
    n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
    n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
    n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
    n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036,
    n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045,
    n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
    n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
    n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
    n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
    n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
    n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
    n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
    n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117,
    n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
    n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
    n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
    n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
    n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
    n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
    n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180,
    n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189,
    n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
    n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
    n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
    n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
    n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
    n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
    n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
    n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261,
    n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
    n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
    n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
    n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
    n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
    n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324,
    n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
    n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
    n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
    n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
    n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
    n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
    n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
    n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405,
    n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
    n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
    n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
    n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
    n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
    n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
    n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468,
    n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477,
    n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
    n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
    n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
    n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
    n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
    n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
    n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
    n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549,
    n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
    n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
    n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
    n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
    n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
    n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
    n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621,
    n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
    n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
    n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
    n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
    n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
    n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693,
    n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
    n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
    n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720,
    n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
    n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
    n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
    n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756,
    n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765,
    n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
    n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
    n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
    n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
    n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837,
    n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
    n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
    n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
    n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900,
    n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909,
    n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
    n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
    n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
    n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
    n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
    n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
    n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972,
    n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981,
    n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
    n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
    n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008,
    n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
    n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
    n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
    n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044,
    n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053,
    n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
    n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080,
    n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
    n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
    n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
    n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116,
    n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125,
    n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143,
    n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
    n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
    n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
    n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188,
    n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197,
    n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
    n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
    n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
    n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260,
    n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269,
    n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
    n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296,
    n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
    n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
    n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
    n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332,
    n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341,
    n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
    n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359,
    n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368,
    n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
    n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
    n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
    n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404,
    n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413,
    n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
    n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431,
    n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
    n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
    n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
    n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
    n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476,
    n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485,
    n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
    n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
    n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512,
    n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
    n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
    n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
    n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548,
    n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557,
    n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
    n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
    n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584,
    n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
    n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
    n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629,
    n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
    n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
    n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
    n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
    n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692,
    n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701,
    n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
    n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719,
    n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728,
    n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
    n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
    n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
    n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764,
    n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773,
    n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
    n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791,
    n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800,
    n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
    n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
    n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
    n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836,
    n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845,
    n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
    n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863,
    n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
    n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
    n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
    n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
    n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908,
    n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917,
    n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
    n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935,
    n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
    n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980,
    n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989,
    n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
    n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007,
    n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
    n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
    n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
    n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
    n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052,
    n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061,
    n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
    n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079,
    n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
    n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
    n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
    n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133,
    n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151,
    n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
    n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
    n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196,
    n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205,
    n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
    n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223,
    n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
    n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
    n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
    n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
    n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268,
    n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277,
    n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
    n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
    n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
    n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
    n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
    n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
    n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340,
    n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349,
    n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
    n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367,
    n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
    n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
    n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
    n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
    n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412,
    n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421,
    n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
    n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439,
    n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
    n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
    n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
    n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
    n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484,
    n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493,
    n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
    n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511,
    n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
    n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
    n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
    n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556,
    n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565,
    n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
    n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583,
    n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
    n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
    n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
    n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
    n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628,
    n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637,
    n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
    n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
    n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
    n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
    n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
    n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
    n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709,
    n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
    n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
    n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
    n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
    n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
    n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
    n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772,
    n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781,
    n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
    n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799,
    n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
    n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
    n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
    n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
    n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844,
    n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853,
    n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
    n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871,
    n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
    n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
    n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
    n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
    n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916,
    n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925,
    n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
    n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
    n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
    n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
    n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
    n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
    n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997,
    n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
    n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
    n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
    n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
    n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
    n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
    n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
    n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
    n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
    n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
    n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
    n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
    n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
    n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
    n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204,
    n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
    n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
    n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276,
    n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285,
    n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
    n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
    n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
    n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
    n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348,
    n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
    n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
    n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
    n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420,
    n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
    n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
    n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
    n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483,
    n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492,
    n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501,
    n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
    n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519,
    n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
    n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
    n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
    n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
    n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564,
    n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573,
    n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
    n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591,
    n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
    n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
    n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
    n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
    n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636,
    n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645,
    n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
    n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663,
    n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
    n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
    n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
    n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699,
    n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708,
    n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717,
    n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
    n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735,
    n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
    n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
    n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
    n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771,
    n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780,
    n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789,
    n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
    n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
    n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
    n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
    n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
    n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
    n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852,
    n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861,
    n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
    n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879,
    n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
    n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
    n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
    n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
    n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924,
    n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933,
    n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
    n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951,
    n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
    n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
    n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
    n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
    n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996,
    n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005,
    n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
    n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
    n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
    n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
    n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
    n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
    n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068,
    n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077,
    n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
    n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
    n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
    n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
    n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
    n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
    n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140,
    n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149,
    n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
    n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167,
    n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
    n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
    n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
    n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
    n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212,
    n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221,
    n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
    n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239,
    n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
    n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
    n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
    n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
    n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284,
    n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293,
    n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
    n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
    n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
    n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
    n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
    n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
    n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356,
    n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365,
    n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
    n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383,
    n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
    n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
    n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
    n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
    n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428,
    n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437,
    n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
    n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
    n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
    n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
    n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
    n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
    n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500,
    n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509,
    n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
    n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527,
    n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
    n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
    n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
    n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
    n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572,
    n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581,
    n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
    n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
    n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
    n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
    n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
    n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
    n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644,
    n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653,
    n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
    n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671,
    n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
    n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
    n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
    n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
    n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
    n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725,
    n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
    n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743,
    n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
    n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
    n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
    n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788,
    n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797,
    n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
    n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815,
    n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
    n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
    n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
    n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
    n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860,
    n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869,
    n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
    n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887,
    n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
    n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
    n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
    n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
    n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932,
    n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941,
    n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
    n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
    n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
    n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
    n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
    n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
    n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004,
    n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013,
    n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
    n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
    n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
    n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
    n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
    n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
    n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085,
    n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
    n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
    n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
    n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
    n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
    n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148,
    n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157,
    n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
    n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
    n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
    n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
    n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
    n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
    n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220,
    n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229,
    n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
    n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
    n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
    n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
    n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
    n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
    n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301,
    n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
    n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
    n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
    n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
    n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373,
    n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
    n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
    n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
    n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
    n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
    n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445,
    n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
    n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
    n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
    n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
    n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
    n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508,
    n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517,
    n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
    n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
    n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
    n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
    n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
    n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
    n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580,
    n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589,
    n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
    n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607,
    n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
    n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
    n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
    n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652,
    n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661,
    n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
    n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679,
    n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
    n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
    n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
    n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
    n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
    n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733,
    n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
    n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751,
    n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
    n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
    n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
    n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
    n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796,
    n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805,
    n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
    n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823,
    n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
    n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
    n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
    n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
    n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868,
    n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877,
    n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
    n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895,
    n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
    n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
    n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949,
    n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
    n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967,
    n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
    n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
    n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
    n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
    n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021,
    n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
    n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
    n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
    n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
    n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
    n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
    n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093,
    n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102,
    n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
    n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
    n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
    n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
    n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
    n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156,
    n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165,
    n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174,
    n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183,
    n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
    n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
    n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
    n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
    n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228,
    n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237,
    n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246,
    n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255,
    n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
    n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
    n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
    n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
    n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300,
    n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309,
    n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318,
    n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327,
    n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
    n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
    n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
    n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
    n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
    n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381,
    n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390,
    n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
    n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
    n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
    n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
    n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
    n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444,
    n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453,
    n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462,
    n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
    n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
    n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
    n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
    n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525,
    n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
    n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
    n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
    n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
    n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
    n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588,
    n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597,
    n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606,
    n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615,
    n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
    n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
    n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
    n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
    n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660,
    n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669,
    n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
    n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687,
    n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
    n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
    n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
    n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
    n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732,
    n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741,
    n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
    n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759,
    n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
    n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
    n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
    n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
    n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804,
    n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813,
    n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
    n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831,
    n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
    n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
    n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
    n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
    n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876,
    n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885,
    n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903,
    n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
    n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
    n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
    n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
    n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948,
    n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957,
    n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
    n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975,
    n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
    n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
    n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
    n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
    n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020,
    n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029,
    n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047,
    n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
    n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
    n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
    n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
    n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092,
    n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101,
    n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
    n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119,
    n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
    n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
    n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
    n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173,
    n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
    n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191,
    n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
    n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
    n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
    n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
    n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
    n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245,
    n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
    n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263,
    n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
    n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
    n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
    n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
    n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
    n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317,
    n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
    n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335,
    n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
    n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
    n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
    n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
    n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380,
    n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389,
    n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
    n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407,
    n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
    n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
    n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
    n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
    n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452,
    n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461,
    n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
    n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479,
    n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488,
    n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
    n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
    n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
    n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524,
    n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533,
    n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
    n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551,
    n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560,
    n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
    n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
    n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596,
    n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605,
    n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623,
    n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
    n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
    n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
    n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668,
    n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677,
    n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
    n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695,
    n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704,
    n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
    n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
    n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
    n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740,
    n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749,
    n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
    n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767,
    n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
    n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
    n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
    n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
    n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812,
    n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821,
    n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
    n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839,
    n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848,
    n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
    n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
    n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
    n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884,
    n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893,
    n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
    n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911,
    n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920,
    n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
    n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
    n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
    n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956,
    n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965,
    n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
    n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983,
    n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992,
    n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
    n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
    n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
    n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028,
    n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037,
    n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
    n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055,
    n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
    n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
    n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
    n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
    n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100,
    n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109,
    n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
    n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127,
    n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
    n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
    n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
    n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
    n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172,
    n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181,
    n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
    n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199,
    n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
    n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
    n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
    n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
    n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244,
    n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253,
    n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
    n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271,
    n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
    n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
    n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
    n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
    n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316,
    n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325,
    n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
    n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343,
    n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
    n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
    n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397,
    n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415,
    n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
    n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
    n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469,
    n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487,
    n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
    n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
    n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541,
    n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
    n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559,
    n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568,
    n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
    n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
    n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
    n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604,
    n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613,
    n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
    n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631,
    n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640,
    n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
    n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
    n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
    n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676,
    n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685,
    n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
    n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703,
    n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712,
    n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
    n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
    n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
    n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748,
    n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757,
    n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
    n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775,
    n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
    n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
    n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
    n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
    n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820,
    n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829,
    n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847,
    n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856,
    n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
    n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
    n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
    n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892,
    n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901,
    n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
    n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919,
    n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928,
    n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
    n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
    n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
    n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964,
    n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973,
    n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
    n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991,
    n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000,
    n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
    n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
    n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
    n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036,
    n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045,
    n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
    n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063,
    n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072,
    n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
    n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
    n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
    n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108,
    n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117,
    n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
    n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135,
    n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144,
    n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
    n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
    n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
    n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180,
    n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189,
    n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
    n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207,
    n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216,
    n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
    n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
    n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
    n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252,
    n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261,
    n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
    n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279,
    n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288,
    n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
    n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
    n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
    n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324,
    n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333,
    n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
    n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351,
    n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
    n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
    n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
    n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
    n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396,
    n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405,
    n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
    n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423,
    n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
    n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
    n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
    n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468,
    n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477,
    n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
    n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495,
    n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504,
    n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
    n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
    n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
    n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540,
    n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549,
    n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
    n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567,
    n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
    n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
    n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
    n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
    n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612,
    n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621,
    n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
    n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639,
    n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648,
    n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
    n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
    n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
    n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684,
    n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693,
    n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
    n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711,
    n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720,
    n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729,
    n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
    n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
    n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756,
    n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765,
    n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
    n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783,
    n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792,
    n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801,
    n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
    n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
    n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828,
    n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837,
    n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
    n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855,
    n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
    n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873,
    n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
    n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
    n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900,
    n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909,
    n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
    n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927,
    n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936,
    n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945,
    n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
    n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
    n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972,
    n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
    n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999,
    n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008,
    n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
    n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
    n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
    n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044,
    n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053,
    n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
    n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071,
    n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080,
    n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089,
    n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
    n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
    n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116,
    n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125,
    n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
    n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143,
    n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
    n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161,
    n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
    n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
    n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188,
    n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197,
    n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
    n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215,
    n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224,
    n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233,
    n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
    n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
    n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260,
    n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269,
    n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
    n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287,
    n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296,
    n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
    n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
    n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
    n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332,
    n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341,
    n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
    n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359,
    n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
    n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
    n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
    n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
    n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404,
    n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413,
    n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
    n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431,
    n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440,
    n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
    n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
    n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
    n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476,
    n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485,
    n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503,
    n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521,
    n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
    n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539,
    n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548,
    n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557,
    n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
    n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575,
    n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584,
    n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593,
    n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
    n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611,
    n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620,
    n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629,
    n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
    n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647,
    n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656,
    n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665,
    n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
    n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683,
    n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692,
    n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701,
    n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
    n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719,
    n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
    n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737,
    n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
    n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755,
    n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764,
    n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773,
    n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
    n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791,
    n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
    n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
    n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
    n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
    n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836,
    n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845,
    n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
    n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863,
    n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
    n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
    n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
    n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
    n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908,
    n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917,
    n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
    n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935,
    n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
    n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
    n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
    n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989,
    n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
    n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007,
    n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
    n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
    n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
    n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
    n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052,
    n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061,
    n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
    n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079,
    n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
    n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
    n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
    n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
    n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124,
    n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133,
    n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
    n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151,
    n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
    n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
    n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
    n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
    n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196,
    n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205,
    n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
    n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223,
    n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
    n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
    n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
    n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
    n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268,
    n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277,
    n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
    n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295,
    n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
    n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
    n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
    n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
    n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340,
    n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349,
    n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
    n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367,
    n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
    n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
    n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
    n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
    n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412,
    n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
    n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
    n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439,
    n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
    n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
    n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
    n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
    n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484,
    n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493,
    n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
    n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511,
    n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
    n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
    n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
    n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
    n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556,
    n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565,
    n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
    n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583,
    n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
    n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
    n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
    n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
    n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628,
    n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637,
    n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
    n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655,
    n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
    n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
    n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
    n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
    n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700,
    n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709,
    n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
    n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727,
    n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736,
    n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
    n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
    n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
    n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772,
    n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781,
    n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790,
    n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799,
    n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808,
    n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
    n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
    n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835,
    n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844,
    n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853,
    n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862,
    n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871,
    n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
    n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
    n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
    n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
    n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916,
    n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925,
    n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934,
    n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943,
    n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952,
    n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
    n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
    n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
    n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988,
    n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997,
    n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
    n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015,
    n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
    n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
    n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
    n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051,
    n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060,
    n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069,
    n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078,
    n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087,
    n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096,
    n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
    n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
    n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123,
    n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132,
    n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141,
    n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150,
    n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159,
    n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168,
    n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
    n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
    n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195,
    n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204,
    n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213,
    n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222,
    n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231,
    n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240,
    n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
    n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
    n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267,
    n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276,
    n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285,
    n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
    n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303,
    n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
    n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
    n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
    n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
    n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348,
    n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357,
    n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366,
    n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375,
    n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384,
    n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
    n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
    n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
    n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420,
    n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429,
    n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438,
    n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447,
    n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456,
    n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
    n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
    n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
    n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492,
    n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501,
    n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510,
    n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519,
    n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528,
    n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537,
    n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
    n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
    n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564,
    n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573,
    n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
    n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591,
    n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600,
    n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609,
    n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
    n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
    n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636,
    n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645,
    n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
    n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663,
    n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
    n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
    n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
    n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
    n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708,
    n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
    n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735,
    n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744,
    n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753,
    n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
    n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
    n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780,
    n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789,
    n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798,
    n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807,
    n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816,
    n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825,
    n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
    n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
    n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852,
    n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861,
    n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
    n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879,
    n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888,
    n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897,
    n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
    n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915,
    n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924,
    n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933,
    n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942,
    n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951,
    n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960,
    n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969,
    n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
    n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
    n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996,
    n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005,
    n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014,
    n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023,
    n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032,
    n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041,
    n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
    n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059,
    n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068,
    n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077,
    n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
    n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095,
    n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104,
    n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113,
    n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
    n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131,
    n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140,
    n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149,
    n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
    n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167,
    n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176,
    n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185,
    n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
    n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203,
    n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212,
    n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221,
    n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
    n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239,
    n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
    n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
    n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
    n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
    n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284,
    n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293,
    n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
    n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311,
    n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
    n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329,
    n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
    n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347,
    n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356,
    n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365,
    n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374,
    n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383,
    n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392,
    n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401,
    n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
    n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419,
    n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428,
    n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437,
    n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446,
    n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455,
    n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
    n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473,
    n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
    n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491,
    n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500,
    n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509,
    n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
    n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527,
    n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536,
    n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545,
    n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
    n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563,
    n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572,
    n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581,
    n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
    n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599,
    n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608,
    n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617,
    n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
    n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635,
    n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644,
    n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653,
    n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
    n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671,
    n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680,
    n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689,
    n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
    n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707,
    n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716,
    n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725,
    n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734,
    n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743,
    n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752,
    n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761,
    n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
    n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
    n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788,
    n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797,
    n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806,
    n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815,
    n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824,
    n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833,
    n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
    n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851,
    n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860,
    n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869,
    n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
    n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887,
    n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896,
    n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905,
    n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
    n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923,
    n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932,
    n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941,
    n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
    n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959,
    n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
    n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977,
    n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
    n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
    n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004,
    n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013,
    n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
    n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031,
    n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
    n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049,
    n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
    n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067,
    n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076,
    n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085,
    n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094,
    n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103,
    n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112,
    n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121,
    n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
    n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139,
    n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148,
    n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157,
    n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166,
    n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175,
    n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
    n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193,
    n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
    n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211,
    n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220,
    n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229,
    n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238,
    n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247,
    n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256,
    n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265,
    n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
    n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283,
    n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292,
    n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301,
    n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310,
    n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319,
    n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
    n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337,
    n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
    n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355,
    n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364,
    n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373,
    n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382,
    n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391,
    n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400,
    n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409,
    n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
    n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
    n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436,
    n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445,
    n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
    n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463,
    n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472,
    n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481,
    n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
    n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499,
    n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508,
    n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517,
    n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
    n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535,
    n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544,
    n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553,
    n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
    n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571,
    n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580,
    n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589,
    n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
    n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607,
    n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616,
    n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625,
    n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
    n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
    n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652,
    n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661,
    n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
    n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679,
    n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688,
    n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697,
    n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
    n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715,
    n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724,
    n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733,
    n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
    n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751,
    n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
    n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769,
    n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
    n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787,
    n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796,
    n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805,
    n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
    n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823,
    n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
    n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841,
    n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
    n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859,
    n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868,
    n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877,
    n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
    n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895,
    n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904,
    n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913,
    n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
    n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
    n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940,
    n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949,
    n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
    n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967,
    n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976,
    n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985,
    n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
    n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003,
    n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012,
    n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021,
    n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
    n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039,
    n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
    n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057,
    n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
    n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
    n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084,
    n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093,
    n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
    n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111,
    n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
    n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129,
    n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
    n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147,
    n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156,
    n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165,
    n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174,
    n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183,
    n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
    n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201,
    n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
    n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219,
    n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228,
    n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237,
    n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
    n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255,
    n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
    n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273,
    n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
    n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
    n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300,
    n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309,
    n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
    n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327,
    n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
    n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345,
    n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
    n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363,
    n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372,
    n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381,
    n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390,
    n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399,
    n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
    n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417,
    n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
    n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435,
    n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444,
    n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453,
    n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462,
    n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471,
    n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
    n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489,
    n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
    n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
    n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
    n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525,
    n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534,
    n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543,
    n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
    n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561,
    n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
    n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
    n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588,
    n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597,
    n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606,
    n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615,
    n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
    n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633,
    n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
    n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
    n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660,
    n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669,
    n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678,
    n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687,
    n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696,
    n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705,
    n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
    n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723,
    n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732,
    n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741,
    n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
    n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759,
    n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768,
    n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777,
    n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
    n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795,
    n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804,
    n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813,
    n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822,
    n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831,
    n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840,
    n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
    n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
    n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867,
    n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876,
    n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885,
    n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894,
    n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903,
    n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
    n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921,
    n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
    n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939,
    n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948,
    n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957,
    n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966,
    n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975,
    n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984,
    n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993,
    n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
    n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011,
    n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020,
    n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029,
    n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
    n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047,
    n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
    n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065,
    n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
    n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083,
    n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092,
    n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101,
    n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
    n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119,
    n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
    n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137,
    n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
    n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155,
    n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164,
    n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173,
    n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182,
    n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191,
    n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200,
    n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209,
    n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
    n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227,
    n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236,
    n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245,
    n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254,
    n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263,
    n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272,
    n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281,
    n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
    n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299,
    n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308,
    n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317,
    n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326,
    n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335,
    n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
    n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353,
    n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
    n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371,
    n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380,
    n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389,
    n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398,
    n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407,
    n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
    n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425,
    n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
    n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443,
    n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452,
    n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461,
    n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470,
    n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479,
    n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488,
    n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497,
    n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
    n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515,
    n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524,
    n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533,
    n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542,
    n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551,
    n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560,
    n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569,
    n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
    n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587,
    n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
    n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605,
    n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614,
    n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623,
    n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
    n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641,
    n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
    n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659,
    n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
    n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677,
    n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686,
    n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695,
    n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704,
    n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713,
    n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
    n51723, n51724, n51725, n51726, n51727;
  assign n112 = reg_i_StoB_REQ1_out & reg_controllable_BtoS_ACK1_out;
  assign n113 = ~reg_controllable_BtoS_ACK2_out & n112;
  assign n114 = ~reg_controllable_BtoS_ACK2_out & ~n113;
  assign n115 = reg_i_StoB_REQ2_out & ~n114;
  assign n116 = ~reg_i_StoB_REQ2_out & n112;
  assign n117 = ~n115 & ~n116;
  assign n118 = sys_fair2done_out & ~n117;
  assign n119 = reg_controllable_BtoS_ACK2_out & n112;
  assign n120 = reg_controllable_BtoS_ACK2_out & ~n119;
  assign n121 = ~reg_i_StoB_REQ2_out & ~n120;
  assign n122 = ~n115 & ~n121;
  assign n123 = ~sys_fair2done_out & ~n122;
  assign n124 = ~n118 & ~n123;
  assign n125 = sys_fair1done_out & ~n124;
  assign n126 = ~reg_i_StoB_REQ1_out & ~reg_controllable_BtoS_ACK1_out;
  assign n127 = ~n112 & ~n126;
  assign n128 = ~reg_controllable_BtoS_ACK2_out & ~n127;
  assign n129 = ~reg_controllable_BtoS_ACK2_out & ~n128;
  assign n130 = reg_i_StoB_REQ2_out & ~n129;
  assign n131 = ~reg_i_StoB_REQ2_out & ~n127;
  assign n132 = ~n130 & ~n131;
  assign n133 = sys_fair2done_out & ~n132;
  assign n134 = ~n119 & ~n128;
  assign n135 = ~reg_i_StoB_REQ2_out & ~n134;
  assign n136 = ~n115 & ~n135;
  assign n137 = ~sys_fair2done_out & ~n136;
  assign n138 = ~n133 & ~n137;
  assign n139 = ~sys_fair1done_out & ~n138;
  assign n140 = ~n125 & ~n139;
  assign n141 = ~reg_controllable_BtoS_ACK3_out & ~n140;
  assign n142 = ~reg_controllable_BtoS_ACK3_out & ~n141;
  assign n143 = reg_i_StoB_REQ3_out & ~n142;
  assign n144 = ~reg_i_StoB_REQ3_out & ~n140;
  assign n145 = ~n143 & ~n144;
  assign n146 = sys_fair3done_out & ~n145;
  assign n147 = ~reg_controllable_BtoS_ACK3_out & ~n117;
  assign n148 = ~reg_controllable_BtoS_ACK3_out & ~n147;
  assign n149 = reg_i_StoB_REQ3_out & ~n148;
  assign n150 = reg_controllable_BtoS_ACK3_out & ~n117;
  assign n151 = ~sys_fair2done_out & ~n123;
  assign n152 = sys_fair1done_out & ~n151;
  assign n153 = ~n139 & ~n152;
  assign n154 = ~reg_controllable_BtoS_ACK3_out & ~n153;
  assign n155 = ~n150 & ~n154;
  assign n156 = ~reg_i_StoB_REQ3_out & ~n155;
  assign n157 = ~n149 & ~n156;
  assign n158 = ~sys_fair3done_out & ~n157;
  assign n159 = ~n146 & ~n158;
  assign n160 = ~reg_controllable_BtoS_ACK4_out & ~n159;
  assign n161 = ~reg_controllable_BtoS_ACK4_out & ~n160;
  assign n162 = reg_i_StoB_REQ4_out & ~n161;
  assign n163 = ~reg_i_StoB_REQ4_out & ~n159;
  assign n164 = ~n162 & ~n163;
  assign n165 = sys_fair4done_out & ~n164;
  assign n166 = ~reg_i_StoB_REQ3_out & ~n117;
  assign n167 = ~n149 & ~n166;
  assign n168 = ~reg_controllable_BtoS_ACK4_out & ~n167;
  assign n169 = ~reg_controllable_BtoS_ACK4_out & ~n168;
  assign n170 = reg_i_StoB_REQ4_out & ~n169;
  assign n171 = reg_controllable_BtoS_ACK4_out & ~n167;
  assign n172 = ~reg_controllable_BtoS_ACK3_out & ~n154;
  assign n173 = reg_i_StoB_REQ3_out & ~n172;
  assign n174 = ~reg_i_StoB_REQ3_out & ~n153;
  assign n175 = ~n173 & ~n174;
  assign n176 = sys_fair3done_out & ~n175;
  assign n177 = ~n158 & ~n176;
  assign n178 = ~reg_controllable_BtoS_ACK4_out & ~n177;
  assign n179 = ~n171 & ~n178;
  assign n180 = ~reg_i_StoB_REQ4_out & ~n179;
  assign n181 = ~n170 & ~n180;
  assign n182 = ~sys_fair4done_out & ~n181;
  assign n183 = ~n165 & ~n182;
  assign n184 = ~reg_controllable_BtoS_ACK5_out & ~n183;
  assign n185 = ~reg_controllable_BtoS_ACK5_out & ~n184;
  assign n186 = reg_i_StoB_REQ5_out & ~n185;
  assign n187 = ~reg_i_StoB_REQ5_out & ~n183;
  assign n188 = ~n186 & ~n187;
  assign n189 = sys_fair5done_out & ~n188;
  assign n190 = ~reg_i_StoB_REQ4_out & ~n167;
  assign n191 = ~n170 & ~n190;
  assign n192 = ~reg_controllable_BtoS_ACK5_out & ~n191;
  assign n193 = ~reg_controllable_BtoS_ACK5_out & ~n192;
  assign n194 = reg_i_StoB_REQ5_out & ~n193;
  assign n195 = reg_controllable_BtoS_ACK5_out & ~n191;
  assign n196 = ~reg_controllable_BtoS_ACK4_out & ~n178;
  assign n197 = reg_i_StoB_REQ4_out & ~n196;
  assign n198 = ~reg_i_StoB_REQ4_out & ~n177;
  assign n199 = ~n197 & ~n198;
  assign n200 = sys_fair4done_out & ~n199;
  assign n201 = ~n182 & ~n200;
  assign n202 = ~reg_controllable_BtoS_ACK5_out & ~n201;
  assign n203 = ~n195 & ~n202;
  assign n204 = ~reg_i_StoB_REQ5_out & ~n203;
  assign n205 = ~n194 & ~n204;
  assign n206 = ~sys_fair5done_out & ~n205;
  assign n207 = ~n189 & ~n206;
  assign n208 = ~reg_controllable_BtoS_ACK8_out & ~n207;
  assign n209 = ~reg_controllable_BtoS_ACK8_out & ~n208;
  assign n210 = reg_i_StoB_REQ8_out & ~n209;
  assign n211 = ~reg_i_StoB_REQ8_out & ~n207;
  assign n212 = ~n210 & ~n211;
  assign n213 = sys_fair8done_out & ~n212;
  assign n214 = ~reg_i_StoB_REQ5_out & ~n191;
  assign n215 = ~n194 & ~n214;
  assign n216 = ~reg_controllable_BtoS_ACK8_out & ~n215;
  assign n217 = ~reg_controllable_BtoS_ACK8_out & ~n216;
  assign n218 = reg_i_StoB_REQ8_out & ~n217;
  assign n219 = reg_controllable_BtoS_ACK8_out & ~n215;
  assign n220 = ~reg_controllable_BtoS_ACK5_out & ~n202;
  assign n221 = reg_i_StoB_REQ5_out & ~n220;
  assign n222 = ~reg_i_StoB_REQ5_out & ~n201;
  assign n223 = ~n221 & ~n222;
  assign n224 = sys_fair5done_out & ~n223;
  assign n225 = ~n206 & ~n224;
  assign n226 = ~reg_controllable_BtoS_ACK8_out & ~n225;
  assign n227 = ~n219 & ~n226;
  assign n228 = ~reg_i_StoB_REQ8_out & ~n227;
  assign n229 = ~n218 & ~n228;
  assign n230 = ~sys_fair8done_out & ~n229;
  assign n231 = ~n213 & ~n230;
  assign n232 = ~reg_controllable_BtoS_ACK6_out & ~n231;
  assign n233 = ~reg_controllable_BtoS_ACK6_out & ~n232;
  assign n234 = reg_i_StoB_REQ6_out & ~n233;
  assign n235 = ~reg_i_StoB_REQ6_out & ~n231;
  assign n236 = ~n234 & ~n235;
  assign n237 = sys_fair6done_out & ~n236;
  assign n238 = ~reg_i_StoB_REQ8_out & ~n215;
  assign n239 = ~n218 & ~n238;
  assign n240 = ~reg_controllable_BtoS_ACK6_out & ~n239;
  assign n241 = ~reg_controllable_BtoS_ACK6_out & ~n240;
  assign n242 = reg_i_StoB_REQ6_out & ~n241;
  assign n243 = reg_controllable_BtoS_ACK6_out & ~n239;
  assign n244 = ~reg_controllable_BtoS_ACK8_out & ~n226;
  assign n245 = reg_i_StoB_REQ8_out & ~n244;
  assign n246 = ~reg_i_StoB_REQ8_out & ~n225;
  assign n247 = ~n245 & ~n246;
  assign n248 = sys_fair8done_out & ~n247;
  assign n249 = ~n230 & ~n248;
  assign n250 = ~reg_controllable_BtoS_ACK6_out & ~n249;
  assign n251 = ~n243 & ~n250;
  assign n252 = ~reg_i_StoB_REQ6_out & ~n251;
  assign n253 = ~n242 & ~n252;
  assign n254 = ~sys_fair6done_out & ~n253;
  assign n255 = ~n237 & ~n254;
  assign n256 = sys_fair7done_out & ~n255;
  assign n257 = ~reg_i_StoB_REQ6_out & ~n239;
  assign n258 = ~n242 & ~n257;
  assign n259 = ~sys_fair7done_out & ~n258;
  assign n260 = ~n256 & ~n259;
  assign n261 = ~reg_controllable_BtoS_ACK7_out & ~n260;
  assign n262 = ~reg_controllable_BtoS_ACK7_out & ~n261;
  assign n263 = reg_i_StoB_REQ7_out & ~n262;
  assign n264 = reg_controllable_BtoS_ACK7_out & ~n260;
  assign n265 = ~reg_controllable_BtoS_ACK6_out & ~n250;
  assign n266 = reg_i_StoB_REQ6_out & ~n265;
  assign n267 = ~reg_i_StoB_REQ6_out & ~n249;
  assign n268 = ~n266 & ~n267;
  assign n269 = sys_fair6done_out & ~n268;
  assign n270 = ~n254 & ~n269;
  assign n271 = ~sys_fair7done_out & ~n270;
  assign n272 = ~n256 & ~n271;
  assign n273 = ~reg_controllable_BtoS_ACK7_out & ~n272;
  assign n274 = ~n264 & ~n273;
  assign n275 = ~reg_i_StoB_REQ7_out & ~n274;
  assign n276 = ~n263 & ~n275;
  assign n277 = ~reg_controllable_BtoS_ACK9_out & ~n276;
  assign n278 = ~reg_controllable_BtoS_ACK9_out & ~n277;
  assign n279 = reg_i_StoB_REQ9_out & ~n278;
  assign n280 = ~reg_i_StoB_REQ9_out & ~n276;
  assign n281 = ~n279 & ~n280;
  assign n282 = sys_fair9done_out & ~n281;
  assign n283 = ~reg_controllable_BtoS_ACK7_out & ~n258;
  assign n284 = ~reg_controllable_BtoS_ACK7_out & ~n283;
  assign n285 = reg_i_StoB_REQ7_out & ~n284;
  assign n286 = ~reg_i_StoB_REQ7_out & ~n258;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~reg_controllable_BtoS_ACK9_out & ~n287;
  assign n289 = ~reg_controllable_BtoS_ACK9_out & ~n288;
  assign n290 = reg_i_StoB_REQ9_out & ~n289;
  assign n291 = reg_controllable_BtoS_ACK9_out & ~n287;
  assign n292 = sys_fair7done_out & ~n270;
  assign n293 = ~n259 & ~n292;
  assign n294 = ~reg_controllable_BtoS_ACK7_out & ~n293;
  assign n295 = ~reg_controllable_BtoS_ACK7_out & ~n294;
  assign n296 = reg_i_StoB_REQ7_out & ~n295;
  assign n297 = reg_controllable_BtoS_ACK7_out & ~n293;
  assign n298 = ~reg_controllable_BtoS_ACK7_out & ~n270;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~reg_i_StoB_REQ7_out & ~n299;
  assign n301 = ~n296 & ~n300;
  assign n302 = ~reg_controllable_BtoS_ACK9_out & ~n301;
  assign n303 = ~n291 & ~n302;
  assign n304 = ~reg_i_StoB_REQ9_out & ~n303;
  assign n305 = ~n290 & ~n304;
  assign n306 = ~sys_fair9done_out & ~n305;
  assign n307 = ~n282 & ~n306;
  assign n308 = ~reg_controllable_BtoS_ACK11_out & ~n307;
  assign n309 = ~reg_controllable_BtoS_ACK11_out & ~n308;
  assign n310 = reg_i_StoB_REQ11_out & ~n309;
  assign n311 = ~reg_i_StoB_REQ11_out & ~n307;
  assign n312 = ~n310 & ~n311;
  assign n313 = sys_fair11done_out & ~n312;
  assign n314 = ~reg_i_StoB_REQ9_out & ~n287;
  assign n315 = ~n290 & ~n314;
  assign n316 = ~reg_controllable_BtoS_ACK11_out & ~n315;
  assign n317 = ~reg_controllable_BtoS_ACK11_out & ~n316;
  assign n318 = reg_i_StoB_REQ11_out & ~n317;
  assign n319 = reg_controllable_BtoS_ACK11_out & ~n315;
  assign n320 = ~reg_controllable_BtoS_ACK9_out & ~n302;
  assign n321 = reg_i_StoB_REQ9_out & ~n320;
  assign n322 = ~reg_i_StoB_REQ9_out & ~n301;
  assign n323 = ~n321 & ~n322;
  assign n324 = sys_fair9done_out & ~n323;
  assign n325 = ~n306 & ~n324;
  assign n326 = ~reg_controllable_BtoS_ACK11_out & ~n325;
  assign n327 = ~n319 & ~n326;
  assign n328 = ~reg_i_StoB_REQ11_out & ~n327;
  assign n329 = ~n318 & ~n328;
  assign n330 = ~sys_fair11done_out & ~n329;
  assign n331 = ~n313 & ~n330;
  assign n332 = sys_fair12done_out & ~n331;
  assign n333 = ~reg_i_StoB_REQ11_out & ~n315;
  assign n334 = ~n318 & ~n333;
  assign n335 = ~sys_fair12done_out & ~n334;
  assign n336 = ~n332 & ~n335;
  assign n337 = ~reg_controllable_BtoS_ACK12_out & ~n336;
  assign n338 = ~reg_controllable_BtoS_ACK12_out & ~n337;
  assign n339 = reg_i_StoB_REQ12_out & ~n338;
  assign n340 = reg_controllable_BtoS_ACK12_out & ~n336;
  assign n341 = ~reg_controllable_BtoS_ACK11_out & ~n326;
  assign n342 = reg_i_StoB_REQ11_out & ~n341;
  assign n343 = ~reg_i_StoB_REQ11_out & ~n325;
  assign n344 = ~n342 & ~n343;
  assign n345 = sys_fair11done_out & ~n344;
  assign n346 = ~n330 & ~n345;
  assign n347 = ~sys_fair12done_out & ~n346;
  assign n348 = ~n332 & ~n347;
  assign n349 = ~reg_controllable_BtoS_ACK12_out & ~n348;
  assign n350 = ~n340 & ~n349;
  assign n351 = ~reg_i_StoB_REQ12_out & ~n350;
  assign n352 = ~n339 & ~n351;
  assign n353 = ~reg_controllable_BtoS_ACK13_out & ~n352;
  assign n354 = ~reg_controllable_BtoS_ACK13_out & ~n353;
  assign n355 = reg_i_StoB_REQ13_out & ~n354;
  assign n356 = ~reg_i_StoB_REQ13_out & ~n352;
  assign n357 = ~n355 & ~n356;
  assign n358 = sys_fair13done_out & ~n357;
  assign n359 = ~reg_controllable_BtoS_ACK12_out & ~n334;
  assign n360 = ~reg_controllable_BtoS_ACK12_out & ~n359;
  assign n361 = reg_i_StoB_REQ12_out & ~n360;
  assign n362 = ~reg_i_StoB_REQ12_out & ~n334;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~reg_controllable_BtoS_ACK13_out & ~n363;
  assign n365 = ~reg_controllable_BtoS_ACK13_out & ~n364;
  assign n366 = reg_i_StoB_REQ13_out & ~n365;
  assign n367 = reg_controllable_BtoS_ACK13_out & ~n363;
  assign n368 = sys_fair12done_out & ~n346;
  assign n369 = ~n335 & ~n368;
  assign n370 = ~reg_controllable_BtoS_ACK12_out & ~n369;
  assign n371 = ~reg_controllable_BtoS_ACK12_out & ~n370;
  assign n372 = reg_i_StoB_REQ12_out & ~n371;
  assign n373 = reg_controllable_BtoS_ACK12_out & ~n369;
  assign n374 = ~reg_controllable_BtoS_ACK12_out & ~n346;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~reg_i_StoB_REQ12_out & ~n375;
  assign n377 = ~n372 & ~n376;
  assign n378 = ~reg_controllable_BtoS_ACK13_out & ~n377;
  assign n379 = ~n367 & ~n378;
  assign n380 = ~reg_i_StoB_REQ13_out & ~n379;
  assign n381 = ~n366 & ~n380;
  assign n382 = ~sys_fair13done_out & ~n381;
  assign n383 = ~n358 & ~n382;
  assign n384 = sys_fair0done_out & ~n383;
  assign n385 = ~reg_i_StoB_REQ13_out & ~n363;
  assign n386 = ~n366 & ~n385;
  assign n387 = ~sys_fair0done_out & ~n386;
  assign n388 = ~n384 & ~n387;
  assign n389 = ~reg_controllable_BtoS_ACK0_out & ~n388;
  assign n390 = ~reg_controllable_BtoS_ACK0_out & ~n389;
  assign n391 = reg_i_StoB_REQ0_out & ~n390;
  assign n392 = reg_controllable_BtoS_ACK0_out & ~n388;
  assign n393 = ~reg_controllable_BtoS_ACK13_out & ~n378;
  assign n394 = reg_i_StoB_REQ13_out & ~n393;
  assign n395 = ~reg_i_StoB_REQ13_out & ~n377;
  assign n396 = ~n394 & ~n395;
  assign n397 = sys_fair13done_out & ~n396;
  assign n398 = ~n382 & ~n397;
  assign n399 = ~sys_fair0done_out & ~n398;
  assign n400 = ~n384 & ~n399;
  assign n401 = ~reg_controllable_BtoS_ACK0_out & ~n400;
  assign n402 = ~n392 & ~n401;
  assign n403 = ~reg_i_StoB_REQ0_out & ~n402;
  assign n404 = ~n391 & ~n403;
  assign n405 = ~reg_controllable_BtoS_ACK10_out & ~n404;
  assign n406 = ~reg_controllable_BtoS_ACK10_out & ~n405;
  assign n407 = reg_i_StoB_REQ10_out & ~n406;
  assign n408 = ~reg_i_StoB_REQ10_out & ~n404;
  assign n409 = ~n407 & ~n408;
  assign n410 = sys_fair10done_out & ~n409;
  assign n411 = ~reg_controllable_BtoS_ACK0_out & ~n386;
  assign n412 = ~reg_controllable_BtoS_ACK0_out & ~n411;
  assign n413 = reg_i_StoB_REQ0_out & ~n412;
  assign n414 = ~reg_i_StoB_REQ0_out & ~n386;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~reg_controllable_BtoS_ACK10_out & ~n415;
  assign n417 = ~reg_controllable_BtoS_ACK10_out & ~n416;
  assign n418 = reg_i_StoB_REQ10_out & ~n417;
  assign n419 = reg_controllable_BtoS_ACK10_out & ~n415;
  assign n420 = sys_fair0done_out & ~n398;
  assign n421 = ~n387 & ~n420;
  assign n422 = ~reg_controllable_BtoS_ACK0_out & ~n421;
  assign n423 = ~reg_controllable_BtoS_ACK0_out & ~n422;
  assign n424 = reg_i_StoB_REQ0_out & ~n423;
  assign n425 = reg_controllable_BtoS_ACK0_out & ~n421;
  assign n426 = ~reg_controllable_BtoS_ACK0_out & ~n398;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~reg_i_StoB_REQ0_out & ~n427;
  assign n429 = ~n424 & ~n428;
  assign n430 = ~reg_controllable_BtoS_ACK10_out & ~n429;
  assign n431 = ~n419 & ~n430;
  assign n432 = ~reg_i_StoB_REQ10_out & ~n431;
  assign n433 = ~n418 & ~n432;
  assign n434 = ~sys_fair10done_out & ~n433;
  assign n435 = ~n410 & ~n434;
  assign n436 = ~reg_controllable_BtoS_ACK14_out & ~n435;
  assign n437 = ~reg_controllable_BtoS_ACK14_out & ~n436;
  assign n438 = reg_i_StoB_REQ14_out & ~n437;
  assign n439 = ~reg_controllable_BtoS_ACK1_out & ~n126;
  assign n440 = ~reg_i_StoB_REQ2_out & ~n439;
  assign n441 = ~n115 & ~n440;
  assign n442 = sys_fair2done_out & ~n441;
  assign n443 = reg_controllable_BtoS_ACK2_out & ~n439;
  assign n444 = reg_controllable_BtoS_ACK2_out & ~n443;
  assign n445 = ~reg_i_StoB_REQ2_out & ~n444;
  assign n446 = ~n115 & ~n445;
  assign n447 = ~sys_fair2done_out & ~n446;
  assign n448 = ~n442 & ~n447;
  assign n449 = sys_fair1done_out & ~n448;
  assign n450 = ~n130 & ~n440;
  assign n451 = sys_fair2done_out & ~n450;
  assign n452 = ~sys_fair2done_out & ~n441;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~sys_fair1done_out & ~n453;
  assign n455 = ~n449 & ~n454;
  assign n456 = ~reg_i_StoB_REQ3_out & ~n455;
  assign n457 = ~n143 & ~n456;
  assign n458 = sys_fair3done_out & ~n457;
  assign n459 = reg_controllable_BtoS_ACK3_out & ~n441;
  assign n460 = ~sys_fair2done_out & ~n447;
  assign n461 = sys_fair1done_out & ~n460;
  assign n462 = ~n454 & ~n461;
  assign n463 = ~reg_controllable_BtoS_ACK3_out & ~n462;
  assign n464 = ~n459 & ~n463;
  assign n465 = ~reg_i_StoB_REQ3_out & ~n464;
  assign n466 = ~n149 & ~n465;
  assign n467 = ~sys_fair3done_out & ~n466;
  assign n468 = ~n458 & ~n467;
  assign n469 = ~reg_i_StoB_REQ4_out & ~n468;
  assign n470 = ~n162 & ~n469;
  assign n471 = sys_fair4done_out & ~n470;
  assign n472 = ~reg_i_StoB_REQ3_out & ~n441;
  assign n473 = ~n149 & ~n472;
  assign n474 = reg_controllable_BtoS_ACK4_out & ~n473;
  assign n475 = ~reg_i_StoB_REQ3_out & ~n462;
  assign n476 = ~n173 & ~n475;
  assign n477 = sys_fair3done_out & ~n476;
  assign n478 = ~n467 & ~n477;
  assign n479 = ~reg_controllable_BtoS_ACK4_out & ~n478;
  assign n480 = ~n474 & ~n479;
  assign n481 = ~reg_i_StoB_REQ4_out & ~n480;
  assign n482 = ~n170 & ~n481;
  assign n483 = ~sys_fair4done_out & ~n482;
  assign n484 = ~n471 & ~n483;
  assign n485 = ~reg_i_StoB_REQ5_out & ~n484;
  assign n486 = ~n186 & ~n485;
  assign n487 = sys_fair5done_out & ~n486;
  assign n488 = ~reg_i_StoB_REQ4_out & ~n473;
  assign n489 = ~n170 & ~n488;
  assign n490 = reg_controllable_BtoS_ACK5_out & ~n489;
  assign n491 = ~reg_i_StoB_REQ4_out & ~n478;
  assign n492 = ~n197 & ~n491;
  assign n493 = sys_fair4done_out & ~n492;
  assign n494 = ~n483 & ~n493;
  assign n495 = ~reg_controllable_BtoS_ACK5_out & ~n494;
  assign n496 = ~n490 & ~n495;
  assign n497 = ~reg_i_StoB_REQ5_out & ~n496;
  assign n498 = ~n194 & ~n497;
  assign n499 = ~sys_fair5done_out & ~n498;
  assign n500 = ~n487 & ~n499;
  assign n501 = ~reg_i_StoB_REQ8_out & ~n500;
  assign n502 = ~n210 & ~n501;
  assign n503 = sys_fair8done_out & ~n502;
  assign n504 = ~reg_i_StoB_REQ5_out & ~n489;
  assign n505 = ~n194 & ~n504;
  assign n506 = reg_controllable_BtoS_ACK8_out & ~n505;
  assign n507 = ~reg_i_StoB_REQ5_out & ~n494;
  assign n508 = ~n221 & ~n507;
  assign n509 = sys_fair5done_out & ~n508;
  assign n510 = ~n499 & ~n509;
  assign n511 = ~reg_controllable_BtoS_ACK8_out & ~n510;
  assign n512 = ~n506 & ~n511;
  assign n513 = ~reg_i_StoB_REQ8_out & ~n512;
  assign n514 = ~n218 & ~n513;
  assign n515 = ~sys_fair8done_out & ~n514;
  assign n516 = ~n503 & ~n515;
  assign n517 = ~reg_i_StoB_REQ6_out & ~n516;
  assign n518 = ~n234 & ~n517;
  assign n519 = sys_fair6done_out & ~n518;
  assign n520 = ~reg_i_StoB_REQ8_out & ~n505;
  assign n521 = ~n218 & ~n520;
  assign n522 = reg_controllable_BtoS_ACK6_out & ~n521;
  assign n523 = ~reg_i_StoB_REQ8_out & ~n510;
  assign n524 = ~n245 & ~n523;
  assign n525 = sys_fair8done_out & ~n524;
  assign n526 = ~n515 & ~n525;
  assign n527 = ~reg_controllable_BtoS_ACK6_out & ~n526;
  assign n528 = ~n522 & ~n527;
  assign n529 = ~reg_i_StoB_REQ6_out & ~n528;
  assign n530 = ~n242 & ~n529;
  assign n531 = ~sys_fair6done_out & ~n530;
  assign n532 = ~n519 & ~n531;
  assign n533 = sys_fair7done_out & ~n532;
  assign n534 = ~reg_i_StoB_REQ6_out & ~n521;
  assign n535 = ~n242 & ~n534;
  assign n536 = ~sys_fair7done_out & ~n535;
  assign n537 = ~n533 & ~n536;
  assign n538 = reg_controllable_BtoS_ACK7_out & ~n537;
  assign n539 = ~reg_i_StoB_REQ6_out & ~n526;
  assign n540 = ~n266 & ~n539;
  assign n541 = sys_fair6done_out & ~n540;
  assign n542 = ~n531 & ~n541;
  assign n543 = ~sys_fair7done_out & ~n542;
  assign n544 = ~n533 & ~n543;
  assign n545 = ~reg_controllable_BtoS_ACK7_out & ~n544;
  assign n546 = ~n538 & ~n545;
  assign n547 = ~reg_i_StoB_REQ7_out & ~n546;
  assign n548 = ~n263 & ~n547;
  assign n549 = ~reg_i_StoB_REQ9_out & ~n548;
  assign n550 = ~n279 & ~n549;
  assign n551 = sys_fair9done_out & ~n550;
  assign n552 = ~reg_i_StoB_REQ7_out & ~n535;
  assign n553 = ~n285 & ~n552;
  assign n554 = reg_controllable_BtoS_ACK9_out & ~n553;
  assign n555 = sys_fair7done_out & ~n542;
  assign n556 = ~n536 & ~n555;
  assign n557 = reg_controllable_BtoS_ACK7_out & ~n556;
  assign n558 = ~reg_controllable_BtoS_ACK7_out & ~n542;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~reg_i_StoB_REQ7_out & ~n559;
  assign n561 = ~n296 & ~n560;
  assign n562 = ~reg_controllable_BtoS_ACK9_out & ~n561;
  assign n563 = ~n554 & ~n562;
  assign n564 = ~reg_i_StoB_REQ9_out & ~n563;
  assign n565 = ~n290 & ~n564;
  assign n566 = ~sys_fair9done_out & ~n565;
  assign n567 = ~n551 & ~n566;
  assign n568 = ~reg_i_StoB_REQ11_out & ~n567;
  assign n569 = ~n310 & ~n568;
  assign n570 = sys_fair11done_out & ~n569;
  assign n571 = ~reg_i_StoB_REQ9_out & ~n553;
  assign n572 = ~n290 & ~n571;
  assign n573 = reg_controllable_BtoS_ACK11_out & ~n572;
  assign n574 = ~reg_i_StoB_REQ9_out & ~n561;
  assign n575 = ~n321 & ~n574;
  assign n576 = sys_fair9done_out & ~n575;
  assign n577 = ~n566 & ~n576;
  assign n578 = ~reg_controllable_BtoS_ACK11_out & ~n577;
  assign n579 = ~n573 & ~n578;
  assign n580 = ~reg_i_StoB_REQ11_out & ~n579;
  assign n581 = ~n318 & ~n580;
  assign n582 = ~sys_fair11done_out & ~n581;
  assign n583 = ~n570 & ~n582;
  assign n584 = sys_fair12done_out & ~n583;
  assign n585 = ~reg_i_StoB_REQ11_out & ~n572;
  assign n586 = ~n318 & ~n585;
  assign n587 = ~sys_fair12done_out & ~n586;
  assign n588 = ~n584 & ~n587;
  assign n589 = reg_controllable_BtoS_ACK12_out & ~n588;
  assign n590 = ~reg_i_StoB_REQ11_out & ~n577;
  assign n591 = ~n342 & ~n590;
  assign n592 = sys_fair11done_out & ~n591;
  assign n593 = ~n582 & ~n592;
  assign n594 = ~sys_fair12done_out & ~n593;
  assign n595 = ~n584 & ~n594;
  assign n596 = ~reg_controllable_BtoS_ACK12_out & ~n595;
  assign n597 = ~n589 & ~n596;
  assign n598 = ~reg_i_StoB_REQ12_out & ~n597;
  assign n599 = ~n339 & ~n598;
  assign n600 = ~reg_i_StoB_REQ13_out & ~n599;
  assign n601 = ~n355 & ~n600;
  assign n602 = sys_fair13done_out & ~n601;
  assign n603 = ~reg_i_StoB_REQ12_out & ~n586;
  assign n604 = ~n361 & ~n603;
  assign n605 = reg_controllable_BtoS_ACK13_out & ~n604;
  assign n606 = sys_fair12done_out & ~n593;
  assign n607 = ~n587 & ~n606;
  assign n608 = reg_controllable_BtoS_ACK12_out & ~n607;
  assign n609 = ~reg_controllable_BtoS_ACK12_out & ~n593;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~reg_i_StoB_REQ12_out & ~n610;
  assign n612 = ~n372 & ~n611;
  assign n613 = ~reg_controllable_BtoS_ACK13_out & ~n612;
  assign n614 = ~n605 & ~n613;
  assign n615 = ~reg_i_StoB_REQ13_out & ~n614;
  assign n616 = ~n366 & ~n615;
  assign n617 = ~sys_fair13done_out & ~n616;
  assign n618 = ~n602 & ~n617;
  assign n619 = sys_fair0done_out & ~n618;
  assign n620 = ~reg_i_StoB_REQ13_out & ~n604;
  assign n621 = ~n366 & ~n620;
  assign n622 = ~sys_fair0done_out & ~n621;
  assign n623 = ~n619 & ~n622;
  assign n624 = reg_controllable_BtoS_ACK0_out & ~n623;
  assign n625 = ~reg_i_StoB_REQ13_out & ~n612;
  assign n626 = ~n394 & ~n625;
  assign n627 = sys_fair13done_out & ~n626;
  assign n628 = ~n617 & ~n627;
  assign n629 = ~sys_fair0done_out & ~n628;
  assign n630 = ~n619 & ~n629;
  assign n631 = ~reg_controllable_BtoS_ACK0_out & ~n630;
  assign n632 = ~n624 & ~n631;
  assign n633 = ~reg_i_StoB_REQ0_out & ~n632;
  assign n634 = ~n391 & ~n633;
  assign n635 = ~reg_i_StoB_REQ10_out & ~n634;
  assign n636 = ~n407 & ~n635;
  assign n637 = sys_fair10done_out & ~n636;
  assign n638 = ~reg_i_StoB_REQ0_out & ~n621;
  assign n639 = ~n413 & ~n638;
  assign n640 = reg_controllable_BtoS_ACK10_out & ~n639;
  assign n641 = sys_fair0done_out & ~n628;
  assign n642 = ~n622 & ~n641;
  assign n643 = reg_controllable_BtoS_ACK0_out & ~n642;
  assign n644 = ~reg_controllable_BtoS_ACK0_out & ~n628;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~reg_i_StoB_REQ0_out & ~n645;
  assign n647 = ~n424 & ~n646;
  assign n648 = ~reg_controllable_BtoS_ACK10_out & ~n647;
  assign n649 = ~n640 & ~n648;
  assign n650 = ~reg_i_StoB_REQ10_out & ~n649;
  assign n651 = ~n418 & ~n650;
  assign n652 = ~sys_fair10done_out & ~n651;
  assign n653 = ~n637 & ~n652;
  assign n654 = ~reg_i_StoB_REQ14_out & ~n653;
  assign n655 = ~n438 & ~n654;
  assign n656 = sys_fair14done_out & ~n655;
  assign n657 = ~reg_i_StoB_REQ10_out & ~n415;
  assign n658 = ~n418 & ~n657;
  assign n659 = ~reg_controllable_BtoS_ACK14_out & ~n658;
  assign n660 = ~reg_controllable_BtoS_ACK14_out & ~n659;
  assign n661 = reg_i_StoB_REQ14_out & ~n660;
  assign n662 = ~reg_i_StoB_REQ10_out & ~n639;
  assign n663 = ~n418 & ~n662;
  assign n664 = reg_controllable_BtoS_ACK14_out & ~n663;
  assign n665 = ~reg_controllable_BtoS_ACK10_out & ~n430;
  assign n666 = reg_i_StoB_REQ10_out & ~n665;
  assign n667 = ~reg_i_StoB_REQ10_out & ~n647;
  assign n668 = ~n666 & ~n667;
  assign n669 = sys_fair10done_out & ~n668;
  assign n670 = ~n652 & ~n669;
  assign n671 = ~reg_controllable_BtoS_ACK14_out & ~n670;
  assign n672 = ~n664 & ~n671;
  assign n673 = ~reg_i_StoB_REQ14_out & ~n672;
  assign n674 = ~n661 & ~n673;
  assign n675 = ~sys_fair14done_out & ~n674;
  assign n676 = ~n656 & ~n675;
  assign n677 = sys_fair15done_out & ~n676;
  assign n678 = ~reg_i_StoB_REQ10_out & ~n429;
  assign n679 = ~n666 & ~n678;
  assign n680 = sys_fair10done_out & ~n679;
  assign n681 = ~n434 & ~n680;
  assign n682 = ~reg_controllable_BtoS_ACK14_out & ~n681;
  assign n683 = ~reg_controllable_BtoS_ACK14_out & ~n682;
  assign n684 = reg_i_StoB_REQ14_out & ~n683;
  assign n685 = ~reg_i_StoB_REQ14_out & ~n670;
  assign n686 = ~n684 & ~n685;
  assign n687 = sys_fair14done_out & ~n686;
  assign n688 = ~n675 & ~n687;
  assign n689 = reg_stateG12_out & ~n688;
  assign n690 = ~reg_i_StoB_REQ14_out & ~n663;
  assign n691 = ~n661 & ~n690;
  assign n692 = ~reg_stateG12_out & ~n691;
  assign n693 = ~n689 & ~n692;
  assign n694 = ~sys_fair15done_out & ~n693;
  assign n695 = ~n677 & ~n694;
  assign n696 = fair_cnt<1>_out  & ~n695;
  assign n697 = ~fair_cnt<1>_out  & ~n691;
  assign n698 = ~n696 & ~n697;
  assign n699 = fair_cnt<0>_out  & ~n698;
  assign n700 = ~fair_cnt<0>_out  & ~n691;
  assign n701 = ~n699 & ~n700;
  assign n702 = env_fair1done_out & ~n701;
  assign n703 = ~sys_fair15done_out & ~n691;
  assign n704 = ~n677 & ~n703;
  assign n705 = fair_cnt<1>_out  & ~n704;
  assign n706 = ~n697 & ~n705;
  assign n707 = fair_cnt<0>_out  & ~n706;
  assign n708 = ~n700 & ~n707;
  assign n709 = ~env_fair1done_out & ~n708;
  assign n710 = ~n702 & ~n709;
  assign n711 = reg_i_RtoB_ACK1_out & ~n710;
  assign n712 = ~reg_i_StoB_REQ2_out & ~n121;
  assign n713 = ~sys_fair2done_out & ~n712;
  assign n714 = ~n118 & ~n713;
  assign n715 = sys_fair1done_out & ~n714;
  assign n716 = reg_controllable_BtoS_ACK1_out & ~n112;
  assign n717 = ~reg_controllable_BtoS_ACK2_out & ~n716;
  assign n718 = ~reg_controllable_BtoS_ACK2_out & ~n717;
  assign n719 = reg_i_StoB_REQ2_out & ~n718;
  assign n720 = ~reg_i_StoB_REQ2_out & ~n716;
  assign n721 = ~n719 & ~n720;
  assign n722 = sys_fair2done_out & ~n721;
  assign n723 = ~n119 & ~n717;
  assign n724 = ~reg_i_StoB_REQ2_out & ~n723;
  assign n725 = ~n719 & ~n724;
  assign n726 = ~sys_fair2done_out & ~n725;
  assign n727 = ~n722 & ~n726;
  assign n728 = ~sys_fair1done_out & ~n727;
  assign n729 = ~n715 & ~n728;
  assign n730 = ~reg_controllable_BtoS_ACK3_out & ~n729;
  assign n731 = ~reg_controllable_BtoS_ACK3_out & ~n730;
  assign n732 = reg_i_StoB_REQ3_out & ~n731;
  assign n733 = ~reg_i_StoB_REQ3_out & ~n729;
  assign n734 = ~n732 & ~n733;
  assign n735 = sys_fair3done_out & ~n734;
  assign n736 = ~sys_fair2done_out & ~n713;
  assign n737 = sys_fair1done_out & ~n736;
  assign n738 = ~n728 & ~n737;
  assign n739 = ~reg_controllable_BtoS_ACK3_out & ~n738;
  assign n740 = ~reg_controllable_BtoS_ACK3_out & ~n739;
  assign n741 = reg_i_StoB_REQ3_out & ~n740;
  assign n742 = ~n150 & ~n739;
  assign n743 = ~reg_i_StoB_REQ3_out & ~n742;
  assign n744 = ~n741 & ~n743;
  assign n745 = ~sys_fair3done_out & ~n744;
  assign n746 = ~n735 & ~n745;
  assign n747 = ~reg_controllable_BtoS_ACK4_out & ~n746;
  assign n748 = ~reg_controllable_BtoS_ACK4_out & ~n747;
  assign n749 = reg_i_StoB_REQ4_out & ~n748;
  assign n750 = ~reg_i_StoB_REQ4_out & ~n746;
  assign n751 = ~n749 & ~n750;
  assign n752 = sys_fair4done_out & ~n751;
  assign n753 = ~reg_i_StoB_REQ3_out & ~n738;
  assign n754 = ~n741 & ~n753;
  assign n755 = sys_fair3done_out & ~n754;
  assign n756 = ~n745 & ~n755;
  assign n757 = ~reg_controllable_BtoS_ACK4_out & ~n756;
  assign n758 = ~reg_controllable_BtoS_ACK4_out & ~n757;
  assign n759 = reg_i_StoB_REQ4_out & ~n758;
  assign n760 = ~n171 & ~n757;
  assign n761 = ~reg_i_StoB_REQ4_out & ~n760;
  assign n762 = ~n759 & ~n761;
  assign n763 = ~sys_fair4done_out & ~n762;
  assign n764 = ~n752 & ~n763;
  assign n765 = ~reg_controllable_BtoS_ACK5_out & ~n764;
  assign n766 = ~reg_controllable_BtoS_ACK5_out & ~n765;
  assign n767 = reg_i_StoB_REQ5_out & ~n766;
  assign n768 = ~reg_i_StoB_REQ5_out & ~n764;
  assign n769 = ~n767 & ~n768;
  assign n770 = sys_fair5done_out & ~n769;
  assign n771 = ~reg_i_StoB_REQ4_out & ~n756;
  assign n772 = ~n759 & ~n771;
  assign n773 = sys_fair4done_out & ~n772;
  assign n774 = ~n763 & ~n773;
  assign n775 = ~reg_controllable_BtoS_ACK5_out & ~n774;
  assign n776 = ~reg_controllable_BtoS_ACK5_out & ~n775;
  assign n777 = reg_i_StoB_REQ5_out & ~n776;
  assign n778 = ~n195 & ~n775;
  assign n779 = ~reg_i_StoB_REQ5_out & ~n778;
  assign n780 = ~n777 & ~n779;
  assign n781 = ~sys_fair5done_out & ~n780;
  assign n782 = ~n770 & ~n781;
  assign n783 = ~reg_controllable_BtoS_ACK8_out & ~n782;
  assign n784 = ~reg_controllable_BtoS_ACK8_out & ~n783;
  assign n785 = reg_i_StoB_REQ8_out & ~n784;
  assign n786 = ~reg_i_StoB_REQ8_out & ~n782;
  assign n787 = ~n785 & ~n786;
  assign n788 = sys_fair8done_out & ~n787;
  assign n789 = ~reg_i_StoB_REQ5_out & ~n774;
  assign n790 = ~n777 & ~n789;
  assign n791 = sys_fair5done_out & ~n790;
  assign n792 = ~n781 & ~n791;
  assign n793 = ~reg_controllable_BtoS_ACK8_out & ~n792;
  assign n794 = ~reg_controllable_BtoS_ACK8_out & ~n793;
  assign n795 = reg_i_StoB_REQ8_out & ~n794;
  assign n796 = ~n219 & ~n793;
  assign n797 = ~reg_i_StoB_REQ8_out & ~n796;
  assign n798 = ~n795 & ~n797;
  assign n799 = ~sys_fair8done_out & ~n798;
  assign n800 = ~n788 & ~n799;
  assign n801 = ~reg_controllable_BtoS_ACK6_out & ~n800;
  assign n802 = ~reg_controllable_BtoS_ACK6_out & ~n801;
  assign n803 = reg_i_StoB_REQ6_out & ~n802;
  assign n804 = ~reg_i_StoB_REQ6_out & ~n800;
  assign n805 = ~n803 & ~n804;
  assign n806 = sys_fair6done_out & ~n805;
  assign n807 = ~reg_i_StoB_REQ8_out & ~n792;
  assign n808 = ~n795 & ~n807;
  assign n809 = sys_fair8done_out & ~n808;
  assign n810 = ~n799 & ~n809;
  assign n811 = ~reg_controllable_BtoS_ACK6_out & ~n810;
  assign n812 = ~reg_controllable_BtoS_ACK6_out & ~n811;
  assign n813 = reg_i_StoB_REQ6_out & ~n812;
  assign n814 = ~n243 & ~n811;
  assign n815 = ~reg_i_StoB_REQ6_out & ~n814;
  assign n816 = ~n813 & ~n815;
  assign n817 = ~sys_fair6done_out & ~n816;
  assign n818 = ~n806 & ~n817;
  assign n819 = sys_fair7done_out & ~n818;
  assign n820 = ~reg_i_StoB_REQ6_out & ~n810;
  assign n821 = ~n813 & ~n820;
  assign n822 = sys_fair6done_out & ~n821;
  assign n823 = ~n817 & ~n822;
  assign n824 = ~sys_fair7done_out & ~n823;
  assign n825 = ~n819 & ~n824;
  assign n826 = ~reg_controllable_BtoS_ACK7_out & ~n825;
  assign n827 = ~reg_controllable_BtoS_ACK7_out & ~n826;
  assign n828 = reg_i_StoB_REQ7_out & ~n827;
  assign n829 = ~n259 & ~n819;
  assign n830 = reg_controllable_BtoS_ACK7_out & ~n829;
  assign n831 = ~n826 & ~n830;
  assign n832 = ~reg_i_StoB_REQ7_out & ~n831;
  assign n833 = ~n828 & ~n832;
  assign n834 = ~reg_controllable_BtoS_ACK9_out & ~n833;
  assign n835 = ~reg_controllable_BtoS_ACK9_out & ~n834;
  assign n836 = reg_i_StoB_REQ9_out & ~n835;
  assign n837 = ~reg_i_StoB_REQ9_out & ~n833;
  assign n838 = ~n836 & ~n837;
  assign n839 = sys_fair9done_out & ~n838;
  assign n840 = ~reg_controllable_BtoS_ACK7_out & ~n823;
  assign n841 = ~reg_controllable_BtoS_ACK7_out & ~n840;
  assign n842 = reg_i_StoB_REQ7_out & ~n841;
  assign n843 = sys_fair7done_out & ~n823;
  assign n844 = ~n259 & ~n843;
  assign n845 = reg_controllable_BtoS_ACK7_out & ~n844;
  assign n846 = ~n840 & ~n845;
  assign n847 = ~reg_i_StoB_REQ7_out & ~n846;
  assign n848 = ~n842 & ~n847;
  assign n849 = ~reg_controllable_BtoS_ACK9_out & ~n848;
  assign n850 = ~reg_controllable_BtoS_ACK9_out & ~n849;
  assign n851 = reg_i_StoB_REQ9_out & ~n850;
  assign n852 = ~n291 & ~n849;
  assign n853 = ~reg_i_StoB_REQ9_out & ~n852;
  assign n854 = ~n851 & ~n853;
  assign n855 = ~sys_fair9done_out & ~n854;
  assign n856 = ~n839 & ~n855;
  assign n857 = ~reg_controllable_BtoS_ACK11_out & ~n856;
  assign n858 = ~reg_controllable_BtoS_ACK11_out & ~n857;
  assign n859 = reg_i_StoB_REQ11_out & ~n858;
  assign n860 = ~reg_i_StoB_REQ11_out & ~n856;
  assign n861 = ~n859 & ~n860;
  assign n862 = sys_fair11done_out & ~n861;
  assign n863 = ~reg_i_StoB_REQ9_out & ~n848;
  assign n864 = ~n851 & ~n863;
  assign n865 = sys_fair9done_out & ~n864;
  assign n866 = ~n855 & ~n865;
  assign n867 = ~reg_controllable_BtoS_ACK11_out & ~n866;
  assign n868 = ~reg_controllable_BtoS_ACK11_out & ~n867;
  assign n869 = reg_i_StoB_REQ11_out & ~n868;
  assign n870 = ~n319 & ~n867;
  assign n871 = ~reg_i_StoB_REQ11_out & ~n870;
  assign n872 = ~n869 & ~n871;
  assign n873 = ~sys_fair11done_out & ~n872;
  assign n874 = ~n862 & ~n873;
  assign n875 = sys_fair12done_out & ~n874;
  assign n876 = ~reg_i_StoB_REQ11_out & ~n866;
  assign n877 = ~n869 & ~n876;
  assign n878 = sys_fair11done_out & ~n877;
  assign n879 = ~n873 & ~n878;
  assign n880 = ~sys_fair12done_out & ~n879;
  assign n881 = ~n875 & ~n880;
  assign n882 = ~reg_controllable_BtoS_ACK12_out & ~n881;
  assign n883 = ~reg_controllable_BtoS_ACK12_out & ~n882;
  assign n884 = reg_i_StoB_REQ12_out & ~n883;
  assign n885 = ~n335 & ~n875;
  assign n886 = reg_controllable_BtoS_ACK12_out & ~n885;
  assign n887 = ~n882 & ~n886;
  assign n888 = ~reg_i_StoB_REQ12_out & ~n887;
  assign n889 = ~n884 & ~n888;
  assign n890 = ~reg_controllable_BtoS_ACK13_out & ~n889;
  assign n891 = ~reg_controllable_BtoS_ACK13_out & ~n890;
  assign n892 = reg_i_StoB_REQ13_out & ~n891;
  assign n893 = ~reg_i_StoB_REQ13_out & ~n889;
  assign n894 = ~n892 & ~n893;
  assign n895 = sys_fair13done_out & ~n894;
  assign n896 = ~reg_controllable_BtoS_ACK12_out & ~n879;
  assign n897 = ~reg_controllable_BtoS_ACK12_out & ~n896;
  assign n898 = reg_i_StoB_REQ12_out & ~n897;
  assign n899 = sys_fair12done_out & ~n879;
  assign n900 = ~n335 & ~n899;
  assign n901 = reg_controllable_BtoS_ACK12_out & ~n900;
  assign n902 = ~n896 & ~n901;
  assign n903 = ~reg_i_StoB_REQ12_out & ~n902;
  assign n904 = ~n898 & ~n903;
  assign n905 = ~reg_controllable_BtoS_ACK13_out & ~n904;
  assign n906 = ~reg_controllable_BtoS_ACK13_out & ~n905;
  assign n907 = reg_i_StoB_REQ13_out & ~n906;
  assign n908 = ~n367 & ~n905;
  assign n909 = ~reg_i_StoB_REQ13_out & ~n908;
  assign n910 = ~n907 & ~n909;
  assign n911 = ~sys_fair13done_out & ~n910;
  assign n912 = ~n895 & ~n911;
  assign n913 = sys_fair0done_out & ~n912;
  assign n914 = ~reg_i_StoB_REQ13_out & ~n904;
  assign n915 = ~n907 & ~n914;
  assign n916 = sys_fair13done_out & ~n915;
  assign n917 = ~n911 & ~n916;
  assign n918 = ~sys_fair0done_out & ~n917;
  assign n919 = ~n913 & ~n918;
  assign n920 = ~reg_controllable_BtoS_ACK0_out & ~n919;
  assign n921 = ~reg_controllable_BtoS_ACK0_out & ~n920;
  assign n922 = reg_i_StoB_REQ0_out & ~n921;
  assign n923 = ~n387 & ~n913;
  assign n924 = reg_controllable_BtoS_ACK0_out & ~n923;
  assign n925 = ~n920 & ~n924;
  assign n926 = ~reg_i_StoB_REQ0_out & ~n925;
  assign n927 = ~n922 & ~n926;
  assign n928 = ~reg_controllable_BtoS_ACK10_out & ~n927;
  assign n929 = ~reg_controllable_BtoS_ACK10_out & ~n928;
  assign n930 = reg_i_StoB_REQ10_out & ~n929;
  assign n931 = ~reg_i_StoB_REQ2_out & ~n445;
  assign n932 = ~sys_fair2done_out & ~n931;
  assign n933 = ~n442 & ~n932;
  assign n934 = sys_fair1done_out & ~n933;
  assign n935 = reg_i_StoB_REQ2_out & ~n719;
  assign n936 = sys_fair2done_out & ~n935;
  assign n937 = ~n445 & ~n719;
  assign n938 = ~sys_fair2done_out & ~n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~sys_fair1done_out & ~n939;
  assign n941 = ~n934 & ~n940;
  assign n942 = ~reg_i_StoB_REQ3_out & ~n941;
  assign n943 = ~n732 & ~n942;
  assign n944 = sys_fair3done_out & ~n943;
  assign n945 = ~sys_fair2done_out & ~n932;
  assign n946 = sys_fair1done_out & ~n945;
  assign n947 = ~n940 & ~n946;
  assign n948 = ~reg_controllable_BtoS_ACK3_out & ~n947;
  assign n949 = ~n459 & ~n948;
  assign n950 = ~reg_i_StoB_REQ3_out & ~n949;
  assign n951 = ~n741 & ~n950;
  assign n952 = ~sys_fair3done_out & ~n951;
  assign n953 = ~n944 & ~n952;
  assign n954 = ~reg_i_StoB_REQ4_out & ~n953;
  assign n955 = ~n749 & ~n954;
  assign n956 = sys_fair4done_out & ~n955;
  assign n957 = ~reg_i_StoB_REQ3_out & ~n947;
  assign n958 = ~n741 & ~n957;
  assign n959 = sys_fair3done_out & ~n958;
  assign n960 = ~n952 & ~n959;
  assign n961 = ~reg_controllable_BtoS_ACK4_out & ~n960;
  assign n962 = ~n474 & ~n961;
  assign n963 = ~reg_i_StoB_REQ4_out & ~n962;
  assign n964 = ~n759 & ~n963;
  assign n965 = ~sys_fair4done_out & ~n964;
  assign n966 = ~n956 & ~n965;
  assign n967 = ~reg_i_StoB_REQ5_out & ~n966;
  assign n968 = ~n767 & ~n967;
  assign n969 = sys_fair5done_out & ~n968;
  assign n970 = ~reg_i_StoB_REQ4_out & ~n960;
  assign n971 = ~n759 & ~n970;
  assign n972 = sys_fair4done_out & ~n971;
  assign n973 = ~n965 & ~n972;
  assign n974 = ~reg_controllable_BtoS_ACK5_out & ~n973;
  assign n975 = ~n490 & ~n974;
  assign n976 = ~reg_i_StoB_REQ5_out & ~n975;
  assign n977 = ~n777 & ~n976;
  assign n978 = ~sys_fair5done_out & ~n977;
  assign n979 = ~n969 & ~n978;
  assign n980 = ~reg_i_StoB_REQ8_out & ~n979;
  assign n981 = ~n785 & ~n980;
  assign n982 = sys_fair8done_out & ~n981;
  assign n983 = ~reg_i_StoB_REQ5_out & ~n973;
  assign n984 = ~n777 & ~n983;
  assign n985 = sys_fair5done_out & ~n984;
  assign n986 = ~n978 & ~n985;
  assign n987 = ~reg_controllable_BtoS_ACK8_out & ~n986;
  assign n988 = ~n506 & ~n987;
  assign n989 = ~reg_i_StoB_REQ8_out & ~n988;
  assign n990 = ~n795 & ~n989;
  assign n991 = ~sys_fair8done_out & ~n990;
  assign n992 = ~n982 & ~n991;
  assign n993 = ~reg_i_StoB_REQ6_out & ~n992;
  assign n994 = ~n803 & ~n993;
  assign n995 = sys_fair6done_out & ~n994;
  assign n996 = ~reg_i_StoB_REQ8_out & ~n986;
  assign n997 = ~n795 & ~n996;
  assign n998 = sys_fair8done_out & ~n997;
  assign n999 = ~n991 & ~n998;
  assign n1000 = ~reg_controllable_BtoS_ACK6_out & ~n999;
  assign n1001 = ~n522 & ~n1000;
  assign n1002 = ~reg_i_StoB_REQ6_out & ~n1001;
  assign n1003 = ~n813 & ~n1002;
  assign n1004 = ~sys_fair6done_out & ~n1003;
  assign n1005 = ~n995 & ~n1004;
  assign n1006 = sys_fair7done_out & ~n1005;
  assign n1007 = ~n536 & ~n1006;
  assign n1008 = reg_controllable_BtoS_ACK7_out & ~n1007;
  assign n1009 = ~reg_i_StoB_REQ6_out & ~n999;
  assign n1010 = ~n813 & ~n1009;
  assign n1011 = sys_fair6done_out & ~n1010;
  assign n1012 = ~n1004 & ~n1011;
  assign n1013 = ~sys_fair7done_out & ~n1012;
  assign n1014 = ~n1006 & ~n1013;
  assign n1015 = ~reg_controllable_BtoS_ACK7_out & ~n1014;
  assign n1016 = ~n1008 & ~n1015;
  assign n1017 = ~reg_i_StoB_REQ7_out & ~n1016;
  assign n1018 = ~n828 & ~n1017;
  assign n1019 = ~reg_i_StoB_REQ9_out & ~n1018;
  assign n1020 = ~n836 & ~n1019;
  assign n1021 = sys_fair9done_out & ~n1020;
  assign n1022 = sys_fair7done_out & ~n1012;
  assign n1023 = ~n536 & ~n1022;
  assign n1024 = reg_controllable_BtoS_ACK7_out & ~n1023;
  assign n1025 = ~reg_controllable_BtoS_ACK7_out & ~n1012;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~reg_i_StoB_REQ7_out & ~n1026;
  assign n1028 = ~n842 & ~n1027;
  assign n1029 = ~reg_controllable_BtoS_ACK9_out & ~n1028;
  assign n1030 = ~n554 & ~n1029;
  assign n1031 = ~reg_i_StoB_REQ9_out & ~n1030;
  assign n1032 = ~n851 & ~n1031;
  assign n1033 = ~sys_fair9done_out & ~n1032;
  assign n1034 = ~n1021 & ~n1033;
  assign n1035 = ~reg_i_StoB_REQ11_out & ~n1034;
  assign n1036 = ~n859 & ~n1035;
  assign n1037 = sys_fair11done_out & ~n1036;
  assign n1038 = ~reg_i_StoB_REQ9_out & ~n1028;
  assign n1039 = ~n851 & ~n1038;
  assign n1040 = sys_fair9done_out & ~n1039;
  assign n1041 = ~n1033 & ~n1040;
  assign n1042 = ~reg_controllable_BtoS_ACK11_out & ~n1041;
  assign n1043 = ~n573 & ~n1042;
  assign n1044 = ~reg_i_StoB_REQ11_out & ~n1043;
  assign n1045 = ~n869 & ~n1044;
  assign n1046 = ~sys_fair11done_out & ~n1045;
  assign n1047 = ~n1037 & ~n1046;
  assign n1048 = sys_fair12done_out & ~n1047;
  assign n1049 = ~n587 & ~n1048;
  assign n1050 = reg_controllable_BtoS_ACK12_out & ~n1049;
  assign n1051 = ~reg_i_StoB_REQ11_out & ~n1041;
  assign n1052 = ~n869 & ~n1051;
  assign n1053 = sys_fair11done_out & ~n1052;
  assign n1054 = ~n1046 & ~n1053;
  assign n1055 = ~sys_fair12done_out & ~n1054;
  assign n1056 = ~n1048 & ~n1055;
  assign n1057 = ~reg_controllable_BtoS_ACK12_out & ~n1056;
  assign n1058 = ~n1050 & ~n1057;
  assign n1059 = ~reg_i_StoB_REQ12_out & ~n1058;
  assign n1060 = ~n884 & ~n1059;
  assign n1061 = ~reg_i_StoB_REQ13_out & ~n1060;
  assign n1062 = ~n892 & ~n1061;
  assign n1063 = sys_fair13done_out & ~n1062;
  assign n1064 = sys_fair12done_out & ~n1054;
  assign n1065 = ~n587 & ~n1064;
  assign n1066 = reg_controllable_BtoS_ACK12_out & ~n1065;
  assign n1067 = ~reg_controllable_BtoS_ACK12_out & ~n1054;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~reg_i_StoB_REQ12_out & ~n1068;
  assign n1070 = ~n898 & ~n1069;
  assign n1071 = ~reg_controllable_BtoS_ACK13_out & ~n1070;
  assign n1072 = ~n605 & ~n1071;
  assign n1073 = ~reg_i_StoB_REQ13_out & ~n1072;
  assign n1074 = ~n907 & ~n1073;
  assign n1075 = ~sys_fair13done_out & ~n1074;
  assign n1076 = ~n1063 & ~n1075;
  assign n1077 = sys_fair0done_out & ~n1076;
  assign n1078 = ~n622 & ~n1077;
  assign n1079 = reg_controllable_BtoS_ACK0_out & ~n1078;
  assign n1080 = ~reg_i_StoB_REQ13_out & ~n1070;
  assign n1081 = ~n907 & ~n1080;
  assign n1082 = sys_fair13done_out & ~n1081;
  assign n1083 = ~n1075 & ~n1082;
  assign n1084 = ~sys_fair0done_out & ~n1083;
  assign n1085 = ~n1077 & ~n1084;
  assign n1086 = ~reg_controllable_BtoS_ACK0_out & ~n1085;
  assign n1087 = ~n1079 & ~n1086;
  assign n1088 = ~reg_i_StoB_REQ0_out & ~n1087;
  assign n1089 = ~n922 & ~n1088;
  assign n1090 = ~reg_i_StoB_REQ10_out & ~n1089;
  assign n1091 = ~n930 & ~n1090;
  assign n1092 = sys_fair10done_out & ~n1091;
  assign n1093 = ~reg_controllable_BtoS_ACK0_out & ~n917;
  assign n1094 = ~reg_controllable_BtoS_ACK0_out & ~n1093;
  assign n1095 = reg_i_StoB_REQ0_out & ~n1094;
  assign n1096 = sys_fair0done_out & ~n917;
  assign n1097 = ~n387 & ~n1096;
  assign n1098 = reg_controllable_BtoS_ACK0_out & ~n1097;
  assign n1099 = ~n1093 & ~n1098;
  assign n1100 = ~reg_i_StoB_REQ0_out & ~n1099;
  assign n1101 = ~n1095 & ~n1100;
  assign n1102 = ~reg_controllable_BtoS_ACK10_out & ~n1101;
  assign n1103 = ~reg_controllable_BtoS_ACK10_out & ~n1102;
  assign n1104 = reg_i_StoB_REQ10_out & ~n1103;
  assign n1105 = sys_fair0done_out & ~n1083;
  assign n1106 = ~n622 & ~n1105;
  assign n1107 = reg_controllable_BtoS_ACK0_out & ~n1106;
  assign n1108 = ~reg_controllable_BtoS_ACK0_out & ~n1083;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~reg_i_StoB_REQ0_out & ~n1109;
  assign n1111 = ~n1095 & ~n1110;
  assign n1112 = ~reg_controllable_BtoS_ACK10_out & ~n1111;
  assign n1113 = ~n640 & ~n1112;
  assign n1114 = ~reg_i_StoB_REQ10_out & ~n1113;
  assign n1115 = ~n1104 & ~n1114;
  assign n1116 = ~sys_fair10done_out & ~n1115;
  assign n1117 = ~n1092 & ~n1116;
  assign n1118 = reg_controllable_BtoS_ACK14_out & ~n1117;
  assign n1119 = reg_controllable_BtoS_ACK10_out & ~n927;
  assign n1120 = reg_controllable_BtoS_ACK0_out & ~n919;
  assign n1121 = reg_controllable_BtoS_ACK13_out & ~n889;
  assign n1122 = reg_controllable_BtoS_ACK12_out & ~n881;
  assign n1123 = reg_controllable_BtoS_ACK11_out & ~n856;
  assign n1124 = reg_controllable_BtoS_ACK9_out & ~n833;
  assign n1125 = reg_controllable_BtoS_ACK7_out & ~n825;
  assign n1126 = reg_controllable_BtoS_ACK6_out & ~n800;
  assign n1127 = reg_controllable_BtoS_ACK8_out & ~n782;
  assign n1128 = reg_controllable_BtoS_ACK5_out & ~n764;
  assign n1129 = reg_controllable_BtoS_ACK4_out & ~n746;
  assign n1130 = reg_controllable_BtoS_ACK3_out & ~n729;
  assign n1131 = reg_i_StoB_REQ2_out & n119;
  assign n1132 = sys_fair2done_out & n1131;
  assign n1133 = ~reg_i_StoB_REQ2_out & ~reg_controllable_BtoS_ACK2_out;
  assign n1134 = ~n115 & ~n1133;
  assign n1135 = ~sys_fair2done_out & ~n1134;
  assign n1136 = ~n1132 & ~n1135;
  assign n1137 = sys_fair1done_out & ~n1136;
  assign n1138 = reg_controllable_BtoS_ACK2_out & ~n716;
  assign n1139 = ~n128 & ~n1138;
  assign n1140 = reg_i_StoB_REQ2_out & ~n1139;
  assign n1141 = ~n131 & ~n1140;
  assign n1142 = sys_fair2done_out & ~n1141;
  assign n1143 = ~n113 & ~n1138;
  assign n1144 = reg_i_StoB_REQ2_out & ~n1143;
  assign n1145 = ~reg_controllable_BtoS_ACK2_out & n127;
  assign n1146 = ~reg_controllable_BtoS_ACK2_out & ~n1145;
  assign n1147 = ~reg_i_StoB_REQ2_out & n1146;
  assign n1148 = ~n1144 & ~n1147;
  assign n1149 = ~sys_fair2done_out & ~n1148;
  assign n1150 = ~n1142 & ~n1149;
  assign n1151 = ~sys_fair1done_out & ~n1150;
  assign n1152 = ~n1137 & ~n1151;
  assign n1153 = ~reg_controllable_BtoS_ACK3_out & ~n1152;
  assign n1154 = ~n1130 & ~n1153;
  assign n1155 = reg_i_StoB_REQ3_out & ~n1154;
  assign n1156 = ~reg_i_StoB_REQ3_out & ~n1152;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = sys_fair3done_out & ~n1157;
  assign n1159 = reg_controllable_BtoS_ACK3_out & ~n738;
  assign n1160 = ~reg_controllable_BtoS_ACK2_out & ~n112;
  assign n1161 = ~reg_controllable_BtoS_ACK2_out & ~n1160;
  assign n1162 = ~reg_i_StoB_REQ2_out & n1161;
  assign n1163 = ~n115 & ~n1162;
  assign n1164 = ~sys_fair2done_out & ~n1163;
  assign n1165 = ~n118 & ~n1164;
  assign n1166 = sys_fair1done_out & ~n1165;
  assign n1167 = ~n116 & ~n1144;
  assign n1168 = sys_fair2done_out & ~n1167;
  assign n1169 = ~n1144 & ~n1162;
  assign n1170 = ~sys_fair2done_out & ~n1169;
  assign n1171 = ~n1168 & ~n1170;
  assign n1172 = ~sys_fair1done_out & ~n1171;
  assign n1173 = ~n1166 & ~n1172;
  assign n1174 = ~reg_controllable_BtoS_ACK3_out & ~n1173;
  assign n1175 = ~n1159 & ~n1174;
  assign n1176 = reg_i_StoB_REQ3_out & ~n1175;
  assign n1177 = reg_controllable_BtoS_ACK3_out & n1131;
  assign n1178 = ~sys_fair2done_out & ~n1135;
  assign n1179 = sys_fair1done_out & ~n1178;
  assign n1180 = ~n1151 & ~n1179;
  assign n1181 = ~reg_controllable_BtoS_ACK3_out & ~n1180;
  assign n1182 = ~n1177 & ~n1181;
  assign n1183 = ~reg_i_StoB_REQ3_out & ~n1182;
  assign n1184 = ~n1176 & ~n1183;
  assign n1185 = ~sys_fair3done_out & ~n1184;
  assign n1186 = ~n1158 & ~n1185;
  assign n1187 = ~reg_controllable_BtoS_ACK4_out & ~n1186;
  assign n1188 = ~n1129 & ~n1187;
  assign n1189 = reg_i_StoB_REQ4_out & ~n1188;
  assign n1190 = ~reg_i_StoB_REQ4_out & ~n1186;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = sys_fair4done_out & ~n1191;
  assign n1193 = reg_controllable_BtoS_ACK4_out & ~n756;
  assign n1194 = ~reg_i_StoB_REQ3_out & ~n1173;
  assign n1195 = ~n1176 & ~n1194;
  assign n1196 = sys_fair3done_out & ~n1195;
  assign n1197 = ~n1174 & ~n1177;
  assign n1198 = ~reg_i_StoB_REQ3_out & ~n1197;
  assign n1199 = ~n1176 & ~n1198;
  assign n1200 = ~sys_fair3done_out & ~n1199;
  assign n1201 = ~n1196 & ~n1200;
  assign n1202 = ~reg_controllable_BtoS_ACK4_out & ~n1201;
  assign n1203 = ~n1193 & ~n1202;
  assign n1204 = reg_i_StoB_REQ4_out & ~n1203;
  assign n1205 = ~reg_controllable_BtoS_ACK3_out & n1131;
  assign n1206 = ~n150 & ~n1205;
  assign n1207 = reg_i_StoB_REQ3_out & ~n1206;
  assign n1208 = ~reg_i_StoB_REQ3_out & n1131;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = reg_controllable_BtoS_ACK4_out & ~n1209;
  assign n1211 = ~n1159 & ~n1181;
  assign n1212 = reg_i_StoB_REQ3_out & ~n1211;
  assign n1213 = ~reg_i_StoB_REQ3_out & ~n1180;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = sys_fair3done_out & ~n1214;
  assign n1216 = ~n1185 & ~n1215;
  assign n1217 = ~reg_controllable_BtoS_ACK4_out & ~n1216;
  assign n1218 = ~n1210 & ~n1217;
  assign n1219 = ~reg_i_StoB_REQ4_out & ~n1218;
  assign n1220 = ~n1204 & ~n1219;
  assign n1221 = ~sys_fair4done_out & ~n1220;
  assign n1222 = ~n1192 & ~n1221;
  assign n1223 = ~reg_controllable_BtoS_ACK5_out & ~n1222;
  assign n1224 = ~n1128 & ~n1223;
  assign n1225 = reg_i_StoB_REQ5_out & ~n1224;
  assign n1226 = ~reg_i_StoB_REQ5_out & ~n1222;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = sys_fair5done_out & ~n1227;
  assign n1229 = reg_controllable_BtoS_ACK5_out & ~n774;
  assign n1230 = ~reg_i_StoB_REQ4_out & ~n1201;
  assign n1231 = ~n1204 & ~n1230;
  assign n1232 = sys_fair4done_out & ~n1231;
  assign n1233 = ~n1202 & ~n1210;
  assign n1234 = ~reg_i_StoB_REQ4_out & ~n1233;
  assign n1235 = ~n1204 & ~n1234;
  assign n1236 = ~sys_fair4done_out & ~n1235;
  assign n1237 = ~n1232 & ~n1236;
  assign n1238 = ~reg_controllable_BtoS_ACK5_out & ~n1237;
  assign n1239 = ~n1229 & ~n1238;
  assign n1240 = reg_i_StoB_REQ5_out & ~n1239;
  assign n1241 = ~reg_controllable_BtoS_ACK4_out & ~n1209;
  assign n1242 = ~n171 & ~n1241;
  assign n1243 = reg_i_StoB_REQ4_out & ~n1242;
  assign n1244 = ~reg_i_StoB_REQ4_out & ~n1209;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = reg_controllable_BtoS_ACK5_out & ~n1245;
  assign n1247 = ~n1193 & ~n1217;
  assign n1248 = reg_i_StoB_REQ4_out & ~n1247;
  assign n1249 = ~reg_i_StoB_REQ4_out & ~n1216;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = sys_fair4done_out & ~n1250;
  assign n1252 = ~n1221 & ~n1251;
  assign n1253 = ~reg_controllable_BtoS_ACK5_out & ~n1252;
  assign n1254 = ~n1246 & ~n1253;
  assign n1255 = ~reg_i_StoB_REQ5_out & ~n1254;
  assign n1256 = ~n1240 & ~n1255;
  assign n1257 = ~sys_fair5done_out & ~n1256;
  assign n1258 = ~n1228 & ~n1257;
  assign n1259 = ~reg_controllable_BtoS_ACK8_out & ~n1258;
  assign n1260 = ~n1127 & ~n1259;
  assign n1261 = reg_i_StoB_REQ8_out & ~n1260;
  assign n1262 = ~reg_i_StoB_REQ8_out & ~n1258;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = sys_fair8done_out & ~n1263;
  assign n1265 = reg_controllable_BtoS_ACK8_out & ~n792;
  assign n1266 = ~reg_i_StoB_REQ5_out & ~n1237;
  assign n1267 = ~n1240 & ~n1266;
  assign n1268 = sys_fair5done_out & ~n1267;
  assign n1269 = ~n1238 & ~n1246;
  assign n1270 = ~reg_i_StoB_REQ5_out & ~n1269;
  assign n1271 = ~n1240 & ~n1270;
  assign n1272 = ~sys_fair5done_out & ~n1271;
  assign n1273 = ~n1268 & ~n1272;
  assign n1274 = ~reg_controllable_BtoS_ACK8_out & ~n1273;
  assign n1275 = ~n1265 & ~n1274;
  assign n1276 = reg_i_StoB_REQ8_out & ~n1275;
  assign n1277 = ~reg_controllable_BtoS_ACK5_out & ~n1245;
  assign n1278 = ~n195 & ~n1277;
  assign n1279 = reg_i_StoB_REQ5_out & ~n1278;
  assign n1280 = ~reg_i_StoB_REQ5_out & ~n1245;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = reg_controllable_BtoS_ACK8_out & ~n1281;
  assign n1283 = ~n1229 & ~n1253;
  assign n1284 = reg_i_StoB_REQ5_out & ~n1283;
  assign n1285 = ~reg_i_StoB_REQ5_out & ~n1252;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = sys_fair5done_out & ~n1286;
  assign n1288 = ~n1257 & ~n1287;
  assign n1289 = ~reg_controllable_BtoS_ACK8_out & ~n1288;
  assign n1290 = ~n1282 & ~n1289;
  assign n1291 = ~reg_i_StoB_REQ8_out & ~n1290;
  assign n1292 = ~n1276 & ~n1291;
  assign n1293 = ~sys_fair8done_out & ~n1292;
  assign n1294 = ~n1264 & ~n1293;
  assign n1295 = ~reg_controllable_BtoS_ACK6_out & ~n1294;
  assign n1296 = ~n1126 & ~n1295;
  assign n1297 = reg_i_StoB_REQ6_out & ~n1296;
  assign n1298 = ~reg_i_StoB_REQ6_out & ~n1294;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = sys_fair6done_out & ~n1299;
  assign n1301 = reg_controllable_BtoS_ACK6_out & ~n810;
  assign n1302 = ~reg_i_StoB_REQ8_out & ~n1273;
  assign n1303 = ~n1276 & ~n1302;
  assign n1304 = sys_fair8done_out & ~n1303;
  assign n1305 = ~n1274 & ~n1282;
  assign n1306 = ~reg_i_StoB_REQ8_out & ~n1305;
  assign n1307 = ~n1276 & ~n1306;
  assign n1308 = ~sys_fair8done_out & ~n1307;
  assign n1309 = ~n1304 & ~n1308;
  assign n1310 = ~reg_controllable_BtoS_ACK6_out & ~n1309;
  assign n1311 = ~n1301 & ~n1310;
  assign n1312 = reg_i_StoB_REQ6_out & ~n1311;
  assign n1313 = ~reg_controllable_BtoS_ACK8_out & ~n1281;
  assign n1314 = ~n219 & ~n1313;
  assign n1315 = reg_i_StoB_REQ8_out & ~n1314;
  assign n1316 = ~reg_i_StoB_REQ8_out & ~n1281;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = reg_controllable_BtoS_ACK6_out & ~n1317;
  assign n1319 = ~n1265 & ~n1289;
  assign n1320 = reg_i_StoB_REQ8_out & ~n1319;
  assign n1321 = ~reg_i_StoB_REQ8_out & ~n1288;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = sys_fair8done_out & ~n1322;
  assign n1324 = ~n1293 & ~n1323;
  assign n1325 = ~reg_controllable_BtoS_ACK6_out & ~n1324;
  assign n1326 = ~n1318 & ~n1325;
  assign n1327 = ~reg_i_StoB_REQ6_out & ~n1326;
  assign n1328 = ~n1312 & ~n1327;
  assign n1329 = ~sys_fair6done_out & ~n1328;
  assign n1330 = ~n1300 & ~n1329;
  assign n1331 = sys_fair7done_out & ~n1330;
  assign n1332 = ~reg_i_StoB_REQ6_out & ~n1309;
  assign n1333 = ~n1312 & ~n1332;
  assign n1334 = sys_fair6done_out & ~n1333;
  assign n1335 = ~n1310 & ~n1318;
  assign n1336 = ~reg_i_StoB_REQ6_out & ~n1335;
  assign n1337 = ~n1312 & ~n1336;
  assign n1338 = ~sys_fair6done_out & ~n1337;
  assign n1339 = ~n1334 & ~n1338;
  assign n1340 = ~sys_fair7done_out & ~n1339;
  assign n1341 = ~n1331 & ~n1340;
  assign n1342 = ~reg_controllable_BtoS_ACK7_out & ~n1341;
  assign n1343 = ~n1125 & ~n1342;
  assign n1344 = reg_i_StoB_REQ7_out & ~n1343;
  assign n1345 = ~reg_controllable_BtoS_ACK6_out & ~n1317;
  assign n1346 = ~n243 & ~n1345;
  assign n1347 = reg_i_StoB_REQ6_out & ~n1346;
  assign n1348 = ~reg_i_StoB_REQ6_out & ~n1317;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~sys_fair7done_out & ~n1349;
  assign n1351 = ~n1331 & ~n1350;
  assign n1352 = reg_controllable_BtoS_ACK7_out & ~n1351;
  assign n1353 = ~n1301 & ~n1325;
  assign n1354 = reg_i_StoB_REQ6_out & ~n1353;
  assign n1355 = ~reg_i_StoB_REQ6_out & ~n1324;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = sys_fair6done_out & ~n1356;
  assign n1358 = ~n1329 & ~n1357;
  assign n1359 = ~sys_fair7done_out & ~n1358;
  assign n1360 = ~n1331 & ~n1359;
  assign n1361 = ~reg_controllable_BtoS_ACK7_out & ~n1360;
  assign n1362 = ~n1352 & ~n1361;
  assign n1363 = ~reg_i_StoB_REQ7_out & ~n1362;
  assign n1364 = ~n1344 & ~n1363;
  assign n1365 = ~reg_controllable_BtoS_ACK9_out & ~n1364;
  assign n1366 = ~n1124 & ~n1365;
  assign n1367 = reg_i_StoB_REQ9_out & ~n1366;
  assign n1368 = ~reg_i_StoB_REQ9_out & ~n1364;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = sys_fair9done_out & ~n1369;
  assign n1371 = reg_controllable_BtoS_ACK9_out & ~n848;
  assign n1372 = reg_controllable_BtoS_ACK7_out & ~n823;
  assign n1373 = ~reg_controllable_BtoS_ACK7_out & ~n1339;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = reg_i_StoB_REQ7_out & ~n1374;
  assign n1376 = sys_fair7done_out & ~n1339;
  assign n1377 = ~n1350 & ~n1376;
  assign n1378 = reg_controllable_BtoS_ACK7_out & ~n1377;
  assign n1379 = ~n1373 & ~n1378;
  assign n1380 = ~reg_i_StoB_REQ7_out & ~n1379;
  assign n1381 = ~n1375 & ~n1380;
  assign n1382 = ~reg_controllable_BtoS_ACK9_out & ~n1381;
  assign n1383 = ~n1371 & ~n1382;
  assign n1384 = reg_i_StoB_REQ9_out & ~n1383;
  assign n1385 = reg_controllable_BtoS_ACK7_out & ~n258;
  assign n1386 = ~reg_controllable_BtoS_ACK7_out & ~n1349;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = reg_i_StoB_REQ7_out & ~n1387;
  assign n1389 = ~reg_i_StoB_REQ7_out & ~n1349;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = reg_controllable_BtoS_ACK9_out & ~n1390;
  assign n1392 = sys_fair7done_out & ~n1358;
  assign n1393 = ~n1340 & ~n1392;
  assign n1394 = ~reg_controllable_BtoS_ACK7_out & ~n1393;
  assign n1395 = ~n1372 & ~n1394;
  assign n1396 = reg_i_StoB_REQ7_out & ~n1395;
  assign n1397 = ~n1350 & ~n1392;
  assign n1398 = reg_controllable_BtoS_ACK7_out & ~n1397;
  assign n1399 = ~reg_controllable_BtoS_ACK7_out & ~n1358;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = ~reg_i_StoB_REQ7_out & ~n1400;
  assign n1402 = ~n1396 & ~n1401;
  assign n1403 = ~reg_controllable_BtoS_ACK9_out & ~n1402;
  assign n1404 = ~n1391 & ~n1403;
  assign n1405 = ~reg_i_StoB_REQ9_out & ~n1404;
  assign n1406 = ~n1384 & ~n1405;
  assign n1407 = ~sys_fair9done_out & ~n1406;
  assign n1408 = ~n1370 & ~n1407;
  assign n1409 = ~reg_controllable_BtoS_ACK11_out & ~n1408;
  assign n1410 = ~n1123 & ~n1409;
  assign n1411 = reg_i_StoB_REQ11_out & ~n1410;
  assign n1412 = ~reg_i_StoB_REQ11_out & ~n1408;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = sys_fair11done_out & ~n1413;
  assign n1415 = reg_controllable_BtoS_ACK11_out & ~n866;
  assign n1416 = ~reg_i_StoB_REQ9_out & ~n1381;
  assign n1417 = ~n1384 & ~n1416;
  assign n1418 = sys_fair9done_out & ~n1417;
  assign n1419 = ~n1382 & ~n1391;
  assign n1420 = ~reg_i_StoB_REQ9_out & ~n1419;
  assign n1421 = ~n1384 & ~n1420;
  assign n1422 = ~sys_fair9done_out & ~n1421;
  assign n1423 = ~n1418 & ~n1422;
  assign n1424 = ~reg_controllable_BtoS_ACK11_out & ~n1423;
  assign n1425 = ~n1415 & ~n1424;
  assign n1426 = reg_i_StoB_REQ11_out & ~n1425;
  assign n1427 = ~reg_controllable_BtoS_ACK9_out & ~n1390;
  assign n1428 = ~n291 & ~n1427;
  assign n1429 = reg_i_StoB_REQ9_out & ~n1428;
  assign n1430 = ~reg_i_StoB_REQ9_out & ~n1390;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = reg_controllable_BtoS_ACK11_out & ~n1431;
  assign n1433 = ~n1371 & ~n1403;
  assign n1434 = reg_i_StoB_REQ9_out & ~n1433;
  assign n1435 = ~reg_i_StoB_REQ9_out & ~n1402;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = sys_fair9done_out & ~n1436;
  assign n1438 = ~n1407 & ~n1437;
  assign n1439 = ~reg_controllable_BtoS_ACK11_out & ~n1438;
  assign n1440 = ~n1432 & ~n1439;
  assign n1441 = ~reg_i_StoB_REQ11_out & ~n1440;
  assign n1442 = ~n1426 & ~n1441;
  assign n1443 = ~sys_fair11done_out & ~n1442;
  assign n1444 = ~n1414 & ~n1443;
  assign n1445 = sys_fair12done_out & ~n1444;
  assign n1446 = ~reg_i_StoB_REQ11_out & ~n1423;
  assign n1447 = ~n1426 & ~n1446;
  assign n1448 = sys_fair11done_out & ~n1447;
  assign n1449 = ~n1424 & ~n1432;
  assign n1450 = ~reg_i_StoB_REQ11_out & ~n1449;
  assign n1451 = ~n1426 & ~n1450;
  assign n1452 = ~sys_fair11done_out & ~n1451;
  assign n1453 = ~n1448 & ~n1452;
  assign n1454 = ~sys_fair12done_out & ~n1453;
  assign n1455 = ~n1445 & ~n1454;
  assign n1456 = ~reg_controllable_BtoS_ACK12_out & ~n1455;
  assign n1457 = ~n1122 & ~n1456;
  assign n1458 = reg_i_StoB_REQ12_out & ~n1457;
  assign n1459 = ~reg_controllable_BtoS_ACK11_out & ~n1431;
  assign n1460 = ~n319 & ~n1459;
  assign n1461 = reg_i_StoB_REQ11_out & ~n1460;
  assign n1462 = ~reg_i_StoB_REQ11_out & ~n1431;
  assign n1463 = ~n1461 & ~n1462;
  assign n1464 = ~sys_fair12done_out & ~n1463;
  assign n1465 = ~n1445 & ~n1464;
  assign n1466 = reg_controllable_BtoS_ACK12_out & ~n1465;
  assign n1467 = ~n1415 & ~n1439;
  assign n1468 = reg_i_StoB_REQ11_out & ~n1467;
  assign n1469 = ~reg_i_StoB_REQ11_out & ~n1438;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = sys_fair11done_out & ~n1470;
  assign n1472 = ~n1443 & ~n1471;
  assign n1473 = ~sys_fair12done_out & ~n1472;
  assign n1474 = ~n1445 & ~n1473;
  assign n1475 = ~reg_controllable_BtoS_ACK12_out & ~n1474;
  assign n1476 = ~n1466 & ~n1475;
  assign n1477 = ~reg_i_StoB_REQ12_out & ~n1476;
  assign n1478 = ~n1458 & ~n1477;
  assign n1479 = ~reg_controllable_BtoS_ACK13_out & ~n1478;
  assign n1480 = ~n1121 & ~n1479;
  assign n1481 = reg_i_StoB_REQ13_out & ~n1480;
  assign n1482 = ~reg_i_StoB_REQ13_out & ~n1478;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = sys_fair13done_out & ~n1483;
  assign n1485 = reg_controllable_BtoS_ACK13_out & ~n904;
  assign n1486 = reg_controllable_BtoS_ACK12_out & ~n879;
  assign n1487 = ~reg_controllable_BtoS_ACK12_out & ~n1453;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = reg_i_StoB_REQ12_out & ~n1488;
  assign n1490 = sys_fair12done_out & ~n1453;
  assign n1491 = ~n1464 & ~n1490;
  assign n1492 = reg_controllable_BtoS_ACK12_out & ~n1491;
  assign n1493 = ~n1487 & ~n1492;
  assign n1494 = ~reg_i_StoB_REQ12_out & ~n1493;
  assign n1495 = ~n1489 & ~n1494;
  assign n1496 = ~reg_controllable_BtoS_ACK13_out & ~n1495;
  assign n1497 = ~n1485 & ~n1496;
  assign n1498 = reg_i_StoB_REQ13_out & ~n1497;
  assign n1499 = reg_controllable_BtoS_ACK12_out & ~n334;
  assign n1500 = ~reg_controllable_BtoS_ACK12_out & ~n1463;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = reg_i_StoB_REQ12_out & ~n1501;
  assign n1503 = ~reg_i_StoB_REQ12_out & ~n1463;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = reg_controllable_BtoS_ACK13_out & ~n1504;
  assign n1506 = sys_fair12done_out & ~n1472;
  assign n1507 = ~n1454 & ~n1506;
  assign n1508 = ~reg_controllable_BtoS_ACK12_out & ~n1507;
  assign n1509 = ~n1486 & ~n1508;
  assign n1510 = reg_i_StoB_REQ12_out & ~n1509;
  assign n1511 = ~n1464 & ~n1506;
  assign n1512 = reg_controllable_BtoS_ACK12_out & ~n1511;
  assign n1513 = ~reg_controllable_BtoS_ACK12_out & ~n1472;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~reg_i_StoB_REQ12_out & ~n1514;
  assign n1516 = ~n1510 & ~n1515;
  assign n1517 = ~reg_controllable_BtoS_ACK13_out & ~n1516;
  assign n1518 = ~n1505 & ~n1517;
  assign n1519 = ~reg_i_StoB_REQ13_out & ~n1518;
  assign n1520 = ~n1498 & ~n1519;
  assign n1521 = ~sys_fair13done_out & ~n1520;
  assign n1522 = ~n1484 & ~n1521;
  assign n1523 = sys_fair0done_out & ~n1522;
  assign n1524 = ~reg_i_StoB_REQ13_out & ~n1495;
  assign n1525 = ~n1498 & ~n1524;
  assign n1526 = sys_fair13done_out & ~n1525;
  assign n1527 = ~n1496 & ~n1505;
  assign n1528 = ~reg_i_StoB_REQ13_out & ~n1527;
  assign n1529 = ~n1498 & ~n1528;
  assign n1530 = ~sys_fair13done_out & ~n1529;
  assign n1531 = ~n1526 & ~n1530;
  assign n1532 = ~sys_fair0done_out & ~n1531;
  assign n1533 = ~n1523 & ~n1532;
  assign n1534 = ~reg_controllable_BtoS_ACK0_out & ~n1533;
  assign n1535 = ~n1120 & ~n1534;
  assign n1536 = reg_i_StoB_REQ0_out & ~n1535;
  assign n1537 = ~reg_controllable_BtoS_ACK13_out & ~n1504;
  assign n1538 = ~n367 & ~n1537;
  assign n1539 = reg_i_StoB_REQ13_out & ~n1538;
  assign n1540 = ~reg_i_StoB_REQ13_out & ~n1504;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~sys_fair0done_out & ~n1541;
  assign n1543 = ~n1523 & ~n1542;
  assign n1544 = reg_controllable_BtoS_ACK0_out & ~n1543;
  assign n1545 = ~n1485 & ~n1517;
  assign n1546 = reg_i_StoB_REQ13_out & ~n1545;
  assign n1547 = ~reg_i_StoB_REQ13_out & ~n1516;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = sys_fair13done_out & ~n1548;
  assign n1550 = ~n1521 & ~n1549;
  assign n1551 = ~sys_fair0done_out & ~n1550;
  assign n1552 = ~n1523 & ~n1551;
  assign n1553 = ~reg_controllable_BtoS_ACK0_out & ~n1552;
  assign n1554 = ~n1544 & ~n1553;
  assign n1555 = ~reg_i_StoB_REQ0_out & ~n1554;
  assign n1556 = ~n1536 & ~n1555;
  assign n1557 = ~reg_controllable_BtoS_ACK10_out & ~n1556;
  assign n1558 = ~n1119 & ~n1557;
  assign n1559 = reg_i_StoB_REQ10_out & ~n1558;
  assign n1560 = ~reg_i_StoB_REQ10_out & ~n1556;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = sys_fair10done_out & ~n1561;
  assign n1563 = reg_controllable_BtoS_ACK10_out & ~n1101;
  assign n1564 = reg_controllable_BtoS_ACK0_out & ~n917;
  assign n1565 = ~reg_controllable_BtoS_ACK0_out & ~n1531;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = reg_i_StoB_REQ0_out & ~n1566;
  assign n1568 = sys_fair0done_out & ~n1531;
  assign n1569 = ~n1542 & ~n1568;
  assign n1570 = reg_controllable_BtoS_ACK0_out & ~n1569;
  assign n1571 = ~n1565 & ~n1570;
  assign n1572 = ~reg_i_StoB_REQ0_out & ~n1571;
  assign n1573 = ~n1567 & ~n1572;
  assign n1574 = ~reg_controllable_BtoS_ACK10_out & ~n1573;
  assign n1575 = ~n1563 & ~n1574;
  assign n1576 = reg_i_StoB_REQ10_out & ~n1575;
  assign n1577 = reg_controllable_BtoS_ACK0_out & ~n386;
  assign n1578 = ~reg_controllable_BtoS_ACK0_out & ~n1541;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = reg_i_StoB_REQ0_out & ~n1579;
  assign n1581 = ~reg_i_StoB_REQ0_out & ~n1541;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = reg_controllable_BtoS_ACK10_out & ~n1582;
  assign n1584 = sys_fair0done_out & ~n1550;
  assign n1585 = ~n1532 & ~n1584;
  assign n1586 = ~reg_controllable_BtoS_ACK0_out & ~n1585;
  assign n1587 = ~n1564 & ~n1586;
  assign n1588 = reg_i_StoB_REQ0_out & ~n1587;
  assign n1589 = ~n1542 & ~n1584;
  assign n1590 = reg_controllable_BtoS_ACK0_out & ~n1589;
  assign n1591 = ~reg_controllable_BtoS_ACK0_out & ~n1550;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~reg_i_StoB_REQ0_out & ~n1592;
  assign n1594 = ~n1588 & ~n1593;
  assign n1595 = ~reg_controllable_BtoS_ACK10_out & ~n1594;
  assign n1596 = ~n1583 & ~n1595;
  assign n1597 = ~reg_i_StoB_REQ10_out & ~n1596;
  assign n1598 = ~n1576 & ~n1597;
  assign n1599 = ~sys_fair10done_out & ~n1598;
  assign n1600 = ~n1562 & ~n1599;
  assign n1601 = ~reg_controllable_BtoS_ACK14_out & ~n1600;
  assign n1602 = ~n1118 & ~n1601;
  assign n1603 = reg_i_StoB_REQ14_out & ~n1602;
  assign n1604 = reg_controllable_BtoS_ACK10_out & ~n1089;
  assign n1605 = ~n1557 & ~n1604;
  assign n1606 = reg_i_StoB_REQ10_out & ~n1605;
  assign n1607 = reg_controllable_BtoS_ACK0_out & ~n1085;
  assign n1608 = ~n1534 & ~n1607;
  assign n1609 = reg_i_StoB_REQ0_out & ~n1608;
  assign n1610 = reg_controllable_BtoS_ACK13_out & ~n1060;
  assign n1611 = ~n1479 & ~n1610;
  assign n1612 = reg_i_StoB_REQ13_out & ~n1611;
  assign n1613 = reg_controllable_BtoS_ACK12_out & ~n1056;
  assign n1614 = ~n1456 & ~n1613;
  assign n1615 = reg_i_StoB_REQ12_out & ~n1614;
  assign n1616 = reg_controllable_BtoS_ACK11_out & ~n1034;
  assign n1617 = ~n1409 & ~n1616;
  assign n1618 = reg_i_StoB_REQ11_out & ~n1617;
  assign n1619 = reg_controllable_BtoS_ACK9_out & ~n1018;
  assign n1620 = ~n1365 & ~n1619;
  assign n1621 = reg_i_StoB_REQ9_out & ~n1620;
  assign n1622 = reg_controllable_BtoS_ACK7_out & ~n1014;
  assign n1623 = ~n1342 & ~n1622;
  assign n1624 = reg_i_StoB_REQ7_out & ~n1623;
  assign n1625 = reg_controllable_BtoS_ACK6_out & ~n992;
  assign n1626 = ~n1295 & ~n1625;
  assign n1627 = reg_i_StoB_REQ6_out & ~n1626;
  assign n1628 = reg_controllable_BtoS_ACK8_out & ~n979;
  assign n1629 = ~n1259 & ~n1628;
  assign n1630 = reg_i_StoB_REQ8_out & ~n1629;
  assign n1631 = reg_controllable_BtoS_ACK5_out & ~n966;
  assign n1632 = ~n1223 & ~n1631;
  assign n1633 = reg_i_StoB_REQ5_out & ~n1632;
  assign n1634 = reg_controllable_BtoS_ACK4_out & ~n953;
  assign n1635 = ~n1187 & ~n1634;
  assign n1636 = reg_i_StoB_REQ4_out & ~n1635;
  assign n1637 = reg_controllable_BtoS_ACK3_out & ~n941;
  assign n1638 = ~n1153 & ~n1637;
  assign n1639 = reg_i_StoB_REQ3_out & ~n1638;
  assign n1640 = reg_i_StoB_REQ2_out & n443;
  assign n1641 = ~n440 & ~n1640;
  assign n1642 = sys_fair2done_out & ~n1641;
  assign n1643 = ~n447 & ~n1642;
  assign n1644 = sys_fair1done_out & ~n1643;
  assign n1645 = ~n454 & ~n1644;
  assign n1646 = ~reg_i_StoB_REQ3_out & ~n1645;
  assign n1647 = ~n1639 & ~n1646;
  assign n1648 = sys_fair3done_out & ~n1647;
  assign n1649 = reg_controllable_BtoS_ACK3_out & ~n947;
  assign n1650 = ~n1174 & ~n1649;
  assign n1651 = reg_i_StoB_REQ3_out & ~n1650;
  assign n1652 = reg_controllable_BtoS_ACK3_out & ~n1641;
  assign n1653 = ~n463 & ~n1652;
  assign n1654 = ~reg_i_StoB_REQ3_out & ~n1653;
  assign n1655 = ~n1651 & ~n1654;
  assign n1656 = ~sys_fair3done_out & ~n1655;
  assign n1657 = ~n1648 & ~n1656;
  assign n1658 = ~reg_i_StoB_REQ4_out & ~n1657;
  assign n1659 = ~n1636 & ~n1658;
  assign n1660 = sys_fair4done_out & ~n1659;
  assign n1661 = reg_controllable_BtoS_ACK4_out & ~n960;
  assign n1662 = ~n1202 & ~n1661;
  assign n1663 = reg_i_StoB_REQ4_out & ~n1662;
  assign n1664 = ~n459 & ~n1205;
  assign n1665 = reg_i_StoB_REQ3_out & ~n1664;
  assign n1666 = ~reg_i_StoB_REQ3_out & ~n1641;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = reg_controllable_BtoS_ACK4_out & ~n1667;
  assign n1669 = ~n1181 & ~n1649;
  assign n1670 = reg_i_StoB_REQ3_out & ~n1669;
  assign n1671 = ~n475 & ~n1670;
  assign n1672 = sys_fair3done_out & ~n1671;
  assign n1673 = ~n1656 & ~n1672;
  assign n1674 = ~reg_controllable_BtoS_ACK4_out & ~n1673;
  assign n1675 = ~n1668 & ~n1674;
  assign n1676 = ~reg_i_StoB_REQ4_out & ~n1675;
  assign n1677 = ~n1663 & ~n1676;
  assign n1678 = ~sys_fair4done_out & ~n1677;
  assign n1679 = ~n1660 & ~n1678;
  assign n1680 = ~reg_i_StoB_REQ5_out & ~n1679;
  assign n1681 = ~n1633 & ~n1680;
  assign n1682 = sys_fair5done_out & ~n1681;
  assign n1683 = reg_controllable_BtoS_ACK5_out & ~n973;
  assign n1684 = ~n1238 & ~n1683;
  assign n1685 = reg_i_StoB_REQ5_out & ~n1684;
  assign n1686 = ~n474 & ~n1241;
  assign n1687 = reg_i_StoB_REQ4_out & ~n1686;
  assign n1688 = ~reg_i_StoB_REQ4_out & ~n1667;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = reg_controllable_BtoS_ACK5_out & ~n1689;
  assign n1691 = ~n1217 & ~n1661;
  assign n1692 = reg_i_StoB_REQ4_out & ~n1691;
  assign n1693 = ~reg_i_StoB_REQ4_out & ~n1673;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = sys_fair4done_out & ~n1694;
  assign n1696 = ~n1678 & ~n1695;
  assign n1697 = ~reg_controllable_BtoS_ACK5_out & ~n1696;
  assign n1698 = ~n1690 & ~n1697;
  assign n1699 = ~reg_i_StoB_REQ5_out & ~n1698;
  assign n1700 = ~n1685 & ~n1699;
  assign n1701 = ~sys_fair5done_out & ~n1700;
  assign n1702 = ~n1682 & ~n1701;
  assign n1703 = ~reg_i_StoB_REQ8_out & ~n1702;
  assign n1704 = ~n1630 & ~n1703;
  assign n1705 = sys_fair8done_out & ~n1704;
  assign n1706 = reg_controllable_BtoS_ACK8_out & ~n986;
  assign n1707 = ~n1274 & ~n1706;
  assign n1708 = reg_i_StoB_REQ8_out & ~n1707;
  assign n1709 = ~n490 & ~n1277;
  assign n1710 = reg_i_StoB_REQ5_out & ~n1709;
  assign n1711 = ~reg_i_StoB_REQ5_out & ~n1689;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = reg_controllable_BtoS_ACK8_out & ~n1712;
  assign n1714 = ~n1253 & ~n1683;
  assign n1715 = reg_i_StoB_REQ5_out & ~n1714;
  assign n1716 = ~reg_i_StoB_REQ5_out & ~n1696;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = sys_fair5done_out & ~n1717;
  assign n1719 = ~n1701 & ~n1718;
  assign n1720 = ~reg_controllable_BtoS_ACK8_out & ~n1719;
  assign n1721 = ~n1713 & ~n1720;
  assign n1722 = ~reg_i_StoB_REQ8_out & ~n1721;
  assign n1723 = ~n1708 & ~n1722;
  assign n1724 = ~sys_fair8done_out & ~n1723;
  assign n1725 = ~n1705 & ~n1724;
  assign n1726 = ~reg_i_StoB_REQ6_out & ~n1725;
  assign n1727 = ~n1627 & ~n1726;
  assign n1728 = sys_fair6done_out & ~n1727;
  assign n1729 = reg_controllable_BtoS_ACK6_out & ~n999;
  assign n1730 = ~n1310 & ~n1729;
  assign n1731 = reg_i_StoB_REQ6_out & ~n1730;
  assign n1732 = ~n506 & ~n1313;
  assign n1733 = reg_i_StoB_REQ8_out & ~n1732;
  assign n1734 = ~reg_i_StoB_REQ8_out & ~n1712;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = reg_controllable_BtoS_ACK6_out & ~n1735;
  assign n1737 = ~n1289 & ~n1706;
  assign n1738 = reg_i_StoB_REQ8_out & ~n1737;
  assign n1739 = ~reg_i_StoB_REQ8_out & ~n1719;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = sys_fair8done_out & ~n1740;
  assign n1742 = ~n1724 & ~n1741;
  assign n1743 = ~reg_controllable_BtoS_ACK6_out & ~n1742;
  assign n1744 = ~n1736 & ~n1743;
  assign n1745 = ~reg_i_StoB_REQ6_out & ~n1744;
  assign n1746 = ~n1731 & ~n1745;
  assign n1747 = ~sys_fair6done_out & ~n1746;
  assign n1748 = ~n1728 & ~n1747;
  assign n1749 = sys_fair7done_out & ~n1748;
  assign n1750 = ~n522 & ~n1345;
  assign n1751 = reg_i_StoB_REQ6_out & ~n1750;
  assign n1752 = ~reg_i_StoB_REQ6_out & ~n1735;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~sys_fair7done_out & ~n1753;
  assign n1755 = ~n1749 & ~n1754;
  assign n1756 = reg_controllable_BtoS_ACK7_out & ~n1755;
  assign n1757 = ~n1325 & ~n1729;
  assign n1758 = reg_i_StoB_REQ6_out & ~n1757;
  assign n1759 = ~reg_i_StoB_REQ6_out & ~n1742;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = sys_fair6done_out & ~n1760;
  assign n1762 = ~n1747 & ~n1761;
  assign n1763 = ~sys_fair7done_out & ~n1762;
  assign n1764 = ~n1749 & ~n1763;
  assign n1765 = ~reg_controllable_BtoS_ACK7_out & ~n1764;
  assign n1766 = ~n1756 & ~n1765;
  assign n1767 = ~reg_i_StoB_REQ7_out & ~n1766;
  assign n1768 = ~n1624 & ~n1767;
  assign n1769 = ~reg_i_StoB_REQ9_out & ~n1768;
  assign n1770 = ~n1621 & ~n1769;
  assign n1771 = sys_fair9done_out & ~n1770;
  assign n1772 = reg_controllable_BtoS_ACK9_out & ~n1028;
  assign n1773 = ~n1382 & ~n1772;
  assign n1774 = reg_i_StoB_REQ9_out & ~n1773;
  assign n1775 = reg_controllable_BtoS_ACK7_out & ~n535;
  assign n1776 = ~n1386 & ~n1775;
  assign n1777 = reg_i_StoB_REQ7_out & ~n1776;
  assign n1778 = ~reg_i_StoB_REQ7_out & ~n1753;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = reg_controllable_BtoS_ACK9_out & ~n1779;
  assign n1781 = reg_controllable_BtoS_ACK7_out & ~n1012;
  assign n1782 = ~n1394 & ~n1781;
  assign n1783 = reg_i_StoB_REQ7_out & ~n1782;
  assign n1784 = sys_fair7done_out & ~n1762;
  assign n1785 = ~n1754 & ~n1784;
  assign n1786 = reg_controllable_BtoS_ACK7_out & ~n1785;
  assign n1787 = ~reg_controllable_BtoS_ACK7_out & ~n1762;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = ~reg_i_StoB_REQ7_out & ~n1788;
  assign n1790 = ~n1783 & ~n1789;
  assign n1791 = ~reg_controllable_BtoS_ACK9_out & ~n1790;
  assign n1792 = ~n1780 & ~n1791;
  assign n1793 = ~reg_i_StoB_REQ9_out & ~n1792;
  assign n1794 = ~n1774 & ~n1793;
  assign n1795 = ~sys_fair9done_out & ~n1794;
  assign n1796 = ~n1771 & ~n1795;
  assign n1797 = ~reg_i_StoB_REQ11_out & ~n1796;
  assign n1798 = ~n1618 & ~n1797;
  assign n1799 = sys_fair11done_out & ~n1798;
  assign n1800 = reg_controllable_BtoS_ACK11_out & ~n1041;
  assign n1801 = ~n1424 & ~n1800;
  assign n1802 = reg_i_StoB_REQ11_out & ~n1801;
  assign n1803 = ~n554 & ~n1427;
  assign n1804 = reg_i_StoB_REQ9_out & ~n1803;
  assign n1805 = ~reg_i_StoB_REQ9_out & ~n1779;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = reg_controllable_BtoS_ACK11_out & ~n1806;
  assign n1808 = ~n1403 & ~n1772;
  assign n1809 = reg_i_StoB_REQ9_out & ~n1808;
  assign n1810 = ~reg_i_StoB_REQ9_out & ~n1790;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = sys_fair9done_out & ~n1811;
  assign n1813 = ~n1795 & ~n1812;
  assign n1814 = ~reg_controllable_BtoS_ACK11_out & ~n1813;
  assign n1815 = ~n1807 & ~n1814;
  assign n1816 = ~reg_i_StoB_REQ11_out & ~n1815;
  assign n1817 = ~n1802 & ~n1816;
  assign n1818 = ~sys_fair11done_out & ~n1817;
  assign n1819 = ~n1799 & ~n1818;
  assign n1820 = sys_fair12done_out & ~n1819;
  assign n1821 = ~n573 & ~n1459;
  assign n1822 = reg_i_StoB_REQ11_out & ~n1821;
  assign n1823 = ~reg_i_StoB_REQ11_out & ~n1806;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~sys_fair12done_out & ~n1824;
  assign n1826 = ~n1820 & ~n1825;
  assign n1827 = reg_controllable_BtoS_ACK12_out & ~n1826;
  assign n1828 = ~n1439 & ~n1800;
  assign n1829 = reg_i_StoB_REQ11_out & ~n1828;
  assign n1830 = ~reg_i_StoB_REQ11_out & ~n1813;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = sys_fair11done_out & ~n1831;
  assign n1833 = ~n1818 & ~n1832;
  assign n1834 = ~sys_fair12done_out & ~n1833;
  assign n1835 = ~n1820 & ~n1834;
  assign n1836 = ~reg_controllable_BtoS_ACK12_out & ~n1835;
  assign n1837 = ~n1827 & ~n1836;
  assign n1838 = ~reg_i_StoB_REQ12_out & ~n1837;
  assign n1839 = ~n1615 & ~n1838;
  assign n1840 = ~reg_i_StoB_REQ13_out & ~n1839;
  assign n1841 = ~n1612 & ~n1840;
  assign n1842 = sys_fair13done_out & ~n1841;
  assign n1843 = reg_controllable_BtoS_ACK13_out & ~n1070;
  assign n1844 = ~n1496 & ~n1843;
  assign n1845 = reg_i_StoB_REQ13_out & ~n1844;
  assign n1846 = reg_controllable_BtoS_ACK12_out & ~n586;
  assign n1847 = ~n1500 & ~n1846;
  assign n1848 = reg_i_StoB_REQ12_out & ~n1847;
  assign n1849 = ~reg_i_StoB_REQ12_out & ~n1824;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = reg_controllable_BtoS_ACK13_out & ~n1850;
  assign n1852 = reg_controllable_BtoS_ACK12_out & ~n1054;
  assign n1853 = ~n1508 & ~n1852;
  assign n1854 = reg_i_StoB_REQ12_out & ~n1853;
  assign n1855 = sys_fair12done_out & ~n1833;
  assign n1856 = ~n1825 & ~n1855;
  assign n1857 = reg_controllable_BtoS_ACK12_out & ~n1856;
  assign n1858 = ~reg_controllable_BtoS_ACK12_out & ~n1833;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~reg_i_StoB_REQ12_out & ~n1859;
  assign n1861 = ~n1854 & ~n1860;
  assign n1862 = ~reg_controllable_BtoS_ACK13_out & ~n1861;
  assign n1863 = ~n1851 & ~n1862;
  assign n1864 = ~reg_i_StoB_REQ13_out & ~n1863;
  assign n1865 = ~n1845 & ~n1864;
  assign n1866 = ~sys_fair13done_out & ~n1865;
  assign n1867 = ~n1842 & ~n1866;
  assign n1868 = sys_fair0done_out & ~n1867;
  assign n1869 = ~n605 & ~n1537;
  assign n1870 = reg_i_StoB_REQ13_out & ~n1869;
  assign n1871 = ~reg_i_StoB_REQ13_out & ~n1850;
  assign n1872 = ~n1870 & ~n1871;
  assign n1873 = ~sys_fair0done_out & ~n1872;
  assign n1874 = ~n1868 & ~n1873;
  assign n1875 = reg_controllable_BtoS_ACK0_out & ~n1874;
  assign n1876 = ~n1517 & ~n1843;
  assign n1877 = reg_i_StoB_REQ13_out & ~n1876;
  assign n1878 = ~reg_i_StoB_REQ13_out & ~n1861;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = sys_fair13done_out & ~n1879;
  assign n1881 = ~n1866 & ~n1880;
  assign n1882 = ~sys_fair0done_out & ~n1881;
  assign n1883 = ~n1868 & ~n1882;
  assign n1884 = ~reg_controllable_BtoS_ACK0_out & ~n1883;
  assign n1885 = ~n1875 & ~n1884;
  assign n1886 = ~reg_i_StoB_REQ0_out & ~n1885;
  assign n1887 = ~n1609 & ~n1886;
  assign n1888 = ~reg_i_StoB_REQ10_out & ~n1887;
  assign n1889 = ~n1606 & ~n1888;
  assign n1890 = sys_fair10done_out & ~n1889;
  assign n1891 = reg_controllable_BtoS_ACK10_out & ~n1111;
  assign n1892 = ~n1574 & ~n1891;
  assign n1893 = reg_i_StoB_REQ10_out & ~n1892;
  assign n1894 = reg_controllable_BtoS_ACK0_out & ~n621;
  assign n1895 = ~n1578 & ~n1894;
  assign n1896 = reg_i_StoB_REQ0_out & ~n1895;
  assign n1897 = ~reg_i_StoB_REQ0_out & ~n1872;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = reg_controllable_BtoS_ACK10_out & ~n1898;
  assign n1900 = reg_controllable_BtoS_ACK0_out & ~n1083;
  assign n1901 = ~n1586 & ~n1900;
  assign n1902 = reg_i_StoB_REQ0_out & ~n1901;
  assign n1903 = sys_fair0done_out & ~n1881;
  assign n1904 = ~n1873 & ~n1903;
  assign n1905 = reg_controllable_BtoS_ACK0_out & ~n1904;
  assign n1906 = ~reg_controllable_BtoS_ACK0_out & ~n1881;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~reg_i_StoB_REQ0_out & ~n1907;
  assign n1909 = ~n1902 & ~n1908;
  assign n1910 = ~reg_controllable_BtoS_ACK10_out & ~n1909;
  assign n1911 = ~n1899 & ~n1910;
  assign n1912 = ~reg_i_StoB_REQ10_out & ~n1911;
  assign n1913 = ~n1893 & ~n1912;
  assign n1914 = ~sys_fair10done_out & ~n1913;
  assign n1915 = ~n1890 & ~n1914;
  assign n1916 = ~reg_i_StoB_REQ14_out & ~n1915;
  assign n1917 = ~n1603 & ~n1916;
  assign n1918 = sys_fair14done_out & ~n1917;
  assign n1919 = ~reg_i_StoB_REQ10_out & ~n1111;
  assign n1920 = ~n1104 & ~n1919;
  assign n1921 = sys_fair10done_out & ~n1920;
  assign n1922 = ~n1116 & ~n1921;
  assign n1923 = reg_controllable_BtoS_ACK14_out & ~n1922;
  assign n1924 = ~reg_i_StoB_REQ10_out & ~n1573;
  assign n1925 = ~n1576 & ~n1924;
  assign n1926 = sys_fair10done_out & ~n1925;
  assign n1927 = ~n1574 & ~n1583;
  assign n1928 = ~reg_i_StoB_REQ10_out & ~n1927;
  assign n1929 = ~n1576 & ~n1928;
  assign n1930 = ~sys_fair10done_out & ~n1929;
  assign n1931 = ~n1926 & ~n1930;
  assign n1932 = ~reg_controllable_BtoS_ACK14_out & ~n1931;
  assign n1933 = ~n1923 & ~n1932;
  assign n1934 = reg_i_StoB_REQ14_out & ~n1933;
  assign n1935 = ~reg_controllable_BtoS_ACK10_out & ~n1582;
  assign n1936 = ~n640 & ~n1935;
  assign n1937 = reg_i_StoB_REQ10_out & ~n1936;
  assign n1938 = ~reg_i_StoB_REQ10_out & ~n1898;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = reg_controllable_BtoS_ACK14_out & ~n1939;
  assign n1941 = ~n1595 & ~n1891;
  assign n1942 = reg_i_StoB_REQ10_out & ~n1941;
  assign n1943 = ~reg_i_StoB_REQ10_out & ~n1909;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = sys_fair10done_out & ~n1944;
  assign n1946 = ~n1914 & ~n1945;
  assign n1947 = ~reg_controllable_BtoS_ACK14_out & ~n1946;
  assign n1948 = ~n1940 & ~n1947;
  assign n1949 = ~reg_i_StoB_REQ14_out & ~n1948;
  assign n1950 = ~n1934 & ~n1949;
  assign n1951 = ~sys_fair14done_out & ~n1950;
  assign n1952 = ~n1918 & ~n1951;
  assign n1953 = sys_fair15done_out & ~n1952;
  assign n1954 = ~n1563 & ~n1595;
  assign n1955 = reg_i_StoB_REQ10_out & ~n1954;
  assign n1956 = ~reg_i_StoB_REQ10_out & ~n1594;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = sys_fair10done_out & ~n1957;
  assign n1959 = ~n1599 & ~n1958;
  assign n1960 = ~reg_controllable_BtoS_ACK14_out & ~n1959;
  assign n1961 = ~n1923 & ~n1960;
  assign n1962 = reg_i_StoB_REQ14_out & ~n1961;
  assign n1963 = ~reg_i_StoB_REQ14_out & ~n1946;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = sys_fair14done_out & ~n1964;
  assign n1966 = ~n1951 & ~n1965;
  assign n1967 = reg_stateG12_out & ~n1966;
  assign n1968 = ~n419 & ~n1935;
  assign n1969 = reg_i_StoB_REQ10_out & ~n1968;
  assign n1970 = ~reg_i_StoB_REQ10_out & ~n1582;
  assign n1971 = ~n1969 & ~n1970;
  assign n1972 = ~reg_controllable_BtoS_ACK14_out & ~n1971;
  assign n1973 = ~n664 & ~n1972;
  assign n1974 = reg_i_StoB_REQ14_out & ~n1973;
  assign n1975 = ~reg_i_StoB_REQ14_out & ~n1939;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~reg_stateG12_out & ~n1976;
  assign n1978 = ~n1967 & ~n1977;
  assign n1979 = ~sys_fair15done_out & ~n1978;
  assign n1980 = ~n1953 & ~n1979;
  assign n1981 = fair_cnt<1>_out  & ~n1980;
  assign n1982 = ~fair_cnt<1>_out  & ~n1976;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = fair_cnt<0>_out  & ~n1983;
  assign n1985 = ~fair_cnt<0>_out  & ~n1976;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~reg_i_RtoB_ACK1_out & ~n1986;
  assign n1988 = ~n711 & ~n1987;
  assign n1989 = reg_i_RtoB_ACK0_out & ~n1988;
  assign n1990 = ~reg_i_StoB_REQ10_out & ~n927;
  assign n1991 = ~n930 & ~n1990;
  assign n1992 = sys_fair10done_out & ~n1991;
  assign n1993 = ~n419 & ~n1102;
  assign n1994 = ~reg_i_StoB_REQ10_out & ~n1993;
  assign n1995 = ~n1104 & ~n1994;
  assign n1996 = ~sys_fair10done_out & ~n1995;
  assign n1997 = ~n1992 & ~n1996;
  assign n1998 = reg_controllable_BtoS_ACK14_out & ~n1997;
  assign n1999 = ~reg_i_StoB_REQ2_out & ~n1133;
  assign n2000 = ~sys_fair2done_out & ~n1999;
  assign n2001 = ~n1132 & ~n2000;
  assign n2002 = sys_fair1done_out & ~n2001;
  assign n2003 = sys_fair2done_out & ~n716;
  assign n2004 = reg_i_StoB_REQ2_out & ~n716;
  assign n2005 = ~reg_controllable_BtoS_ACK2_out & n716;
  assign n2006 = ~reg_controllable_BtoS_ACK2_out & ~n2005;
  assign n2007 = ~reg_i_StoB_REQ2_out & n2006;
  assign n2008 = ~n2004 & ~n2007;
  assign n2009 = ~sys_fair2done_out & ~n2008;
  assign n2010 = ~n2003 & ~n2009;
  assign n2011 = ~sys_fair1done_out & ~n2010;
  assign n2012 = ~n2002 & ~n2011;
  assign n2013 = ~reg_controllable_BtoS_ACK3_out & ~n2012;
  assign n2014 = ~n1130 & ~n2013;
  assign n2015 = reg_i_StoB_REQ3_out & ~n2014;
  assign n2016 = ~reg_i_StoB_REQ3_out & ~n2012;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = sys_fair3done_out & ~n2017;
  assign n2019 = ~sys_fair2done_out & ~n2000;
  assign n2020 = sys_fair1done_out & ~n2019;
  assign n2021 = ~n2011 & ~n2020;
  assign n2022 = ~reg_controllable_BtoS_ACK3_out & ~n2021;
  assign n2023 = ~n1159 & ~n2022;
  assign n2024 = reg_i_StoB_REQ3_out & ~n2023;
  assign n2025 = ~n1177 & ~n2022;
  assign n2026 = ~reg_i_StoB_REQ3_out & ~n2025;
  assign n2027 = ~n2024 & ~n2026;
  assign n2028 = ~sys_fair3done_out & ~n2027;
  assign n2029 = ~n2018 & ~n2028;
  assign n2030 = ~reg_controllable_BtoS_ACK4_out & ~n2029;
  assign n2031 = ~n1129 & ~n2030;
  assign n2032 = reg_i_StoB_REQ4_out & ~n2031;
  assign n2033 = ~reg_i_StoB_REQ4_out & ~n2029;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = sys_fair4done_out & ~n2034;
  assign n2036 = ~reg_i_StoB_REQ3_out & ~n2021;
  assign n2037 = ~n2024 & ~n2036;
  assign n2038 = sys_fair3done_out & ~n2037;
  assign n2039 = ~n2028 & ~n2038;
  assign n2040 = ~reg_controllable_BtoS_ACK4_out & ~n2039;
  assign n2041 = ~n1193 & ~n2040;
  assign n2042 = reg_i_StoB_REQ4_out & ~n2041;
  assign n2043 = ~n1210 & ~n2040;
  assign n2044 = ~reg_i_StoB_REQ4_out & ~n2043;
  assign n2045 = ~n2042 & ~n2044;
  assign n2046 = ~sys_fair4done_out & ~n2045;
  assign n2047 = ~n2035 & ~n2046;
  assign n2048 = ~reg_controllable_BtoS_ACK5_out & ~n2047;
  assign n2049 = ~n1128 & ~n2048;
  assign n2050 = reg_i_StoB_REQ5_out & ~n2049;
  assign n2051 = ~reg_i_StoB_REQ5_out & ~n2047;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = sys_fair5done_out & ~n2052;
  assign n2054 = ~reg_i_StoB_REQ4_out & ~n2039;
  assign n2055 = ~n2042 & ~n2054;
  assign n2056 = sys_fair4done_out & ~n2055;
  assign n2057 = ~n2046 & ~n2056;
  assign n2058 = ~reg_controllable_BtoS_ACK5_out & ~n2057;
  assign n2059 = ~n1229 & ~n2058;
  assign n2060 = reg_i_StoB_REQ5_out & ~n2059;
  assign n2061 = ~n1246 & ~n2058;
  assign n2062 = ~reg_i_StoB_REQ5_out & ~n2061;
  assign n2063 = ~n2060 & ~n2062;
  assign n2064 = ~sys_fair5done_out & ~n2063;
  assign n2065 = ~n2053 & ~n2064;
  assign n2066 = ~reg_controllable_BtoS_ACK8_out & ~n2065;
  assign n2067 = ~n1127 & ~n2066;
  assign n2068 = reg_i_StoB_REQ8_out & ~n2067;
  assign n2069 = ~reg_i_StoB_REQ8_out & ~n2065;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = sys_fair8done_out & ~n2070;
  assign n2072 = ~reg_i_StoB_REQ5_out & ~n2057;
  assign n2073 = ~n2060 & ~n2072;
  assign n2074 = sys_fair5done_out & ~n2073;
  assign n2075 = ~n2064 & ~n2074;
  assign n2076 = ~reg_controllable_BtoS_ACK8_out & ~n2075;
  assign n2077 = ~n1265 & ~n2076;
  assign n2078 = reg_i_StoB_REQ8_out & ~n2077;
  assign n2079 = ~n1282 & ~n2076;
  assign n2080 = ~reg_i_StoB_REQ8_out & ~n2079;
  assign n2081 = ~n2078 & ~n2080;
  assign n2082 = ~sys_fair8done_out & ~n2081;
  assign n2083 = ~n2071 & ~n2082;
  assign n2084 = ~reg_controllable_BtoS_ACK6_out & ~n2083;
  assign n2085 = ~n1126 & ~n2084;
  assign n2086 = reg_i_StoB_REQ6_out & ~n2085;
  assign n2087 = ~reg_i_StoB_REQ6_out & ~n2083;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = sys_fair6done_out & ~n2088;
  assign n2090 = ~reg_i_StoB_REQ8_out & ~n2075;
  assign n2091 = ~n2078 & ~n2090;
  assign n2092 = sys_fair8done_out & ~n2091;
  assign n2093 = ~n2082 & ~n2092;
  assign n2094 = ~reg_controllable_BtoS_ACK6_out & ~n2093;
  assign n2095 = ~n1301 & ~n2094;
  assign n2096 = reg_i_StoB_REQ6_out & ~n2095;
  assign n2097 = ~n1318 & ~n2094;
  assign n2098 = ~reg_i_StoB_REQ6_out & ~n2097;
  assign n2099 = ~n2096 & ~n2098;
  assign n2100 = ~sys_fair6done_out & ~n2099;
  assign n2101 = ~n2089 & ~n2100;
  assign n2102 = sys_fair7done_out & ~n2101;
  assign n2103 = ~reg_i_StoB_REQ6_out & ~n2093;
  assign n2104 = ~n2096 & ~n2103;
  assign n2105 = sys_fair6done_out & ~n2104;
  assign n2106 = ~n2100 & ~n2105;
  assign n2107 = ~sys_fair7done_out & ~n2106;
  assign n2108 = ~n2102 & ~n2107;
  assign n2109 = ~reg_controllable_BtoS_ACK7_out & ~n2108;
  assign n2110 = ~n1125 & ~n2109;
  assign n2111 = reg_i_StoB_REQ7_out & ~n2110;
  assign n2112 = ~n1350 & ~n2102;
  assign n2113 = reg_controllable_BtoS_ACK7_out & ~n2112;
  assign n2114 = ~n2109 & ~n2113;
  assign n2115 = ~reg_i_StoB_REQ7_out & ~n2114;
  assign n2116 = ~n2111 & ~n2115;
  assign n2117 = ~reg_controllable_BtoS_ACK9_out & ~n2116;
  assign n2118 = ~n1124 & ~n2117;
  assign n2119 = reg_i_StoB_REQ9_out & ~n2118;
  assign n2120 = ~reg_i_StoB_REQ9_out & ~n2116;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = sys_fair9done_out & ~n2121;
  assign n2123 = ~reg_controllable_BtoS_ACK7_out & ~n2106;
  assign n2124 = ~n1372 & ~n2123;
  assign n2125 = reg_i_StoB_REQ7_out & ~n2124;
  assign n2126 = sys_fair7done_out & ~n2106;
  assign n2127 = ~n1350 & ~n2126;
  assign n2128 = reg_controllable_BtoS_ACK7_out & ~n2127;
  assign n2129 = ~n2123 & ~n2128;
  assign n2130 = ~reg_i_StoB_REQ7_out & ~n2129;
  assign n2131 = ~n2125 & ~n2130;
  assign n2132 = ~reg_controllable_BtoS_ACK9_out & ~n2131;
  assign n2133 = ~n1371 & ~n2132;
  assign n2134 = reg_i_StoB_REQ9_out & ~n2133;
  assign n2135 = ~n1391 & ~n2132;
  assign n2136 = ~reg_i_StoB_REQ9_out & ~n2135;
  assign n2137 = ~n2134 & ~n2136;
  assign n2138 = ~sys_fair9done_out & ~n2137;
  assign n2139 = ~n2122 & ~n2138;
  assign n2140 = ~reg_controllable_BtoS_ACK11_out & ~n2139;
  assign n2141 = ~n1123 & ~n2140;
  assign n2142 = reg_i_StoB_REQ11_out & ~n2141;
  assign n2143 = ~reg_i_StoB_REQ11_out & ~n2139;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = sys_fair11done_out & ~n2144;
  assign n2146 = ~reg_i_StoB_REQ9_out & ~n2131;
  assign n2147 = ~n2134 & ~n2146;
  assign n2148 = sys_fair9done_out & ~n2147;
  assign n2149 = ~n2138 & ~n2148;
  assign n2150 = ~reg_controllable_BtoS_ACK11_out & ~n2149;
  assign n2151 = ~n1415 & ~n2150;
  assign n2152 = reg_i_StoB_REQ11_out & ~n2151;
  assign n2153 = ~n1432 & ~n2150;
  assign n2154 = ~reg_i_StoB_REQ11_out & ~n2153;
  assign n2155 = ~n2152 & ~n2154;
  assign n2156 = ~sys_fair11done_out & ~n2155;
  assign n2157 = ~n2145 & ~n2156;
  assign n2158 = sys_fair12done_out & ~n2157;
  assign n2159 = ~reg_i_StoB_REQ11_out & ~n2149;
  assign n2160 = ~n2152 & ~n2159;
  assign n2161 = sys_fair11done_out & ~n2160;
  assign n2162 = ~n2156 & ~n2161;
  assign n2163 = ~sys_fair12done_out & ~n2162;
  assign n2164 = ~n2158 & ~n2163;
  assign n2165 = ~reg_controllable_BtoS_ACK12_out & ~n2164;
  assign n2166 = ~n1122 & ~n2165;
  assign n2167 = reg_i_StoB_REQ12_out & ~n2166;
  assign n2168 = ~n1464 & ~n2158;
  assign n2169 = reg_controllable_BtoS_ACK12_out & ~n2168;
  assign n2170 = ~n2165 & ~n2169;
  assign n2171 = ~reg_i_StoB_REQ12_out & ~n2170;
  assign n2172 = ~n2167 & ~n2171;
  assign n2173 = ~reg_controllable_BtoS_ACK13_out & ~n2172;
  assign n2174 = ~n1121 & ~n2173;
  assign n2175 = reg_i_StoB_REQ13_out & ~n2174;
  assign n2176 = ~reg_i_StoB_REQ13_out & ~n2172;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = sys_fair13done_out & ~n2177;
  assign n2179 = ~reg_controllable_BtoS_ACK12_out & ~n2162;
  assign n2180 = ~n1486 & ~n2179;
  assign n2181 = reg_i_StoB_REQ12_out & ~n2180;
  assign n2182 = sys_fair12done_out & ~n2162;
  assign n2183 = ~n1464 & ~n2182;
  assign n2184 = reg_controllable_BtoS_ACK12_out & ~n2183;
  assign n2185 = ~n2179 & ~n2184;
  assign n2186 = ~reg_i_StoB_REQ12_out & ~n2185;
  assign n2187 = ~n2181 & ~n2186;
  assign n2188 = ~reg_controllable_BtoS_ACK13_out & ~n2187;
  assign n2189 = ~n1485 & ~n2188;
  assign n2190 = reg_i_StoB_REQ13_out & ~n2189;
  assign n2191 = ~n1505 & ~n2188;
  assign n2192 = ~reg_i_StoB_REQ13_out & ~n2191;
  assign n2193 = ~n2190 & ~n2192;
  assign n2194 = ~sys_fair13done_out & ~n2193;
  assign n2195 = ~n2178 & ~n2194;
  assign n2196 = sys_fair0done_out & ~n2195;
  assign n2197 = ~reg_i_StoB_REQ13_out & ~n2187;
  assign n2198 = ~n2190 & ~n2197;
  assign n2199 = sys_fair13done_out & ~n2198;
  assign n2200 = ~n2194 & ~n2199;
  assign n2201 = ~sys_fair0done_out & ~n2200;
  assign n2202 = ~n2196 & ~n2201;
  assign n2203 = ~reg_controllable_BtoS_ACK0_out & ~n2202;
  assign n2204 = ~n1120 & ~n2203;
  assign n2205 = reg_i_StoB_REQ0_out & ~n2204;
  assign n2206 = ~n1542 & ~n2196;
  assign n2207 = reg_controllable_BtoS_ACK0_out & ~n2206;
  assign n2208 = ~n2203 & ~n2207;
  assign n2209 = ~reg_i_StoB_REQ0_out & ~n2208;
  assign n2210 = ~n2205 & ~n2209;
  assign n2211 = ~reg_controllable_BtoS_ACK10_out & ~n2210;
  assign n2212 = ~n1119 & ~n2211;
  assign n2213 = reg_i_StoB_REQ10_out & ~n2212;
  assign n2214 = ~reg_i_StoB_REQ10_out & ~n2210;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = sys_fair10done_out & ~n2215;
  assign n2217 = ~reg_controllable_BtoS_ACK0_out & ~n2200;
  assign n2218 = ~n1564 & ~n2217;
  assign n2219 = reg_i_StoB_REQ0_out & ~n2218;
  assign n2220 = sys_fair0done_out & ~n2200;
  assign n2221 = ~n1542 & ~n2220;
  assign n2222 = reg_controllable_BtoS_ACK0_out & ~n2221;
  assign n2223 = ~n2217 & ~n2222;
  assign n2224 = ~reg_i_StoB_REQ0_out & ~n2223;
  assign n2225 = ~n2219 & ~n2224;
  assign n2226 = ~reg_controllable_BtoS_ACK10_out & ~n2225;
  assign n2227 = ~n1563 & ~n2226;
  assign n2228 = reg_i_StoB_REQ10_out & ~n2227;
  assign n2229 = ~n1583 & ~n2226;
  assign n2230 = ~reg_i_StoB_REQ10_out & ~n2229;
  assign n2231 = ~n2228 & ~n2230;
  assign n2232 = ~sys_fair10done_out & ~n2231;
  assign n2233 = ~n2216 & ~n2232;
  assign n2234 = ~reg_controllable_BtoS_ACK14_out & ~n2233;
  assign n2235 = ~n1998 & ~n2234;
  assign n2236 = reg_i_StoB_REQ14_out & ~n2235;
  assign n2237 = ~reg_i_StoB_REQ14_out & ~n2233;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = sys_fair14done_out & ~n2238;
  assign n2240 = ~reg_i_StoB_REQ10_out & ~n1101;
  assign n2241 = ~n1104 & ~n2240;
  assign n2242 = sys_fair10done_out & ~n2241;
  assign n2243 = ~n1996 & ~n2242;
  assign n2244 = reg_controllable_BtoS_ACK14_out & ~n2243;
  assign n2245 = ~reg_i_StoB_REQ10_out & ~n2225;
  assign n2246 = ~n2228 & ~n2245;
  assign n2247 = sys_fair10done_out & ~n2246;
  assign n2248 = ~n2232 & ~n2247;
  assign n2249 = ~reg_controllable_BtoS_ACK14_out & ~n2248;
  assign n2250 = ~n2244 & ~n2249;
  assign n2251 = reg_i_StoB_REQ14_out & ~n2250;
  assign n2252 = reg_controllable_BtoS_ACK14_out & ~n1971;
  assign n2253 = ~n2249 & ~n2252;
  assign n2254 = ~reg_i_StoB_REQ14_out & ~n2253;
  assign n2255 = ~n2251 & ~n2254;
  assign n2256 = ~sys_fair14done_out & ~n2255;
  assign n2257 = ~n2239 & ~n2256;
  assign n2258 = sys_fair15done_out & ~n2257;
  assign n2259 = ~reg_i_StoB_REQ14_out & ~n2248;
  assign n2260 = ~n2251 & ~n2259;
  assign n2261 = sys_fair14done_out & ~n2260;
  assign n2262 = ~n2256 & ~n2261;
  assign n2263 = reg_stateG12_out & ~n2262;
  assign n2264 = reg_controllable_BtoS_ACK14_out & ~n658;
  assign n2265 = ~n1972 & ~n2264;
  assign n2266 = reg_i_StoB_REQ14_out & ~n2265;
  assign n2267 = ~reg_i_StoB_REQ14_out & ~n1971;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = ~reg_stateG12_out & ~n2268;
  assign n2270 = ~n2263 & ~n2269;
  assign n2271 = ~sys_fair15done_out & ~n2270;
  assign n2272 = ~n2258 & ~n2271;
  assign n2273 = fair_cnt<1>_out  & ~n2272;
  assign n2274 = ~fair_cnt<1>_out  & ~n2268;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = fair_cnt<0>_out  & ~n2275;
  assign n2277 = ~fair_cnt<0>_out  & ~n2268;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = env_fair1done_out & ~n2278;
  assign n2280 = ~env_fair1done_out & ~n2268;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = env_fair0done_out & ~n2281;
  assign n2283 = sys_fair0done_out & ~n386;
  assign n2284 = ~sys_fair2done_out & ~n117;
  assign n2285 = ~n442 & ~n2284;
  assign n2286 = sys_fair1done_out & ~n2285;
  assign n2287 = ~sys_fair1done_out & ~n117;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~reg_i_StoB_REQ3_out & ~n2288;
  assign n2290 = ~n149 & ~n2289;
  assign n2291 = sys_fair3done_out & ~n2290;
  assign n2292 = ~sys_fair3done_out & ~n167;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~reg_i_StoB_REQ4_out & ~n2293;
  assign n2295 = ~n170 & ~n2294;
  assign n2296 = sys_fair4done_out & ~n2295;
  assign n2297 = ~sys_fair4done_out & ~n191;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = ~reg_i_StoB_REQ5_out & ~n2298;
  assign n2300 = ~n194 & ~n2299;
  assign n2301 = sys_fair5done_out & ~n2300;
  assign n2302 = ~sys_fair5done_out & ~n215;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~reg_i_StoB_REQ8_out & ~n2303;
  assign n2305 = ~n218 & ~n2304;
  assign n2306 = sys_fair8done_out & ~n2305;
  assign n2307 = ~sys_fair8done_out & ~n239;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~reg_i_StoB_REQ6_out & ~n2308;
  assign n2310 = ~n242 & ~n2309;
  assign n2311 = sys_fair6done_out & ~n2310;
  assign n2312 = ~sys_fair6done_out & ~n258;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = sys_fair7done_out & ~n2313;
  assign n2315 = ~n259 & ~n2314;
  assign n2316 = ~reg_i_StoB_REQ7_out & ~n2315;
  assign n2317 = ~n285 & ~n2316;
  assign n2318 = ~reg_i_StoB_REQ9_out & ~n2317;
  assign n2319 = ~n290 & ~n2318;
  assign n2320 = sys_fair9done_out & ~n2319;
  assign n2321 = ~sys_fair9done_out & ~n315;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = ~reg_i_StoB_REQ11_out & ~n2322;
  assign n2324 = ~n318 & ~n2323;
  assign n2325 = sys_fair11done_out & ~n2324;
  assign n2326 = ~sys_fair11done_out & ~n334;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = sys_fair12done_out & ~n2327;
  assign n2329 = ~n335 & ~n2328;
  assign n2330 = ~reg_i_StoB_REQ12_out & ~n2329;
  assign n2331 = ~n361 & ~n2330;
  assign n2332 = ~reg_i_StoB_REQ13_out & ~n2331;
  assign n2333 = ~n366 & ~n2332;
  assign n2334 = sys_fair13done_out & ~n2333;
  assign n2335 = ~sys_fair13done_out & ~n386;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = ~sys_fair0done_out & ~n2336;
  assign n2338 = ~n2283 & ~n2337;
  assign n2339 = reg_controllable_BtoS_ACK0_out & ~n2338;
  assign n2340 = ~n1578 & ~n2339;
  assign n2341 = reg_i_StoB_REQ0_out & ~n2340;
  assign n2342 = sys_fair12done_out & ~n334;
  assign n2343 = ~sys_fair12done_out & ~n2327;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = reg_controllable_BtoS_ACK12_out & ~n2344;
  assign n2346 = ~n1500 & ~n2345;
  assign n2347 = reg_i_StoB_REQ12_out & ~n2346;
  assign n2348 = sys_fair7done_out & ~n258;
  assign n2349 = ~sys_fair7done_out & ~n2313;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = reg_controllable_BtoS_ACK7_out & ~n2350;
  assign n2352 = ~n1386 & ~n2351;
  assign n2353 = reg_i_StoB_REQ7_out & ~n2352;
  assign n2354 = ~sys_fair2done_out & n1640;
  assign n2355 = ~n1132 & ~n2354;
  assign n2356 = sys_fair1done_out & ~n2355;
  assign n2357 = ~n116 & ~n1131;
  assign n2358 = sys_fair2done_out & ~n2357;
  assign n2359 = ~sys_fair2done_out & n1131;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~sys_fair1done_out & ~n2360;
  assign n2362 = ~n2356 & ~n2361;
  assign n2363 = ~reg_i_StoB_REQ3_out & ~n2362;
  assign n2364 = ~n1207 & ~n2363;
  assign n2365 = sys_fair3done_out & ~n2364;
  assign n2366 = reg_controllable_BtoS_ACK3_out & ~n2288;
  assign n2367 = ~n1205 & ~n2366;
  assign n2368 = reg_i_StoB_REQ3_out & ~n2367;
  assign n2369 = ~n1208 & ~n2368;
  assign n2370 = ~sys_fair3done_out & ~n2369;
  assign n2371 = ~n2365 & ~n2370;
  assign n2372 = ~reg_i_StoB_REQ4_out & ~n2371;
  assign n2373 = ~n1243 & ~n2372;
  assign n2374 = sys_fair4done_out & ~n2373;
  assign n2375 = reg_controllable_BtoS_ACK4_out & ~n2293;
  assign n2376 = ~n1241 & ~n2375;
  assign n2377 = reg_i_StoB_REQ4_out & ~n2376;
  assign n2378 = ~n1244 & ~n2377;
  assign n2379 = ~sys_fair4done_out & ~n2378;
  assign n2380 = ~n2374 & ~n2379;
  assign n2381 = ~reg_i_StoB_REQ5_out & ~n2380;
  assign n2382 = ~n1279 & ~n2381;
  assign n2383 = sys_fair5done_out & ~n2382;
  assign n2384 = reg_controllable_BtoS_ACK5_out & ~n2298;
  assign n2385 = ~n1277 & ~n2384;
  assign n2386 = reg_i_StoB_REQ5_out & ~n2385;
  assign n2387 = ~n1280 & ~n2386;
  assign n2388 = ~sys_fair5done_out & ~n2387;
  assign n2389 = ~n2383 & ~n2388;
  assign n2390 = ~reg_i_StoB_REQ8_out & ~n2389;
  assign n2391 = ~n1315 & ~n2390;
  assign n2392 = sys_fair8done_out & ~n2391;
  assign n2393 = reg_controllable_BtoS_ACK8_out & ~n2303;
  assign n2394 = ~n1313 & ~n2393;
  assign n2395 = reg_i_StoB_REQ8_out & ~n2394;
  assign n2396 = ~n1316 & ~n2395;
  assign n2397 = ~sys_fair8done_out & ~n2396;
  assign n2398 = ~n2392 & ~n2397;
  assign n2399 = ~reg_i_StoB_REQ6_out & ~n2398;
  assign n2400 = ~n1347 & ~n2399;
  assign n2401 = sys_fair6done_out & ~n2400;
  assign n2402 = reg_controllable_BtoS_ACK6_out & ~n2308;
  assign n2403 = ~n1345 & ~n2402;
  assign n2404 = reg_i_StoB_REQ6_out & ~n2403;
  assign n2405 = ~n1348 & ~n2404;
  assign n2406 = ~sys_fair6done_out & ~n2405;
  assign n2407 = ~n2401 & ~n2406;
  assign n2408 = sys_fair7done_out & ~n2407;
  assign n2409 = ~n1350 & ~n2408;
  assign n2410 = ~reg_i_StoB_REQ7_out & ~n2409;
  assign n2411 = ~n2353 & ~n2410;
  assign n2412 = ~reg_i_StoB_REQ9_out & ~n2411;
  assign n2413 = ~n1429 & ~n2412;
  assign n2414 = sys_fair9done_out & ~n2413;
  assign n2415 = reg_controllable_BtoS_ACK9_out & ~n2317;
  assign n2416 = ~n1427 & ~n2415;
  assign n2417 = reg_i_StoB_REQ9_out & ~n2416;
  assign n2418 = ~n1430 & ~n2417;
  assign n2419 = ~sys_fair9done_out & ~n2418;
  assign n2420 = ~n2414 & ~n2419;
  assign n2421 = ~reg_i_StoB_REQ11_out & ~n2420;
  assign n2422 = ~n1461 & ~n2421;
  assign n2423 = sys_fair11done_out & ~n2422;
  assign n2424 = reg_controllable_BtoS_ACK11_out & ~n2322;
  assign n2425 = ~n1459 & ~n2424;
  assign n2426 = reg_i_StoB_REQ11_out & ~n2425;
  assign n2427 = ~n1462 & ~n2426;
  assign n2428 = ~sys_fair11done_out & ~n2427;
  assign n2429 = ~n2423 & ~n2428;
  assign n2430 = sys_fair12done_out & ~n2429;
  assign n2431 = ~n1464 & ~n2430;
  assign n2432 = ~reg_i_StoB_REQ12_out & ~n2431;
  assign n2433 = ~n2347 & ~n2432;
  assign n2434 = ~reg_i_StoB_REQ13_out & ~n2433;
  assign n2435 = ~n1539 & ~n2434;
  assign n2436 = sys_fair13done_out & ~n2435;
  assign n2437 = reg_controllable_BtoS_ACK13_out & ~n2331;
  assign n2438 = ~n1537 & ~n2437;
  assign n2439 = reg_i_StoB_REQ13_out & ~n2438;
  assign n2440 = ~n1540 & ~n2439;
  assign n2441 = ~sys_fair13done_out & ~n2440;
  assign n2442 = ~n2436 & ~n2441;
  assign n2443 = sys_fair0done_out & ~n2442;
  assign n2444 = ~n1542 & ~n2443;
  assign n2445 = ~reg_i_StoB_REQ0_out & ~n2444;
  assign n2446 = ~n2341 & ~n2445;
  assign n2447 = ~reg_i_StoB_REQ10_out & ~n2446;
  assign n2448 = ~n1969 & ~n2447;
  assign n2449 = sys_fair10done_out & ~n2448;
  assign n2450 = sys_fair0done_out & ~n2336;
  assign n2451 = ~n387 & ~n2450;
  assign n2452 = ~reg_i_StoB_REQ0_out & ~n2451;
  assign n2453 = ~n413 & ~n2452;
  assign n2454 = reg_controllable_BtoS_ACK10_out & ~n2453;
  assign n2455 = ~n1935 & ~n2454;
  assign n2456 = reg_i_StoB_REQ10_out & ~n2455;
  assign n2457 = ~n1970 & ~n2456;
  assign n2458 = ~sys_fair10done_out & ~n2457;
  assign n2459 = ~n2449 & ~n2458;
  assign n2460 = ~reg_i_StoB_REQ14_out & ~n2459;
  assign n2461 = ~n2266 & ~n2460;
  assign n2462 = sys_fair14done_out & ~n2461;
  assign n2463 = ~reg_i_StoB_REQ10_out & ~n2453;
  assign n2464 = ~n418 & ~n2463;
  assign n2465 = sys_fair10done_out & ~n2464;
  assign n2466 = ~sys_fair10done_out & ~n658;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = reg_controllable_BtoS_ACK14_out & ~n2467;
  assign n2469 = ~n1972 & ~n2468;
  assign n2470 = reg_i_StoB_REQ14_out & ~n2469;
  assign n2471 = ~n2267 & ~n2470;
  assign n2472 = ~sys_fair14done_out & ~n2471;
  assign n2473 = ~n2462 & ~n2472;
  assign n2474 = sys_fair15done_out & ~n2473;
  assign n2475 = reg_controllable_BtoS_ACK0_out & ~n2336;
  assign n2476 = ~n1578 & ~n2475;
  assign n2477 = reg_i_StoB_REQ0_out & ~n2476;
  assign n2478 = reg_controllable_BtoS_ACK12_out & ~n2327;
  assign n2479 = ~n1500 & ~n2478;
  assign n2480 = reg_i_StoB_REQ12_out & ~n2479;
  assign n2481 = reg_controllable_BtoS_ACK7_out & ~n2313;
  assign n2482 = ~n1386 & ~n2481;
  assign n2483 = reg_i_StoB_REQ7_out & ~n2482;
  assign n2484 = ~n1642 & ~n2354;
  assign n2485 = sys_fair1done_out & ~n2484;
  assign n2486 = ~n2361 & ~n2485;
  assign n2487 = ~reg_i_StoB_REQ3_out & ~n2486;
  assign n2488 = ~n2368 & ~n2487;
  assign n2489 = sys_fair3done_out & ~n2488;
  assign n2490 = ~n2370 & ~n2489;
  assign n2491 = ~reg_i_StoB_REQ4_out & ~n2490;
  assign n2492 = ~n2377 & ~n2491;
  assign n2493 = sys_fair4done_out & ~n2492;
  assign n2494 = ~n2379 & ~n2493;
  assign n2495 = ~reg_i_StoB_REQ5_out & ~n2494;
  assign n2496 = ~n2386 & ~n2495;
  assign n2497 = sys_fair5done_out & ~n2496;
  assign n2498 = ~n2388 & ~n2497;
  assign n2499 = ~reg_i_StoB_REQ8_out & ~n2498;
  assign n2500 = ~n2395 & ~n2499;
  assign n2501 = sys_fair8done_out & ~n2500;
  assign n2502 = ~n2397 & ~n2501;
  assign n2503 = ~reg_i_StoB_REQ6_out & ~n2502;
  assign n2504 = ~n2404 & ~n2503;
  assign n2505 = sys_fair6done_out & ~n2504;
  assign n2506 = ~n2406 & ~n2505;
  assign n2507 = sys_fair7done_out & ~n2506;
  assign n2508 = ~n1350 & ~n2507;
  assign n2509 = ~reg_i_StoB_REQ7_out & ~n2508;
  assign n2510 = ~n2483 & ~n2509;
  assign n2511 = ~reg_i_StoB_REQ9_out & ~n2510;
  assign n2512 = ~n2417 & ~n2511;
  assign n2513 = sys_fair9done_out & ~n2512;
  assign n2514 = ~n2419 & ~n2513;
  assign n2515 = ~reg_i_StoB_REQ11_out & ~n2514;
  assign n2516 = ~n2426 & ~n2515;
  assign n2517 = sys_fair11done_out & ~n2516;
  assign n2518 = ~n2428 & ~n2517;
  assign n2519 = sys_fair12done_out & ~n2518;
  assign n2520 = ~n1464 & ~n2519;
  assign n2521 = ~reg_i_StoB_REQ12_out & ~n2520;
  assign n2522 = ~n2480 & ~n2521;
  assign n2523 = ~reg_i_StoB_REQ13_out & ~n2522;
  assign n2524 = ~n2439 & ~n2523;
  assign n2525 = sys_fair13done_out & ~n2524;
  assign n2526 = ~n2441 & ~n2525;
  assign n2527 = sys_fair0done_out & ~n2526;
  assign n2528 = ~n1542 & ~n2527;
  assign n2529 = ~reg_i_StoB_REQ0_out & ~n2528;
  assign n2530 = ~n2477 & ~n2529;
  assign n2531 = ~reg_i_StoB_REQ10_out & ~n2530;
  assign n2532 = ~n2456 & ~n2531;
  assign n2533 = sys_fair10done_out & ~n2532;
  assign n2534 = ~n2458 & ~n2533;
  assign n2535 = ~reg_i_StoB_REQ14_out & ~n2534;
  assign n2536 = ~n2470 & ~n2535;
  assign n2537 = sys_fair14done_out & ~n2536;
  assign n2538 = ~n2472 & ~n2537;
  assign n2539 = reg_stateG12_out & ~n2538;
  assign n2540 = ~n2269 & ~n2539;
  assign n2541 = ~sys_fair15done_out & ~n2540;
  assign n2542 = ~n2474 & ~n2541;
  assign n2543 = fair_cnt<1>_out  & ~n2542;
  assign n2544 = ~n2274 & ~n2543;
  assign n2545 = fair_cnt<0>_out  & ~n2544;
  assign n2546 = ~n2277 & ~n2545;
  assign n2547 = env_fair1done_out & ~n2546;
  assign n2548 = ~n2280 & ~n2547;
  assign n2549 = ~env_fair0done_out & ~n2548;
  assign n2550 = ~n2282 & ~n2549;
  assign n2551 = reg_i_RtoB_ACK1_out & ~n2550;
  assign n2552 = reg_i_StoB_REQ2_out & ~n120;
  assign n2553 = ~n1133 & ~n2552;
  assign n2554 = ~sys_fair2done_out & ~n2553;
  assign n2555 = ~n1132 & ~n2554;
  assign n2556 = sys_fair1done_out & ~n2555;
  assign n2557 = ~reg_controllable_BtoS_ACK1_out & ~reg_controllable_BtoS_ACK2_out;
  assign n2558 = ~n1138 & ~n2557;
  assign n2559 = reg_i_StoB_REQ2_out & ~n2558;
  assign n2560 = ~reg_i_StoB_REQ2_out & ~reg_controllable_BtoS_ACK1_out;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = sys_fair2done_out & ~n2561;
  assign n2563 = ~n119 & ~n2557;
  assign n2564 = reg_i_StoB_REQ2_out & ~n2563;
  assign n2565 = reg_controllable_BtoS_ACK1_out & ~reg_controllable_BtoS_ACK2_out;
  assign n2566 = ~reg_controllable_BtoS_ACK2_out & ~n2565;
  assign n2567 = ~reg_i_StoB_REQ2_out & n2566;
  assign n2568 = ~n2564 & ~n2567;
  assign n2569 = ~sys_fair2done_out & ~n2568;
  assign n2570 = ~n2562 & ~n2569;
  assign n2571 = ~sys_fair1done_out & ~n2570;
  assign n2572 = ~n2556 & ~n2571;
  assign n2573 = ~reg_controllable_BtoS_ACK3_out & ~n2572;
  assign n2574 = ~n1130 & ~n2573;
  assign n2575 = reg_i_StoB_REQ3_out & ~n2574;
  assign n2576 = ~reg_i_StoB_REQ3_out & ~n2572;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = sys_fair3done_out & ~n2577;
  assign n2579 = ~sys_fair2done_out & ~n2554;
  assign n2580 = sys_fair1done_out & ~n2579;
  assign n2581 = ~n2571 & ~n2580;
  assign n2582 = ~reg_controllable_BtoS_ACK3_out & ~n2581;
  assign n2583 = ~n150 & ~n2582;
  assign n2584 = reg_i_StoB_REQ3_out & ~n2583;
  assign n2585 = ~n1177 & ~n2582;
  assign n2586 = ~reg_i_StoB_REQ3_out & ~n2585;
  assign n2587 = ~n2584 & ~n2586;
  assign n2588 = ~sys_fair3done_out & ~n2587;
  assign n2589 = ~n2578 & ~n2588;
  assign n2590 = ~reg_controllable_BtoS_ACK4_out & ~n2589;
  assign n2591 = ~n1129 & ~n2590;
  assign n2592 = reg_i_StoB_REQ4_out & ~n2591;
  assign n2593 = ~reg_i_StoB_REQ4_out & ~n2589;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = sys_fair4done_out & ~n2594;
  assign n2596 = ~n1159 & ~n2582;
  assign n2597 = reg_i_StoB_REQ3_out & ~n2596;
  assign n2598 = ~reg_i_StoB_REQ3_out & ~n2581;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = sys_fair3done_out & ~n2599;
  assign n2601 = ~n2588 & ~n2600;
  assign n2602 = ~reg_controllable_BtoS_ACK4_out & ~n2601;
  assign n2603 = ~n171 & ~n2602;
  assign n2604 = reg_i_StoB_REQ4_out & ~n2603;
  assign n2605 = ~n1210 & ~n2602;
  assign n2606 = ~reg_i_StoB_REQ4_out & ~n2605;
  assign n2607 = ~n2604 & ~n2606;
  assign n2608 = ~sys_fair4done_out & ~n2607;
  assign n2609 = ~n2595 & ~n2608;
  assign n2610 = ~reg_controllable_BtoS_ACK5_out & ~n2609;
  assign n2611 = ~n1128 & ~n2610;
  assign n2612 = reg_i_StoB_REQ5_out & ~n2611;
  assign n2613 = ~reg_i_StoB_REQ5_out & ~n2609;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = sys_fair5done_out & ~n2614;
  assign n2616 = ~n1193 & ~n2602;
  assign n2617 = reg_i_StoB_REQ4_out & ~n2616;
  assign n2618 = ~reg_i_StoB_REQ4_out & ~n2601;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = sys_fair4done_out & ~n2619;
  assign n2621 = ~n2608 & ~n2620;
  assign n2622 = ~reg_controllable_BtoS_ACK5_out & ~n2621;
  assign n2623 = ~n195 & ~n2622;
  assign n2624 = reg_i_StoB_REQ5_out & ~n2623;
  assign n2625 = ~n1246 & ~n2622;
  assign n2626 = ~reg_i_StoB_REQ5_out & ~n2625;
  assign n2627 = ~n2624 & ~n2626;
  assign n2628 = ~sys_fair5done_out & ~n2627;
  assign n2629 = ~n2615 & ~n2628;
  assign n2630 = ~reg_controllable_BtoS_ACK8_out & ~n2629;
  assign n2631 = ~n1127 & ~n2630;
  assign n2632 = reg_i_StoB_REQ8_out & ~n2631;
  assign n2633 = ~reg_i_StoB_REQ8_out & ~n2629;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = sys_fair8done_out & ~n2634;
  assign n2636 = ~n1229 & ~n2622;
  assign n2637 = reg_i_StoB_REQ5_out & ~n2636;
  assign n2638 = ~reg_i_StoB_REQ5_out & ~n2621;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = sys_fair5done_out & ~n2639;
  assign n2641 = ~n2628 & ~n2640;
  assign n2642 = ~reg_controllable_BtoS_ACK8_out & ~n2641;
  assign n2643 = ~n219 & ~n2642;
  assign n2644 = reg_i_StoB_REQ8_out & ~n2643;
  assign n2645 = ~n1282 & ~n2642;
  assign n2646 = ~reg_i_StoB_REQ8_out & ~n2645;
  assign n2647 = ~n2644 & ~n2646;
  assign n2648 = ~sys_fair8done_out & ~n2647;
  assign n2649 = ~n2635 & ~n2648;
  assign n2650 = ~reg_controllable_BtoS_ACK6_out & ~n2649;
  assign n2651 = ~n1126 & ~n2650;
  assign n2652 = reg_i_StoB_REQ6_out & ~n2651;
  assign n2653 = ~reg_i_StoB_REQ6_out & ~n2649;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = sys_fair6done_out & ~n2654;
  assign n2656 = ~n1265 & ~n2642;
  assign n2657 = reg_i_StoB_REQ8_out & ~n2656;
  assign n2658 = ~reg_i_StoB_REQ8_out & ~n2641;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = sys_fair8done_out & ~n2659;
  assign n2661 = ~n2648 & ~n2660;
  assign n2662 = ~reg_controllable_BtoS_ACK6_out & ~n2661;
  assign n2663 = ~n243 & ~n2662;
  assign n2664 = reg_i_StoB_REQ6_out & ~n2663;
  assign n2665 = ~n1318 & ~n2662;
  assign n2666 = ~reg_i_StoB_REQ6_out & ~n2665;
  assign n2667 = ~n2664 & ~n2666;
  assign n2668 = ~sys_fair6done_out & ~n2667;
  assign n2669 = ~n2655 & ~n2668;
  assign n2670 = sys_fair7done_out & ~n2669;
  assign n2671 = ~n1301 & ~n2662;
  assign n2672 = reg_i_StoB_REQ6_out & ~n2671;
  assign n2673 = ~reg_i_StoB_REQ6_out & ~n2661;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = sys_fair6done_out & ~n2674;
  assign n2676 = ~n2668 & ~n2675;
  assign n2677 = ~sys_fair7done_out & ~n2676;
  assign n2678 = ~n2670 & ~n2677;
  assign n2679 = ~reg_controllable_BtoS_ACK7_out & ~n2678;
  assign n2680 = ~n830 & ~n2679;
  assign n2681 = reg_i_StoB_REQ7_out & ~n2680;
  assign n2682 = ~n1350 & ~n2670;
  assign n2683 = reg_controllable_BtoS_ACK7_out & ~n2682;
  assign n2684 = ~n2679 & ~n2683;
  assign n2685 = ~reg_i_StoB_REQ7_out & ~n2684;
  assign n2686 = ~n2681 & ~n2685;
  assign n2687 = ~reg_controllable_BtoS_ACK9_out & ~n2686;
  assign n2688 = ~n1124 & ~n2687;
  assign n2689 = reg_i_StoB_REQ9_out & ~n2688;
  assign n2690 = ~reg_i_StoB_REQ9_out & ~n2686;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = sys_fair9done_out & ~n2691;
  assign n2693 = ~reg_controllable_BtoS_ACK7_out & ~n2676;
  assign n2694 = ~n845 & ~n2693;
  assign n2695 = reg_i_StoB_REQ7_out & ~n2694;
  assign n2696 = sys_fair7done_out & ~n2676;
  assign n2697 = ~n1350 & ~n2696;
  assign n2698 = reg_controllable_BtoS_ACK7_out & ~n2697;
  assign n2699 = ~n2693 & ~n2698;
  assign n2700 = ~reg_i_StoB_REQ7_out & ~n2699;
  assign n2701 = ~n2695 & ~n2700;
  assign n2702 = ~reg_controllable_BtoS_ACK9_out & ~n2701;
  assign n2703 = ~n291 & ~n2702;
  assign n2704 = reg_i_StoB_REQ9_out & ~n2703;
  assign n2705 = ~n1391 & ~n2702;
  assign n2706 = ~reg_i_StoB_REQ9_out & ~n2705;
  assign n2707 = ~n2704 & ~n2706;
  assign n2708 = ~sys_fair9done_out & ~n2707;
  assign n2709 = ~n2692 & ~n2708;
  assign n2710 = ~reg_controllable_BtoS_ACK11_out & ~n2709;
  assign n2711 = ~n1123 & ~n2710;
  assign n2712 = reg_i_StoB_REQ11_out & ~n2711;
  assign n2713 = ~reg_i_StoB_REQ11_out & ~n2709;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = sys_fair11done_out & ~n2714;
  assign n2716 = ~n1371 & ~n2702;
  assign n2717 = reg_i_StoB_REQ9_out & ~n2716;
  assign n2718 = ~reg_i_StoB_REQ9_out & ~n2701;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = sys_fair9done_out & ~n2719;
  assign n2721 = ~n2708 & ~n2720;
  assign n2722 = ~reg_controllable_BtoS_ACK11_out & ~n2721;
  assign n2723 = ~n319 & ~n2722;
  assign n2724 = reg_i_StoB_REQ11_out & ~n2723;
  assign n2725 = ~n1432 & ~n2722;
  assign n2726 = ~reg_i_StoB_REQ11_out & ~n2725;
  assign n2727 = ~n2724 & ~n2726;
  assign n2728 = ~sys_fair11done_out & ~n2727;
  assign n2729 = ~n2715 & ~n2728;
  assign n2730 = sys_fair12done_out & ~n2729;
  assign n2731 = ~n1415 & ~n2722;
  assign n2732 = reg_i_StoB_REQ11_out & ~n2731;
  assign n2733 = ~reg_i_StoB_REQ11_out & ~n2721;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = sys_fair11done_out & ~n2734;
  assign n2736 = ~n2728 & ~n2735;
  assign n2737 = ~sys_fair12done_out & ~n2736;
  assign n2738 = ~n2730 & ~n2737;
  assign n2739 = ~reg_controllable_BtoS_ACK12_out & ~n2738;
  assign n2740 = ~n886 & ~n2739;
  assign n2741 = reg_i_StoB_REQ12_out & ~n2740;
  assign n2742 = ~n1464 & ~n2730;
  assign n2743 = reg_controllable_BtoS_ACK12_out & ~n2742;
  assign n2744 = ~n2739 & ~n2743;
  assign n2745 = ~reg_i_StoB_REQ12_out & ~n2744;
  assign n2746 = ~n2741 & ~n2745;
  assign n2747 = ~reg_controllable_BtoS_ACK13_out & ~n2746;
  assign n2748 = ~n1121 & ~n2747;
  assign n2749 = reg_i_StoB_REQ13_out & ~n2748;
  assign n2750 = ~reg_i_StoB_REQ13_out & ~n2746;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = sys_fair13done_out & ~n2751;
  assign n2753 = ~reg_controllable_BtoS_ACK12_out & ~n2736;
  assign n2754 = ~n901 & ~n2753;
  assign n2755 = reg_i_StoB_REQ12_out & ~n2754;
  assign n2756 = sys_fair12done_out & ~n2736;
  assign n2757 = ~n1464 & ~n2756;
  assign n2758 = reg_controllable_BtoS_ACK12_out & ~n2757;
  assign n2759 = ~n2753 & ~n2758;
  assign n2760 = ~reg_i_StoB_REQ12_out & ~n2759;
  assign n2761 = ~n2755 & ~n2760;
  assign n2762 = ~reg_controllable_BtoS_ACK13_out & ~n2761;
  assign n2763 = ~n367 & ~n2762;
  assign n2764 = reg_i_StoB_REQ13_out & ~n2763;
  assign n2765 = ~n1505 & ~n2762;
  assign n2766 = ~reg_i_StoB_REQ13_out & ~n2765;
  assign n2767 = ~n2764 & ~n2766;
  assign n2768 = ~sys_fair13done_out & ~n2767;
  assign n2769 = ~n2752 & ~n2768;
  assign n2770 = sys_fair0done_out & ~n2769;
  assign n2771 = ~n1485 & ~n2762;
  assign n2772 = reg_i_StoB_REQ13_out & ~n2771;
  assign n2773 = ~reg_i_StoB_REQ13_out & ~n2761;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = sys_fair13done_out & ~n2774;
  assign n2776 = ~n2768 & ~n2775;
  assign n2777 = ~sys_fair0done_out & ~n2776;
  assign n2778 = ~n2770 & ~n2777;
  assign n2779 = ~reg_controllable_BtoS_ACK0_out & ~n2778;
  assign n2780 = ~n924 & ~n2779;
  assign n2781 = reg_i_StoB_REQ0_out & ~n2780;
  assign n2782 = ~n1542 & ~n2770;
  assign n2783 = reg_controllable_BtoS_ACK0_out & ~n2782;
  assign n2784 = ~n2779 & ~n2783;
  assign n2785 = ~reg_i_StoB_REQ0_out & ~n2784;
  assign n2786 = ~n2781 & ~n2785;
  assign n2787 = ~reg_controllable_BtoS_ACK10_out & ~n2786;
  assign n2788 = ~n1119 & ~n2787;
  assign n2789 = reg_i_StoB_REQ10_out & ~n2788;
  assign n2790 = ~reg_i_StoB_REQ10_out & ~n2786;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = sys_fair10done_out & ~n2791;
  assign n2793 = ~reg_controllable_BtoS_ACK0_out & ~n2776;
  assign n2794 = ~n1098 & ~n2793;
  assign n2795 = reg_i_StoB_REQ0_out & ~n2794;
  assign n2796 = sys_fair0done_out & ~n2776;
  assign n2797 = ~n1542 & ~n2796;
  assign n2798 = reg_controllable_BtoS_ACK0_out & ~n2797;
  assign n2799 = ~n2793 & ~n2798;
  assign n2800 = ~reg_i_StoB_REQ0_out & ~n2799;
  assign n2801 = ~n2795 & ~n2800;
  assign n2802 = ~reg_controllable_BtoS_ACK10_out & ~n2801;
  assign n2803 = ~n419 & ~n2802;
  assign n2804 = reg_i_StoB_REQ10_out & ~n2803;
  assign n2805 = ~n1583 & ~n2802;
  assign n2806 = ~reg_i_StoB_REQ10_out & ~n2805;
  assign n2807 = ~n2804 & ~n2806;
  assign n2808 = ~sys_fair10done_out & ~n2807;
  assign n2809 = ~n2792 & ~n2808;
  assign n2810 = ~reg_controllable_BtoS_ACK14_out & ~n2809;
  assign n2811 = ~n1998 & ~n2810;
  assign n2812 = reg_i_StoB_REQ14_out & ~n2811;
  assign n2813 = ~reg_i_StoB_REQ14_out & ~n2809;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = sys_fair14done_out & ~n2814;
  assign n2816 = ~n1563 & ~n2802;
  assign n2817 = reg_i_StoB_REQ10_out & ~n2816;
  assign n2818 = ~reg_i_StoB_REQ10_out & ~n2801;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = sys_fair10done_out & ~n2819;
  assign n2821 = ~n2808 & ~n2820;
  assign n2822 = ~reg_controllable_BtoS_ACK14_out & ~n2821;
  assign n2823 = ~n2264 & ~n2822;
  assign n2824 = reg_i_StoB_REQ14_out & ~n2823;
  assign n2825 = ~n2252 & ~n2822;
  assign n2826 = ~reg_i_StoB_REQ14_out & ~n2825;
  assign n2827 = ~n2824 & ~n2826;
  assign n2828 = ~sys_fair14done_out & ~n2827;
  assign n2829 = ~n2815 & ~n2828;
  assign n2830 = sys_fair15done_out & ~n2829;
  assign n2831 = ~sys_fair15done_out & ~n2268;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = fair_cnt<1>_out  & ~n2832;
  assign n2834 = ~n2274 & ~n2833;
  assign n2835 = ~fair_cnt<0>_out  & ~n2834;
  assign n2836 = ~n2276 & ~n2835;
  assign n2837 = env_fair1done_out & ~n2836;
  assign n2838 = ~env_fair1done_out & ~n2278;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = ~reg_i_RtoB_ACK1_out & ~n2839;
  assign n2841 = ~n2551 & ~n2840;
  assign n2842 = ~reg_i_RtoB_ACK0_out & ~n2841;
  assign n2843 = ~n1989 & ~n2842;
  assign n2844 = reg_nstateG7_1_out & ~n2843;
  assign n2845 = reg_nstateG7_1_out & ~n2844;
  assign n2846 = reg_stateG7_0_out & ~n2845;
  assign n2847 = ~reg_stateG7_0_out & ~n2843;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = ~reg_controllable_BtoR_REQ0_out & ~n2848;
  assign n2850 = ~reg_controllable_BtoR_REQ0_out & ~n2849;
  assign n2851 = reg_controllable_BtoR_REQ1_out & ~n2850;
  assign n2852 = env_fair0done_out & ~n701;
  assign n2853 = ~env_fair0done_out & ~n708;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = reg_i_RtoB_ACK1_out & ~n2854;
  assign n2856 = ~env_fair1done_out & ~n2546;
  assign n2857 = ~n2279 & ~n2856;
  assign n2858 = env_fair0done_out & ~n2857;
  assign n2859 = ~env_fair0done_out & ~n2268;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = ~reg_i_RtoB_ACK1_out & ~n2860;
  assign n2862 = ~n2855 & ~n2861;
  assign n2863 = reg_i_RtoB_ACK0_out & ~n2862;
  assign n2864 = reg_i_RtoB_ACK1_out & ~n1986;
  assign n2865 = env_fair0done_out & ~n2836;
  assign n2866 = ~env_fair0done_out & ~n2278;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = ~reg_i_RtoB_ACK1_out & ~n2867;
  assign n2869 = ~n2864 & ~n2868;
  assign n2870 = ~reg_i_RtoB_ACK0_out & ~n2869;
  assign n2871 = ~n2863 & ~n2870;
  assign n2872 = ~reg_nstateG7_1_out & ~n2871;
  assign n2873 = ~reg_nstateG7_1_out & ~n2872;
  assign n2874 = reg_stateG7_0_out & ~n2873;
  assign n2875 = ~reg_stateG7_0_out & ~n2871;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = reg_controllable_BtoR_REQ0_out & ~n2876;
  assign n2878 = ~n1601 & ~n1998;
  assign n2879 = reg_i_StoB_REQ14_out & ~n2878;
  assign n2880 = ~reg_i_StoB_REQ14_out & ~n1600;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = sys_fair14done_out & ~n2881;
  assign n2883 = ~n1932 & ~n2244;
  assign n2884 = reg_i_StoB_REQ14_out & ~n2883;
  assign n2885 = ~n1960 & ~n2252;
  assign n2886 = ~reg_i_StoB_REQ14_out & ~n2885;
  assign n2887 = ~n2884 & ~n2886;
  assign n2888 = ~sys_fair14done_out & ~n2887;
  assign n2889 = ~n2882 & ~n2888;
  assign n2890 = sys_fair15done_out & ~n2889;
  assign n2891 = ~n1960 & ~n2244;
  assign n2892 = reg_i_StoB_REQ14_out & ~n2891;
  assign n2893 = ~reg_i_StoB_REQ14_out & ~n1959;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = sys_fair14done_out & ~n2894;
  assign n2896 = ~n2888 & ~n2895;
  assign n2897 = reg_stateG12_out & ~n2896;
  assign n2898 = ~n2269 & ~n2897;
  assign n2899 = ~sys_fair15done_out & ~n2898;
  assign n2900 = ~n2890 & ~n2899;
  assign n2901 = fair_cnt<1>_out  & ~n2900;
  assign n2902 = ~n2274 & ~n2901;
  assign n2903 = fair_cnt<0>_out  & ~n2902;
  assign n2904 = ~n2277 & ~n2903;
  assign n2905 = reg_i_RtoB_ACK1_out & ~n2904;
  assign n2906 = env_fair1done_out & ~n2904;
  assign n2907 = ~n2856 & ~n2906;
  assign n2908 = ~reg_i_RtoB_ACK1_out & ~n2907;
  assign n2909 = ~n2905 & ~n2908;
  assign n2910 = reg_i_RtoB_ACK0_out & ~n2909;
  assign n2911 = fair_cnt<0>_out  & ~n2834;
  assign n2912 = ~n2277 & ~n2911;
  assign n2913 = ~env_fair1done_out & ~n2912;
  assign n2914 = ~n2837 & ~n2913;
  assign n2915 = ~reg_i_RtoB_ACK1_out & ~n2914;
  assign n2916 = ~n2905 & ~n2915;
  assign n2917 = ~reg_i_RtoB_ACK0_out & ~n2916;
  assign n2918 = ~n2910 & ~n2917;
  assign n2919 = reg_nstateG7_1_out & ~n2918;
  assign n2920 = reg_i_RtoB_ACK0_out & ~n2904;
  assign n2921 = env_fair0done_out & ~n2904;
  assign n2922 = ~env_fair0done_out & ~n2546;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = reg_i_RtoB_ACK1_out & ~n2923;
  assign n2925 = ~env_fair0done_out & ~n2912;
  assign n2926 = ~n2865 & ~n2925;
  assign n2927 = ~reg_i_RtoB_ACK1_out & ~n2926;
  assign n2928 = ~n2924 & ~n2927;
  assign n2929 = ~reg_i_RtoB_ACK0_out & ~n2928;
  assign n2930 = ~n2920 & ~n2929;
  assign n2931 = ~reg_nstateG7_1_out & ~n2930;
  assign n2932 = ~n2919 & ~n2931;
  assign n2933 = ~reg_controllable_BtoR_REQ0_out & ~n2932;
  assign n2934 = ~n2877 & ~n2933;
  assign n2935 = ~reg_controllable_BtoR_REQ1_out & ~n2934;
  assign n2936 = ~n2851 & ~n2935;
  assign n2937 = reg_controllable_ENQ_out & ~n2936;
  assign n2938 = env_fair0done_out & ~n710;
  assign n2939 = ~reg_controllable_BtoS_ACK14_out & ~n2467;
  assign n2940 = ~reg_controllable_BtoS_ACK14_out & ~n2939;
  assign n2941 = reg_i_StoB_REQ14_out & ~n2940;
  assign n2942 = ~reg_controllable_BtoS_ACK10_out & ~n2453;
  assign n2943 = ~reg_controllable_BtoS_ACK10_out & ~n2942;
  assign n2944 = reg_i_StoB_REQ10_out & ~n2943;
  assign n2945 = ~reg_controllable_BtoS_ACK0_out & ~n2451;
  assign n2946 = ~reg_controllable_BtoS_ACK0_out & ~n2945;
  assign n2947 = reg_i_StoB_REQ0_out & ~n2946;
  assign n2948 = ~reg_controllable_BtoS_ACK13_out & ~n2331;
  assign n2949 = ~reg_controllable_BtoS_ACK13_out & ~n2948;
  assign n2950 = reg_i_StoB_REQ13_out & ~n2949;
  assign n2951 = ~reg_controllable_BtoS_ACK12_out & ~n2329;
  assign n2952 = ~reg_controllable_BtoS_ACK12_out & ~n2951;
  assign n2953 = reg_i_StoB_REQ12_out & ~n2952;
  assign n2954 = ~reg_controllable_BtoS_ACK11_out & ~n2322;
  assign n2955 = ~reg_controllable_BtoS_ACK11_out & ~n2954;
  assign n2956 = reg_i_StoB_REQ11_out & ~n2955;
  assign n2957 = ~reg_controllable_BtoS_ACK9_out & ~n2317;
  assign n2958 = ~reg_controllable_BtoS_ACK9_out & ~n2957;
  assign n2959 = reg_i_StoB_REQ9_out & ~n2958;
  assign n2960 = ~reg_controllable_BtoS_ACK7_out & ~n2315;
  assign n2961 = ~reg_controllable_BtoS_ACK7_out & ~n2960;
  assign n2962 = reg_i_StoB_REQ7_out & ~n2961;
  assign n2963 = ~reg_controllable_BtoS_ACK6_out & ~n2308;
  assign n2964 = ~reg_controllable_BtoS_ACK6_out & ~n2963;
  assign n2965 = reg_i_StoB_REQ6_out & ~n2964;
  assign n2966 = ~reg_controllable_BtoS_ACK8_out & ~n2303;
  assign n2967 = ~reg_controllable_BtoS_ACK8_out & ~n2966;
  assign n2968 = reg_i_StoB_REQ8_out & ~n2967;
  assign n2969 = ~reg_controllable_BtoS_ACK5_out & ~n2298;
  assign n2970 = ~reg_controllable_BtoS_ACK5_out & ~n2969;
  assign n2971 = reg_i_StoB_REQ5_out & ~n2970;
  assign n2972 = ~reg_controllable_BtoS_ACK4_out & ~n2293;
  assign n2973 = ~reg_controllable_BtoS_ACK4_out & ~n2972;
  assign n2974 = reg_i_StoB_REQ4_out & ~n2973;
  assign n2975 = ~reg_controllable_BtoS_ACK3_out & ~n2288;
  assign n2976 = ~reg_controllable_BtoS_ACK3_out & ~n2975;
  assign n2977 = reg_i_StoB_REQ3_out & ~n2976;
  assign n2978 = ~reg_controllable_BtoS_ACK2_out & ~n439;
  assign n2979 = ~reg_controllable_BtoS_ACK2_out & ~n2978;
  assign n2980 = reg_i_StoB_REQ2_out & ~n2979;
  assign n2981 = reg_i_StoB_REQ2_out & ~n2980;
  assign n2982 = sys_fair2done_out & ~n2981;
  assign n2983 = ~n452 & ~n2982;
  assign n2984 = sys_fair1done_out & ~n2983;
  assign n2985 = ~sys_fair1done_out & ~n441;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = ~reg_i_StoB_REQ3_out & ~n2986;
  assign n2988 = ~n2977 & ~n2987;
  assign n2989 = sys_fair3done_out & ~n2988;
  assign n2990 = ~sys_fair3done_out & ~n473;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = ~reg_i_StoB_REQ4_out & ~n2991;
  assign n2993 = ~n2974 & ~n2992;
  assign n2994 = sys_fair4done_out & ~n2993;
  assign n2995 = ~sys_fair4done_out & ~n489;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = ~reg_i_StoB_REQ5_out & ~n2996;
  assign n2998 = ~n2971 & ~n2997;
  assign n2999 = sys_fair5done_out & ~n2998;
  assign n3000 = ~sys_fair5done_out & ~n505;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = ~reg_i_StoB_REQ8_out & ~n3001;
  assign n3003 = ~n2968 & ~n3002;
  assign n3004 = sys_fair8done_out & ~n3003;
  assign n3005 = ~sys_fair8done_out & ~n521;
  assign n3006 = ~n3004 & ~n3005;
  assign n3007 = ~reg_i_StoB_REQ6_out & ~n3006;
  assign n3008 = ~n2965 & ~n3007;
  assign n3009 = sys_fair6done_out & ~n3008;
  assign n3010 = ~sys_fair6done_out & ~n535;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = sys_fair7done_out & ~n3011;
  assign n3013 = ~n536 & ~n3012;
  assign n3014 = ~reg_i_StoB_REQ7_out & ~n3013;
  assign n3015 = ~n2962 & ~n3014;
  assign n3016 = ~reg_i_StoB_REQ9_out & ~n3015;
  assign n3017 = ~n2959 & ~n3016;
  assign n3018 = sys_fair9done_out & ~n3017;
  assign n3019 = ~sys_fair9done_out & ~n572;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = ~reg_i_StoB_REQ11_out & ~n3020;
  assign n3022 = ~n2956 & ~n3021;
  assign n3023 = sys_fair11done_out & ~n3022;
  assign n3024 = ~sys_fair11done_out & ~n586;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = sys_fair12done_out & ~n3025;
  assign n3027 = ~n587 & ~n3026;
  assign n3028 = ~reg_i_StoB_REQ12_out & ~n3027;
  assign n3029 = ~n2953 & ~n3028;
  assign n3030 = ~reg_i_StoB_REQ13_out & ~n3029;
  assign n3031 = ~n2950 & ~n3030;
  assign n3032 = sys_fair13done_out & ~n3031;
  assign n3033 = ~sys_fair13done_out & ~n621;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = sys_fair0done_out & ~n3034;
  assign n3036 = ~n622 & ~n3035;
  assign n3037 = ~reg_i_StoB_REQ0_out & ~n3036;
  assign n3038 = ~n2947 & ~n3037;
  assign n3039 = ~reg_i_StoB_REQ10_out & ~n3038;
  assign n3040 = ~n2944 & ~n3039;
  assign n3041 = sys_fair10done_out & ~n3040;
  assign n3042 = ~sys_fair10done_out & ~n663;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = ~reg_i_StoB_REQ14_out & ~n3043;
  assign n3045 = ~n2941 & ~n3044;
  assign n3046 = sys_fair14done_out & ~n3045;
  assign n3047 = ~sys_fair14done_out & ~n691;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = reg_stateG12_out & ~n3048;
  assign n3050 = ~n692 & ~n3049;
  assign n3051 = ~sys_fair15done_out & ~n3050;
  assign n3052 = ~n677 & ~n3051;
  assign n3053 = fair_cnt<1>_out  & ~n3052;
  assign n3054 = ~n697 & ~n3053;
  assign n3055 = fair_cnt<0>_out  & ~n3054;
  assign n3056 = ~n700 & ~n3055;
  assign n3057 = env_fair1done_out & ~n3056;
  assign n3058 = ~n709 & ~n3057;
  assign n3059 = ~env_fair0done_out & ~n3058;
  assign n3060 = ~n2938 & ~n3059;
  assign n3061 = reg_i_RtoB_ACK1_out & ~n3060;
  assign n3062 = ~n1987 & ~n3061;
  assign n3063 = ~reg_i_RtoB_ACK0_out & ~n3062;
  assign n3064 = ~reg_i_RtoB_ACK0_out & ~n3063;
  assign n3065 = reg_nstateG7_1_out & ~n3064;
  assign n3066 = reg_nstateG7_1_out & ~n3065;
  assign n3067 = reg_stateG7_0_out & ~n3066;
  assign n3068 = ~reg_stateG7_0_out & ~n3064;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = ~reg_controllable_BtoR_REQ0_out & ~n3069;
  assign n3071 = ~reg_controllable_BtoR_REQ0_out & ~n3070;
  assign n3072 = reg_controllable_BtoR_REQ1_out & ~n3071;
  assign n3073 = ~env_fair1done_out & ~n3056;
  assign n3074 = ~n702 & ~n3073;
  assign n3075 = env_fair0done_out & ~n3074;
  assign n3076 = ~n2853 & ~n3075;
  assign n3077 = ~reg_i_RtoB_ACK1_out & ~n3076;
  assign n3078 = ~reg_i_RtoB_ACK1_out & ~n3077;
  assign n3079 = reg_i_RtoB_ACK0_out & ~n3078;
  assign n3080 = ~reg_i_RtoB_ACK1_out & ~n1987;
  assign n3081 = ~reg_i_RtoB_ACK0_out & ~n3080;
  assign n3082 = ~n3079 & ~n3081;
  assign n3083 = ~reg_nstateG7_1_out & ~n3082;
  assign n3084 = ~reg_nstateG7_1_out & ~n3083;
  assign n3085 = reg_stateG7_0_out & ~n3084;
  assign n3086 = ~reg_stateG7_0_out & ~n3082;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = reg_controllable_BtoR_REQ0_out & ~n3087;
  assign n3089 = ~reg_i_RtoB_ACK1_out & ~n2908;
  assign n3090 = ~reg_i_RtoB_ACK0_out & ~n3089;
  assign n3091 = ~reg_i_RtoB_ACK0_out & ~n3090;
  assign n3092 = reg_nstateG7_1_out & ~n3091;
  assign n3093 = ~reg_i_RtoB_ACK1_out & ~n2923;
  assign n3094 = ~reg_i_RtoB_ACK1_out & ~n3093;
  assign n3095 = ~reg_i_RtoB_ACK0_out & ~n3094;
  assign n3096 = ~reg_i_RtoB_ACK0_out & ~n3095;
  assign n3097 = ~reg_nstateG7_1_out & ~n3096;
  assign n3098 = ~n3092 & ~n3097;
  assign n3099 = ~reg_controllable_BtoR_REQ0_out & ~n3098;
  assign n3100 = ~n3088 & ~n3099;
  assign n3101 = ~reg_controllable_BtoR_REQ1_out & ~n3100;
  assign n3102 = ~n3072 & ~n3101;
  assign n3103 = ~reg_controllable_ENQ_out & ~n3102;
  assign n3104 = ~n2937 & ~n3103;
  assign n3105 = reg_controllable_DEQ_out & ~n3104;
  assign n3106 = sys_fair15done_out & ~n691;
  assign n3107 = ~n3051 & ~n3106;
  assign n3108 = fair_cnt<1>_out  & ~n3107;
  assign n3109 = ~n697 & ~n3108;
  assign n3110 = ~fair_cnt<0>_out  & ~n3109;
  assign n3111 = ~n699 & ~n3110;
  assign n3112 = env_fair1done_out & ~n3111;
  assign n3113 = ~env_fair1done_out & ~n701;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = reg_i_RtoB_ACK1_out & ~n3114;
  assign n3116 = sys_fair15done_out & ~n1976;
  assign n3117 = ~sys_fair2done_out & ~n2284;
  assign n3118 = sys_fair1done_out & ~n3117;
  assign n3119 = ~n2287 & ~n3118;
  assign n3120 = ~reg_controllable_BtoS_ACK3_out & ~n3119;
  assign n3121 = ~reg_controllable_BtoS_ACK3_out & ~n3120;
  assign n3122 = reg_i_StoB_REQ3_out & ~n3121;
  assign n3123 = ~reg_i_StoB_REQ3_out & ~n3119;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = sys_fair3done_out & ~n3124;
  assign n3126 = ~n2292 & ~n3125;
  assign n3127 = ~reg_controllable_BtoS_ACK4_out & ~n3126;
  assign n3128 = ~reg_controllable_BtoS_ACK4_out & ~n3127;
  assign n3129 = reg_i_StoB_REQ4_out & ~n3128;
  assign n3130 = ~reg_i_StoB_REQ4_out & ~n3126;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = sys_fair4done_out & ~n3131;
  assign n3133 = ~n2297 & ~n3132;
  assign n3134 = ~reg_controllable_BtoS_ACK5_out & ~n3133;
  assign n3135 = ~reg_controllable_BtoS_ACK5_out & ~n3134;
  assign n3136 = reg_i_StoB_REQ5_out & ~n3135;
  assign n3137 = ~reg_i_StoB_REQ5_out & ~n3133;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = sys_fair5done_out & ~n3138;
  assign n3140 = ~n2302 & ~n3139;
  assign n3141 = ~reg_controllable_BtoS_ACK8_out & ~n3140;
  assign n3142 = ~reg_controllable_BtoS_ACK8_out & ~n3141;
  assign n3143 = reg_i_StoB_REQ8_out & ~n3142;
  assign n3144 = ~reg_i_StoB_REQ8_out & ~n3140;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = sys_fair8done_out & ~n3145;
  assign n3147 = ~n2307 & ~n3146;
  assign n3148 = ~reg_controllable_BtoS_ACK6_out & ~n3147;
  assign n3149 = ~reg_controllable_BtoS_ACK6_out & ~n3148;
  assign n3150 = reg_i_StoB_REQ6_out & ~n3149;
  assign n3151 = ~reg_i_StoB_REQ6_out & ~n3147;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = sys_fair6done_out & ~n3152;
  assign n3154 = ~n2312 & ~n3153;
  assign n3155 = sys_fair7done_out & ~n3154;
  assign n3156 = ~n259 & ~n3155;
  assign n3157 = ~reg_controllable_BtoS_ACK7_out & ~n3156;
  assign n3158 = ~reg_controllable_BtoS_ACK7_out & ~n3157;
  assign n3159 = reg_i_StoB_REQ7_out & ~n3158;
  assign n3160 = ~reg_i_StoB_REQ7_out & ~n3156;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = ~reg_controllable_BtoS_ACK9_out & ~n3161;
  assign n3163 = ~reg_controllable_BtoS_ACK9_out & ~n3162;
  assign n3164 = reg_i_StoB_REQ9_out & ~n3163;
  assign n3165 = ~reg_i_StoB_REQ9_out & ~n3161;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = sys_fair9done_out & ~n3166;
  assign n3168 = ~n2321 & ~n3167;
  assign n3169 = ~reg_controllable_BtoS_ACK11_out & ~n3168;
  assign n3170 = ~reg_controllable_BtoS_ACK11_out & ~n3169;
  assign n3171 = reg_i_StoB_REQ11_out & ~n3170;
  assign n3172 = ~reg_i_StoB_REQ11_out & ~n3168;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = sys_fair11done_out & ~n3173;
  assign n3175 = ~n2326 & ~n3174;
  assign n3176 = sys_fair12done_out & ~n3175;
  assign n3177 = ~n335 & ~n3176;
  assign n3178 = ~reg_controllable_BtoS_ACK12_out & ~n3177;
  assign n3179 = ~reg_controllable_BtoS_ACK12_out & ~n3178;
  assign n3180 = reg_i_StoB_REQ12_out & ~n3179;
  assign n3181 = ~reg_i_StoB_REQ12_out & ~n3177;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = ~reg_controllable_BtoS_ACK13_out & ~n3182;
  assign n3184 = ~reg_controllable_BtoS_ACK13_out & ~n3183;
  assign n3185 = reg_i_StoB_REQ13_out & ~n3184;
  assign n3186 = ~reg_i_StoB_REQ13_out & ~n3182;
  assign n3187 = ~n3185 & ~n3186;
  assign n3188 = sys_fair13done_out & ~n3187;
  assign n3189 = ~n2335 & ~n3188;
  assign n3190 = sys_fair0done_out & ~n3189;
  assign n3191 = ~n387 & ~n3190;
  assign n3192 = ~reg_controllable_BtoS_ACK0_out & ~n3191;
  assign n3193 = ~reg_controllable_BtoS_ACK0_out & ~n3192;
  assign n3194 = reg_i_StoB_REQ0_out & ~n3193;
  assign n3195 = ~reg_i_StoB_REQ0_out & ~n3191;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = ~reg_controllable_BtoS_ACK10_out & ~n3196;
  assign n3198 = ~reg_controllable_BtoS_ACK10_out & ~n3197;
  assign n3199 = reg_i_StoB_REQ10_out & ~n3198;
  assign n3200 = ~sys_fair2done_out & ~n452;
  assign n3201 = sys_fair1done_out & ~n3200;
  assign n3202 = ~n2985 & ~n3201;
  assign n3203 = ~reg_i_StoB_REQ3_out & ~n3202;
  assign n3204 = ~n3122 & ~n3203;
  assign n3205 = sys_fair3done_out & ~n3204;
  assign n3206 = ~n2990 & ~n3205;
  assign n3207 = ~reg_i_StoB_REQ4_out & ~n3206;
  assign n3208 = ~n3129 & ~n3207;
  assign n3209 = sys_fair4done_out & ~n3208;
  assign n3210 = ~n2995 & ~n3209;
  assign n3211 = ~reg_i_StoB_REQ5_out & ~n3210;
  assign n3212 = ~n3136 & ~n3211;
  assign n3213 = sys_fair5done_out & ~n3212;
  assign n3214 = ~n3000 & ~n3213;
  assign n3215 = ~reg_i_StoB_REQ8_out & ~n3214;
  assign n3216 = ~n3143 & ~n3215;
  assign n3217 = sys_fair8done_out & ~n3216;
  assign n3218 = ~n3005 & ~n3217;
  assign n3219 = ~reg_i_StoB_REQ6_out & ~n3218;
  assign n3220 = ~n3150 & ~n3219;
  assign n3221 = sys_fair6done_out & ~n3220;
  assign n3222 = ~n3010 & ~n3221;
  assign n3223 = sys_fair7done_out & ~n3222;
  assign n3224 = ~n536 & ~n3223;
  assign n3225 = ~reg_i_StoB_REQ7_out & ~n3224;
  assign n3226 = ~n3159 & ~n3225;
  assign n3227 = ~reg_i_StoB_REQ9_out & ~n3226;
  assign n3228 = ~n3164 & ~n3227;
  assign n3229 = sys_fair9done_out & ~n3228;
  assign n3230 = ~n3019 & ~n3229;
  assign n3231 = ~reg_i_StoB_REQ11_out & ~n3230;
  assign n3232 = ~n3171 & ~n3231;
  assign n3233 = sys_fair11done_out & ~n3232;
  assign n3234 = ~n3024 & ~n3233;
  assign n3235 = sys_fair12done_out & ~n3234;
  assign n3236 = ~n587 & ~n3235;
  assign n3237 = ~reg_i_StoB_REQ12_out & ~n3236;
  assign n3238 = ~n3180 & ~n3237;
  assign n3239 = ~reg_i_StoB_REQ13_out & ~n3238;
  assign n3240 = ~n3185 & ~n3239;
  assign n3241 = sys_fair13done_out & ~n3240;
  assign n3242 = ~n3033 & ~n3241;
  assign n3243 = sys_fair0done_out & ~n3242;
  assign n3244 = ~n622 & ~n3243;
  assign n3245 = ~reg_i_StoB_REQ0_out & ~n3244;
  assign n3246 = ~n3194 & ~n3245;
  assign n3247 = ~reg_i_StoB_REQ10_out & ~n3246;
  assign n3248 = ~n3199 & ~n3247;
  assign n3249 = sys_fair10done_out & ~n3248;
  assign n3250 = ~n3042 & ~n3249;
  assign n3251 = reg_controllable_BtoS_ACK14_out & ~n3250;
  assign n3252 = reg_controllable_BtoS_ACK10_out & ~n3196;
  assign n3253 = reg_controllable_BtoS_ACK0_out & ~n3191;
  assign n3254 = reg_controllable_BtoS_ACK13_out & ~n3182;
  assign n3255 = reg_controllable_BtoS_ACK12_out & ~n3177;
  assign n3256 = reg_controllable_BtoS_ACK11_out & ~n3168;
  assign n3257 = reg_controllable_BtoS_ACK9_out & ~n3161;
  assign n3258 = reg_controllable_BtoS_ACK7_out & ~n3156;
  assign n3259 = reg_controllable_BtoS_ACK6_out & ~n3147;
  assign n3260 = reg_controllable_BtoS_ACK8_out & ~n3140;
  assign n3261 = reg_controllable_BtoS_ACK5_out & ~n3133;
  assign n3262 = reg_controllable_BtoS_ACK4_out & ~n3126;
  assign n3263 = reg_controllable_BtoS_ACK3_out & ~n3119;
  assign n3264 = ~sys_fair2done_out & ~n2359;
  assign n3265 = sys_fair1done_out & ~n3264;
  assign n3266 = ~sys_fair1done_out & n1131;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = ~reg_controllable_BtoS_ACK3_out & ~n3267;
  assign n3269 = ~n3263 & ~n3268;
  assign n3270 = reg_i_StoB_REQ3_out & ~n3269;
  assign n3271 = ~reg_i_StoB_REQ3_out & ~n3267;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = sys_fair3done_out & ~n3272;
  assign n3274 = ~sys_fair3done_out & ~n1209;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = ~reg_controllable_BtoS_ACK4_out & ~n3275;
  assign n3277 = ~n3262 & ~n3276;
  assign n3278 = reg_i_StoB_REQ4_out & ~n3277;
  assign n3279 = ~reg_i_StoB_REQ4_out & ~n3275;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = sys_fair4done_out & ~n3280;
  assign n3282 = ~sys_fair4done_out & ~n1245;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~reg_controllable_BtoS_ACK5_out & ~n3283;
  assign n3285 = ~n3261 & ~n3284;
  assign n3286 = reg_i_StoB_REQ5_out & ~n3285;
  assign n3287 = ~reg_i_StoB_REQ5_out & ~n3283;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = sys_fair5done_out & ~n3288;
  assign n3290 = ~sys_fair5done_out & ~n1281;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = ~reg_controllable_BtoS_ACK8_out & ~n3291;
  assign n3293 = ~n3260 & ~n3292;
  assign n3294 = reg_i_StoB_REQ8_out & ~n3293;
  assign n3295 = ~reg_i_StoB_REQ8_out & ~n3291;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = sys_fair8done_out & ~n3296;
  assign n3298 = ~sys_fair8done_out & ~n1317;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~reg_controllable_BtoS_ACK6_out & ~n3299;
  assign n3301 = ~n3259 & ~n3300;
  assign n3302 = reg_i_StoB_REQ6_out & ~n3301;
  assign n3303 = ~reg_i_StoB_REQ6_out & ~n3299;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = sys_fair6done_out & ~n3304;
  assign n3306 = ~sys_fair6done_out & ~n1349;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = sys_fair7done_out & ~n3307;
  assign n3309 = ~n1350 & ~n3308;
  assign n3310 = ~reg_controllable_BtoS_ACK7_out & ~n3309;
  assign n3311 = ~n3258 & ~n3310;
  assign n3312 = reg_i_StoB_REQ7_out & ~n3311;
  assign n3313 = ~reg_i_StoB_REQ7_out & ~n3309;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~reg_controllable_BtoS_ACK9_out & ~n3314;
  assign n3316 = ~n3257 & ~n3315;
  assign n3317 = reg_i_StoB_REQ9_out & ~n3316;
  assign n3318 = ~reg_i_StoB_REQ9_out & ~n3314;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = sys_fair9done_out & ~n3319;
  assign n3321 = ~sys_fair9done_out & ~n1431;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = ~reg_controllable_BtoS_ACK11_out & ~n3322;
  assign n3324 = ~n3256 & ~n3323;
  assign n3325 = reg_i_StoB_REQ11_out & ~n3324;
  assign n3326 = ~reg_i_StoB_REQ11_out & ~n3322;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = sys_fair11done_out & ~n3327;
  assign n3329 = ~sys_fair11done_out & ~n1463;
  assign n3330 = ~n3328 & ~n3329;
  assign n3331 = sys_fair12done_out & ~n3330;
  assign n3332 = ~n1464 & ~n3331;
  assign n3333 = ~reg_controllable_BtoS_ACK12_out & ~n3332;
  assign n3334 = ~n3255 & ~n3333;
  assign n3335 = reg_i_StoB_REQ12_out & ~n3334;
  assign n3336 = ~reg_i_StoB_REQ12_out & ~n3332;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = ~reg_controllable_BtoS_ACK13_out & ~n3337;
  assign n3339 = ~n3254 & ~n3338;
  assign n3340 = reg_i_StoB_REQ13_out & ~n3339;
  assign n3341 = ~reg_i_StoB_REQ13_out & ~n3337;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = sys_fair13done_out & ~n3342;
  assign n3344 = ~sys_fair13done_out & ~n1541;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = sys_fair0done_out & ~n3345;
  assign n3347 = ~n1542 & ~n3346;
  assign n3348 = ~reg_controllable_BtoS_ACK0_out & ~n3347;
  assign n3349 = ~n3253 & ~n3348;
  assign n3350 = reg_i_StoB_REQ0_out & ~n3349;
  assign n3351 = ~reg_i_StoB_REQ0_out & ~n3347;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = ~reg_controllable_BtoS_ACK10_out & ~n3352;
  assign n3354 = ~n3252 & ~n3353;
  assign n3355 = reg_i_StoB_REQ10_out & ~n3354;
  assign n3356 = ~reg_i_StoB_REQ10_out & ~n3352;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = sys_fair10done_out & ~n3357;
  assign n3359 = ~sys_fair10done_out & ~n1971;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~reg_controllable_BtoS_ACK14_out & ~n3360;
  assign n3362 = ~n3251 & ~n3361;
  assign n3363 = reg_i_StoB_REQ14_out & ~n3362;
  assign n3364 = reg_controllable_BtoS_ACK10_out & ~n3246;
  assign n3365 = ~n3353 & ~n3364;
  assign n3366 = reg_i_StoB_REQ10_out & ~n3365;
  assign n3367 = reg_controllable_BtoS_ACK0_out & ~n3244;
  assign n3368 = ~n3348 & ~n3367;
  assign n3369 = reg_i_StoB_REQ0_out & ~n3368;
  assign n3370 = reg_controllable_BtoS_ACK13_out & ~n3238;
  assign n3371 = ~n3338 & ~n3370;
  assign n3372 = reg_i_StoB_REQ13_out & ~n3371;
  assign n3373 = reg_controllable_BtoS_ACK12_out & ~n3236;
  assign n3374 = ~n3333 & ~n3373;
  assign n3375 = reg_i_StoB_REQ12_out & ~n3374;
  assign n3376 = reg_controllable_BtoS_ACK11_out & ~n3230;
  assign n3377 = ~n3323 & ~n3376;
  assign n3378 = reg_i_StoB_REQ11_out & ~n3377;
  assign n3379 = reg_controllable_BtoS_ACK9_out & ~n3226;
  assign n3380 = ~n3315 & ~n3379;
  assign n3381 = reg_i_StoB_REQ9_out & ~n3380;
  assign n3382 = reg_controllable_BtoS_ACK7_out & ~n3224;
  assign n3383 = ~n3310 & ~n3382;
  assign n3384 = reg_i_StoB_REQ7_out & ~n3383;
  assign n3385 = reg_controllable_BtoS_ACK6_out & ~n3218;
  assign n3386 = ~n3300 & ~n3385;
  assign n3387 = reg_i_StoB_REQ6_out & ~n3386;
  assign n3388 = reg_controllable_BtoS_ACK8_out & ~n3214;
  assign n3389 = ~n3292 & ~n3388;
  assign n3390 = reg_i_StoB_REQ8_out & ~n3389;
  assign n3391 = reg_controllable_BtoS_ACK5_out & ~n3210;
  assign n3392 = ~n3284 & ~n3391;
  assign n3393 = reg_i_StoB_REQ5_out & ~n3392;
  assign n3394 = reg_controllable_BtoS_ACK4_out & ~n3206;
  assign n3395 = ~n3276 & ~n3394;
  assign n3396 = reg_i_StoB_REQ4_out & ~n3395;
  assign n3397 = reg_controllable_BtoS_ACK3_out & ~n3202;
  assign n3398 = ~n3268 & ~n3397;
  assign n3399 = reg_i_StoB_REQ3_out & ~n3398;
  assign n3400 = ~sys_fair2done_out & ~n1641;
  assign n3401 = ~sys_fair2done_out & ~n3400;
  assign n3402 = sys_fair1done_out & ~n3401;
  assign n3403 = ~sys_fair1done_out & ~n1641;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = ~reg_i_StoB_REQ3_out & ~n3404;
  assign n3406 = ~n3399 & ~n3405;
  assign n3407 = sys_fair3done_out & ~n3406;
  assign n3408 = ~sys_fair3done_out & ~n1667;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~reg_i_StoB_REQ4_out & ~n3409;
  assign n3411 = ~n3396 & ~n3410;
  assign n3412 = sys_fair4done_out & ~n3411;
  assign n3413 = ~sys_fair4done_out & ~n1689;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~reg_i_StoB_REQ5_out & ~n3414;
  assign n3416 = ~n3393 & ~n3415;
  assign n3417 = sys_fair5done_out & ~n3416;
  assign n3418 = ~sys_fair5done_out & ~n1712;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = ~reg_i_StoB_REQ8_out & ~n3419;
  assign n3421 = ~n3390 & ~n3420;
  assign n3422 = sys_fair8done_out & ~n3421;
  assign n3423 = ~sys_fair8done_out & ~n1735;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~reg_i_StoB_REQ6_out & ~n3424;
  assign n3426 = ~n3387 & ~n3425;
  assign n3427 = sys_fair6done_out & ~n3426;
  assign n3428 = ~sys_fair6done_out & ~n1753;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = sys_fair7done_out & ~n3429;
  assign n3431 = ~n1754 & ~n3430;
  assign n3432 = ~reg_i_StoB_REQ7_out & ~n3431;
  assign n3433 = ~n3384 & ~n3432;
  assign n3434 = ~reg_i_StoB_REQ9_out & ~n3433;
  assign n3435 = ~n3381 & ~n3434;
  assign n3436 = sys_fair9done_out & ~n3435;
  assign n3437 = ~sys_fair9done_out & ~n1806;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = ~reg_i_StoB_REQ11_out & ~n3438;
  assign n3440 = ~n3378 & ~n3439;
  assign n3441 = sys_fair11done_out & ~n3440;
  assign n3442 = ~sys_fair11done_out & ~n1824;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = sys_fair12done_out & ~n3443;
  assign n3445 = ~n1825 & ~n3444;
  assign n3446 = ~reg_i_StoB_REQ12_out & ~n3445;
  assign n3447 = ~n3375 & ~n3446;
  assign n3448 = ~reg_i_StoB_REQ13_out & ~n3447;
  assign n3449 = ~n3372 & ~n3448;
  assign n3450 = sys_fair13done_out & ~n3449;
  assign n3451 = ~sys_fair13done_out & ~n1872;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = sys_fair0done_out & ~n3452;
  assign n3454 = ~n1873 & ~n3453;
  assign n3455 = ~reg_i_StoB_REQ0_out & ~n3454;
  assign n3456 = ~n3369 & ~n3455;
  assign n3457 = ~reg_i_StoB_REQ10_out & ~n3456;
  assign n3458 = ~n3366 & ~n3457;
  assign n3459 = sys_fair10done_out & ~n3458;
  assign n3460 = ~sys_fair10done_out & ~n1939;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = ~reg_i_StoB_REQ14_out & ~n3461;
  assign n3463 = ~n3363 & ~n3462;
  assign n3464 = sys_fair14done_out & ~n3463;
  assign n3465 = ~sys_fair14done_out & ~n1976;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = reg_stateG12_out & ~n3466;
  assign n3468 = ~n1977 & ~n3467;
  assign n3469 = ~sys_fair15done_out & ~n3468;
  assign n3470 = ~n3116 & ~n3469;
  assign n3471 = fair_cnt<1>_out  & ~n3470;
  assign n3472 = ~n1982 & ~n3471;
  assign n3473 = ~fair_cnt<0>_out  & ~n3472;
  assign n3474 = ~n1984 & ~n3473;
  assign n3475 = env_fair1done_out & ~n3474;
  assign n3476 = ~env_fair1done_out & ~n1986;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = ~reg_i_RtoB_ACK1_out & ~n3477;
  assign n3479 = ~n3115 & ~n3478;
  assign n3480 = reg_i_RtoB_ACK0_out & ~n3479;
  assign n3481 = sys_fair15done_out & ~n2268;
  assign n3482 = reg_controllable_BtoS_ACK0_out & ~n2451;
  assign n3483 = ~n1578 & ~n3482;
  assign n3484 = reg_i_StoB_REQ0_out & ~n3483;
  assign n3485 = reg_controllable_BtoS_ACK12_out & ~n2329;
  assign n3486 = ~n1500 & ~n3485;
  assign n3487 = reg_i_StoB_REQ12_out & ~n3486;
  assign n3488 = reg_controllable_BtoS_ACK7_out & ~n2315;
  assign n3489 = ~n1386 & ~n3488;
  assign n3490 = reg_i_StoB_REQ7_out & ~n3489;
  assign n3491 = ~n1642 & ~n2359;
  assign n3492 = sys_fair1done_out & ~n3491;
  assign n3493 = ~n3266 & ~n3492;
  assign n3494 = ~reg_i_StoB_REQ3_out & ~n3493;
  assign n3495 = ~n2368 & ~n3494;
  assign n3496 = sys_fair3done_out & ~n3495;
  assign n3497 = ~n3274 & ~n3496;
  assign n3498 = ~reg_i_StoB_REQ4_out & ~n3497;
  assign n3499 = ~n2377 & ~n3498;
  assign n3500 = sys_fair4done_out & ~n3499;
  assign n3501 = ~n3282 & ~n3500;
  assign n3502 = ~reg_i_StoB_REQ5_out & ~n3501;
  assign n3503 = ~n2386 & ~n3502;
  assign n3504 = sys_fair5done_out & ~n3503;
  assign n3505 = ~n3290 & ~n3504;
  assign n3506 = ~reg_i_StoB_REQ8_out & ~n3505;
  assign n3507 = ~n2395 & ~n3506;
  assign n3508 = sys_fair8done_out & ~n3507;
  assign n3509 = ~n3298 & ~n3508;
  assign n3510 = ~reg_i_StoB_REQ6_out & ~n3509;
  assign n3511 = ~n2404 & ~n3510;
  assign n3512 = sys_fair6done_out & ~n3511;
  assign n3513 = ~n3306 & ~n3512;
  assign n3514 = sys_fair7done_out & ~n3513;
  assign n3515 = ~n1350 & ~n3514;
  assign n3516 = ~reg_i_StoB_REQ7_out & ~n3515;
  assign n3517 = ~n3490 & ~n3516;
  assign n3518 = ~reg_i_StoB_REQ9_out & ~n3517;
  assign n3519 = ~n2417 & ~n3518;
  assign n3520 = sys_fair9done_out & ~n3519;
  assign n3521 = ~n3321 & ~n3520;
  assign n3522 = ~reg_i_StoB_REQ11_out & ~n3521;
  assign n3523 = ~n2426 & ~n3522;
  assign n3524 = sys_fair11done_out & ~n3523;
  assign n3525 = ~n3329 & ~n3524;
  assign n3526 = sys_fair12done_out & ~n3525;
  assign n3527 = ~n1464 & ~n3526;
  assign n3528 = ~reg_i_StoB_REQ12_out & ~n3527;
  assign n3529 = ~n3487 & ~n3528;
  assign n3530 = ~reg_i_StoB_REQ13_out & ~n3529;
  assign n3531 = ~n2439 & ~n3530;
  assign n3532 = sys_fair13done_out & ~n3531;
  assign n3533 = ~n3344 & ~n3532;
  assign n3534 = sys_fair0done_out & ~n3533;
  assign n3535 = ~n1542 & ~n3534;
  assign n3536 = ~reg_i_StoB_REQ0_out & ~n3535;
  assign n3537 = ~n3484 & ~n3536;
  assign n3538 = ~reg_i_StoB_REQ10_out & ~n3537;
  assign n3539 = ~n2456 & ~n3538;
  assign n3540 = sys_fair10done_out & ~n3539;
  assign n3541 = ~n3359 & ~n3540;
  assign n3542 = ~reg_i_StoB_REQ14_out & ~n3541;
  assign n3543 = ~n2470 & ~n3542;
  assign n3544 = sys_fair14done_out & ~n3543;
  assign n3545 = ~sys_fair14done_out & ~n2268;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = reg_stateG12_out & ~n3546;
  assign n3548 = ~n2269 & ~n3547;
  assign n3549 = ~sys_fair15done_out & ~n3548;
  assign n3550 = ~n3481 & ~n3549;
  assign n3551 = ~fair_cnt<1>_out  & ~n3550;
  assign n3552 = ~n2273 & ~n3551;
  assign n3553 = fair_cnt<0>_out  & ~n3552;
  assign n3554 = ~reg_i_StoB_REQ10_out & ~n3196;
  assign n3555 = ~n3199 & ~n3554;
  assign n3556 = sys_fair10done_out & ~n3555;
  assign n3557 = ~n2466 & ~n3556;
  assign n3558 = reg_controllable_BtoS_ACK14_out & ~n3557;
  assign n3559 = ~n3361 & ~n3558;
  assign n3560 = reg_i_StoB_REQ14_out & ~n3559;
  assign n3561 = ~reg_i_StoB_REQ14_out & ~n3360;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = sys_fair14done_out & ~n3562;
  assign n3564 = ~n3545 & ~n3563;
  assign n3565 = reg_stateG12_out & ~n3564;
  assign n3566 = ~n2269 & ~n3565;
  assign n3567 = ~sys_fair15done_out & ~n3566;
  assign n3568 = ~n3481 & ~n3567;
  assign n3569 = fair_cnt<1>_out  & ~n3568;
  assign n3570 = ~n2274 & ~n3569;
  assign n3571 = ~fair_cnt<0>_out  & ~n3570;
  assign n3572 = ~n3553 & ~n3571;
  assign n3573 = env_fair1done_out & ~n3572;
  assign n3574 = fair_cnt<0>_out  & ~n3570;
  assign n3575 = fair_cnt<1>_out  & ~n3550;
  assign n3576 = ~n2274 & ~n3575;
  assign n3577 = ~fair_cnt<0>_out  & ~n3576;
  assign n3578 = ~n3574 & ~n3577;
  assign n3579 = ~env_fair1done_out & ~n3578;
  assign n3580 = ~n3573 & ~n3579;
  assign n3581 = env_fair0done_out & ~n3580;
  assign n3582 = ~n2337 & ~n3190;
  assign n3583 = reg_controllable_BtoS_ACK0_out & ~n3582;
  assign n3584 = ~n3348 & ~n3583;
  assign n3585 = reg_i_StoB_REQ0_out & ~n3584;
  assign n3586 = ~n2343 & ~n3176;
  assign n3587 = reg_controllable_BtoS_ACK12_out & ~n3586;
  assign n3588 = ~n3333 & ~n3587;
  assign n3589 = reg_i_StoB_REQ12_out & ~n3588;
  assign n3590 = ~n2349 & ~n3155;
  assign n3591 = reg_controllable_BtoS_ACK7_out & ~n3590;
  assign n3592 = ~n3310 & ~n3591;
  assign n3593 = reg_i_StoB_REQ7_out & ~n3592;
  assign n3594 = ~sys_fair2done_out & ~n2354;
  assign n3595 = sys_fair1done_out & ~n3594;
  assign n3596 = ~n2361 & ~n3595;
  assign n3597 = ~reg_i_StoB_REQ3_out & ~n3596;
  assign n3598 = ~n3270 & ~n3597;
  assign n3599 = sys_fair3done_out & ~n3598;
  assign n3600 = ~n2370 & ~n3599;
  assign n3601 = ~reg_i_StoB_REQ4_out & ~n3600;
  assign n3602 = ~n3278 & ~n3601;
  assign n3603 = sys_fair4done_out & ~n3602;
  assign n3604 = ~n2379 & ~n3603;
  assign n3605 = ~reg_i_StoB_REQ5_out & ~n3604;
  assign n3606 = ~n3286 & ~n3605;
  assign n3607 = sys_fair5done_out & ~n3606;
  assign n3608 = ~n2388 & ~n3607;
  assign n3609 = ~reg_i_StoB_REQ8_out & ~n3608;
  assign n3610 = ~n3294 & ~n3609;
  assign n3611 = sys_fair8done_out & ~n3610;
  assign n3612 = ~n2397 & ~n3611;
  assign n3613 = ~reg_i_StoB_REQ6_out & ~n3612;
  assign n3614 = ~n3302 & ~n3613;
  assign n3615 = sys_fair6done_out & ~n3614;
  assign n3616 = ~n2406 & ~n3615;
  assign n3617 = sys_fair7done_out & ~n3616;
  assign n3618 = ~n1350 & ~n3617;
  assign n3619 = ~reg_i_StoB_REQ7_out & ~n3618;
  assign n3620 = ~n3593 & ~n3619;
  assign n3621 = ~reg_i_StoB_REQ9_out & ~n3620;
  assign n3622 = ~n3317 & ~n3621;
  assign n3623 = sys_fair9done_out & ~n3622;
  assign n3624 = ~n2419 & ~n3623;
  assign n3625 = ~reg_i_StoB_REQ11_out & ~n3624;
  assign n3626 = ~n3325 & ~n3625;
  assign n3627 = sys_fair11done_out & ~n3626;
  assign n3628 = ~n2428 & ~n3627;
  assign n3629 = sys_fair12done_out & ~n3628;
  assign n3630 = ~n1464 & ~n3629;
  assign n3631 = ~reg_i_StoB_REQ12_out & ~n3630;
  assign n3632 = ~n3589 & ~n3631;
  assign n3633 = ~reg_i_StoB_REQ13_out & ~n3632;
  assign n3634 = ~n3340 & ~n3633;
  assign n3635 = sys_fair13done_out & ~n3634;
  assign n3636 = ~n2441 & ~n3635;
  assign n3637 = sys_fair0done_out & ~n3636;
  assign n3638 = ~n1542 & ~n3637;
  assign n3639 = ~reg_i_StoB_REQ0_out & ~n3638;
  assign n3640 = ~n3585 & ~n3639;
  assign n3641 = ~reg_i_StoB_REQ10_out & ~n3640;
  assign n3642 = ~n3355 & ~n3641;
  assign n3643 = sys_fair10done_out & ~n3642;
  assign n3644 = ~n2458 & ~n3643;
  assign n3645 = ~reg_i_StoB_REQ14_out & ~n3644;
  assign n3646 = ~n3560 & ~n3645;
  assign n3647 = sys_fair14done_out & ~n3646;
  assign n3648 = ~n2472 & ~n3647;
  assign n3649 = reg_stateG12_out & ~n3648;
  assign n3650 = ~n2269 & ~n3649;
  assign n3651 = ~sys_fair15done_out & ~n3650;
  assign n3652 = ~n2474 & ~n3651;
  assign n3653 = fair_cnt<1>_out  & ~n3652;
  assign n3654 = ~n3551 & ~n3653;
  assign n3655 = fair_cnt<0>_out  & ~n3654;
  assign n3656 = ~n3577 & ~n3655;
  assign n3657 = env_fair1done_out & ~n3656;
  assign n3658 = ~n3579 & ~n3657;
  assign n3659 = ~env_fair0done_out & ~n3658;
  assign n3660 = ~n3581 & ~n3659;
  assign n3661 = reg_i_RtoB_ACK1_out & ~n3660;
  assign n3662 = ~fair_cnt<1>_out  & ~n3568;
  assign n3663 = ~n2273 & ~n3662;
  assign n3664 = fair_cnt<0>_out  & ~n3663;
  assign n3665 = ~n2244 & ~n2822;
  assign n3666 = reg_i_StoB_REQ14_out & ~n3665;
  assign n3667 = ~reg_i_StoB_REQ14_out & ~n2821;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = sys_fair14done_out & ~n3668;
  assign n3670 = ~n2828 & ~n3669;
  assign n3671 = reg_stateG12_out & ~n3670;
  assign n3672 = ~n2269 & ~n3671;
  assign n3673 = ~sys_fair15done_out & ~n3672;
  assign n3674 = ~n2830 & ~n3673;
  assign n3675 = fair_cnt<1>_out  & ~n3674;
  assign n3676 = ~n3551 & ~n3675;
  assign n3677 = ~fair_cnt<0>_out  & ~n3676;
  assign n3678 = ~n3664 & ~n3677;
  assign n3679 = env_fair1done_out & ~n3678;
  assign n3680 = ~env_fair1done_out & ~n3572;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = ~reg_i_RtoB_ACK1_out & ~n3681;
  assign n3683 = ~n3661 & ~n3682;
  assign n3684 = ~reg_i_RtoB_ACK0_out & ~n3683;
  assign n3685 = ~n3480 & ~n3684;
  assign n3686 = reg_nstateG7_1_out & ~n3685;
  assign n3687 = reg_nstateG7_1_out & ~n3686;
  assign n3688 = reg_stateG7_0_out & ~n3687;
  assign n3689 = ~reg_stateG7_0_out & ~n3685;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = ~reg_controllable_BtoR_REQ0_out & ~n3690;
  assign n3692 = ~reg_controllable_BtoR_REQ0_out & ~n3691;
  assign n3693 = reg_controllable_BtoR_REQ1_out & ~n3692;
  assign n3694 = env_fair0done_out & ~n3111;
  assign n3695 = ~env_fair0done_out & ~n701;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = reg_i_RtoB_ACK1_out & ~n3696;
  assign n3698 = ~env_fair1done_out & ~n3656;
  assign n3699 = ~n3573 & ~n3698;
  assign n3700 = env_fair0done_out & ~n3699;
  assign n3701 = ~env_fair0done_out & ~n3578;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = ~reg_i_RtoB_ACK1_out & ~n3702;
  assign n3704 = ~n3697 & ~n3703;
  assign n3705 = reg_i_RtoB_ACK0_out & ~n3704;
  assign n3706 = env_fair0done_out & ~n3474;
  assign n3707 = ~env_fair0done_out & ~n1986;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = reg_i_RtoB_ACK1_out & ~n3708;
  assign n3710 = env_fair0done_out & ~n3678;
  assign n3711 = ~env_fair0done_out & ~n3572;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~reg_i_RtoB_ACK1_out & ~n3712;
  assign n3714 = ~n3709 & ~n3713;
  assign n3715 = ~reg_i_RtoB_ACK0_out & ~n3714;
  assign n3716 = ~n3705 & ~n3715;
  assign n3717 = ~reg_nstateG7_1_out & ~n3716;
  assign n3718 = ~reg_nstateG7_1_out & ~n3717;
  assign n3719 = reg_stateG7_0_out & ~n3718;
  assign n3720 = ~reg_stateG7_0_out & ~n3716;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = reg_controllable_BtoR_REQ0_out & ~n3721;
  assign n3723 = ~n2903 & ~n3577;
  assign n3724 = reg_i_RtoB_ACK1_out & ~n3723;
  assign n3725 = env_fair1done_out & ~n3723;
  assign n3726 = ~n2274 & ~n3653;
  assign n3727 = fair_cnt<0>_out  & ~n3726;
  assign n3728 = ~n3577 & ~n3727;
  assign n3729 = ~env_fair1done_out & ~n3728;
  assign n3730 = ~n3725 & ~n3729;
  assign n3731 = ~reg_i_RtoB_ACK1_out & ~n3730;
  assign n3732 = ~n3724 & ~n3731;
  assign n3733 = reg_i_RtoB_ACK0_out & ~n3732;
  assign n3734 = fair_cnt<0>_out  & ~n3676;
  assign n3735 = ~n3571 & ~n3734;
  assign n3736 = ~env_fair1done_out & ~n3735;
  assign n3737 = ~n3679 & ~n3736;
  assign n3738 = ~reg_i_RtoB_ACK1_out & ~n3737;
  assign n3739 = ~n3724 & ~n3738;
  assign n3740 = ~reg_i_RtoB_ACK0_out & ~n3739;
  assign n3741 = ~n3733 & ~n3740;
  assign n3742 = reg_nstateG7_1_out & ~n3741;
  assign n3743 = reg_i_RtoB_ACK0_out & ~n3723;
  assign n3744 = env_fair0done_out & ~n3723;
  assign n3745 = ~env_fair0done_out & ~n3728;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = reg_i_RtoB_ACK1_out & ~n3746;
  assign n3748 = ~env_fair0done_out & ~n3735;
  assign n3749 = ~n3710 & ~n3748;
  assign n3750 = ~reg_i_RtoB_ACK1_out & ~n3749;
  assign n3751 = ~n3747 & ~n3750;
  assign n3752 = ~reg_i_RtoB_ACK0_out & ~n3751;
  assign n3753 = ~n3743 & ~n3752;
  assign n3754 = ~reg_nstateG7_1_out & ~n3753;
  assign n3755 = ~n3742 & ~n3754;
  assign n3756 = ~reg_controllable_BtoR_REQ0_out & ~n3755;
  assign n3757 = ~n3722 & ~n3756;
  assign n3758 = ~reg_controllable_BtoR_REQ1_out & ~n3757;
  assign n3759 = ~n3693 & ~n3758;
  assign n3760 = ~reg_controllable_DEQ_out & ~n3759;
  assign n3761 = ~n3105 & ~n3760;
  assign n3762 = reg_i_nEMPTY_out & ~n3761;
  assign n3763 = ~reg_controllable_ENQ_out & ~n3103;
  assign n3764 = reg_controllable_DEQ_out & ~n3763;
  assign n3765 = reg_controllable_ENQ_out & ~n3759;
  assign n3766 = reg_controllable_ENQ_out & ~n3765;
  assign n3767 = ~reg_controllable_DEQ_out & ~n3766;
  assign n3768 = ~n3764 & ~n3767;
  assign n3769 = ~reg_i_nEMPTY_out & ~n3768;
  assign n3770 = ~n3762 & ~n3769;
  assign n3771 = reg_i_FULL_out & ~n3770;
  assign n3772 = ~n2280 & ~n2906;
  assign n3773 = env_fair0done_out & ~n3772;
  assign n3774 = ~n2549 & ~n3773;
  assign n3775 = reg_i_RtoB_ACK1_out & ~n3774;
  assign n3776 = ~reg_i_RtoB_ACK1_out & ~n2904;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = ~reg_i_RtoB_ACK0_out & ~n3777;
  assign n3779 = ~n1989 & ~n3778;
  assign n3780 = reg_nstateG7_1_out & ~n3779;
  assign n3781 = reg_nstateG7_1_out & ~n3780;
  assign n3782 = reg_stateG7_0_out & ~n3781;
  assign n3783 = ~reg_stateG7_0_out & ~n3779;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~reg_controllable_BtoR_REQ0_out & ~n3784;
  assign n3786 = ~reg_controllable_BtoR_REQ0_out & ~n3785;
  assign n3787 = reg_controllable_BtoR_REQ1_out & ~n3786;
  assign n3788 = env_fair0done_out & ~n2907;
  assign n3789 = ~n2859 & ~n3788;
  assign n3790 = ~reg_i_RtoB_ACK1_out & ~n3789;
  assign n3791 = ~n2855 & ~n3790;
  assign n3792 = reg_i_RtoB_ACK0_out & ~n3791;
  assign n3793 = ~n2864 & ~n3776;
  assign n3794 = ~reg_i_RtoB_ACK0_out & ~n3793;
  assign n3795 = ~n3792 & ~n3794;
  assign n3796 = ~reg_nstateG7_1_out & ~n3795;
  assign n3797 = ~reg_nstateG7_1_out & ~n3796;
  assign n3798 = reg_stateG7_0_out & ~n3797;
  assign n3799 = ~reg_stateG7_0_out & ~n3795;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = reg_controllable_BtoR_REQ0_out & ~n3800;
  assign n3802 = ~reg_i_RtoB_ACK1_out & ~n3772;
  assign n3803 = ~n2905 & ~n3802;
  assign n3804 = ~reg_i_RtoB_ACK0_out & ~n3803;
  assign n3805 = ~n2910 & ~n3804;
  assign n3806 = reg_nstateG7_1_out & ~n3805;
  assign n3807 = ~n2859 & ~n2921;
  assign n3808 = ~reg_i_RtoB_ACK1_out & ~n3807;
  assign n3809 = ~n2924 & ~n3808;
  assign n3810 = ~reg_i_RtoB_ACK0_out & ~n3809;
  assign n3811 = ~n2920 & ~n3810;
  assign n3812 = ~reg_nstateG7_1_out & ~n3811;
  assign n3813 = ~n3806 & ~n3812;
  assign n3814 = ~reg_controllable_BtoR_REQ0_out & ~n3813;
  assign n3815 = ~n3801 & ~n3814;
  assign n3816 = ~reg_controllable_BtoR_REQ1_out & ~n3815;
  assign n3817 = ~n3787 & ~n3816;
  assign n3818 = reg_controllable_ENQ_out & ~n3817;
  assign n3819 = ~n3103 & ~n3818;
  assign n3820 = reg_controllable_DEQ_out & ~n3819;
  assign n3821 = ~n2901 & ~n3551;
  assign n3822 = fair_cnt<0>_out  & ~n3821;
  assign n3823 = ~n3571 & ~n3822;
  assign n3824 = env_fair1done_out & ~n3823;
  assign n3825 = ~n3579 & ~n3824;
  assign n3826 = env_fair0done_out & ~n3825;
  assign n3827 = ~n3659 & ~n3826;
  assign n3828 = reg_i_RtoB_ACK1_out & ~n3827;
  assign n3829 = ~n2901 & ~n3662;
  assign n3830 = fair_cnt<0>_out  & ~n3829;
  assign n3831 = ~n3551 & ~n3569;
  assign n3832 = ~fair_cnt<0>_out  & ~n3831;
  assign n3833 = ~n3830 & ~n3832;
  assign n3834 = env_fair1done_out & ~n3833;
  assign n3835 = ~env_fair1done_out & ~n3823;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~reg_i_RtoB_ACK1_out & ~n3836;
  assign n3838 = ~n3828 & ~n3837;
  assign n3839 = ~reg_i_RtoB_ACK0_out & ~n3838;
  assign n3840 = ~n3480 & ~n3839;
  assign n3841 = reg_nstateG7_1_out & ~n3840;
  assign n3842 = reg_nstateG7_1_out & ~n3841;
  assign n3843 = reg_stateG7_0_out & ~n3842;
  assign n3844 = ~reg_stateG7_0_out & ~n3840;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~reg_controllable_BtoR_REQ0_out & ~n3845;
  assign n3847 = ~reg_controllable_BtoR_REQ0_out & ~n3846;
  assign n3848 = reg_controllable_BtoR_REQ1_out & ~n3847;
  assign n3849 = ~n3698 & ~n3824;
  assign n3850 = env_fair0done_out & ~n3849;
  assign n3851 = ~n3701 & ~n3850;
  assign n3852 = ~reg_i_RtoB_ACK1_out & ~n3851;
  assign n3853 = ~n3697 & ~n3852;
  assign n3854 = reg_i_RtoB_ACK0_out & ~n3853;
  assign n3855 = env_fair0done_out & ~n3833;
  assign n3856 = ~env_fair0done_out & ~n3823;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = ~reg_i_RtoB_ACK1_out & ~n3857;
  assign n3859 = ~n3709 & ~n3858;
  assign n3860 = ~reg_i_RtoB_ACK0_out & ~n3859;
  assign n3861 = ~n3854 & ~n3860;
  assign n3862 = ~reg_nstateG7_1_out & ~n3861;
  assign n3863 = ~reg_nstateG7_1_out & ~n3862;
  assign n3864 = reg_stateG7_0_out & ~n3863;
  assign n3865 = ~reg_stateG7_0_out & ~n3861;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = reg_controllable_BtoR_REQ0_out & ~n3866;
  assign n3868 = fair_cnt<0>_out  & ~n3831;
  assign n3869 = ~n3571 & ~n3868;
  assign n3870 = ~env_fair1done_out & ~n3869;
  assign n3871 = ~n3834 & ~n3870;
  assign n3872 = ~reg_i_RtoB_ACK1_out & ~n3871;
  assign n3873 = ~n3724 & ~n3872;
  assign n3874 = ~reg_i_RtoB_ACK0_out & ~n3873;
  assign n3875 = ~n3733 & ~n3874;
  assign n3876 = reg_nstateG7_1_out & ~n3875;
  assign n3877 = ~env_fair0done_out & ~n3869;
  assign n3878 = ~n3855 & ~n3877;
  assign n3879 = ~reg_i_RtoB_ACK1_out & ~n3878;
  assign n3880 = ~n3747 & ~n3879;
  assign n3881 = ~reg_i_RtoB_ACK0_out & ~n3880;
  assign n3882 = ~n3743 & ~n3881;
  assign n3883 = ~reg_nstateG7_1_out & ~n3882;
  assign n3884 = ~n3876 & ~n3883;
  assign n3885 = ~reg_controllable_BtoR_REQ0_out & ~n3884;
  assign n3886 = ~n3867 & ~n3885;
  assign n3887 = ~reg_controllable_BtoR_REQ1_out & ~n3886;
  assign n3888 = ~n3848 & ~n3887;
  assign n3889 = ~reg_controllable_ENQ_out & ~n3888;
  assign n3890 = ~n3765 & ~n3889;
  assign n3891 = ~reg_controllable_DEQ_out & ~n3890;
  assign n3892 = ~n3820 & ~n3891;
  assign n3893 = reg_i_nEMPTY_out & ~n3892;
  assign n3894 = reg_controllable_DEQ_out & ~n3102;
  assign n3895 = ~fair_cnt<1>_out  & ~n3107;
  assign n3896 = ~n696 & ~n3895;
  assign n3897 = fair_cnt<0>_out  & ~n3896;
  assign n3898 = ~reg_controllable_BtoS_ACK14_out & ~n3557;
  assign n3899 = ~reg_controllable_BtoS_ACK14_out & ~n3898;
  assign n3900 = reg_i_StoB_REQ14_out & ~n3899;
  assign n3901 = ~reg_i_StoB_REQ14_out & ~n3250;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = sys_fair14done_out & ~n3902;
  assign n3904 = ~n3047 & ~n3903;
  assign n3905 = reg_stateG12_out & ~n3904;
  assign n3906 = ~n692 & ~n3905;
  assign n3907 = ~sys_fair15done_out & ~n3906;
  assign n3908 = ~n3106 & ~n3907;
  assign n3909 = fair_cnt<1>_out  & ~n3908;
  assign n3910 = ~n697 & ~n3909;
  assign n3911 = ~fair_cnt<0>_out  & ~n3910;
  assign n3912 = ~n3897 & ~n3911;
  assign n3913 = env_fair1done_out & ~n3912;
  assign n3914 = ~env_fair1done_out & ~n3111;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = env_fair0done_out & ~n3915;
  assign n3917 = ~n3110 & ~n3897;
  assign n3918 = env_fair1done_out & ~n3917;
  assign n3919 = ~n3914 & ~n3918;
  assign n3920 = ~env_fair0done_out & ~n3919;
  assign n3921 = ~n3916 & ~n3920;
  assign n3922 = reg_i_RtoB_ACK1_out & ~n3921;
  assign n3923 = ~fair_cnt<1>_out  & ~n3470;
  assign n3924 = ~n1981 & ~n3923;
  assign n3925 = fair_cnt<0>_out  & ~n3924;
  assign n3926 = reg_controllable_BtoS_ACK14_out & ~n3043;
  assign n3927 = ~reg_controllable_BtoS_ACK14_out & ~n3541;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = reg_i_StoB_REQ14_out & ~n3928;
  assign n3930 = reg_controllable_BtoS_ACK10_out & ~n3038;
  assign n3931 = ~reg_controllable_BtoS_ACK10_out & ~n3537;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = reg_i_StoB_REQ10_out & ~n3932;
  assign n3934 = reg_controllable_BtoS_ACK0_out & ~n3036;
  assign n3935 = ~reg_controllable_BtoS_ACK0_out & ~n3535;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = reg_i_StoB_REQ0_out & ~n3936;
  assign n3938 = reg_controllable_BtoS_ACK13_out & ~n3029;
  assign n3939 = ~reg_controllable_BtoS_ACK13_out & ~n3529;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = reg_i_StoB_REQ13_out & ~n3940;
  assign n3942 = reg_controllable_BtoS_ACK12_out & ~n3027;
  assign n3943 = ~reg_controllable_BtoS_ACK12_out & ~n3527;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = reg_i_StoB_REQ12_out & ~n3944;
  assign n3946 = reg_controllable_BtoS_ACK11_out & ~n3020;
  assign n3947 = ~reg_controllable_BtoS_ACK11_out & ~n3521;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = reg_i_StoB_REQ11_out & ~n3948;
  assign n3950 = reg_controllable_BtoS_ACK9_out & ~n3015;
  assign n3951 = ~reg_controllable_BtoS_ACK9_out & ~n3517;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = reg_i_StoB_REQ9_out & ~n3952;
  assign n3954 = reg_controllable_BtoS_ACK7_out & ~n3013;
  assign n3955 = ~reg_controllable_BtoS_ACK7_out & ~n3515;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = reg_i_StoB_REQ7_out & ~n3956;
  assign n3958 = reg_controllable_BtoS_ACK6_out & ~n3006;
  assign n3959 = ~reg_controllable_BtoS_ACK6_out & ~n3509;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = reg_i_StoB_REQ6_out & ~n3960;
  assign n3962 = reg_controllable_BtoS_ACK8_out & ~n3001;
  assign n3963 = ~reg_controllable_BtoS_ACK8_out & ~n3505;
  assign n3964 = ~n3962 & ~n3963;
  assign n3965 = reg_i_StoB_REQ8_out & ~n3964;
  assign n3966 = reg_controllable_BtoS_ACK5_out & ~n2996;
  assign n3967 = ~reg_controllable_BtoS_ACK5_out & ~n3501;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = reg_i_StoB_REQ5_out & ~n3968;
  assign n3970 = reg_controllable_BtoS_ACK4_out & ~n2991;
  assign n3971 = ~reg_controllable_BtoS_ACK4_out & ~n3497;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = reg_i_StoB_REQ4_out & ~n3972;
  assign n3974 = reg_controllable_BtoS_ACK3_out & ~n2986;
  assign n3975 = ~reg_controllable_BtoS_ACK3_out & ~n3493;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = reg_i_StoB_REQ3_out & ~n3976;
  assign n3978 = ~n2982 & ~n3400;
  assign n3979 = sys_fair1done_out & ~n3978;
  assign n3980 = ~n3403 & ~n3979;
  assign n3981 = ~reg_i_StoB_REQ3_out & ~n3980;
  assign n3982 = ~n3977 & ~n3981;
  assign n3983 = sys_fair3done_out & ~n3982;
  assign n3984 = ~n3408 & ~n3983;
  assign n3985 = ~reg_i_StoB_REQ4_out & ~n3984;
  assign n3986 = ~n3973 & ~n3985;
  assign n3987 = sys_fair4done_out & ~n3986;
  assign n3988 = ~n3413 & ~n3987;
  assign n3989 = ~reg_i_StoB_REQ5_out & ~n3988;
  assign n3990 = ~n3969 & ~n3989;
  assign n3991 = sys_fair5done_out & ~n3990;
  assign n3992 = ~n3418 & ~n3991;
  assign n3993 = ~reg_i_StoB_REQ8_out & ~n3992;
  assign n3994 = ~n3965 & ~n3993;
  assign n3995 = sys_fair8done_out & ~n3994;
  assign n3996 = ~n3423 & ~n3995;
  assign n3997 = ~reg_i_StoB_REQ6_out & ~n3996;
  assign n3998 = ~n3961 & ~n3997;
  assign n3999 = sys_fair6done_out & ~n3998;
  assign n4000 = ~n3428 & ~n3999;
  assign n4001 = sys_fair7done_out & ~n4000;
  assign n4002 = ~n1754 & ~n4001;
  assign n4003 = ~reg_i_StoB_REQ7_out & ~n4002;
  assign n4004 = ~n3957 & ~n4003;
  assign n4005 = ~reg_i_StoB_REQ9_out & ~n4004;
  assign n4006 = ~n3953 & ~n4005;
  assign n4007 = sys_fair9done_out & ~n4006;
  assign n4008 = ~n3437 & ~n4007;
  assign n4009 = ~reg_i_StoB_REQ11_out & ~n4008;
  assign n4010 = ~n3949 & ~n4009;
  assign n4011 = sys_fair11done_out & ~n4010;
  assign n4012 = ~n3442 & ~n4011;
  assign n4013 = sys_fair12done_out & ~n4012;
  assign n4014 = ~n1825 & ~n4013;
  assign n4015 = ~reg_i_StoB_REQ12_out & ~n4014;
  assign n4016 = ~n3945 & ~n4015;
  assign n4017 = ~reg_i_StoB_REQ13_out & ~n4016;
  assign n4018 = ~n3941 & ~n4017;
  assign n4019 = sys_fair13done_out & ~n4018;
  assign n4020 = ~n3451 & ~n4019;
  assign n4021 = sys_fair0done_out & ~n4020;
  assign n4022 = ~n1873 & ~n4021;
  assign n4023 = ~reg_i_StoB_REQ0_out & ~n4022;
  assign n4024 = ~n3937 & ~n4023;
  assign n4025 = ~reg_i_StoB_REQ10_out & ~n4024;
  assign n4026 = ~n3933 & ~n4025;
  assign n4027 = sys_fair10done_out & ~n4026;
  assign n4028 = ~n3460 & ~n4027;
  assign n4029 = ~reg_i_StoB_REQ14_out & ~n4028;
  assign n4030 = ~n3929 & ~n4029;
  assign n4031 = sys_fair14done_out & ~n4030;
  assign n4032 = ~n3465 & ~n4031;
  assign n4033 = reg_stateG12_out & ~n4032;
  assign n4034 = ~n1977 & ~n4033;
  assign n4035 = ~sys_fair15done_out & ~n4034;
  assign n4036 = ~n3116 & ~n4035;
  assign n4037 = ~fair_cnt<1>_out  & ~n4036;
  assign n4038 = ~n3471 & ~n4037;
  assign n4039 = ~fair_cnt<0>_out  & ~n4038;
  assign n4040 = ~n3925 & ~n4039;
  assign n4041 = env_fair1done_out & ~n4040;
  assign n4042 = ~n1981 & ~n4037;
  assign n4043 = fair_cnt<0>_out  & ~n4042;
  assign n4044 = ~n3473 & ~n4043;
  assign n4045 = ~env_fair1done_out & ~n4044;
  assign n4046 = ~n4041 & ~n4045;
  assign n4047 = ~reg_i_RtoB_ACK1_out & ~n4046;
  assign n4048 = ~n3922 & ~n4047;
  assign n4049 = ~reg_i_RtoB_ACK0_out & ~n4048;
  assign n4050 = ~reg_i_RtoB_ACK0_out & ~n4049;
  assign n4051 = reg_nstateG7_1_out & ~n4050;
  assign n4052 = reg_nstateG7_1_out & ~n4051;
  assign n4053 = reg_stateG7_0_out & ~n4052;
  assign n4054 = ~reg_stateG7_0_out & ~n4050;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~reg_controllable_BtoR_REQ0_out & ~n4055;
  assign n4057 = ~reg_controllable_BtoR_REQ0_out & ~n4056;
  assign n4058 = reg_controllable_BtoR_REQ1_out & ~n4057;
  assign n4059 = ~env_fair1done_out & ~n3917;
  assign n4060 = ~n3913 & ~n4059;
  assign n4061 = env_fair0done_out & ~n4060;
  assign n4062 = ~env_fair0done_out & ~n3111;
  assign n4063 = ~n4061 & ~n4062;
  assign n4064 = ~reg_i_RtoB_ACK1_out & ~n4063;
  assign n4065 = ~reg_i_RtoB_ACK1_out & ~n4064;
  assign n4066 = reg_i_RtoB_ACK0_out & ~n4065;
  assign n4067 = env_fair0done_out & ~n4040;
  assign n4068 = ~env_fair0done_out & ~n4044;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~reg_i_RtoB_ACK1_out & ~n4069;
  assign n4071 = ~reg_i_RtoB_ACK1_out & ~n4070;
  assign n4072 = ~reg_i_RtoB_ACK0_out & ~n4071;
  assign n4073 = ~n4066 & ~n4072;
  assign n4074 = ~reg_nstateG7_1_out & ~n4073;
  assign n4075 = ~reg_nstateG7_1_out & ~n4074;
  assign n4076 = reg_stateG7_0_out & ~n4075;
  assign n4077 = ~reg_stateG7_0_out & ~n4073;
  assign n4078 = ~n4076 & ~n4077;
  assign n4079 = reg_controllable_BtoR_REQ0_out & ~n4078;
  assign n4080 = reg_stateG12_out & ~n1952;
  assign n4081 = ~reg_stateG12_out & ~n2889;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = sys_fair15done_out & ~n4082;
  assign n4084 = ~n1967 & ~n2269;
  assign n4085 = ~sys_fair15done_out & ~n4084;
  assign n4086 = ~n4083 & ~n4085;
  assign n4087 = fair_cnt<1>_out  & ~n4086;
  assign n4088 = reg_stateG12_out & ~n1976;
  assign n4089 = ~n2269 & ~n4088;
  assign n4090 = sys_fair15done_out & ~n4089;
  assign n4091 = ~n2269 & ~n3467;
  assign n4092 = ~sys_fair15done_out & ~n4091;
  assign n4093 = ~n4090 & ~n4092;
  assign n4094 = ~fair_cnt<1>_out  & ~n4093;
  assign n4095 = ~n4087 & ~n4094;
  assign n4096 = fair_cnt<0>_out  & ~n4095;
  assign n4097 = fair_cnt<1>_out  & ~n4093;
  assign n4098 = ~n2269 & ~n4033;
  assign n4099 = ~sys_fair15done_out & ~n4098;
  assign n4100 = ~n4090 & ~n4099;
  assign n4101 = ~fair_cnt<1>_out  & ~n4100;
  assign n4102 = ~n4097 & ~n4101;
  assign n4103 = ~fair_cnt<0>_out  & ~n4102;
  assign n4104 = ~n4096 & ~n4103;
  assign n4105 = env_fair1done_out & ~n4104;
  assign n4106 = ~reg_stateG12_out & ~n2473;
  assign n4107 = ~n4088 & ~n4106;
  assign n4108 = sys_fair15done_out & ~n4107;
  assign n4109 = ~n4092 & ~n4108;
  assign n4110 = fair_cnt<1>_out  & ~n4109;
  assign n4111 = ~n4101 & ~n4110;
  assign n4112 = fair_cnt<0>_out  & ~n4111;
  assign n4113 = ~fair_cnt<1>_out  & ~n4089;
  assign n4114 = ~n4097 & ~n4113;
  assign n4115 = ~fair_cnt<0>_out  & ~n4114;
  assign n4116 = ~n4112 & ~n4115;
  assign n4117 = ~env_fair1done_out & ~n4116;
  assign n4118 = ~n4105 & ~n4117;
  assign n4119 = ~reg_i_RtoB_ACK1_out & ~n4118;
  assign n4120 = ~reg_i_RtoB_ACK1_out & ~n4119;
  assign n4121 = ~reg_i_RtoB_ACK0_out & ~n4120;
  assign n4122 = ~reg_i_RtoB_ACK0_out & ~n4121;
  assign n4123 = reg_nstateG7_1_out & ~n4122;
  assign n4124 = env_fair0done_out & ~n4104;
  assign n4125 = ~env_fair0done_out & ~n4116;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~reg_i_RtoB_ACK1_out & ~n4126;
  assign n4128 = ~reg_i_RtoB_ACK1_out & ~n4127;
  assign n4129 = ~reg_i_RtoB_ACK0_out & ~n4128;
  assign n4130 = ~reg_i_RtoB_ACK0_out & ~n4129;
  assign n4131 = ~reg_nstateG7_1_out & ~n4130;
  assign n4132 = ~n4123 & ~n4131;
  assign n4133 = ~reg_controllable_BtoR_REQ0_out & ~n4132;
  assign n4134 = ~n4079 & ~n4133;
  assign n4135 = ~reg_controllable_BtoR_REQ1_out & ~n4134;
  assign n4136 = ~n4058 & ~n4135;
  assign n4137 = ~reg_controllable_ENQ_out & ~n4136;
  assign n4138 = ~n3765 & ~n4137;
  assign n4139 = ~reg_controllable_DEQ_out & ~n4138;
  assign n4140 = ~n3894 & ~n4139;
  assign n4141 = ~reg_i_nEMPTY_out & ~n4140;
  assign n4142 = ~n3893 & ~n4141;
  assign n4143 = ~reg_i_FULL_out & ~n4142;
  assign n4144 = ~n3771 & ~n4143;
  assign n4145 = ~fair_cnt<2>_out  & ~n4144;
  assign n4146 = ~fair_cnt<2>_out  & ~n4145;
  assign n4147 = ~env_safe_err_happened_out & n4146;
  assign n4148 = ~env_safe_err_happened_out & ~n4147;
  assign n4149 = n87 & ~n4148;
  assign n4150 = n87 & ~n4149;
  assign n4151 = n87 & reg_stateG12_out;
  assign n4152 = n87 & sys_fair15done_out;
  assign n4153 = n4151 & ~n4152;
  assign n4154 = n87 & sys_fair8done_out;
  assign n4155 = ~i_StoB_REQ8 & controllable_BtoS_ACK8;
  assign n4156 = i_StoB_REQ8 & ~controllable_BtoS_ACK8;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4154 & ~n4157;
  assign n4159 = ~i_StoB_REQ0 & controllable_BtoS_ACK0;
  assign n4160 = i_StoB_REQ0 & ~controllable_BtoS_ACK0;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = n87 & sys_fair0done_out;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~i_StoB_REQ1 & controllable_BtoS_ACK1;
  assign n4165 = i_StoB_REQ1 & ~controllable_BtoS_ACK1;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = n87 & sys_fair1done_out;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = ~n4163 & ~n4168;
  assign n4170 = ~i_StoB_REQ2 & controllable_BtoS_ACK2;
  assign n4171 = i_StoB_REQ2 & ~controllable_BtoS_ACK2;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = n87 & sys_fair2done_out;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = n4169 & ~n4174;
  assign n4176 = ~i_StoB_REQ3 & controllable_BtoS_ACK3;
  assign n4177 = i_StoB_REQ3 & ~controllable_BtoS_ACK3;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = n87 & sys_fair3done_out;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = n4175 & ~n4180;
  assign n4182 = ~i_StoB_REQ4 & controllable_BtoS_ACK4;
  assign n4183 = i_StoB_REQ4 & ~controllable_BtoS_ACK4;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = n87 & sys_fair4done_out;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = n4181 & ~n4186;
  assign n4188 = ~i_StoB_REQ5 & controllable_BtoS_ACK5;
  assign n4189 = i_StoB_REQ5 & ~controllable_BtoS_ACK5;
  assign n4190 = ~n4188 & ~n4189;
  assign n4191 = n87 & sys_fair5done_out;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = n4187 & ~n4192;
  assign n4194 = ~i_StoB_REQ6 & controllable_BtoS_ACK6;
  assign n4195 = i_StoB_REQ6 & ~controllable_BtoS_ACK6;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = n87 & sys_fair6done_out;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = n4193 & ~n4198;
  assign n4200 = ~i_StoB_REQ7 & controllable_BtoS_ACK7;
  assign n4201 = i_StoB_REQ7 & ~controllable_BtoS_ACK7;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = n87 & sys_fair7done_out;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = n4199 & ~n4204;
  assign n4206 = ~n4158 & n4205;
  assign n4207 = ~i_StoB_REQ9 & controllable_BtoS_ACK9;
  assign n4208 = i_StoB_REQ9 & ~controllable_BtoS_ACK9;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = n87 & sys_fair9done_out;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = n4206 & ~n4211;
  assign n4213 = ~i_StoB_REQ10 & controllable_BtoS_ACK10;
  assign n4214 = i_StoB_REQ10 & ~controllable_BtoS_ACK10;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = n87 & sys_fair10done_out;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = n4212 & ~n4217;
  assign n4219 = ~i_StoB_REQ11 & controllable_BtoS_ACK11;
  assign n4220 = i_StoB_REQ11 & ~controllable_BtoS_ACK11;
  assign n4221 = ~n4219 & ~n4220;
  assign n4222 = n87 & sys_fair11done_out;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = n4218 & ~n4223;
  assign n4225 = ~i_StoB_REQ12 & controllable_BtoS_ACK12;
  assign n4226 = i_StoB_REQ12 & ~controllable_BtoS_ACK12;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = n87 & sys_fair12done_out;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = n4224 & ~n4229;
  assign n4231 = ~i_StoB_REQ13 & controllable_BtoS_ACK13;
  assign n4232 = i_StoB_REQ13 & ~controllable_BtoS_ACK13;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = n87 & sys_fair13done_out;
  assign n4235 = ~n4233 & ~n4234;
  assign n4236 = n4230 & ~n4235;
  assign n4237 = ~i_StoB_REQ14 & controllable_BtoS_ACK14;
  assign n4238 = i_StoB_REQ14 & ~controllable_BtoS_ACK14;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = n87 & sys_fair14done_out;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = n4236 & ~n4241;
  assign n4243 = ~n4153 & n4242;
  assign n4244 = ~n4153 & ~n4243;
  assign n4245 = n87 & reg_i_StoB_REQ1_out;
  assign n4246 = n87 & reg_controllable_BtoS_ACK1_out;
  assign n4247 = n4245 & ~n4246;
  assign n4248 = ~i_StoB_REQ1 & n4247;
  assign n4249 = n87 & reg_controllable_BtoS_ACK0_out;
  assign n4250 = ~i_StoB_REQ0 & n4249;
  assign n4251 = n87 & reg_i_StoB_REQ0_out;
  assign n4252 = ~i_StoB_REQ0 & n4251;
  assign n4253 = ~n4249 & ~n4252;
  assign n4254 = ~n4250 & ~n4253;
  assign n4255 = ~n4248 & ~n4254;
  assign n4256 = i_StoB_REQ1 & n4246;
  assign n4257 = n4255 & ~n4256;
  assign n4258 = n87 & reg_i_StoB_REQ2_out;
  assign n4259 = n87 & reg_controllable_BtoS_ACK2_out;
  assign n4260 = n4258 & ~n4259;
  assign n4261 = ~i_StoB_REQ2 & n4260;
  assign n4262 = n4257 & ~n4261;
  assign n4263 = i_StoB_REQ2 & n4259;
  assign n4264 = n4262 & ~n4263;
  assign n4265 = n87 & reg_i_StoB_REQ3_out;
  assign n4266 = n87 & reg_controllable_BtoS_ACK3_out;
  assign n4267 = n4265 & ~n4266;
  assign n4268 = ~i_StoB_REQ3 & n4267;
  assign n4269 = n4264 & ~n4268;
  assign n4270 = i_StoB_REQ3 & n4266;
  assign n4271 = n4269 & ~n4270;
  assign n4272 = n87 & reg_i_StoB_REQ4_out;
  assign n4273 = n87 & reg_controllable_BtoS_ACK4_out;
  assign n4274 = n4272 & ~n4273;
  assign n4275 = ~i_StoB_REQ4 & n4274;
  assign n4276 = n4271 & ~n4275;
  assign n4277 = i_StoB_REQ4 & n4273;
  assign n4278 = n4276 & ~n4277;
  assign n4279 = n87 & reg_i_StoB_REQ5_out;
  assign n4280 = n87 & reg_controllable_BtoS_ACK5_out;
  assign n4281 = n4279 & ~n4280;
  assign n4282 = ~i_StoB_REQ5 & n4281;
  assign n4283 = n4278 & ~n4282;
  assign n4284 = i_StoB_REQ5 & n4280;
  assign n4285 = n4283 & ~n4284;
  assign n4286 = n87 & reg_i_StoB_REQ6_out;
  assign n4287 = n87 & reg_controllable_BtoS_ACK6_out;
  assign n4288 = n4286 & ~n4287;
  assign n4289 = ~i_StoB_REQ6 & n4288;
  assign n4290 = n4285 & ~n4289;
  assign n4291 = i_StoB_REQ6 & n4287;
  assign n4292 = n4290 & ~n4291;
  assign n4293 = n87 & reg_i_StoB_REQ7_out;
  assign n4294 = n87 & reg_controllable_BtoS_ACK7_out;
  assign n4295 = n4293 & ~n4294;
  assign n4296 = ~i_StoB_REQ7 & n4295;
  assign n4297 = n4292 & ~n4296;
  assign n4298 = i_StoB_REQ7 & n4294;
  assign n4299 = n4297 & ~n4298;
  assign n4300 = n87 & reg_i_StoB_REQ8_out;
  assign n4301 = n87 & reg_controllable_BtoS_ACK8_out;
  assign n4302 = n4300 & ~n4301;
  assign n4303 = ~i_StoB_REQ8 & n4302;
  assign n4304 = n4299 & ~n4303;
  assign n4305 = i_StoB_REQ8 & n4301;
  assign n4306 = n4304 & ~n4305;
  assign n4307 = n87 & reg_i_StoB_REQ9_out;
  assign n4308 = n87 & reg_controllable_BtoS_ACK9_out;
  assign n4309 = n4307 & ~n4308;
  assign n4310 = ~i_StoB_REQ9 & n4309;
  assign n4311 = n4306 & ~n4310;
  assign n4312 = i_StoB_REQ9 & n4308;
  assign n4313 = n4311 & ~n4312;
  assign n4314 = n87 & reg_i_StoB_REQ10_out;
  assign n4315 = n87 & reg_controllable_BtoS_ACK10_out;
  assign n4316 = n4314 & ~n4315;
  assign n4317 = ~i_StoB_REQ10 & n4316;
  assign n4318 = n4313 & ~n4317;
  assign n4319 = i_StoB_REQ10 & n4315;
  assign n4320 = n4318 & ~n4319;
  assign n4321 = n87 & reg_i_StoB_REQ11_out;
  assign n4322 = n87 & reg_controllable_BtoS_ACK11_out;
  assign n4323 = n4321 & ~n4322;
  assign n4324 = ~i_StoB_REQ11 & n4323;
  assign n4325 = n4320 & ~n4324;
  assign n4326 = i_StoB_REQ11 & n4322;
  assign n4327 = n4325 & ~n4326;
  assign n4328 = n87 & reg_i_StoB_REQ12_out;
  assign n4329 = n87 & reg_controllable_BtoS_ACK12_out;
  assign n4330 = n4328 & ~n4329;
  assign n4331 = ~i_StoB_REQ12 & n4330;
  assign n4332 = n4327 & ~n4331;
  assign n4333 = i_StoB_REQ12 & n4329;
  assign n4334 = n4332 & ~n4333;
  assign n4335 = n87 & reg_i_StoB_REQ13_out;
  assign n4336 = n87 & reg_controllable_BtoS_ACK13_out;
  assign n4337 = n4335 & ~n4336;
  assign n4338 = ~i_StoB_REQ13 & n4337;
  assign n4339 = n4334 & ~n4338;
  assign n4340 = i_StoB_REQ13 & n4336;
  assign n4341 = n4339 & ~n4340;
  assign n4342 = n87 & reg_i_StoB_REQ14_out;
  assign n4343 = n87 & reg_controllable_BtoS_ACK14_out;
  assign n4344 = n4342 & ~n4343;
  assign n4345 = ~i_StoB_REQ14 & n4344;
  assign n4346 = n4341 & ~n4345;
  assign n4347 = i_StoB_REQ14 & n4343;
  assign n4348 = n4346 & ~n4347;
  assign n4349 = n87 & reg_controllable_BtoR_REQ0_out;
  assign n4350 = i_RtoB_ACK0 & ~n4349;
  assign n4351 = n4348 & ~n4350;
  assign n4352 = n87 & reg_i_RtoB_ACK0_out;
  assign n4353 = ~i_RtoB_ACK0 & n4352;
  assign n4354 = n4349 & n4353;
  assign n4355 = n4351 & ~n4354;
  assign n4356 = n87 & reg_controllable_BtoR_REQ1_out;
  assign n4357 = i_RtoB_ACK1 & ~n4356;
  assign n4358 = n4355 & ~n4357;
  assign n4359 = n87 & reg_i_RtoB_ACK1_out;
  assign n4360 = ~i_RtoB_ACK1 & n4359;
  assign n4361 = n4356 & n4360;
  assign n4362 = n4358 & ~n4361;
  assign n4363 = n87 & reg_controllable_DEQ_out;
  assign n4364 = n87 & reg_controllable_ENQ_out;
  assign n4365 = ~n4363 & n4364;
  assign n4366 = ~i_nEMPTY & n4365;
  assign n4367 = n4362 & ~n4366;
  assign n4368 = n4363 & ~n4364;
  assign n4369 = i_FULL & n4368;
  assign n4370 = n4367 & ~n4369;
  assign n4371 = ~n4365 & ~n4368;
  assign n4372 = n87 & reg_i_FULL_out;
  assign n4373 = i_FULL & ~n4372;
  assign n4374 = ~i_FULL & n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = n87 & reg_i_nEMPTY_out;
  assign n4377 = i_nEMPTY & ~n4376;
  assign n4378 = ~i_nEMPTY & n4376;
  assign n4379 = ~n4377 & ~n4378;
  assign n4380 = n4375 & n4379;
  assign n4381 = n4371 & ~n4380;
  assign n4382 = n4370 & ~n4381;
  assign n4383 = n87 & env_safe_err_happened_out;
  assign n4384 = n4382 & ~n4383;
  assign n4385 = ~n4151 & ~n4376;
  assign n4386 = ~n4363 & ~n4385;
  assign n4387 = n4161 & ~n4162;
  assign n4388 = n4166 & ~n4167;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390 = n4172 & ~n4173;
  assign n4391 = n4389 & ~n4390;
  assign n4392 = n4178 & ~n4179;
  assign n4393 = n4391 & ~n4392;
  assign n4394 = n4184 & ~n4185;
  assign n4395 = n4393 & ~n4394;
  assign n4396 = n4190 & ~n4191;
  assign n4397 = n4395 & ~n4396;
  assign n4398 = n4196 & ~n4197;
  assign n4399 = n4397 & ~n4398;
  assign n4400 = n4202 & ~n4203;
  assign n4401 = n4399 & ~n4400;
  assign n4402 = ~n4154 & n4157;
  assign n4403 = n4401 & ~n4402;
  assign n4404 = n4209 & ~n4210;
  assign n4405 = n4403 & ~n4404;
  assign n4406 = n4215 & ~n4216;
  assign n4407 = n4405 & ~n4406;
  assign n4408 = n4221 & ~n4222;
  assign n4409 = n4407 & ~n4408;
  assign n4410 = n4227 & ~n4228;
  assign n4411 = n4409 & ~n4410;
  assign n4412 = n4233 & ~n4234;
  assign n4413 = n4411 & ~n4412;
  assign n4414 = n4239 & ~n4240;
  assign n4415 = n4413 & ~n4414;
  assign n4416 = ~n4151 & ~n4152;
  assign n4417 = n4415 & ~n4416;
  assign n4418 = ~n4243 & n4417;
  assign n4419 = n87 & fair_cnt<2>_out ;
  assign n4420 = i_RtoB_ACK1 & ~controllable_BtoR_REQ1;
  assign n4421 = ~i_RtoB_ACK1 & controllable_BtoR_REQ1;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = n87 & env_fair1done_out;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = i_RtoB_ACK0 & ~controllable_BtoR_REQ0;
  assign n4426 = ~i_RtoB_ACK0 & controllable_BtoR_REQ0;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = n87 & env_fair0done_out;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = ~n4424 & ~n4429;
  assign n4431 = n87 & fair_cnt<0>_out ;
  assign n4432 = n4430 & n4431;
  assign n4433 = n87 & fair_cnt<1>_out ;
  assign n4434 = n4432 & n4433;
  assign n4435 = ~n4419 & ~n4434;
  assign n4436 = n4419 & n4434;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = n4418 & n4437;
  assign n4439 = ~n4432 & n4433;
  assign n4440 = n4432 & ~n4433;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = n4418 & ~n4441;
  assign n4443 = ~n4430 & ~n4431;
  assign n4444 = ~n4432 & ~n4443;
  assign n4445 = n4418 & n4444;
  assign n4446 = n87 & reg_nstateG7_1_out;
  assign n4447 = ~n4349 & n4446;
  assign n4448 = n4356 & n4447;
  assign n4449 = n4349 & ~n4446;
  assign n4450 = ~n4356 & n4449;
  assign n4451 = ~n4448 & ~n4450;
  assign n4452 = n87 & reg_stateG7_0_out;
  assign n4453 = ~n4349 & ~n4356;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = n4451 & ~n4454;
  assign n4456 = ~n4447 & ~n4449;
  assign n4457 = ~n4356 & ~n4456;
  assign n4458 = n4349 & n4446;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = n4418 & ~n4430;
  assign n4461 = ~n4429 & n4460;
  assign n4462 = ~n4217 & ~n4243;
  assign n4463 = ~n4424 & n4460;
  assign n4464 = ~n4241 & ~n4243;
  assign n4465 = ~n4163 & ~n4243;
  assign n4466 = ~n4235 & ~n4243;
  assign n4467 = ~n4229 & ~n4243;
  assign n4468 = ~n4223 & ~n4243;
  assign n4469 = ~n4211 & ~n4243;
  assign n4470 = ~n4204 & ~n4243;
  assign n4471 = ~n4198 & ~n4243;
  assign n4472 = ~n4158 & ~n4243;
  assign n4473 = ~n4192 & ~n4243;
  assign n4474 = ~n4186 & ~n4243;
  assign n4475 = ~n4180 & ~n4243;
  assign n4476 = ~n4168 & ~n4243;
  assign n4477 = ~n4174 & ~n4243;
  assign n4478 = i_StoB_REQ1 & controllable_BtoS_ACK1;
  assign n4479 = ~i_StoB_REQ2 & n4478;
  assign n4480 = ~i_StoB_REQ2 & ~n4479;
  assign n4481 = controllable_BtoS_ACK2 & ~n4480;
  assign n4482 = ~controllable_BtoS_ACK2 & n4478;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = n4477 & ~n4483;
  assign n4485 = controllable_BtoS_ACK2 & ~n4481;
  assign n4486 = ~n4477 & ~n4485;
  assign n4487 = ~n4484 & ~n4486;
  assign n4488 = n4476 & ~n4487;
  assign n4489 = ~i_StoB_REQ1 & ~controllable_BtoS_ACK1;
  assign n4490 = ~i_StoB_REQ1 & ~n4489;
  assign n4491 = ~i_StoB_REQ2 & ~n4490;
  assign n4492 = ~i_StoB_REQ2 & ~n4491;
  assign n4493 = controllable_BtoS_ACK2 & ~n4492;
  assign n4494 = ~controllable_BtoS_ACK2 & ~n4490;
  assign n4495 = ~n4493 & ~n4494;
  assign n4496 = n4477 & ~n4495;
  assign n4497 = ~n4481 & ~n4494;
  assign n4498 = ~n4477 & ~n4497;
  assign n4499 = ~n4496 & ~n4498;
  assign n4500 = ~n4476 & ~n4499;
  assign n4501 = ~n4488 & ~n4500;
  assign n4502 = ~i_StoB_REQ3 & ~n4501;
  assign n4503 = ~i_StoB_REQ3 & ~n4502;
  assign n4504 = controllable_BtoS_ACK3 & ~n4503;
  assign n4505 = ~controllable_BtoS_ACK3 & ~n4501;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = n4475 & ~n4506;
  assign n4508 = ~i_StoB_REQ3 & ~n4483;
  assign n4509 = ~i_StoB_REQ3 & ~n4508;
  assign n4510 = controllable_BtoS_ACK3 & ~n4509;
  assign n4511 = ~n4477 & ~n4486;
  assign n4512 = n4476 & ~n4511;
  assign n4513 = ~n4500 & ~n4512;
  assign n4514 = ~controllable_BtoS_ACK3 & ~n4513;
  assign n4515 = ~n4510 & ~n4514;
  assign n4516 = ~n4475 & ~n4515;
  assign n4517 = ~n4507 & ~n4516;
  assign n4518 = ~i_StoB_REQ4 & ~n4517;
  assign n4519 = ~i_StoB_REQ4 & ~n4518;
  assign n4520 = controllable_BtoS_ACK4 & ~n4519;
  assign n4521 = ~controllable_BtoS_ACK4 & ~n4517;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = n4474 & ~n4522;
  assign n4524 = ~controllable_BtoS_ACK3 & ~n4483;
  assign n4525 = ~n4510 & ~n4524;
  assign n4526 = ~i_StoB_REQ4 & ~n4525;
  assign n4527 = ~i_StoB_REQ4 & ~n4526;
  assign n4528 = controllable_BtoS_ACK4 & ~n4527;
  assign n4529 = ~i_StoB_REQ3 & ~n4513;
  assign n4530 = ~i_StoB_REQ3 & ~n4529;
  assign n4531 = controllable_BtoS_ACK3 & ~n4530;
  assign n4532 = ~n4514 & ~n4531;
  assign n4533 = n4475 & ~n4532;
  assign n4534 = ~n4516 & ~n4533;
  assign n4535 = ~controllable_BtoS_ACK4 & ~n4534;
  assign n4536 = ~n4528 & ~n4535;
  assign n4537 = ~n4474 & ~n4536;
  assign n4538 = ~n4523 & ~n4537;
  assign n4539 = ~i_StoB_REQ5 & ~n4538;
  assign n4540 = ~i_StoB_REQ5 & ~n4539;
  assign n4541 = controllable_BtoS_ACK5 & ~n4540;
  assign n4542 = ~controllable_BtoS_ACK5 & ~n4538;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = n4473 & ~n4543;
  assign n4545 = ~controllable_BtoS_ACK4 & ~n4525;
  assign n4546 = ~n4528 & ~n4545;
  assign n4547 = ~i_StoB_REQ5 & ~n4546;
  assign n4548 = ~i_StoB_REQ5 & ~n4547;
  assign n4549 = controllable_BtoS_ACK5 & ~n4548;
  assign n4550 = ~i_StoB_REQ4 & ~n4534;
  assign n4551 = ~i_StoB_REQ4 & ~n4550;
  assign n4552 = controllable_BtoS_ACK4 & ~n4551;
  assign n4553 = ~n4535 & ~n4552;
  assign n4554 = n4474 & ~n4553;
  assign n4555 = ~n4537 & ~n4554;
  assign n4556 = ~controllable_BtoS_ACK5 & ~n4555;
  assign n4557 = ~n4549 & ~n4556;
  assign n4558 = ~n4473 & ~n4557;
  assign n4559 = ~n4544 & ~n4558;
  assign n4560 = ~i_StoB_REQ8 & ~n4559;
  assign n4561 = ~i_StoB_REQ8 & ~n4560;
  assign n4562 = controllable_BtoS_ACK8 & ~n4561;
  assign n4563 = ~controllable_BtoS_ACK8 & ~n4559;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = n4472 & ~n4564;
  assign n4566 = ~controllable_BtoS_ACK5 & ~n4546;
  assign n4567 = ~n4549 & ~n4566;
  assign n4568 = ~i_StoB_REQ8 & ~n4567;
  assign n4569 = ~i_StoB_REQ8 & ~n4568;
  assign n4570 = controllable_BtoS_ACK8 & ~n4569;
  assign n4571 = ~i_StoB_REQ5 & ~n4555;
  assign n4572 = ~i_StoB_REQ5 & ~n4571;
  assign n4573 = controllable_BtoS_ACK5 & ~n4572;
  assign n4574 = ~n4556 & ~n4573;
  assign n4575 = n4473 & ~n4574;
  assign n4576 = ~n4558 & ~n4575;
  assign n4577 = ~controllable_BtoS_ACK8 & ~n4576;
  assign n4578 = ~n4570 & ~n4577;
  assign n4579 = ~n4472 & ~n4578;
  assign n4580 = ~n4565 & ~n4579;
  assign n4581 = n4471 & ~n4580;
  assign n4582 = ~controllable_BtoS_ACK8 & ~n4567;
  assign n4583 = ~n4570 & ~n4582;
  assign n4584 = ~n4471 & ~n4583;
  assign n4585 = ~n4581 & ~n4584;
  assign n4586 = ~i_StoB_REQ6 & ~n4585;
  assign n4587 = ~i_StoB_REQ6 & ~n4586;
  assign n4588 = controllable_BtoS_ACK6 & ~n4587;
  assign n4589 = ~i_StoB_REQ8 & ~n4576;
  assign n4590 = ~i_StoB_REQ8 & ~n4589;
  assign n4591 = controllable_BtoS_ACK8 & ~n4590;
  assign n4592 = ~n4577 & ~n4591;
  assign n4593 = n4472 & ~n4592;
  assign n4594 = ~n4579 & ~n4593;
  assign n4595 = ~n4471 & ~n4594;
  assign n4596 = ~n4581 & ~n4595;
  assign n4597 = ~controllable_BtoS_ACK6 & ~n4596;
  assign n4598 = ~n4588 & ~n4597;
  assign n4599 = ~i_StoB_REQ7 & ~n4598;
  assign n4600 = ~i_StoB_REQ7 & ~n4599;
  assign n4601 = controllable_BtoS_ACK7 & ~n4600;
  assign n4602 = ~controllable_BtoS_ACK7 & ~n4598;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = n4470 & ~n4603;
  assign n4605 = ~i_StoB_REQ6 & ~n4583;
  assign n4606 = ~i_StoB_REQ6 & ~n4605;
  assign n4607 = controllable_BtoS_ACK6 & ~n4606;
  assign n4608 = ~controllable_BtoS_ACK6 & ~n4583;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = ~i_StoB_REQ7 & ~n4609;
  assign n4611 = ~i_StoB_REQ7 & ~n4610;
  assign n4612 = controllable_BtoS_ACK7 & ~n4611;
  assign n4613 = n4471 & ~n4594;
  assign n4614 = ~n4584 & ~n4613;
  assign n4615 = ~i_StoB_REQ6 & ~n4614;
  assign n4616 = ~i_StoB_REQ6 & ~n4615;
  assign n4617 = controllable_BtoS_ACK6 & ~n4616;
  assign n4618 = ~controllable_BtoS_ACK6 & ~n4594;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~controllable_BtoS_ACK7 & ~n4619;
  assign n4621 = ~n4612 & ~n4620;
  assign n4622 = ~n4470 & ~n4621;
  assign n4623 = ~n4604 & ~n4622;
  assign n4624 = n4469 & ~n4623;
  assign n4625 = ~controllable_BtoS_ACK7 & ~n4609;
  assign n4626 = ~n4612 & ~n4625;
  assign n4627 = ~n4469 & ~n4626;
  assign n4628 = ~n4624 & ~n4627;
  assign n4629 = ~i_StoB_REQ9 & ~n4628;
  assign n4630 = ~i_StoB_REQ9 & ~n4629;
  assign n4631 = controllable_BtoS_ACK9 & ~n4630;
  assign n4632 = ~i_StoB_REQ7 & ~n4619;
  assign n4633 = ~i_StoB_REQ7 & ~n4632;
  assign n4634 = controllable_BtoS_ACK7 & ~n4633;
  assign n4635 = ~n4620 & ~n4634;
  assign n4636 = n4470 & ~n4635;
  assign n4637 = ~n4622 & ~n4636;
  assign n4638 = ~n4469 & ~n4637;
  assign n4639 = ~n4624 & ~n4638;
  assign n4640 = ~controllable_BtoS_ACK9 & ~n4639;
  assign n4641 = ~n4631 & ~n4640;
  assign n4642 = n4468 & ~n4641;
  assign n4643 = ~i_StoB_REQ9 & ~n4626;
  assign n4644 = ~i_StoB_REQ9 & ~n4643;
  assign n4645 = controllable_BtoS_ACK9 & ~n4644;
  assign n4646 = ~controllable_BtoS_ACK9 & ~n4626;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~n4468 & ~n4647;
  assign n4649 = ~n4642 & ~n4648;
  assign n4650 = ~i_StoB_REQ11 & ~n4649;
  assign n4651 = ~i_StoB_REQ11 & ~n4650;
  assign n4652 = controllable_BtoS_ACK11 & ~n4651;
  assign n4653 = n4469 & ~n4637;
  assign n4654 = ~n4627 & ~n4653;
  assign n4655 = ~i_StoB_REQ9 & ~n4654;
  assign n4656 = ~i_StoB_REQ9 & ~n4655;
  assign n4657 = controllable_BtoS_ACK9 & ~n4656;
  assign n4658 = ~controllable_BtoS_ACK9 & ~n4637;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n4468 & ~n4659;
  assign n4661 = ~n4642 & ~n4660;
  assign n4662 = ~controllable_BtoS_ACK11 & ~n4661;
  assign n4663 = ~n4652 & ~n4662;
  assign n4664 = n4467 & ~n4663;
  assign n4665 = ~i_StoB_REQ11 & ~n4647;
  assign n4666 = ~i_StoB_REQ11 & ~n4665;
  assign n4667 = controllable_BtoS_ACK11 & ~n4666;
  assign n4668 = ~controllable_BtoS_ACK11 & ~n4647;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = ~n4467 & ~n4669;
  assign n4671 = ~n4664 & ~n4670;
  assign n4672 = ~i_StoB_REQ12 & ~n4671;
  assign n4673 = ~i_StoB_REQ12 & ~n4672;
  assign n4674 = controllable_BtoS_ACK12 & ~n4673;
  assign n4675 = n4468 & ~n4659;
  assign n4676 = ~n4648 & ~n4675;
  assign n4677 = ~i_StoB_REQ11 & ~n4676;
  assign n4678 = ~i_StoB_REQ11 & ~n4677;
  assign n4679 = controllable_BtoS_ACK11 & ~n4678;
  assign n4680 = ~controllable_BtoS_ACK11 & ~n4659;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = ~n4467 & ~n4681;
  assign n4683 = ~n4664 & ~n4682;
  assign n4684 = ~controllable_BtoS_ACK12 & ~n4683;
  assign n4685 = ~n4674 & ~n4684;
  assign n4686 = ~controllable_BtoS_ACK13 & ~n4685;
  assign n4687 = ~controllable_BtoS_ACK13 & ~n4686;
  assign n4688 = i_StoB_REQ13 & ~n4687;
  assign n4689 = i_StoB_REQ1 & ~n4478;
  assign n4690 = ~i_StoB_REQ2 & ~n4689;
  assign n4691 = ~i_StoB_REQ2 & ~n4690;
  assign n4692 = controllable_BtoS_ACK2 & ~n4691;
  assign n4693 = i_StoB_REQ2 & n4478;
  assign n4694 = ~n4690 & ~n4693;
  assign n4695 = ~controllable_BtoS_ACK2 & ~n4694;
  assign n4696 = ~n4692 & ~n4695;
  assign n4697 = n4477 & ~n4696;
  assign n4698 = controllable_BtoS_ACK2 & ~n4692;
  assign n4699 = ~n4477 & ~n4698;
  assign n4700 = ~n4697 & ~n4699;
  assign n4701 = n4476 & ~n4700;
  assign n4702 = i_StoB_REQ2 & ~n4490;
  assign n4703 = i_StoB_REQ2 & ~n4702;
  assign n4704 = ~controllable_BtoS_ACK2 & ~n4703;
  assign n4705 = ~controllable_BtoS_ACK2 & ~n4704;
  assign n4706 = n4477 & ~n4705;
  assign n4707 = ~n4692 & ~n4704;
  assign n4708 = ~n4477 & ~n4707;
  assign n4709 = ~n4706 & ~n4708;
  assign n4710 = ~n4476 & ~n4709;
  assign n4711 = ~n4701 & ~n4710;
  assign n4712 = ~i_StoB_REQ3 & ~n4711;
  assign n4713 = ~i_StoB_REQ3 & ~n4712;
  assign n4714 = controllable_BtoS_ACK3 & ~n4713;
  assign n4715 = i_StoB_REQ3 & ~n4501;
  assign n4716 = ~n4712 & ~n4715;
  assign n4717 = ~controllable_BtoS_ACK3 & ~n4716;
  assign n4718 = ~n4714 & ~n4717;
  assign n4719 = n4475 & ~n4718;
  assign n4720 = ~i_StoB_REQ3 & ~n4696;
  assign n4721 = ~i_StoB_REQ3 & ~n4720;
  assign n4722 = controllable_BtoS_ACK3 & ~n4721;
  assign n4723 = i_StoB_REQ3 & ~n4513;
  assign n4724 = ~n4477 & ~n4699;
  assign n4725 = n4476 & ~n4724;
  assign n4726 = ~n4710 & ~n4725;
  assign n4727 = ~i_StoB_REQ3 & ~n4726;
  assign n4728 = ~n4723 & ~n4727;
  assign n4729 = ~controllable_BtoS_ACK3 & ~n4728;
  assign n4730 = ~n4722 & ~n4729;
  assign n4731 = ~n4475 & ~n4730;
  assign n4732 = ~n4719 & ~n4731;
  assign n4733 = ~i_StoB_REQ4 & ~n4732;
  assign n4734 = ~i_StoB_REQ4 & ~n4733;
  assign n4735 = controllable_BtoS_ACK4 & ~n4734;
  assign n4736 = i_StoB_REQ4 & ~n4517;
  assign n4737 = ~n4733 & ~n4736;
  assign n4738 = ~controllable_BtoS_ACK4 & ~n4737;
  assign n4739 = ~n4735 & ~n4738;
  assign n4740 = n4474 & ~n4739;
  assign n4741 = i_StoB_REQ3 & ~n4483;
  assign n4742 = ~n4720 & ~n4741;
  assign n4743 = ~controllable_BtoS_ACK3 & ~n4742;
  assign n4744 = ~n4722 & ~n4743;
  assign n4745 = ~i_StoB_REQ4 & ~n4744;
  assign n4746 = ~i_StoB_REQ4 & ~n4745;
  assign n4747 = controllable_BtoS_ACK4 & ~n4746;
  assign n4748 = i_StoB_REQ4 & ~n4534;
  assign n4749 = ~i_StoB_REQ3 & ~n4727;
  assign n4750 = controllable_BtoS_ACK3 & ~n4749;
  assign n4751 = ~n4729 & ~n4750;
  assign n4752 = n4475 & ~n4751;
  assign n4753 = ~n4731 & ~n4752;
  assign n4754 = ~i_StoB_REQ4 & ~n4753;
  assign n4755 = ~n4748 & ~n4754;
  assign n4756 = ~controllable_BtoS_ACK4 & ~n4755;
  assign n4757 = ~n4747 & ~n4756;
  assign n4758 = ~n4474 & ~n4757;
  assign n4759 = ~n4740 & ~n4758;
  assign n4760 = ~i_StoB_REQ5 & ~n4759;
  assign n4761 = ~i_StoB_REQ5 & ~n4760;
  assign n4762 = controllable_BtoS_ACK5 & ~n4761;
  assign n4763 = i_StoB_REQ5 & ~n4538;
  assign n4764 = ~n4760 & ~n4763;
  assign n4765 = ~controllable_BtoS_ACK5 & ~n4764;
  assign n4766 = ~n4762 & ~n4765;
  assign n4767 = n4473 & ~n4766;
  assign n4768 = i_StoB_REQ4 & ~n4525;
  assign n4769 = ~n4745 & ~n4768;
  assign n4770 = ~controllable_BtoS_ACK4 & ~n4769;
  assign n4771 = ~n4747 & ~n4770;
  assign n4772 = ~i_StoB_REQ5 & ~n4771;
  assign n4773 = ~i_StoB_REQ5 & ~n4772;
  assign n4774 = controllable_BtoS_ACK5 & ~n4773;
  assign n4775 = i_StoB_REQ5 & ~n4555;
  assign n4776 = ~i_StoB_REQ4 & ~n4754;
  assign n4777 = controllable_BtoS_ACK4 & ~n4776;
  assign n4778 = ~n4756 & ~n4777;
  assign n4779 = n4474 & ~n4778;
  assign n4780 = ~n4758 & ~n4779;
  assign n4781 = ~i_StoB_REQ5 & ~n4780;
  assign n4782 = ~n4775 & ~n4781;
  assign n4783 = ~controllable_BtoS_ACK5 & ~n4782;
  assign n4784 = ~n4774 & ~n4783;
  assign n4785 = ~n4473 & ~n4784;
  assign n4786 = ~n4767 & ~n4785;
  assign n4787 = ~i_StoB_REQ8 & ~n4786;
  assign n4788 = ~i_StoB_REQ8 & ~n4787;
  assign n4789 = controllable_BtoS_ACK8 & ~n4788;
  assign n4790 = i_StoB_REQ8 & ~n4559;
  assign n4791 = ~n4787 & ~n4790;
  assign n4792 = ~controllable_BtoS_ACK8 & ~n4791;
  assign n4793 = ~n4789 & ~n4792;
  assign n4794 = n4472 & ~n4793;
  assign n4795 = i_StoB_REQ5 & ~n4546;
  assign n4796 = ~n4772 & ~n4795;
  assign n4797 = ~controllable_BtoS_ACK5 & ~n4796;
  assign n4798 = ~n4774 & ~n4797;
  assign n4799 = ~i_StoB_REQ8 & ~n4798;
  assign n4800 = ~i_StoB_REQ8 & ~n4799;
  assign n4801 = controllable_BtoS_ACK8 & ~n4800;
  assign n4802 = i_StoB_REQ8 & ~n4576;
  assign n4803 = ~i_StoB_REQ5 & ~n4781;
  assign n4804 = controllable_BtoS_ACK5 & ~n4803;
  assign n4805 = ~n4783 & ~n4804;
  assign n4806 = n4473 & ~n4805;
  assign n4807 = ~n4785 & ~n4806;
  assign n4808 = ~i_StoB_REQ8 & ~n4807;
  assign n4809 = ~n4802 & ~n4808;
  assign n4810 = ~controllable_BtoS_ACK8 & ~n4809;
  assign n4811 = ~n4801 & ~n4810;
  assign n4812 = ~n4472 & ~n4811;
  assign n4813 = ~n4794 & ~n4812;
  assign n4814 = n4471 & ~n4813;
  assign n4815 = i_StoB_REQ8 & ~n4567;
  assign n4816 = ~n4799 & ~n4815;
  assign n4817 = ~controllable_BtoS_ACK8 & ~n4816;
  assign n4818 = ~n4801 & ~n4817;
  assign n4819 = ~n4471 & ~n4818;
  assign n4820 = ~n4814 & ~n4819;
  assign n4821 = ~i_StoB_REQ6 & ~n4820;
  assign n4822 = ~i_StoB_REQ6 & ~n4821;
  assign n4823 = controllable_BtoS_ACK6 & ~n4822;
  assign n4824 = i_StoB_REQ6 & ~n4596;
  assign n4825 = ~i_StoB_REQ8 & ~n4808;
  assign n4826 = controllable_BtoS_ACK8 & ~n4825;
  assign n4827 = ~n4810 & ~n4826;
  assign n4828 = n4472 & ~n4827;
  assign n4829 = ~n4812 & ~n4828;
  assign n4830 = ~n4471 & ~n4829;
  assign n4831 = ~n4814 & ~n4830;
  assign n4832 = ~i_StoB_REQ6 & ~n4831;
  assign n4833 = ~n4824 & ~n4832;
  assign n4834 = ~controllable_BtoS_ACK6 & ~n4833;
  assign n4835 = ~n4823 & ~n4834;
  assign n4836 = ~i_StoB_REQ7 & ~n4835;
  assign n4837 = ~i_StoB_REQ7 & ~n4836;
  assign n4838 = controllable_BtoS_ACK7 & ~n4837;
  assign n4839 = i_StoB_REQ7 & ~n4598;
  assign n4840 = ~n4836 & ~n4839;
  assign n4841 = ~controllable_BtoS_ACK7 & ~n4840;
  assign n4842 = ~n4838 & ~n4841;
  assign n4843 = n4470 & ~n4842;
  assign n4844 = ~i_StoB_REQ6 & ~n4818;
  assign n4845 = ~i_StoB_REQ6 & ~n4844;
  assign n4846 = controllable_BtoS_ACK6 & ~n4845;
  assign n4847 = i_StoB_REQ6 & ~n4583;
  assign n4848 = ~n4844 & ~n4847;
  assign n4849 = ~controllable_BtoS_ACK6 & ~n4848;
  assign n4850 = ~n4846 & ~n4849;
  assign n4851 = ~i_StoB_REQ7 & ~n4850;
  assign n4852 = ~i_StoB_REQ7 & ~n4851;
  assign n4853 = controllable_BtoS_ACK7 & ~n4852;
  assign n4854 = i_StoB_REQ7 & ~n4619;
  assign n4855 = n4471 & ~n4829;
  assign n4856 = ~n4819 & ~n4855;
  assign n4857 = ~i_StoB_REQ6 & ~n4856;
  assign n4858 = ~i_StoB_REQ6 & ~n4857;
  assign n4859 = controllable_BtoS_ACK6 & ~n4858;
  assign n4860 = i_StoB_REQ6 & ~n4594;
  assign n4861 = ~i_StoB_REQ6 & ~n4829;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~controllable_BtoS_ACK6 & ~n4862;
  assign n4864 = ~n4859 & ~n4863;
  assign n4865 = ~i_StoB_REQ7 & ~n4864;
  assign n4866 = ~n4854 & ~n4865;
  assign n4867 = ~controllable_BtoS_ACK7 & ~n4866;
  assign n4868 = ~n4853 & ~n4867;
  assign n4869 = ~n4470 & ~n4868;
  assign n4870 = ~n4843 & ~n4869;
  assign n4871 = n4469 & ~n4870;
  assign n4872 = i_StoB_REQ7 & ~n4609;
  assign n4873 = ~n4851 & ~n4872;
  assign n4874 = ~controllable_BtoS_ACK7 & ~n4873;
  assign n4875 = ~n4853 & ~n4874;
  assign n4876 = ~n4469 & ~n4875;
  assign n4877 = ~n4871 & ~n4876;
  assign n4878 = ~i_StoB_REQ9 & ~n4877;
  assign n4879 = ~i_StoB_REQ9 & ~n4878;
  assign n4880 = controllable_BtoS_ACK9 & ~n4879;
  assign n4881 = i_StoB_REQ9 & ~n4639;
  assign n4882 = ~i_StoB_REQ7 & ~n4865;
  assign n4883 = controllable_BtoS_ACK7 & ~n4882;
  assign n4884 = ~n4867 & ~n4883;
  assign n4885 = n4470 & ~n4884;
  assign n4886 = ~n4869 & ~n4885;
  assign n4887 = ~n4469 & ~n4886;
  assign n4888 = ~n4871 & ~n4887;
  assign n4889 = ~i_StoB_REQ9 & ~n4888;
  assign n4890 = ~n4881 & ~n4889;
  assign n4891 = ~controllable_BtoS_ACK9 & ~n4890;
  assign n4892 = ~n4880 & ~n4891;
  assign n4893 = n4468 & ~n4892;
  assign n4894 = ~i_StoB_REQ9 & ~n4875;
  assign n4895 = ~i_StoB_REQ9 & ~n4894;
  assign n4896 = controllable_BtoS_ACK9 & ~n4895;
  assign n4897 = i_StoB_REQ9 & ~n4626;
  assign n4898 = ~n4894 & ~n4897;
  assign n4899 = ~controllable_BtoS_ACK9 & ~n4898;
  assign n4900 = ~n4896 & ~n4899;
  assign n4901 = ~n4468 & ~n4900;
  assign n4902 = ~n4893 & ~n4901;
  assign n4903 = ~i_StoB_REQ11 & ~n4902;
  assign n4904 = ~i_StoB_REQ11 & ~n4903;
  assign n4905 = controllable_BtoS_ACK11 & ~n4904;
  assign n4906 = i_StoB_REQ11 & ~n4661;
  assign n4907 = n4469 & ~n4886;
  assign n4908 = ~n4876 & ~n4907;
  assign n4909 = ~i_StoB_REQ9 & ~n4908;
  assign n4910 = ~i_StoB_REQ9 & ~n4909;
  assign n4911 = controllable_BtoS_ACK9 & ~n4910;
  assign n4912 = i_StoB_REQ9 & ~n4637;
  assign n4913 = ~i_StoB_REQ9 & ~n4886;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = ~controllable_BtoS_ACK9 & ~n4914;
  assign n4916 = ~n4911 & ~n4915;
  assign n4917 = ~n4468 & ~n4916;
  assign n4918 = ~n4893 & ~n4917;
  assign n4919 = ~i_StoB_REQ11 & ~n4918;
  assign n4920 = ~n4906 & ~n4919;
  assign n4921 = ~controllable_BtoS_ACK11 & ~n4920;
  assign n4922 = ~n4905 & ~n4921;
  assign n4923 = n4467 & ~n4922;
  assign n4924 = ~i_StoB_REQ11 & ~n4900;
  assign n4925 = ~i_StoB_REQ11 & ~n4924;
  assign n4926 = controllable_BtoS_ACK11 & ~n4925;
  assign n4927 = i_StoB_REQ11 & ~n4647;
  assign n4928 = ~n4924 & ~n4927;
  assign n4929 = ~controllable_BtoS_ACK11 & ~n4928;
  assign n4930 = ~n4926 & ~n4929;
  assign n4931 = ~n4467 & ~n4930;
  assign n4932 = ~n4923 & ~n4931;
  assign n4933 = ~i_StoB_REQ12 & ~n4932;
  assign n4934 = ~i_StoB_REQ12 & ~n4933;
  assign n4935 = controllable_BtoS_ACK12 & ~n4934;
  assign n4936 = i_StoB_REQ12 & ~n4683;
  assign n4937 = n4468 & ~n4916;
  assign n4938 = ~n4901 & ~n4937;
  assign n4939 = ~i_StoB_REQ11 & ~n4938;
  assign n4940 = ~i_StoB_REQ11 & ~n4939;
  assign n4941 = controllable_BtoS_ACK11 & ~n4940;
  assign n4942 = i_StoB_REQ11 & ~n4659;
  assign n4943 = ~i_StoB_REQ11 & ~n4916;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~controllable_BtoS_ACK11 & ~n4944;
  assign n4946 = ~n4941 & ~n4945;
  assign n4947 = ~n4467 & ~n4946;
  assign n4948 = ~n4923 & ~n4947;
  assign n4949 = ~i_StoB_REQ12 & ~n4948;
  assign n4950 = ~n4936 & ~n4949;
  assign n4951 = ~controllable_BtoS_ACK12 & ~n4950;
  assign n4952 = ~n4935 & ~n4951;
  assign n4953 = ~i_StoB_REQ13 & ~n4952;
  assign n4954 = ~n4688 & ~n4953;
  assign n4955 = n4466 & ~n4954;
  assign n4956 = n4467 & ~n4681;
  assign n4957 = ~n4670 & ~n4956;
  assign n4958 = ~i_StoB_REQ12 & ~n4957;
  assign n4959 = ~i_StoB_REQ12 & ~n4958;
  assign n4960 = controllable_BtoS_ACK12 & ~n4959;
  assign n4961 = ~controllable_BtoS_ACK12 & ~n4681;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~controllable_BtoS_ACK13 & ~n4962;
  assign n4964 = ~controllable_BtoS_ACK13 & ~n4963;
  assign n4965 = i_StoB_REQ13 & ~n4964;
  assign n4966 = ~i_StoB_REQ12 & ~n4930;
  assign n4967 = ~i_StoB_REQ12 & ~n4966;
  assign n4968 = controllable_BtoS_ACK12 & ~n4967;
  assign n4969 = i_StoB_REQ12 & ~n4669;
  assign n4970 = ~n4966 & ~n4969;
  assign n4971 = ~controllable_BtoS_ACK12 & ~n4970;
  assign n4972 = ~n4968 & ~n4971;
  assign n4973 = controllable_BtoS_ACK13 & ~n4972;
  assign n4974 = n4467 & ~n4946;
  assign n4975 = ~n4931 & ~n4974;
  assign n4976 = ~i_StoB_REQ12 & ~n4975;
  assign n4977 = ~i_StoB_REQ12 & ~n4976;
  assign n4978 = controllable_BtoS_ACK12 & ~n4977;
  assign n4979 = i_StoB_REQ12 & ~n4681;
  assign n4980 = ~i_StoB_REQ12 & ~n4946;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = ~controllable_BtoS_ACK12 & ~n4981;
  assign n4983 = ~n4978 & ~n4982;
  assign n4984 = ~controllable_BtoS_ACK13 & ~n4983;
  assign n4985 = ~n4973 & ~n4984;
  assign n4986 = ~i_StoB_REQ13 & ~n4985;
  assign n4987 = ~n4965 & ~n4986;
  assign n4988 = ~n4466 & ~n4987;
  assign n4989 = ~n4955 & ~n4988;
  assign n4990 = ~i_StoB_REQ0 & ~n4989;
  assign n4991 = ~i_StoB_REQ0 & ~n4990;
  assign n4992 = ~i_StoB_REQ14 & ~n4991;
  assign n4993 = ~i_StoB_REQ14 & ~n4992;
  assign n4994 = controllable_BtoS_ACK14 & ~n4993;
  assign n4995 = ~i_StoB_REQ13 & ~n4685;
  assign n4996 = ~n4688 & ~n4995;
  assign n4997 = n4466 & ~n4996;
  assign n4998 = ~i_StoB_REQ12 & ~n4669;
  assign n4999 = ~i_StoB_REQ12 & ~n4998;
  assign n5000 = controllable_BtoS_ACK12 & ~n4999;
  assign n5001 = ~controllable_BtoS_ACK12 & ~n4669;
  assign n5002 = ~n5000 & ~n5001;
  assign n5003 = controllable_BtoS_ACK13 & ~n5002;
  assign n5004 = ~n4963 & ~n5003;
  assign n5005 = ~i_StoB_REQ13 & ~n5004;
  assign n5006 = ~n4965 & ~n5005;
  assign n5007 = ~n4466 & ~n5006;
  assign n5008 = ~n4997 & ~n5007;
  assign n5009 = ~i_StoB_REQ0 & ~n5008;
  assign n5010 = ~i_StoB_REQ0 & ~n5009;
  assign n5011 = i_StoB_REQ14 & ~n5010;
  assign n5012 = ~n4992 & ~n5011;
  assign n5013 = ~controllable_BtoS_ACK14 & ~n5012;
  assign n5014 = ~n4994 & ~n5013;
  assign n5015 = controllable_ENQ & ~n5014;
  assign n5016 = controllable_ENQ & ~n5015;
  assign n5017 = ~i_RtoB_ACK1 & ~n5016;
  assign n5018 = ~i_RtoB_ACK1 & ~n5017;
  assign n5019 = controllable_BtoR_REQ1 & ~n5018;
  assign n5020 = ~i_StoB_REQ14 & ~n5010;
  assign n5021 = ~i_StoB_REQ14 & ~n5020;
  assign n5022 = controllable_BtoS_ACK14 & ~n5021;
  assign n5023 = ~controllable_BtoS_ACK14 & ~n5010;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = controllable_ENQ & ~n5024;
  assign n5026 = controllable_ENQ & ~n5025;
  assign n5027 = ~controllable_BtoR_REQ1 & ~n5026;
  assign n5028 = ~n5019 & ~n5027;
  assign n5029 = ~controllable_BtoR_REQ0 & ~n5028;
  assign n5030 = ~controllable_BtoR_REQ0 & ~n5029;
  assign n5031 = i_RtoB_ACK0 & ~n5030;
  assign n5032 = i_RtoB_ACK1 & ~n5026;
  assign n5033 = ~controllable_ENQ & ~n5014;
  assign n5034 = ~n5025 & ~n5033;
  assign n5035 = ~i_RtoB_ACK1 & ~n5034;
  assign n5036 = ~n5032 & ~n5035;
  assign n5037 = controllable_BtoR_REQ1 & ~n5036;
  assign n5038 = ~i_RtoB_ACK1 & ~n5024;
  assign n5039 = ~n5032 & ~n5038;
  assign n5040 = ~controllable_BtoR_REQ1 & ~n5039;
  assign n5041 = ~n5037 & ~n5040;
  assign n5042 = ~controllable_BtoR_REQ0 & ~n5041;
  assign n5043 = ~controllable_BtoR_REQ0 & ~n5042;
  assign n5044 = ~i_RtoB_ACK0 & ~n5043;
  assign n5045 = ~n5031 & ~n5044;
  assign n5046 = controllable_DEQ & ~n5045;
  assign n5047 = ~i_RtoB_ACK1 & ~n5014;
  assign n5048 = ~i_RtoB_ACK1 & ~n5047;
  assign n5049 = controllable_BtoR_REQ1 & ~n5048;
  assign n5050 = ~controllable_BtoR_REQ1 & ~n5024;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = ~controllable_BtoR_REQ0 & ~n5051;
  assign n5053 = ~controllable_BtoR_REQ0 & ~n5052;
  assign n5054 = i_RtoB_ACK0 & ~n5053;
  assign n5055 = ~controllable_BtoR_REQ0 & ~n5024;
  assign n5056 = ~controllable_BtoR_REQ0 & ~n5055;
  assign n5057 = ~i_RtoB_ACK0 & ~n5056;
  assign n5058 = ~n5054 & ~n5057;
  assign n5059 = ~controllable_DEQ & ~n5058;
  assign n5060 = ~n5046 & ~n5059;
  assign n5061 = i_nEMPTY & ~n5060;
  assign n5062 = ~controllable_ENQ & ~n5033;
  assign n5063 = ~i_RtoB_ACK1 & ~n5062;
  assign n5064 = ~i_RtoB_ACK1 & ~n5063;
  assign n5065 = controllable_BtoR_REQ1 & ~n5064;
  assign n5066 = ~controllable_ENQ & ~n5024;
  assign n5067 = ~controllable_ENQ & ~n5066;
  assign n5068 = ~i_RtoB_ACK1 & ~n5067;
  assign n5069 = ~i_RtoB_ACK1 & ~n5068;
  assign n5070 = ~controllable_BtoR_REQ1 & ~n5069;
  assign n5071 = ~n5065 & ~n5070;
  assign n5072 = ~controllable_BtoR_REQ0 & ~n5071;
  assign n5073 = ~controllable_BtoR_REQ0 & ~n5072;
  assign n5074 = ~i_RtoB_ACK0 & ~n5073;
  assign n5075 = ~i_RtoB_ACK0 & ~n5074;
  assign n5076 = controllable_DEQ & ~n5075;
  assign n5077 = ~controllable_BtoR_REQ0 & ~n5026;
  assign n5078 = ~controllable_BtoR_REQ0 & ~n5077;
  assign n5079 = ~i_RtoB_ACK0 & ~n5078;
  assign n5080 = ~n5031 & ~n5079;
  assign n5081 = ~controllable_DEQ & ~n5080;
  assign n5082 = ~n5076 & ~n5081;
  assign n5083 = i_FULL & ~n5082;
  assign n5084 = ~i_RtoB_ACK1 & ~n5038;
  assign n5085 = ~controllable_BtoR_REQ1 & ~n5084;
  assign n5086 = ~n5049 & ~n5085;
  assign n5087 = ~controllable_BtoR_REQ0 & ~n5086;
  assign n5088 = ~controllable_BtoR_REQ0 & ~n5087;
  assign n5089 = ~i_RtoB_ACK0 & ~n5088;
  assign n5090 = ~i_RtoB_ACK0 & ~n5089;
  assign n5091 = controllable_DEQ & ~n5090;
  assign n5092 = ~controllable_BtoR_REQ0 & ~n5036;
  assign n5093 = ~controllable_BtoR_REQ0 & ~n5092;
  assign n5094 = ~i_RtoB_ACK0 & ~n5093;
  assign n5095 = ~n5031 & ~n5094;
  assign n5096 = ~controllable_DEQ & ~n5095;
  assign n5097 = ~n5091 & ~n5096;
  assign n5098 = ~i_FULL & ~n5097;
  assign n5099 = ~n5083 & ~n5098;
  assign n5100 = ~i_nEMPTY & ~n5099;
  assign n5101 = ~n5061 & ~n5100;
  assign n5102 = controllable_BtoS_ACK0 & ~n5101;
  assign n5103 = i_StoB_REQ0 & ~n5008;
  assign n5104 = ~n4990 & ~n5103;
  assign n5105 = ~i_StoB_REQ14 & ~n5104;
  assign n5106 = ~i_StoB_REQ14 & ~n5105;
  assign n5107 = controllable_BtoS_ACK14 & ~n5106;
  assign n5108 = i_StoB_REQ14 & ~n5008;
  assign n5109 = ~n5105 & ~n5108;
  assign n5110 = ~controllable_BtoS_ACK14 & ~n5109;
  assign n5111 = ~n5107 & ~n5110;
  assign n5112 = controllable_ENQ & ~n5111;
  assign n5113 = controllable_ENQ & ~n5112;
  assign n5114 = ~i_RtoB_ACK1 & ~n5113;
  assign n5115 = ~i_RtoB_ACK1 & ~n5114;
  assign n5116 = controllable_BtoR_REQ1 & ~n5115;
  assign n5117 = ~i_StoB_REQ14 & ~n5008;
  assign n5118 = ~i_StoB_REQ14 & ~n5117;
  assign n5119 = controllable_BtoS_ACK14 & ~n5118;
  assign n5120 = ~controllable_BtoS_ACK14 & ~n5008;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = controllable_ENQ & ~n5121;
  assign n5123 = controllable_ENQ & ~n5122;
  assign n5124 = ~controllable_BtoR_REQ1 & ~n5123;
  assign n5125 = ~n5116 & ~n5124;
  assign n5126 = ~controllable_BtoR_REQ0 & ~n5125;
  assign n5127 = ~controllable_BtoR_REQ0 & ~n5126;
  assign n5128 = i_RtoB_ACK0 & ~n5127;
  assign n5129 = i_RtoB_ACK1 & ~n5123;
  assign n5130 = ~controllable_ENQ & ~n5111;
  assign n5131 = ~n5122 & ~n5130;
  assign n5132 = ~i_RtoB_ACK1 & ~n5131;
  assign n5133 = ~n5129 & ~n5132;
  assign n5134 = controllable_BtoR_REQ1 & ~n5133;
  assign n5135 = ~i_RtoB_ACK1 & ~n5121;
  assign n5136 = ~n5129 & ~n5135;
  assign n5137 = ~controllable_BtoR_REQ1 & ~n5136;
  assign n5138 = ~n5134 & ~n5137;
  assign n5139 = ~controllable_BtoR_REQ0 & ~n5138;
  assign n5140 = ~controllable_BtoR_REQ0 & ~n5139;
  assign n5141 = ~i_RtoB_ACK0 & ~n5140;
  assign n5142 = ~n5128 & ~n5141;
  assign n5143 = controllable_DEQ & ~n5142;
  assign n5144 = ~i_RtoB_ACK1 & ~n5111;
  assign n5145 = ~i_RtoB_ACK1 & ~n5144;
  assign n5146 = controllable_BtoR_REQ1 & ~n5145;
  assign n5147 = ~controllable_BtoR_REQ1 & ~n5121;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = ~controllable_BtoR_REQ0 & ~n5148;
  assign n5150 = ~controllable_BtoR_REQ0 & ~n5149;
  assign n5151 = i_RtoB_ACK0 & ~n5150;
  assign n5152 = ~controllable_BtoR_REQ0 & ~n5121;
  assign n5153 = ~controllable_BtoR_REQ0 & ~n5152;
  assign n5154 = ~i_RtoB_ACK0 & ~n5153;
  assign n5155 = ~n5151 & ~n5154;
  assign n5156 = ~controllable_DEQ & ~n5155;
  assign n5157 = ~n5143 & ~n5156;
  assign n5158 = i_nEMPTY & ~n5157;
  assign n5159 = ~controllable_ENQ & ~n5130;
  assign n5160 = ~i_RtoB_ACK1 & ~n5159;
  assign n5161 = ~i_RtoB_ACK1 & ~n5160;
  assign n5162 = controllable_BtoR_REQ1 & ~n5161;
  assign n5163 = ~controllable_ENQ & ~n5121;
  assign n5164 = ~controllable_ENQ & ~n5163;
  assign n5165 = ~i_RtoB_ACK1 & ~n5164;
  assign n5166 = ~i_RtoB_ACK1 & ~n5165;
  assign n5167 = ~controllable_BtoR_REQ1 & ~n5166;
  assign n5168 = ~n5162 & ~n5167;
  assign n5169 = ~controllable_BtoR_REQ0 & ~n5168;
  assign n5170 = ~controllable_BtoR_REQ0 & ~n5169;
  assign n5171 = ~i_RtoB_ACK0 & ~n5170;
  assign n5172 = ~i_RtoB_ACK0 & ~n5171;
  assign n5173 = controllable_DEQ & ~n5172;
  assign n5174 = ~controllable_BtoR_REQ0 & ~n5123;
  assign n5175 = ~controllable_BtoR_REQ0 & ~n5174;
  assign n5176 = ~i_RtoB_ACK0 & ~n5175;
  assign n5177 = ~n5128 & ~n5176;
  assign n5178 = ~controllable_DEQ & ~n5177;
  assign n5179 = ~n5173 & ~n5178;
  assign n5180 = i_FULL & ~n5179;
  assign n5181 = ~i_RtoB_ACK1 & ~n5135;
  assign n5182 = ~controllable_BtoR_REQ1 & ~n5181;
  assign n5183 = ~n5146 & ~n5182;
  assign n5184 = ~controllable_BtoR_REQ0 & ~n5183;
  assign n5185 = ~controllable_BtoR_REQ0 & ~n5184;
  assign n5186 = ~i_RtoB_ACK0 & ~n5185;
  assign n5187 = ~i_RtoB_ACK0 & ~n5186;
  assign n5188 = controllable_DEQ & ~n5187;
  assign n5189 = ~controllable_BtoR_REQ0 & ~n5133;
  assign n5190 = ~controllable_BtoR_REQ0 & ~n5189;
  assign n5191 = ~i_RtoB_ACK0 & ~n5190;
  assign n5192 = ~n5128 & ~n5191;
  assign n5193 = ~controllable_DEQ & ~n5192;
  assign n5194 = ~n5188 & ~n5193;
  assign n5195 = ~i_FULL & ~n5194;
  assign n5196 = ~n5180 & ~n5195;
  assign n5197 = ~i_nEMPTY & ~n5196;
  assign n5198 = ~n5158 & ~n5197;
  assign n5199 = ~controllable_BtoS_ACK0 & ~n5198;
  assign n5200 = ~n5102 & ~n5199;
  assign n5201 = n4465 & ~n5200;
  assign n5202 = ~controllable_BtoS_ACK13 & ~n5002;
  assign n5203 = ~controllable_BtoS_ACK13 & ~n5202;
  assign n5204 = i_StoB_REQ13 & ~n5203;
  assign n5205 = ~i_StoB_REQ13 & ~n4972;
  assign n5206 = ~n5204 & ~n5205;
  assign n5207 = ~i_StoB_REQ0 & ~n5206;
  assign n5208 = ~i_StoB_REQ0 & ~n5207;
  assign n5209 = ~i_StoB_REQ14 & ~n5208;
  assign n5210 = ~i_StoB_REQ14 & ~n5209;
  assign n5211 = controllable_BtoS_ACK14 & ~n5210;
  assign n5212 = ~i_StoB_REQ13 & ~n5002;
  assign n5213 = ~n5204 & ~n5212;
  assign n5214 = ~i_StoB_REQ0 & ~n5213;
  assign n5215 = ~i_StoB_REQ0 & ~n5214;
  assign n5216 = i_StoB_REQ14 & ~n5215;
  assign n5217 = ~n5209 & ~n5216;
  assign n5218 = ~controllable_BtoS_ACK14 & ~n5217;
  assign n5219 = ~n5211 & ~n5218;
  assign n5220 = controllable_ENQ & ~n5219;
  assign n5221 = controllable_ENQ & ~n5220;
  assign n5222 = ~i_RtoB_ACK1 & ~n5221;
  assign n5223 = ~i_RtoB_ACK1 & ~n5222;
  assign n5224 = controllable_BtoR_REQ1 & ~n5223;
  assign n5225 = ~i_StoB_REQ14 & ~n5215;
  assign n5226 = ~i_StoB_REQ14 & ~n5225;
  assign n5227 = controllable_BtoS_ACK14 & ~n5226;
  assign n5228 = ~controllable_BtoS_ACK14 & ~n5215;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = controllable_ENQ & ~n5229;
  assign n5231 = controllable_ENQ & ~n5230;
  assign n5232 = ~controllable_BtoR_REQ1 & ~n5231;
  assign n5233 = ~n5224 & ~n5232;
  assign n5234 = ~controllable_BtoR_REQ0 & ~n5233;
  assign n5235 = ~controllable_BtoR_REQ0 & ~n5234;
  assign n5236 = i_RtoB_ACK0 & ~n5235;
  assign n5237 = i_RtoB_ACK1 & ~n5231;
  assign n5238 = ~controllable_ENQ & ~n5219;
  assign n5239 = ~n5230 & ~n5238;
  assign n5240 = ~i_RtoB_ACK1 & ~n5239;
  assign n5241 = ~n5237 & ~n5240;
  assign n5242 = controllable_BtoR_REQ1 & ~n5241;
  assign n5243 = ~i_RtoB_ACK1 & ~n5229;
  assign n5244 = ~n5237 & ~n5243;
  assign n5245 = ~controllable_BtoR_REQ1 & ~n5244;
  assign n5246 = ~n5242 & ~n5245;
  assign n5247 = ~controllable_BtoR_REQ0 & ~n5246;
  assign n5248 = ~controllable_BtoR_REQ0 & ~n5247;
  assign n5249 = ~i_RtoB_ACK0 & ~n5248;
  assign n5250 = ~n5236 & ~n5249;
  assign n5251 = controllable_DEQ & ~n5250;
  assign n5252 = ~i_RtoB_ACK1 & ~n5219;
  assign n5253 = ~i_RtoB_ACK1 & ~n5252;
  assign n5254 = controllable_BtoR_REQ1 & ~n5253;
  assign n5255 = ~controllable_BtoR_REQ1 & ~n5229;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = ~controllable_BtoR_REQ0 & ~n5256;
  assign n5258 = ~controllable_BtoR_REQ0 & ~n5257;
  assign n5259 = i_RtoB_ACK0 & ~n5258;
  assign n5260 = ~controllable_BtoR_REQ0 & ~n5229;
  assign n5261 = ~controllable_BtoR_REQ0 & ~n5260;
  assign n5262 = ~i_RtoB_ACK0 & ~n5261;
  assign n5263 = ~n5259 & ~n5262;
  assign n5264 = ~controllable_DEQ & ~n5263;
  assign n5265 = ~n5251 & ~n5264;
  assign n5266 = i_nEMPTY & ~n5265;
  assign n5267 = ~controllable_ENQ & ~n5238;
  assign n5268 = ~i_RtoB_ACK1 & ~n5267;
  assign n5269 = ~i_RtoB_ACK1 & ~n5268;
  assign n5270 = controllable_BtoR_REQ1 & ~n5269;
  assign n5271 = ~controllable_ENQ & ~n5229;
  assign n5272 = ~controllable_ENQ & ~n5271;
  assign n5273 = ~i_RtoB_ACK1 & ~n5272;
  assign n5274 = ~i_RtoB_ACK1 & ~n5273;
  assign n5275 = ~controllable_BtoR_REQ1 & ~n5274;
  assign n5276 = ~n5270 & ~n5275;
  assign n5277 = ~controllable_BtoR_REQ0 & ~n5276;
  assign n5278 = ~controllable_BtoR_REQ0 & ~n5277;
  assign n5279 = ~i_RtoB_ACK0 & ~n5278;
  assign n5280 = ~i_RtoB_ACK0 & ~n5279;
  assign n5281 = controllable_DEQ & ~n5280;
  assign n5282 = ~controllable_BtoR_REQ0 & ~n5231;
  assign n5283 = ~controllable_BtoR_REQ0 & ~n5282;
  assign n5284 = ~i_RtoB_ACK0 & ~n5283;
  assign n5285 = ~n5236 & ~n5284;
  assign n5286 = ~controllable_DEQ & ~n5285;
  assign n5287 = ~n5281 & ~n5286;
  assign n5288 = i_FULL & ~n5287;
  assign n5289 = ~i_RtoB_ACK1 & ~n5243;
  assign n5290 = ~controllable_BtoR_REQ1 & ~n5289;
  assign n5291 = ~n5254 & ~n5290;
  assign n5292 = ~controllable_BtoR_REQ0 & ~n5291;
  assign n5293 = ~controllable_BtoR_REQ0 & ~n5292;
  assign n5294 = ~i_RtoB_ACK0 & ~n5293;
  assign n5295 = ~i_RtoB_ACK0 & ~n5294;
  assign n5296 = controllable_DEQ & ~n5295;
  assign n5297 = ~controllable_BtoR_REQ0 & ~n5241;
  assign n5298 = ~controllable_BtoR_REQ0 & ~n5297;
  assign n5299 = ~i_RtoB_ACK0 & ~n5298;
  assign n5300 = ~n5236 & ~n5299;
  assign n5301 = ~controllable_DEQ & ~n5300;
  assign n5302 = ~n5296 & ~n5301;
  assign n5303 = ~i_FULL & ~n5302;
  assign n5304 = ~n5288 & ~n5303;
  assign n5305 = ~i_nEMPTY & ~n5304;
  assign n5306 = ~n5266 & ~n5305;
  assign n5307 = controllable_BtoS_ACK0 & ~n5306;
  assign n5308 = ~i_StoB_REQ13 & ~n4962;
  assign n5309 = ~n4965 & ~n5308;
  assign n5310 = n4466 & ~n5309;
  assign n5311 = ~n5007 & ~n5310;
  assign n5312 = i_StoB_REQ0 & ~n5311;
  assign n5313 = ~i_StoB_REQ13 & ~n4983;
  assign n5314 = ~n4965 & ~n5313;
  assign n5315 = n4466 & ~n5314;
  assign n5316 = ~n4988 & ~n5315;
  assign n5317 = ~i_StoB_REQ0 & ~n5316;
  assign n5318 = ~n5312 & ~n5317;
  assign n5319 = ~i_StoB_REQ14 & ~n5318;
  assign n5320 = ~i_StoB_REQ14 & ~n5319;
  assign n5321 = controllable_BtoS_ACK14 & ~n5320;
  assign n5322 = i_StoB_REQ14 & ~n5311;
  assign n5323 = ~n5319 & ~n5322;
  assign n5324 = ~controllable_BtoS_ACK14 & ~n5323;
  assign n5325 = ~n5321 & ~n5324;
  assign n5326 = controllable_ENQ & ~n5325;
  assign n5327 = controllable_ENQ & ~n5326;
  assign n5328 = ~i_RtoB_ACK1 & ~n5327;
  assign n5329 = ~i_RtoB_ACK1 & ~n5328;
  assign n5330 = controllable_BtoR_REQ1 & ~n5329;
  assign n5331 = ~i_StoB_REQ14 & ~n5311;
  assign n5332 = ~i_StoB_REQ14 & ~n5331;
  assign n5333 = controllable_BtoS_ACK14 & ~n5332;
  assign n5334 = ~controllable_BtoS_ACK14 & ~n5311;
  assign n5335 = ~n5333 & ~n5334;
  assign n5336 = controllable_ENQ & ~n5335;
  assign n5337 = controllable_ENQ & ~n5336;
  assign n5338 = ~controllable_BtoR_REQ1 & ~n5337;
  assign n5339 = ~n5330 & ~n5338;
  assign n5340 = ~controllable_BtoR_REQ0 & ~n5339;
  assign n5341 = ~controllable_BtoR_REQ0 & ~n5340;
  assign n5342 = i_RtoB_ACK0 & ~n5341;
  assign n5343 = i_RtoB_ACK1 & ~n5337;
  assign n5344 = ~controllable_ENQ & ~n5325;
  assign n5345 = ~n5336 & ~n5344;
  assign n5346 = ~i_RtoB_ACK1 & ~n5345;
  assign n5347 = ~n5343 & ~n5346;
  assign n5348 = controllable_BtoR_REQ1 & ~n5347;
  assign n5349 = ~i_RtoB_ACK1 & ~n5335;
  assign n5350 = ~n5343 & ~n5349;
  assign n5351 = ~controllable_BtoR_REQ1 & ~n5350;
  assign n5352 = ~n5348 & ~n5351;
  assign n5353 = ~controllable_BtoR_REQ0 & ~n5352;
  assign n5354 = ~controllable_BtoR_REQ0 & ~n5353;
  assign n5355 = ~i_RtoB_ACK0 & ~n5354;
  assign n5356 = ~n5342 & ~n5355;
  assign n5357 = controllable_DEQ & ~n5356;
  assign n5358 = ~i_RtoB_ACK1 & ~n5325;
  assign n5359 = ~i_RtoB_ACK1 & ~n5358;
  assign n5360 = controllable_BtoR_REQ1 & ~n5359;
  assign n5361 = ~controllable_BtoR_REQ1 & ~n5335;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = ~controllable_BtoR_REQ0 & ~n5362;
  assign n5364 = ~controllable_BtoR_REQ0 & ~n5363;
  assign n5365 = i_RtoB_ACK0 & ~n5364;
  assign n5366 = ~controllable_BtoR_REQ0 & ~n5335;
  assign n5367 = ~controllable_BtoR_REQ0 & ~n5366;
  assign n5368 = ~i_RtoB_ACK0 & ~n5367;
  assign n5369 = ~n5365 & ~n5368;
  assign n5370 = ~controllable_DEQ & ~n5369;
  assign n5371 = ~n5357 & ~n5370;
  assign n5372 = i_nEMPTY & ~n5371;
  assign n5373 = ~controllable_ENQ & ~n5344;
  assign n5374 = ~i_RtoB_ACK1 & ~n5373;
  assign n5375 = ~i_RtoB_ACK1 & ~n5374;
  assign n5376 = controllable_BtoR_REQ1 & ~n5375;
  assign n5377 = ~controllable_ENQ & ~n5335;
  assign n5378 = ~controllable_ENQ & ~n5377;
  assign n5379 = ~i_RtoB_ACK1 & ~n5378;
  assign n5380 = ~i_RtoB_ACK1 & ~n5379;
  assign n5381 = ~controllable_BtoR_REQ1 & ~n5380;
  assign n5382 = ~n5376 & ~n5381;
  assign n5383 = ~controllable_BtoR_REQ0 & ~n5382;
  assign n5384 = ~controllable_BtoR_REQ0 & ~n5383;
  assign n5385 = ~i_RtoB_ACK0 & ~n5384;
  assign n5386 = ~i_RtoB_ACK0 & ~n5385;
  assign n5387 = controllable_DEQ & ~n5386;
  assign n5388 = ~controllable_BtoR_REQ0 & ~n5337;
  assign n5389 = ~controllable_BtoR_REQ0 & ~n5388;
  assign n5390 = ~i_RtoB_ACK0 & ~n5389;
  assign n5391 = ~n5342 & ~n5390;
  assign n5392 = ~controllable_DEQ & ~n5391;
  assign n5393 = ~n5387 & ~n5392;
  assign n5394 = i_FULL & ~n5393;
  assign n5395 = ~i_RtoB_ACK1 & ~n5349;
  assign n5396 = ~controllable_BtoR_REQ1 & ~n5395;
  assign n5397 = ~n5360 & ~n5396;
  assign n5398 = ~controllable_BtoR_REQ0 & ~n5397;
  assign n5399 = ~controllable_BtoR_REQ0 & ~n5398;
  assign n5400 = ~i_RtoB_ACK0 & ~n5399;
  assign n5401 = ~i_RtoB_ACK0 & ~n5400;
  assign n5402 = controllable_DEQ & ~n5401;
  assign n5403 = ~controllable_BtoR_REQ0 & ~n5347;
  assign n5404 = ~controllable_BtoR_REQ0 & ~n5403;
  assign n5405 = ~i_RtoB_ACK0 & ~n5404;
  assign n5406 = ~n5342 & ~n5405;
  assign n5407 = ~controllable_DEQ & ~n5406;
  assign n5408 = ~n5402 & ~n5407;
  assign n5409 = ~i_FULL & ~n5408;
  assign n5410 = ~n5394 & ~n5409;
  assign n5411 = ~i_nEMPTY & ~n5410;
  assign n5412 = ~n5372 & ~n5411;
  assign n5413 = ~controllable_BtoS_ACK0 & ~n5412;
  assign n5414 = ~n5307 & ~n5413;
  assign n5415 = ~n4465 & ~n5414;
  assign n5416 = ~n5201 & ~n5415;
  assign n5417 = i_StoB_REQ10 & ~n5416;
  assign n5418 = i_StoB_REQ2 & ~n4693;
  assign n5419 = ~controllable_BtoS_ACK2 & ~n5418;
  assign n5420 = ~n4481 & ~n5419;
  assign n5421 = ~n4477 & ~n5420;
  assign n5422 = ~n4484 & ~n5421;
  assign n5423 = n4476 & ~n5422;
  assign n5424 = ~n4478 & ~n4489;
  assign n5425 = ~i_StoB_REQ2 & ~n5424;
  assign n5426 = ~i_StoB_REQ2 & ~n5425;
  assign n5427 = controllable_BtoS_ACK2 & ~n5426;
  assign n5428 = ~controllable_BtoS_ACK2 & ~n5424;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = n4477 & ~n5429;
  assign n5431 = ~n4693 & ~n5425;
  assign n5432 = ~controllable_BtoS_ACK2 & ~n5431;
  assign n5433 = ~n4481 & ~n5432;
  assign n5434 = ~n4477 & ~n5433;
  assign n5435 = ~n5430 & ~n5434;
  assign n5436 = ~n4476 & ~n5435;
  assign n5437 = ~n5423 & ~n5436;
  assign n5438 = ~i_StoB_REQ3 & ~n5437;
  assign n5439 = ~i_StoB_REQ3 & ~n5438;
  assign n5440 = controllable_BtoS_ACK3 & ~n5439;
  assign n5441 = ~controllable_BtoS_ACK3 & ~n5437;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = n4475 & ~n5442;
  assign n5444 = ~n4477 & ~n5421;
  assign n5445 = n4476 & ~n5444;
  assign n5446 = ~n5436 & ~n5445;
  assign n5447 = ~i_StoB_REQ3 & ~n5446;
  assign n5448 = ~n4741 & ~n5447;
  assign n5449 = ~controllable_BtoS_ACK3 & ~n5448;
  assign n5450 = ~n4510 & ~n5449;
  assign n5451 = ~n4475 & ~n5450;
  assign n5452 = ~n5443 & ~n5451;
  assign n5453 = ~i_StoB_REQ4 & ~n5452;
  assign n5454 = ~i_StoB_REQ4 & ~n5453;
  assign n5455 = controllable_BtoS_ACK4 & ~n5454;
  assign n5456 = ~controllable_BtoS_ACK4 & ~n5452;
  assign n5457 = ~n5455 & ~n5456;
  assign n5458 = n4474 & ~n5457;
  assign n5459 = ~i_StoB_REQ3 & ~n5447;
  assign n5460 = controllable_BtoS_ACK3 & ~n5459;
  assign n5461 = ~controllable_BtoS_ACK3 & ~n5446;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n4475 & ~n5462;
  assign n5464 = ~n5451 & ~n5463;
  assign n5465 = ~i_StoB_REQ4 & ~n5464;
  assign n5466 = ~n4768 & ~n5465;
  assign n5467 = ~controllable_BtoS_ACK4 & ~n5466;
  assign n5468 = ~n4528 & ~n5467;
  assign n5469 = ~n4474 & ~n5468;
  assign n5470 = ~n5458 & ~n5469;
  assign n5471 = ~i_StoB_REQ5 & ~n5470;
  assign n5472 = ~i_StoB_REQ5 & ~n5471;
  assign n5473 = controllable_BtoS_ACK5 & ~n5472;
  assign n5474 = ~controllable_BtoS_ACK5 & ~n5470;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = n4473 & ~n5475;
  assign n5477 = ~i_StoB_REQ4 & ~n5465;
  assign n5478 = controllable_BtoS_ACK4 & ~n5477;
  assign n5479 = ~controllable_BtoS_ACK4 & ~n5464;
  assign n5480 = ~n5478 & ~n5479;
  assign n5481 = n4474 & ~n5480;
  assign n5482 = ~n5469 & ~n5481;
  assign n5483 = ~i_StoB_REQ5 & ~n5482;
  assign n5484 = ~n4795 & ~n5483;
  assign n5485 = ~controllable_BtoS_ACK5 & ~n5484;
  assign n5486 = ~n4549 & ~n5485;
  assign n5487 = ~n4473 & ~n5486;
  assign n5488 = ~n5476 & ~n5487;
  assign n5489 = ~i_StoB_REQ8 & ~n5488;
  assign n5490 = ~i_StoB_REQ8 & ~n5489;
  assign n5491 = controllable_BtoS_ACK8 & ~n5490;
  assign n5492 = ~controllable_BtoS_ACK8 & ~n5488;
  assign n5493 = ~n5491 & ~n5492;
  assign n5494 = n4472 & ~n5493;
  assign n5495 = ~i_StoB_REQ5 & ~n5483;
  assign n5496 = controllable_BtoS_ACK5 & ~n5495;
  assign n5497 = ~controllable_BtoS_ACK5 & ~n5482;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = n4473 & ~n5498;
  assign n5500 = ~n5487 & ~n5499;
  assign n5501 = ~i_StoB_REQ8 & ~n5500;
  assign n5502 = ~n4815 & ~n5501;
  assign n5503 = ~controllable_BtoS_ACK8 & ~n5502;
  assign n5504 = ~n4570 & ~n5503;
  assign n5505 = ~n4472 & ~n5504;
  assign n5506 = ~n5494 & ~n5505;
  assign n5507 = n4471 & ~n5506;
  assign n5508 = ~n4584 & ~n5507;
  assign n5509 = ~i_StoB_REQ6 & ~n5508;
  assign n5510 = ~i_StoB_REQ6 & ~n5509;
  assign n5511 = controllable_BtoS_ACK6 & ~n5510;
  assign n5512 = i_StoB_REQ6 & ~n5508;
  assign n5513 = ~i_StoB_REQ8 & ~n5501;
  assign n5514 = controllable_BtoS_ACK8 & ~n5513;
  assign n5515 = ~controllable_BtoS_ACK8 & ~n5500;
  assign n5516 = ~n5514 & ~n5515;
  assign n5517 = n4472 & ~n5516;
  assign n5518 = ~n5505 & ~n5517;
  assign n5519 = ~n4471 & ~n5518;
  assign n5520 = ~n5507 & ~n5519;
  assign n5521 = ~i_StoB_REQ6 & ~n5520;
  assign n5522 = ~n5512 & ~n5521;
  assign n5523 = ~controllable_BtoS_ACK6 & ~n5522;
  assign n5524 = ~n5511 & ~n5523;
  assign n5525 = ~i_StoB_REQ7 & ~n5524;
  assign n5526 = ~i_StoB_REQ7 & ~n5525;
  assign n5527 = controllable_BtoS_ACK7 & ~n5526;
  assign n5528 = ~controllable_BtoS_ACK7 & ~n5524;
  assign n5529 = ~n5527 & ~n5528;
  assign n5530 = n4470 & ~n5529;
  assign n5531 = n4471 & ~n5518;
  assign n5532 = ~n4584 & ~n5531;
  assign n5533 = ~i_StoB_REQ6 & ~n5532;
  assign n5534 = ~i_StoB_REQ6 & ~n5533;
  assign n5535 = controllable_BtoS_ACK6 & ~n5534;
  assign n5536 = i_StoB_REQ6 & ~n5532;
  assign n5537 = ~i_StoB_REQ6 & ~n5518;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~controllable_BtoS_ACK6 & ~n5538;
  assign n5540 = ~n5535 & ~n5539;
  assign n5541 = ~i_StoB_REQ7 & ~n5540;
  assign n5542 = ~n4872 & ~n5541;
  assign n5543 = ~controllable_BtoS_ACK7 & ~n5542;
  assign n5544 = ~n4612 & ~n5543;
  assign n5545 = ~n4470 & ~n5544;
  assign n5546 = ~n5530 & ~n5545;
  assign n5547 = n4469 & ~n5546;
  assign n5548 = ~n4627 & ~n5547;
  assign n5549 = ~i_StoB_REQ9 & ~n5548;
  assign n5550 = ~i_StoB_REQ9 & ~n5549;
  assign n5551 = controllable_BtoS_ACK9 & ~n5550;
  assign n5552 = i_StoB_REQ9 & ~n5548;
  assign n5553 = ~i_StoB_REQ7 & ~n5541;
  assign n5554 = controllable_BtoS_ACK7 & ~n5553;
  assign n5555 = ~controllable_BtoS_ACK7 & ~n5540;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = n4470 & ~n5556;
  assign n5558 = ~n5545 & ~n5557;
  assign n5559 = ~n4469 & ~n5558;
  assign n5560 = ~n5547 & ~n5559;
  assign n5561 = ~i_StoB_REQ9 & ~n5560;
  assign n5562 = ~n5552 & ~n5561;
  assign n5563 = ~controllable_BtoS_ACK9 & ~n5562;
  assign n5564 = ~n5551 & ~n5563;
  assign n5565 = n4468 & ~n5564;
  assign n5566 = ~n4648 & ~n5565;
  assign n5567 = ~i_StoB_REQ11 & ~n5566;
  assign n5568 = ~i_StoB_REQ11 & ~n5567;
  assign n5569 = controllable_BtoS_ACK11 & ~n5568;
  assign n5570 = i_StoB_REQ11 & ~n5566;
  assign n5571 = n4469 & ~n5558;
  assign n5572 = ~n4627 & ~n5571;
  assign n5573 = ~i_StoB_REQ9 & ~n5572;
  assign n5574 = ~i_StoB_REQ9 & ~n5573;
  assign n5575 = controllable_BtoS_ACK9 & ~n5574;
  assign n5576 = i_StoB_REQ9 & ~n5572;
  assign n5577 = ~i_StoB_REQ9 & ~n5558;
  assign n5578 = ~n5576 & ~n5577;
  assign n5579 = ~controllable_BtoS_ACK9 & ~n5578;
  assign n5580 = ~n5575 & ~n5579;
  assign n5581 = ~n4468 & ~n5580;
  assign n5582 = ~n5565 & ~n5581;
  assign n5583 = ~i_StoB_REQ11 & ~n5582;
  assign n5584 = ~n5570 & ~n5583;
  assign n5585 = ~controllable_BtoS_ACK11 & ~n5584;
  assign n5586 = ~n5569 & ~n5585;
  assign n5587 = n4467 & ~n5586;
  assign n5588 = ~n4670 & ~n5587;
  assign n5589 = ~i_StoB_REQ12 & ~n5588;
  assign n5590 = ~i_StoB_REQ12 & ~n5589;
  assign n5591 = controllable_BtoS_ACK12 & ~n5590;
  assign n5592 = i_StoB_REQ12 & ~n5588;
  assign n5593 = n4468 & ~n5580;
  assign n5594 = ~n4648 & ~n5593;
  assign n5595 = ~i_StoB_REQ11 & ~n5594;
  assign n5596 = ~i_StoB_REQ11 & ~n5595;
  assign n5597 = controllable_BtoS_ACK11 & ~n5596;
  assign n5598 = i_StoB_REQ11 & ~n5594;
  assign n5599 = ~i_StoB_REQ11 & ~n5580;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = ~controllable_BtoS_ACK11 & ~n5600;
  assign n5602 = ~n5597 & ~n5601;
  assign n5603 = ~n4467 & ~n5602;
  assign n5604 = ~n5587 & ~n5603;
  assign n5605 = ~i_StoB_REQ12 & ~n5604;
  assign n5606 = ~n5592 & ~n5605;
  assign n5607 = ~controllable_BtoS_ACK12 & ~n5606;
  assign n5608 = ~n5591 & ~n5607;
  assign n5609 = ~controllable_BtoS_ACK13 & ~n5608;
  assign n5610 = ~controllable_BtoS_ACK13 & ~n5609;
  assign n5611 = i_StoB_REQ13 & ~n5610;
  assign n5612 = ~n4692 & ~n5419;
  assign n5613 = ~n4477 & ~n5612;
  assign n5614 = ~n4697 & ~n5613;
  assign n5615 = n4476 & ~n5614;
  assign n5616 = i_StoB_REQ2 & ~n5424;
  assign n5617 = ~n4690 & ~n5616;
  assign n5618 = ~controllable_BtoS_ACK2 & ~n5617;
  assign n5619 = ~n4692 & ~n5618;
  assign n5620 = n4477 & ~n5619;
  assign n5621 = ~n4477 & ~n4696;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~n4476 & ~n5622;
  assign n5624 = ~n5615 & ~n5623;
  assign n5625 = ~i_StoB_REQ3 & ~n5624;
  assign n5626 = ~i_StoB_REQ3 & ~n5625;
  assign n5627 = controllable_BtoS_ACK3 & ~n5626;
  assign n5628 = i_StoB_REQ3 & ~n5437;
  assign n5629 = ~n5625 & ~n5628;
  assign n5630 = ~controllable_BtoS_ACK3 & ~n5629;
  assign n5631 = ~n5627 & ~n5630;
  assign n5632 = n4475 & ~n5631;
  assign n5633 = ~n4477 & ~n5613;
  assign n5634 = n4476 & ~n5633;
  assign n5635 = ~n5623 & ~n5634;
  assign n5636 = ~i_StoB_REQ3 & ~n5635;
  assign n5637 = ~n4741 & ~n5636;
  assign n5638 = ~controllable_BtoS_ACK3 & ~n5637;
  assign n5639 = ~n4722 & ~n5638;
  assign n5640 = ~n4475 & ~n5639;
  assign n5641 = ~n5632 & ~n5640;
  assign n5642 = ~i_StoB_REQ4 & ~n5641;
  assign n5643 = ~i_StoB_REQ4 & ~n5642;
  assign n5644 = controllable_BtoS_ACK4 & ~n5643;
  assign n5645 = i_StoB_REQ4 & ~n5452;
  assign n5646 = ~n5642 & ~n5645;
  assign n5647 = ~controllable_BtoS_ACK4 & ~n5646;
  assign n5648 = ~n5644 & ~n5647;
  assign n5649 = n4474 & ~n5648;
  assign n5650 = ~i_StoB_REQ3 & ~n5636;
  assign n5651 = controllable_BtoS_ACK3 & ~n5650;
  assign n5652 = i_StoB_REQ3 & ~n5446;
  assign n5653 = ~n5636 & ~n5652;
  assign n5654 = ~controllable_BtoS_ACK3 & ~n5653;
  assign n5655 = ~n5651 & ~n5654;
  assign n5656 = n4475 & ~n5655;
  assign n5657 = ~n5640 & ~n5656;
  assign n5658 = ~i_StoB_REQ4 & ~n5657;
  assign n5659 = ~n4768 & ~n5658;
  assign n5660 = ~controllable_BtoS_ACK4 & ~n5659;
  assign n5661 = ~n4747 & ~n5660;
  assign n5662 = ~n4474 & ~n5661;
  assign n5663 = ~n5649 & ~n5662;
  assign n5664 = ~i_StoB_REQ5 & ~n5663;
  assign n5665 = ~i_StoB_REQ5 & ~n5664;
  assign n5666 = controllable_BtoS_ACK5 & ~n5665;
  assign n5667 = i_StoB_REQ5 & ~n5470;
  assign n5668 = ~n5664 & ~n5667;
  assign n5669 = ~controllable_BtoS_ACK5 & ~n5668;
  assign n5670 = ~n5666 & ~n5669;
  assign n5671 = n4473 & ~n5670;
  assign n5672 = ~i_StoB_REQ4 & ~n5658;
  assign n5673 = controllable_BtoS_ACK4 & ~n5672;
  assign n5674 = i_StoB_REQ4 & ~n5464;
  assign n5675 = ~n5658 & ~n5674;
  assign n5676 = ~controllable_BtoS_ACK4 & ~n5675;
  assign n5677 = ~n5673 & ~n5676;
  assign n5678 = n4474 & ~n5677;
  assign n5679 = ~n5662 & ~n5678;
  assign n5680 = ~i_StoB_REQ5 & ~n5679;
  assign n5681 = ~n4795 & ~n5680;
  assign n5682 = ~controllable_BtoS_ACK5 & ~n5681;
  assign n5683 = ~n4774 & ~n5682;
  assign n5684 = ~n4473 & ~n5683;
  assign n5685 = ~n5671 & ~n5684;
  assign n5686 = ~i_StoB_REQ8 & ~n5685;
  assign n5687 = ~i_StoB_REQ8 & ~n5686;
  assign n5688 = controllable_BtoS_ACK8 & ~n5687;
  assign n5689 = i_StoB_REQ8 & ~n5488;
  assign n5690 = ~n5686 & ~n5689;
  assign n5691 = ~controllable_BtoS_ACK8 & ~n5690;
  assign n5692 = ~n5688 & ~n5691;
  assign n5693 = n4472 & ~n5692;
  assign n5694 = ~i_StoB_REQ5 & ~n5680;
  assign n5695 = controllable_BtoS_ACK5 & ~n5694;
  assign n5696 = i_StoB_REQ5 & ~n5482;
  assign n5697 = ~n5680 & ~n5696;
  assign n5698 = ~controllable_BtoS_ACK5 & ~n5697;
  assign n5699 = ~n5695 & ~n5698;
  assign n5700 = n4473 & ~n5699;
  assign n5701 = ~n5684 & ~n5700;
  assign n5702 = ~i_StoB_REQ8 & ~n5701;
  assign n5703 = ~n4815 & ~n5702;
  assign n5704 = ~controllable_BtoS_ACK8 & ~n5703;
  assign n5705 = ~n4801 & ~n5704;
  assign n5706 = ~n4472 & ~n5705;
  assign n5707 = ~n5693 & ~n5706;
  assign n5708 = n4471 & ~n5707;
  assign n5709 = ~n4819 & ~n5708;
  assign n5710 = ~i_StoB_REQ6 & ~n5709;
  assign n5711 = ~i_StoB_REQ6 & ~n5710;
  assign n5712 = controllable_BtoS_ACK6 & ~n5711;
  assign n5713 = ~i_StoB_REQ8 & ~n5702;
  assign n5714 = controllable_BtoS_ACK8 & ~n5713;
  assign n5715 = i_StoB_REQ8 & ~n5500;
  assign n5716 = ~n5702 & ~n5715;
  assign n5717 = ~controllable_BtoS_ACK8 & ~n5716;
  assign n5718 = ~n5714 & ~n5717;
  assign n5719 = n4472 & ~n5718;
  assign n5720 = ~n5706 & ~n5719;
  assign n5721 = ~n4471 & ~n5720;
  assign n5722 = ~n5708 & ~n5721;
  assign n5723 = ~i_StoB_REQ6 & ~n5722;
  assign n5724 = ~n5512 & ~n5723;
  assign n5725 = ~controllable_BtoS_ACK6 & ~n5724;
  assign n5726 = ~n5712 & ~n5725;
  assign n5727 = ~i_StoB_REQ7 & ~n5726;
  assign n5728 = ~i_StoB_REQ7 & ~n5727;
  assign n5729 = controllable_BtoS_ACK7 & ~n5728;
  assign n5730 = i_StoB_REQ7 & ~n5524;
  assign n5731 = ~n5727 & ~n5730;
  assign n5732 = ~controllable_BtoS_ACK7 & ~n5731;
  assign n5733 = ~n5729 & ~n5732;
  assign n5734 = n4470 & ~n5733;
  assign n5735 = n4471 & ~n5720;
  assign n5736 = ~n4819 & ~n5735;
  assign n5737 = ~i_StoB_REQ6 & ~n5736;
  assign n5738 = ~i_StoB_REQ6 & ~n5737;
  assign n5739 = controllable_BtoS_ACK6 & ~n5738;
  assign n5740 = ~i_StoB_REQ6 & ~n5720;
  assign n5741 = ~n5536 & ~n5740;
  assign n5742 = ~controllable_BtoS_ACK6 & ~n5741;
  assign n5743 = ~n5739 & ~n5742;
  assign n5744 = ~i_StoB_REQ7 & ~n5743;
  assign n5745 = ~n4872 & ~n5744;
  assign n5746 = ~controllable_BtoS_ACK7 & ~n5745;
  assign n5747 = ~n4853 & ~n5746;
  assign n5748 = ~n4470 & ~n5747;
  assign n5749 = ~n5734 & ~n5748;
  assign n5750 = n4469 & ~n5749;
  assign n5751 = ~n4876 & ~n5750;
  assign n5752 = ~i_StoB_REQ9 & ~n5751;
  assign n5753 = ~i_StoB_REQ9 & ~n5752;
  assign n5754 = controllable_BtoS_ACK9 & ~n5753;
  assign n5755 = ~i_StoB_REQ7 & ~n5744;
  assign n5756 = controllable_BtoS_ACK7 & ~n5755;
  assign n5757 = i_StoB_REQ7 & ~n5540;
  assign n5758 = ~n5744 & ~n5757;
  assign n5759 = ~controllable_BtoS_ACK7 & ~n5758;
  assign n5760 = ~n5756 & ~n5759;
  assign n5761 = n4470 & ~n5760;
  assign n5762 = ~n5748 & ~n5761;
  assign n5763 = ~n4469 & ~n5762;
  assign n5764 = ~n5750 & ~n5763;
  assign n5765 = ~i_StoB_REQ9 & ~n5764;
  assign n5766 = ~n5552 & ~n5765;
  assign n5767 = ~controllable_BtoS_ACK9 & ~n5766;
  assign n5768 = ~n5754 & ~n5767;
  assign n5769 = n4468 & ~n5768;
  assign n5770 = ~n4901 & ~n5769;
  assign n5771 = ~i_StoB_REQ11 & ~n5770;
  assign n5772 = ~i_StoB_REQ11 & ~n5771;
  assign n5773 = controllable_BtoS_ACK11 & ~n5772;
  assign n5774 = n4469 & ~n5762;
  assign n5775 = ~n4876 & ~n5774;
  assign n5776 = ~i_StoB_REQ9 & ~n5775;
  assign n5777 = ~i_StoB_REQ9 & ~n5776;
  assign n5778 = controllable_BtoS_ACK9 & ~n5777;
  assign n5779 = ~i_StoB_REQ9 & ~n5762;
  assign n5780 = ~n5576 & ~n5779;
  assign n5781 = ~controllable_BtoS_ACK9 & ~n5780;
  assign n5782 = ~n5778 & ~n5781;
  assign n5783 = ~n4468 & ~n5782;
  assign n5784 = ~n5769 & ~n5783;
  assign n5785 = ~i_StoB_REQ11 & ~n5784;
  assign n5786 = ~n5570 & ~n5785;
  assign n5787 = ~controllable_BtoS_ACK11 & ~n5786;
  assign n5788 = ~n5773 & ~n5787;
  assign n5789 = n4467 & ~n5788;
  assign n5790 = ~n4931 & ~n5789;
  assign n5791 = ~i_StoB_REQ12 & ~n5790;
  assign n5792 = ~i_StoB_REQ12 & ~n5791;
  assign n5793 = controllable_BtoS_ACK12 & ~n5792;
  assign n5794 = n4468 & ~n5782;
  assign n5795 = ~n4901 & ~n5794;
  assign n5796 = ~i_StoB_REQ11 & ~n5795;
  assign n5797 = ~i_StoB_REQ11 & ~n5796;
  assign n5798 = controllable_BtoS_ACK11 & ~n5797;
  assign n5799 = ~i_StoB_REQ11 & ~n5782;
  assign n5800 = ~n5598 & ~n5799;
  assign n5801 = ~controllable_BtoS_ACK11 & ~n5800;
  assign n5802 = ~n5798 & ~n5801;
  assign n5803 = ~n4467 & ~n5802;
  assign n5804 = ~n5789 & ~n5803;
  assign n5805 = ~i_StoB_REQ12 & ~n5804;
  assign n5806 = ~n5592 & ~n5805;
  assign n5807 = ~controllable_BtoS_ACK12 & ~n5806;
  assign n5808 = ~n5793 & ~n5807;
  assign n5809 = ~i_StoB_REQ13 & ~n5808;
  assign n5810 = ~n5611 & ~n5809;
  assign n5811 = n4466 & ~n5810;
  assign n5812 = n4467 & ~n5802;
  assign n5813 = ~n4931 & ~n5812;
  assign n5814 = ~i_StoB_REQ12 & ~n5813;
  assign n5815 = ~i_StoB_REQ12 & ~n5814;
  assign n5816 = controllable_BtoS_ACK12 & ~n5815;
  assign n5817 = n4467 & ~n5602;
  assign n5818 = ~n4670 & ~n5817;
  assign n5819 = i_StoB_REQ12 & ~n5818;
  assign n5820 = ~i_StoB_REQ12 & ~n5802;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = ~controllable_BtoS_ACK12 & ~n5821;
  assign n5823 = ~n5816 & ~n5822;
  assign n5824 = ~controllable_BtoS_ACK13 & ~n5823;
  assign n5825 = ~n4973 & ~n5824;
  assign n5826 = ~i_StoB_REQ13 & ~n5825;
  assign n5827 = ~n5204 & ~n5826;
  assign n5828 = ~n4466 & ~n5827;
  assign n5829 = ~n5811 & ~n5828;
  assign n5830 = ~i_StoB_REQ0 & ~n5829;
  assign n5831 = ~i_StoB_REQ0 & ~n5830;
  assign n5832 = ~i_StoB_REQ14 & ~n5831;
  assign n5833 = ~i_StoB_REQ14 & ~n5832;
  assign n5834 = controllable_BtoS_ACK14 & ~n5833;
  assign n5835 = ~i_StoB_REQ13 & ~n5608;
  assign n5836 = ~n5611 & ~n5835;
  assign n5837 = n4466 & ~n5836;
  assign n5838 = ~i_StoB_REQ12 & ~n5818;
  assign n5839 = ~i_StoB_REQ12 & ~n5838;
  assign n5840 = controllable_BtoS_ACK12 & ~n5839;
  assign n5841 = ~i_StoB_REQ12 & ~n5602;
  assign n5842 = ~n5819 & ~n5841;
  assign n5843 = ~controllable_BtoS_ACK12 & ~n5842;
  assign n5844 = ~n5840 & ~n5843;
  assign n5845 = ~controllable_BtoS_ACK13 & ~n5844;
  assign n5846 = ~n5003 & ~n5845;
  assign n5847 = ~i_StoB_REQ13 & ~n5846;
  assign n5848 = ~n5204 & ~n5847;
  assign n5849 = ~n4466 & ~n5848;
  assign n5850 = ~n5837 & ~n5849;
  assign n5851 = ~i_StoB_REQ0 & ~n5850;
  assign n5852 = ~i_StoB_REQ0 & ~n5851;
  assign n5853 = i_StoB_REQ14 & ~n5852;
  assign n5854 = ~n5832 & ~n5853;
  assign n5855 = ~controllable_BtoS_ACK14 & ~n5854;
  assign n5856 = ~n5834 & ~n5855;
  assign n5857 = controllable_ENQ & ~n5856;
  assign n5858 = controllable_ENQ & ~n5857;
  assign n5859 = i_RtoB_ACK1 & ~n5858;
  assign n5860 = i_StoB_REQ14 & ~n4991;
  assign n5861 = i_StoB_REQ0 & ~n4989;
  assign n5862 = controllable_BtoS_ACK13 & ~n4952;
  assign n5863 = controllable_BtoS_ACK2 & n4693;
  assign n5864 = n4477 & n5863;
  assign n5865 = i_StoB_REQ2 & controllable_BtoS_ACK2;
  assign n5866 = ~n5419 & ~n5865;
  assign n5867 = ~n4477 & ~n5866;
  assign n5868 = ~n5864 & ~n5867;
  assign n5869 = n4476 & ~n5868;
  assign n5870 = ~n4702 & ~n5425;
  assign n5871 = controllable_BtoS_ACK2 & ~n5870;
  assign n5872 = ~n5428 & ~n5871;
  assign n5873 = n4477 & ~n5872;
  assign n5874 = controllable_BtoS_ACK2 & n4702;
  assign n5875 = ~n5432 & ~n5874;
  assign n5876 = ~n4477 & ~n5875;
  assign n5877 = ~n5873 & ~n5876;
  assign n5878 = ~n4476 & ~n5877;
  assign n5879 = ~n5869 & ~n5878;
  assign n5880 = ~i_StoB_REQ3 & ~n5879;
  assign n5881 = ~n4715 & ~n5880;
  assign n5882 = controllable_BtoS_ACK3 & ~n5881;
  assign n5883 = ~controllable_BtoS_ACK3 & ~n5879;
  assign n5884 = ~n5882 & ~n5883;
  assign n5885 = n4475 & ~n5884;
  assign n5886 = ~i_StoB_REQ3 & n5863;
  assign n5887 = ~n4723 & ~n5886;
  assign n5888 = controllable_BtoS_ACK3 & ~n5887;
  assign n5889 = ~n4482 & ~n5865;
  assign n5890 = ~n4477 & ~n5889;
  assign n5891 = ~n4484 & ~n5890;
  assign n5892 = n4476 & ~n5891;
  assign n5893 = ~n4479 & ~n4702;
  assign n5894 = controllable_BtoS_ACK2 & ~n5893;
  assign n5895 = ~n4482 & ~n5894;
  assign n5896 = n4477 & ~n5895;
  assign n5897 = ~n4482 & ~n5874;
  assign n5898 = ~n4477 & ~n5897;
  assign n5899 = ~n5896 & ~n5898;
  assign n5900 = ~n4476 & ~n5899;
  assign n5901 = ~n5892 & ~n5900;
  assign n5902 = i_StoB_REQ3 & ~n5901;
  assign n5903 = ~n4477 & ~n5867;
  assign n5904 = n4476 & ~n5903;
  assign n5905 = ~n5878 & ~n5904;
  assign n5906 = ~i_StoB_REQ3 & ~n5905;
  assign n5907 = ~n5902 & ~n5906;
  assign n5908 = ~controllable_BtoS_ACK3 & ~n5907;
  assign n5909 = ~n5888 & ~n5908;
  assign n5910 = ~n4475 & ~n5909;
  assign n5911 = ~n5885 & ~n5910;
  assign n5912 = ~i_StoB_REQ4 & ~n5911;
  assign n5913 = ~n4736 & ~n5912;
  assign n5914 = controllable_BtoS_ACK4 & ~n5913;
  assign n5915 = ~controllable_BtoS_ACK4 & ~n5911;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = n4474 & ~n5916;
  assign n5918 = ~n4741 & ~n5886;
  assign n5919 = controllable_BtoS_ACK3 & ~n5918;
  assign n5920 = ~controllable_BtoS_ACK3 & n5863;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = ~i_StoB_REQ4 & ~n5921;
  assign n5923 = ~n4748 & ~n5922;
  assign n5924 = controllable_BtoS_ACK4 & ~n5923;
  assign n5925 = ~i_StoB_REQ3 & ~n5901;
  assign n5926 = ~n4723 & ~n5925;
  assign n5927 = controllable_BtoS_ACK3 & ~n5926;
  assign n5928 = ~controllable_BtoS_ACK3 & ~n5901;
  assign n5929 = ~n5927 & ~n5928;
  assign n5930 = n4475 & ~n5929;
  assign n5931 = ~n5888 & ~n5928;
  assign n5932 = ~n4475 & ~n5931;
  assign n5933 = ~n5930 & ~n5932;
  assign n5934 = i_StoB_REQ4 & ~n5933;
  assign n5935 = ~n4723 & ~n5906;
  assign n5936 = controllable_BtoS_ACK3 & ~n5935;
  assign n5937 = ~controllable_BtoS_ACK3 & ~n5905;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = n4475 & ~n5938;
  assign n5940 = ~n5910 & ~n5939;
  assign n5941 = ~i_StoB_REQ4 & ~n5940;
  assign n5942 = ~n5934 & ~n5941;
  assign n5943 = ~controllable_BtoS_ACK4 & ~n5942;
  assign n5944 = ~n5924 & ~n5943;
  assign n5945 = ~n4474 & ~n5944;
  assign n5946 = ~n5917 & ~n5945;
  assign n5947 = ~i_StoB_REQ5 & ~n5946;
  assign n5948 = ~n4763 & ~n5947;
  assign n5949 = controllable_BtoS_ACK5 & ~n5948;
  assign n5950 = ~controllable_BtoS_ACK5 & ~n5946;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = n4473 & ~n5951;
  assign n5953 = ~n4768 & ~n5922;
  assign n5954 = controllable_BtoS_ACK4 & ~n5953;
  assign n5955 = ~controllable_BtoS_ACK4 & ~n5921;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~i_StoB_REQ5 & ~n5956;
  assign n5958 = ~n4775 & ~n5957;
  assign n5959 = controllable_BtoS_ACK5 & ~n5958;
  assign n5960 = ~i_StoB_REQ4 & ~n5933;
  assign n5961 = ~n4748 & ~n5960;
  assign n5962 = controllable_BtoS_ACK4 & ~n5961;
  assign n5963 = ~controllable_BtoS_ACK4 & ~n5933;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = n4474 & ~n5964;
  assign n5966 = ~n5924 & ~n5963;
  assign n5967 = ~n4474 & ~n5966;
  assign n5968 = ~n5965 & ~n5967;
  assign n5969 = i_StoB_REQ5 & ~n5968;
  assign n5970 = ~n4748 & ~n5941;
  assign n5971 = controllable_BtoS_ACK4 & ~n5970;
  assign n5972 = ~controllable_BtoS_ACK4 & ~n5940;
  assign n5973 = ~n5971 & ~n5972;
  assign n5974 = n4474 & ~n5973;
  assign n5975 = ~n5945 & ~n5974;
  assign n5976 = ~i_StoB_REQ5 & ~n5975;
  assign n5977 = ~n5969 & ~n5976;
  assign n5978 = ~controllable_BtoS_ACK5 & ~n5977;
  assign n5979 = ~n5959 & ~n5978;
  assign n5980 = ~n4473 & ~n5979;
  assign n5981 = ~n5952 & ~n5980;
  assign n5982 = ~i_StoB_REQ8 & ~n5981;
  assign n5983 = ~n4790 & ~n5982;
  assign n5984 = controllable_BtoS_ACK8 & ~n5983;
  assign n5985 = ~controllable_BtoS_ACK8 & ~n5981;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = n4472 & ~n5986;
  assign n5988 = ~n4795 & ~n5957;
  assign n5989 = controllable_BtoS_ACK5 & ~n5988;
  assign n5990 = ~controllable_BtoS_ACK5 & ~n5956;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = ~i_StoB_REQ8 & ~n5991;
  assign n5993 = ~n4802 & ~n5992;
  assign n5994 = controllable_BtoS_ACK8 & ~n5993;
  assign n5995 = ~i_StoB_REQ5 & ~n5968;
  assign n5996 = ~n4775 & ~n5995;
  assign n5997 = controllable_BtoS_ACK5 & ~n5996;
  assign n5998 = ~controllable_BtoS_ACK5 & ~n5968;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = n4473 & ~n5999;
  assign n6001 = ~n5959 & ~n5998;
  assign n6002 = ~n4473 & ~n6001;
  assign n6003 = ~n6000 & ~n6002;
  assign n6004 = i_StoB_REQ8 & ~n6003;
  assign n6005 = ~n4775 & ~n5976;
  assign n6006 = controllable_BtoS_ACK5 & ~n6005;
  assign n6007 = ~controllable_BtoS_ACK5 & ~n5975;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = n4473 & ~n6008;
  assign n6010 = ~n5980 & ~n6009;
  assign n6011 = ~i_StoB_REQ8 & ~n6010;
  assign n6012 = ~n6004 & ~n6011;
  assign n6013 = ~controllable_BtoS_ACK8 & ~n6012;
  assign n6014 = ~n5994 & ~n6013;
  assign n6015 = ~n4472 & ~n6014;
  assign n6016 = ~n5987 & ~n6015;
  assign n6017 = n4471 & ~n6016;
  assign n6018 = ~n4815 & ~n5992;
  assign n6019 = controllable_BtoS_ACK8 & ~n6018;
  assign n6020 = ~controllable_BtoS_ACK8 & ~n5991;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n4471 & ~n6021;
  assign n6023 = ~n6017 & ~n6022;
  assign n6024 = ~i_StoB_REQ6 & ~n6023;
  assign n6025 = ~n4824 & ~n6024;
  assign n6026 = controllable_BtoS_ACK6 & ~n6025;
  assign n6027 = ~i_StoB_REQ8 & ~n6003;
  assign n6028 = ~n4802 & ~n6027;
  assign n6029 = controllable_BtoS_ACK8 & ~n6028;
  assign n6030 = ~controllable_BtoS_ACK8 & ~n6003;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = n4472 & ~n6031;
  assign n6033 = ~n5994 & ~n6030;
  assign n6034 = ~n4472 & ~n6033;
  assign n6035 = ~n6032 & ~n6034;
  assign n6036 = ~n4471 & ~n6035;
  assign n6037 = ~n6017 & ~n6036;
  assign n6038 = i_StoB_REQ6 & ~n6037;
  assign n6039 = ~n4802 & ~n6011;
  assign n6040 = controllable_BtoS_ACK8 & ~n6039;
  assign n6041 = ~controllable_BtoS_ACK8 & ~n6010;
  assign n6042 = ~n6040 & ~n6041;
  assign n6043 = n4472 & ~n6042;
  assign n6044 = ~n6015 & ~n6043;
  assign n6045 = ~n4471 & ~n6044;
  assign n6046 = ~n6017 & ~n6045;
  assign n6047 = ~i_StoB_REQ6 & ~n6046;
  assign n6048 = ~n6038 & ~n6047;
  assign n6049 = ~controllable_BtoS_ACK6 & ~n6048;
  assign n6050 = ~n6026 & ~n6049;
  assign n6051 = ~i_StoB_REQ7 & ~n6050;
  assign n6052 = ~n4839 & ~n6051;
  assign n6053 = controllable_BtoS_ACK7 & ~n6052;
  assign n6054 = ~controllable_BtoS_ACK7 & ~n6050;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = n4470 & ~n6055;
  assign n6057 = ~i_StoB_REQ6 & ~n6021;
  assign n6058 = ~n4847 & ~n6057;
  assign n6059 = controllable_BtoS_ACK6 & ~n6058;
  assign n6060 = ~controllable_BtoS_ACK6 & ~n6021;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~i_StoB_REQ7 & ~n6061;
  assign n6063 = ~n4854 & ~n6062;
  assign n6064 = controllable_BtoS_ACK7 & ~n6063;
  assign n6065 = n4471 & ~n6035;
  assign n6066 = ~n6022 & ~n6065;
  assign n6067 = ~i_StoB_REQ6 & ~n6066;
  assign n6068 = ~n4860 & ~n6067;
  assign n6069 = controllable_BtoS_ACK6 & ~n6068;
  assign n6070 = ~controllable_BtoS_ACK6 & ~n6035;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = i_StoB_REQ7 & ~n6071;
  assign n6073 = n4471 & ~n6044;
  assign n6074 = ~n6022 & ~n6073;
  assign n6075 = ~i_StoB_REQ6 & ~n6074;
  assign n6076 = ~n4860 & ~n6075;
  assign n6077 = controllable_BtoS_ACK6 & ~n6076;
  assign n6078 = ~n6036 & ~n6073;
  assign n6079 = i_StoB_REQ6 & ~n6078;
  assign n6080 = ~i_StoB_REQ6 & ~n6044;
  assign n6081 = ~n6079 & ~n6080;
  assign n6082 = ~controllable_BtoS_ACK6 & ~n6081;
  assign n6083 = ~n6077 & ~n6082;
  assign n6084 = ~i_StoB_REQ7 & ~n6083;
  assign n6085 = ~n6072 & ~n6084;
  assign n6086 = ~controllable_BtoS_ACK7 & ~n6085;
  assign n6087 = ~n6064 & ~n6086;
  assign n6088 = ~n4470 & ~n6087;
  assign n6089 = ~n6056 & ~n6088;
  assign n6090 = n4469 & ~n6089;
  assign n6091 = ~n4872 & ~n6062;
  assign n6092 = controllable_BtoS_ACK7 & ~n6091;
  assign n6093 = ~controllable_BtoS_ACK7 & ~n6061;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = ~n4469 & ~n6094;
  assign n6096 = ~n6090 & ~n6095;
  assign n6097 = ~i_StoB_REQ9 & ~n6096;
  assign n6098 = ~n4881 & ~n6097;
  assign n6099 = controllable_BtoS_ACK9 & ~n6098;
  assign n6100 = ~i_StoB_REQ7 & ~n6071;
  assign n6101 = ~n4854 & ~n6100;
  assign n6102 = controllable_BtoS_ACK7 & ~n6101;
  assign n6103 = ~controllable_BtoS_ACK7 & ~n6071;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = n4470 & ~n6104;
  assign n6106 = ~n6064 & ~n6103;
  assign n6107 = ~n4470 & ~n6106;
  assign n6108 = ~n6105 & ~n6107;
  assign n6109 = ~n4469 & ~n6108;
  assign n6110 = ~n6090 & ~n6109;
  assign n6111 = i_StoB_REQ9 & ~n6110;
  assign n6112 = ~n4854 & ~n6084;
  assign n6113 = controllable_BtoS_ACK7 & ~n6112;
  assign n6114 = ~controllable_BtoS_ACK7 & ~n6083;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = n4470 & ~n6115;
  assign n6117 = ~n6088 & ~n6116;
  assign n6118 = ~n4469 & ~n6117;
  assign n6119 = ~n6090 & ~n6118;
  assign n6120 = ~i_StoB_REQ9 & ~n6119;
  assign n6121 = ~n6111 & ~n6120;
  assign n6122 = ~controllable_BtoS_ACK9 & ~n6121;
  assign n6123 = ~n6099 & ~n6122;
  assign n6124 = n4468 & ~n6123;
  assign n6125 = ~i_StoB_REQ9 & ~n6094;
  assign n6126 = ~n4897 & ~n6125;
  assign n6127 = controllable_BtoS_ACK9 & ~n6126;
  assign n6128 = ~controllable_BtoS_ACK9 & ~n6094;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = ~n4468 & ~n6129;
  assign n6131 = ~n6124 & ~n6130;
  assign n6132 = ~i_StoB_REQ11 & ~n6131;
  assign n6133 = ~n4906 & ~n6132;
  assign n6134 = controllable_BtoS_ACK11 & ~n6133;
  assign n6135 = n4469 & ~n6108;
  assign n6136 = ~n6095 & ~n6135;
  assign n6137 = ~i_StoB_REQ9 & ~n6136;
  assign n6138 = ~n4912 & ~n6137;
  assign n6139 = controllable_BtoS_ACK9 & ~n6138;
  assign n6140 = ~controllable_BtoS_ACK9 & ~n6108;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = ~n4468 & ~n6141;
  assign n6143 = ~n6124 & ~n6142;
  assign n6144 = i_StoB_REQ11 & ~n6143;
  assign n6145 = n4469 & ~n6117;
  assign n6146 = ~n6095 & ~n6145;
  assign n6147 = ~i_StoB_REQ9 & ~n6146;
  assign n6148 = ~n4912 & ~n6147;
  assign n6149 = controllable_BtoS_ACK9 & ~n6148;
  assign n6150 = ~n6109 & ~n6145;
  assign n6151 = i_StoB_REQ9 & ~n6150;
  assign n6152 = ~i_StoB_REQ9 & ~n6117;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = ~controllable_BtoS_ACK9 & ~n6153;
  assign n6155 = ~n6149 & ~n6154;
  assign n6156 = ~n4468 & ~n6155;
  assign n6157 = ~n6124 & ~n6156;
  assign n6158 = ~i_StoB_REQ11 & ~n6157;
  assign n6159 = ~n6144 & ~n6158;
  assign n6160 = ~controllable_BtoS_ACK11 & ~n6159;
  assign n6161 = ~n6134 & ~n6160;
  assign n6162 = n4467 & ~n6161;
  assign n6163 = ~i_StoB_REQ11 & ~n6129;
  assign n6164 = ~n4927 & ~n6163;
  assign n6165 = controllable_BtoS_ACK11 & ~n6164;
  assign n6166 = ~controllable_BtoS_ACK11 & ~n6129;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = ~n4467 & ~n6167;
  assign n6169 = ~n6162 & ~n6168;
  assign n6170 = ~i_StoB_REQ12 & ~n6169;
  assign n6171 = ~n4936 & ~n6170;
  assign n6172 = controllable_BtoS_ACK12 & ~n6171;
  assign n6173 = n4468 & ~n6141;
  assign n6174 = ~n6130 & ~n6173;
  assign n6175 = ~i_StoB_REQ11 & ~n6174;
  assign n6176 = ~n4942 & ~n6175;
  assign n6177 = controllable_BtoS_ACK11 & ~n6176;
  assign n6178 = ~controllable_BtoS_ACK11 & ~n6141;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = ~n4467 & ~n6179;
  assign n6181 = ~n6162 & ~n6180;
  assign n6182 = i_StoB_REQ12 & ~n6181;
  assign n6183 = n4468 & ~n6155;
  assign n6184 = ~n6130 & ~n6183;
  assign n6185 = ~i_StoB_REQ11 & ~n6184;
  assign n6186 = ~n4942 & ~n6185;
  assign n6187 = controllable_BtoS_ACK11 & ~n6186;
  assign n6188 = ~n6142 & ~n6183;
  assign n6189 = i_StoB_REQ11 & ~n6188;
  assign n6190 = ~i_StoB_REQ11 & ~n6155;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = ~controllable_BtoS_ACK11 & ~n6191;
  assign n6193 = ~n6187 & ~n6192;
  assign n6194 = ~n4467 & ~n6193;
  assign n6195 = ~n6162 & ~n6194;
  assign n6196 = ~i_StoB_REQ12 & ~n6195;
  assign n6197 = ~n6182 & ~n6196;
  assign n6198 = ~controllable_BtoS_ACK12 & ~n6197;
  assign n6199 = ~n6172 & ~n6198;
  assign n6200 = ~controllable_BtoS_ACK13 & ~n6199;
  assign n6201 = ~n5862 & ~n6200;
  assign n6202 = i_StoB_REQ13 & ~n6201;
  assign n6203 = i_StoB_REQ12 & ~n4948;
  assign n6204 = i_StoB_REQ11 & ~n4918;
  assign n6205 = i_StoB_REQ9 & ~n4888;
  assign n6206 = i_StoB_REQ7 & ~n4835;
  assign n6207 = i_StoB_REQ6 & ~n4831;
  assign n6208 = i_StoB_REQ8 & ~n4786;
  assign n6209 = i_StoB_REQ5 & ~n4759;
  assign n6210 = i_StoB_REQ4 & ~n4732;
  assign n6211 = i_StoB_REQ3 & ~n4711;
  assign n6212 = controllable_BtoS_ACK2 & ~n4689;
  assign n6213 = ~i_StoB_REQ2 & n4689;
  assign n6214 = ~i_StoB_REQ2 & ~n6213;
  assign n6215 = ~controllable_BtoS_ACK2 & n6214;
  assign n6216 = ~n6212 & ~n6215;
  assign n6217 = n4477 & ~n6216;
  assign n6218 = ~n5613 & ~n6217;
  assign n6219 = n4476 & ~n6218;
  assign n6220 = ~n5623 & ~n6219;
  assign n6221 = ~i_StoB_REQ3 & ~n6220;
  assign n6222 = ~n6211 & ~n6221;
  assign n6223 = controllable_BtoS_ACK3 & ~n6222;
  assign n6224 = i_StoB_REQ3 & ~n5879;
  assign n6225 = ~n6221 & ~n6224;
  assign n6226 = ~controllable_BtoS_ACK3 & ~n6225;
  assign n6227 = ~n6223 & ~n6226;
  assign n6228 = n4475 & ~n6227;
  assign n6229 = i_StoB_REQ3 & ~n4726;
  assign n6230 = ~i_StoB_REQ3 & ~n6216;
  assign n6231 = ~n6229 & ~n6230;
  assign n6232 = controllable_BtoS_ACK3 & ~n6231;
  assign n6233 = ~n5636 & ~n5902;
  assign n6234 = ~controllable_BtoS_ACK3 & ~n6233;
  assign n6235 = ~n6232 & ~n6234;
  assign n6236 = ~n4475 & ~n6235;
  assign n6237 = ~n6228 & ~n6236;
  assign n6238 = ~i_StoB_REQ4 & ~n6237;
  assign n6239 = ~n6210 & ~n6238;
  assign n6240 = controllable_BtoS_ACK4 & ~n6239;
  assign n6241 = i_StoB_REQ4 & ~n5911;
  assign n6242 = ~n6238 & ~n6241;
  assign n6243 = ~controllable_BtoS_ACK4 & ~n6242;
  assign n6244 = ~n6240 & ~n6243;
  assign n6245 = n4474 & ~n6244;
  assign n6246 = i_StoB_REQ4 & ~n4753;
  assign n6247 = i_StoB_REQ3 & ~n4696;
  assign n6248 = ~n6230 & ~n6247;
  assign n6249 = controllable_BtoS_ACK3 & ~n6248;
  assign n6250 = i_StoB_REQ3 & n5863;
  assign n6251 = ~n6230 & ~n6250;
  assign n6252 = ~controllable_BtoS_ACK3 & ~n6251;
  assign n6253 = ~n6249 & ~n6252;
  assign n6254 = ~i_StoB_REQ4 & ~n6253;
  assign n6255 = ~n6246 & ~n6254;
  assign n6256 = controllable_BtoS_ACK4 & ~n6255;
  assign n6257 = ~n5636 & ~n6229;
  assign n6258 = controllable_BtoS_ACK3 & ~n6257;
  assign n6259 = i_StoB_REQ3 & ~n5905;
  assign n6260 = ~n5636 & ~n6259;
  assign n6261 = ~controllable_BtoS_ACK3 & ~n6260;
  assign n6262 = ~n6258 & ~n6261;
  assign n6263 = n4475 & ~n6262;
  assign n6264 = ~n6236 & ~n6263;
  assign n6265 = ~i_StoB_REQ4 & ~n6264;
  assign n6266 = ~n5934 & ~n6265;
  assign n6267 = ~controllable_BtoS_ACK4 & ~n6266;
  assign n6268 = ~n6256 & ~n6267;
  assign n6269 = ~n4474 & ~n6268;
  assign n6270 = ~n6245 & ~n6269;
  assign n6271 = ~i_StoB_REQ5 & ~n6270;
  assign n6272 = ~n6209 & ~n6271;
  assign n6273 = controllable_BtoS_ACK5 & ~n6272;
  assign n6274 = i_StoB_REQ5 & ~n5946;
  assign n6275 = ~n6271 & ~n6274;
  assign n6276 = ~controllable_BtoS_ACK5 & ~n6275;
  assign n6277 = ~n6273 & ~n6276;
  assign n6278 = n4473 & ~n6277;
  assign n6279 = i_StoB_REQ5 & ~n4780;
  assign n6280 = i_StoB_REQ4 & ~n4744;
  assign n6281 = ~n6254 & ~n6280;
  assign n6282 = controllable_BtoS_ACK4 & ~n6281;
  assign n6283 = i_StoB_REQ4 & ~n5921;
  assign n6284 = ~n6254 & ~n6283;
  assign n6285 = ~controllable_BtoS_ACK4 & ~n6284;
  assign n6286 = ~n6282 & ~n6285;
  assign n6287 = ~i_StoB_REQ5 & ~n6286;
  assign n6288 = ~n6279 & ~n6287;
  assign n6289 = controllable_BtoS_ACK5 & ~n6288;
  assign n6290 = ~n6246 & ~n6265;
  assign n6291 = controllable_BtoS_ACK4 & ~n6290;
  assign n6292 = i_StoB_REQ4 & ~n5940;
  assign n6293 = ~n6265 & ~n6292;
  assign n6294 = ~controllable_BtoS_ACK4 & ~n6293;
  assign n6295 = ~n6291 & ~n6294;
  assign n6296 = n4474 & ~n6295;
  assign n6297 = ~n6269 & ~n6296;
  assign n6298 = ~i_StoB_REQ5 & ~n6297;
  assign n6299 = ~n5969 & ~n6298;
  assign n6300 = ~controllable_BtoS_ACK5 & ~n6299;
  assign n6301 = ~n6289 & ~n6300;
  assign n6302 = ~n4473 & ~n6301;
  assign n6303 = ~n6278 & ~n6302;
  assign n6304 = ~i_StoB_REQ8 & ~n6303;
  assign n6305 = ~n6208 & ~n6304;
  assign n6306 = controllable_BtoS_ACK8 & ~n6305;
  assign n6307 = i_StoB_REQ8 & ~n5981;
  assign n6308 = ~n6304 & ~n6307;
  assign n6309 = ~controllable_BtoS_ACK8 & ~n6308;
  assign n6310 = ~n6306 & ~n6309;
  assign n6311 = n4472 & ~n6310;
  assign n6312 = i_StoB_REQ8 & ~n4807;
  assign n6313 = i_StoB_REQ5 & ~n4771;
  assign n6314 = ~n6287 & ~n6313;
  assign n6315 = controllable_BtoS_ACK5 & ~n6314;
  assign n6316 = i_StoB_REQ5 & ~n5956;
  assign n6317 = ~n6287 & ~n6316;
  assign n6318 = ~controllable_BtoS_ACK5 & ~n6317;
  assign n6319 = ~n6315 & ~n6318;
  assign n6320 = ~i_StoB_REQ8 & ~n6319;
  assign n6321 = ~n6312 & ~n6320;
  assign n6322 = controllable_BtoS_ACK8 & ~n6321;
  assign n6323 = ~n6279 & ~n6298;
  assign n6324 = controllable_BtoS_ACK5 & ~n6323;
  assign n6325 = i_StoB_REQ5 & ~n5975;
  assign n6326 = ~n6298 & ~n6325;
  assign n6327 = ~controllable_BtoS_ACK5 & ~n6326;
  assign n6328 = ~n6324 & ~n6327;
  assign n6329 = n4473 & ~n6328;
  assign n6330 = ~n6302 & ~n6329;
  assign n6331 = ~i_StoB_REQ8 & ~n6330;
  assign n6332 = ~n6004 & ~n6331;
  assign n6333 = ~controllable_BtoS_ACK8 & ~n6332;
  assign n6334 = ~n6322 & ~n6333;
  assign n6335 = ~n4472 & ~n6334;
  assign n6336 = ~n6311 & ~n6335;
  assign n6337 = n4471 & ~n6336;
  assign n6338 = i_StoB_REQ8 & ~n4798;
  assign n6339 = ~n6320 & ~n6338;
  assign n6340 = controllable_BtoS_ACK8 & ~n6339;
  assign n6341 = i_StoB_REQ8 & ~n5991;
  assign n6342 = ~n6320 & ~n6341;
  assign n6343 = ~controllable_BtoS_ACK8 & ~n6342;
  assign n6344 = ~n6340 & ~n6343;
  assign n6345 = ~n4471 & ~n6344;
  assign n6346 = ~n6337 & ~n6345;
  assign n6347 = ~i_StoB_REQ6 & ~n6346;
  assign n6348 = ~n6207 & ~n6347;
  assign n6349 = controllable_BtoS_ACK6 & ~n6348;
  assign n6350 = ~n6312 & ~n6331;
  assign n6351 = controllable_BtoS_ACK8 & ~n6350;
  assign n6352 = i_StoB_REQ8 & ~n6010;
  assign n6353 = ~n6331 & ~n6352;
  assign n6354 = ~controllable_BtoS_ACK8 & ~n6353;
  assign n6355 = ~n6351 & ~n6354;
  assign n6356 = n4472 & ~n6355;
  assign n6357 = ~n6335 & ~n6356;
  assign n6358 = ~n4471 & ~n6357;
  assign n6359 = ~n6337 & ~n6358;
  assign n6360 = ~i_StoB_REQ6 & ~n6359;
  assign n6361 = ~n6038 & ~n6360;
  assign n6362 = ~controllable_BtoS_ACK6 & ~n6361;
  assign n6363 = ~n6349 & ~n6362;
  assign n6364 = ~i_StoB_REQ7 & ~n6363;
  assign n6365 = ~n6206 & ~n6364;
  assign n6366 = controllable_BtoS_ACK7 & ~n6365;
  assign n6367 = i_StoB_REQ7 & ~n6050;
  assign n6368 = ~n6364 & ~n6367;
  assign n6369 = ~controllable_BtoS_ACK7 & ~n6368;
  assign n6370 = ~n6366 & ~n6369;
  assign n6371 = n4470 & ~n6370;
  assign n6372 = i_StoB_REQ7 & ~n4864;
  assign n6373 = i_StoB_REQ6 & ~n4818;
  assign n6374 = ~i_StoB_REQ6 & ~n6344;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = controllable_BtoS_ACK6 & ~n6375;
  assign n6377 = i_StoB_REQ6 & ~n6021;
  assign n6378 = ~n6374 & ~n6377;
  assign n6379 = ~controllable_BtoS_ACK6 & ~n6378;
  assign n6380 = ~n6376 & ~n6379;
  assign n6381 = ~i_StoB_REQ7 & ~n6380;
  assign n6382 = ~n6372 & ~n6381;
  assign n6383 = controllable_BtoS_ACK7 & ~n6382;
  assign n6384 = i_StoB_REQ6 & ~n4829;
  assign n6385 = n4471 & ~n6357;
  assign n6386 = ~n6345 & ~n6385;
  assign n6387 = ~i_StoB_REQ6 & ~n6386;
  assign n6388 = ~n6384 & ~n6387;
  assign n6389 = controllable_BtoS_ACK6 & ~n6388;
  assign n6390 = ~i_StoB_REQ6 & ~n6357;
  assign n6391 = ~n6079 & ~n6390;
  assign n6392 = ~controllable_BtoS_ACK6 & ~n6391;
  assign n6393 = ~n6389 & ~n6392;
  assign n6394 = ~i_StoB_REQ7 & ~n6393;
  assign n6395 = ~n6072 & ~n6394;
  assign n6396 = ~controllable_BtoS_ACK7 & ~n6395;
  assign n6397 = ~n6383 & ~n6396;
  assign n6398 = ~n4470 & ~n6397;
  assign n6399 = ~n6371 & ~n6398;
  assign n6400 = n4469 & ~n6399;
  assign n6401 = i_StoB_REQ7 & ~n4850;
  assign n6402 = ~n6381 & ~n6401;
  assign n6403 = controllable_BtoS_ACK7 & ~n6402;
  assign n6404 = i_StoB_REQ7 & ~n6061;
  assign n6405 = ~n6381 & ~n6404;
  assign n6406 = ~controllable_BtoS_ACK7 & ~n6405;
  assign n6407 = ~n6403 & ~n6406;
  assign n6408 = ~n4469 & ~n6407;
  assign n6409 = ~n6400 & ~n6408;
  assign n6410 = ~i_StoB_REQ9 & ~n6409;
  assign n6411 = ~n6205 & ~n6410;
  assign n6412 = controllable_BtoS_ACK9 & ~n6411;
  assign n6413 = ~n6372 & ~n6394;
  assign n6414 = controllable_BtoS_ACK7 & ~n6413;
  assign n6415 = i_StoB_REQ7 & ~n6083;
  assign n6416 = ~n6394 & ~n6415;
  assign n6417 = ~controllable_BtoS_ACK7 & ~n6416;
  assign n6418 = ~n6414 & ~n6417;
  assign n6419 = n4470 & ~n6418;
  assign n6420 = ~n6398 & ~n6419;
  assign n6421 = ~n4469 & ~n6420;
  assign n6422 = ~n6400 & ~n6421;
  assign n6423 = ~i_StoB_REQ9 & ~n6422;
  assign n6424 = ~n6111 & ~n6423;
  assign n6425 = ~controllable_BtoS_ACK9 & ~n6424;
  assign n6426 = ~n6412 & ~n6425;
  assign n6427 = n4468 & ~n6426;
  assign n6428 = i_StoB_REQ9 & ~n4875;
  assign n6429 = ~i_StoB_REQ9 & ~n6407;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = controllable_BtoS_ACK9 & ~n6430;
  assign n6432 = i_StoB_REQ9 & ~n6094;
  assign n6433 = ~n6429 & ~n6432;
  assign n6434 = ~controllable_BtoS_ACK9 & ~n6433;
  assign n6435 = ~n6431 & ~n6434;
  assign n6436 = ~n4468 & ~n6435;
  assign n6437 = ~n6427 & ~n6436;
  assign n6438 = ~i_StoB_REQ11 & ~n6437;
  assign n6439 = ~n6204 & ~n6438;
  assign n6440 = controllable_BtoS_ACK11 & ~n6439;
  assign n6441 = i_StoB_REQ9 & ~n4886;
  assign n6442 = n4469 & ~n6420;
  assign n6443 = ~n6408 & ~n6442;
  assign n6444 = ~i_StoB_REQ9 & ~n6443;
  assign n6445 = ~n6441 & ~n6444;
  assign n6446 = controllable_BtoS_ACK9 & ~n6445;
  assign n6447 = ~i_StoB_REQ9 & ~n6420;
  assign n6448 = ~n6151 & ~n6447;
  assign n6449 = ~controllable_BtoS_ACK9 & ~n6448;
  assign n6450 = ~n6446 & ~n6449;
  assign n6451 = ~n4468 & ~n6450;
  assign n6452 = ~n6427 & ~n6451;
  assign n6453 = ~i_StoB_REQ11 & ~n6452;
  assign n6454 = ~n6144 & ~n6453;
  assign n6455 = ~controllable_BtoS_ACK11 & ~n6454;
  assign n6456 = ~n6440 & ~n6455;
  assign n6457 = n4467 & ~n6456;
  assign n6458 = i_StoB_REQ11 & ~n4900;
  assign n6459 = ~i_StoB_REQ11 & ~n6435;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = controllable_BtoS_ACK11 & ~n6460;
  assign n6462 = i_StoB_REQ11 & ~n6129;
  assign n6463 = ~n6459 & ~n6462;
  assign n6464 = ~controllable_BtoS_ACK11 & ~n6463;
  assign n6465 = ~n6461 & ~n6464;
  assign n6466 = ~n4467 & ~n6465;
  assign n6467 = ~n6457 & ~n6466;
  assign n6468 = ~i_StoB_REQ12 & ~n6467;
  assign n6469 = ~n6203 & ~n6468;
  assign n6470 = controllable_BtoS_ACK12 & ~n6469;
  assign n6471 = i_StoB_REQ11 & ~n4916;
  assign n6472 = n4468 & ~n6450;
  assign n6473 = ~n6436 & ~n6472;
  assign n6474 = ~i_StoB_REQ11 & ~n6473;
  assign n6475 = ~n6471 & ~n6474;
  assign n6476 = controllable_BtoS_ACK11 & ~n6475;
  assign n6477 = ~i_StoB_REQ11 & ~n6450;
  assign n6478 = ~n6189 & ~n6477;
  assign n6479 = ~controllable_BtoS_ACK11 & ~n6478;
  assign n6480 = ~n6476 & ~n6479;
  assign n6481 = ~n4467 & ~n6480;
  assign n6482 = ~n6457 & ~n6481;
  assign n6483 = ~i_StoB_REQ12 & ~n6482;
  assign n6484 = ~n6182 & ~n6483;
  assign n6485 = ~controllable_BtoS_ACK12 & ~n6484;
  assign n6486 = ~n6470 & ~n6485;
  assign n6487 = ~i_StoB_REQ13 & ~n6486;
  assign n6488 = ~n6202 & ~n6487;
  assign n6489 = n4466 & ~n6488;
  assign n6490 = controllable_BtoS_ACK13 & ~n4983;
  assign n6491 = n4467 & ~n6179;
  assign n6492 = ~n6168 & ~n6491;
  assign n6493 = ~i_StoB_REQ12 & ~n6492;
  assign n6494 = ~n4979 & ~n6493;
  assign n6495 = controllable_BtoS_ACK12 & ~n6494;
  assign n6496 = ~controllable_BtoS_ACK12 & ~n6179;
  assign n6497 = ~n6495 & ~n6496;
  assign n6498 = ~controllable_BtoS_ACK13 & ~n6497;
  assign n6499 = ~n6490 & ~n6498;
  assign n6500 = i_StoB_REQ13 & ~n6499;
  assign n6501 = i_StoB_REQ12 & ~n4930;
  assign n6502 = ~i_StoB_REQ12 & ~n6465;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = controllable_BtoS_ACK12 & ~n6503;
  assign n6505 = i_StoB_REQ12 & ~n6167;
  assign n6506 = ~n6502 & ~n6505;
  assign n6507 = ~controllable_BtoS_ACK12 & ~n6506;
  assign n6508 = ~n6504 & ~n6507;
  assign n6509 = controllable_BtoS_ACK13 & ~n6508;
  assign n6510 = i_StoB_REQ12 & ~n4946;
  assign n6511 = n4467 & ~n6480;
  assign n6512 = ~n6466 & ~n6511;
  assign n6513 = ~i_StoB_REQ12 & ~n6512;
  assign n6514 = ~n6510 & ~n6513;
  assign n6515 = controllable_BtoS_ACK12 & ~n6514;
  assign n6516 = n4467 & ~n6193;
  assign n6517 = ~n6180 & ~n6516;
  assign n6518 = i_StoB_REQ12 & ~n6517;
  assign n6519 = ~i_StoB_REQ12 & ~n6480;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = ~controllable_BtoS_ACK12 & ~n6520;
  assign n6522 = ~n6515 & ~n6521;
  assign n6523 = ~controllable_BtoS_ACK13 & ~n6522;
  assign n6524 = ~n6509 & ~n6523;
  assign n6525 = ~i_StoB_REQ13 & ~n6524;
  assign n6526 = ~n6500 & ~n6525;
  assign n6527 = ~n4466 & ~n6526;
  assign n6528 = ~n6489 & ~n6527;
  assign n6529 = ~i_StoB_REQ0 & ~n6528;
  assign n6530 = ~n5861 & ~n6529;
  assign n6531 = ~i_StoB_REQ14 & ~n6530;
  assign n6532 = ~n5860 & ~n6531;
  assign n6533 = controllable_BtoS_ACK14 & ~n6532;
  assign n6534 = controllable_BtoS_ACK13 & ~n4685;
  assign n6535 = ~n6200 & ~n6534;
  assign n6536 = i_StoB_REQ13 & ~n6535;
  assign n6537 = ~i_StoB_REQ13 & ~n6199;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = n4466 & ~n6538;
  assign n6540 = controllable_BtoS_ACK13 & ~n4962;
  assign n6541 = ~n6498 & ~n6540;
  assign n6542 = i_StoB_REQ13 & ~n6541;
  assign n6543 = ~i_StoB_REQ12 & ~n6167;
  assign n6544 = ~n4969 & ~n6543;
  assign n6545 = controllable_BtoS_ACK12 & ~n6544;
  assign n6546 = ~controllable_BtoS_ACK12 & ~n6167;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = controllable_BtoS_ACK13 & ~n6547;
  assign n6549 = ~n6168 & ~n6516;
  assign n6550 = ~i_StoB_REQ12 & ~n6549;
  assign n6551 = ~n4979 & ~n6550;
  assign n6552 = controllable_BtoS_ACK12 & ~n6551;
  assign n6553 = ~i_StoB_REQ12 & ~n6193;
  assign n6554 = ~n6518 & ~n6553;
  assign n6555 = ~controllable_BtoS_ACK12 & ~n6554;
  assign n6556 = ~n6552 & ~n6555;
  assign n6557 = ~controllable_BtoS_ACK13 & ~n6556;
  assign n6558 = ~n6548 & ~n6557;
  assign n6559 = ~i_StoB_REQ13 & ~n6558;
  assign n6560 = ~n6542 & ~n6559;
  assign n6561 = ~n4466 & ~n6560;
  assign n6562 = ~n6539 & ~n6561;
  assign n6563 = ~i_StoB_REQ0 & ~n6562;
  assign n6564 = ~n5103 & ~n6563;
  assign n6565 = i_StoB_REQ14 & ~n6564;
  assign n6566 = ~n6531 & ~n6565;
  assign n6567 = ~controllable_BtoS_ACK14 & ~n6566;
  assign n6568 = ~n6533 & ~n6567;
  assign n6569 = controllable_ENQ & ~n6568;
  assign n6570 = controllable_ENQ & ~n6569;
  assign n6571 = ~i_RtoB_ACK1 & ~n6570;
  assign n6572 = ~n5859 & ~n6571;
  assign n6573 = controllable_BtoR_REQ1 & ~n6572;
  assign n6574 = ~i_StoB_REQ14 & ~n6564;
  assign n6575 = ~n5011 & ~n6574;
  assign n6576 = controllable_BtoS_ACK14 & ~n6575;
  assign n6577 = ~controllable_BtoS_ACK14 & ~n6564;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = controllable_ENQ & ~n6578;
  assign n6580 = controllable_ENQ & ~n6579;
  assign n6581 = ~controllable_BtoR_REQ1 & ~n6580;
  assign n6582 = ~n6573 & ~n6581;
  assign n6583 = ~controllable_BtoR_REQ0 & ~n6582;
  assign n6584 = ~controllable_BtoR_REQ0 & ~n6583;
  assign n6585 = i_RtoB_ACK0 & ~n6584;
  assign n6586 = controllable_BtoS_ACK2 & ~n5865;
  assign n6587 = ~n4477 & ~n6586;
  assign n6588 = ~n5864 & ~n6587;
  assign n6589 = n4476 & ~n6588;
  assign n6590 = n4477 & ~n4490;
  assign n6591 = ~n4494 & ~n5874;
  assign n6592 = ~n4477 & ~n6591;
  assign n6593 = ~n6590 & ~n6592;
  assign n6594 = ~n4476 & ~n6593;
  assign n6595 = ~n6589 & ~n6594;
  assign n6596 = ~i_StoB_REQ3 & ~n6595;
  assign n6597 = ~n4715 & ~n6596;
  assign n6598 = controllable_BtoS_ACK3 & ~n6597;
  assign n6599 = ~controllable_BtoS_ACK3 & ~n6595;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = n4475 & ~n6600;
  assign n6602 = ~n4477 & ~n6587;
  assign n6603 = n4476 & ~n6602;
  assign n6604 = ~n6594 & ~n6603;
  assign n6605 = ~controllable_BtoS_ACK3 & ~n6604;
  assign n6606 = ~n5888 & ~n6605;
  assign n6607 = ~n4475 & ~n6606;
  assign n6608 = ~n6601 & ~n6607;
  assign n6609 = ~i_StoB_REQ4 & ~n6608;
  assign n6610 = ~n4736 & ~n6609;
  assign n6611 = controllable_BtoS_ACK4 & ~n6610;
  assign n6612 = ~controllable_BtoS_ACK4 & ~n6608;
  assign n6613 = ~n6611 & ~n6612;
  assign n6614 = n4474 & ~n6613;
  assign n6615 = ~i_StoB_REQ3 & ~n6604;
  assign n6616 = ~n4723 & ~n6615;
  assign n6617 = controllable_BtoS_ACK3 & ~n6616;
  assign n6618 = ~n6605 & ~n6617;
  assign n6619 = n4475 & ~n6618;
  assign n6620 = ~n6607 & ~n6619;
  assign n6621 = ~controllable_BtoS_ACK4 & ~n6620;
  assign n6622 = ~n5924 & ~n6621;
  assign n6623 = ~n4474 & ~n6622;
  assign n6624 = ~n6614 & ~n6623;
  assign n6625 = ~i_StoB_REQ5 & ~n6624;
  assign n6626 = ~n4763 & ~n6625;
  assign n6627 = controllable_BtoS_ACK5 & ~n6626;
  assign n6628 = ~controllable_BtoS_ACK5 & ~n6624;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = n4473 & ~n6629;
  assign n6631 = ~i_StoB_REQ4 & ~n6620;
  assign n6632 = ~n4748 & ~n6631;
  assign n6633 = controllable_BtoS_ACK4 & ~n6632;
  assign n6634 = ~n6621 & ~n6633;
  assign n6635 = n4474 & ~n6634;
  assign n6636 = ~n6623 & ~n6635;
  assign n6637 = ~controllable_BtoS_ACK5 & ~n6636;
  assign n6638 = ~n5959 & ~n6637;
  assign n6639 = ~n4473 & ~n6638;
  assign n6640 = ~n6630 & ~n6639;
  assign n6641 = ~i_StoB_REQ8 & ~n6640;
  assign n6642 = ~n4790 & ~n6641;
  assign n6643 = controllable_BtoS_ACK8 & ~n6642;
  assign n6644 = ~controllable_BtoS_ACK8 & ~n6640;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = n4472 & ~n6645;
  assign n6647 = ~i_StoB_REQ5 & ~n6636;
  assign n6648 = ~n4775 & ~n6647;
  assign n6649 = controllable_BtoS_ACK5 & ~n6648;
  assign n6650 = ~n6637 & ~n6649;
  assign n6651 = n4473 & ~n6650;
  assign n6652 = ~n6639 & ~n6651;
  assign n6653 = ~controllable_BtoS_ACK8 & ~n6652;
  assign n6654 = ~n5994 & ~n6653;
  assign n6655 = ~n4472 & ~n6654;
  assign n6656 = ~n6646 & ~n6655;
  assign n6657 = n4471 & ~n6656;
  assign n6658 = ~n6022 & ~n6657;
  assign n6659 = ~i_StoB_REQ6 & ~n6658;
  assign n6660 = ~n4824 & ~n6659;
  assign n6661 = controllable_BtoS_ACK6 & ~n6660;
  assign n6662 = ~i_StoB_REQ8 & ~n6652;
  assign n6663 = ~n4802 & ~n6662;
  assign n6664 = controllable_BtoS_ACK8 & ~n6663;
  assign n6665 = ~n6653 & ~n6664;
  assign n6666 = n4472 & ~n6665;
  assign n6667 = ~n6655 & ~n6666;
  assign n6668 = ~n4471 & ~n6667;
  assign n6669 = ~n6657 & ~n6668;
  assign n6670 = ~controllable_BtoS_ACK6 & ~n6669;
  assign n6671 = ~n6661 & ~n6670;
  assign n6672 = ~i_StoB_REQ7 & ~n6671;
  assign n6673 = ~n4839 & ~n6672;
  assign n6674 = controllable_BtoS_ACK7 & ~n6673;
  assign n6675 = ~controllable_BtoS_ACK7 & ~n6671;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = n4470 & ~n6676;
  assign n6678 = n4471 & ~n6667;
  assign n6679 = ~n6022 & ~n6678;
  assign n6680 = ~i_StoB_REQ6 & ~n6679;
  assign n6681 = ~n4860 & ~n6680;
  assign n6682 = controllable_BtoS_ACK6 & ~n6681;
  assign n6683 = ~controllable_BtoS_ACK6 & ~n6667;
  assign n6684 = ~n6682 & ~n6683;
  assign n6685 = ~controllable_BtoS_ACK7 & ~n6684;
  assign n6686 = ~n6064 & ~n6685;
  assign n6687 = ~n4470 & ~n6686;
  assign n6688 = ~n6677 & ~n6687;
  assign n6689 = n4469 & ~n6688;
  assign n6690 = ~n6095 & ~n6689;
  assign n6691 = ~i_StoB_REQ9 & ~n6690;
  assign n6692 = ~n4881 & ~n6691;
  assign n6693 = controllable_BtoS_ACK9 & ~n6692;
  assign n6694 = ~i_StoB_REQ7 & ~n6684;
  assign n6695 = ~n4854 & ~n6694;
  assign n6696 = controllable_BtoS_ACK7 & ~n6695;
  assign n6697 = ~n6685 & ~n6696;
  assign n6698 = n4470 & ~n6697;
  assign n6699 = ~n6687 & ~n6698;
  assign n6700 = ~n4469 & ~n6699;
  assign n6701 = ~n6689 & ~n6700;
  assign n6702 = ~controllable_BtoS_ACK9 & ~n6701;
  assign n6703 = ~n6693 & ~n6702;
  assign n6704 = n4468 & ~n6703;
  assign n6705 = ~n6130 & ~n6704;
  assign n6706 = ~i_StoB_REQ11 & ~n6705;
  assign n6707 = ~n4906 & ~n6706;
  assign n6708 = controllable_BtoS_ACK11 & ~n6707;
  assign n6709 = n4469 & ~n6699;
  assign n6710 = ~n6095 & ~n6709;
  assign n6711 = ~i_StoB_REQ9 & ~n6710;
  assign n6712 = ~n4912 & ~n6711;
  assign n6713 = controllable_BtoS_ACK9 & ~n6712;
  assign n6714 = ~controllable_BtoS_ACK9 & ~n6699;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = ~n4468 & ~n6715;
  assign n6717 = ~n6704 & ~n6716;
  assign n6718 = ~controllable_BtoS_ACK11 & ~n6717;
  assign n6719 = ~n6708 & ~n6718;
  assign n6720 = n4467 & ~n6719;
  assign n6721 = ~n6168 & ~n6720;
  assign n6722 = ~i_StoB_REQ12 & ~n6721;
  assign n6723 = ~n4936 & ~n6722;
  assign n6724 = controllable_BtoS_ACK12 & ~n6723;
  assign n6725 = n4468 & ~n6715;
  assign n6726 = ~n6130 & ~n6725;
  assign n6727 = ~i_StoB_REQ11 & ~n6726;
  assign n6728 = ~n4942 & ~n6727;
  assign n6729 = controllable_BtoS_ACK11 & ~n6728;
  assign n6730 = ~controllable_BtoS_ACK11 & ~n6715;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = ~n4467 & ~n6731;
  assign n6733 = ~n6720 & ~n6732;
  assign n6734 = ~controllable_BtoS_ACK12 & ~n6733;
  assign n6735 = ~n6724 & ~n6734;
  assign n6736 = ~controllable_BtoS_ACK13 & ~n6735;
  assign n6737 = ~n6534 & ~n6736;
  assign n6738 = i_StoB_REQ13 & ~n6737;
  assign n6739 = ~i_StoB_REQ13 & ~n6735;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = n4466 & ~n6740;
  assign n6742 = n4467 & ~n6731;
  assign n6743 = ~n6168 & ~n6742;
  assign n6744 = ~i_StoB_REQ12 & ~n6743;
  assign n6745 = ~n4979 & ~n6744;
  assign n6746 = controllable_BtoS_ACK12 & ~n6745;
  assign n6747 = ~controllable_BtoS_ACK12 & ~n6731;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = ~controllable_BtoS_ACK13 & ~n6748;
  assign n6750 = ~n6540 & ~n6749;
  assign n6751 = i_StoB_REQ13 & ~n6750;
  assign n6752 = ~n6548 & ~n6749;
  assign n6753 = ~i_StoB_REQ13 & ~n6752;
  assign n6754 = ~n6751 & ~n6753;
  assign n6755 = ~n4466 & ~n6754;
  assign n6756 = ~n6741 & ~n6755;
  assign n6757 = ~i_StoB_REQ0 & ~n6756;
  assign n6758 = ~n5103 & ~n6757;
  assign n6759 = ~i_StoB_REQ14 & ~n6758;
  assign n6760 = ~n5011 & ~n6759;
  assign n6761 = controllable_BtoS_ACK14 & ~n6760;
  assign n6762 = ~controllable_BtoS_ACK14 & ~n6758;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = controllable_ENQ & ~n6763;
  assign n6765 = ~controllable_ENQ & ~n5856;
  assign n6766 = ~n6764 & ~n6765;
  assign n6767 = i_RtoB_ACK1 & ~n6766;
  assign n6768 = ~controllable_ENQ & ~n6568;
  assign n6769 = ~n6764 & ~n6768;
  assign n6770 = ~i_RtoB_ACK1 & ~n6769;
  assign n6771 = ~n6767 & ~n6770;
  assign n6772 = controllable_BtoR_REQ1 & ~n6771;
  assign n6773 = i_RtoB_ACK1 & ~n6580;
  assign n6774 = ~controllable_ENQ & ~n6578;
  assign n6775 = ~n6764 & ~n6774;
  assign n6776 = ~i_RtoB_ACK1 & ~n6775;
  assign n6777 = ~n6773 & ~n6776;
  assign n6778 = ~controllable_BtoR_REQ1 & ~n6777;
  assign n6779 = ~n6772 & ~n6778;
  assign n6780 = ~controllable_BtoR_REQ0 & ~n6779;
  assign n6781 = ~controllable_BtoR_REQ0 & ~n6780;
  assign n6782 = ~i_RtoB_ACK0 & ~n6781;
  assign n6783 = ~n6585 & ~n6782;
  assign n6784 = controllable_DEQ & ~n6783;
  assign n6785 = i_RtoB_ACK1 & ~n5856;
  assign n6786 = ~i_RtoB_ACK1 & ~n6568;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = controllable_BtoR_REQ1 & ~n6787;
  assign n6789 = ~controllable_BtoR_REQ1 & ~n6578;
  assign n6790 = ~n6788 & ~n6789;
  assign n6791 = ~controllable_BtoR_REQ0 & ~n6790;
  assign n6792 = ~controllable_BtoR_REQ0 & ~n6791;
  assign n6793 = i_RtoB_ACK0 & ~n6792;
  assign n6794 = controllable_BtoR_REQ1 & ~n6763;
  assign n6795 = i_RtoB_ACK1 & ~n6578;
  assign n6796 = ~i_RtoB_ACK1 & ~n6763;
  assign n6797 = ~n6795 & ~n6796;
  assign n6798 = ~controllable_BtoR_REQ1 & ~n6797;
  assign n6799 = ~n6794 & ~n6798;
  assign n6800 = ~controllable_BtoR_REQ0 & ~n6799;
  assign n6801 = ~controllable_BtoR_REQ0 & ~n6800;
  assign n6802 = ~i_RtoB_ACK0 & ~n6801;
  assign n6803 = ~n6793 & ~n6802;
  assign n6804 = ~controllable_DEQ & ~n6803;
  assign n6805 = ~n6784 & ~n6804;
  assign n6806 = i_FULL & ~n6805;
  assign n6807 = ~n6579 & ~n6765;
  assign n6808 = i_RtoB_ACK1 & ~n6807;
  assign n6809 = ~n6579 & ~n6768;
  assign n6810 = ~i_RtoB_ACK1 & ~n6809;
  assign n6811 = ~n6808 & ~n6810;
  assign n6812 = controllable_BtoR_REQ1 & ~n6811;
  assign n6813 = ~i_RtoB_ACK1 & ~n6578;
  assign n6814 = ~n6773 & ~n6813;
  assign n6815 = ~controllable_BtoR_REQ1 & ~n6814;
  assign n6816 = ~n6812 & ~n6815;
  assign n6817 = ~controllable_BtoR_REQ0 & ~n6816;
  assign n6818 = ~controllable_BtoR_REQ0 & ~n6817;
  assign n6819 = ~i_RtoB_ACK0 & ~n6818;
  assign n6820 = ~n6585 & ~n6819;
  assign n6821 = controllable_DEQ & ~n6820;
  assign n6822 = controllable_BtoR_REQ1 & ~n6775;
  assign n6823 = ~n6776 & ~n6795;
  assign n6824 = ~controllable_BtoR_REQ1 & ~n6823;
  assign n6825 = ~n6822 & ~n6824;
  assign n6826 = ~controllable_BtoR_REQ0 & ~n6825;
  assign n6827 = ~controllable_BtoR_REQ0 & ~n6826;
  assign n6828 = ~i_RtoB_ACK0 & ~n6827;
  assign n6829 = ~n6793 & ~n6828;
  assign n6830 = ~controllable_DEQ & ~n6829;
  assign n6831 = ~n6821 & ~n6830;
  assign n6832 = ~i_FULL & ~n6831;
  assign n6833 = ~n6806 & ~n6832;
  assign n6834 = i_nEMPTY & ~n6833;
  assign n6835 = ~controllable_ENQ & ~n6765;
  assign n6836 = i_RtoB_ACK1 & ~n6835;
  assign n6837 = ~controllable_ENQ & ~n6768;
  assign n6838 = ~i_RtoB_ACK1 & ~n6837;
  assign n6839 = ~n6836 & ~n6838;
  assign n6840 = controllable_BtoR_REQ1 & ~n6839;
  assign n6841 = ~controllable_ENQ & ~n6774;
  assign n6842 = ~i_RtoB_ACK1 & ~n6841;
  assign n6843 = ~i_RtoB_ACK1 & ~n6842;
  assign n6844 = ~controllable_BtoR_REQ1 & ~n6843;
  assign n6845 = ~n6840 & ~n6844;
  assign n6846 = ~controllable_BtoR_REQ0 & ~n6845;
  assign n6847 = ~controllable_BtoR_REQ0 & ~n6846;
  assign n6848 = ~i_RtoB_ACK0 & ~n6847;
  assign n6849 = ~i_RtoB_ACK0 & ~n6848;
  assign n6850 = controllable_DEQ & ~n6849;
  assign n6851 = controllable_ENQ & ~n6764;
  assign n6852 = controllable_BtoR_REQ1 & ~n6851;
  assign n6853 = ~i_RtoB_ACK1 & ~n6851;
  assign n6854 = ~n6773 & ~n6853;
  assign n6855 = ~controllable_BtoR_REQ1 & ~n6854;
  assign n6856 = ~n6852 & ~n6855;
  assign n6857 = ~controllable_BtoR_REQ0 & ~n6856;
  assign n6858 = ~controllable_BtoR_REQ0 & ~n6857;
  assign n6859 = ~i_RtoB_ACK0 & ~n6858;
  assign n6860 = ~n6585 & ~n6859;
  assign n6861 = ~controllable_DEQ & ~n6860;
  assign n6862 = ~n6850 & ~n6861;
  assign n6863 = i_FULL & ~n6862;
  assign n6864 = ~i_RtoB_ACK1 & ~n6813;
  assign n6865 = ~controllable_BtoR_REQ1 & ~n6864;
  assign n6866 = ~n6788 & ~n6865;
  assign n6867 = ~controllable_BtoR_REQ0 & ~n6866;
  assign n6868 = ~controllable_BtoR_REQ0 & ~n6867;
  assign n6869 = ~i_RtoB_ACK0 & ~n6868;
  assign n6870 = ~i_RtoB_ACK0 & ~n6869;
  assign n6871 = controllable_DEQ & ~n6870;
  assign n6872 = ~n6770 & ~n6773;
  assign n6873 = ~controllable_BtoR_REQ1 & ~n6872;
  assign n6874 = ~n6772 & ~n6873;
  assign n6875 = ~controllable_BtoR_REQ0 & ~n6874;
  assign n6876 = ~controllable_BtoR_REQ0 & ~n6875;
  assign n6877 = ~i_RtoB_ACK0 & ~n6876;
  assign n6878 = ~n6585 & ~n6877;
  assign n6879 = ~controllable_DEQ & ~n6878;
  assign n6880 = ~n6871 & ~n6879;
  assign n6881 = ~i_FULL & ~n6880;
  assign n6882 = ~n6863 & ~n6881;
  assign n6883 = ~i_nEMPTY & ~n6882;
  assign n6884 = ~n6834 & ~n6883;
  assign n6885 = controllable_BtoS_ACK0 & ~n6884;
  assign n6886 = i_StoB_REQ0 & ~n5850;
  assign n6887 = ~n5830 & ~n6886;
  assign n6888 = ~i_StoB_REQ14 & ~n6887;
  assign n6889 = ~i_StoB_REQ14 & ~n6888;
  assign n6890 = controllable_BtoS_ACK14 & ~n6889;
  assign n6891 = i_StoB_REQ14 & ~n5850;
  assign n6892 = ~n6888 & ~n6891;
  assign n6893 = ~controllable_BtoS_ACK14 & ~n6892;
  assign n6894 = ~n6890 & ~n6893;
  assign n6895 = controllable_ENQ & ~n6894;
  assign n6896 = controllable_ENQ & ~n6895;
  assign n6897 = i_RtoB_ACK1 & ~n6896;
  assign n6898 = i_StoB_REQ14 & ~n5104;
  assign n6899 = i_StoB_REQ0 & ~n6562;
  assign n6900 = ~n6529 & ~n6899;
  assign n6901 = ~i_StoB_REQ14 & ~n6900;
  assign n6902 = ~n6898 & ~n6901;
  assign n6903 = controllable_BtoS_ACK14 & ~n6902;
  assign n6904 = i_StoB_REQ14 & ~n6562;
  assign n6905 = ~n6901 & ~n6904;
  assign n6906 = ~controllable_BtoS_ACK14 & ~n6905;
  assign n6907 = ~n6903 & ~n6906;
  assign n6908 = controllable_ENQ & ~n6907;
  assign n6909 = controllable_ENQ & ~n6908;
  assign n6910 = ~i_RtoB_ACK1 & ~n6909;
  assign n6911 = ~n6897 & ~n6910;
  assign n6912 = controllable_BtoR_REQ1 & ~n6911;
  assign n6913 = ~i_StoB_REQ14 & ~n6562;
  assign n6914 = ~n5108 & ~n6913;
  assign n6915 = controllable_BtoS_ACK14 & ~n6914;
  assign n6916 = ~controllable_BtoS_ACK14 & ~n6562;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = controllable_ENQ & ~n6917;
  assign n6919 = controllable_ENQ & ~n6918;
  assign n6920 = ~controllable_BtoR_REQ1 & ~n6919;
  assign n6921 = ~n6912 & ~n6920;
  assign n6922 = ~controllable_BtoR_REQ0 & ~n6921;
  assign n6923 = ~controllable_BtoR_REQ0 & ~n6922;
  assign n6924 = i_RtoB_ACK0 & ~n6923;
  assign n6925 = ~i_StoB_REQ14 & ~n6756;
  assign n6926 = ~n5108 & ~n6925;
  assign n6927 = controllable_BtoS_ACK14 & ~n6926;
  assign n6928 = ~controllable_BtoS_ACK14 & ~n6756;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = controllable_ENQ & ~n6929;
  assign n6931 = ~controllable_ENQ & ~n6894;
  assign n6932 = ~n6930 & ~n6931;
  assign n6933 = i_RtoB_ACK1 & ~n6932;
  assign n6934 = ~controllable_ENQ & ~n6907;
  assign n6935 = ~n6930 & ~n6934;
  assign n6936 = ~i_RtoB_ACK1 & ~n6935;
  assign n6937 = ~n6933 & ~n6936;
  assign n6938 = controllable_BtoR_REQ1 & ~n6937;
  assign n6939 = i_RtoB_ACK1 & ~n6919;
  assign n6940 = ~controllable_ENQ & ~n6917;
  assign n6941 = ~n6930 & ~n6940;
  assign n6942 = ~i_RtoB_ACK1 & ~n6941;
  assign n6943 = ~n6939 & ~n6942;
  assign n6944 = ~controllable_BtoR_REQ1 & ~n6943;
  assign n6945 = ~n6938 & ~n6944;
  assign n6946 = ~controllable_BtoR_REQ0 & ~n6945;
  assign n6947 = ~controllable_BtoR_REQ0 & ~n6946;
  assign n6948 = ~i_RtoB_ACK0 & ~n6947;
  assign n6949 = ~n6924 & ~n6948;
  assign n6950 = controllable_DEQ & ~n6949;
  assign n6951 = i_RtoB_ACK1 & ~n6894;
  assign n6952 = ~i_RtoB_ACK1 & ~n6907;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = controllable_BtoR_REQ1 & ~n6953;
  assign n6955 = ~controllable_BtoR_REQ1 & ~n6917;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~controllable_BtoR_REQ0 & ~n6956;
  assign n6958 = ~controllable_BtoR_REQ0 & ~n6957;
  assign n6959 = i_RtoB_ACK0 & ~n6958;
  assign n6960 = controllable_BtoR_REQ1 & ~n6929;
  assign n6961 = i_RtoB_ACK1 & ~n6917;
  assign n6962 = ~i_RtoB_ACK1 & ~n6929;
  assign n6963 = ~n6961 & ~n6962;
  assign n6964 = ~controllable_BtoR_REQ1 & ~n6963;
  assign n6965 = ~n6960 & ~n6964;
  assign n6966 = ~controllable_BtoR_REQ0 & ~n6965;
  assign n6967 = ~controllable_BtoR_REQ0 & ~n6966;
  assign n6968 = ~i_RtoB_ACK0 & ~n6967;
  assign n6969 = ~n6959 & ~n6968;
  assign n6970 = ~controllable_DEQ & ~n6969;
  assign n6971 = ~n6950 & ~n6970;
  assign n6972 = i_FULL & ~n6971;
  assign n6973 = ~n6918 & ~n6931;
  assign n6974 = i_RtoB_ACK1 & ~n6973;
  assign n6975 = ~n6918 & ~n6934;
  assign n6976 = ~i_RtoB_ACK1 & ~n6975;
  assign n6977 = ~n6974 & ~n6976;
  assign n6978 = controllable_BtoR_REQ1 & ~n6977;
  assign n6979 = ~i_RtoB_ACK1 & ~n6917;
  assign n6980 = ~n6939 & ~n6979;
  assign n6981 = ~controllable_BtoR_REQ1 & ~n6980;
  assign n6982 = ~n6978 & ~n6981;
  assign n6983 = ~controllable_BtoR_REQ0 & ~n6982;
  assign n6984 = ~controllable_BtoR_REQ0 & ~n6983;
  assign n6985 = ~i_RtoB_ACK0 & ~n6984;
  assign n6986 = ~n6924 & ~n6985;
  assign n6987 = controllable_DEQ & ~n6986;
  assign n6988 = controllable_BtoR_REQ1 & ~n6941;
  assign n6989 = ~n6942 & ~n6961;
  assign n6990 = ~controllable_BtoR_REQ1 & ~n6989;
  assign n6991 = ~n6988 & ~n6990;
  assign n6992 = ~controllable_BtoR_REQ0 & ~n6991;
  assign n6993 = ~controllable_BtoR_REQ0 & ~n6992;
  assign n6994 = ~i_RtoB_ACK0 & ~n6993;
  assign n6995 = ~n6959 & ~n6994;
  assign n6996 = ~controllable_DEQ & ~n6995;
  assign n6997 = ~n6987 & ~n6996;
  assign n6998 = ~i_FULL & ~n6997;
  assign n6999 = ~n6972 & ~n6998;
  assign n7000 = i_nEMPTY & ~n6999;
  assign n7001 = ~controllable_ENQ & ~n6931;
  assign n7002 = i_RtoB_ACK1 & ~n7001;
  assign n7003 = ~controllable_ENQ & ~n6934;
  assign n7004 = ~i_RtoB_ACK1 & ~n7003;
  assign n7005 = ~n7002 & ~n7004;
  assign n7006 = controllable_BtoR_REQ1 & ~n7005;
  assign n7007 = ~controllable_ENQ & ~n6940;
  assign n7008 = ~i_RtoB_ACK1 & ~n7007;
  assign n7009 = ~i_RtoB_ACK1 & ~n7008;
  assign n7010 = ~controllable_BtoR_REQ1 & ~n7009;
  assign n7011 = ~n7006 & ~n7010;
  assign n7012 = ~controllable_BtoR_REQ0 & ~n7011;
  assign n7013 = ~controllable_BtoR_REQ0 & ~n7012;
  assign n7014 = ~i_RtoB_ACK0 & ~n7013;
  assign n7015 = ~i_RtoB_ACK0 & ~n7014;
  assign n7016 = controllable_DEQ & ~n7015;
  assign n7017 = controllable_ENQ & ~n6930;
  assign n7018 = controllable_BtoR_REQ1 & ~n7017;
  assign n7019 = ~i_RtoB_ACK1 & ~n7017;
  assign n7020 = ~n6939 & ~n7019;
  assign n7021 = ~controllable_BtoR_REQ1 & ~n7020;
  assign n7022 = ~n7018 & ~n7021;
  assign n7023 = ~controllable_BtoR_REQ0 & ~n7022;
  assign n7024 = ~controllable_BtoR_REQ0 & ~n7023;
  assign n7025 = ~i_RtoB_ACK0 & ~n7024;
  assign n7026 = ~n6924 & ~n7025;
  assign n7027 = ~controllable_DEQ & ~n7026;
  assign n7028 = ~n7016 & ~n7027;
  assign n7029 = i_FULL & ~n7028;
  assign n7030 = ~i_RtoB_ACK1 & ~n6979;
  assign n7031 = ~controllable_BtoR_REQ1 & ~n7030;
  assign n7032 = ~n6954 & ~n7031;
  assign n7033 = ~controllable_BtoR_REQ0 & ~n7032;
  assign n7034 = ~controllable_BtoR_REQ0 & ~n7033;
  assign n7035 = ~i_RtoB_ACK0 & ~n7034;
  assign n7036 = ~i_RtoB_ACK0 & ~n7035;
  assign n7037 = controllable_DEQ & ~n7036;
  assign n7038 = ~n6936 & ~n6939;
  assign n7039 = ~controllable_BtoR_REQ1 & ~n7038;
  assign n7040 = ~n6938 & ~n7039;
  assign n7041 = ~controllable_BtoR_REQ0 & ~n7040;
  assign n7042 = ~controllable_BtoR_REQ0 & ~n7041;
  assign n7043 = ~i_RtoB_ACK0 & ~n7042;
  assign n7044 = ~n6924 & ~n7043;
  assign n7045 = ~controllable_DEQ & ~n7044;
  assign n7046 = ~n7037 & ~n7045;
  assign n7047 = ~i_FULL & ~n7046;
  assign n7048 = ~n7029 & ~n7047;
  assign n7049 = ~i_nEMPTY & ~n7048;
  assign n7050 = ~n7000 & ~n7049;
  assign n7051 = ~controllable_BtoS_ACK0 & ~n7050;
  assign n7052 = ~n6885 & ~n7051;
  assign n7053 = n4465 & ~n7052;
  assign n7054 = i_RtoB_ACK1 & ~n5221;
  assign n7055 = i_StoB_REQ14 & ~n5208;
  assign n7056 = i_StoB_REQ0 & ~n5316;
  assign n7057 = ~controllable_BtoS_ACK13 & ~n6547;
  assign n7058 = ~n4973 & ~n7057;
  assign n7059 = i_StoB_REQ13 & ~n7058;
  assign n7060 = ~i_StoB_REQ13 & ~n6508;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = ~i_StoB_REQ0 & ~n7061;
  assign n7063 = ~n7056 & ~n7062;
  assign n7064 = ~i_StoB_REQ14 & ~n7063;
  assign n7065 = ~n7055 & ~n7064;
  assign n7066 = controllable_BtoS_ACK14 & ~n7065;
  assign n7067 = ~n5003 & ~n7057;
  assign n7068 = i_StoB_REQ13 & ~n7067;
  assign n7069 = ~i_StoB_REQ13 & ~n6547;
  assign n7070 = ~n7068 & ~n7069;
  assign n7071 = ~i_StoB_REQ0 & ~n7070;
  assign n7072 = ~n5312 & ~n7071;
  assign n7073 = i_StoB_REQ14 & ~n7072;
  assign n7074 = ~n7064 & ~n7073;
  assign n7075 = ~controllable_BtoS_ACK14 & ~n7074;
  assign n7076 = ~n7066 & ~n7075;
  assign n7077 = controllable_ENQ & ~n7076;
  assign n7078 = controllable_ENQ & ~n7077;
  assign n7079 = ~i_RtoB_ACK1 & ~n7078;
  assign n7080 = ~n7054 & ~n7079;
  assign n7081 = controllable_BtoR_REQ1 & ~n7080;
  assign n7082 = ~i_StoB_REQ14 & ~n7072;
  assign n7083 = ~n5216 & ~n7082;
  assign n7084 = controllable_BtoS_ACK14 & ~n7083;
  assign n7085 = ~controllable_BtoS_ACK14 & ~n7072;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = controllable_ENQ & ~n7086;
  assign n7088 = controllable_ENQ & ~n7087;
  assign n7089 = ~controllable_BtoR_REQ1 & ~n7088;
  assign n7090 = ~n7081 & ~n7089;
  assign n7091 = ~controllable_BtoR_REQ0 & ~n7090;
  assign n7092 = ~controllable_BtoR_REQ0 & ~n7091;
  assign n7093 = i_RtoB_ACK0 & ~n7092;
  assign n7094 = ~n5238 & ~n7087;
  assign n7095 = i_RtoB_ACK1 & ~n7094;
  assign n7096 = ~controllable_ENQ & ~n7076;
  assign n7097 = ~n7087 & ~n7096;
  assign n7098 = ~i_RtoB_ACK1 & ~n7097;
  assign n7099 = ~n7095 & ~n7098;
  assign n7100 = controllable_BtoR_REQ1 & ~n7099;
  assign n7101 = i_RtoB_ACK1 & ~n7088;
  assign n7102 = ~i_RtoB_ACK1 & ~n7086;
  assign n7103 = ~n7101 & ~n7102;
  assign n7104 = ~controllable_BtoR_REQ1 & ~n7103;
  assign n7105 = ~n7100 & ~n7104;
  assign n7106 = ~controllable_BtoR_REQ0 & ~n7105;
  assign n7107 = ~controllable_BtoR_REQ0 & ~n7106;
  assign n7108 = ~i_RtoB_ACK0 & ~n7107;
  assign n7109 = ~n7093 & ~n7108;
  assign n7110 = controllable_DEQ & ~n7109;
  assign n7111 = i_RtoB_ACK1 & ~n5219;
  assign n7112 = ~i_RtoB_ACK1 & ~n7076;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = controllable_BtoR_REQ1 & ~n7113;
  assign n7115 = ~controllable_BtoR_REQ1 & ~n7086;
  assign n7116 = ~n7114 & ~n7115;
  assign n7117 = ~controllable_BtoR_REQ0 & ~n7116;
  assign n7118 = ~controllable_BtoR_REQ0 & ~n7117;
  assign n7119 = i_RtoB_ACK0 & ~n7118;
  assign n7120 = ~controllable_BtoR_REQ0 & ~n7086;
  assign n7121 = ~controllable_BtoR_REQ0 & ~n7120;
  assign n7122 = ~i_RtoB_ACK0 & ~n7121;
  assign n7123 = ~n7119 & ~n7122;
  assign n7124 = ~controllable_DEQ & ~n7123;
  assign n7125 = ~n7110 & ~n7124;
  assign n7126 = i_nEMPTY & ~n7125;
  assign n7127 = i_RtoB_ACK1 & ~n5267;
  assign n7128 = ~controllable_ENQ & ~n7096;
  assign n7129 = ~i_RtoB_ACK1 & ~n7128;
  assign n7130 = ~n7127 & ~n7129;
  assign n7131 = controllable_BtoR_REQ1 & ~n7130;
  assign n7132 = ~controllable_ENQ & ~n7086;
  assign n7133 = ~controllable_ENQ & ~n7132;
  assign n7134 = ~i_RtoB_ACK1 & ~n7133;
  assign n7135 = ~i_RtoB_ACK1 & ~n7134;
  assign n7136 = ~controllable_BtoR_REQ1 & ~n7135;
  assign n7137 = ~n7131 & ~n7136;
  assign n7138 = ~controllable_BtoR_REQ0 & ~n7137;
  assign n7139 = ~controllable_BtoR_REQ0 & ~n7138;
  assign n7140 = ~i_RtoB_ACK0 & ~n7139;
  assign n7141 = ~i_RtoB_ACK0 & ~n7140;
  assign n7142 = controllable_DEQ & ~n7141;
  assign n7143 = ~controllable_BtoR_REQ0 & ~n7088;
  assign n7144 = ~controllable_BtoR_REQ0 & ~n7143;
  assign n7145 = ~i_RtoB_ACK0 & ~n7144;
  assign n7146 = ~n7093 & ~n7145;
  assign n7147 = ~controllable_DEQ & ~n7146;
  assign n7148 = ~n7142 & ~n7147;
  assign n7149 = i_FULL & ~n7148;
  assign n7150 = ~i_RtoB_ACK1 & ~n7102;
  assign n7151 = ~controllable_BtoR_REQ1 & ~n7150;
  assign n7152 = ~n7114 & ~n7151;
  assign n7153 = ~controllable_BtoR_REQ0 & ~n7152;
  assign n7154 = ~controllable_BtoR_REQ0 & ~n7153;
  assign n7155 = ~i_RtoB_ACK0 & ~n7154;
  assign n7156 = ~i_RtoB_ACK0 & ~n7155;
  assign n7157 = controllable_DEQ & ~n7156;
  assign n7158 = ~n7098 & ~n7101;
  assign n7159 = ~controllable_BtoR_REQ1 & ~n7158;
  assign n7160 = ~n7100 & ~n7159;
  assign n7161 = ~controllable_BtoR_REQ0 & ~n7160;
  assign n7162 = ~controllable_BtoR_REQ0 & ~n7161;
  assign n7163 = ~i_RtoB_ACK0 & ~n7162;
  assign n7164 = ~n7093 & ~n7163;
  assign n7165 = ~controllable_DEQ & ~n7164;
  assign n7166 = ~n7157 & ~n7165;
  assign n7167 = ~i_FULL & ~n7166;
  assign n7168 = ~n7149 & ~n7167;
  assign n7169 = ~i_nEMPTY & ~n7168;
  assign n7170 = ~n7126 & ~n7169;
  assign n7171 = controllable_BtoS_ACK0 & ~n7170;
  assign n7172 = i_StoB_REQ0 & ~n5213;
  assign n7173 = ~controllable_BtoS_ACK13 & ~n5845;
  assign n7174 = i_StoB_REQ13 & ~n7173;
  assign n7175 = ~i_StoB_REQ13 & ~n5823;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = n4466 & ~n7176;
  assign n7178 = ~n5828 & ~n7177;
  assign n7179 = ~i_StoB_REQ0 & ~n7178;
  assign n7180 = ~n7172 & ~n7179;
  assign n7181 = ~i_StoB_REQ14 & ~n7180;
  assign n7182 = ~i_StoB_REQ14 & ~n7181;
  assign n7183 = controllable_BtoS_ACK14 & ~n7182;
  assign n7184 = ~i_StoB_REQ13 & ~n5844;
  assign n7185 = ~n7174 & ~n7184;
  assign n7186 = n4466 & ~n7185;
  assign n7187 = ~n5849 & ~n7186;
  assign n7188 = ~i_StoB_REQ0 & ~n7187;
  assign n7189 = ~n7172 & ~n7188;
  assign n7190 = i_StoB_REQ14 & ~n7189;
  assign n7191 = ~n7181 & ~n7190;
  assign n7192 = ~controllable_BtoS_ACK14 & ~n7191;
  assign n7193 = ~n7183 & ~n7192;
  assign n7194 = controllable_ENQ & ~n7193;
  assign n7195 = controllable_ENQ & ~n7194;
  assign n7196 = i_RtoB_ACK1 & ~n7195;
  assign n7197 = i_StoB_REQ14 & ~n5318;
  assign n7198 = ~i_StoB_REQ13 & ~n6497;
  assign n7199 = ~n6542 & ~n7198;
  assign n7200 = n4466 & ~n7199;
  assign n7201 = ~n6498 & ~n6548;
  assign n7202 = ~i_StoB_REQ13 & ~n7201;
  assign n7203 = ~n6542 & ~n7202;
  assign n7204 = ~n4466 & ~n7203;
  assign n7205 = ~n7200 & ~n7204;
  assign n7206 = i_StoB_REQ0 & ~n7205;
  assign n7207 = ~n6490 & ~n6557;
  assign n7208 = i_StoB_REQ13 & ~n7207;
  assign n7209 = ~i_StoB_REQ13 & ~n6522;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = n4466 & ~n7210;
  assign n7212 = ~n6527 & ~n7211;
  assign n7213 = ~i_StoB_REQ0 & ~n7212;
  assign n7214 = ~n7206 & ~n7213;
  assign n7215 = ~i_StoB_REQ14 & ~n7214;
  assign n7216 = ~n7197 & ~n7215;
  assign n7217 = controllable_BtoS_ACK14 & ~n7216;
  assign n7218 = ~n6540 & ~n6557;
  assign n7219 = i_StoB_REQ13 & ~n7218;
  assign n7220 = ~i_StoB_REQ13 & ~n6556;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = n4466 & ~n7221;
  assign n7223 = ~n6561 & ~n7222;
  assign n7224 = ~i_StoB_REQ0 & ~n7223;
  assign n7225 = ~n7206 & ~n7224;
  assign n7226 = i_StoB_REQ14 & ~n7225;
  assign n7227 = ~n7215 & ~n7226;
  assign n7228 = ~controllable_BtoS_ACK14 & ~n7227;
  assign n7229 = ~n7217 & ~n7228;
  assign n7230 = controllable_ENQ & ~n7229;
  assign n7231 = controllable_ENQ & ~n7230;
  assign n7232 = ~i_RtoB_ACK1 & ~n7231;
  assign n7233 = ~n7196 & ~n7232;
  assign n7234 = controllable_BtoR_REQ1 & ~n7233;
  assign n7235 = ~i_StoB_REQ14 & ~n7225;
  assign n7236 = ~n5322 & ~n7235;
  assign n7237 = controllable_BtoS_ACK14 & ~n7236;
  assign n7238 = ~controllable_BtoS_ACK14 & ~n7225;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = controllable_ENQ & ~n7239;
  assign n7241 = controllable_ENQ & ~n7240;
  assign n7242 = ~controllable_BtoR_REQ1 & ~n7241;
  assign n7243 = ~n7234 & ~n7242;
  assign n7244 = ~controllable_BtoR_REQ0 & ~n7243;
  assign n7245 = ~controllable_BtoR_REQ0 & ~n7244;
  assign n7246 = i_RtoB_ACK0 & ~n7245;
  assign n7247 = ~i_StoB_REQ13 & ~n6748;
  assign n7248 = ~n6751 & ~n7247;
  assign n7249 = n4466 & ~n7248;
  assign n7250 = ~n6755 & ~n7249;
  assign n7251 = ~i_StoB_REQ14 & ~n7250;
  assign n7252 = ~n5322 & ~n7251;
  assign n7253 = controllable_BtoS_ACK14 & ~n7252;
  assign n7254 = ~controllable_BtoS_ACK14 & ~n7250;
  assign n7255 = ~n7253 & ~n7254;
  assign n7256 = controllable_ENQ & ~n7255;
  assign n7257 = ~controllable_ENQ & ~n7193;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = i_RtoB_ACK1 & ~n7258;
  assign n7260 = ~controllable_ENQ & ~n7229;
  assign n7261 = ~n7256 & ~n7260;
  assign n7262 = ~i_RtoB_ACK1 & ~n7261;
  assign n7263 = ~n7259 & ~n7262;
  assign n7264 = controllable_BtoR_REQ1 & ~n7263;
  assign n7265 = i_RtoB_ACK1 & ~n7241;
  assign n7266 = ~controllable_ENQ & ~n7239;
  assign n7267 = ~n7256 & ~n7266;
  assign n7268 = ~i_RtoB_ACK1 & ~n7267;
  assign n7269 = ~n7265 & ~n7268;
  assign n7270 = ~controllable_BtoR_REQ1 & ~n7269;
  assign n7271 = ~n7264 & ~n7270;
  assign n7272 = ~controllable_BtoR_REQ0 & ~n7271;
  assign n7273 = ~controllable_BtoR_REQ0 & ~n7272;
  assign n7274 = ~i_RtoB_ACK0 & ~n7273;
  assign n7275 = ~n7246 & ~n7274;
  assign n7276 = controllable_DEQ & ~n7275;
  assign n7277 = i_RtoB_ACK1 & ~n7193;
  assign n7278 = ~i_RtoB_ACK1 & ~n7229;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = controllable_BtoR_REQ1 & ~n7279;
  assign n7281 = ~controllable_BtoR_REQ1 & ~n7239;
  assign n7282 = ~n7280 & ~n7281;
  assign n7283 = ~controllable_BtoR_REQ0 & ~n7282;
  assign n7284 = ~controllable_BtoR_REQ0 & ~n7283;
  assign n7285 = i_RtoB_ACK0 & ~n7284;
  assign n7286 = controllable_BtoR_REQ1 & ~n7255;
  assign n7287 = i_RtoB_ACK1 & ~n7239;
  assign n7288 = ~i_RtoB_ACK1 & ~n7255;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = ~controllable_BtoR_REQ1 & ~n7289;
  assign n7291 = ~n7286 & ~n7290;
  assign n7292 = ~controllable_BtoR_REQ0 & ~n7291;
  assign n7293 = ~controllable_BtoR_REQ0 & ~n7292;
  assign n7294 = ~i_RtoB_ACK0 & ~n7293;
  assign n7295 = ~n7285 & ~n7294;
  assign n7296 = ~controllable_DEQ & ~n7295;
  assign n7297 = ~n7276 & ~n7296;
  assign n7298 = i_FULL & ~n7297;
  assign n7299 = ~n7240 & ~n7257;
  assign n7300 = i_RtoB_ACK1 & ~n7299;
  assign n7301 = ~n7240 & ~n7260;
  assign n7302 = ~i_RtoB_ACK1 & ~n7301;
  assign n7303 = ~n7300 & ~n7302;
  assign n7304 = controllable_BtoR_REQ1 & ~n7303;
  assign n7305 = ~i_RtoB_ACK1 & ~n7239;
  assign n7306 = ~n7265 & ~n7305;
  assign n7307 = ~controllable_BtoR_REQ1 & ~n7306;
  assign n7308 = ~n7304 & ~n7307;
  assign n7309 = ~controllable_BtoR_REQ0 & ~n7308;
  assign n7310 = ~controllable_BtoR_REQ0 & ~n7309;
  assign n7311 = ~i_RtoB_ACK0 & ~n7310;
  assign n7312 = ~n7246 & ~n7311;
  assign n7313 = controllable_DEQ & ~n7312;
  assign n7314 = controllable_BtoR_REQ1 & ~n7267;
  assign n7315 = ~n7268 & ~n7287;
  assign n7316 = ~controllable_BtoR_REQ1 & ~n7315;
  assign n7317 = ~n7314 & ~n7316;
  assign n7318 = ~controllable_BtoR_REQ0 & ~n7317;
  assign n7319 = ~controllable_BtoR_REQ0 & ~n7318;
  assign n7320 = ~i_RtoB_ACK0 & ~n7319;
  assign n7321 = ~n7285 & ~n7320;
  assign n7322 = ~controllable_DEQ & ~n7321;
  assign n7323 = ~n7313 & ~n7322;
  assign n7324 = ~i_FULL & ~n7323;
  assign n7325 = ~n7298 & ~n7324;
  assign n7326 = i_nEMPTY & ~n7325;
  assign n7327 = ~controllable_ENQ & ~n7257;
  assign n7328 = i_RtoB_ACK1 & ~n7327;
  assign n7329 = ~controllable_ENQ & ~n7260;
  assign n7330 = ~i_RtoB_ACK1 & ~n7329;
  assign n7331 = ~n7328 & ~n7330;
  assign n7332 = controllable_BtoR_REQ1 & ~n7331;
  assign n7333 = ~controllable_ENQ & ~n7266;
  assign n7334 = ~i_RtoB_ACK1 & ~n7333;
  assign n7335 = ~i_RtoB_ACK1 & ~n7334;
  assign n7336 = ~controllable_BtoR_REQ1 & ~n7335;
  assign n7337 = ~n7332 & ~n7336;
  assign n7338 = ~controllable_BtoR_REQ0 & ~n7337;
  assign n7339 = ~controllable_BtoR_REQ0 & ~n7338;
  assign n7340 = ~i_RtoB_ACK0 & ~n7339;
  assign n7341 = ~i_RtoB_ACK0 & ~n7340;
  assign n7342 = controllable_DEQ & ~n7341;
  assign n7343 = controllable_ENQ & ~n7256;
  assign n7344 = controllable_BtoR_REQ1 & ~n7343;
  assign n7345 = ~i_RtoB_ACK1 & ~n7343;
  assign n7346 = ~n7265 & ~n7345;
  assign n7347 = ~controllable_BtoR_REQ1 & ~n7346;
  assign n7348 = ~n7344 & ~n7347;
  assign n7349 = ~controllable_BtoR_REQ0 & ~n7348;
  assign n7350 = ~controllable_BtoR_REQ0 & ~n7349;
  assign n7351 = ~i_RtoB_ACK0 & ~n7350;
  assign n7352 = ~n7246 & ~n7351;
  assign n7353 = ~controllable_DEQ & ~n7352;
  assign n7354 = ~n7342 & ~n7353;
  assign n7355 = i_FULL & ~n7354;
  assign n7356 = ~i_RtoB_ACK1 & ~n7305;
  assign n7357 = ~controllable_BtoR_REQ1 & ~n7356;
  assign n7358 = ~n7280 & ~n7357;
  assign n7359 = ~controllable_BtoR_REQ0 & ~n7358;
  assign n7360 = ~controllable_BtoR_REQ0 & ~n7359;
  assign n7361 = ~i_RtoB_ACK0 & ~n7360;
  assign n7362 = ~i_RtoB_ACK0 & ~n7361;
  assign n7363 = controllable_DEQ & ~n7362;
  assign n7364 = ~n7262 & ~n7265;
  assign n7365 = ~controllable_BtoR_REQ1 & ~n7364;
  assign n7366 = ~n7264 & ~n7365;
  assign n7367 = ~controllable_BtoR_REQ0 & ~n7366;
  assign n7368 = ~controllable_BtoR_REQ0 & ~n7367;
  assign n7369 = ~i_RtoB_ACK0 & ~n7368;
  assign n7370 = ~n7246 & ~n7369;
  assign n7371 = ~controllable_DEQ & ~n7370;
  assign n7372 = ~n7363 & ~n7371;
  assign n7373 = ~i_FULL & ~n7372;
  assign n7374 = ~n7355 & ~n7373;
  assign n7375 = ~i_nEMPTY & ~n7374;
  assign n7376 = ~n7326 & ~n7375;
  assign n7377 = ~controllable_BtoS_ACK0 & ~n7376;
  assign n7378 = ~n7171 & ~n7377;
  assign n7379 = ~n4465 & ~n7378;
  assign n7380 = ~n7053 & ~n7379;
  assign n7381 = ~i_StoB_REQ10 & ~n7380;
  assign n7382 = ~n5417 & ~n7381;
  assign n7383 = controllable_BtoS_ACK10 & ~n7382;
  assign n7384 = ~i_StoB_REQ14 & ~n5852;
  assign n7385 = ~i_StoB_REQ14 & ~n7384;
  assign n7386 = controllable_BtoS_ACK14 & ~n7385;
  assign n7387 = ~controllable_BtoS_ACK14 & ~n5852;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = controllable_ENQ & ~n7388;
  assign n7390 = controllable_ENQ & ~n7389;
  assign n7391 = i_RtoB_ACK1 & ~n7390;
  assign n7392 = ~i_RtoB_ACK1 & ~n6580;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 = controllable_BtoR_REQ1 & ~n7393;
  assign n7395 = ~n6581 & ~n7394;
  assign n7396 = ~controllable_BtoR_REQ0 & ~n7395;
  assign n7397 = ~controllable_BtoR_REQ0 & ~n7396;
  assign n7398 = i_RtoB_ACK0 & ~n7397;
  assign n7399 = ~controllable_ENQ & ~n7388;
  assign n7400 = ~n6764 & ~n7399;
  assign n7401 = i_RtoB_ACK1 & ~n7400;
  assign n7402 = ~n6776 & ~n7401;
  assign n7403 = controllable_BtoR_REQ1 & ~n7402;
  assign n7404 = ~n6778 & ~n7403;
  assign n7405 = ~controllable_BtoR_REQ0 & ~n7404;
  assign n7406 = ~controllable_BtoR_REQ0 & ~n7405;
  assign n7407 = ~i_RtoB_ACK0 & ~n7406;
  assign n7408 = ~n7398 & ~n7407;
  assign n7409 = controllable_DEQ & ~n7408;
  assign n7410 = i_RtoB_ACK1 & ~n7388;
  assign n7411 = ~n6813 & ~n7410;
  assign n7412 = controllable_BtoR_REQ1 & ~n7411;
  assign n7413 = ~n6789 & ~n7412;
  assign n7414 = ~controllable_BtoR_REQ0 & ~n7413;
  assign n7415 = ~controllable_BtoR_REQ0 & ~n7414;
  assign n7416 = i_RtoB_ACK0 & ~n7415;
  assign n7417 = ~n6802 & ~n7416;
  assign n7418 = ~controllable_DEQ & ~n7417;
  assign n7419 = ~n7409 & ~n7418;
  assign n7420 = i_FULL & ~n7419;
  assign n7421 = ~n6579 & ~n7399;
  assign n7422 = i_RtoB_ACK1 & ~n7421;
  assign n7423 = ~n6813 & ~n7422;
  assign n7424 = controllable_BtoR_REQ1 & ~n7423;
  assign n7425 = ~n6815 & ~n7424;
  assign n7426 = ~controllable_BtoR_REQ0 & ~n7425;
  assign n7427 = ~controllable_BtoR_REQ0 & ~n7426;
  assign n7428 = ~i_RtoB_ACK0 & ~n7427;
  assign n7429 = ~n7398 & ~n7428;
  assign n7430 = controllable_DEQ & ~n7429;
  assign n7431 = ~n6828 & ~n7416;
  assign n7432 = ~controllable_DEQ & ~n7431;
  assign n7433 = ~n7430 & ~n7432;
  assign n7434 = ~i_FULL & ~n7433;
  assign n7435 = ~n7420 & ~n7434;
  assign n7436 = i_nEMPTY & ~n7435;
  assign n7437 = ~controllable_ENQ & ~n7399;
  assign n7438 = i_RtoB_ACK1 & ~n7437;
  assign n7439 = ~n6842 & ~n7438;
  assign n7440 = controllable_BtoR_REQ1 & ~n7439;
  assign n7441 = ~n6844 & ~n7440;
  assign n7442 = ~controllable_BtoR_REQ0 & ~n7441;
  assign n7443 = ~controllable_BtoR_REQ0 & ~n7442;
  assign n7444 = ~i_RtoB_ACK0 & ~n7443;
  assign n7445 = ~i_RtoB_ACK0 & ~n7444;
  assign n7446 = controllable_DEQ & ~n7445;
  assign n7447 = ~n6859 & ~n7398;
  assign n7448 = ~controllable_DEQ & ~n7447;
  assign n7449 = ~n7446 & ~n7448;
  assign n7450 = i_FULL & ~n7449;
  assign n7451 = ~n6865 & ~n7412;
  assign n7452 = ~controllable_BtoR_REQ0 & ~n7451;
  assign n7453 = ~controllable_BtoR_REQ0 & ~n7452;
  assign n7454 = ~i_RtoB_ACK0 & ~n7453;
  assign n7455 = ~i_RtoB_ACK0 & ~n7454;
  assign n7456 = controllable_DEQ & ~n7455;
  assign n7457 = ~controllable_DEQ & ~n7408;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = ~i_FULL & ~n7458;
  assign n7460 = ~n7450 & ~n7459;
  assign n7461 = ~i_nEMPTY & ~n7460;
  assign n7462 = ~n7436 & ~n7461;
  assign n7463 = controllable_BtoS_ACK0 & ~n7462;
  assign n7464 = ~i_StoB_REQ14 & ~n5850;
  assign n7465 = ~i_StoB_REQ14 & ~n7464;
  assign n7466 = controllable_BtoS_ACK14 & ~n7465;
  assign n7467 = ~controllable_BtoS_ACK14 & ~n5850;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = controllable_ENQ & ~n7468;
  assign n7470 = controllable_ENQ & ~n7469;
  assign n7471 = i_RtoB_ACK1 & ~n7470;
  assign n7472 = ~i_RtoB_ACK1 & ~n6919;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = controllable_BtoR_REQ1 & ~n7473;
  assign n7475 = ~n6920 & ~n7474;
  assign n7476 = ~controllable_BtoR_REQ0 & ~n7475;
  assign n7477 = ~controllable_BtoR_REQ0 & ~n7476;
  assign n7478 = i_RtoB_ACK0 & ~n7477;
  assign n7479 = ~controllable_ENQ & ~n7468;
  assign n7480 = ~n6930 & ~n7479;
  assign n7481 = i_RtoB_ACK1 & ~n7480;
  assign n7482 = ~n6942 & ~n7481;
  assign n7483 = controllable_BtoR_REQ1 & ~n7482;
  assign n7484 = ~n6944 & ~n7483;
  assign n7485 = ~controllable_BtoR_REQ0 & ~n7484;
  assign n7486 = ~controllable_BtoR_REQ0 & ~n7485;
  assign n7487 = ~i_RtoB_ACK0 & ~n7486;
  assign n7488 = ~n7478 & ~n7487;
  assign n7489 = controllable_DEQ & ~n7488;
  assign n7490 = i_RtoB_ACK1 & ~n7468;
  assign n7491 = ~n6979 & ~n7490;
  assign n7492 = controllable_BtoR_REQ1 & ~n7491;
  assign n7493 = ~n6955 & ~n7492;
  assign n7494 = ~controllable_BtoR_REQ0 & ~n7493;
  assign n7495 = ~controllable_BtoR_REQ0 & ~n7494;
  assign n7496 = i_RtoB_ACK0 & ~n7495;
  assign n7497 = ~n6968 & ~n7496;
  assign n7498 = ~controllable_DEQ & ~n7497;
  assign n7499 = ~n7489 & ~n7498;
  assign n7500 = i_FULL & ~n7499;
  assign n7501 = ~n6918 & ~n7479;
  assign n7502 = i_RtoB_ACK1 & ~n7501;
  assign n7503 = ~n6979 & ~n7502;
  assign n7504 = controllable_BtoR_REQ1 & ~n7503;
  assign n7505 = ~n6981 & ~n7504;
  assign n7506 = ~controllable_BtoR_REQ0 & ~n7505;
  assign n7507 = ~controllable_BtoR_REQ0 & ~n7506;
  assign n7508 = ~i_RtoB_ACK0 & ~n7507;
  assign n7509 = ~n7478 & ~n7508;
  assign n7510 = controllable_DEQ & ~n7509;
  assign n7511 = ~n6994 & ~n7496;
  assign n7512 = ~controllable_DEQ & ~n7511;
  assign n7513 = ~n7510 & ~n7512;
  assign n7514 = ~i_FULL & ~n7513;
  assign n7515 = ~n7500 & ~n7514;
  assign n7516 = i_nEMPTY & ~n7515;
  assign n7517 = ~controllable_ENQ & ~n7479;
  assign n7518 = i_RtoB_ACK1 & ~n7517;
  assign n7519 = ~n7008 & ~n7518;
  assign n7520 = controllable_BtoR_REQ1 & ~n7519;
  assign n7521 = ~n7010 & ~n7520;
  assign n7522 = ~controllable_BtoR_REQ0 & ~n7521;
  assign n7523 = ~controllable_BtoR_REQ0 & ~n7522;
  assign n7524 = ~i_RtoB_ACK0 & ~n7523;
  assign n7525 = ~i_RtoB_ACK0 & ~n7524;
  assign n7526 = controllable_DEQ & ~n7525;
  assign n7527 = ~n7025 & ~n7478;
  assign n7528 = ~controllable_DEQ & ~n7527;
  assign n7529 = ~n7526 & ~n7528;
  assign n7530 = i_FULL & ~n7529;
  assign n7531 = ~n7031 & ~n7492;
  assign n7532 = ~controllable_BtoR_REQ0 & ~n7531;
  assign n7533 = ~controllable_BtoR_REQ0 & ~n7532;
  assign n7534 = ~i_RtoB_ACK0 & ~n7533;
  assign n7535 = ~i_RtoB_ACK0 & ~n7534;
  assign n7536 = controllable_DEQ & ~n7535;
  assign n7537 = ~controllable_DEQ & ~n7488;
  assign n7538 = ~n7536 & ~n7537;
  assign n7539 = ~i_FULL & ~n7538;
  assign n7540 = ~n7530 & ~n7539;
  assign n7541 = ~i_nEMPTY & ~n7540;
  assign n7542 = ~n7516 & ~n7541;
  assign n7543 = ~controllable_BtoS_ACK0 & ~n7542;
  assign n7544 = ~n7463 & ~n7543;
  assign n7545 = n4465 & ~n7544;
  assign n7546 = ~i_RtoB_ACK1 & ~n7088;
  assign n7547 = ~n5237 & ~n7546;
  assign n7548 = controllable_BtoR_REQ1 & ~n7547;
  assign n7549 = ~n7089 & ~n7548;
  assign n7550 = ~controllable_BtoR_REQ0 & ~n7549;
  assign n7551 = ~controllable_BtoR_REQ0 & ~n7550;
  assign n7552 = i_RtoB_ACK0 & ~n7551;
  assign n7553 = ~n5271 & ~n7087;
  assign n7554 = i_RtoB_ACK1 & ~n7553;
  assign n7555 = ~n7102 & ~n7554;
  assign n7556 = controllable_BtoR_REQ1 & ~n7555;
  assign n7557 = ~n7104 & ~n7556;
  assign n7558 = ~controllable_BtoR_REQ0 & ~n7557;
  assign n7559 = ~controllable_BtoR_REQ0 & ~n7558;
  assign n7560 = ~i_RtoB_ACK0 & ~n7559;
  assign n7561 = ~n7552 & ~n7560;
  assign n7562 = controllable_DEQ & ~n7561;
  assign n7563 = i_RtoB_ACK1 & ~n5229;
  assign n7564 = ~n7102 & ~n7563;
  assign n7565 = controllable_BtoR_REQ1 & ~n7564;
  assign n7566 = ~n7115 & ~n7565;
  assign n7567 = ~controllable_BtoR_REQ0 & ~n7566;
  assign n7568 = ~controllable_BtoR_REQ0 & ~n7567;
  assign n7569 = i_RtoB_ACK0 & ~n7568;
  assign n7570 = ~n7122 & ~n7569;
  assign n7571 = ~controllable_DEQ & ~n7570;
  assign n7572 = ~n7562 & ~n7571;
  assign n7573 = i_nEMPTY & ~n7572;
  assign n7574 = i_RtoB_ACK1 & ~n5272;
  assign n7575 = ~n7134 & ~n7574;
  assign n7576 = controllable_BtoR_REQ1 & ~n7575;
  assign n7577 = ~n7136 & ~n7576;
  assign n7578 = ~controllable_BtoR_REQ0 & ~n7577;
  assign n7579 = ~controllable_BtoR_REQ0 & ~n7578;
  assign n7580 = ~i_RtoB_ACK0 & ~n7579;
  assign n7581 = ~i_RtoB_ACK0 & ~n7580;
  assign n7582 = controllable_DEQ & ~n7581;
  assign n7583 = ~n7145 & ~n7552;
  assign n7584 = ~controllable_DEQ & ~n7583;
  assign n7585 = ~n7582 & ~n7584;
  assign n7586 = i_FULL & ~n7585;
  assign n7587 = ~n7151 & ~n7565;
  assign n7588 = ~controllable_BtoR_REQ0 & ~n7587;
  assign n7589 = ~controllable_BtoR_REQ0 & ~n7588;
  assign n7590 = ~i_RtoB_ACK0 & ~n7589;
  assign n7591 = ~i_RtoB_ACK0 & ~n7590;
  assign n7592 = controllable_DEQ & ~n7591;
  assign n7593 = ~controllable_DEQ & ~n7561;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = ~i_FULL & ~n7594;
  assign n7596 = ~n7586 & ~n7595;
  assign n7597 = ~i_nEMPTY & ~n7596;
  assign n7598 = ~n7573 & ~n7597;
  assign n7599 = controllable_BtoS_ACK0 & ~n7598;
  assign n7600 = ~i_StoB_REQ14 & ~n7189;
  assign n7601 = ~i_StoB_REQ14 & ~n7600;
  assign n7602 = controllable_BtoS_ACK14 & ~n7601;
  assign n7603 = ~controllable_BtoS_ACK14 & ~n7189;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = controllable_ENQ & ~n7604;
  assign n7606 = controllable_ENQ & ~n7605;
  assign n7607 = i_RtoB_ACK1 & ~n7606;
  assign n7608 = ~i_RtoB_ACK1 & ~n7241;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = controllable_BtoR_REQ1 & ~n7609;
  assign n7611 = ~n7242 & ~n7610;
  assign n7612 = ~controllable_BtoR_REQ0 & ~n7611;
  assign n7613 = ~controllable_BtoR_REQ0 & ~n7612;
  assign n7614 = i_RtoB_ACK0 & ~n7613;
  assign n7615 = ~controllable_ENQ & ~n7604;
  assign n7616 = ~n7256 & ~n7615;
  assign n7617 = i_RtoB_ACK1 & ~n7616;
  assign n7618 = ~n7268 & ~n7617;
  assign n7619 = controllable_BtoR_REQ1 & ~n7618;
  assign n7620 = ~n7270 & ~n7619;
  assign n7621 = ~controllable_BtoR_REQ0 & ~n7620;
  assign n7622 = ~controllable_BtoR_REQ0 & ~n7621;
  assign n7623 = ~i_RtoB_ACK0 & ~n7622;
  assign n7624 = ~n7614 & ~n7623;
  assign n7625 = controllable_DEQ & ~n7624;
  assign n7626 = i_RtoB_ACK1 & ~n7604;
  assign n7627 = ~n7305 & ~n7626;
  assign n7628 = controllable_BtoR_REQ1 & ~n7627;
  assign n7629 = ~n7281 & ~n7628;
  assign n7630 = ~controllable_BtoR_REQ0 & ~n7629;
  assign n7631 = ~controllable_BtoR_REQ0 & ~n7630;
  assign n7632 = i_RtoB_ACK0 & ~n7631;
  assign n7633 = ~n7294 & ~n7632;
  assign n7634 = ~controllable_DEQ & ~n7633;
  assign n7635 = ~n7625 & ~n7634;
  assign n7636 = i_FULL & ~n7635;
  assign n7637 = ~n7240 & ~n7615;
  assign n7638 = i_RtoB_ACK1 & ~n7637;
  assign n7639 = ~n7305 & ~n7638;
  assign n7640 = controllable_BtoR_REQ1 & ~n7639;
  assign n7641 = ~n7307 & ~n7640;
  assign n7642 = ~controllable_BtoR_REQ0 & ~n7641;
  assign n7643 = ~controllable_BtoR_REQ0 & ~n7642;
  assign n7644 = ~i_RtoB_ACK0 & ~n7643;
  assign n7645 = ~n7614 & ~n7644;
  assign n7646 = controllable_DEQ & ~n7645;
  assign n7647 = ~n7320 & ~n7632;
  assign n7648 = ~controllable_DEQ & ~n7647;
  assign n7649 = ~n7646 & ~n7648;
  assign n7650 = ~i_FULL & ~n7649;
  assign n7651 = ~n7636 & ~n7650;
  assign n7652 = i_nEMPTY & ~n7651;
  assign n7653 = ~controllable_ENQ & ~n7615;
  assign n7654 = i_RtoB_ACK1 & ~n7653;
  assign n7655 = ~n7334 & ~n7654;
  assign n7656 = controllable_BtoR_REQ1 & ~n7655;
  assign n7657 = ~n7336 & ~n7656;
  assign n7658 = ~controllable_BtoR_REQ0 & ~n7657;
  assign n7659 = ~controllable_BtoR_REQ0 & ~n7658;
  assign n7660 = ~i_RtoB_ACK0 & ~n7659;
  assign n7661 = ~i_RtoB_ACK0 & ~n7660;
  assign n7662 = controllable_DEQ & ~n7661;
  assign n7663 = ~n7351 & ~n7614;
  assign n7664 = ~controllable_DEQ & ~n7663;
  assign n7665 = ~n7662 & ~n7664;
  assign n7666 = i_FULL & ~n7665;
  assign n7667 = ~n7357 & ~n7628;
  assign n7668 = ~controllable_BtoR_REQ0 & ~n7667;
  assign n7669 = ~controllable_BtoR_REQ0 & ~n7668;
  assign n7670 = ~i_RtoB_ACK0 & ~n7669;
  assign n7671 = ~i_RtoB_ACK0 & ~n7670;
  assign n7672 = controllable_DEQ & ~n7671;
  assign n7673 = ~controllable_DEQ & ~n7624;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = ~i_FULL & ~n7674;
  assign n7676 = ~n7666 & ~n7675;
  assign n7677 = ~i_nEMPTY & ~n7676;
  assign n7678 = ~n7652 & ~n7677;
  assign n7679 = ~controllable_BtoS_ACK0 & ~n7678;
  assign n7680 = ~n7599 & ~n7679;
  assign n7681 = ~n4465 & ~n7680;
  assign n7682 = ~n7545 & ~n7681;
  assign n7683 = i_StoB_REQ10 & ~n7682;
  assign n7684 = ~n7381 & ~n7683;
  assign n7685 = ~controllable_BtoS_ACK10 & ~n7684;
  assign n7686 = ~n7383 & ~n7685;
  assign n7687 = n4464 & ~n7686;
  assign n7688 = ~i_StoB_REQ0 & ~n5311;
  assign n7689 = ~i_StoB_REQ0 & ~n7688;
  assign n7690 = i_StoB_REQ14 & ~n7689;
  assign n7691 = ~i_StoB_REQ0 & ~n5317;
  assign n7692 = ~i_StoB_REQ14 & ~n7691;
  assign n7693 = ~n7690 & ~n7692;
  assign n7694 = ~controllable_BtoS_ACK14 & ~n7693;
  assign n7695 = ~n5211 & ~n7694;
  assign n7696 = controllable_ENQ & ~n7695;
  assign n7697 = controllable_ENQ & ~n7696;
  assign n7698 = ~i_RtoB_ACK1 & ~n7697;
  assign n7699 = ~i_RtoB_ACK1 & ~n7698;
  assign n7700 = controllable_BtoR_REQ1 & ~n7699;
  assign n7701 = ~controllable_BtoS_ACK14 & ~n7689;
  assign n7702 = ~n5227 & ~n7701;
  assign n7703 = controllable_ENQ & ~n7702;
  assign n7704 = controllable_ENQ & ~n7703;
  assign n7705 = ~controllable_BtoR_REQ1 & ~n7704;
  assign n7706 = ~n7700 & ~n7705;
  assign n7707 = ~controllable_BtoR_REQ0 & ~n7706;
  assign n7708 = ~controllable_BtoR_REQ0 & ~n7707;
  assign n7709 = i_RtoB_ACK0 & ~n7708;
  assign n7710 = i_RtoB_ACK1 & ~n7704;
  assign n7711 = ~controllable_ENQ & ~n7695;
  assign n7712 = ~n7703 & ~n7711;
  assign n7713 = ~i_RtoB_ACK1 & ~n7712;
  assign n7714 = ~n7710 & ~n7713;
  assign n7715 = controllable_BtoR_REQ1 & ~n7714;
  assign n7716 = ~i_RtoB_ACK1 & ~n7702;
  assign n7717 = ~n7710 & ~n7716;
  assign n7718 = ~controllable_BtoR_REQ1 & ~n7717;
  assign n7719 = ~n7715 & ~n7718;
  assign n7720 = ~controllable_BtoR_REQ0 & ~n7719;
  assign n7721 = ~controllable_BtoR_REQ0 & ~n7720;
  assign n7722 = ~i_RtoB_ACK0 & ~n7721;
  assign n7723 = ~n7709 & ~n7722;
  assign n7724 = controllable_DEQ & ~n7723;
  assign n7725 = ~i_RtoB_ACK1 & ~n7695;
  assign n7726 = ~i_RtoB_ACK1 & ~n7725;
  assign n7727 = controllable_BtoR_REQ1 & ~n7726;
  assign n7728 = ~controllable_BtoR_REQ1 & ~n7702;
  assign n7729 = ~n7727 & ~n7728;
  assign n7730 = ~controllable_BtoR_REQ0 & ~n7729;
  assign n7731 = ~controllable_BtoR_REQ0 & ~n7730;
  assign n7732 = i_RtoB_ACK0 & ~n7731;
  assign n7733 = ~controllable_BtoR_REQ0 & ~n7702;
  assign n7734 = ~controllable_BtoR_REQ0 & ~n7733;
  assign n7735 = ~i_RtoB_ACK0 & ~n7734;
  assign n7736 = ~n7732 & ~n7735;
  assign n7737 = ~controllable_DEQ & ~n7736;
  assign n7738 = ~n7724 & ~n7737;
  assign n7739 = i_nEMPTY & ~n7738;
  assign n7740 = ~controllable_ENQ & ~n7711;
  assign n7741 = ~i_RtoB_ACK1 & ~n7740;
  assign n7742 = ~i_RtoB_ACK1 & ~n7741;
  assign n7743 = controllable_BtoR_REQ1 & ~n7742;
  assign n7744 = ~controllable_ENQ & ~n7702;
  assign n7745 = ~controllable_ENQ & ~n7744;
  assign n7746 = ~i_RtoB_ACK1 & ~n7745;
  assign n7747 = ~i_RtoB_ACK1 & ~n7746;
  assign n7748 = ~controllable_BtoR_REQ1 & ~n7747;
  assign n7749 = ~n7743 & ~n7748;
  assign n7750 = ~controllable_BtoR_REQ0 & ~n7749;
  assign n7751 = ~controllable_BtoR_REQ0 & ~n7750;
  assign n7752 = ~i_RtoB_ACK0 & ~n7751;
  assign n7753 = ~i_RtoB_ACK0 & ~n7752;
  assign n7754 = controllable_DEQ & ~n7753;
  assign n7755 = ~controllable_BtoR_REQ0 & ~n7704;
  assign n7756 = ~controllable_BtoR_REQ0 & ~n7755;
  assign n7757 = ~i_RtoB_ACK0 & ~n7756;
  assign n7758 = ~n7709 & ~n7757;
  assign n7759 = ~controllable_DEQ & ~n7758;
  assign n7760 = ~n7754 & ~n7759;
  assign n7761 = i_FULL & ~n7760;
  assign n7762 = ~i_RtoB_ACK1 & ~n7716;
  assign n7763 = ~controllable_BtoR_REQ1 & ~n7762;
  assign n7764 = ~n7727 & ~n7763;
  assign n7765 = ~controllable_BtoR_REQ0 & ~n7764;
  assign n7766 = ~controllable_BtoR_REQ0 & ~n7765;
  assign n7767 = ~i_RtoB_ACK0 & ~n7766;
  assign n7768 = ~i_RtoB_ACK0 & ~n7767;
  assign n7769 = controllable_DEQ & ~n7768;
  assign n7770 = ~controllable_BtoR_REQ0 & ~n7714;
  assign n7771 = ~controllable_BtoR_REQ0 & ~n7770;
  assign n7772 = ~i_RtoB_ACK0 & ~n7771;
  assign n7773 = ~n7709 & ~n7772;
  assign n7774 = ~controllable_DEQ & ~n7773;
  assign n7775 = ~n7769 & ~n7774;
  assign n7776 = ~i_FULL & ~n7775;
  assign n7777 = ~n7761 & ~n7776;
  assign n7778 = ~i_nEMPTY & ~n7777;
  assign n7779 = ~n7739 & ~n7778;
  assign n7780 = controllable_BtoS_ACK0 & ~n7779;
  assign n7781 = ~n5207 & ~n7172;
  assign n7782 = ~i_StoB_REQ14 & ~n7781;
  assign n7783 = ~i_StoB_REQ14 & ~n7782;
  assign n7784 = controllable_BtoS_ACK14 & ~n7783;
  assign n7785 = ~n5324 & ~n7784;
  assign n7786 = controllable_ENQ & ~n7785;
  assign n7787 = controllable_ENQ & ~n7786;
  assign n7788 = ~i_RtoB_ACK1 & ~n7787;
  assign n7789 = ~i_RtoB_ACK1 & ~n7788;
  assign n7790 = controllable_BtoR_REQ1 & ~n7789;
  assign n7791 = ~i_StoB_REQ14 & ~n5213;
  assign n7792 = ~i_StoB_REQ14 & ~n7791;
  assign n7793 = controllable_BtoS_ACK14 & ~n7792;
  assign n7794 = ~n5334 & ~n7793;
  assign n7795 = controllable_ENQ & ~n7794;
  assign n7796 = controllable_ENQ & ~n7795;
  assign n7797 = ~controllable_BtoR_REQ1 & ~n7796;
  assign n7798 = ~n7790 & ~n7797;
  assign n7799 = ~controllable_BtoR_REQ0 & ~n7798;
  assign n7800 = ~controllable_BtoR_REQ0 & ~n7799;
  assign n7801 = i_RtoB_ACK0 & ~n7800;
  assign n7802 = i_RtoB_ACK1 & ~n7796;
  assign n7803 = ~controllable_ENQ & ~n7785;
  assign n7804 = ~n7795 & ~n7803;
  assign n7805 = ~i_RtoB_ACK1 & ~n7804;
  assign n7806 = ~n7802 & ~n7805;
  assign n7807 = controllable_BtoR_REQ1 & ~n7806;
  assign n7808 = ~i_RtoB_ACK1 & ~n7794;
  assign n7809 = ~n7802 & ~n7808;
  assign n7810 = ~controllable_BtoR_REQ1 & ~n7809;
  assign n7811 = ~n7807 & ~n7810;
  assign n7812 = ~controllable_BtoR_REQ0 & ~n7811;
  assign n7813 = ~controllable_BtoR_REQ0 & ~n7812;
  assign n7814 = ~i_RtoB_ACK0 & ~n7813;
  assign n7815 = ~n7801 & ~n7814;
  assign n7816 = controllable_DEQ & ~n7815;
  assign n7817 = ~i_RtoB_ACK1 & ~n7785;
  assign n7818 = ~i_RtoB_ACK1 & ~n7817;
  assign n7819 = controllable_BtoR_REQ1 & ~n7818;
  assign n7820 = ~controllable_BtoR_REQ1 & ~n7794;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~controllable_BtoR_REQ0 & ~n7821;
  assign n7823 = ~controllable_BtoR_REQ0 & ~n7822;
  assign n7824 = i_RtoB_ACK0 & ~n7823;
  assign n7825 = ~controllable_BtoR_REQ0 & ~n7794;
  assign n7826 = ~controllable_BtoR_REQ0 & ~n7825;
  assign n7827 = ~i_RtoB_ACK0 & ~n7826;
  assign n7828 = ~n7824 & ~n7827;
  assign n7829 = ~controllable_DEQ & ~n7828;
  assign n7830 = ~n7816 & ~n7829;
  assign n7831 = i_nEMPTY & ~n7830;
  assign n7832 = ~controllable_ENQ & ~n7803;
  assign n7833 = ~i_RtoB_ACK1 & ~n7832;
  assign n7834 = ~i_RtoB_ACK1 & ~n7833;
  assign n7835 = controllable_BtoR_REQ1 & ~n7834;
  assign n7836 = ~controllable_ENQ & ~n7794;
  assign n7837 = ~controllable_ENQ & ~n7836;
  assign n7838 = ~i_RtoB_ACK1 & ~n7837;
  assign n7839 = ~i_RtoB_ACK1 & ~n7838;
  assign n7840 = ~controllable_BtoR_REQ1 & ~n7839;
  assign n7841 = ~n7835 & ~n7840;
  assign n7842 = ~controllable_BtoR_REQ0 & ~n7841;
  assign n7843 = ~controllable_BtoR_REQ0 & ~n7842;
  assign n7844 = ~i_RtoB_ACK0 & ~n7843;
  assign n7845 = ~i_RtoB_ACK0 & ~n7844;
  assign n7846 = controllable_DEQ & ~n7845;
  assign n7847 = ~controllable_BtoR_REQ0 & ~n7796;
  assign n7848 = ~controllable_BtoR_REQ0 & ~n7847;
  assign n7849 = ~i_RtoB_ACK0 & ~n7848;
  assign n7850 = ~n7801 & ~n7849;
  assign n7851 = ~controllable_DEQ & ~n7850;
  assign n7852 = ~n7846 & ~n7851;
  assign n7853 = i_FULL & ~n7852;
  assign n7854 = ~i_RtoB_ACK1 & ~n7808;
  assign n7855 = ~controllable_BtoR_REQ1 & ~n7854;
  assign n7856 = ~n7819 & ~n7855;
  assign n7857 = ~controllable_BtoR_REQ0 & ~n7856;
  assign n7858 = ~controllable_BtoR_REQ0 & ~n7857;
  assign n7859 = ~i_RtoB_ACK0 & ~n7858;
  assign n7860 = ~i_RtoB_ACK0 & ~n7859;
  assign n7861 = controllable_DEQ & ~n7860;
  assign n7862 = ~controllable_BtoR_REQ0 & ~n7806;
  assign n7863 = ~controllable_BtoR_REQ0 & ~n7862;
  assign n7864 = ~i_RtoB_ACK0 & ~n7863;
  assign n7865 = ~n7801 & ~n7864;
  assign n7866 = ~controllable_DEQ & ~n7865;
  assign n7867 = ~n7861 & ~n7866;
  assign n7868 = ~i_FULL & ~n7867;
  assign n7869 = ~n7853 & ~n7868;
  assign n7870 = ~i_nEMPTY & ~n7869;
  assign n7871 = ~n7831 & ~n7870;
  assign n7872 = ~controllable_BtoS_ACK0 & ~n7871;
  assign n7873 = ~n7780 & ~n7872;
  assign n7874 = n4465 & ~n7873;
  assign n7875 = ~n5307 & ~n7872;
  assign n7876 = ~n4465 & ~n7875;
  assign n7877 = ~n7874 & ~n7876;
  assign n7878 = i_StoB_REQ10 & ~n7877;
  assign n7879 = ~i_StoB_REQ0 & ~n7179;
  assign n7880 = ~i_StoB_REQ14 & ~n7879;
  assign n7881 = ~n5216 & ~n7880;
  assign n7882 = ~controllable_BtoS_ACK14 & ~n7881;
  assign n7883 = ~n5211 & ~n7882;
  assign n7884 = controllable_ENQ & ~n7883;
  assign n7885 = controllable_ENQ & ~n7884;
  assign n7886 = i_RtoB_ACK1 & ~n7885;
  assign n7887 = i_StoB_REQ14 & ~n7691;
  assign n7888 = i_StoB_REQ0 & ~n5206;
  assign n7889 = ~n7062 & ~n7888;
  assign n7890 = ~i_StoB_REQ14 & ~n7889;
  assign n7891 = ~n7887 & ~n7890;
  assign n7892 = controllable_BtoS_ACK14 & ~n7891;
  assign n7893 = ~i_StoB_REQ0 & ~n7205;
  assign n7894 = ~n5312 & ~n7893;
  assign n7895 = i_StoB_REQ14 & ~n7894;
  assign n7896 = ~n7056 & ~n7213;
  assign n7897 = ~i_StoB_REQ14 & ~n7896;
  assign n7898 = ~n7895 & ~n7897;
  assign n7899 = ~controllable_BtoS_ACK14 & ~n7898;
  assign n7900 = ~n7892 & ~n7899;
  assign n7901 = controllable_ENQ & ~n7900;
  assign n7902 = controllable_ENQ & ~n7901;
  assign n7903 = ~i_RtoB_ACK1 & ~n7902;
  assign n7904 = ~n7886 & ~n7903;
  assign n7905 = controllable_BtoR_REQ1 & ~n7904;
  assign n7906 = ~n7071 & ~n7172;
  assign n7907 = ~i_StoB_REQ14 & ~n7906;
  assign n7908 = ~n7690 & ~n7907;
  assign n7909 = controllable_BtoS_ACK14 & ~n7908;
  assign n7910 = ~n5312 & ~n7224;
  assign n7911 = ~i_StoB_REQ14 & ~n7910;
  assign n7912 = ~n7895 & ~n7911;
  assign n7913 = ~controllable_BtoS_ACK14 & ~n7912;
  assign n7914 = ~n7909 & ~n7913;
  assign n7915 = controllable_ENQ & ~n7914;
  assign n7916 = controllable_ENQ & ~n7915;
  assign n7917 = ~controllable_BtoR_REQ1 & ~n7916;
  assign n7918 = ~n7905 & ~n7917;
  assign n7919 = ~controllable_BtoR_REQ0 & ~n7918;
  assign n7920 = ~controllable_BtoR_REQ0 & ~n7919;
  assign n7921 = i_RtoB_ACK0 & ~n7920;
  assign n7922 = ~i_StoB_REQ0 & ~n7250;
  assign n7923 = ~n5312 & ~n7922;
  assign n7924 = ~controllable_BtoS_ACK14 & ~n7923;
  assign n7925 = ~n7909 & ~n7924;
  assign n7926 = controllable_ENQ & ~n7925;
  assign n7927 = ~controllable_ENQ & ~n7883;
  assign n7928 = ~n7926 & ~n7927;
  assign n7929 = i_RtoB_ACK1 & ~n7928;
  assign n7930 = ~controllable_ENQ & ~n7900;
  assign n7931 = ~n7926 & ~n7930;
  assign n7932 = ~i_RtoB_ACK1 & ~n7931;
  assign n7933 = ~n7929 & ~n7932;
  assign n7934 = controllable_BtoR_REQ1 & ~n7933;
  assign n7935 = i_RtoB_ACK1 & ~n7916;
  assign n7936 = ~controllable_ENQ & ~n7914;
  assign n7937 = ~n7926 & ~n7936;
  assign n7938 = ~i_RtoB_ACK1 & ~n7937;
  assign n7939 = ~n7935 & ~n7938;
  assign n7940 = ~controllable_BtoR_REQ1 & ~n7939;
  assign n7941 = ~n7934 & ~n7940;
  assign n7942 = ~controllable_BtoR_REQ0 & ~n7941;
  assign n7943 = ~controllable_BtoR_REQ0 & ~n7942;
  assign n7944 = ~i_RtoB_ACK0 & ~n7943;
  assign n7945 = ~n7921 & ~n7944;
  assign n7946 = controllable_DEQ & ~n7945;
  assign n7947 = i_RtoB_ACK1 & ~n7883;
  assign n7948 = ~i_RtoB_ACK1 & ~n7900;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = controllable_BtoR_REQ1 & ~n7949;
  assign n7951 = ~controllable_BtoR_REQ1 & ~n7914;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~controllable_BtoR_REQ0 & ~n7952;
  assign n7954 = ~controllable_BtoR_REQ0 & ~n7953;
  assign n7955 = i_RtoB_ACK0 & ~n7954;
  assign n7956 = controllable_BtoR_REQ1 & ~n7925;
  assign n7957 = i_RtoB_ACK1 & ~n7914;
  assign n7958 = ~i_RtoB_ACK1 & ~n7925;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = ~controllable_BtoR_REQ1 & ~n7959;
  assign n7961 = ~n7956 & ~n7960;
  assign n7962 = ~controllable_BtoR_REQ0 & ~n7961;
  assign n7963 = ~controllable_BtoR_REQ0 & ~n7962;
  assign n7964 = ~i_RtoB_ACK0 & ~n7963;
  assign n7965 = ~n7955 & ~n7964;
  assign n7966 = ~controllable_DEQ & ~n7965;
  assign n7967 = ~n7946 & ~n7966;
  assign n7968 = i_FULL & ~n7967;
  assign n7969 = ~n7915 & ~n7927;
  assign n7970 = i_RtoB_ACK1 & ~n7969;
  assign n7971 = ~n7915 & ~n7930;
  assign n7972 = ~i_RtoB_ACK1 & ~n7971;
  assign n7973 = ~n7970 & ~n7972;
  assign n7974 = controllable_BtoR_REQ1 & ~n7973;
  assign n7975 = ~i_RtoB_ACK1 & ~n7914;
  assign n7976 = ~n7935 & ~n7975;
  assign n7977 = ~controllable_BtoR_REQ1 & ~n7976;
  assign n7978 = ~n7974 & ~n7977;
  assign n7979 = ~controllable_BtoR_REQ0 & ~n7978;
  assign n7980 = ~controllable_BtoR_REQ0 & ~n7979;
  assign n7981 = ~i_RtoB_ACK0 & ~n7980;
  assign n7982 = ~n7921 & ~n7981;
  assign n7983 = controllable_DEQ & ~n7982;
  assign n7984 = controllable_BtoR_REQ1 & ~n7937;
  assign n7985 = ~n7938 & ~n7957;
  assign n7986 = ~controllable_BtoR_REQ1 & ~n7985;
  assign n7987 = ~n7984 & ~n7986;
  assign n7988 = ~controllable_BtoR_REQ0 & ~n7987;
  assign n7989 = ~controllable_BtoR_REQ0 & ~n7988;
  assign n7990 = ~i_RtoB_ACK0 & ~n7989;
  assign n7991 = ~n7955 & ~n7990;
  assign n7992 = ~controllable_DEQ & ~n7991;
  assign n7993 = ~n7983 & ~n7992;
  assign n7994 = ~i_FULL & ~n7993;
  assign n7995 = ~n7968 & ~n7994;
  assign n7996 = i_nEMPTY & ~n7995;
  assign n7997 = ~controllable_ENQ & ~n7927;
  assign n7998 = i_RtoB_ACK1 & ~n7997;
  assign n7999 = ~controllable_ENQ & ~n7930;
  assign n8000 = ~i_RtoB_ACK1 & ~n7999;
  assign n8001 = ~n7998 & ~n8000;
  assign n8002 = controllable_BtoR_REQ1 & ~n8001;
  assign n8003 = ~controllable_ENQ & ~n7936;
  assign n8004 = ~i_RtoB_ACK1 & ~n8003;
  assign n8005 = ~i_RtoB_ACK1 & ~n8004;
  assign n8006 = ~controllable_BtoR_REQ1 & ~n8005;
  assign n8007 = ~n8002 & ~n8006;
  assign n8008 = ~controllable_BtoR_REQ0 & ~n8007;
  assign n8009 = ~controllable_BtoR_REQ0 & ~n8008;
  assign n8010 = ~i_RtoB_ACK0 & ~n8009;
  assign n8011 = ~i_RtoB_ACK0 & ~n8010;
  assign n8012 = controllable_DEQ & ~n8011;
  assign n8013 = controllable_ENQ & ~n7926;
  assign n8014 = controllable_BtoR_REQ1 & ~n8013;
  assign n8015 = ~i_RtoB_ACK1 & ~n8013;
  assign n8016 = ~n7935 & ~n8015;
  assign n8017 = ~controllable_BtoR_REQ1 & ~n8016;
  assign n8018 = ~n8014 & ~n8017;
  assign n8019 = ~controllable_BtoR_REQ0 & ~n8018;
  assign n8020 = ~controllable_BtoR_REQ0 & ~n8019;
  assign n8021 = ~i_RtoB_ACK0 & ~n8020;
  assign n8022 = ~n7921 & ~n8021;
  assign n8023 = ~controllable_DEQ & ~n8022;
  assign n8024 = ~n8012 & ~n8023;
  assign n8025 = i_FULL & ~n8024;
  assign n8026 = ~i_RtoB_ACK1 & ~n7975;
  assign n8027 = ~controllable_BtoR_REQ1 & ~n8026;
  assign n8028 = ~n7950 & ~n8027;
  assign n8029 = ~controllable_BtoR_REQ0 & ~n8028;
  assign n8030 = ~controllable_BtoR_REQ0 & ~n8029;
  assign n8031 = ~i_RtoB_ACK0 & ~n8030;
  assign n8032 = ~i_RtoB_ACK0 & ~n8031;
  assign n8033 = controllable_DEQ & ~n8032;
  assign n8034 = ~n7932 & ~n7935;
  assign n8035 = ~controllable_BtoR_REQ1 & ~n8034;
  assign n8036 = ~n7934 & ~n8035;
  assign n8037 = ~controllable_BtoR_REQ0 & ~n8036;
  assign n8038 = ~controllable_BtoR_REQ0 & ~n8037;
  assign n8039 = ~i_RtoB_ACK0 & ~n8038;
  assign n8040 = ~n7921 & ~n8039;
  assign n8041 = ~controllable_DEQ & ~n8040;
  assign n8042 = ~n8033 & ~n8041;
  assign n8043 = ~i_FULL & ~n8042;
  assign n8044 = ~n8025 & ~n8043;
  assign n8045 = ~i_nEMPTY & ~n8044;
  assign n8046 = ~n7996 & ~n8045;
  assign n8047 = controllable_BtoS_ACK0 & ~n8046;
  assign n8048 = i_StoB_REQ14 & ~n5213;
  assign n8049 = i_StoB_REQ0 & ~n7187;
  assign n8050 = ~n7179 & ~n8049;
  assign n8051 = ~i_StoB_REQ14 & ~n8050;
  assign n8052 = ~n8048 & ~n8051;
  assign n8053 = ~controllable_BtoS_ACK14 & ~n8052;
  assign n8054 = ~n7784 & ~n8053;
  assign n8055 = controllable_ENQ & ~n8054;
  assign n8056 = controllable_ENQ & ~n8055;
  assign n8057 = i_RtoB_ACK1 & ~n8056;
  assign n8058 = i_StoB_REQ0 & ~n7070;
  assign n8059 = ~n7062 & ~n8058;
  assign n8060 = ~i_StoB_REQ14 & ~n8059;
  assign n8061 = ~n7197 & ~n8060;
  assign n8062 = controllable_BtoS_ACK14 & ~n8061;
  assign n8063 = i_StoB_REQ14 & ~n7205;
  assign n8064 = i_StoB_REQ0 & ~n7223;
  assign n8065 = ~n7213 & ~n8064;
  assign n8066 = ~i_StoB_REQ14 & ~n8065;
  assign n8067 = ~n8063 & ~n8066;
  assign n8068 = ~controllable_BtoS_ACK14 & ~n8067;
  assign n8069 = ~n8062 & ~n8068;
  assign n8070 = controllable_ENQ & ~n8069;
  assign n8071 = controllable_ENQ & ~n8070;
  assign n8072 = ~i_RtoB_ACK1 & ~n8071;
  assign n8073 = ~n8057 & ~n8072;
  assign n8074 = controllable_BtoR_REQ1 & ~n8073;
  assign n8075 = ~i_StoB_REQ14 & ~n7070;
  assign n8076 = ~n5322 & ~n8075;
  assign n8077 = controllable_BtoS_ACK14 & ~n8076;
  assign n8078 = ~i_StoB_REQ14 & ~n7223;
  assign n8079 = ~n8063 & ~n8078;
  assign n8080 = ~controllable_BtoS_ACK14 & ~n8079;
  assign n8081 = ~n8077 & ~n8080;
  assign n8082 = controllable_ENQ & ~n8081;
  assign n8083 = controllable_ENQ & ~n8082;
  assign n8084 = ~controllable_BtoR_REQ1 & ~n8083;
  assign n8085 = ~n8074 & ~n8084;
  assign n8086 = ~controllable_BtoR_REQ0 & ~n8085;
  assign n8087 = ~controllable_BtoR_REQ0 & ~n8086;
  assign n8088 = i_RtoB_ACK0 & ~n8087;
  assign n8089 = ~n7254 & ~n8077;
  assign n8090 = controllable_ENQ & ~n8089;
  assign n8091 = ~controllable_ENQ & ~n8054;
  assign n8092 = ~n8090 & ~n8091;
  assign n8093 = i_RtoB_ACK1 & ~n8092;
  assign n8094 = ~controllable_ENQ & ~n8069;
  assign n8095 = ~n8090 & ~n8094;
  assign n8096 = ~i_RtoB_ACK1 & ~n8095;
  assign n8097 = ~n8093 & ~n8096;
  assign n8098 = controllable_BtoR_REQ1 & ~n8097;
  assign n8099 = i_RtoB_ACK1 & ~n8083;
  assign n8100 = ~controllable_ENQ & ~n8081;
  assign n8101 = ~n8090 & ~n8100;
  assign n8102 = ~i_RtoB_ACK1 & ~n8101;
  assign n8103 = ~n8099 & ~n8102;
  assign n8104 = ~controllable_BtoR_REQ1 & ~n8103;
  assign n8105 = ~n8098 & ~n8104;
  assign n8106 = ~controllable_BtoR_REQ0 & ~n8105;
  assign n8107 = ~controllable_BtoR_REQ0 & ~n8106;
  assign n8108 = ~i_RtoB_ACK0 & ~n8107;
  assign n8109 = ~n8088 & ~n8108;
  assign n8110 = controllable_DEQ & ~n8109;
  assign n8111 = i_RtoB_ACK1 & ~n8054;
  assign n8112 = ~i_RtoB_ACK1 & ~n8069;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = controllable_BtoR_REQ1 & ~n8113;
  assign n8115 = ~controllable_BtoR_REQ1 & ~n8081;
  assign n8116 = ~n8114 & ~n8115;
  assign n8117 = ~controllable_BtoR_REQ0 & ~n8116;
  assign n8118 = ~controllable_BtoR_REQ0 & ~n8117;
  assign n8119 = i_RtoB_ACK0 & ~n8118;
  assign n8120 = controllable_BtoR_REQ1 & ~n8089;
  assign n8121 = i_RtoB_ACK1 & ~n8081;
  assign n8122 = ~i_RtoB_ACK1 & ~n8089;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = ~controllable_BtoR_REQ1 & ~n8123;
  assign n8125 = ~n8120 & ~n8124;
  assign n8126 = ~controllable_BtoR_REQ0 & ~n8125;
  assign n8127 = ~controllable_BtoR_REQ0 & ~n8126;
  assign n8128 = ~i_RtoB_ACK0 & ~n8127;
  assign n8129 = ~n8119 & ~n8128;
  assign n8130 = ~controllable_DEQ & ~n8129;
  assign n8131 = ~n8110 & ~n8130;
  assign n8132 = i_FULL & ~n8131;
  assign n8133 = ~n8082 & ~n8091;
  assign n8134 = i_RtoB_ACK1 & ~n8133;
  assign n8135 = ~n8082 & ~n8094;
  assign n8136 = ~i_RtoB_ACK1 & ~n8135;
  assign n8137 = ~n8134 & ~n8136;
  assign n8138 = controllable_BtoR_REQ1 & ~n8137;
  assign n8139 = ~i_RtoB_ACK1 & ~n8081;
  assign n8140 = ~n8099 & ~n8139;
  assign n8141 = ~controllable_BtoR_REQ1 & ~n8140;
  assign n8142 = ~n8138 & ~n8141;
  assign n8143 = ~controllable_BtoR_REQ0 & ~n8142;
  assign n8144 = ~controllable_BtoR_REQ0 & ~n8143;
  assign n8145 = ~i_RtoB_ACK0 & ~n8144;
  assign n8146 = ~n8088 & ~n8145;
  assign n8147 = controllable_DEQ & ~n8146;
  assign n8148 = controllable_BtoR_REQ1 & ~n8101;
  assign n8149 = ~n8102 & ~n8121;
  assign n8150 = ~controllable_BtoR_REQ1 & ~n8149;
  assign n8151 = ~n8148 & ~n8150;
  assign n8152 = ~controllable_BtoR_REQ0 & ~n8151;
  assign n8153 = ~controllable_BtoR_REQ0 & ~n8152;
  assign n8154 = ~i_RtoB_ACK0 & ~n8153;
  assign n8155 = ~n8119 & ~n8154;
  assign n8156 = ~controllable_DEQ & ~n8155;
  assign n8157 = ~n8147 & ~n8156;
  assign n8158 = ~i_FULL & ~n8157;
  assign n8159 = ~n8132 & ~n8158;
  assign n8160 = i_nEMPTY & ~n8159;
  assign n8161 = ~controllable_ENQ & ~n8091;
  assign n8162 = i_RtoB_ACK1 & ~n8161;
  assign n8163 = ~controllable_ENQ & ~n8094;
  assign n8164 = ~i_RtoB_ACK1 & ~n8163;
  assign n8165 = ~n8162 & ~n8164;
  assign n8166 = controllable_BtoR_REQ1 & ~n8165;
  assign n8167 = ~controllable_ENQ & ~n8100;
  assign n8168 = ~i_RtoB_ACK1 & ~n8167;
  assign n8169 = ~i_RtoB_ACK1 & ~n8168;
  assign n8170 = ~controllable_BtoR_REQ1 & ~n8169;
  assign n8171 = ~n8166 & ~n8170;
  assign n8172 = ~controllable_BtoR_REQ0 & ~n8171;
  assign n8173 = ~controllable_BtoR_REQ0 & ~n8172;
  assign n8174 = ~i_RtoB_ACK0 & ~n8173;
  assign n8175 = ~i_RtoB_ACK0 & ~n8174;
  assign n8176 = controllable_DEQ & ~n8175;
  assign n8177 = controllable_ENQ & ~n8090;
  assign n8178 = controllable_BtoR_REQ1 & ~n8177;
  assign n8179 = ~i_RtoB_ACK1 & ~n8177;
  assign n8180 = ~n8099 & ~n8179;
  assign n8181 = ~controllable_BtoR_REQ1 & ~n8180;
  assign n8182 = ~n8178 & ~n8181;
  assign n8183 = ~controllable_BtoR_REQ0 & ~n8182;
  assign n8184 = ~controllable_BtoR_REQ0 & ~n8183;
  assign n8185 = ~i_RtoB_ACK0 & ~n8184;
  assign n8186 = ~n8088 & ~n8185;
  assign n8187 = ~controllable_DEQ & ~n8186;
  assign n8188 = ~n8176 & ~n8187;
  assign n8189 = i_FULL & ~n8188;
  assign n8190 = ~i_RtoB_ACK1 & ~n8139;
  assign n8191 = ~controllable_BtoR_REQ1 & ~n8190;
  assign n8192 = ~n8114 & ~n8191;
  assign n8193 = ~controllable_BtoR_REQ0 & ~n8192;
  assign n8194 = ~controllable_BtoR_REQ0 & ~n8193;
  assign n8195 = ~i_RtoB_ACK0 & ~n8194;
  assign n8196 = ~i_RtoB_ACK0 & ~n8195;
  assign n8197 = controllable_DEQ & ~n8196;
  assign n8198 = ~n8096 & ~n8099;
  assign n8199 = ~controllable_BtoR_REQ1 & ~n8198;
  assign n8200 = ~n8098 & ~n8199;
  assign n8201 = ~controllable_BtoR_REQ0 & ~n8200;
  assign n8202 = ~controllable_BtoR_REQ0 & ~n8201;
  assign n8203 = ~i_RtoB_ACK0 & ~n8202;
  assign n8204 = ~n8088 & ~n8203;
  assign n8205 = ~controllable_DEQ & ~n8204;
  assign n8206 = ~n8197 & ~n8205;
  assign n8207 = ~i_FULL & ~n8206;
  assign n8208 = ~n8189 & ~n8207;
  assign n8209 = ~i_nEMPTY & ~n8208;
  assign n8210 = ~n8160 & ~n8209;
  assign n8211 = ~controllable_BtoS_ACK0 & ~n8210;
  assign n8212 = ~n8047 & ~n8211;
  assign n8213 = n4465 & ~n8212;
  assign n8214 = ~n7055 & ~n7890;
  assign n8215 = controllable_BtoS_ACK14 & ~n8214;
  assign n8216 = ~n7075 & ~n8215;
  assign n8217 = controllable_ENQ & ~n8216;
  assign n8218 = controllable_ENQ & ~n8217;
  assign n8219 = ~i_RtoB_ACK1 & ~n8218;
  assign n8220 = ~n7054 & ~n8219;
  assign n8221 = controllable_BtoR_REQ1 & ~n8220;
  assign n8222 = ~n5216 & ~n7907;
  assign n8223 = controllable_BtoS_ACK14 & ~n8222;
  assign n8224 = ~n7085 & ~n8223;
  assign n8225 = controllable_ENQ & ~n8224;
  assign n8226 = controllable_ENQ & ~n8225;
  assign n8227 = ~controllable_BtoR_REQ1 & ~n8226;
  assign n8228 = ~n8221 & ~n8227;
  assign n8229 = ~controllable_BtoR_REQ0 & ~n8228;
  assign n8230 = ~controllable_BtoR_REQ0 & ~n8229;
  assign n8231 = i_RtoB_ACK0 & ~n8230;
  assign n8232 = ~n5238 & ~n8225;
  assign n8233 = i_RtoB_ACK1 & ~n8232;
  assign n8234 = ~controllable_ENQ & ~n8216;
  assign n8235 = ~n8225 & ~n8234;
  assign n8236 = ~i_RtoB_ACK1 & ~n8235;
  assign n8237 = ~n8233 & ~n8236;
  assign n8238 = controllable_BtoR_REQ1 & ~n8237;
  assign n8239 = i_RtoB_ACK1 & ~n8226;
  assign n8240 = ~i_RtoB_ACK1 & ~n8224;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~controllable_BtoR_REQ1 & ~n8241;
  assign n8243 = ~n8238 & ~n8242;
  assign n8244 = ~controllable_BtoR_REQ0 & ~n8243;
  assign n8245 = ~controllable_BtoR_REQ0 & ~n8244;
  assign n8246 = ~i_RtoB_ACK0 & ~n8245;
  assign n8247 = ~n8231 & ~n8246;
  assign n8248 = controllable_DEQ & ~n8247;
  assign n8249 = ~i_RtoB_ACK1 & ~n8216;
  assign n8250 = ~n7111 & ~n8249;
  assign n8251 = controllable_BtoR_REQ1 & ~n8250;
  assign n8252 = ~controllable_BtoR_REQ1 & ~n8224;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = ~controllable_BtoR_REQ0 & ~n8253;
  assign n8255 = ~controllable_BtoR_REQ0 & ~n8254;
  assign n8256 = i_RtoB_ACK0 & ~n8255;
  assign n8257 = ~controllable_BtoR_REQ0 & ~n8224;
  assign n8258 = ~controllable_BtoR_REQ0 & ~n8257;
  assign n8259 = ~i_RtoB_ACK0 & ~n8258;
  assign n8260 = ~n8256 & ~n8259;
  assign n8261 = ~controllable_DEQ & ~n8260;
  assign n8262 = ~n8248 & ~n8261;
  assign n8263 = i_nEMPTY & ~n8262;
  assign n8264 = ~controllable_ENQ & ~n8234;
  assign n8265 = ~i_RtoB_ACK1 & ~n8264;
  assign n8266 = ~n7127 & ~n8265;
  assign n8267 = controllable_BtoR_REQ1 & ~n8266;
  assign n8268 = ~controllable_ENQ & ~n8224;
  assign n8269 = ~controllable_ENQ & ~n8268;
  assign n8270 = ~i_RtoB_ACK1 & ~n8269;
  assign n8271 = ~i_RtoB_ACK1 & ~n8270;
  assign n8272 = ~controllable_BtoR_REQ1 & ~n8271;
  assign n8273 = ~n8267 & ~n8272;
  assign n8274 = ~controllable_BtoR_REQ0 & ~n8273;
  assign n8275 = ~controllable_BtoR_REQ0 & ~n8274;
  assign n8276 = ~i_RtoB_ACK0 & ~n8275;
  assign n8277 = ~i_RtoB_ACK0 & ~n8276;
  assign n8278 = controllable_DEQ & ~n8277;
  assign n8279 = ~controllable_BtoR_REQ0 & ~n8226;
  assign n8280 = ~controllable_BtoR_REQ0 & ~n8279;
  assign n8281 = ~i_RtoB_ACK0 & ~n8280;
  assign n8282 = ~n8231 & ~n8281;
  assign n8283 = ~controllable_DEQ & ~n8282;
  assign n8284 = ~n8278 & ~n8283;
  assign n8285 = i_FULL & ~n8284;
  assign n8286 = ~i_RtoB_ACK1 & ~n8240;
  assign n8287 = ~controllable_BtoR_REQ1 & ~n8286;
  assign n8288 = ~n8251 & ~n8287;
  assign n8289 = ~controllable_BtoR_REQ0 & ~n8288;
  assign n8290 = ~controllable_BtoR_REQ0 & ~n8289;
  assign n8291 = ~i_RtoB_ACK0 & ~n8290;
  assign n8292 = ~i_RtoB_ACK0 & ~n8291;
  assign n8293 = controllable_DEQ & ~n8292;
  assign n8294 = ~n8236 & ~n8239;
  assign n8295 = ~controllable_BtoR_REQ1 & ~n8294;
  assign n8296 = ~n8238 & ~n8295;
  assign n8297 = ~controllable_BtoR_REQ0 & ~n8296;
  assign n8298 = ~controllable_BtoR_REQ0 & ~n8297;
  assign n8299 = ~i_RtoB_ACK0 & ~n8298;
  assign n8300 = ~n8231 & ~n8299;
  assign n8301 = ~controllable_DEQ & ~n8300;
  assign n8302 = ~n8293 & ~n8301;
  assign n8303 = ~i_FULL & ~n8302;
  assign n8304 = ~n8285 & ~n8303;
  assign n8305 = ~i_nEMPTY & ~n8304;
  assign n8306 = ~n8263 & ~n8305;
  assign n8307 = controllable_BtoS_ACK0 & ~n8306;
  assign n8308 = ~n7181 & ~n8048;
  assign n8309 = ~controllable_BtoS_ACK14 & ~n8308;
  assign n8310 = ~n7784 & ~n8309;
  assign n8311 = controllable_ENQ & ~n8310;
  assign n8312 = controllable_ENQ & ~n8311;
  assign n8313 = i_RtoB_ACK1 & ~n8312;
  assign n8314 = ~n7215 & ~n8063;
  assign n8315 = ~controllable_BtoS_ACK14 & ~n8314;
  assign n8316 = ~n8062 & ~n8315;
  assign n8317 = controllable_ENQ & ~n8316;
  assign n8318 = controllable_ENQ & ~n8317;
  assign n8319 = ~i_RtoB_ACK1 & ~n8318;
  assign n8320 = ~n8313 & ~n8319;
  assign n8321 = controllable_BtoR_REQ1 & ~n8320;
  assign n8322 = ~n7235 & ~n8063;
  assign n8323 = ~controllable_BtoS_ACK14 & ~n8322;
  assign n8324 = ~n8077 & ~n8323;
  assign n8325 = controllable_ENQ & ~n8324;
  assign n8326 = controllable_ENQ & ~n8325;
  assign n8327 = ~controllable_BtoR_REQ1 & ~n8326;
  assign n8328 = ~n8321 & ~n8327;
  assign n8329 = ~controllable_BtoR_REQ0 & ~n8328;
  assign n8330 = ~controllable_BtoR_REQ0 & ~n8329;
  assign n8331 = i_RtoB_ACK0 & ~n8330;
  assign n8332 = ~controllable_ENQ & ~n8310;
  assign n8333 = ~n8090 & ~n8332;
  assign n8334 = i_RtoB_ACK1 & ~n8333;
  assign n8335 = ~controllable_ENQ & ~n8316;
  assign n8336 = ~n8090 & ~n8335;
  assign n8337 = ~i_RtoB_ACK1 & ~n8336;
  assign n8338 = ~n8334 & ~n8337;
  assign n8339 = controllable_BtoR_REQ1 & ~n8338;
  assign n8340 = i_RtoB_ACK1 & ~n8326;
  assign n8341 = ~controllable_ENQ & ~n8324;
  assign n8342 = ~n8090 & ~n8341;
  assign n8343 = ~i_RtoB_ACK1 & ~n8342;
  assign n8344 = ~n8340 & ~n8343;
  assign n8345 = ~controllable_BtoR_REQ1 & ~n8344;
  assign n8346 = ~n8339 & ~n8345;
  assign n8347 = ~controllable_BtoR_REQ0 & ~n8346;
  assign n8348 = ~controllable_BtoR_REQ0 & ~n8347;
  assign n8349 = ~i_RtoB_ACK0 & ~n8348;
  assign n8350 = ~n8331 & ~n8349;
  assign n8351 = controllable_DEQ & ~n8350;
  assign n8352 = i_RtoB_ACK1 & ~n8310;
  assign n8353 = ~i_RtoB_ACK1 & ~n8316;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = controllable_BtoR_REQ1 & ~n8354;
  assign n8356 = ~controllable_BtoR_REQ1 & ~n8324;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~controllable_BtoR_REQ0 & ~n8357;
  assign n8359 = ~controllable_BtoR_REQ0 & ~n8358;
  assign n8360 = i_RtoB_ACK0 & ~n8359;
  assign n8361 = i_RtoB_ACK1 & ~n8324;
  assign n8362 = ~n8122 & ~n8361;
  assign n8363 = ~controllable_BtoR_REQ1 & ~n8362;
  assign n8364 = ~n8120 & ~n8363;
  assign n8365 = ~controllable_BtoR_REQ0 & ~n8364;
  assign n8366 = ~controllable_BtoR_REQ0 & ~n8365;
  assign n8367 = ~i_RtoB_ACK0 & ~n8366;
  assign n8368 = ~n8360 & ~n8367;
  assign n8369 = ~controllable_DEQ & ~n8368;
  assign n8370 = ~n8351 & ~n8369;
  assign n8371 = i_FULL & ~n8370;
  assign n8372 = ~n8325 & ~n8332;
  assign n8373 = i_RtoB_ACK1 & ~n8372;
  assign n8374 = ~n8325 & ~n8335;
  assign n8375 = ~i_RtoB_ACK1 & ~n8374;
  assign n8376 = ~n8373 & ~n8375;
  assign n8377 = controllable_BtoR_REQ1 & ~n8376;
  assign n8378 = ~i_RtoB_ACK1 & ~n8324;
  assign n8379 = ~n8340 & ~n8378;
  assign n8380 = ~controllable_BtoR_REQ1 & ~n8379;
  assign n8381 = ~n8377 & ~n8380;
  assign n8382 = ~controllable_BtoR_REQ0 & ~n8381;
  assign n8383 = ~controllable_BtoR_REQ0 & ~n8382;
  assign n8384 = ~i_RtoB_ACK0 & ~n8383;
  assign n8385 = ~n8331 & ~n8384;
  assign n8386 = controllable_DEQ & ~n8385;
  assign n8387 = controllable_BtoR_REQ1 & ~n8342;
  assign n8388 = ~n8343 & ~n8361;
  assign n8389 = ~controllable_BtoR_REQ1 & ~n8388;
  assign n8390 = ~n8387 & ~n8389;
  assign n8391 = ~controllable_BtoR_REQ0 & ~n8390;
  assign n8392 = ~controllable_BtoR_REQ0 & ~n8391;
  assign n8393 = ~i_RtoB_ACK0 & ~n8392;
  assign n8394 = ~n8360 & ~n8393;
  assign n8395 = ~controllable_DEQ & ~n8394;
  assign n8396 = ~n8386 & ~n8395;
  assign n8397 = ~i_FULL & ~n8396;
  assign n8398 = ~n8371 & ~n8397;
  assign n8399 = i_nEMPTY & ~n8398;
  assign n8400 = ~controllable_ENQ & ~n8332;
  assign n8401 = i_RtoB_ACK1 & ~n8400;
  assign n8402 = ~controllable_ENQ & ~n8335;
  assign n8403 = ~i_RtoB_ACK1 & ~n8402;
  assign n8404 = ~n8401 & ~n8403;
  assign n8405 = controllable_BtoR_REQ1 & ~n8404;
  assign n8406 = ~controllable_ENQ & ~n8341;
  assign n8407 = ~i_RtoB_ACK1 & ~n8406;
  assign n8408 = ~i_RtoB_ACK1 & ~n8407;
  assign n8409 = ~controllable_BtoR_REQ1 & ~n8408;
  assign n8410 = ~n8405 & ~n8409;
  assign n8411 = ~controllable_BtoR_REQ0 & ~n8410;
  assign n8412 = ~controllable_BtoR_REQ0 & ~n8411;
  assign n8413 = ~i_RtoB_ACK0 & ~n8412;
  assign n8414 = ~i_RtoB_ACK0 & ~n8413;
  assign n8415 = controllable_DEQ & ~n8414;
  assign n8416 = ~n8179 & ~n8340;
  assign n8417 = ~controllable_BtoR_REQ1 & ~n8416;
  assign n8418 = ~n8178 & ~n8417;
  assign n8419 = ~controllable_BtoR_REQ0 & ~n8418;
  assign n8420 = ~controllable_BtoR_REQ0 & ~n8419;
  assign n8421 = ~i_RtoB_ACK0 & ~n8420;
  assign n8422 = ~n8331 & ~n8421;
  assign n8423 = ~controllable_DEQ & ~n8422;
  assign n8424 = ~n8415 & ~n8423;
  assign n8425 = i_FULL & ~n8424;
  assign n8426 = ~i_RtoB_ACK1 & ~n8378;
  assign n8427 = ~controllable_BtoR_REQ1 & ~n8426;
  assign n8428 = ~n8355 & ~n8427;
  assign n8429 = ~controllable_BtoR_REQ0 & ~n8428;
  assign n8430 = ~controllable_BtoR_REQ0 & ~n8429;
  assign n8431 = ~i_RtoB_ACK0 & ~n8430;
  assign n8432 = ~i_RtoB_ACK0 & ~n8431;
  assign n8433 = controllable_DEQ & ~n8432;
  assign n8434 = ~n8337 & ~n8340;
  assign n8435 = ~controllable_BtoR_REQ1 & ~n8434;
  assign n8436 = ~n8339 & ~n8435;
  assign n8437 = ~controllable_BtoR_REQ0 & ~n8436;
  assign n8438 = ~controllable_BtoR_REQ0 & ~n8437;
  assign n8439 = ~i_RtoB_ACK0 & ~n8438;
  assign n8440 = ~n8331 & ~n8439;
  assign n8441 = ~controllable_DEQ & ~n8440;
  assign n8442 = ~n8433 & ~n8441;
  assign n8443 = ~i_FULL & ~n8442;
  assign n8444 = ~n8425 & ~n8443;
  assign n8445 = ~i_nEMPTY & ~n8444;
  assign n8446 = ~n8399 & ~n8445;
  assign n8447 = ~controllable_BtoS_ACK0 & ~n8446;
  assign n8448 = ~n8307 & ~n8447;
  assign n8449 = ~n4465 & ~n8448;
  assign n8450 = ~n8213 & ~n8449;
  assign n8451 = ~i_StoB_REQ10 & ~n8450;
  assign n8452 = ~n7878 & ~n8451;
  assign n8453 = controllable_BtoS_ACK10 & ~n8452;
  assign n8454 = ~i_StoB_REQ0 & ~n7188;
  assign n8455 = ~i_StoB_REQ14 & ~n8454;
  assign n8456 = ~n5216 & ~n8455;
  assign n8457 = ~controllable_BtoS_ACK14 & ~n8456;
  assign n8458 = ~n5227 & ~n8457;
  assign n8459 = controllable_ENQ & ~n8458;
  assign n8460 = controllable_ENQ & ~n8459;
  assign n8461 = i_RtoB_ACK1 & ~n8460;
  assign n8462 = ~i_RtoB_ACK1 & ~n7916;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = controllable_BtoR_REQ1 & ~n8463;
  assign n8465 = ~n7917 & ~n8464;
  assign n8466 = ~controllable_BtoR_REQ0 & ~n8465;
  assign n8467 = ~controllable_BtoR_REQ0 & ~n8466;
  assign n8468 = i_RtoB_ACK0 & ~n8467;
  assign n8469 = ~controllable_ENQ & ~n8458;
  assign n8470 = ~n7926 & ~n8469;
  assign n8471 = i_RtoB_ACK1 & ~n8470;
  assign n8472 = ~n7938 & ~n8471;
  assign n8473 = controllable_BtoR_REQ1 & ~n8472;
  assign n8474 = ~n7940 & ~n8473;
  assign n8475 = ~controllable_BtoR_REQ0 & ~n8474;
  assign n8476 = ~controllable_BtoR_REQ0 & ~n8475;
  assign n8477 = ~i_RtoB_ACK0 & ~n8476;
  assign n8478 = ~n8468 & ~n8477;
  assign n8479 = controllable_DEQ & ~n8478;
  assign n8480 = i_RtoB_ACK1 & ~n8458;
  assign n8481 = ~n7975 & ~n8480;
  assign n8482 = controllable_BtoR_REQ1 & ~n8481;
  assign n8483 = ~n7951 & ~n8482;
  assign n8484 = ~controllable_BtoR_REQ0 & ~n8483;
  assign n8485 = ~controllable_BtoR_REQ0 & ~n8484;
  assign n8486 = i_RtoB_ACK0 & ~n8485;
  assign n8487 = ~n7964 & ~n8486;
  assign n8488 = ~controllable_DEQ & ~n8487;
  assign n8489 = ~n8479 & ~n8488;
  assign n8490 = i_FULL & ~n8489;
  assign n8491 = ~n7915 & ~n8469;
  assign n8492 = i_RtoB_ACK1 & ~n8491;
  assign n8493 = ~n7975 & ~n8492;
  assign n8494 = controllable_BtoR_REQ1 & ~n8493;
  assign n8495 = ~n7977 & ~n8494;
  assign n8496 = ~controllable_BtoR_REQ0 & ~n8495;
  assign n8497 = ~controllable_BtoR_REQ0 & ~n8496;
  assign n8498 = ~i_RtoB_ACK0 & ~n8497;
  assign n8499 = ~n8468 & ~n8498;
  assign n8500 = controllable_DEQ & ~n8499;
  assign n8501 = ~n7990 & ~n8486;
  assign n8502 = ~controllable_DEQ & ~n8501;
  assign n8503 = ~n8500 & ~n8502;
  assign n8504 = ~i_FULL & ~n8503;
  assign n8505 = ~n8490 & ~n8504;
  assign n8506 = i_nEMPTY & ~n8505;
  assign n8507 = ~controllable_ENQ & ~n8469;
  assign n8508 = i_RtoB_ACK1 & ~n8507;
  assign n8509 = ~n8004 & ~n8508;
  assign n8510 = controllable_BtoR_REQ1 & ~n8509;
  assign n8511 = ~n8006 & ~n8510;
  assign n8512 = ~controllable_BtoR_REQ0 & ~n8511;
  assign n8513 = ~controllable_BtoR_REQ0 & ~n8512;
  assign n8514 = ~i_RtoB_ACK0 & ~n8513;
  assign n8515 = ~i_RtoB_ACK0 & ~n8514;
  assign n8516 = controllable_DEQ & ~n8515;
  assign n8517 = ~n8021 & ~n8468;
  assign n8518 = ~controllable_DEQ & ~n8517;
  assign n8519 = ~n8516 & ~n8518;
  assign n8520 = i_FULL & ~n8519;
  assign n8521 = ~n8027 & ~n8482;
  assign n8522 = ~controllable_BtoR_REQ0 & ~n8521;
  assign n8523 = ~controllable_BtoR_REQ0 & ~n8522;
  assign n8524 = ~i_RtoB_ACK0 & ~n8523;
  assign n8525 = ~i_RtoB_ACK0 & ~n8524;
  assign n8526 = controllable_DEQ & ~n8525;
  assign n8527 = ~controllable_DEQ & ~n8478;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = ~i_FULL & ~n8528;
  assign n8530 = ~n8520 & ~n8529;
  assign n8531 = ~i_nEMPTY & ~n8530;
  assign n8532 = ~n8506 & ~n8531;
  assign n8533 = controllable_BtoS_ACK0 & ~n8532;
  assign n8534 = ~i_StoB_REQ14 & ~n7187;
  assign n8535 = ~n8048 & ~n8534;
  assign n8536 = ~controllable_BtoS_ACK14 & ~n8535;
  assign n8537 = ~n7793 & ~n8536;
  assign n8538 = controllable_ENQ & ~n8537;
  assign n8539 = controllable_ENQ & ~n8538;
  assign n8540 = i_RtoB_ACK1 & ~n8539;
  assign n8541 = ~i_RtoB_ACK1 & ~n8083;
  assign n8542 = ~n8540 & ~n8541;
  assign n8543 = controllable_BtoR_REQ1 & ~n8542;
  assign n8544 = ~n8084 & ~n8543;
  assign n8545 = ~controllable_BtoR_REQ0 & ~n8544;
  assign n8546 = ~controllable_BtoR_REQ0 & ~n8545;
  assign n8547 = i_RtoB_ACK0 & ~n8546;
  assign n8548 = ~controllable_ENQ & ~n8537;
  assign n8549 = ~n8090 & ~n8548;
  assign n8550 = i_RtoB_ACK1 & ~n8549;
  assign n8551 = ~n8102 & ~n8550;
  assign n8552 = controllable_BtoR_REQ1 & ~n8551;
  assign n8553 = ~n8104 & ~n8552;
  assign n8554 = ~controllable_BtoR_REQ0 & ~n8553;
  assign n8555 = ~controllable_BtoR_REQ0 & ~n8554;
  assign n8556 = ~i_RtoB_ACK0 & ~n8555;
  assign n8557 = ~n8547 & ~n8556;
  assign n8558 = controllable_DEQ & ~n8557;
  assign n8559 = i_RtoB_ACK1 & ~n8537;
  assign n8560 = ~n8139 & ~n8559;
  assign n8561 = controllable_BtoR_REQ1 & ~n8560;
  assign n8562 = ~n8115 & ~n8561;
  assign n8563 = ~controllable_BtoR_REQ0 & ~n8562;
  assign n8564 = ~controllable_BtoR_REQ0 & ~n8563;
  assign n8565 = i_RtoB_ACK0 & ~n8564;
  assign n8566 = ~n8128 & ~n8565;
  assign n8567 = ~controllable_DEQ & ~n8566;
  assign n8568 = ~n8558 & ~n8567;
  assign n8569 = i_FULL & ~n8568;
  assign n8570 = ~n8082 & ~n8548;
  assign n8571 = i_RtoB_ACK1 & ~n8570;
  assign n8572 = ~n8139 & ~n8571;
  assign n8573 = controllable_BtoR_REQ1 & ~n8572;
  assign n8574 = ~n8141 & ~n8573;
  assign n8575 = ~controllable_BtoR_REQ0 & ~n8574;
  assign n8576 = ~controllable_BtoR_REQ0 & ~n8575;
  assign n8577 = ~i_RtoB_ACK0 & ~n8576;
  assign n8578 = ~n8547 & ~n8577;
  assign n8579 = controllable_DEQ & ~n8578;
  assign n8580 = ~n8154 & ~n8565;
  assign n8581 = ~controllable_DEQ & ~n8580;
  assign n8582 = ~n8579 & ~n8581;
  assign n8583 = ~i_FULL & ~n8582;
  assign n8584 = ~n8569 & ~n8583;
  assign n8585 = i_nEMPTY & ~n8584;
  assign n8586 = ~controllable_ENQ & ~n8548;
  assign n8587 = i_RtoB_ACK1 & ~n8586;
  assign n8588 = ~n8168 & ~n8587;
  assign n8589 = controllable_BtoR_REQ1 & ~n8588;
  assign n8590 = ~n8170 & ~n8589;
  assign n8591 = ~controllable_BtoR_REQ0 & ~n8590;
  assign n8592 = ~controllable_BtoR_REQ0 & ~n8591;
  assign n8593 = ~i_RtoB_ACK0 & ~n8592;
  assign n8594 = ~i_RtoB_ACK0 & ~n8593;
  assign n8595 = controllable_DEQ & ~n8594;
  assign n8596 = ~n8185 & ~n8547;
  assign n8597 = ~controllable_DEQ & ~n8596;
  assign n8598 = ~n8595 & ~n8597;
  assign n8599 = i_FULL & ~n8598;
  assign n8600 = ~n8191 & ~n8561;
  assign n8601 = ~controllable_BtoR_REQ0 & ~n8600;
  assign n8602 = ~controllable_BtoR_REQ0 & ~n8601;
  assign n8603 = ~i_RtoB_ACK0 & ~n8602;
  assign n8604 = ~i_RtoB_ACK0 & ~n8603;
  assign n8605 = controllable_DEQ & ~n8604;
  assign n8606 = ~controllable_DEQ & ~n8557;
  assign n8607 = ~n8605 & ~n8606;
  assign n8608 = ~i_FULL & ~n8607;
  assign n8609 = ~n8599 & ~n8608;
  assign n8610 = ~i_nEMPTY & ~n8609;
  assign n8611 = ~n8585 & ~n8610;
  assign n8612 = ~controllable_BtoS_ACK0 & ~n8611;
  assign n8613 = ~n8533 & ~n8612;
  assign n8614 = n4465 & ~n8613;
  assign n8615 = ~i_RtoB_ACK1 & ~n8226;
  assign n8616 = ~n5237 & ~n8615;
  assign n8617 = controllable_BtoR_REQ1 & ~n8616;
  assign n8618 = ~n8227 & ~n8617;
  assign n8619 = ~controllable_BtoR_REQ0 & ~n8618;
  assign n8620 = ~controllable_BtoR_REQ0 & ~n8619;
  assign n8621 = i_RtoB_ACK0 & ~n8620;
  assign n8622 = ~n5271 & ~n8225;
  assign n8623 = i_RtoB_ACK1 & ~n8622;
  assign n8624 = ~n8240 & ~n8623;
  assign n8625 = controllable_BtoR_REQ1 & ~n8624;
  assign n8626 = ~n8242 & ~n8625;
  assign n8627 = ~controllable_BtoR_REQ0 & ~n8626;
  assign n8628 = ~controllable_BtoR_REQ0 & ~n8627;
  assign n8629 = ~i_RtoB_ACK0 & ~n8628;
  assign n8630 = ~n8621 & ~n8629;
  assign n8631 = controllable_DEQ & ~n8630;
  assign n8632 = ~n7563 & ~n8240;
  assign n8633 = controllable_BtoR_REQ1 & ~n8632;
  assign n8634 = ~n8252 & ~n8633;
  assign n8635 = ~controllable_BtoR_REQ0 & ~n8634;
  assign n8636 = ~controllable_BtoR_REQ0 & ~n8635;
  assign n8637 = i_RtoB_ACK0 & ~n8636;
  assign n8638 = ~n8259 & ~n8637;
  assign n8639 = ~controllable_DEQ & ~n8638;
  assign n8640 = ~n8631 & ~n8639;
  assign n8641 = i_nEMPTY & ~n8640;
  assign n8642 = ~n7574 & ~n8270;
  assign n8643 = controllable_BtoR_REQ1 & ~n8642;
  assign n8644 = ~n8272 & ~n8643;
  assign n8645 = ~controllable_BtoR_REQ0 & ~n8644;
  assign n8646 = ~controllable_BtoR_REQ0 & ~n8645;
  assign n8647 = ~i_RtoB_ACK0 & ~n8646;
  assign n8648 = ~i_RtoB_ACK0 & ~n8647;
  assign n8649 = controllable_DEQ & ~n8648;
  assign n8650 = ~n8281 & ~n8621;
  assign n8651 = ~controllable_DEQ & ~n8650;
  assign n8652 = ~n8649 & ~n8651;
  assign n8653 = i_FULL & ~n8652;
  assign n8654 = ~n8287 & ~n8633;
  assign n8655 = ~controllable_BtoR_REQ0 & ~n8654;
  assign n8656 = ~controllable_BtoR_REQ0 & ~n8655;
  assign n8657 = ~i_RtoB_ACK0 & ~n8656;
  assign n8658 = ~i_RtoB_ACK0 & ~n8657;
  assign n8659 = controllable_DEQ & ~n8658;
  assign n8660 = ~controllable_DEQ & ~n8630;
  assign n8661 = ~n8659 & ~n8660;
  assign n8662 = ~i_FULL & ~n8661;
  assign n8663 = ~n8653 & ~n8662;
  assign n8664 = ~i_nEMPTY & ~n8663;
  assign n8665 = ~n8641 & ~n8664;
  assign n8666 = controllable_BtoS_ACK0 & ~n8665;
  assign n8667 = ~n7600 & ~n8048;
  assign n8668 = ~controllable_BtoS_ACK14 & ~n8667;
  assign n8669 = ~n7793 & ~n8668;
  assign n8670 = controllable_ENQ & ~n8669;
  assign n8671 = controllable_ENQ & ~n8670;
  assign n8672 = i_RtoB_ACK1 & ~n8671;
  assign n8673 = ~i_RtoB_ACK1 & ~n8326;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = controllable_BtoR_REQ1 & ~n8674;
  assign n8676 = ~n8327 & ~n8675;
  assign n8677 = ~controllable_BtoR_REQ0 & ~n8676;
  assign n8678 = ~controllable_BtoR_REQ0 & ~n8677;
  assign n8679 = i_RtoB_ACK0 & ~n8678;
  assign n8680 = ~controllable_ENQ & ~n8669;
  assign n8681 = ~n8090 & ~n8680;
  assign n8682 = i_RtoB_ACK1 & ~n8681;
  assign n8683 = ~n8343 & ~n8682;
  assign n8684 = controllable_BtoR_REQ1 & ~n8683;
  assign n8685 = ~n8345 & ~n8684;
  assign n8686 = ~controllable_BtoR_REQ0 & ~n8685;
  assign n8687 = ~controllable_BtoR_REQ0 & ~n8686;
  assign n8688 = ~i_RtoB_ACK0 & ~n8687;
  assign n8689 = ~n8679 & ~n8688;
  assign n8690 = controllable_DEQ & ~n8689;
  assign n8691 = i_RtoB_ACK1 & ~n8669;
  assign n8692 = ~n8378 & ~n8691;
  assign n8693 = controllable_BtoR_REQ1 & ~n8692;
  assign n8694 = ~n8356 & ~n8693;
  assign n8695 = ~controllable_BtoR_REQ0 & ~n8694;
  assign n8696 = ~controllable_BtoR_REQ0 & ~n8695;
  assign n8697 = i_RtoB_ACK0 & ~n8696;
  assign n8698 = ~n8367 & ~n8697;
  assign n8699 = ~controllable_DEQ & ~n8698;
  assign n8700 = ~n8690 & ~n8699;
  assign n8701 = i_FULL & ~n8700;
  assign n8702 = ~n8325 & ~n8680;
  assign n8703 = i_RtoB_ACK1 & ~n8702;
  assign n8704 = ~n8378 & ~n8703;
  assign n8705 = controllable_BtoR_REQ1 & ~n8704;
  assign n8706 = ~n8380 & ~n8705;
  assign n8707 = ~controllable_BtoR_REQ0 & ~n8706;
  assign n8708 = ~controllable_BtoR_REQ0 & ~n8707;
  assign n8709 = ~i_RtoB_ACK0 & ~n8708;
  assign n8710 = ~n8679 & ~n8709;
  assign n8711 = controllable_DEQ & ~n8710;
  assign n8712 = ~n8393 & ~n8697;
  assign n8713 = ~controllable_DEQ & ~n8712;
  assign n8714 = ~n8711 & ~n8713;
  assign n8715 = ~i_FULL & ~n8714;
  assign n8716 = ~n8701 & ~n8715;
  assign n8717 = i_nEMPTY & ~n8716;
  assign n8718 = ~controllable_ENQ & ~n8680;
  assign n8719 = i_RtoB_ACK1 & ~n8718;
  assign n8720 = ~n8407 & ~n8719;
  assign n8721 = controllable_BtoR_REQ1 & ~n8720;
  assign n8722 = ~n8409 & ~n8721;
  assign n8723 = ~controllable_BtoR_REQ0 & ~n8722;
  assign n8724 = ~controllable_BtoR_REQ0 & ~n8723;
  assign n8725 = ~i_RtoB_ACK0 & ~n8724;
  assign n8726 = ~i_RtoB_ACK0 & ~n8725;
  assign n8727 = controllable_DEQ & ~n8726;
  assign n8728 = ~n8421 & ~n8679;
  assign n8729 = ~controllable_DEQ & ~n8728;
  assign n8730 = ~n8727 & ~n8729;
  assign n8731 = i_FULL & ~n8730;
  assign n8732 = ~n8427 & ~n8693;
  assign n8733 = ~controllable_BtoR_REQ0 & ~n8732;
  assign n8734 = ~controllable_BtoR_REQ0 & ~n8733;
  assign n8735 = ~i_RtoB_ACK0 & ~n8734;
  assign n8736 = ~i_RtoB_ACK0 & ~n8735;
  assign n8737 = controllable_DEQ & ~n8736;
  assign n8738 = ~controllable_DEQ & ~n8689;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = ~i_FULL & ~n8739;
  assign n8741 = ~n8731 & ~n8740;
  assign n8742 = ~i_nEMPTY & ~n8741;
  assign n8743 = ~n8717 & ~n8742;
  assign n8744 = ~controllable_BtoS_ACK0 & ~n8743;
  assign n8745 = ~n8666 & ~n8744;
  assign n8746 = ~n4465 & ~n8745;
  assign n8747 = ~n8614 & ~n8746;
  assign n8748 = i_StoB_REQ10 & ~n8747;
  assign n8749 = ~n8451 & ~n8748;
  assign n8750 = ~controllable_BtoS_ACK10 & ~n8749;
  assign n8751 = ~n8453 & ~n8750;
  assign n8752 = ~n4464 & ~n8751;
  assign n8753 = ~n7687 & ~n8752;
  assign n8754 = n4463 & ~n8753;
  assign n8755 = ~i_RtoB_ACK1 & ~n5231;
  assign n8756 = ~n5032 & ~n8755;
  assign n8757 = ~controllable_BtoR_REQ1 & ~n8756;
  assign n8758 = ~n5019 & ~n8757;
  assign n8759 = ~controllable_BtoR_REQ0 & ~n8758;
  assign n8760 = ~controllable_BtoR_REQ0 & ~n8759;
  assign n8761 = i_RtoB_ACK0 & ~n8760;
  assign n8762 = ~n5035 & ~n5237;
  assign n8763 = controllable_BtoR_REQ1 & ~n8762;
  assign n8764 = ~n5025 & ~n5271;
  assign n8765 = ~i_RtoB_ACK1 & ~n8764;
  assign n8766 = ~n5032 & ~n8765;
  assign n8767 = ~controllable_BtoR_REQ1 & ~n8766;
  assign n8768 = ~n8763 & ~n8767;
  assign n8769 = ~controllable_BtoR_REQ0 & ~n8768;
  assign n8770 = ~controllable_BtoR_REQ0 & ~n8769;
  assign n8771 = ~i_RtoB_ACK0 & ~n8770;
  assign n8772 = ~n8761 & ~n8771;
  assign n8773 = controllable_DEQ & ~n8772;
  assign n8774 = i_RtoB_ACK1 & ~n5024;
  assign n8775 = ~n5243 & ~n8774;
  assign n8776 = ~controllable_BtoR_REQ1 & ~n8775;
  assign n8777 = ~n5049 & ~n8776;
  assign n8778 = ~controllable_BtoR_REQ0 & ~n8777;
  assign n8779 = ~controllable_BtoR_REQ0 & ~n8778;
  assign n8780 = i_RtoB_ACK0 & ~n8779;
  assign n8781 = ~n5038 & ~n7563;
  assign n8782 = controllable_BtoR_REQ1 & ~n8781;
  assign n8783 = ~n5050 & ~n8782;
  assign n8784 = ~controllable_BtoR_REQ0 & ~n8783;
  assign n8785 = ~controllable_BtoR_REQ0 & ~n8784;
  assign n8786 = ~i_RtoB_ACK0 & ~n8785;
  assign n8787 = ~n8780 & ~n8786;
  assign n8788 = ~controllable_DEQ & ~n8787;
  assign n8789 = ~n8773 & ~n8788;
  assign n8790 = i_FULL & ~n8789;
  assign n8791 = ~n5032 & ~n5243;
  assign n8792 = ~controllable_BtoR_REQ1 & ~n8791;
  assign n8793 = ~n8763 & ~n8792;
  assign n8794 = ~controllable_BtoR_REQ0 & ~n8793;
  assign n8795 = ~controllable_BtoR_REQ0 & ~n8794;
  assign n8796 = ~i_RtoB_ACK0 & ~n8795;
  assign n8797 = ~n8761 & ~n8796;
  assign n8798 = controllable_DEQ & ~n8797;
  assign n8799 = ~n8765 & ~n8774;
  assign n8800 = ~controllable_BtoR_REQ1 & ~n8799;
  assign n8801 = ~n8782 & ~n8800;
  assign n8802 = ~controllable_BtoR_REQ0 & ~n8801;
  assign n8803 = ~controllable_BtoR_REQ0 & ~n8802;
  assign n8804 = ~i_RtoB_ACK0 & ~n8803;
  assign n8805 = ~n8780 & ~n8804;
  assign n8806 = ~controllable_DEQ & ~n8805;
  assign n8807 = ~n8798 & ~n8806;
  assign n8808 = ~i_FULL & ~n8807;
  assign n8809 = ~n8790 & ~n8808;
  assign n8810 = i_nEMPTY & ~n8809;
  assign n8811 = ~n5065 & ~n5275;
  assign n8812 = ~controllable_BtoR_REQ0 & ~n8811;
  assign n8813 = ~controllable_BtoR_REQ0 & ~n8812;
  assign n8814 = ~i_RtoB_ACK0 & ~n8813;
  assign n8815 = ~i_RtoB_ACK0 & ~n8814;
  assign n8816 = controllable_DEQ & ~n8815;
  assign n8817 = ~i_RtoB_ACK1 & ~n5026;
  assign n8818 = ~n5237 & ~n8817;
  assign n8819 = controllable_BtoR_REQ1 & ~n8818;
  assign n8820 = ~n5027 & ~n8819;
  assign n8821 = ~controllable_BtoR_REQ0 & ~n8820;
  assign n8822 = ~controllable_BtoR_REQ0 & ~n8821;
  assign n8823 = ~i_RtoB_ACK0 & ~n8822;
  assign n8824 = ~n8761 & ~n8823;
  assign n8825 = ~controllable_DEQ & ~n8824;
  assign n8826 = ~n8816 & ~n8825;
  assign n8827 = i_FULL & ~n8826;
  assign n8828 = ~n5049 & ~n5290;
  assign n8829 = ~controllable_BtoR_REQ0 & ~n8828;
  assign n8830 = ~controllable_BtoR_REQ0 & ~n8829;
  assign n8831 = ~i_RtoB_ACK0 & ~n8830;
  assign n8832 = ~i_RtoB_ACK0 & ~n8831;
  assign n8833 = controllable_DEQ & ~n8832;
  assign n8834 = ~n5025 & ~n5238;
  assign n8835 = ~i_RtoB_ACK1 & ~n8834;
  assign n8836 = ~n5032 & ~n8835;
  assign n8837 = ~controllable_BtoR_REQ1 & ~n8836;
  assign n8838 = ~n8763 & ~n8837;
  assign n8839 = ~controllable_BtoR_REQ0 & ~n8838;
  assign n8840 = ~controllable_BtoR_REQ0 & ~n8839;
  assign n8841 = ~i_RtoB_ACK0 & ~n8840;
  assign n8842 = ~n8761 & ~n8841;
  assign n8843 = ~controllable_DEQ & ~n8842;
  assign n8844 = ~n8833 & ~n8843;
  assign n8845 = ~i_FULL & ~n8844;
  assign n8846 = ~n8827 & ~n8845;
  assign n8847 = ~i_nEMPTY & ~n8846;
  assign n8848 = ~n8810 & ~n8847;
  assign n8849 = controllable_BtoS_ACK0 & ~n8848;
  assign n8850 = ~controllable_BtoS_ACK14 & ~n5213;
  assign n8851 = ~n7793 & ~n8850;
  assign n8852 = controllable_ENQ & ~n8851;
  assign n8853 = controllable_ENQ & ~n8852;
  assign n8854 = ~i_RtoB_ACK1 & ~n8853;
  assign n8855 = ~n5129 & ~n8854;
  assign n8856 = ~controllable_BtoR_REQ1 & ~n8855;
  assign n8857 = ~n5116 & ~n8856;
  assign n8858 = ~controllable_BtoR_REQ0 & ~n8857;
  assign n8859 = ~controllable_BtoR_REQ0 & ~n8858;
  assign n8860 = i_RtoB_ACK0 & ~n8859;
  assign n8861 = i_RtoB_ACK1 & ~n8853;
  assign n8862 = ~n5132 & ~n8861;
  assign n8863 = controllable_BtoR_REQ1 & ~n8862;
  assign n8864 = ~controllable_ENQ & ~n8851;
  assign n8865 = ~n5122 & ~n8864;
  assign n8866 = ~i_RtoB_ACK1 & ~n8865;
  assign n8867 = ~n5129 & ~n8866;
  assign n8868 = ~controllable_BtoR_REQ1 & ~n8867;
  assign n8869 = ~n8863 & ~n8868;
  assign n8870 = ~controllable_BtoR_REQ0 & ~n8869;
  assign n8871 = ~controllable_BtoR_REQ0 & ~n8870;
  assign n8872 = ~i_RtoB_ACK0 & ~n8871;
  assign n8873 = ~n8860 & ~n8872;
  assign n8874 = controllable_DEQ & ~n8873;
  assign n8875 = i_RtoB_ACK1 & ~n5121;
  assign n8876 = ~i_RtoB_ACK1 & ~n8851;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~controllable_BtoR_REQ1 & ~n8877;
  assign n8879 = ~n5146 & ~n8878;
  assign n8880 = ~controllable_BtoR_REQ0 & ~n8879;
  assign n8881 = ~controllable_BtoR_REQ0 & ~n8880;
  assign n8882 = i_RtoB_ACK0 & ~n8881;
  assign n8883 = i_RtoB_ACK1 & ~n8851;
  assign n8884 = ~n5135 & ~n8883;
  assign n8885 = controllable_BtoR_REQ1 & ~n8884;
  assign n8886 = ~n5147 & ~n8885;
  assign n8887 = ~controllable_BtoR_REQ0 & ~n8886;
  assign n8888 = ~controllable_BtoR_REQ0 & ~n8887;
  assign n8889 = ~i_RtoB_ACK0 & ~n8888;
  assign n8890 = ~n8882 & ~n8889;
  assign n8891 = ~controllable_DEQ & ~n8890;
  assign n8892 = ~n8874 & ~n8891;
  assign n8893 = i_FULL & ~n8892;
  assign n8894 = ~n5129 & ~n8876;
  assign n8895 = ~controllable_BtoR_REQ1 & ~n8894;
  assign n8896 = ~n8863 & ~n8895;
  assign n8897 = ~controllable_BtoR_REQ0 & ~n8896;
  assign n8898 = ~controllable_BtoR_REQ0 & ~n8897;
  assign n8899 = ~i_RtoB_ACK0 & ~n8898;
  assign n8900 = ~n8860 & ~n8899;
  assign n8901 = controllable_DEQ & ~n8900;
  assign n8902 = ~n8866 & ~n8875;
  assign n8903 = ~controllable_BtoR_REQ1 & ~n8902;
  assign n8904 = ~n8885 & ~n8903;
  assign n8905 = ~controllable_BtoR_REQ0 & ~n8904;
  assign n8906 = ~controllable_BtoR_REQ0 & ~n8905;
  assign n8907 = ~i_RtoB_ACK0 & ~n8906;
  assign n8908 = ~n8882 & ~n8907;
  assign n8909 = ~controllable_DEQ & ~n8908;
  assign n8910 = ~n8901 & ~n8909;
  assign n8911 = ~i_FULL & ~n8910;
  assign n8912 = ~n8893 & ~n8911;
  assign n8913 = i_nEMPTY & ~n8912;
  assign n8914 = ~controllable_ENQ & ~n8864;
  assign n8915 = ~i_RtoB_ACK1 & ~n8914;
  assign n8916 = ~i_RtoB_ACK1 & ~n8915;
  assign n8917 = ~controllable_BtoR_REQ1 & ~n8916;
  assign n8918 = ~n5162 & ~n8917;
  assign n8919 = ~controllable_BtoR_REQ0 & ~n8918;
  assign n8920 = ~controllable_BtoR_REQ0 & ~n8919;
  assign n8921 = ~i_RtoB_ACK0 & ~n8920;
  assign n8922 = ~i_RtoB_ACK0 & ~n8921;
  assign n8923 = controllable_DEQ & ~n8922;
  assign n8924 = ~i_RtoB_ACK1 & ~n5123;
  assign n8925 = ~n8861 & ~n8924;
  assign n8926 = controllable_BtoR_REQ1 & ~n8925;
  assign n8927 = ~n5124 & ~n8926;
  assign n8928 = ~controllable_BtoR_REQ0 & ~n8927;
  assign n8929 = ~controllable_BtoR_REQ0 & ~n8928;
  assign n8930 = ~i_RtoB_ACK0 & ~n8929;
  assign n8931 = ~n8860 & ~n8930;
  assign n8932 = ~controllable_DEQ & ~n8931;
  assign n8933 = ~n8923 & ~n8932;
  assign n8934 = i_FULL & ~n8933;
  assign n8935 = ~i_RtoB_ACK1 & ~n8876;
  assign n8936 = ~controllable_BtoR_REQ1 & ~n8935;
  assign n8937 = ~n5146 & ~n8936;
  assign n8938 = ~controllable_BtoR_REQ0 & ~n8937;
  assign n8939 = ~controllable_BtoR_REQ0 & ~n8938;
  assign n8940 = ~i_RtoB_ACK0 & ~n8939;
  assign n8941 = ~i_RtoB_ACK0 & ~n8940;
  assign n8942 = controllable_DEQ & ~n8941;
  assign n8943 = ~n7782 & ~n8048;
  assign n8944 = ~controllable_BtoS_ACK14 & ~n8943;
  assign n8945 = ~n7784 & ~n8944;
  assign n8946 = ~controllable_ENQ & ~n8945;
  assign n8947 = ~n5122 & ~n8946;
  assign n8948 = ~i_RtoB_ACK1 & ~n8947;
  assign n8949 = ~n5129 & ~n8948;
  assign n8950 = ~controllable_BtoR_REQ1 & ~n8949;
  assign n8951 = ~n8863 & ~n8950;
  assign n8952 = ~controllable_BtoR_REQ0 & ~n8951;
  assign n8953 = ~controllable_BtoR_REQ0 & ~n8952;
  assign n8954 = ~i_RtoB_ACK0 & ~n8953;
  assign n8955 = ~n8860 & ~n8954;
  assign n8956 = ~controllable_DEQ & ~n8955;
  assign n8957 = ~n8942 & ~n8956;
  assign n8958 = ~i_FULL & ~n8957;
  assign n8959 = ~n8934 & ~n8958;
  assign n8960 = ~i_nEMPTY & ~n8959;
  assign n8961 = ~n8913 & ~n8960;
  assign n8962 = ~controllable_BtoS_ACK0 & ~n8961;
  assign n8963 = ~n8849 & ~n8962;
  assign n8964 = n4465 & ~n8963;
  assign n8965 = ~n5343 & ~n8854;
  assign n8966 = ~controllable_BtoR_REQ1 & ~n8965;
  assign n8967 = ~n5330 & ~n8966;
  assign n8968 = ~controllable_BtoR_REQ0 & ~n8967;
  assign n8969 = ~controllable_BtoR_REQ0 & ~n8968;
  assign n8970 = i_RtoB_ACK0 & ~n8969;
  assign n8971 = ~n5346 & ~n8861;
  assign n8972 = controllable_BtoR_REQ1 & ~n8971;
  assign n8973 = ~n5336 & ~n8864;
  assign n8974 = ~i_RtoB_ACK1 & ~n8973;
  assign n8975 = ~n5343 & ~n8974;
  assign n8976 = ~controllable_BtoR_REQ1 & ~n8975;
  assign n8977 = ~n8972 & ~n8976;
  assign n8978 = ~controllable_BtoR_REQ0 & ~n8977;
  assign n8979 = ~controllable_BtoR_REQ0 & ~n8978;
  assign n8980 = ~i_RtoB_ACK0 & ~n8979;
  assign n8981 = ~n8970 & ~n8980;
  assign n8982 = controllable_DEQ & ~n8981;
  assign n8983 = i_RtoB_ACK1 & ~n5335;
  assign n8984 = ~n8876 & ~n8983;
  assign n8985 = ~controllable_BtoR_REQ1 & ~n8984;
  assign n8986 = ~n5360 & ~n8985;
  assign n8987 = ~controllable_BtoR_REQ0 & ~n8986;
  assign n8988 = ~controllable_BtoR_REQ0 & ~n8987;
  assign n8989 = i_RtoB_ACK0 & ~n8988;
  assign n8990 = ~n5349 & ~n8883;
  assign n8991 = controllable_BtoR_REQ1 & ~n8990;
  assign n8992 = ~n5361 & ~n8991;
  assign n8993 = ~controllable_BtoR_REQ0 & ~n8992;
  assign n8994 = ~controllable_BtoR_REQ0 & ~n8993;
  assign n8995 = ~i_RtoB_ACK0 & ~n8994;
  assign n8996 = ~n8989 & ~n8995;
  assign n8997 = ~controllable_DEQ & ~n8996;
  assign n8998 = ~n8982 & ~n8997;
  assign n8999 = i_FULL & ~n8998;
  assign n9000 = ~n5343 & ~n8876;
  assign n9001 = ~controllable_BtoR_REQ1 & ~n9000;
  assign n9002 = ~n8972 & ~n9001;
  assign n9003 = ~controllable_BtoR_REQ0 & ~n9002;
  assign n9004 = ~controllable_BtoR_REQ0 & ~n9003;
  assign n9005 = ~i_RtoB_ACK0 & ~n9004;
  assign n9006 = ~n8970 & ~n9005;
  assign n9007 = controllable_DEQ & ~n9006;
  assign n9008 = ~n8974 & ~n8983;
  assign n9009 = ~controllable_BtoR_REQ1 & ~n9008;
  assign n9010 = ~n8991 & ~n9009;
  assign n9011 = ~controllable_BtoR_REQ0 & ~n9010;
  assign n9012 = ~controllable_BtoR_REQ0 & ~n9011;
  assign n9013 = ~i_RtoB_ACK0 & ~n9012;
  assign n9014 = ~n8989 & ~n9013;
  assign n9015 = ~controllable_DEQ & ~n9014;
  assign n9016 = ~n9007 & ~n9015;
  assign n9017 = ~i_FULL & ~n9016;
  assign n9018 = ~n8999 & ~n9017;
  assign n9019 = i_nEMPTY & ~n9018;
  assign n9020 = ~n5376 & ~n8917;
  assign n9021 = ~controllable_BtoR_REQ0 & ~n9020;
  assign n9022 = ~controllable_BtoR_REQ0 & ~n9021;
  assign n9023 = ~i_RtoB_ACK0 & ~n9022;
  assign n9024 = ~i_RtoB_ACK0 & ~n9023;
  assign n9025 = controllable_DEQ & ~n9024;
  assign n9026 = ~i_RtoB_ACK1 & ~n5337;
  assign n9027 = ~n8861 & ~n9026;
  assign n9028 = controllable_BtoR_REQ1 & ~n9027;
  assign n9029 = ~n5338 & ~n9028;
  assign n9030 = ~controllable_BtoR_REQ0 & ~n9029;
  assign n9031 = ~controllable_BtoR_REQ0 & ~n9030;
  assign n9032 = ~i_RtoB_ACK0 & ~n9031;
  assign n9033 = ~n8970 & ~n9032;
  assign n9034 = ~controllable_DEQ & ~n9033;
  assign n9035 = ~n9025 & ~n9034;
  assign n9036 = i_FULL & ~n9035;
  assign n9037 = ~n5360 & ~n8936;
  assign n9038 = ~controllable_BtoR_REQ0 & ~n9037;
  assign n9039 = ~controllable_BtoR_REQ0 & ~n9038;
  assign n9040 = ~i_RtoB_ACK0 & ~n9039;
  assign n9041 = ~i_RtoB_ACK0 & ~n9040;
  assign n9042 = controllable_DEQ & ~n9041;
  assign n9043 = ~n5336 & ~n8946;
  assign n9044 = ~i_RtoB_ACK1 & ~n9043;
  assign n9045 = ~n5343 & ~n9044;
  assign n9046 = ~controllable_BtoR_REQ1 & ~n9045;
  assign n9047 = ~n8972 & ~n9046;
  assign n9048 = ~controllable_BtoR_REQ0 & ~n9047;
  assign n9049 = ~controllable_BtoR_REQ0 & ~n9048;
  assign n9050 = ~i_RtoB_ACK0 & ~n9049;
  assign n9051 = ~n8970 & ~n9050;
  assign n9052 = ~controllable_DEQ & ~n9051;
  assign n9053 = ~n9042 & ~n9052;
  assign n9054 = ~i_FULL & ~n9053;
  assign n9055 = ~n9036 & ~n9054;
  assign n9056 = ~i_nEMPTY & ~n9055;
  assign n9057 = ~n9019 & ~n9056;
  assign n9058 = ~controllable_BtoS_ACK0 & ~n9057;
  assign n9059 = ~n5307 & ~n9058;
  assign n9060 = ~n4465 & ~n9059;
  assign n9061 = ~n8964 & ~n9060;
  assign n9062 = i_StoB_REQ10 & ~n9061;
  assign n9063 = n4467 & ~n4669;
  assign n9064 = ~n4477 & ~n4483;
  assign n9065 = ~n4697 & ~n9064;
  assign n9066 = n4476 & ~n9065;
  assign n9067 = ~n4476 & ~n4483;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = ~i_StoB_REQ3 & ~n9068;
  assign n9070 = ~i_StoB_REQ3 & ~n9069;
  assign n9071 = controllable_BtoS_ACK3 & ~n9070;
  assign n9072 = ~n4741 & ~n9069;
  assign n9073 = ~controllable_BtoS_ACK3 & ~n9072;
  assign n9074 = ~n9071 & ~n9073;
  assign n9075 = n4475 & ~n9074;
  assign n9076 = ~n4475 & ~n4525;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = ~i_StoB_REQ4 & ~n9077;
  assign n9079 = ~i_StoB_REQ4 & ~n9078;
  assign n9080 = controllable_BtoS_ACK4 & ~n9079;
  assign n9081 = ~n4768 & ~n9078;
  assign n9082 = ~controllable_BtoS_ACK4 & ~n9081;
  assign n9083 = ~n9080 & ~n9082;
  assign n9084 = n4474 & ~n9083;
  assign n9085 = ~n4474 & ~n4546;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = ~i_StoB_REQ5 & ~n9086;
  assign n9088 = ~i_StoB_REQ5 & ~n9087;
  assign n9089 = controllable_BtoS_ACK5 & ~n9088;
  assign n9090 = ~n4795 & ~n9087;
  assign n9091 = ~controllable_BtoS_ACK5 & ~n9090;
  assign n9092 = ~n9089 & ~n9091;
  assign n9093 = n4473 & ~n9092;
  assign n9094 = ~n4473 & ~n4567;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~i_StoB_REQ8 & ~n9095;
  assign n9097 = ~i_StoB_REQ8 & ~n9096;
  assign n9098 = controllable_BtoS_ACK8 & ~n9097;
  assign n9099 = ~n4815 & ~n9096;
  assign n9100 = ~controllable_BtoS_ACK8 & ~n9099;
  assign n9101 = ~n9098 & ~n9100;
  assign n9102 = n4472 & ~n9101;
  assign n9103 = ~n4472 & ~n4583;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = n4471 & ~n9104;
  assign n9106 = ~n4584 & ~n9105;
  assign n9107 = ~i_StoB_REQ6 & ~n9106;
  assign n9108 = ~i_StoB_REQ6 & ~n9107;
  assign n9109 = controllable_BtoS_ACK6 & ~n9108;
  assign n9110 = ~n4847 & ~n9107;
  assign n9111 = ~controllable_BtoS_ACK6 & ~n9110;
  assign n9112 = ~n9109 & ~n9111;
  assign n9113 = ~i_StoB_REQ7 & ~n9112;
  assign n9114 = ~i_StoB_REQ7 & ~n9113;
  assign n9115 = controllable_BtoS_ACK7 & ~n9114;
  assign n9116 = ~n4872 & ~n9113;
  assign n9117 = ~controllable_BtoS_ACK7 & ~n9116;
  assign n9118 = ~n9115 & ~n9117;
  assign n9119 = n4470 & ~n9118;
  assign n9120 = ~n4470 & ~n4626;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = n4469 & ~n9121;
  assign n9123 = ~n4627 & ~n9122;
  assign n9124 = ~i_StoB_REQ9 & ~n9123;
  assign n9125 = ~i_StoB_REQ9 & ~n9124;
  assign n9126 = controllable_BtoS_ACK9 & ~n9125;
  assign n9127 = ~n4897 & ~n9124;
  assign n9128 = ~controllable_BtoS_ACK9 & ~n9127;
  assign n9129 = ~n9126 & ~n9128;
  assign n9130 = n4468 & ~n9129;
  assign n9131 = ~n4648 & ~n9130;
  assign n9132 = ~i_StoB_REQ11 & ~n9131;
  assign n9133 = ~i_StoB_REQ11 & ~n9132;
  assign n9134 = controllable_BtoS_ACK11 & ~n9133;
  assign n9135 = ~n4927 & ~n9132;
  assign n9136 = ~controllable_BtoS_ACK11 & ~n9135;
  assign n9137 = ~n9134 & ~n9136;
  assign n9138 = ~n4467 & ~n9137;
  assign n9139 = ~n9063 & ~n9138;
  assign n9140 = i_StoB_REQ12 & ~n9139;
  assign n9141 = n4468 & ~n4647;
  assign n9142 = ~n4468 & ~n9129;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 = i_StoB_REQ11 & ~n9143;
  assign n9145 = n4469 & ~n4626;
  assign n9146 = ~n4469 & ~n9121;
  assign n9147 = ~n9145 & ~n9146;
  assign n9148 = i_StoB_REQ9 & ~n9147;
  assign n9149 = n4471 & ~n4583;
  assign n9150 = ~n4471 & ~n9104;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = i_StoB_REQ6 & ~n9151;
  assign n9153 = i_StoB_REQ2 & ~n4689;
  assign n9154 = controllable_BtoS_ACK2 & n9153;
  assign n9155 = ~n4477 & n9154;
  assign n9156 = ~n5864 & ~n9155;
  assign n9157 = n4476 & ~n9156;
  assign n9158 = controllable_BtoS_ACK2 & n4478;
  assign n9159 = ~i_StoB_REQ2 & ~n4478;
  assign n9160 = ~i_StoB_REQ2 & ~n9159;
  assign n9161 = ~controllable_BtoS_ACK2 & n9160;
  assign n9162 = ~n9158 & ~n9161;
  assign n9163 = n4477 & ~n9162;
  assign n9164 = ~n4477 & n5863;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~n4476 & ~n9165;
  assign n9167 = ~n9157 & ~n9166;
  assign n9168 = ~i_StoB_REQ3 & ~n9167;
  assign n9169 = ~n4741 & ~n9168;
  assign n9170 = controllable_BtoS_ACK3 & ~n9169;
  assign n9171 = ~n6250 & ~n9168;
  assign n9172 = ~controllable_BtoS_ACK3 & ~n9171;
  assign n9173 = ~n9170 & ~n9172;
  assign n9174 = n4475 & ~n9173;
  assign n9175 = i_StoB_REQ3 & ~n9068;
  assign n9176 = ~n5886 & ~n9175;
  assign n9177 = controllable_BtoS_ACK3 & ~n9176;
  assign n9178 = ~n5920 & ~n9177;
  assign n9179 = ~n4475 & ~n9178;
  assign n9180 = ~n9174 & ~n9179;
  assign n9181 = ~i_StoB_REQ4 & ~n9180;
  assign n9182 = ~n4768 & ~n9181;
  assign n9183 = controllable_BtoS_ACK4 & ~n9182;
  assign n9184 = ~n6283 & ~n9181;
  assign n9185 = ~controllable_BtoS_ACK4 & ~n9184;
  assign n9186 = ~n9183 & ~n9185;
  assign n9187 = n4474 & ~n9186;
  assign n9188 = i_StoB_REQ4 & ~n9077;
  assign n9189 = ~n5922 & ~n9188;
  assign n9190 = controllable_BtoS_ACK4 & ~n9189;
  assign n9191 = ~n5955 & ~n9190;
  assign n9192 = ~n4474 & ~n9191;
  assign n9193 = ~n9187 & ~n9192;
  assign n9194 = ~i_StoB_REQ5 & ~n9193;
  assign n9195 = ~n4795 & ~n9194;
  assign n9196 = controllable_BtoS_ACK5 & ~n9195;
  assign n9197 = ~n6316 & ~n9194;
  assign n9198 = ~controllable_BtoS_ACK5 & ~n9197;
  assign n9199 = ~n9196 & ~n9198;
  assign n9200 = n4473 & ~n9199;
  assign n9201 = i_StoB_REQ5 & ~n9086;
  assign n9202 = ~n5957 & ~n9201;
  assign n9203 = controllable_BtoS_ACK5 & ~n9202;
  assign n9204 = ~n5990 & ~n9203;
  assign n9205 = ~n4473 & ~n9204;
  assign n9206 = ~n9200 & ~n9205;
  assign n9207 = ~i_StoB_REQ8 & ~n9206;
  assign n9208 = ~n4815 & ~n9207;
  assign n9209 = controllable_BtoS_ACK8 & ~n9208;
  assign n9210 = ~n6341 & ~n9207;
  assign n9211 = ~controllable_BtoS_ACK8 & ~n9210;
  assign n9212 = ~n9209 & ~n9211;
  assign n9213 = n4472 & ~n9212;
  assign n9214 = i_StoB_REQ8 & ~n9095;
  assign n9215 = ~n5992 & ~n9214;
  assign n9216 = controllable_BtoS_ACK8 & ~n9215;
  assign n9217 = ~n6020 & ~n9216;
  assign n9218 = ~n4472 & ~n9217;
  assign n9219 = ~n9213 & ~n9218;
  assign n9220 = n4471 & ~n9219;
  assign n9221 = ~n6022 & ~n9220;
  assign n9222 = ~i_StoB_REQ6 & ~n9221;
  assign n9223 = ~n9152 & ~n9222;
  assign n9224 = controllable_BtoS_ACK6 & ~n9223;
  assign n9225 = ~n6377 & ~n9222;
  assign n9226 = ~controllable_BtoS_ACK6 & ~n9225;
  assign n9227 = ~n9224 & ~n9226;
  assign n9228 = ~i_StoB_REQ7 & ~n9227;
  assign n9229 = ~n4872 & ~n9228;
  assign n9230 = controllable_BtoS_ACK7 & ~n9229;
  assign n9231 = ~n6404 & ~n9228;
  assign n9232 = ~controllable_BtoS_ACK7 & ~n9231;
  assign n9233 = ~n9230 & ~n9232;
  assign n9234 = n4470 & ~n9233;
  assign n9235 = i_StoB_REQ7 & ~n9112;
  assign n9236 = ~n6062 & ~n9235;
  assign n9237 = controllable_BtoS_ACK7 & ~n9236;
  assign n9238 = ~n6093 & ~n9237;
  assign n9239 = ~n4470 & ~n9238;
  assign n9240 = ~n9234 & ~n9239;
  assign n9241 = n4469 & ~n9240;
  assign n9242 = ~n6095 & ~n9241;
  assign n9243 = ~i_StoB_REQ9 & ~n9242;
  assign n9244 = ~n9148 & ~n9243;
  assign n9245 = controllable_BtoS_ACK9 & ~n9244;
  assign n9246 = ~n6432 & ~n9243;
  assign n9247 = ~controllable_BtoS_ACK9 & ~n9246;
  assign n9248 = ~n9245 & ~n9247;
  assign n9249 = n4468 & ~n9248;
  assign n9250 = ~n6130 & ~n9249;
  assign n9251 = ~i_StoB_REQ11 & ~n9250;
  assign n9252 = ~n9144 & ~n9251;
  assign n9253 = controllable_BtoS_ACK11 & ~n9252;
  assign n9254 = ~n6462 & ~n9251;
  assign n9255 = ~controllable_BtoS_ACK11 & ~n9254;
  assign n9256 = ~n9253 & ~n9255;
  assign n9257 = n4467 & ~n9256;
  assign n9258 = ~n6168 & ~n9257;
  assign n9259 = ~i_StoB_REQ12 & ~n9258;
  assign n9260 = ~n9140 & ~n9259;
  assign n9261 = controllable_BtoS_ACK12 & ~n9260;
  assign n9262 = ~n6505 & ~n9259;
  assign n9263 = ~controllable_BtoS_ACK12 & ~n9262;
  assign n9264 = ~n9261 & ~n9263;
  assign n9265 = ~i_StoB_REQ13 & ~n9264;
  assign n9266 = ~n7068 & ~n9265;
  assign n9267 = n4466 & ~n9266;
  assign n9268 = n4467 & ~n9137;
  assign n9269 = ~n4670 & ~n9268;
  assign n9270 = ~i_StoB_REQ12 & ~n9269;
  assign n9271 = ~i_StoB_REQ12 & ~n9270;
  assign n9272 = controllable_BtoS_ACK12 & ~n9271;
  assign n9273 = ~n4969 & ~n9270;
  assign n9274 = ~controllable_BtoS_ACK12 & ~n9273;
  assign n9275 = ~n9272 & ~n9274;
  assign n9276 = controllable_BtoS_ACK13 & ~n9275;
  assign n9277 = ~n7057 & ~n9276;
  assign n9278 = i_StoB_REQ13 & ~n9277;
  assign n9279 = ~n7069 & ~n9278;
  assign n9280 = ~n4466 & ~n9279;
  assign n9281 = ~n9267 & ~n9280;
  assign n9282 = ~i_StoB_REQ0 & ~n9281;
  assign n9283 = ~n7172 & ~n9282;
  assign n9284 = ~i_StoB_REQ14 & ~n9283;
  assign n9285 = ~n5216 & ~n9284;
  assign n9286 = controllable_BtoS_ACK14 & ~n9285;
  assign n9287 = i_StoB_REQ14 & ~n7906;
  assign n9288 = ~n9284 & ~n9287;
  assign n9289 = ~controllable_BtoS_ACK14 & ~n9288;
  assign n9290 = ~n9286 & ~n9289;
  assign n9291 = controllable_ENQ & ~n9290;
  assign n9292 = controllable_ENQ & ~n9291;
  assign n9293 = ~i_RtoB_ACK1 & ~n9292;
  assign n9294 = ~n6773 & ~n9293;
  assign n9295 = ~controllable_BtoR_REQ1 & ~n9294;
  assign n9296 = ~n6573 & ~n9295;
  assign n9297 = ~controllable_BtoR_REQ0 & ~n9296;
  assign n9298 = ~controllable_BtoR_REQ0 & ~n9297;
  assign n9299 = i_RtoB_ACK0 & ~n9298;
  assign n9300 = ~controllable_BtoS_ACK14 & ~n7906;
  assign n9301 = ~n8223 & ~n9300;
  assign n9302 = controllable_ENQ & ~n9301;
  assign n9303 = ~n6765 & ~n9302;
  assign n9304 = i_RtoB_ACK1 & ~n9303;
  assign n9305 = ~n6770 & ~n9304;
  assign n9306 = controllable_BtoR_REQ1 & ~n9305;
  assign n9307 = i_StoB_REQ12 & ~n4671;
  assign n9308 = i_StoB_REQ11 & ~n4649;
  assign n9309 = i_StoB_REQ9 & ~n4628;
  assign n9310 = i_StoB_REQ6 & ~n4585;
  assign n9311 = controllable_BtoS_ACK2 & ~n5863;
  assign n9312 = ~n4477 & ~n9311;
  assign n9313 = ~n5864 & ~n9312;
  assign n9314 = n4476 & ~n9313;
  assign n9315 = ~i_StoB_REQ2 & ~controllable_BtoS_ACK1;
  assign n9316 = ~n4702 & ~n9315;
  assign n9317 = controllable_BtoS_ACK2 & ~n9316;
  assign n9318 = ~controllable_BtoS_ACK1 & ~controllable_BtoS_ACK2;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = n4477 & ~n9319;
  assign n9321 = ~n5863 & ~n9318;
  assign n9322 = ~n4477 & ~n9321;
  assign n9323 = ~n9320 & ~n9322;
  assign n9324 = ~n4476 & ~n9323;
  assign n9325 = ~n9314 & ~n9324;
  assign n9326 = ~i_StoB_REQ3 & ~n9325;
  assign n9327 = ~n4715 & ~n9326;
  assign n9328 = controllable_BtoS_ACK3 & ~n9327;
  assign n9329 = ~controllable_BtoS_ACK3 & ~n9325;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = n4475 & ~n9330;
  assign n9332 = ~n4477 & ~n9312;
  assign n9333 = n4476 & ~n9332;
  assign n9334 = ~n9324 & ~n9333;
  assign n9335 = ~controllable_BtoS_ACK3 & ~n9334;
  assign n9336 = ~n5919 & ~n9335;
  assign n9337 = ~n4475 & ~n9336;
  assign n9338 = ~n9331 & ~n9337;
  assign n9339 = ~i_StoB_REQ4 & ~n9338;
  assign n9340 = ~n4736 & ~n9339;
  assign n9341 = controllable_BtoS_ACK4 & ~n9340;
  assign n9342 = ~controllable_BtoS_ACK4 & ~n9338;
  assign n9343 = ~n9341 & ~n9342;
  assign n9344 = n4474 & ~n9343;
  assign n9345 = ~i_StoB_REQ3 & ~n9334;
  assign n9346 = ~n4723 & ~n9345;
  assign n9347 = controllable_BtoS_ACK3 & ~n9346;
  assign n9348 = ~n9335 & ~n9347;
  assign n9349 = n4475 & ~n9348;
  assign n9350 = ~n9337 & ~n9349;
  assign n9351 = ~controllable_BtoS_ACK4 & ~n9350;
  assign n9352 = ~n5954 & ~n9351;
  assign n9353 = ~n4474 & ~n9352;
  assign n9354 = ~n9344 & ~n9353;
  assign n9355 = ~i_StoB_REQ5 & ~n9354;
  assign n9356 = ~n4763 & ~n9355;
  assign n9357 = controllable_BtoS_ACK5 & ~n9356;
  assign n9358 = ~controllable_BtoS_ACK5 & ~n9354;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = n4473 & ~n9359;
  assign n9361 = ~i_StoB_REQ4 & ~n9350;
  assign n9362 = ~n4748 & ~n9361;
  assign n9363 = controllable_BtoS_ACK4 & ~n9362;
  assign n9364 = ~n9351 & ~n9363;
  assign n9365 = n4474 & ~n9364;
  assign n9366 = ~n9353 & ~n9365;
  assign n9367 = ~controllable_BtoS_ACK5 & ~n9366;
  assign n9368 = ~n5989 & ~n9367;
  assign n9369 = ~n4473 & ~n9368;
  assign n9370 = ~n9360 & ~n9369;
  assign n9371 = ~i_StoB_REQ8 & ~n9370;
  assign n9372 = ~n4790 & ~n9371;
  assign n9373 = controllable_BtoS_ACK8 & ~n9372;
  assign n9374 = ~controllable_BtoS_ACK8 & ~n9370;
  assign n9375 = ~n9373 & ~n9374;
  assign n9376 = n4472 & ~n9375;
  assign n9377 = ~i_StoB_REQ5 & ~n9366;
  assign n9378 = ~n4775 & ~n9377;
  assign n9379 = controllable_BtoS_ACK5 & ~n9378;
  assign n9380 = ~n9367 & ~n9379;
  assign n9381 = n4473 & ~n9380;
  assign n9382 = ~n9369 & ~n9381;
  assign n9383 = ~controllable_BtoS_ACK8 & ~n9382;
  assign n9384 = ~n6019 & ~n9383;
  assign n9385 = ~n4472 & ~n9384;
  assign n9386 = ~n9376 & ~n9385;
  assign n9387 = n4471 & ~n9386;
  assign n9388 = ~n6022 & ~n9387;
  assign n9389 = ~i_StoB_REQ6 & ~n9388;
  assign n9390 = ~n9310 & ~n9389;
  assign n9391 = controllable_BtoS_ACK6 & ~n9390;
  assign n9392 = ~i_StoB_REQ8 & ~n9382;
  assign n9393 = ~n4802 & ~n9392;
  assign n9394 = controllable_BtoS_ACK8 & ~n9393;
  assign n9395 = ~n9383 & ~n9394;
  assign n9396 = n4472 & ~n9395;
  assign n9397 = ~n9385 & ~n9396;
  assign n9398 = ~n4471 & ~n9397;
  assign n9399 = ~n9387 & ~n9398;
  assign n9400 = ~controllable_BtoS_ACK6 & ~n9399;
  assign n9401 = ~n9391 & ~n9400;
  assign n9402 = ~i_StoB_REQ7 & ~n9401;
  assign n9403 = ~n4839 & ~n9402;
  assign n9404 = controllable_BtoS_ACK7 & ~n9403;
  assign n9405 = ~controllable_BtoS_ACK7 & ~n9401;
  assign n9406 = ~n9404 & ~n9405;
  assign n9407 = n4470 & ~n9406;
  assign n9408 = i_StoB_REQ6 & ~n4614;
  assign n9409 = n4471 & ~n9397;
  assign n9410 = ~n6022 & ~n9409;
  assign n9411 = ~i_StoB_REQ6 & ~n9410;
  assign n9412 = ~n9408 & ~n9411;
  assign n9413 = controllable_BtoS_ACK6 & ~n9412;
  assign n9414 = ~controllable_BtoS_ACK6 & ~n9397;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = ~controllable_BtoS_ACK7 & ~n9415;
  assign n9417 = ~n6092 & ~n9416;
  assign n9418 = ~n4470 & ~n9417;
  assign n9419 = ~n9407 & ~n9418;
  assign n9420 = n4469 & ~n9419;
  assign n9421 = ~n6095 & ~n9420;
  assign n9422 = ~i_StoB_REQ9 & ~n9421;
  assign n9423 = ~n9309 & ~n9422;
  assign n9424 = controllable_BtoS_ACK9 & ~n9423;
  assign n9425 = ~i_StoB_REQ7 & ~n9415;
  assign n9426 = ~n4854 & ~n9425;
  assign n9427 = controllable_BtoS_ACK7 & ~n9426;
  assign n9428 = ~n9416 & ~n9427;
  assign n9429 = n4470 & ~n9428;
  assign n9430 = ~n9418 & ~n9429;
  assign n9431 = ~n4469 & ~n9430;
  assign n9432 = ~n9420 & ~n9431;
  assign n9433 = ~controllable_BtoS_ACK9 & ~n9432;
  assign n9434 = ~n9424 & ~n9433;
  assign n9435 = n4468 & ~n9434;
  assign n9436 = ~n6130 & ~n9435;
  assign n9437 = ~i_StoB_REQ11 & ~n9436;
  assign n9438 = ~n9308 & ~n9437;
  assign n9439 = controllable_BtoS_ACK11 & ~n9438;
  assign n9440 = i_StoB_REQ9 & ~n4654;
  assign n9441 = n4469 & ~n9430;
  assign n9442 = ~n6095 & ~n9441;
  assign n9443 = ~i_StoB_REQ9 & ~n9442;
  assign n9444 = ~n9440 & ~n9443;
  assign n9445 = controllable_BtoS_ACK9 & ~n9444;
  assign n9446 = ~controllable_BtoS_ACK9 & ~n9430;
  assign n9447 = ~n9445 & ~n9446;
  assign n9448 = ~n4468 & ~n9447;
  assign n9449 = ~n9435 & ~n9448;
  assign n9450 = ~controllable_BtoS_ACK11 & ~n9449;
  assign n9451 = ~n9439 & ~n9450;
  assign n9452 = n4467 & ~n9451;
  assign n9453 = ~n6168 & ~n9452;
  assign n9454 = ~i_StoB_REQ12 & ~n9453;
  assign n9455 = ~n9307 & ~n9454;
  assign n9456 = controllable_BtoS_ACK12 & ~n9455;
  assign n9457 = i_StoB_REQ11 & ~n4676;
  assign n9458 = n4468 & ~n9447;
  assign n9459 = ~n6130 & ~n9458;
  assign n9460 = ~i_StoB_REQ11 & ~n9459;
  assign n9461 = ~n9457 & ~n9460;
  assign n9462 = controllable_BtoS_ACK11 & ~n9461;
  assign n9463 = ~controllable_BtoS_ACK11 & ~n9447;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = ~n4467 & ~n9464;
  assign n9466 = ~n9452 & ~n9465;
  assign n9467 = ~controllable_BtoS_ACK12 & ~n9466;
  assign n9468 = ~n9456 & ~n9467;
  assign n9469 = ~controllable_BtoS_ACK13 & ~n9468;
  assign n9470 = ~n6534 & ~n9469;
  assign n9471 = i_StoB_REQ13 & ~n9470;
  assign n9472 = ~i_StoB_REQ13 & ~n9468;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = n4466 & ~n9473;
  assign n9475 = i_StoB_REQ12 & ~n4957;
  assign n9476 = n4467 & ~n9464;
  assign n9477 = ~n6168 & ~n9476;
  assign n9478 = ~i_StoB_REQ12 & ~n9477;
  assign n9479 = ~n9475 & ~n9478;
  assign n9480 = controllable_BtoS_ACK12 & ~n9479;
  assign n9481 = ~controllable_BtoS_ACK12 & ~n9464;
  assign n9482 = ~n9480 & ~n9481;
  assign n9483 = ~controllable_BtoS_ACK13 & ~n9482;
  assign n9484 = ~n5003 & ~n9483;
  assign n9485 = i_StoB_REQ13 & ~n9484;
  assign n9486 = ~n6548 & ~n9483;
  assign n9487 = ~i_StoB_REQ13 & ~n9486;
  assign n9488 = ~n9485 & ~n9487;
  assign n9489 = ~n4466 & ~n9488;
  assign n9490 = ~n9474 & ~n9489;
  assign n9491 = ~i_StoB_REQ0 & ~n9490;
  assign n9492 = ~n5103 & ~n9491;
  assign n9493 = ~i_StoB_REQ14 & ~n9492;
  assign n9494 = ~n5011 & ~n9493;
  assign n9495 = controllable_BtoS_ACK14 & ~n9494;
  assign n9496 = ~controllable_BtoS_ACK14 & ~n9492;
  assign n9497 = ~n9495 & ~n9496;
  assign n9498 = controllable_ENQ & ~n9497;
  assign n9499 = ~controllable_ENQ & ~n9290;
  assign n9500 = ~n9498 & ~n9499;
  assign n9501 = ~i_RtoB_ACK1 & ~n9500;
  assign n9502 = ~n6773 & ~n9501;
  assign n9503 = ~controllable_BtoR_REQ1 & ~n9502;
  assign n9504 = ~n9306 & ~n9503;
  assign n9505 = ~controllable_BtoR_REQ0 & ~n9504;
  assign n9506 = ~controllable_BtoR_REQ0 & ~n9505;
  assign n9507 = ~i_RtoB_ACK0 & ~n9506;
  assign n9508 = ~n9299 & ~n9507;
  assign n9509 = controllable_DEQ & ~n9508;
  assign n9510 = ~i_RtoB_ACK1 & ~n9290;
  assign n9511 = ~n6795 & ~n9510;
  assign n9512 = ~controllable_BtoR_REQ1 & ~n9511;
  assign n9513 = ~n6788 & ~n9512;
  assign n9514 = ~controllable_BtoR_REQ0 & ~n9513;
  assign n9515 = ~controllable_BtoR_REQ0 & ~n9514;
  assign n9516 = i_RtoB_ACK0 & ~n9515;
  assign n9517 = i_RtoB_ACK1 & ~n9301;
  assign n9518 = ~n6796 & ~n9517;
  assign n9519 = controllable_BtoR_REQ1 & ~n9518;
  assign n9520 = ~i_RtoB_ACK1 & ~n9497;
  assign n9521 = ~n6795 & ~n9520;
  assign n9522 = ~controllable_BtoR_REQ1 & ~n9521;
  assign n9523 = ~n9519 & ~n9522;
  assign n9524 = ~controllable_BtoR_REQ0 & ~n9523;
  assign n9525 = ~controllable_BtoR_REQ0 & ~n9524;
  assign n9526 = ~i_RtoB_ACK0 & ~n9525;
  assign n9527 = ~n9516 & ~n9526;
  assign n9528 = ~controllable_DEQ & ~n9527;
  assign n9529 = ~n9509 & ~n9528;
  assign n9530 = i_FULL & ~n9529;
  assign n9531 = ~n6810 & ~n9304;
  assign n9532 = controllable_BtoR_REQ1 & ~n9531;
  assign n9533 = ~n9302 & ~n9499;
  assign n9534 = ~i_RtoB_ACK1 & ~n9533;
  assign n9535 = ~n6773 & ~n9534;
  assign n9536 = ~controllable_BtoR_REQ1 & ~n9535;
  assign n9537 = ~n9532 & ~n9536;
  assign n9538 = ~controllable_BtoR_REQ0 & ~n9537;
  assign n9539 = ~controllable_BtoR_REQ0 & ~n9538;
  assign n9540 = ~i_RtoB_ACK0 & ~n9539;
  assign n9541 = ~n9299 & ~n9540;
  assign n9542 = controllable_DEQ & ~n9541;
  assign n9543 = ~n6776 & ~n9517;
  assign n9544 = controllable_BtoR_REQ1 & ~n9543;
  assign n9545 = ~controllable_ENQ & ~n9301;
  assign n9546 = ~n9498 & ~n9545;
  assign n9547 = ~i_RtoB_ACK1 & ~n9546;
  assign n9548 = ~n6795 & ~n9547;
  assign n9549 = ~controllable_BtoR_REQ1 & ~n9548;
  assign n9550 = ~n9544 & ~n9549;
  assign n9551 = ~controllable_BtoR_REQ0 & ~n9550;
  assign n9552 = ~controllable_BtoR_REQ0 & ~n9551;
  assign n9553 = ~i_RtoB_ACK0 & ~n9552;
  assign n9554 = ~n9516 & ~n9553;
  assign n9555 = ~controllable_DEQ & ~n9554;
  assign n9556 = ~n9542 & ~n9555;
  assign n9557 = ~i_FULL & ~n9556;
  assign n9558 = ~n9530 & ~n9557;
  assign n9559 = i_nEMPTY & ~n9558;
  assign n9560 = ~controllable_ENQ & ~n9499;
  assign n9561 = ~i_RtoB_ACK1 & ~n9560;
  assign n9562 = ~i_RtoB_ACK1 & ~n9561;
  assign n9563 = ~controllable_BtoR_REQ1 & ~n9562;
  assign n9564 = ~n6840 & ~n9563;
  assign n9565 = ~controllable_BtoR_REQ0 & ~n9564;
  assign n9566 = ~controllable_BtoR_REQ0 & ~n9565;
  assign n9567 = ~i_RtoB_ACK0 & ~n9566;
  assign n9568 = ~i_RtoB_ACK0 & ~n9567;
  assign n9569 = controllable_DEQ & ~n9568;
  assign n9570 = controllable_ENQ & ~n9302;
  assign n9571 = i_RtoB_ACK1 & ~n9570;
  assign n9572 = ~n6853 & ~n9571;
  assign n9573 = controllable_BtoR_REQ1 & ~n9572;
  assign n9574 = controllable_ENQ & ~n9498;
  assign n9575 = ~i_RtoB_ACK1 & ~n9574;
  assign n9576 = ~n6773 & ~n9575;
  assign n9577 = ~controllable_BtoR_REQ1 & ~n9576;
  assign n9578 = ~n9573 & ~n9577;
  assign n9579 = ~controllable_BtoR_REQ0 & ~n9578;
  assign n9580 = ~controllable_BtoR_REQ0 & ~n9579;
  assign n9581 = ~i_RtoB_ACK0 & ~n9580;
  assign n9582 = ~n9299 & ~n9581;
  assign n9583 = ~controllable_DEQ & ~n9582;
  assign n9584 = ~n9569 & ~n9583;
  assign n9585 = i_FULL & ~n9584;
  assign n9586 = ~i_RtoB_ACK1 & ~n9510;
  assign n9587 = ~controllable_BtoR_REQ1 & ~n9586;
  assign n9588 = ~n6788 & ~n9587;
  assign n9589 = ~controllable_BtoR_REQ0 & ~n9588;
  assign n9590 = ~controllable_BtoR_REQ0 & ~n9589;
  assign n9591 = ~i_RtoB_ACK0 & ~n9590;
  assign n9592 = ~i_RtoB_ACK0 & ~n9591;
  assign n9593 = controllable_DEQ & ~n9592;
  assign n9594 = ~n7890 & ~n9287;
  assign n9595 = ~controllable_BtoS_ACK14 & ~n9594;
  assign n9596 = ~n8215 & ~n9595;
  assign n9597 = ~controllable_ENQ & ~n9596;
  assign n9598 = ~n9498 & ~n9597;
  assign n9599 = ~i_RtoB_ACK1 & ~n9598;
  assign n9600 = ~n6773 & ~n9599;
  assign n9601 = ~controllable_BtoR_REQ1 & ~n9600;
  assign n9602 = ~n9306 & ~n9601;
  assign n9603 = ~controllable_BtoR_REQ0 & ~n9602;
  assign n9604 = ~controllable_BtoR_REQ0 & ~n9603;
  assign n9605 = ~i_RtoB_ACK0 & ~n9604;
  assign n9606 = ~n9299 & ~n9605;
  assign n9607 = ~controllable_DEQ & ~n9606;
  assign n9608 = ~n9593 & ~n9607;
  assign n9609 = ~i_FULL & ~n9608;
  assign n9610 = ~n9585 & ~n9609;
  assign n9611 = ~i_nEMPTY & ~n9610;
  assign n9612 = ~n9559 & ~n9611;
  assign n9613 = controllable_BtoS_ACK0 & ~n9612;
  assign n9614 = ~n8058 & ~n9282;
  assign n9615 = ~i_StoB_REQ14 & ~n9614;
  assign n9616 = ~n8048 & ~n9615;
  assign n9617 = controllable_BtoS_ACK14 & ~n9616;
  assign n9618 = i_StoB_REQ14 & ~n7070;
  assign n9619 = ~n9615 & ~n9618;
  assign n9620 = ~controllable_BtoS_ACK14 & ~n9619;
  assign n9621 = ~n9617 & ~n9620;
  assign n9622 = controllable_ENQ & ~n9621;
  assign n9623 = controllable_ENQ & ~n9622;
  assign n9624 = ~i_RtoB_ACK1 & ~n9623;
  assign n9625 = ~n6939 & ~n9624;
  assign n9626 = ~controllable_BtoR_REQ1 & ~n9625;
  assign n9627 = ~n6912 & ~n9626;
  assign n9628 = ~controllable_BtoR_REQ0 & ~n9627;
  assign n9629 = ~controllable_BtoR_REQ0 & ~n9628;
  assign n9630 = i_RtoB_ACK0 & ~n9629;
  assign n9631 = ~n8048 & ~n8075;
  assign n9632 = controllable_BtoS_ACK14 & ~n9631;
  assign n9633 = ~controllable_BtoS_ACK14 & ~n7070;
  assign n9634 = ~n9632 & ~n9633;
  assign n9635 = controllable_ENQ & ~n9634;
  assign n9636 = ~n6931 & ~n9635;
  assign n9637 = i_RtoB_ACK1 & ~n9636;
  assign n9638 = ~n6936 & ~n9637;
  assign n9639 = controllable_BtoR_REQ1 & ~n9638;
  assign n9640 = ~i_StoB_REQ14 & ~n9490;
  assign n9641 = ~n5108 & ~n9640;
  assign n9642 = controllable_BtoS_ACK14 & ~n9641;
  assign n9643 = ~controllable_BtoS_ACK14 & ~n9490;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = controllable_ENQ & ~n9644;
  assign n9646 = ~controllable_ENQ & ~n9621;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = ~i_RtoB_ACK1 & ~n9647;
  assign n9649 = ~n6939 & ~n9648;
  assign n9650 = ~controllable_BtoR_REQ1 & ~n9649;
  assign n9651 = ~n9639 & ~n9650;
  assign n9652 = ~controllable_BtoR_REQ0 & ~n9651;
  assign n9653 = ~controllable_BtoR_REQ0 & ~n9652;
  assign n9654 = ~i_RtoB_ACK0 & ~n9653;
  assign n9655 = ~n9630 & ~n9654;
  assign n9656 = controllable_DEQ & ~n9655;
  assign n9657 = ~i_RtoB_ACK1 & ~n9621;
  assign n9658 = ~n6961 & ~n9657;
  assign n9659 = ~controllable_BtoR_REQ1 & ~n9658;
  assign n9660 = ~n6954 & ~n9659;
  assign n9661 = ~controllable_BtoR_REQ0 & ~n9660;
  assign n9662 = ~controllable_BtoR_REQ0 & ~n9661;
  assign n9663 = i_RtoB_ACK0 & ~n9662;
  assign n9664 = i_RtoB_ACK1 & ~n9634;
  assign n9665 = ~n6962 & ~n9664;
  assign n9666 = controllable_BtoR_REQ1 & ~n9665;
  assign n9667 = ~i_RtoB_ACK1 & ~n9644;
  assign n9668 = ~n6961 & ~n9667;
  assign n9669 = ~controllable_BtoR_REQ1 & ~n9668;
  assign n9670 = ~n9666 & ~n9669;
  assign n9671 = ~controllable_BtoR_REQ0 & ~n9670;
  assign n9672 = ~controllable_BtoR_REQ0 & ~n9671;
  assign n9673 = ~i_RtoB_ACK0 & ~n9672;
  assign n9674 = ~n9663 & ~n9673;
  assign n9675 = ~controllable_DEQ & ~n9674;
  assign n9676 = ~n9656 & ~n9675;
  assign n9677 = i_FULL & ~n9676;
  assign n9678 = ~n6976 & ~n9637;
  assign n9679 = controllable_BtoR_REQ1 & ~n9678;
  assign n9680 = ~n9635 & ~n9646;
  assign n9681 = ~i_RtoB_ACK1 & ~n9680;
  assign n9682 = ~n6939 & ~n9681;
  assign n9683 = ~controllable_BtoR_REQ1 & ~n9682;
  assign n9684 = ~n9679 & ~n9683;
  assign n9685 = ~controllable_BtoR_REQ0 & ~n9684;
  assign n9686 = ~controllable_BtoR_REQ0 & ~n9685;
  assign n9687 = ~i_RtoB_ACK0 & ~n9686;
  assign n9688 = ~n9630 & ~n9687;
  assign n9689 = controllable_DEQ & ~n9688;
  assign n9690 = ~n6942 & ~n9664;
  assign n9691 = controllable_BtoR_REQ1 & ~n9690;
  assign n9692 = ~controllable_ENQ & ~n9634;
  assign n9693 = ~n9645 & ~n9692;
  assign n9694 = ~i_RtoB_ACK1 & ~n9693;
  assign n9695 = ~n6961 & ~n9694;
  assign n9696 = ~controllable_BtoR_REQ1 & ~n9695;
  assign n9697 = ~n9691 & ~n9696;
  assign n9698 = ~controllable_BtoR_REQ0 & ~n9697;
  assign n9699 = ~controllable_BtoR_REQ0 & ~n9698;
  assign n9700 = ~i_RtoB_ACK0 & ~n9699;
  assign n9701 = ~n9663 & ~n9700;
  assign n9702 = ~controllable_DEQ & ~n9701;
  assign n9703 = ~n9689 & ~n9702;
  assign n9704 = ~i_FULL & ~n9703;
  assign n9705 = ~n9677 & ~n9704;
  assign n9706 = i_nEMPTY & ~n9705;
  assign n9707 = ~controllable_ENQ & ~n9646;
  assign n9708 = ~i_RtoB_ACK1 & ~n9707;
  assign n9709 = ~i_RtoB_ACK1 & ~n9708;
  assign n9710 = ~controllable_BtoR_REQ1 & ~n9709;
  assign n9711 = ~n7006 & ~n9710;
  assign n9712 = ~controllable_BtoR_REQ0 & ~n9711;
  assign n9713 = ~controllable_BtoR_REQ0 & ~n9712;
  assign n9714 = ~i_RtoB_ACK0 & ~n9713;
  assign n9715 = ~i_RtoB_ACK0 & ~n9714;
  assign n9716 = controllable_DEQ & ~n9715;
  assign n9717 = controllable_ENQ & ~n9635;
  assign n9718 = i_RtoB_ACK1 & ~n9717;
  assign n9719 = ~n7019 & ~n9718;
  assign n9720 = controllable_BtoR_REQ1 & ~n9719;
  assign n9721 = controllable_ENQ & ~n9645;
  assign n9722 = ~i_RtoB_ACK1 & ~n9721;
  assign n9723 = ~n6939 & ~n9722;
  assign n9724 = ~controllable_BtoR_REQ1 & ~n9723;
  assign n9725 = ~n9720 & ~n9724;
  assign n9726 = ~controllable_BtoR_REQ0 & ~n9725;
  assign n9727 = ~controllable_BtoR_REQ0 & ~n9726;
  assign n9728 = ~i_RtoB_ACK0 & ~n9727;
  assign n9729 = ~n9630 & ~n9728;
  assign n9730 = ~controllable_DEQ & ~n9729;
  assign n9731 = ~n9716 & ~n9730;
  assign n9732 = i_FULL & ~n9731;
  assign n9733 = ~i_RtoB_ACK1 & ~n9657;
  assign n9734 = ~controllable_BtoR_REQ1 & ~n9733;
  assign n9735 = ~n6954 & ~n9734;
  assign n9736 = ~controllable_BtoR_REQ0 & ~n9735;
  assign n9737 = ~controllable_BtoR_REQ0 & ~n9736;
  assign n9738 = ~i_RtoB_ACK0 & ~n9737;
  assign n9739 = ~i_RtoB_ACK0 & ~n9738;
  assign n9740 = controllable_DEQ & ~n9739;
  assign n9741 = i_StoB_REQ14 & ~n7781;
  assign n9742 = ~n8060 & ~n9741;
  assign n9743 = controllable_BtoS_ACK14 & ~n9742;
  assign n9744 = ~n8060 & ~n9618;
  assign n9745 = ~controllable_BtoS_ACK14 & ~n9744;
  assign n9746 = ~n9743 & ~n9745;
  assign n9747 = ~controllable_ENQ & ~n9746;
  assign n9748 = ~n9645 & ~n9747;
  assign n9749 = ~i_RtoB_ACK1 & ~n9748;
  assign n9750 = ~n6939 & ~n9749;
  assign n9751 = ~controllable_BtoR_REQ1 & ~n9750;
  assign n9752 = ~n9639 & ~n9751;
  assign n9753 = ~controllable_BtoR_REQ0 & ~n9752;
  assign n9754 = ~controllable_BtoR_REQ0 & ~n9753;
  assign n9755 = ~i_RtoB_ACK0 & ~n9754;
  assign n9756 = ~n9630 & ~n9755;
  assign n9757 = ~controllable_DEQ & ~n9756;
  assign n9758 = ~n9740 & ~n9757;
  assign n9759 = ~i_FULL & ~n9758;
  assign n9760 = ~n9732 & ~n9759;
  assign n9761 = ~i_nEMPTY & ~n9760;
  assign n9762 = ~n9706 & ~n9761;
  assign n9763 = ~controllable_BtoS_ACK0 & ~n9762;
  assign n9764 = ~n9613 & ~n9763;
  assign n9765 = n4465 & ~n9764;
  assign n9766 = ~i_StoB_REQ13 & ~n9275;
  assign n9767 = ~n5204 & ~n9766;
  assign n9768 = n4466 & ~n9767;
  assign n9769 = ~n4466 & ~n5213;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = i_StoB_REQ0 & ~n9770;
  assign n9772 = ~n7071 & ~n9771;
  assign n9773 = ~i_StoB_REQ14 & ~n9772;
  assign n9774 = ~n5216 & ~n9773;
  assign n9775 = controllable_BtoS_ACK14 & ~n9774;
  assign n9776 = ~n9287 & ~n9773;
  assign n9777 = ~controllable_BtoS_ACK14 & ~n9776;
  assign n9778 = ~n9775 & ~n9777;
  assign n9779 = controllable_ENQ & ~n9778;
  assign n9780 = controllable_ENQ & ~n9779;
  assign n9781 = ~i_RtoB_ACK1 & ~n9780;
  assign n9782 = ~n7101 & ~n9781;
  assign n9783 = ~controllable_BtoR_REQ1 & ~n9782;
  assign n9784 = ~n7081 & ~n9783;
  assign n9785 = ~controllable_BtoR_REQ0 & ~n9784;
  assign n9786 = ~controllable_BtoR_REQ0 & ~n9785;
  assign n9787 = i_RtoB_ACK0 & ~n9786;
  assign n9788 = ~n5238 & ~n9302;
  assign n9789 = i_RtoB_ACK1 & ~n9788;
  assign n9790 = ~n7098 & ~n9789;
  assign n9791 = controllable_BtoR_REQ1 & ~n9790;
  assign n9792 = ~controllable_ENQ & ~n9778;
  assign n9793 = ~n9302 & ~n9792;
  assign n9794 = ~i_RtoB_ACK1 & ~n9793;
  assign n9795 = ~n7101 & ~n9794;
  assign n9796 = ~controllable_BtoR_REQ1 & ~n9795;
  assign n9797 = ~n9791 & ~n9796;
  assign n9798 = ~controllable_BtoR_REQ0 & ~n9797;
  assign n9799 = ~controllable_BtoR_REQ0 & ~n9798;
  assign n9800 = ~i_RtoB_ACK0 & ~n9799;
  assign n9801 = ~n9787 & ~n9800;
  assign n9802 = controllable_DEQ & ~n9801;
  assign n9803 = i_RtoB_ACK1 & ~n7086;
  assign n9804 = ~i_RtoB_ACK1 & ~n9778;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~controllable_BtoR_REQ1 & ~n9805;
  assign n9807 = ~n7114 & ~n9806;
  assign n9808 = ~controllable_BtoR_REQ0 & ~n9807;
  assign n9809 = ~controllable_BtoR_REQ0 & ~n9808;
  assign n9810 = i_RtoB_ACK0 & ~n9809;
  assign n9811 = ~n7102 & ~n9517;
  assign n9812 = controllable_BtoR_REQ1 & ~n9811;
  assign n9813 = ~i_RtoB_ACK1 & ~n9301;
  assign n9814 = ~n9803 & ~n9813;
  assign n9815 = ~controllable_BtoR_REQ1 & ~n9814;
  assign n9816 = ~n9812 & ~n9815;
  assign n9817 = ~controllable_BtoR_REQ0 & ~n9816;
  assign n9818 = ~controllable_BtoR_REQ0 & ~n9817;
  assign n9819 = ~i_RtoB_ACK0 & ~n9818;
  assign n9820 = ~n9810 & ~n9819;
  assign n9821 = ~controllable_DEQ & ~n9820;
  assign n9822 = ~n9802 & ~n9821;
  assign n9823 = i_nEMPTY & ~n9822;
  assign n9824 = ~controllable_ENQ & ~n9792;
  assign n9825 = ~i_RtoB_ACK1 & ~n9824;
  assign n9826 = ~i_RtoB_ACK1 & ~n9825;
  assign n9827 = ~controllable_BtoR_REQ1 & ~n9826;
  assign n9828 = ~n7131 & ~n9827;
  assign n9829 = ~controllable_BtoR_REQ0 & ~n9828;
  assign n9830 = ~controllable_BtoR_REQ0 & ~n9829;
  assign n9831 = ~i_RtoB_ACK0 & ~n9830;
  assign n9832 = ~i_RtoB_ACK0 & ~n9831;
  assign n9833 = controllable_DEQ & ~n9832;
  assign n9834 = ~n7546 & ~n9571;
  assign n9835 = controllable_BtoR_REQ1 & ~n9834;
  assign n9836 = ~i_RtoB_ACK1 & ~n9570;
  assign n9837 = ~n7101 & ~n9836;
  assign n9838 = ~controllable_BtoR_REQ1 & ~n9837;
  assign n9839 = ~n9835 & ~n9838;
  assign n9840 = ~controllable_BtoR_REQ0 & ~n9839;
  assign n9841 = ~controllable_BtoR_REQ0 & ~n9840;
  assign n9842 = ~i_RtoB_ACK0 & ~n9841;
  assign n9843 = ~n9787 & ~n9842;
  assign n9844 = ~controllable_DEQ & ~n9843;
  assign n9845 = ~n9833 & ~n9844;
  assign n9846 = i_FULL & ~n9845;
  assign n9847 = ~i_RtoB_ACK1 & ~n9804;
  assign n9848 = ~controllable_BtoR_REQ1 & ~n9847;
  assign n9849 = ~n7114 & ~n9848;
  assign n9850 = ~controllable_BtoR_REQ0 & ~n9849;
  assign n9851 = ~controllable_BtoR_REQ0 & ~n9850;
  assign n9852 = ~i_RtoB_ACK0 & ~n9851;
  assign n9853 = ~i_RtoB_ACK0 & ~n9852;
  assign n9854 = controllable_DEQ & ~n9853;
  assign n9855 = ~n9302 & ~n9597;
  assign n9856 = ~i_RtoB_ACK1 & ~n9855;
  assign n9857 = ~n7101 & ~n9856;
  assign n9858 = ~controllable_BtoR_REQ1 & ~n9857;
  assign n9859 = ~n9791 & ~n9858;
  assign n9860 = ~controllable_BtoR_REQ0 & ~n9859;
  assign n9861 = ~controllable_BtoR_REQ0 & ~n9860;
  assign n9862 = ~i_RtoB_ACK0 & ~n9861;
  assign n9863 = ~n9787 & ~n9862;
  assign n9864 = ~controllable_DEQ & ~n9863;
  assign n9865 = ~n9854 & ~n9864;
  assign n9866 = ~i_FULL & ~n9865;
  assign n9867 = ~n9846 & ~n9866;
  assign n9868 = ~i_nEMPTY & ~n9867;
  assign n9869 = ~n9823 & ~n9868;
  assign n9870 = controllable_BtoS_ACK0 & ~n9869;
  assign n9871 = ~i_RtoB_ACK1 & ~n9717;
  assign n9872 = ~n7265 & ~n9871;
  assign n9873 = ~controllable_BtoR_REQ1 & ~n9872;
  assign n9874 = ~n7234 & ~n9873;
  assign n9875 = ~controllable_BtoR_REQ0 & ~n9874;
  assign n9876 = ~controllable_BtoR_REQ0 & ~n9875;
  assign n9877 = i_RtoB_ACK0 & ~n9876;
  assign n9878 = ~n7257 & ~n9635;
  assign n9879 = i_RtoB_ACK1 & ~n9878;
  assign n9880 = ~n7262 & ~n9879;
  assign n9881 = controllable_BtoR_REQ1 & ~n9880;
  assign n9882 = ~n6540 & ~n9483;
  assign n9883 = i_StoB_REQ13 & ~n9882;
  assign n9884 = ~i_StoB_REQ13 & ~n9482;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = n4466 & ~n9885;
  assign n9887 = ~n9489 & ~n9886;
  assign n9888 = ~i_StoB_REQ14 & ~n9887;
  assign n9889 = ~n5322 & ~n9888;
  assign n9890 = controllable_BtoS_ACK14 & ~n9889;
  assign n9891 = ~controllable_BtoS_ACK14 & ~n9887;
  assign n9892 = ~n9890 & ~n9891;
  assign n9893 = controllable_ENQ & ~n9892;
  assign n9894 = ~n9692 & ~n9893;
  assign n9895 = ~i_RtoB_ACK1 & ~n9894;
  assign n9896 = ~n7265 & ~n9895;
  assign n9897 = ~controllable_BtoR_REQ1 & ~n9896;
  assign n9898 = ~n9881 & ~n9897;
  assign n9899 = ~controllable_BtoR_REQ0 & ~n9898;
  assign n9900 = ~controllable_BtoR_REQ0 & ~n9899;
  assign n9901 = ~i_RtoB_ACK0 & ~n9900;
  assign n9902 = ~n9877 & ~n9901;
  assign n9903 = controllable_DEQ & ~n9902;
  assign n9904 = ~i_RtoB_ACK1 & ~n9634;
  assign n9905 = ~n7287 & ~n9904;
  assign n9906 = ~controllable_BtoR_REQ1 & ~n9905;
  assign n9907 = ~n7280 & ~n9906;
  assign n9908 = ~controllable_BtoR_REQ0 & ~n9907;
  assign n9909 = ~controllable_BtoR_REQ0 & ~n9908;
  assign n9910 = i_RtoB_ACK0 & ~n9909;
  assign n9911 = ~n7288 & ~n9664;
  assign n9912 = controllable_BtoR_REQ1 & ~n9911;
  assign n9913 = ~i_RtoB_ACK1 & ~n9892;
  assign n9914 = ~n7287 & ~n9913;
  assign n9915 = ~controllable_BtoR_REQ1 & ~n9914;
  assign n9916 = ~n9912 & ~n9915;
  assign n9917 = ~controllable_BtoR_REQ0 & ~n9916;
  assign n9918 = ~controllable_BtoR_REQ0 & ~n9917;
  assign n9919 = ~i_RtoB_ACK0 & ~n9918;
  assign n9920 = ~n9910 & ~n9919;
  assign n9921 = ~controllable_DEQ & ~n9920;
  assign n9922 = ~n9903 & ~n9921;
  assign n9923 = i_FULL & ~n9922;
  assign n9924 = ~n7302 & ~n9879;
  assign n9925 = controllable_BtoR_REQ1 & ~n9924;
  assign n9926 = ~n7265 & ~n9904;
  assign n9927 = ~controllable_BtoR_REQ1 & ~n9926;
  assign n9928 = ~n9925 & ~n9927;
  assign n9929 = ~controllable_BtoR_REQ0 & ~n9928;
  assign n9930 = ~controllable_BtoR_REQ0 & ~n9929;
  assign n9931 = ~i_RtoB_ACK0 & ~n9930;
  assign n9932 = ~n9877 & ~n9931;
  assign n9933 = controllable_DEQ & ~n9932;
  assign n9934 = ~n7268 & ~n9664;
  assign n9935 = controllable_BtoR_REQ1 & ~n9934;
  assign n9936 = ~n7287 & ~n9895;
  assign n9937 = ~controllable_BtoR_REQ1 & ~n9936;
  assign n9938 = ~n9935 & ~n9937;
  assign n9939 = ~controllable_BtoR_REQ0 & ~n9938;
  assign n9940 = ~controllable_BtoR_REQ0 & ~n9939;
  assign n9941 = ~i_RtoB_ACK0 & ~n9940;
  assign n9942 = ~n9910 & ~n9941;
  assign n9943 = ~controllable_DEQ & ~n9942;
  assign n9944 = ~n9933 & ~n9943;
  assign n9945 = ~i_FULL & ~n9944;
  assign n9946 = ~n9923 & ~n9945;
  assign n9947 = i_nEMPTY & ~n9946;
  assign n9948 = ~controllable_ENQ & ~n9692;
  assign n9949 = ~i_RtoB_ACK1 & ~n9948;
  assign n9950 = ~i_RtoB_ACK1 & ~n9949;
  assign n9951 = ~controllable_BtoR_REQ1 & ~n9950;
  assign n9952 = ~n7332 & ~n9951;
  assign n9953 = ~controllable_BtoR_REQ0 & ~n9952;
  assign n9954 = ~controllable_BtoR_REQ0 & ~n9953;
  assign n9955 = ~i_RtoB_ACK0 & ~n9954;
  assign n9956 = ~i_RtoB_ACK0 & ~n9955;
  assign n9957 = controllable_DEQ & ~n9956;
  assign n9958 = ~n7345 & ~n9718;
  assign n9959 = controllable_BtoR_REQ1 & ~n9958;
  assign n9960 = controllable_ENQ & ~n9893;
  assign n9961 = ~i_RtoB_ACK1 & ~n9960;
  assign n9962 = ~n7265 & ~n9961;
  assign n9963 = ~controllable_BtoR_REQ1 & ~n9962;
  assign n9964 = ~n9959 & ~n9963;
  assign n9965 = ~controllable_BtoR_REQ0 & ~n9964;
  assign n9966 = ~controllable_BtoR_REQ0 & ~n9965;
  assign n9967 = ~i_RtoB_ACK0 & ~n9966;
  assign n9968 = ~n9877 & ~n9967;
  assign n9969 = ~controllable_DEQ & ~n9968;
  assign n9970 = ~n9957 & ~n9969;
  assign n9971 = i_FULL & ~n9970;
  assign n9972 = ~i_RtoB_ACK1 & ~n9904;
  assign n9973 = ~controllable_BtoR_REQ1 & ~n9972;
  assign n9974 = ~n7280 & ~n9973;
  assign n9975 = ~controllable_BtoR_REQ0 & ~n9974;
  assign n9976 = ~controllable_BtoR_REQ0 & ~n9975;
  assign n9977 = ~i_RtoB_ACK0 & ~n9976;
  assign n9978 = ~i_RtoB_ACK0 & ~n9977;
  assign n9979 = controllable_DEQ & ~n9978;
  assign n9980 = ~n9747 & ~n9893;
  assign n9981 = ~i_RtoB_ACK1 & ~n9980;
  assign n9982 = ~n7265 & ~n9981;
  assign n9983 = ~controllable_BtoR_REQ1 & ~n9982;
  assign n9984 = ~n9881 & ~n9983;
  assign n9985 = ~controllable_BtoR_REQ0 & ~n9984;
  assign n9986 = ~controllable_BtoR_REQ0 & ~n9985;
  assign n9987 = ~i_RtoB_ACK0 & ~n9986;
  assign n9988 = ~n9877 & ~n9987;
  assign n9989 = ~controllable_DEQ & ~n9988;
  assign n9990 = ~n9979 & ~n9989;
  assign n9991 = ~i_FULL & ~n9990;
  assign n9992 = ~n9971 & ~n9991;
  assign n9993 = ~i_nEMPTY & ~n9992;
  assign n9994 = ~n9947 & ~n9993;
  assign n9995 = ~controllable_BtoS_ACK0 & ~n9994;
  assign n9996 = ~n9870 & ~n9995;
  assign n9997 = ~n4465 & ~n9996;
  assign n9998 = ~n9765 & ~n9997;
  assign n9999 = ~i_StoB_REQ10 & ~n9998;
  assign n10000 = ~n9062 & ~n9999;
  assign n10001 = controllable_BtoS_ACK10 & ~n10000;
  assign n10002 = ~n6773 & ~n9836;
  assign n10003 = ~controllable_BtoR_REQ1 & ~n10002;
  assign n10004 = ~n7394 & ~n10003;
  assign n10005 = ~controllable_BtoR_REQ0 & ~n10004;
  assign n10006 = ~controllable_BtoR_REQ0 & ~n10005;
  assign n10007 = i_RtoB_ACK0 & ~n10006;
  assign n10008 = ~n7399 & ~n9302;
  assign n10009 = i_RtoB_ACK1 & ~n10008;
  assign n10010 = ~n6776 & ~n10009;
  assign n10011 = controllable_BtoR_REQ1 & ~n10010;
  assign n10012 = ~n6773 & ~n9547;
  assign n10013 = ~controllable_BtoR_REQ1 & ~n10012;
  assign n10014 = ~n10011 & ~n10013;
  assign n10015 = ~controllable_BtoR_REQ0 & ~n10014;
  assign n10016 = ~controllable_BtoR_REQ0 & ~n10015;
  assign n10017 = ~i_RtoB_ACK0 & ~n10016;
  assign n10018 = ~n10007 & ~n10017;
  assign n10019 = controllable_DEQ & ~n10018;
  assign n10020 = ~n6795 & ~n9813;
  assign n10021 = ~controllable_BtoR_REQ1 & ~n10020;
  assign n10022 = ~n7412 & ~n10021;
  assign n10023 = ~controllable_BtoR_REQ0 & ~n10022;
  assign n10024 = ~controllable_BtoR_REQ0 & ~n10023;
  assign n10025 = i_RtoB_ACK0 & ~n10024;
  assign n10026 = ~n9526 & ~n10025;
  assign n10027 = ~controllable_DEQ & ~n10026;
  assign n10028 = ~n10019 & ~n10027;
  assign n10029 = i_FULL & ~n10028;
  assign n10030 = ~n6813 & ~n10009;
  assign n10031 = controllable_BtoR_REQ1 & ~n10030;
  assign n10032 = ~n6773 & ~n9813;
  assign n10033 = ~controllable_BtoR_REQ1 & ~n10032;
  assign n10034 = ~n10031 & ~n10033;
  assign n10035 = ~controllable_BtoR_REQ0 & ~n10034;
  assign n10036 = ~controllable_BtoR_REQ0 & ~n10035;
  assign n10037 = ~i_RtoB_ACK0 & ~n10036;
  assign n10038 = ~n10007 & ~n10037;
  assign n10039 = controllable_DEQ & ~n10038;
  assign n10040 = ~n9553 & ~n10025;
  assign n10041 = ~controllable_DEQ & ~n10040;
  assign n10042 = ~n10039 & ~n10041;
  assign n10043 = ~i_FULL & ~n10042;
  assign n10044 = ~n10029 & ~n10043;
  assign n10045 = i_nEMPTY & ~n10044;
  assign n10046 = ~controllable_ENQ & ~n9545;
  assign n10047 = ~i_RtoB_ACK1 & ~n10046;
  assign n10048 = ~i_RtoB_ACK1 & ~n10047;
  assign n10049 = ~controllable_BtoR_REQ1 & ~n10048;
  assign n10050 = ~n7440 & ~n10049;
  assign n10051 = ~controllable_BtoR_REQ0 & ~n10050;
  assign n10052 = ~controllable_BtoR_REQ0 & ~n10051;
  assign n10053 = ~i_RtoB_ACK0 & ~n10052;
  assign n10054 = ~i_RtoB_ACK0 & ~n10053;
  assign n10055 = controllable_DEQ & ~n10054;
  assign n10056 = ~n9581 & ~n10007;
  assign n10057 = ~controllable_DEQ & ~n10056;
  assign n10058 = ~n10055 & ~n10057;
  assign n10059 = i_FULL & ~n10058;
  assign n10060 = ~i_RtoB_ACK1 & ~n9813;
  assign n10061 = ~controllable_BtoR_REQ1 & ~n10060;
  assign n10062 = ~n7412 & ~n10061;
  assign n10063 = ~controllable_BtoR_REQ0 & ~n10062;
  assign n10064 = ~controllable_BtoR_REQ0 & ~n10063;
  assign n10065 = ~i_RtoB_ACK0 & ~n10064;
  assign n10066 = ~i_RtoB_ACK0 & ~n10065;
  assign n10067 = controllable_DEQ & ~n10066;
  assign n10068 = ~controllable_DEQ & ~n10018;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = ~i_FULL & ~n10069;
  assign n10071 = ~n10059 & ~n10070;
  assign n10072 = ~i_nEMPTY & ~n10071;
  assign n10073 = ~n10045 & ~n10072;
  assign n10074 = controllable_BtoS_ACK0 & ~n10073;
  assign n10075 = ~n6939 & ~n9871;
  assign n10076 = ~controllable_BtoR_REQ1 & ~n10075;
  assign n10077 = ~n7474 & ~n10076;
  assign n10078 = ~controllable_BtoR_REQ0 & ~n10077;
  assign n10079 = ~controllable_BtoR_REQ0 & ~n10078;
  assign n10080 = i_RtoB_ACK0 & ~n10079;
  assign n10081 = ~n7479 & ~n9635;
  assign n10082 = i_RtoB_ACK1 & ~n10081;
  assign n10083 = ~n6942 & ~n10082;
  assign n10084 = controllable_BtoR_REQ1 & ~n10083;
  assign n10085 = ~n6939 & ~n9694;
  assign n10086 = ~controllable_BtoR_REQ1 & ~n10085;
  assign n10087 = ~n10084 & ~n10086;
  assign n10088 = ~controllable_BtoR_REQ0 & ~n10087;
  assign n10089 = ~controllable_BtoR_REQ0 & ~n10088;
  assign n10090 = ~i_RtoB_ACK0 & ~n10089;
  assign n10091 = ~n10080 & ~n10090;
  assign n10092 = controllable_DEQ & ~n10091;
  assign n10093 = ~n6961 & ~n9904;
  assign n10094 = ~controllable_BtoR_REQ1 & ~n10093;
  assign n10095 = ~n7492 & ~n10094;
  assign n10096 = ~controllable_BtoR_REQ0 & ~n10095;
  assign n10097 = ~controllable_BtoR_REQ0 & ~n10096;
  assign n10098 = i_RtoB_ACK0 & ~n10097;
  assign n10099 = ~n9673 & ~n10098;
  assign n10100 = ~controllable_DEQ & ~n10099;
  assign n10101 = ~n10092 & ~n10100;
  assign n10102 = i_FULL & ~n10101;
  assign n10103 = ~n6979 & ~n10082;
  assign n10104 = controllable_BtoR_REQ1 & ~n10103;
  assign n10105 = ~n6939 & ~n9904;
  assign n10106 = ~controllable_BtoR_REQ1 & ~n10105;
  assign n10107 = ~n10104 & ~n10106;
  assign n10108 = ~controllable_BtoR_REQ0 & ~n10107;
  assign n10109 = ~controllable_BtoR_REQ0 & ~n10108;
  assign n10110 = ~i_RtoB_ACK0 & ~n10109;
  assign n10111 = ~n10080 & ~n10110;
  assign n10112 = controllable_DEQ & ~n10111;
  assign n10113 = ~n9700 & ~n10098;
  assign n10114 = ~controllable_DEQ & ~n10113;
  assign n10115 = ~n10112 & ~n10114;
  assign n10116 = ~i_FULL & ~n10115;
  assign n10117 = ~n10102 & ~n10116;
  assign n10118 = i_nEMPTY & ~n10117;
  assign n10119 = ~n7520 & ~n9951;
  assign n10120 = ~controllable_BtoR_REQ0 & ~n10119;
  assign n10121 = ~controllable_BtoR_REQ0 & ~n10120;
  assign n10122 = ~i_RtoB_ACK0 & ~n10121;
  assign n10123 = ~i_RtoB_ACK0 & ~n10122;
  assign n10124 = controllable_DEQ & ~n10123;
  assign n10125 = ~n9728 & ~n10080;
  assign n10126 = ~controllable_DEQ & ~n10125;
  assign n10127 = ~n10124 & ~n10126;
  assign n10128 = i_FULL & ~n10127;
  assign n10129 = ~n7492 & ~n9973;
  assign n10130 = ~controllable_BtoR_REQ0 & ~n10129;
  assign n10131 = ~controllable_BtoR_REQ0 & ~n10130;
  assign n10132 = ~i_RtoB_ACK0 & ~n10131;
  assign n10133 = ~i_RtoB_ACK0 & ~n10132;
  assign n10134 = controllable_DEQ & ~n10133;
  assign n10135 = ~controllable_DEQ & ~n10091;
  assign n10136 = ~n10134 & ~n10135;
  assign n10137 = ~i_FULL & ~n10136;
  assign n10138 = ~n10128 & ~n10137;
  assign n10139 = ~i_nEMPTY & ~n10138;
  assign n10140 = ~n10118 & ~n10139;
  assign n10141 = ~controllable_BtoS_ACK0 & ~n10140;
  assign n10142 = ~n10074 & ~n10141;
  assign n10143 = n4465 & ~n10142;
  assign n10144 = ~n7548 & ~n9838;
  assign n10145 = ~controllable_BtoR_REQ0 & ~n10144;
  assign n10146 = ~controllable_BtoR_REQ0 & ~n10145;
  assign n10147 = i_RtoB_ACK0 & ~n10146;
  assign n10148 = ~n5271 & ~n9302;
  assign n10149 = i_RtoB_ACK1 & ~n10148;
  assign n10150 = ~n7102 & ~n10149;
  assign n10151 = controllable_BtoR_REQ1 & ~n10150;
  assign n10152 = ~n7101 & ~n9813;
  assign n10153 = ~controllable_BtoR_REQ1 & ~n10152;
  assign n10154 = ~n10151 & ~n10153;
  assign n10155 = ~controllable_BtoR_REQ0 & ~n10154;
  assign n10156 = ~controllable_BtoR_REQ0 & ~n10155;
  assign n10157 = ~i_RtoB_ACK0 & ~n10156;
  assign n10158 = ~n10147 & ~n10157;
  assign n10159 = controllable_DEQ & ~n10158;
  assign n10160 = ~n7565 & ~n9815;
  assign n10161 = ~controllable_BtoR_REQ0 & ~n10160;
  assign n10162 = ~controllable_BtoR_REQ0 & ~n10161;
  assign n10163 = i_RtoB_ACK0 & ~n10162;
  assign n10164 = ~n9819 & ~n10163;
  assign n10165 = ~controllable_DEQ & ~n10164;
  assign n10166 = ~n10159 & ~n10165;
  assign n10167 = i_nEMPTY & ~n10166;
  assign n10168 = ~n7576 & ~n10049;
  assign n10169 = ~controllable_BtoR_REQ0 & ~n10168;
  assign n10170 = ~controllable_BtoR_REQ0 & ~n10169;
  assign n10171 = ~i_RtoB_ACK0 & ~n10170;
  assign n10172 = ~i_RtoB_ACK0 & ~n10171;
  assign n10173 = controllable_DEQ & ~n10172;
  assign n10174 = ~n9842 & ~n10147;
  assign n10175 = ~controllable_DEQ & ~n10174;
  assign n10176 = ~n10173 & ~n10175;
  assign n10177 = i_FULL & ~n10176;
  assign n10178 = ~n7565 & ~n10061;
  assign n10179 = ~controllable_BtoR_REQ0 & ~n10178;
  assign n10180 = ~controllable_BtoR_REQ0 & ~n10179;
  assign n10181 = ~i_RtoB_ACK0 & ~n10180;
  assign n10182 = ~i_RtoB_ACK0 & ~n10181;
  assign n10183 = controllable_DEQ & ~n10182;
  assign n10184 = ~controllable_DEQ & ~n10158;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = ~i_FULL & ~n10185;
  assign n10187 = ~n10177 & ~n10186;
  assign n10188 = ~i_nEMPTY & ~n10187;
  assign n10189 = ~n10167 & ~n10188;
  assign n10190 = controllable_BtoS_ACK0 & ~n10189;
  assign n10191 = ~n7610 & ~n9873;
  assign n10192 = ~controllable_BtoR_REQ0 & ~n10191;
  assign n10193 = ~controllable_BtoR_REQ0 & ~n10192;
  assign n10194 = i_RtoB_ACK0 & ~n10193;
  assign n10195 = ~n7615 & ~n9635;
  assign n10196 = i_RtoB_ACK1 & ~n10195;
  assign n10197 = ~n7268 & ~n10196;
  assign n10198 = controllable_BtoR_REQ1 & ~n10197;
  assign n10199 = ~n9897 & ~n10198;
  assign n10200 = ~controllable_BtoR_REQ0 & ~n10199;
  assign n10201 = ~controllable_BtoR_REQ0 & ~n10200;
  assign n10202 = ~i_RtoB_ACK0 & ~n10201;
  assign n10203 = ~n10194 & ~n10202;
  assign n10204 = controllable_DEQ & ~n10203;
  assign n10205 = ~n7628 & ~n9906;
  assign n10206 = ~controllable_BtoR_REQ0 & ~n10205;
  assign n10207 = ~controllable_BtoR_REQ0 & ~n10206;
  assign n10208 = i_RtoB_ACK0 & ~n10207;
  assign n10209 = ~n9919 & ~n10208;
  assign n10210 = ~controllable_DEQ & ~n10209;
  assign n10211 = ~n10204 & ~n10210;
  assign n10212 = i_FULL & ~n10211;
  assign n10213 = ~n7305 & ~n10196;
  assign n10214 = controllable_BtoR_REQ1 & ~n10213;
  assign n10215 = ~n9927 & ~n10214;
  assign n10216 = ~controllable_BtoR_REQ0 & ~n10215;
  assign n10217 = ~controllable_BtoR_REQ0 & ~n10216;
  assign n10218 = ~i_RtoB_ACK0 & ~n10217;
  assign n10219 = ~n10194 & ~n10218;
  assign n10220 = controllable_DEQ & ~n10219;
  assign n10221 = ~n9941 & ~n10208;
  assign n10222 = ~controllable_DEQ & ~n10221;
  assign n10223 = ~n10220 & ~n10222;
  assign n10224 = ~i_FULL & ~n10223;
  assign n10225 = ~n10212 & ~n10224;
  assign n10226 = i_nEMPTY & ~n10225;
  assign n10227 = ~n7656 & ~n9951;
  assign n10228 = ~controllable_BtoR_REQ0 & ~n10227;
  assign n10229 = ~controllable_BtoR_REQ0 & ~n10228;
  assign n10230 = ~i_RtoB_ACK0 & ~n10229;
  assign n10231 = ~i_RtoB_ACK0 & ~n10230;
  assign n10232 = controllable_DEQ & ~n10231;
  assign n10233 = ~n9967 & ~n10194;
  assign n10234 = ~controllable_DEQ & ~n10233;
  assign n10235 = ~n10232 & ~n10234;
  assign n10236 = i_FULL & ~n10235;
  assign n10237 = ~n7628 & ~n9973;
  assign n10238 = ~controllable_BtoR_REQ0 & ~n10237;
  assign n10239 = ~controllable_BtoR_REQ0 & ~n10238;
  assign n10240 = ~i_RtoB_ACK0 & ~n10239;
  assign n10241 = ~i_RtoB_ACK0 & ~n10240;
  assign n10242 = controllable_DEQ & ~n10241;
  assign n10243 = ~controllable_DEQ & ~n10203;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = ~i_FULL & ~n10244;
  assign n10246 = ~n10236 & ~n10245;
  assign n10247 = ~i_nEMPTY & ~n10246;
  assign n10248 = ~n10226 & ~n10247;
  assign n10249 = ~controllable_BtoS_ACK0 & ~n10248;
  assign n10250 = ~n10190 & ~n10249;
  assign n10251 = ~n4465 & ~n10250;
  assign n10252 = ~n10143 & ~n10251;
  assign n10253 = i_StoB_REQ10 & ~n10252;
  assign n10254 = ~n9999 & ~n10253;
  assign n10255 = ~controllable_BtoS_ACK10 & ~n10254;
  assign n10256 = ~n10001 & ~n10255;
  assign n10257 = n4464 & ~n10256;
  assign n10258 = ~n7710 & ~n8755;
  assign n10259 = ~controllable_BtoR_REQ1 & ~n10258;
  assign n10260 = ~n7700 & ~n10259;
  assign n10261 = ~controllable_BtoR_REQ0 & ~n10260;
  assign n10262 = ~controllable_BtoR_REQ0 & ~n10261;
  assign n10263 = i_RtoB_ACK0 & ~n10262;
  assign n10264 = ~n5237 & ~n7713;
  assign n10265 = controllable_BtoR_REQ1 & ~n10264;
  assign n10266 = ~n5271 & ~n7703;
  assign n10267 = ~i_RtoB_ACK1 & ~n10266;
  assign n10268 = ~n7710 & ~n10267;
  assign n10269 = ~controllable_BtoR_REQ1 & ~n10268;
  assign n10270 = ~n10265 & ~n10269;
  assign n10271 = ~controllable_BtoR_REQ0 & ~n10270;
  assign n10272 = ~controllable_BtoR_REQ0 & ~n10271;
  assign n10273 = ~i_RtoB_ACK0 & ~n10272;
  assign n10274 = ~n10263 & ~n10273;
  assign n10275 = controllable_DEQ & ~n10274;
  assign n10276 = i_RtoB_ACK1 & ~n7702;
  assign n10277 = ~n5243 & ~n10276;
  assign n10278 = ~controllable_BtoR_REQ1 & ~n10277;
  assign n10279 = ~n7727 & ~n10278;
  assign n10280 = ~controllable_BtoR_REQ0 & ~n10279;
  assign n10281 = ~controllable_BtoR_REQ0 & ~n10280;
  assign n10282 = i_RtoB_ACK0 & ~n10281;
  assign n10283 = ~n7563 & ~n7716;
  assign n10284 = controllable_BtoR_REQ1 & ~n10283;
  assign n10285 = ~n7728 & ~n10284;
  assign n10286 = ~controllable_BtoR_REQ0 & ~n10285;
  assign n10287 = ~controllable_BtoR_REQ0 & ~n10286;
  assign n10288 = ~i_RtoB_ACK0 & ~n10287;
  assign n10289 = ~n10282 & ~n10288;
  assign n10290 = ~controllable_DEQ & ~n10289;
  assign n10291 = ~n10275 & ~n10290;
  assign n10292 = i_FULL & ~n10291;
  assign n10293 = ~n5243 & ~n7710;
  assign n10294 = ~controllable_BtoR_REQ1 & ~n10293;
  assign n10295 = ~n10265 & ~n10294;
  assign n10296 = ~controllable_BtoR_REQ0 & ~n10295;
  assign n10297 = ~controllable_BtoR_REQ0 & ~n10296;
  assign n10298 = ~i_RtoB_ACK0 & ~n10297;
  assign n10299 = ~n10263 & ~n10298;
  assign n10300 = controllable_DEQ & ~n10299;
  assign n10301 = ~n10267 & ~n10276;
  assign n10302 = ~controllable_BtoR_REQ1 & ~n10301;
  assign n10303 = ~n10284 & ~n10302;
  assign n10304 = ~controllable_BtoR_REQ0 & ~n10303;
  assign n10305 = ~controllable_BtoR_REQ0 & ~n10304;
  assign n10306 = ~i_RtoB_ACK0 & ~n10305;
  assign n10307 = ~n10282 & ~n10306;
  assign n10308 = ~controllable_DEQ & ~n10307;
  assign n10309 = ~n10300 & ~n10308;
  assign n10310 = ~i_FULL & ~n10309;
  assign n10311 = ~n10292 & ~n10310;
  assign n10312 = i_nEMPTY & ~n10311;
  assign n10313 = ~n5275 & ~n7743;
  assign n10314 = ~controllable_BtoR_REQ0 & ~n10313;
  assign n10315 = ~controllable_BtoR_REQ0 & ~n10314;
  assign n10316 = ~i_RtoB_ACK0 & ~n10315;
  assign n10317 = ~i_RtoB_ACK0 & ~n10316;
  assign n10318 = controllable_DEQ & ~n10317;
  assign n10319 = ~i_RtoB_ACK1 & ~n7704;
  assign n10320 = ~n5237 & ~n10319;
  assign n10321 = controllable_BtoR_REQ1 & ~n10320;
  assign n10322 = ~n7705 & ~n10321;
  assign n10323 = ~controllable_BtoR_REQ0 & ~n10322;
  assign n10324 = ~controllable_BtoR_REQ0 & ~n10323;
  assign n10325 = ~i_RtoB_ACK0 & ~n10324;
  assign n10326 = ~n10263 & ~n10325;
  assign n10327 = ~controllable_DEQ & ~n10326;
  assign n10328 = ~n10318 & ~n10327;
  assign n10329 = i_FULL & ~n10328;
  assign n10330 = ~n5290 & ~n7727;
  assign n10331 = ~controllable_BtoR_REQ0 & ~n10330;
  assign n10332 = ~controllable_BtoR_REQ0 & ~n10331;
  assign n10333 = ~i_RtoB_ACK0 & ~n10332;
  assign n10334 = ~i_RtoB_ACK0 & ~n10333;
  assign n10335 = controllable_DEQ & ~n10334;
  assign n10336 = ~n5238 & ~n7703;
  assign n10337 = ~i_RtoB_ACK1 & ~n10336;
  assign n10338 = ~n7710 & ~n10337;
  assign n10339 = ~controllable_BtoR_REQ1 & ~n10338;
  assign n10340 = ~n10265 & ~n10339;
  assign n10341 = ~controllable_BtoR_REQ0 & ~n10340;
  assign n10342 = ~controllable_BtoR_REQ0 & ~n10341;
  assign n10343 = ~i_RtoB_ACK0 & ~n10342;
  assign n10344 = ~n10263 & ~n10343;
  assign n10345 = ~controllable_DEQ & ~n10344;
  assign n10346 = ~n10335 & ~n10345;
  assign n10347 = ~i_FULL & ~n10346;
  assign n10348 = ~n10329 & ~n10347;
  assign n10349 = ~i_nEMPTY & ~n10348;
  assign n10350 = ~n10312 & ~n10349;
  assign n10351 = controllable_BtoS_ACK0 & ~n10350;
  assign n10352 = ~n7802 & ~n8854;
  assign n10353 = ~controllable_BtoR_REQ1 & ~n10352;
  assign n10354 = ~n7790 & ~n10353;
  assign n10355 = ~controllable_BtoR_REQ0 & ~n10354;
  assign n10356 = ~controllable_BtoR_REQ0 & ~n10355;
  assign n10357 = i_RtoB_ACK0 & ~n10356;
  assign n10358 = ~n7805 & ~n8861;
  assign n10359 = controllable_BtoR_REQ1 & ~n10358;
  assign n10360 = ~n7795 & ~n8864;
  assign n10361 = ~i_RtoB_ACK1 & ~n10360;
  assign n10362 = ~n7802 & ~n10361;
  assign n10363 = ~controllable_BtoR_REQ1 & ~n10362;
  assign n10364 = ~n10359 & ~n10363;
  assign n10365 = ~controllable_BtoR_REQ0 & ~n10364;
  assign n10366 = ~controllable_BtoR_REQ0 & ~n10365;
  assign n10367 = ~i_RtoB_ACK0 & ~n10366;
  assign n10368 = ~n10357 & ~n10367;
  assign n10369 = controllable_DEQ & ~n10368;
  assign n10370 = i_RtoB_ACK1 & ~n7794;
  assign n10371 = ~n8876 & ~n10370;
  assign n10372 = ~controllable_BtoR_REQ1 & ~n10371;
  assign n10373 = ~n7819 & ~n10372;
  assign n10374 = ~controllable_BtoR_REQ0 & ~n10373;
  assign n10375 = ~controllable_BtoR_REQ0 & ~n10374;
  assign n10376 = i_RtoB_ACK0 & ~n10375;
  assign n10377 = ~n7808 & ~n8883;
  assign n10378 = controllable_BtoR_REQ1 & ~n10377;
  assign n10379 = ~n7820 & ~n10378;
  assign n10380 = ~controllable_BtoR_REQ0 & ~n10379;
  assign n10381 = ~controllable_BtoR_REQ0 & ~n10380;
  assign n10382 = ~i_RtoB_ACK0 & ~n10381;
  assign n10383 = ~n10376 & ~n10382;
  assign n10384 = ~controllable_DEQ & ~n10383;
  assign n10385 = ~n10369 & ~n10384;
  assign n10386 = i_FULL & ~n10385;
  assign n10387 = ~n7802 & ~n8876;
  assign n10388 = ~controllable_BtoR_REQ1 & ~n10387;
  assign n10389 = ~n10359 & ~n10388;
  assign n10390 = ~controllable_BtoR_REQ0 & ~n10389;
  assign n10391 = ~controllable_BtoR_REQ0 & ~n10390;
  assign n10392 = ~i_RtoB_ACK0 & ~n10391;
  assign n10393 = ~n10357 & ~n10392;
  assign n10394 = controllable_DEQ & ~n10393;
  assign n10395 = ~n10361 & ~n10370;
  assign n10396 = ~controllable_BtoR_REQ1 & ~n10395;
  assign n10397 = ~n10378 & ~n10396;
  assign n10398 = ~controllable_BtoR_REQ0 & ~n10397;
  assign n10399 = ~controllable_BtoR_REQ0 & ~n10398;
  assign n10400 = ~i_RtoB_ACK0 & ~n10399;
  assign n10401 = ~n10376 & ~n10400;
  assign n10402 = ~controllable_DEQ & ~n10401;
  assign n10403 = ~n10394 & ~n10402;
  assign n10404 = ~i_FULL & ~n10403;
  assign n10405 = ~n10386 & ~n10404;
  assign n10406 = i_nEMPTY & ~n10405;
  assign n10407 = ~n7835 & ~n8917;
  assign n10408 = ~controllable_BtoR_REQ0 & ~n10407;
  assign n10409 = ~controllable_BtoR_REQ0 & ~n10408;
  assign n10410 = ~i_RtoB_ACK0 & ~n10409;
  assign n10411 = ~i_RtoB_ACK0 & ~n10410;
  assign n10412 = controllable_DEQ & ~n10411;
  assign n10413 = ~i_RtoB_ACK1 & ~n7796;
  assign n10414 = ~n8861 & ~n10413;
  assign n10415 = controllable_BtoR_REQ1 & ~n10414;
  assign n10416 = ~n7797 & ~n10415;
  assign n10417 = ~controllable_BtoR_REQ0 & ~n10416;
  assign n10418 = ~controllable_BtoR_REQ0 & ~n10417;
  assign n10419 = ~i_RtoB_ACK0 & ~n10418;
  assign n10420 = ~n10357 & ~n10419;
  assign n10421 = ~controllable_DEQ & ~n10420;
  assign n10422 = ~n10412 & ~n10421;
  assign n10423 = i_FULL & ~n10422;
  assign n10424 = ~n7819 & ~n8936;
  assign n10425 = ~controllable_BtoR_REQ0 & ~n10424;
  assign n10426 = ~controllable_BtoR_REQ0 & ~n10425;
  assign n10427 = ~i_RtoB_ACK0 & ~n10426;
  assign n10428 = ~i_RtoB_ACK0 & ~n10427;
  assign n10429 = controllable_DEQ & ~n10428;
  assign n10430 = ~n7795 & ~n8946;
  assign n10431 = ~i_RtoB_ACK1 & ~n10430;
  assign n10432 = ~n7802 & ~n10431;
  assign n10433 = ~controllable_BtoR_REQ1 & ~n10432;
  assign n10434 = ~n10359 & ~n10433;
  assign n10435 = ~controllable_BtoR_REQ0 & ~n10434;
  assign n10436 = ~controllable_BtoR_REQ0 & ~n10435;
  assign n10437 = ~i_RtoB_ACK0 & ~n10436;
  assign n10438 = ~n10357 & ~n10437;
  assign n10439 = ~controllable_DEQ & ~n10438;
  assign n10440 = ~n10429 & ~n10439;
  assign n10441 = ~i_FULL & ~n10440;
  assign n10442 = ~n10423 & ~n10441;
  assign n10443 = ~i_nEMPTY & ~n10442;
  assign n10444 = ~n10406 & ~n10443;
  assign n10445 = ~controllable_BtoS_ACK0 & ~n10444;
  assign n10446 = ~n10351 & ~n10445;
  assign n10447 = n4465 & ~n10446;
  assign n10448 = ~n5307 & ~n10445;
  assign n10449 = ~n4465 & ~n10448;
  assign n10450 = ~n10447 & ~n10449;
  assign n10451 = i_StoB_REQ10 & ~n10450;
  assign n10452 = ~i_StoB_REQ0 & ~n9770;
  assign n10453 = ~i_StoB_REQ0 & ~n10452;
  assign n10454 = i_StoB_REQ14 & ~n10453;
  assign n10455 = ~n7907 & ~n10454;
  assign n10456 = controllable_BtoS_ACK14 & ~n10455;
  assign n10457 = ~n9300 & ~n10456;
  assign n10458 = controllable_ENQ & ~n10457;
  assign n10459 = controllable_ENQ & ~n10458;
  assign n10460 = ~i_RtoB_ACK1 & ~n10459;
  assign n10461 = ~n7935 & ~n10460;
  assign n10462 = ~controllable_BtoR_REQ1 & ~n10461;
  assign n10463 = ~n7905 & ~n10462;
  assign n10464 = ~controllable_BtoR_REQ0 & ~n10463;
  assign n10465 = ~controllable_BtoR_REQ0 & ~n10464;
  assign n10466 = i_RtoB_ACK0 & ~n10465;
  assign n10467 = ~n7927 & ~n9302;
  assign n10468 = i_RtoB_ACK1 & ~n10467;
  assign n10469 = ~n7932 & ~n10468;
  assign n10470 = controllable_BtoR_REQ1 & ~n10469;
  assign n10471 = ~i_StoB_REQ0 & ~n9887;
  assign n10472 = ~n5312 & ~n10471;
  assign n10473 = ~controllable_BtoS_ACK14 & ~n10472;
  assign n10474 = ~n8223 & ~n10473;
  assign n10475 = controllable_ENQ & ~n10474;
  assign n10476 = ~controllable_ENQ & ~n10457;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = ~i_RtoB_ACK1 & ~n10477;
  assign n10479 = ~n7935 & ~n10478;
  assign n10480 = ~controllable_BtoR_REQ1 & ~n10479;
  assign n10481 = ~n10470 & ~n10480;
  assign n10482 = ~controllable_BtoR_REQ0 & ~n10481;
  assign n10483 = ~controllable_BtoR_REQ0 & ~n10482;
  assign n10484 = ~i_RtoB_ACK0 & ~n10483;
  assign n10485 = ~n10466 & ~n10484;
  assign n10486 = controllable_DEQ & ~n10485;
  assign n10487 = ~i_RtoB_ACK1 & ~n10457;
  assign n10488 = ~n7957 & ~n10487;
  assign n10489 = ~controllable_BtoR_REQ1 & ~n10488;
  assign n10490 = ~n7950 & ~n10489;
  assign n10491 = ~controllable_BtoR_REQ0 & ~n10490;
  assign n10492 = ~controllable_BtoR_REQ0 & ~n10491;
  assign n10493 = i_RtoB_ACK0 & ~n10492;
  assign n10494 = ~n7958 & ~n9517;
  assign n10495 = controllable_BtoR_REQ1 & ~n10494;
  assign n10496 = ~i_RtoB_ACK1 & ~n10474;
  assign n10497 = ~n7957 & ~n10496;
  assign n10498 = ~controllable_BtoR_REQ1 & ~n10497;
  assign n10499 = ~n10495 & ~n10498;
  assign n10500 = ~controllable_BtoR_REQ0 & ~n10499;
  assign n10501 = ~controllable_BtoR_REQ0 & ~n10500;
  assign n10502 = ~i_RtoB_ACK0 & ~n10501;
  assign n10503 = ~n10493 & ~n10502;
  assign n10504 = ~controllable_DEQ & ~n10503;
  assign n10505 = ~n10486 & ~n10504;
  assign n10506 = i_FULL & ~n10505;
  assign n10507 = ~n7972 & ~n10468;
  assign n10508 = controllable_BtoR_REQ1 & ~n10507;
  assign n10509 = ~n9302 & ~n10476;
  assign n10510 = ~i_RtoB_ACK1 & ~n10509;
  assign n10511 = ~n7935 & ~n10510;
  assign n10512 = ~controllable_BtoR_REQ1 & ~n10511;
  assign n10513 = ~n10508 & ~n10512;
  assign n10514 = ~controllable_BtoR_REQ0 & ~n10513;
  assign n10515 = ~controllable_BtoR_REQ0 & ~n10514;
  assign n10516 = ~i_RtoB_ACK0 & ~n10515;
  assign n10517 = ~n10466 & ~n10516;
  assign n10518 = controllable_DEQ & ~n10517;
  assign n10519 = ~n7938 & ~n9517;
  assign n10520 = controllable_BtoR_REQ1 & ~n10519;
  assign n10521 = ~n9545 & ~n10475;
  assign n10522 = ~i_RtoB_ACK1 & ~n10521;
  assign n10523 = ~n7957 & ~n10522;
  assign n10524 = ~controllable_BtoR_REQ1 & ~n10523;
  assign n10525 = ~n10520 & ~n10524;
  assign n10526 = ~controllable_BtoR_REQ0 & ~n10525;
  assign n10527 = ~controllable_BtoR_REQ0 & ~n10526;
  assign n10528 = ~i_RtoB_ACK0 & ~n10527;
  assign n10529 = ~n10493 & ~n10528;
  assign n10530 = ~controllable_DEQ & ~n10529;
  assign n10531 = ~n10518 & ~n10530;
  assign n10532 = ~i_FULL & ~n10531;
  assign n10533 = ~n10506 & ~n10532;
  assign n10534 = i_nEMPTY & ~n10533;
  assign n10535 = ~controllable_ENQ & ~n10476;
  assign n10536 = ~i_RtoB_ACK1 & ~n10535;
  assign n10537 = ~i_RtoB_ACK1 & ~n10536;
  assign n10538 = ~controllable_BtoR_REQ1 & ~n10537;
  assign n10539 = ~n8002 & ~n10538;
  assign n10540 = ~controllable_BtoR_REQ0 & ~n10539;
  assign n10541 = ~controllable_BtoR_REQ0 & ~n10540;
  assign n10542 = ~i_RtoB_ACK0 & ~n10541;
  assign n10543 = ~i_RtoB_ACK0 & ~n10542;
  assign n10544 = controllable_DEQ & ~n10543;
  assign n10545 = ~n8015 & ~n9571;
  assign n10546 = controllable_BtoR_REQ1 & ~n10545;
  assign n10547 = controllable_ENQ & ~n10475;
  assign n10548 = ~i_RtoB_ACK1 & ~n10547;
  assign n10549 = ~n7935 & ~n10548;
  assign n10550 = ~controllable_BtoR_REQ1 & ~n10549;
  assign n10551 = ~n10546 & ~n10550;
  assign n10552 = ~controllable_BtoR_REQ0 & ~n10551;
  assign n10553 = ~controllable_BtoR_REQ0 & ~n10552;
  assign n10554 = ~i_RtoB_ACK0 & ~n10553;
  assign n10555 = ~n10466 & ~n10554;
  assign n10556 = ~controllable_DEQ & ~n10555;
  assign n10557 = ~n10544 & ~n10556;
  assign n10558 = i_FULL & ~n10557;
  assign n10559 = ~i_RtoB_ACK1 & ~n10487;
  assign n10560 = ~controllable_BtoR_REQ1 & ~n10559;
  assign n10561 = ~n7950 & ~n10560;
  assign n10562 = ~controllable_BtoR_REQ0 & ~n10561;
  assign n10563 = ~controllable_BtoR_REQ0 & ~n10562;
  assign n10564 = ~i_RtoB_ACK0 & ~n10563;
  assign n10565 = ~i_RtoB_ACK0 & ~n10564;
  assign n10566 = controllable_DEQ & ~n10565;
  assign n10567 = ~n9597 & ~n10475;
  assign n10568 = ~i_RtoB_ACK1 & ~n10567;
  assign n10569 = ~n7935 & ~n10568;
  assign n10570 = ~controllable_BtoR_REQ1 & ~n10569;
  assign n10571 = ~n10470 & ~n10570;
  assign n10572 = ~controllable_BtoR_REQ0 & ~n10571;
  assign n10573 = ~controllable_BtoR_REQ0 & ~n10572;
  assign n10574 = ~i_RtoB_ACK0 & ~n10573;
  assign n10575 = ~n10466 & ~n10574;
  assign n10576 = ~controllable_DEQ & ~n10575;
  assign n10577 = ~n10566 & ~n10576;
  assign n10578 = ~i_FULL & ~n10577;
  assign n10579 = ~n10558 & ~n10578;
  assign n10580 = ~i_nEMPTY & ~n10579;
  assign n10581 = ~n10534 & ~n10580;
  assign n10582 = controllable_BtoS_ACK0 & ~n10581;
  assign n10583 = ~n7172 & ~n10452;
  assign n10584 = i_StoB_REQ14 & ~n10583;
  assign n10585 = ~n8075 & ~n10584;
  assign n10586 = controllable_BtoS_ACK14 & ~n10585;
  assign n10587 = ~n9633 & ~n10586;
  assign n10588 = controllable_ENQ & ~n10587;
  assign n10589 = controllable_ENQ & ~n10588;
  assign n10590 = ~i_RtoB_ACK1 & ~n10589;
  assign n10591 = ~n8099 & ~n10590;
  assign n10592 = ~controllable_BtoR_REQ1 & ~n10591;
  assign n10593 = ~n8074 & ~n10592;
  assign n10594 = ~controllable_BtoR_REQ0 & ~n10593;
  assign n10595 = ~controllable_BtoR_REQ0 & ~n10594;
  assign n10596 = i_RtoB_ACK0 & ~n10595;
  assign n10597 = ~n8091 & ~n9635;
  assign n10598 = i_RtoB_ACK1 & ~n10597;
  assign n10599 = ~n8096 & ~n10598;
  assign n10600 = controllable_BtoR_REQ1 & ~n10599;
  assign n10601 = ~n9632 & ~n9891;
  assign n10602 = controllable_ENQ & ~n10601;
  assign n10603 = ~controllable_ENQ & ~n10587;
  assign n10604 = ~n10602 & ~n10603;
  assign n10605 = ~i_RtoB_ACK1 & ~n10604;
  assign n10606 = ~n8099 & ~n10605;
  assign n10607 = ~controllable_BtoR_REQ1 & ~n10606;
  assign n10608 = ~n10600 & ~n10607;
  assign n10609 = ~controllable_BtoR_REQ0 & ~n10608;
  assign n10610 = ~controllable_BtoR_REQ0 & ~n10609;
  assign n10611 = ~i_RtoB_ACK0 & ~n10610;
  assign n10612 = ~n10596 & ~n10611;
  assign n10613 = controllable_DEQ & ~n10612;
  assign n10614 = ~i_RtoB_ACK1 & ~n10587;
  assign n10615 = ~n8121 & ~n10614;
  assign n10616 = ~controllable_BtoR_REQ1 & ~n10615;
  assign n10617 = ~n8114 & ~n10616;
  assign n10618 = ~controllable_BtoR_REQ0 & ~n10617;
  assign n10619 = ~controllable_BtoR_REQ0 & ~n10618;
  assign n10620 = i_RtoB_ACK0 & ~n10619;
  assign n10621 = ~n8122 & ~n9664;
  assign n10622 = controllable_BtoR_REQ1 & ~n10621;
  assign n10623 = ~i_RtoB_ACK1 & ~n10601;
  assign n10624 = ~n8121 & ~n10623;
  assign n10625 = ~controllable_BtoR_REQ1 & ~n10624;
  assign n10626 = ~n10622 & ~n10625;
  assign n10627 = ~controllable_BtoR_REQ0 & ~n10626;
  assign n10628 = ~controllable_BtoR_REQ0 & ~n10627;
  assign n10629 = ~i_RtoB_ACK0 & ~n10628;
  assign n10630 = ~n10620 & ~n10629;
  assign n10631 = ~controllable_DEQ & ~n10630;
  assign n10632 = ~n10613 & ~n10631;
  assign n10633 = i_FULL & ~n10632;
  assign n10634 = ~n8136 & ~n10598;
  assign n10635 = controllable_BtoR_REQ1 & ~n10634;
  assign n10636 = ~n9635 & ~n10603;
  assign n10637 = ~i_RtoB_ACK1 & ~n10636;
  assign n10638 = ~n8099 & ~n10637;
  assign n10639 = ~controllable_BtoR_REQ1 & ~n10638;
  assign n10640 = ~n10635 & ~n10639;
  assign n10641 = ~controllable_BtoR_REQ0 & ~n10640;
  assign n10642 = ~controllable_BtoR_REQ0 & ~n10641;
  assign n10643 = ~i_RtoB_ACK0 & ~n10642;
  assign n10644 = ~n10596 & ~n10643;
  assign n10645 = controllable_DEQ & ~n10644;
  assign n10646 = ~n8102 & ~n9664;
  assign n10647 = controllable_BtoR_REQ1 & ~n10646;
  assign n10648 = ~n9692 & ~n10602;
  assign n10649 = ~i_RtoB_ACK1 & ~n10648;
  assign n10650 = ~n8121 & ~n10649;
  assign n10651 = ~controllable_BtoR_REQ1 & ~n10650;
  assign n10652 = ~n10647 & ~n10651;
  assign n10653 = ~controllable_BtoR_REQ0 & ~n10652;
  assign n10654 = ~controllable_BtoR_REQ0 & ~n10653;
  assign n10655 = ~i_RtoB_ACK0 & ~n10654;
  assign n10656 = ~n10620 & ~n10655;
  assign n10657 = ~controllable_DEQ & ~n10656;
  assign n10658 = ~n10645 & ~n10657;
  assign n10659 = ~i_FULL & ~n10658;
  assign n10660 = ~n10633 & ~n10659;
  assign n10661 = i_nEMPTY & ~n10660;
  assign n10662 = ~controllable_ENQ & ~n10603;
  assign n10663 = ~i_RtoB_ACK1 & ~n10662;
  assign n10664 = ~i_RtoB_ACK1 & ~n10663;
  assign n10665 = ~controllable_BtoR_REQ1 & ~n10664;
  assign n10666 = ~n8166 & ~n10665;
  assign n10667 = ~controllable_BtoR_REQ0 & ~n10666;
  assign n10668 = ~controllable_BtoR_REQ0 & ~n10667;
  assign n10669 = ~i_RtoB_ACK0 & ~n10668;
  assign n10670 = ~i_RtoB_ACK0 & ~n10669;
  assign n10671 = controllable_DEQ & ~n10670;
  assign n10672 = ~n8179 & ~n9718;
  assign n10673 = controllable_BtoR_REQ1 & ~n10672;
  assign n10674 = controllable_ENQ & ~n10602;
  assign n10675 = ~i_RtoB_ACK1 & ~n10674;
  assign n10676 = ~n8099 & ~n10675;
  assign n10677 = ~controllable_BtoR_REQ1 & ~n10676;
  assign n10678 = ~n10673 & ~n10677;
  assign n10679 = ~controllable_BtoR_REQ0 & ~n10678;
  assign n10680 = ~controllable_BtoR_REQ0 & ~n10679;
  assign n10681 = ~i_RtoB_ACK0 & ~n10680;
  assign n10682 = ~n10596 & ~n10681;
  assign n10683 = ~controllable_DEQ & ~n10682;
  assign n10684 = ~n10671 & ~n10683;
  assign n10685 = i_FULL & ~n10684;
  assign n10686 = ~i_RtoB_ACK1 & ~n10614;
  assign n10687 = ~controllable_BtoR_REQ1 & ~n10686;
  assign n10688 = ~n8114 & ~n10687;
  assign n10689 = ~controllable_BtoR_REQ0 & ~n10688;
  assign n10690 = ~controllable_BtoR_REQ0 & ~n10689;
  assign n10691 = ~i_RtoB_ACK0 & ~n10690;
  assign n10692 = ~i_RtoB_ACK0 & ~n10691;
  assign n10693 = controllable_DEQ & ~n10692;
  assign n10694 = ~n9747 & ~n10602;
  assign n10695 = ~i_RtoB_ACK1 & ~n10694;
  assign n10696 = ~n8099 & ~n10695;
  assign n10697 = ~controllable_BtoR_REQ1 & ~n10696;
  assign n10698 = ~n10600 & ~n10697;
  assign n10699 = ~controllable_BtoR_REQ0 & ~n10698;
  assign n10700 = ~controllable_BtoR_REQ0 & ~n10699;
  assign n10701 = ~i_RtoB_ACK0 & ~n10700;
  assign n10702 = ~n10596 & ~n10701;
  assign n10703 = ~controllable_DEQ & ~n10702;
  assign n10704 = ~n10693 & ~n10703;
  assign n10705 = ~i_FULL & ~n10704;
  assign n10706 = ~n10685 & ~n10705;
  assign n10707 = ~i_nEMPTY & ~n10706;
  assign n10708 = ~n10661 & ~n10707;
  assign n10709 = ~controllable_BtoS_ACK0 & ~n10708;
  assign n10710 = ~n10582 & ~n10709;
  assign n10711 = n4465 & ~n10710;
  assign n10712 = ~n8239 & ~n9836;
  assign n10713 = ~controllable_BtoR_REQ1 & ~n10712;
  assign n10714 = ~n8221 & ~n10713;
  assign n10715 = ~controllable_BtoR_REQ0 & ~n10714;
  assign n10716 = ~controllable_BtoR_REQ0 & ~n10715;
  assign n10717 = i_RtoB_ACK0 & ~n10716;
  assign n10718 = ~n8236 & ~n9789;
  assign n10719 = controllable_BtoR_REQ1 & ~n10718;
  assign n10720 = ~n8239 & ~n9813;
  assign n10721 = ~controllable_BtoR_REQ1 & ~n10720;
  assign n10722 = ~n10719 & ~n10721;
  assign n10723 = ~controllable_BtoR_REQ0 & ~n10722;
  assign n10724 = ~controllable_BtoR_REQ0 & ~n10723;
  assign n10725 = ~i_RtoB_ACK0 & ~n10724;
  assign n10726 = ~n10717 & ~n10725;
  assign n10727 = controllable_DEQ & ~n10726;
  assign n10728 = i_RtoB_ACK1 & ~n8224;
  assign n10729 = ~n9813 & ~n10728;
  assign n10730 = ~controllable_BtoR_REQ1 & ~n10729;
  assign n10731 = ~n8251 & ~n10730;
  assign n10732 = ~controllable_BtoR_REQ0 & ~n10731;
  assign n10733 = ~controllable_BtoR_REQ0 & ~n10732;
  assign n10734 = i_RtoB_ACK0 & ~n10733;
  assign n10735 = ~n8240 & ~n9517;
  assign n10736 = controllable_BtoR_REQ1 & ~n10735;
  assign n10737 = ~n10730 & ~n10736;
  assign n10738 = ~controllable_BtoR_REQ0 & ~n10737;
  assign n10739 = ~controllable_BtoR_REQ0 & ~n10738;
  assign n10740 = ~i_RtoB_ACK0 & ~n10739;
  assign n10741 = ~n10734 & ~n10740;
  assign n10742 = ~controllable_DEQ & ~n10741;
  assign n10743 = ~n10727 & ~n10742;
  assign n10744 = i_nEMPTY & ~n10743;
  assign n10745 = ~n8267 & ~n10049;
  assign n10746 = ~controllable_BtoR_REQ0 & ~n10745;
  assign n10747 = ~controllable_BtoR_REQ0 & ~n10746;
  assign n10748 = ~i_RtoB_ACK0 & ~n10747;
  assign n10749 = ~i_RtoB_ACK0 & ~n10748;
  assign n10750 = controllable_DEQ & ~n10749;
  assign n10751 = ~n8615 & ~n9571;
  assign n10752 = controllable_BtoR_REQ1 & ~n10751;
  assign n10753 = ~n10713 & ~n10752;
  assign n10754 = ~controllable_BtoR_REQ0 & ~n10753;
  assign n10755 = ~controllable_BtoR_REQ0 & ~n10754;
  assign n10756 = ~i_RtoB_ACK0 & ~n10755;
  assign n10757 = ~n10717 & ~n10756;
  assign n10758 = ~controllable_DEQ & ~n10757;
  assign n10759 = ~n10750 & ~n10758;
  assign n10760 = i_FULL & ~n10759;
  assign n10761 = ~n8251 & ~n10061;
  assign n10762 = ~controllable_BtoR_REQ0 & ~n10761;
  assign n10763 = ~controllable_BtoR_REQ0 & ~n10762;
  assign n10764 = ~i_RtoB_ACK0 & ~n10763;
  assign n10765 = ~i_RtoB_ACK0 & ~n10764;
  assign n10766 = controllable_DEQ & ~n10765;
  assign n10767 = ~n8239 & ~n9856;
  assign n10768 = ~controllable_BtoR_REQ1 & ~n10767;
  assign n10769 = ~n10719 & ~n10768;
  assign n10770 = ~controllable_BtoR_REQ0 & ~n10769;
  assign n10771 = ~controllable_BtoR_REQ0 & ~n10770;
  assign n10772 = ~i_RtoB_ACK0 & ~n10771;
  assign n10773 = ~n10717 & ~n10772;
  assign n10774 = ~controllable_DEQ & ~n10773;
  assign n10775 = ~n10766 & ~n10774;
  assign n10776 = ~i_FULL & ~n10775;
  assign n10777 = ~n10760 & ~n10776;
  assign n10778 = ~i_nEMPTY & ~n10777;
  assign n10779 = ~n10744 & ~n10778;
  assign n10780 = controllable_BtoS_ACK0 & ~n10779;
  assign n10781 = ~n8340 & ~n9871;
  assign n10782 = ~controllable_BtoR_REQ1 & ~n10781;
  assign n10783 = ~n8321 & ~n10782;
  assign n10784 = ~controllable_BtoR_REQ0 & ~n10783;
  assign n10785 = ~controllable_BtoR_REQ0 & ~n10784;
  assign n10786 = i_RtoB_ACK0 & ~n10785;
  assign n10787 = ~n8332 & ~n9635;
  assign n10788 = i_RtoB_ACK1 & ~n10787;
  assign n10789 = ~n8337 & ~n10788;
  assign n10790 = controllable_BtoR_REQ1 & ~n10789;
  assign n10791 = ~n8340 & ~n10649;
  assign n10792 = ~controllable_BtoR_REQ1 & ~n10791;
  assign n10793 = ~n10790 & ~n10792;
  assign n10794 = ~controllable_BtoR_REQ0 & ~n10793;
  assign n10795 = ~controllable_BtoR_REQ0 & ~n10794;
  assign n10796 = ~i_RtoB_ACK0 & ~n10795;
  assign n10797 = ~n10786 & ~n10796;
  assign n10798 = controllable_DEQ & ~n10797;
  assign n10799 = ~n8361 & ~n9904;
  assign n10800 = ~controllable_BtoR_REQ1 & ~n10799;
  assign n10801 = ~n8355 & ~n10800;
  assign n10802 = ~controllable_BtoR_REQ0 & ~n10801;
  assign n10803 = ~controllable_BtoR_REQ0 & ~n10802;
  assign n10804 = i_RtoB_ACK0 & ~n10803;
  assign n10805 = ~n8361 & ~n10623;
  assign n10806 = ~controllable_BtoR_REQ1 & ~n10805;
  assign n10807 = ~n10622 & ~n10806;
  assign n10808 = ~controllable_BtoR_REQ0 & ~n10807;
  assign n10809 = ~controllable_BtoR_REQ0 & ~n10808;
  assign n10810 = ~i_RtoB_ACK0 & ~n10809;
  assign n10811 = ~n10804 & ~n10810;
  assign n10812 = ~controllable_DEQ & ~n10811;
  assign n10813 = ~n10798 & ~n10812;
  assign n10814 = i_FULL & ~n10813;
  assign n10815 = ~n8375 & ~n10788;
  assign n10816 = controllable_BtoR_REQ1 & ~n10815;
  assign n10817 = ~n8340 & ~n9904;
  assign n10818 = ~controllable_BtoR_REQ1 & ~n10817;
  assign n10819 = ~n10816 & ~n10818;
  assign n10820 = ~controllable_BtoR_REQ0 & ~n10819;
  assign n10821 = ~controllable_BtoR_REQ0 & ~n10820;
  assign n10822 = ~i_RtoB_ACK0 & ~n10821;
  assign n10823 = ~n10786 & ~n10822;
  assign n10824 = controllable_DEQ & ~n10823;
  assign n10825 = ~n8343 & ~n9664;
  assign n10826 = controllable_BtoR_REQ1 & ~n10825;
  assign n10827 = ~n8361 & ~n10649;
  assign n10828 = ~controllable_BtoR_REQ1 & ~n10827;
  assign n10829 = ~n10826 & ~n10828;
  assign n10830 = ~controllable_BtoR_REQ0 & ~n10829;
  assign n10831 = ~controllable_BtoR_REQ0 & ~n10830;
  assign n10832 = ~i_RtoB_ACK0 & ~n10831;
  assign n10833 = ~n10804 & ~n10832;
  assign n10834 = ~controllable_DEQ & ~n10833;
  assign n10835 = ~n10824 & ~n10834;
  assign n10836 = ~i_FULL & ~n10835;
  assign n10837 = ~n10814 & ~n10836;
  assign n10838 = i_nEMPTY & ~n10837;
  assign n10839 = ~n8405 & ~n9951;
  assign n10840 = ~controllable_BtoR_REQ0 & ~n10839;
  assign n10841 = ~controllable_BtoR_REQ0 & ~n10840;
  assign n10842 = ~i_RtoB_ACK0 & ~n10841;
  assign n10843 = ~i_RtoB_ACK0 & ~n10842;
  assign n10844 = controllable_DEQ & ~n10843;
  assign n10845 = ~n8340 & ~n10675;
  assign n10846 = ~controllable_BtoR_REQ1 & ~n10845;
  assign n10847 = ~n10673 & ~n10846;
  assign n10848 = ~controllable_BtoR_REQ0 & ~n10847;
  assign n10849 = ~controllable_BtoR_REQ0 & ~n10848;
  assign n10850 = ~i_RtoB_ACK0 & ~n10849;
  assign n10851 = ~n10786 & ~n10850;
  assign n10852 = ~controllable_DEQ & ~n10851;
  assign n10853 = ~n10844 & ~n10852;
  assign n10854 = i_FULL & ~n10853;
  assign n10855 = ~n8355 & ~n9973;
  assign n10856 = ~controllable_BtoR_REQ0 & ~n10855;
  assign n10857 = ~controllable_BtoR_REQ0 & ~n10856;
  assign n10858 = ~i_RtoB_ACK0 & ~n10857;
  assign n10859 = ~i_RtoB_ACK0 & ~n10858;
  assign n10860 = controllable_DEQ & ~n10859;
  assign n10861 = ~n8340 & ~n10695;
  assign n10862 = ~controllable_BtoR_REQ1 & ~n10861;
  assign n10863 = ~n10790 & ~n10862;
  assign n10864 = ~controllable_BtoR_REQ0 & ~n10863;
  assign n10865 = ~controllable_BtoR_REQ0 & ~n10864;
  assign n10866 = ~i_RtoB_ACK0 & ~n10865;
  assign n10867 = ~n10786 & ~n10866;
  assign n10868 = ~controllable_DEQ & ~n10867;
  assign n10869 = ~n10860 & ~n10868;
  assign n10870 = ~i_FULL & ~n10869;
  assign n10871 = ~n10854 & ~n10870;
  assign n10872 = ~i_nEMPTY & ~n10871;
  assign n10873 = ~n10838 & ~n10872;
  assign n10874 = ~controllable_BtoS_ACK0 & ~n10873;
  assign n10875 = ~n10780 & ~n10874;
  assign n10876 = ~n4465 & ~n10875;
  assign n10877 = ~n10711 & ~n10876;
  assign n10878 = ~i_StoB_REQ10 & ~n10877;
  assign n10879 = ~n10451 & ~n10878;
  assign n10880 = controllable_BtoS_ACK10 & ~n10879;
  assign n10881 = ~n7935 & ~n9836;
  assign n10882 = ~controllable_BtoR_REQ1 & ~n10881;
  assign n10883 = ~n8464 & ~n10882;
  assign n10884 = ~controllable_BtoR_REQ0 & ~n10883;
  assign n10885 = ~controllable_BtoR_REQ0 & ~n10884;
  assign n10886 = i_RtoB_ACK0 & ~n10885;
  assign n10887 = ~n8469 & ~n9302;
  assign n10888 = i_RtoB_ACK1 & ~n10887;
  assign n10889 = ~n7938 & ~n10888;
  assign n10890 = controllable_BtoR_REQ1 & ~n10889;
  assign n10891 = ~n7935 & ~n10522;
  assign n10892 = ~controllable_BtoR_REQ1 & ~n10891;
  assign n10893 = ~n10890 & ~n10892;
  assign n10894 = ~controllable_BtoR_REQ0 & ~n10893;
  assign n10895 = ~controllable_BtoR_REQ0 & ~n10894;
  assign n10896 = ~i_RtoB_ACK0 & ~n10895;
  assign n10897 = ~n10886 & ~n10896;
  assign n10898 = controllable_DEQ & ~n10897;
  assign n10899 = ~n7957 & ~n9813;
  assign n10900 = ~controllable_BtoR_REQ1 & ~n10899;
  assign n10901 = ~n8482 & ~n10900;
  assign n10902 = ~controllable_BtoR_REQ0 & ~n10901;
  assign n10903 = ~controllable_BtoR_REQ0 & ~n10902;
  assign n10904 = i_RtoB_ACK0 & ~n10903;
  assign n10905 = ~n10502 & ~n10904;
  assign n10906 = ~controllable_DEQ & ~n10905;
  assign n10907 = ~n10898 & ~n10906;
  assign n10908 = i_FULL & ~n10907;
  assign n10909 = ~n7975 & ~n10888;
  assign n10910 = controllable_BtoR_REQ1 & ~n10909;
  assign n10911 = ~n7935 & ~n9813;
  assign n10912 = ~controllable_BtoR_REQ1 & ~n10911;
  assign n10913 = ~n10910 & ~n10912;
  assign n10914 = ~controllable_BtoR_REQ0 & ~n10913;
  assign n10915 = ~controllable_BtoR_REQ0 & ~n10914;
  assign n10916 = ~i_RtoB_ACK0 & ~n10915;
  assign n10917 = ~n10886 & ~n10916;
  assign n10918 = controllable_DEQ & ~n10917;
  assign n10919 = ~n10528 & ~n10904;
  assign n10920 = ~controllable_DEQ & ~n10919;
  assign n10921 = ~n10918 & ~n10920;
  assign n10922 = ~i_FULL & ~n10921;
  assign n10923 = ~n10908 & ~n10922;
  assign n10924 = i_nEMPTY & ~n10923;
  assign n10925 = ~n8510 & ~n10049;
  assign n10926 = ~controllable_BtoR_REQ0 & ~n10925;
  assign n10927 = ~controllable_BtoR_REQ0 & ~n10926;
  assign n10928 = ~i_RtoB_ACK0 & ~n10927;
  assign n10929 = ~i_RtoB_ACK0 & ~n10928;
  assign n10930 = controllable_DEQ & ~n10929;
  assign n10931 = ~n10554 & ~n10886;
  assign n10932 = ~controllable_DEQ & ~n10931;
  assign n10933 = ~n10930 & ~n10932;
  assign n10934 = i_FULL & ~n10933;
  assign n10935 = ~n8482 & ~n10061;
  assign n10936 = ~controllable_BtoR_REQ0 & ~n10935;
  assign n10937 = ~controllable_BtoR_REQ0 & ~n10936;
  assign n10938 = ~i_RtoB_ACK0 & ~n10937;
  assign n10939 = ~i_RtoB_ACK0 & ~n10938;
  assign n10940 = controllable_DEQ & ~n10939;
  assign n10941 = ~controllable_DEQ & ~n10897;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = ~i_FULL & ~n10942;
  assign n10944 = ~n10934 & ~n10943;
  assign n10945 = ~i_nEMPTY & ~n10944;
  assign n10946 = ~n10924 & ~n10945;
  assign n10947 = controllable_BtoS_ACK0 & ~n10946;
  assign n10948 = ~n8099 & ~n9871;
  assign n10949 = ~controllable_BtoR_REQ1 & ~n10948;
  assign n10950 = ~n8543 & ~n10949;
  assign n10951 = ~controllable_BtoR_REQ0 & ~n10950;
  assign n10952 = ~controllable_BtoR_REQ0 & ~n10951;
  assign n10953 = i_RtoB_ACK0 & ~n10952;
  assign n10954 = ~n8548 & ~n9635;
  assign n10955 = i_RtoB_ACK1 & ~n10954;
  assign n10956 = ~n8102 & ~n10955;
  assign n10957 = controllable_BtoR_REQ1 & ~n10956;
  assign n10958 = ~n8099 & ~n10649;
  assign n10959 = ~controllable_BtoR_REQ1 & ~n10958;
  assign n10960 = ~n10957 & ~n10959;
  assign n10961 = ~controllable_BtoR_REQ0 & ~n10960;
  assign n10962 = ~controllable_BtoR_REQ0 & ~n10961;
  assign n10963 = ~i_RtoB_ACK0 & ~n10962;
  assign n10964 = ~n10953 & ~n10963;
  assign n10965 = controllable_DEQ & ~n10964;
  assign n10966 = ~n8121 & ~n9904;
  assign n10967 = ~controllable_BtoR_REQ1 & ~n10966;
  assign n10968 = ~n8561 & ~n10967;
  assign n10969 = ~controllable_BtoR_REQ0 & ~n10968;
  assign n10970 = ~controllable_BtoR_REQ0 & ~n10969;
  assign n10971 = i_RtoB_ACK0 & ~n10970;
  assign n10972 = ~n10629 & ~n10971;
  assign n10973 = ~controllable_DEQ & ~n10972;
  assign n10974 = ~n10965 & ~n10973;
  assign n10975 = i_FULL & ~n10974;
  assign n10976 = ~n8139 & ~n10955;
  assign n10977 = controllable_BtoR_REQ1 & ~n10976;
  assign n10978 = ~n8099 & ~n9904;
  assign n10979 = ~controllable_BtoR_REQ1 & ~n10978;
  assign n10980 = ~n10977 & ~n10979;
  assign n10981 = ~controllable_BtoR_REQ0 & ~n10980;
  assign n10982 = ~controllable_BtoR_REQ0 & ~n10981;
  assign n10983 = ~i_RtoB_ACK0 & ~n10982;
  assign n10984 = ~n10953 & ~n10983;
  assign n10985 = controllable_DEQ & ~n10984;
  assign n10986 = ~n10655 & ~n10971;
  assign n10987 = ~controllable_DEQ & ~n10986;
  assign n10988 = ~n10985 & ~n10987;
  assign n10989 = ~i_FULL & ~n10988;
  assign n10990 = ~n10975 & ~n10989;
  assign n10991 = i_nEMPTY & ~n10990;
  assign n10992 = ~n8589 & ~n9951;
  assign n10993 = ~controllable_BtoR_REQ0 & ~n10992;
  assign n10994 = ~controllable_BtoR_REQ0 & ~n10993;
  assign n10995 = ~i_RtoB_ACK0 & ~n10994;
  assign n10996 = ~i_RtoB_ACK0 & ~n10995;
  assign n10997 = controllable_DEQ & ~n10996;
  assign n10998 = ~n10681 & ~n10953;
  assign n10999 = ~controllable_DEQ & ~n10998;
  assign n11000 = ~n10997 & ~n10999;
  assign n11001 = i_FULL & ~n11000;
  assign n11002 = ~n8561 & ~n9973;
  assign n11003 = ~controllable_BtoR_REQ0 & ~n11002;
  assign n11004 = ~controllable_BtoR_REQ0 & ~n11003;
  assign n11005 = ~i_RtoB_ACK0 & ~n11004;
  assign n11006 = ~i_RtoB_ACK0 & ~n11005;
  assign n11007 = controllable_DEQ & ~n11006;
  assign n11008 = ~controllable_DEQ & ~n10964;
  assign n11009 = ~n11007 & ~n11008;
  assign n11010 = ~i_FULL & ~n11009;
  assign n11011 = ~n11001 & ~n11010;
  assign n11012 = ~i_nEMPTY & ~n11011;
  assign n11013 = ~n10991 & ~n11012;
  assign n11014 = ~controllable_BtoS_ACK0 & ~n11013;
  assign n11015 = ~n10947 & ~n11014;
  assign n11016 = n4465 & ~n11015;
  assign n11017 = ~n8617 & ~n10713;
  assign n11018 = ~controllable_BtoR_REQ0 & ~n11017;
  assign n11019 = ~controllable_BtoR_REQ0 & ~n11018;
  assign n11020 = i_RtoB_ACK0 & ~n11019;
  assign n11021 = ~n8240 & ~n10149;
  assign n11022 = controllable_BtoR_REQ1 & ~n11021;
  assign n11023 = ~n10721 & ~n11022;
  assign n11024 = ~controllable_BtoR_REQ0 & ~n11023;
  assign n11025 = ~controllable_BtoR_REQ0 & ~n11024;
  assign n11026 = ~i_RtoB_ACK0 & ~n11025;
  assign n11027 = ~n11020 & ~n11026;
  assign n11028 = controllable_DEQ & ~n11027;
  assign n11029 = ~n8633 & ~n10730;
  assign n11030 = ~controllable_BtoR_REQ0 & ~n11029;
  assign n11031 = ~controllable_BtoR_REQ0 & ~n11030;
  assign n11032 = i_RtoB_ACK0 & ~n11031;
  assign n11033 = ~n10740 & ~n11032;
  assign n11034 = ~controllable_DEQ & ~n11033;
  assign n11035 = ~n11028 & ~n11034;
  assign n11036 = i_nEMPTY & ~n11035;
  assign n11037 = ~n8643 & ~n10049;
  assign n11038 = ~controllable_BtoR_REQ0 & ~n11037;
  assign n11039 = ~controllable_BtoR_REQ0 & ~n11038;
  assign n11040 = ~i_RtoB_ACK0 & ~n11039;
  assign n11041 = ~i_RtoB_ACK0 & ~n11040;
  assign n11042 = controllable_DEQ & ~n11041;
  assign n11043 = ~n10756 & ~n11020;
  assign n11044 = ~controllable_DEQ & ~n11043;
  assign n11045 = ~n11042 & ~n11044;
  assign n11046 = i_FULL & ~n11045;
  assign n11047 = ~n8633 & ~n10061;
  assign n11048 = ~controllable_BtoR_REQ0 & ~n11047;
  assign n11049 = ~controllable_BtoR_REQ0 & ~n11048;
  assign n11050 = ~i_RtoB_ACK0 & ~n11049;
  assign n11051 = ~i_RtoB_ACK0 & ~n11050;
  assign n11052 = controllable_DEQ & ~n11051;
  assign n11053 = ~controllable_DEQ & ~n11027;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = ~i_FULL & ~n11054;
  assign n11056 = ~n11046 & ~n11055;
  assign n11057 = ~i_nEMPTY & ~n11056;
  assign n11058 = ~n11036 & ~n11057;
  assign n11059 = controllable_BtoS_ACK0 & ~n11058;
  assign n11060 = ~n8675 & ~n10782;
  assign n11061 = ~controllable_BtoR_REQ0 & ~n11060;
  assign n11062 = ~controllable_BtoR_REQ0 & ~n11061;
  assign n11063 = i_RtoB_ACK0 & ~n11062;
  assign n11064 = ~n8680 & ~n9635;
  assign n11065 = i_RtoB_ACK1 & ~n11064;
  assign n11066 = ~n8343 & ~n11065;
  assign n11067 = controllable_BtoR_REQ1 & ~n11066;
  assign n11068 = ~n10792 & ~n11067;
  assign n11069 = ~controllable_BtoR_REQ0 & ~n11068;
  assign n11070 = ~controllable_BtoR_REQ0 & ~n11069;
  assign n11071 = ~i_RtoB_ACK0 & ~n11070;
  assign n11072 = ~n11063 & ~n11071;
  assign n11073 = controllable_DEQ & ~n11072;
  assign n11074 = ~n8693 & ~n10800;
  assign n11075 = ~controllable_BtoR_REQ0 & ~n11074;
  assign n11076 = ~controllable_BtoR_REQ0 & ~n11075;
  assign n11077 = i_RtoB_ACK0 & ~n11076;
  assign n11078 = ~n10810 & ~n11077;
  assign n11079 = ~controllable_DEQ & ~n11078;
  assign n11080 = ~n11073 & ~n11079;
  assign n11081 = i_FULL & ~n11080;
  assign n11082 = ~n8378 & ~n11065;
  assign n11083 = controllable_BtoR_REQ1 & ~n11082;
  assign n11084 = ~n10818 & ~n11083;
  assign n11085 = ~controllable_BtoR_REQ0 & ~n11084;
  assign n11086 = ~controllable_BtoR_REQ0 & ~n11085;
  assign n11087 = ~i_RtoB_ACK0 & ~n11086;
  assign n11088 = ~n11063 & ~n11087;
  assign n11089 = controllable_DEQ & ~n11088;
  assign n11090 = ~n10832 & ~n11077;
  assign n11091 = ~controllable_DEQ & ~n11090;
  assign n11092 = ~n11089 & ~n11091;
  assign n11093 = ~i_FULL & ~n11092;
  assign n11094 = ~n11081 & ~n11093;
  assign n11095 = i_nEMPTY & ~n11094;
  assign n11096 = ~n8721 & ~n9951;
  assign n11097 = ~controllable_BtoR_REQ0 & ~n11096;
  assign n11098 = ~controllable_BtoR_REQ0 & ~n11097;
  assign n11099 = ~i_RtoB_ACK0 & ~n11098;
  assign n11100 = ~i_RtoB_ACK0 & ~n11099;
  assign n11101 = controllable_DEQ & ~n11100;
  assign n11102 = ~n10850 & ~n11063;
  assign n11103 = ~controllable_DEQ & ~n11102;
  assign n11104 = ~n11101 & ~n11103;
  assign n11105 = i_FULL & ~n11104;
  assign n11106 = ~n8693 & ~n9973;
  assign n11107 = ~controllable_BtoR_REQ0 & ~n11106;
  assign n11108 = ~controllable_BtoR_REQ0 & ~n11107;
  assign n11109 = ~i_RtoB_ACK0 & ~n11108;
  assign n11110 = ~i_RtoB_ACK0 & ~n11109;
  assign n11111 = controllable_DEQ & ~n11110;
  assign n11112 = ~controllable_DEQ & ~n11072;
  assign n11113 = ~n11111 & ~n11112;
  assign n11114 = ~i_FULL & ~n11113;
  assign n11115 = ~n11105 & ~n11114;
  assign n11116 = ~i_nEMPTY & ~n11115;
  assign n11117 = ~n11095 & ~n11116;
  assign n11118 = ~controllable_BtoS_ACK0 & ~n11117;
  assign n11119 = ~n11059 & ~n11118;
  assign n11120 = ~n4465 & ~n11119;
  assign n11121 = ~n11016 & ~n11120;
  assign n11122 = i_StoB_REQ10 & ~n11121;
  assign n11123 = ~n10878 & ~n11122;
  assign n11124 = ~controllable_BtoS_ACK10 & ~n11123;
  assign n11125 = ~n10880 & ~n11124;
  assign n11126 = ~n4464 & ~n11125;
  assign n11127 = ~n10257 & ~n11126;
  assign n11128 = ~n4463 & ~n11127;
  assign n11129 = ~n8754 & ~n11128;
  assign n11130 = n4462 & ~n11129;
  assign n11131 = ~i_StoB_REQ14 & ~n7692;
  assign n11132 = controllable_BtoS_ACK14 & ~n11131;
  assign n11133 = ~n7694 & ~n11132;
  assign n11134 = controllable_ENQ & ~n11133;
  assign n11135 = controllable_ENQ & ~n11134;
  assign n11136 = ~i_RtoB_ACK1 & ~n11135;
  assign n11137 = ~i_RtoB_ACK1 & ~n11136;
  assign n11138 = controllable_BtoR_REQ1 & ~n11137;
  assign n11139 = ~i_StoB_REQ14 & ~n7689;
  assign n11140 = ~i_StoB_REQ14 & ~n11139;
  assign n11141 = controllable_BtoS_ACK14 & ~n11140;
  assign n11142 = ~n7701 & ~n11141;
  assign n11143 = controllable_ENQ & ~n11142;
  assign n11144 = controllable_ENQ & ~n11143;
  assign n11145 = ~controllable_BtoR_REQ1 & ~n11144;
  assign n11146 = ~n11138 & ~n11145;
  assign n11147 = ~controllable_BtoR_REQ0 & ~n11146;
  assign n11148 = ~controllable_BtoR_REQ0 & ~n11147;
  assign n11149 = i_RtoB_ACK0 & ~n11148;
  assign n11150 = i_RtoB_ACK1 & ~n11144;
  assign n11151 = ~controllable_ENQ & ~n11133;
  assign n11152 = ~n11143 & ~n11151;
  assign n11153 = ~i_RtoB_ACK1 & ~n11152;
  assign n11154 = ~n11150 & ~n11153;
  assign n11155 = controllable_BtoR_REQ1 & ~n11154;
  assign n11156 = ~i_RtoB_ACK1 & ~n11142;
  assign n11157 = ~n11150 & ~n11156;
  assign n11158 = ~controllable_BtoR_REQ1 & ~n11157;
  assign n11159 = ~n11155 & ~n11158;
  assign n11160 = ~controllable_BtoR_REQ0 & ~n11159;
  assign n11161 = ~controllable_BtoR_REQ0 & ~n11160;
  assign n11162 = ~i_RtoB_ACK0 & ~n11161;
  assign n11163 = ~n11149 & ~n11162;
  assign n11164 = controllable_DEQ & ~n11163;
  assign n11165 = ~i_RtoB_ACK1 & ~n11133;
  assign n11166 = ~i_RtoB_ACK1 & ~n11165;
  assign n11167 = controllable_BtoR_REQ1 & ~n11166;
  assign n11168 = ~controllable_BtoR_REQ1 & ~n11142;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = ~controllable_BtoR_REQ0 & ~n11169;
  assign n11171 = ~controllable_BtoR_REQ0 & ~n11170;
  assign n11172 = i_RtoB_ACK0 & ~n11171;
  assign n11173 = ~controllable_BtoR_REQ0 & ~n11142;
  assign n11174 = ~controllable_BtoR_REQ0 & ~n11173;
  assign n11175 = ~i_RtoB_ACK0 & ~n11174;
  assign n11176 = ~n11172 & ~n11175;
  assign n11177 = ~controllable_DEQ & ~n11176;
  assign n11178 = ~n11164 & ~n11177;
  assign n11179 = i_nEMPTY & ~n11178;
  assign n11180 = ~controllable_ENQ & ~n11151;
  assign n11181 = ~i_RtoB_ACK1 & ~n11180;
  assign n11182 = ~i_RtoB_ACK1 & ~n11181;
  assign n11183 = controllable_BtoR_REQ1 & ~n11182;
  assign n11184 = ~controllable_ENQ & ~n11142;
  assign n11185 = ~controllable_ENQ & ~n11184;
  assign n11186 = ~i_RtoB_ACK1 & ~n11185;
  assign n11187 = ~i_RtoB_ACK1 & ~n11186;
  assign n11188 = ~controllable_BtoR_REQ1 & ~n11187;
  assign n11189 = ~n11183 & ~n11188;
  assign n11190 = ~controllable_BtoR_REQ0 & ~n11189;
  assign n11191 = ~controllable_BtoR_REQ0 & ~n11190;
  assign n11192 = ~i_RtoB_ACK0 & ~n11191;
  assign n11193 = ~i_RtoB_ACK0 & ~n11192;
  assign n11194 = controllable_DEQ & ~n11193;
  assign n11195 = ~controllable_BtoR_REQ0 & ~n11144;
  assign n11196 = ~controllable_BtoR_REQ0 & ~n11195;
  assign n11197 = ~i_RtoB_ACK0 & ~n11196;
  assign n11198 = ~n11149 & ~n11197;
  assign n11199 = ~controllable_DEQ & ~n11198;
  assign n11200 = ~n11194 & ~n11199;
  assign n11201 = i_FULL & ~n11200;
  assign n11202 = ~i_RtoB_ACK1 & ~n11156;
  assign n11203 = ~controllable_BtoR_REQ1 & ~n11202;
  assign n11204 = ~n11167 & ~n11203;
  assign n11205 = ~controllable_BtoR_REQ0 & ~n11204;
  assign n11206 = ~controllable_BtoR_REQ0 & ~n11205;
  assign n11207 = ~i_RtoB_ACK0 & ~n11206;
  assign n11208 = ~i_RtoB_ACK0 & ~n11207;
  assign n11209 = controllable_DEQ & ~n11208;
  assign n11210 = ~controllable_BtoR_REQ0 & ~n11154;
  assign n11211 = ~controllable_BtoR_REQ0 & ~n11210;
  assign n11212 = ~i_RtoB_ACK0 & ~n11211;
  assign n11213 = ~n11149 & ~n11212;
  assign n11214 = ~controllable_DEQ & ~n11213;
  assign n11215 = ~n11209 & ~n11214;
  assign n11216 = ~i_FULL & ~n11215;
  assign n11217 = ~n11201 & ~n11216;
  assign n11218 = ~i_nEMPTY & ~n11217;
  assign n11219 = ~n11179 & ~n11218;
  assign n11220 = controllable_BtoS_ACK0 & ~n11219;
  assign n11221 = ~n5413 & ~n11220;
  assign n11222 = n4465 & ~n11221;
  assign n11223 = ~n5415 & ~n11222;
  assign n11224 = i_StoB_REQ10 & ~n11223;
  assign n11225 = controllable_ENQ & ~n9596;
  assign n11226 = controllable_ENQ & ~n11225;
  assign n11227 = ~i_RtoB_ACK1 & ~n11226;
  assign n11228 = ~n7054 & ~n11227;
  assign n11229 = controllable_BtoR_REQ1 & ~n11228;
  assign n11230 = ~controllable_BtoR_REQ1 & ~n9570;
  assign n11231 = ~n11229 & ~n11230;
  assign n11232 = ~controllable_BtoR_REQ0 & ~n11231;
  assign n11233 = ~controllable_BtoR_REQ0 & ~n11232;
  assign n11234 = i_RtoB_ACK0 & ~n11233;
  assign n11235 = ~n9789 & ~n9856;
  assign n11236 = controllable_BtoR_REQ1 & ~n11235;
  assign n11237 = ~n9571 & ~n9813;
  assign n11238 = ~controllable_BtoR_REQ1 & ~n11237;
  assign n11239 = ~n11236 & ~n11238;
  assign n11240 = ~controllable_BtoR_REQ0 & ~n11239;
  assign n11241 = ~controllable_BtoR_REQ0 & ~n11240;
  assign n11242 = ~i_RtoB_ACK0 & ~n11241;
  assign n11243 = ~n11234 & ~n11242;
  assign n11244 = controllable_DEQ & ~n11243;
  assign n11245 = ~i_RtoB_ACK1 & ~n9596;
  assign n11246 = ~n7111 & ~n11245;
  assign n11247 = controllable_BtoR_REQ1 & ~n11246;
  assign n11248 = ~controllable_BtoR_REQ1 & ~n9301;
  assign n11249 = ~n11247 & ~n11248;
  assign n11250 = ~controllable_BtoR_REQ0 & ~n11249;
  assign n11251 = ~controllable_BtoR_REQ0 & ~n11250;
  assign n11252 = i_RtoB_ACK0 & ~n11251;
  assign n11253 = ~controllable_BtoR_REQ0 & ~n9301;
  assign n11254 = ~controllable_BtoR_REQ0 & ~n11253;
  assign n11255 = ~i_RtoB_ACK0 & ~n11254;
  assign n11256 = ~n11252 & ~n11255;
  assign n11257 = ~controllable_DEQ & ~n11256;
  assign n11258 = ~n11244 & ~n11257;
  assign n11259 = i_nEMPTY & ~n11258;
  assign n11260 = ~controllable_ENQ & ~n9597;
  assign n11261 = ~i_RtoB_ACK1 & ~n11260;
  assign n11262 = ~n7127 & ~n11261;
  assign n11263 = controllable_BtoR_REQ1 & ~n11262;
  assign n11264 = ~n10049 & ~n11263;
  assign n11265 = ~controllable_BtoR_REQ0 & ~n11264;
  assign n11266 = ~controllable_BtoR_REQ0 & ~n11265;
  assign n11267 = ~i_RtoB_ACK0 & ~n11266;
  assign n11268 = ~i_RtoB_ACK0 & ~n11267;
  assign n11269 = controllable_DEQ & ~n11268;
  assign n11270 = ~controllable_BtoR_REQ0 & ~n9570;
  assign n11271 = ~controllable_BtoR_REQ0 & ~n11270;
  assign n11272 = ~i_RtoB_ACK0 & ~n11271;
  assign n11273 = ~n11234 & ~n11272;
  assign n11274 = ~controllable_DEQ & ~n11273;
  assign n11275 = ~n11269 & ~n11274;
  assign n11276 = i_FULL & ~n11275;
  assign n11277 = ~n10061 & ~n11247;
  assign n11278 = ~controllable_BtoR_REQ0 & ~n11277;
  assign n11279 = ~controllable_BtoR_REQ0 & ~n11278;
  assign n11280 = ~i_RtoB_ACK0 & ~n11279;
  assign n11281 = ~i_RtoB_ACK0 & ~n11280;
  assign n11282 = controllable_DEQ & ~n11281;
  assign n11283 = ~n9571 & ~n9856;
  assign n11284 = ~controllable_BtoR_REQ1 & ~n11283;
  assign n11285 = ~n11236 & ~n11284;
  assign n11286 = ~controllable_BtoR_REQ0 & ~n11285;
  assign n11287 = ~controllable_BtoR_REQ0 & ~n11286;
  assign n11288 = ~i_RtoB_ACK0 & ~n11287;
  assign n11289 = ~n11234 & ~n11288;
  assign n11290 = ~controllable_DEQ & ~n11289;
  assign n11291 = ~n11282 & ~n11290;
  assign n11292 = ~i_FULL & ~n11291;
  assign n11293 = ~n11276 & ~n11292;
  assign n11294 = ~i_nEMPTY & ~n11293;
  assign n11295 = ~n11259 & ~n11294;
  assign n11296 = controllable_BtoS_ACK0 & ~n11295;
  assign n11297 = controllable_ENQ & ~n8945;
  assign n11298 = controllable_ENQ & ~n11297;
  assign n11299 = i_RtoB_ACK1 & ~n11298;
  assign n11300 = controllable_ENQ & ~n9746;
  assign n11301 = controllable_ENQ & ~n11300;
  assign n11302 = ~i_RtoB_ACK1 & ~n11301;
  assign n11303 = ~n11299 & ~n11302;
  assign n11304 = controllable_BtoR_REQ1 & ~n11303;
  assign n11305 = ~controllable_BtoR_REQ1 & ~n9717;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = ~controllable_BtoR_REQ0 & ~n11306;
  assign n11308 = ~controllable_BtoR_REQ0 & ~n11307;
  assign n11309 = i_RtoB_ACK0 & ~n11308;
  assign n11310 = ~n8946 & ~n9635;
  assign n11311 = i_RtoB_ACK1 & ~n11310;
  assign n11312 = ~n9635 & ~n9747;
  assign n11313 = ~i_RtoB_ACK1 & ~n11312;
  assign n11314 = ~n11311 & ~n11313;
  assign n11315 = controllable_BtoR_REQ1 & ~n11314;
  assign n11316 = ~n9718 & ~n9904;
  assign n11317 = ~controllable_BtoR_REQ1 & ~n11316;
  assign n11318 = ~n11315 & ~n11317;
  assign n11319 = ~controllable_BtoR_REQ0 & ~n11318;
  assign n11320 = ~controllable_BtoR_REQ0 & ~n11319;
  assign n11321 = ~i_RtoB_ACK0 & ~n11320;
  assign n11322 = ~n11309 & ~n11321;
  assign n11323 = controllable_DEQ & ~n11322;
  assign n11324 = i_RtoB_ACK1 & ~n8945;
  assign n11325 = ~i_RtoB_ACK1 & ~n9746;
  assign n11326 = ~n11324 & ~n11325;
  assign n11327 = controllable_BtoR_REQ1 & ~n11326;
  assign n11328 = ~controllable_BtoR_REQ1 & ~n9634;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~controllable_BtoR_REQ0 & ~n11329;
  assign n11331 = ~controllable_BtoR_REQ0 & ~n11330;
  assign n11332 = i_RtoB_ACK0 & ~n11331;
  assign n11333 = ~controllable_BtoR_REQ0 & ~n9634;
  assign n11334 = ~controllable_BtoR_REQ0 & ~n11333;
  assign n11335 = ~i_RtoB_ACK0 & ~n11334;
  assign n11336 = ~n11332 & ~n11335;
  assign n11337 = ~controllable_DEQ & ~n11336;
  assign n11338 = ~n11323 & ~n11337;
  assign n11339 = i_nEMPTY & ~n11338;
  assign n11340 = ~controllable_ENQ & ~n8946;
  assign n11341 = i_RtoB_ACK1 & ~n11340;
  assign n11342 = ~controllable_ENQ & ~n9747;
  assign n11343 = ~i_RtoB_ACK1 & ~n11342;
  assign n11344 = ~n11341 & ~n11343;
  assign n11345 = controllable_BtoR_REQ1 & ~n11344;
  assign n11346 = ~n9951 & ~n11345;
  assign n11347 = ~controllable_BtoR_REQ0 & ~n11346;
  assign n11348 = ~controllable_BtoR_REQ0 & ~n11347;
  assign n11349 = ~i_RtoB_ACK0 & ~n11348;
  assign n11350 = ~i_RtoB_ACK0 & ~n11349;
  assign n11351 = controllable_DEQ & ~n11350;
  assign n11352 = ~controllable_BtoR_REQ0 & ~n9717;
  assign n11353 = ~controllable_BtoR_REQ0 & ~n11352;
  assign n11354 = ~i_RtoB_ACK0 & ~n11353;
  assign n11355 = ~n11309 & ~n11354;
  assign n11356 = ~controllable_DEQ & ~n11355;
  assign n11357 = ~n11351 & ~n11356;
  assign n11358 = i_FULL & ~n11357;
  assign n11359 = ~n9973 & ~n11327;
  assign n11360 = ~controllable_BtoR_REQ0 & ~n11359;
  assign n11361 = ~controllable_BtoR_REQ0 & ~n11360;
  assign n11362 = ~i_RtoB_ACK0 & ~n11361;
  assign n11363 = ~i_RtoB_ACK0 & ~n11362;
  assign n11364 = controllable_DEQ & ~n11363;
  assign n11365 = ~n9718 & ~n11313;
  assign n11366 = ~controllable_BtoR_REQ1 & ~n11365;
  assign n11367 = ~n11315 & ~n11366;
  assign n11368 = ~controllable_BtoR_REQ0 & ~n11367;
  assign n11369 = ~controllable_BtoR_REQ0 & ~n11368;
  assign n11370 = ~i_RtoB_ACK0 & ~n11369;
  assign n11371 = ~n11309 & ~n11370;
  assign n11372 = ~controllable_DEQ & ~n11371;
  assign n11373 = ~n11364 & ~n11372;
  assign n11374 = ~i_FULL & ~n11373;
  assign n11375 = ~n11358 & ~n11374;
  assign n11376 = ~i_nEMPTY & ~n11375;
  assign n11377 = ~n11339 & ~n11376;
  assign n11378 = ~controllable_BtoS_ACK0 & ~n11377;
  assign n11379 = ~n11296 & ~n11378;
  assign n11380 = ~i_StoB_REQ10 & ~n11379;
  assign n11381 = ~n11224 & ~n11380;
  assign n11382 = controllable_BtoS_ACK10 & ~n11381;
  assign n11383 = ~i_StoB_REQ14 & ~n7894;
  assign n11384 = ~n7690 & ~n11383;
  assign n11385 = controllable_BtoS_ACK14 & ~n11384;
  assign n11386 = ~controllable_BtoS_ACK14 & ~n7894;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = controllable_ENQ & ~n11387;
  assign n11389 = controllable_ENQ & ~n11388;
  assign n11390 = ~i_RtoB_ACK1 & ~n11389;
  assign n11391 = ~n5237 & ~n11390;
  assign n11392 = controllable_BtoR_REQ1 & ~n11391;
  assign n11393 = ~controllable_BtoR_REQ1 & ~n11389;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = ~controllable_BtoR_REQ0 & ~n11394;
  assign n11396 = ~controllable_BtoR_REQ0 & ~n11395;
  assign n11397 = i_RtoB_ACK0 & ~n11396;
  assign n11398 = ~i_StoB_REQ14 & ~n7923;
  assign n11399 = ~n7690 & ~n11398;
  assign n11400 = controllable_BtoS_ACK14 & ~n11399;
  assign n11401 = ~n7924 & ~n11400;
  assign n11402 = controllable_ENQ & ~n11401;
  assign n11403 = ~n5271 & ~n11402;
  assign n11404 = i_RtoB_ACK1 & ~n11403;
  assign n11405 = ~controllable_ENQ & ~n11387;
  assign n11406 = ~n11402 & ~n11405;
  assign n11407 = ~i_RtoB_ACK1 & ~n11406;
  assign n11408 = ~n11404 & ~n11407;
  assign n11409 = controllable_BtoR_REQ1 & ~n11408;
  assign n11410 = i_RtoB_ACK1 & ~n11389;
  assign n11411 = ~n11407 & ~n11410;
  assign n11412 = ~controllable_BtoR_REQ1 & ~n11411;
  assign n11413 = ~n11409 & ~n11412;
  assign n11414 = ~controllable_BtoR_REQ0 & ~n11413;
  assign n11415 = ~controllable_BtoR_REQ0 & ~n11414;
  assign n11416 = ~i_RtoB_ACK0 & ~n11415;
  assign n11417 = ~n11397 & ~n11416;
  assign n11418 = controllable_DEQ & ~n11417;
  assign n11419 = ~i_RtoB_ACK1 & ~n11387;
  assign n11420 = ~n7563 & ~n11419;
  assign n11421 = controllable_BtoR_REQ1 & ~n11420;
  assign n11422 = ~controllable_BtoR_REQ1 & ~n11387;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = ~controllable_BtoR_REQ0 & ~n11423;
  assign n11425 = ~controllable_BtoR_REQ0 & ~n11424;
  assign n11426 = i_RtoB_ACK0 & ~n11425;
  assign n11427 = controllable_BtoR_REQ1 & ~n11401;
  assign n11428 = i_RtoB_ACK1 & ~n11387;
  assign n11429 = ~i_RtoB_ACK1 & ~n11401;
  assign n11430 = ~n11428 & ~n11429;
  assign n11431 = ~controllable_BtoR_REQ1 & ~n11430;
  assign n11432 = ~n11427 & ~n11431;
  assign n11433 = ~controllable_BtoR_REQ0 & ~n11432;
  assign n11434 = ~controllable_BtoR_REQ0 & ~n11433;
  assign n11435 = ~i_RtoB_ACK0 & ~n11434;
  assign n11436 = ~n11426 & ~n11435;
  assign n11437 = ~controllable_DEQ & ~n11436;
  assign n11438 = ~n11418 & ~n11437;
  assign n11439 = i_FULL & ~n11438;
  assign n11440 = ~n5271 & ~n11388;
  assign n11441 = i_RtoB_ACK1 & ~n11440;
  assign n11442 = ~n11419 & ~n11441;
  assign n11443 = controllable_BtoR_REQ1 & ~n11442;
  assign n11444 = ~n11410 & ~n11419;
  assign n11445 = ~controllable_BtoR_REQ1 & ~n11444;
  assign n11446 = ~n11443 & ~n11445;
  assign n11447 = ~controllable_BtoR_REQ0 & ~n11446;
  assign n11448 = ~controllable_BtoR_REQ0 & ~n11447;
  assign n11449 = ~i_RtoB_ACK0 & ~n11448;
  assign n11450 = ~n11397 & ~n11449;
  assign n11451 = controllable_DEQ & ~n11450;
  assign n11452 = controllable_BtoR_REQ1 & ~n11406;
  assign n11453 = ~n11407 & ~n11428;
  assign n11454 = ~controllable_BtoR_REQ1 & ~n11453;
  assign n11455 = ~n11452 & ~n11454;
  assign n11456 = ~controllable_BtoR_REQ0 & ~n11455;
  assign n11457 = ~controllable_BtoR_REQ0 & ~n11456;
  assign n11458 = ~i_RtoB_ACK0 & ~n11457;
  assign n11459 = ~n11426 & ~n11458;
  assign n11460 = ~controllable_DEQ & ~n11459;
  assign n11461 = ~n11451 & ~n11460;
  assign n11462 = ~i_FULL & ~n11461;
  assign n11463 = ~n11439 & ~n11462;
  assign n11464 = i_nEMPTY & ~n11463;
  assign n11465 = ~controllable_ENQ & ~n11405;
  assign n11466 = ~i_RtoB_ACK1 & ~n11465;
  assign n11467 = ~n7574 & ~n11466;
  assign n11468 = controllable_BtoR_REQ1 & ~n11467;
  assign n11469 = ~i_RtoB_ACK1 & ~n11466;
  assign n11470 = ~controllable_BtoR_REQ1 & ~n11469;
  assign n11471 = ~n11468 & ~n11470;
  assign n11472 = ~controllable_BtoR_REQ0 & ~n11471;
  assign n11473 = ~controllable_BtoR_REQ0 & ~n11472;
  assign n11474 = ~i_RtoB_ACK0 & ~n11473;
  assign n11475 = ~i_RtoB_ACK0 & ~n11474;
  assign n11476 = controllable_DEQ & ~n11475;
  assign n11477 = controllable_ENQ & ~n11402;
  assign n11478 = controllable_BtoR_REQ1 & ~n11477;
  assign n11479 = ~i_RtoB_ACK1 & ~n11477;
  assign n11480 = ~n11410 & ~n11479;
  assign n11481 = ~controllable_BtoR_REQ1 & ~n11480;
  assign n11482 = ~n11478 & ~n11481;
  assign n11483 = ~controllable_BtoR_REQ0 & ~n11482;
  assign n11484 = ~controllable_BtoR_REQ0 & ~n11483;
  assign n11485 = ~i_RtoB_ACK0 & ~n11484;
  assign n11486 = ~n11397 & ~n11485;
  assign n11487 = ~controllable_DEQ & ~n11486;
  assign n11488 = ~n11476 & ~n11487;
  assign n11489 = i_FULL & ~n11488;
  assign n11490 = ~i_RtoB_ACK1 & ~n11419;
  assign n11491 = ~controllable_BtoR_REQ1 & ~n11490;
  assign n11492 = ~n11421 & ~n11491;
  assign n11493 = ~controllable_BtoR_REQ0 & ~n11492;
  assign n11494 = ~controllable_BtoR_REQ0 & ~n11493;
  assign n11495 = ~i_RtoB_ACK0 & ~n11494;
  assign n11496 = ~i_RtoB_ACK0 & ~n11495;
  assign n11497 = controllable_DEQ & ~n11496;
  assign n11498 = ~controllable_DEQ & ~n11417;
  assign n11499 = ~n11497 & ~n11498;
  assign n11500 = ~i_FULL & ~n11499;
  assign n11501 = ~n11489 & ~n11500;
  assign n11502 = ~i_nEMPTY & ~n11501;
  assign n11503 = ~n11464 & ~n11502;
  assign n11504 = controllable_BtoS_ACK0 & ~n11503;
  assign n11505 = ~i_StoB_REQ14 & ~n7205;
  assign n11506 = ~n5322 & ~n11505;
  assign n11507 = controllable_BtoS_ACK14 & ~n11506;
  assign n11508 = ~controllable_BtoS_ACK14 & ~n7205;
  assign n11509 = ~n11507 & ~n11508;
  assign n11510 = controllable_ENQ & ~n11509;
  assign n11511 = controllable_ENQ & ~n11510;
  assign n11512 = ~i_RtoB_ACK1 & ~n11511;
  assign n11513 = ~n8861 & ~n11512;
  assign n11514 = controllable_BtoR_REQ1 & ~n11513;
  assign n11515 = ~controllable_BtoR_REQ1 & ~n11511;
  assign n11516 = ~n11514 & ~n11515;
  assign n11517 = ~controllable_BtoR_REQ0 & ~n11516;
  assign n11518 = ~controllable_BtoR_REQ0 & ~n11517;
  assign n11519 = i_RtoB_ACK0 & ~n11518;
  assign n11520 = ~n7256 & ~n8864;
  assign n11521 = i_RtoB_ACK1 & ~n11520;
  assign n11522 = ~controllable_ENQ & ~n11509;
  assign n11523 = ~n7256 & ~n11522;
  assign n11524 = ~i_RtoB_ACK1 & ~n11523;
  assign n11525 = ~n11521 & ~n11524;
  assign n11526 = controllable_BtoR_REQ1 & ~n11525;
  assign n11527 = i_RtoB_ACK1 & ~n11511;
  assign n11528 = ~n11524 & ~n11527;
  assign n11529 = ~controllable_BtoR_REQ1 & ~n11528;
  assign n11530 = ~n11526 & ~n11529;
  assign n11531 = ~controllable_BtoR_REQ0 & ~n11530;
  assign n11532 = ~controllable_BtoR_REQ0 & ~n11531;
  assign n11533 = ~i_RtoB_ACK0 & ~n11532;
  assign n11534 = ~n11519 & ~n11533;
  assign n11535 = controllable_DEQ & ~n11534;
  assign n11536 = ~i_RtoB_ACK1 & ~n11509;
  assign n11537 = ~n8883 & ~n11536;
  assign n11538 = controllable_BtoR_REQ1 & ~n11537;
  assign n11539 = ~controllable_BtoR_REQ1 & ~n11509;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~controllable_BtoR_REQ0 & ~n11540;
  assign n11542 = ~controllable_BtoR_REQ0 & ~n11541;
  assign n11543 = i_RtoB_ACK0 & ~n11542;
  assign n11544 = i_RtoB_ACK1 & ~n11509;
  assign n11545 = ~n7288 & ~n11544;
  assign n11546 = ~controllable_BtoR_REQ1 & ~n11545;
  assign n11547 = ~n7286 & ~n11546;
  assign n11548 = ~controllable_BtoR_REQ0 & ~n11547;
  assign n11549 = ~controllable_BtoR_REQ0 & ~n11548;
  assign n11550 = ~i_RtoB_ACK0 & ~n11549;
  assign n11551 = ~n11543 & ~n11550;
  assign n11552 = ~controllable_DEQ & ~n11551;
  assign n11553 = ~n11535 & ~n11552;
  assign n11554 = i_FULL & ~n11553;
  assign n11555 = ~n8864 & ~n11510;
  assign n11556 = i_RtoB_ACK1 & ~n11555;
  assign n11557 = ~n11536 & ~n11556;
  assign n11558 = controllable_BtoR_REQ1 & ~n11557;
  assign n11559 = ~n11527 & ~n11536;
  assign n11560 = ~controllable_BtoR_REQ1 & ~n11559;
  assign n11561 = ~n11558 & ~n11560;
  assign n11562 = ~controllable_BtoR_REQ0 & ~n11561;
  assign n11563 = ~controllable_BtoR_REQ0 & ~n11562;
  assign n11564 = ~i_RtoB_ACK0 & ~n11563;
  assign n11565 = ~n11519 & ~n11564;
  assign n11566 = controllable_DEQ & ~n11565;
  assign n11567 = controllable_BtoR_REQ1 & ~n11523;
  assign n11568 = ~n11524 & ~n11544;
  assign n11569 = ~controllable_BtoR_REQ1 & ~n11568;
  assign n11570 = ~n11567 & ~n11569;
  assign n11571 = ~controllable_BtoR_REQ0 & ~n11570;
  assign n11572 = ~controllable_BtoR_REQ0 & ~n11571;
  assign n11573 = ~i_RtoB_ACK0 & ~n11572;
  assign n11574 = ~n11543 & ~n11573;
  assign n11575 = ~controllable_DEQ & ~n11574;
  assign n11576 = ~n11566 & ~n11575;
  assign n11577 = ~i_FULL & ~n11576;
  assign n11578 = ~n11554 & ~n11577;
  assign n11579 = i_nEMPTY & ~n11578;
  assign n11580 = i_RtoB_ACK1 & ~n8914;
  assign n11581 = ~controllable_ENQ & ~n11522;
  assign n11582 = ~i_RtoB_ACK1 & ~n11581;
  assign n11583 = ~n11580 & ~n11582;
  assign n11584 = controllable_BtoR_REQ1 & ~n11583;
  assign n11585 = ~i_RtoB_ACK1 & ~n11582;
  assign n11586 = ~controllable_BtoR_REQ1 & ~n11585;
  assign n11587 = ~n11584 & ~n11586;
  assign n11588 = ~controllable_BtoR_REQ0 & ~n11587;
  assign n11589 = ~controllable_BtoR_REQ0 & ~n11588;
  assign n11590 = ~i_RtoB_ACK0 & ~n11589;
  assign n11591 = ~i_RtoB_ACK0 & ~n11590;
  assign n11592 = controllable_DEQ & ~n11591;
  assign n11593 = ~n7345 & ~n11527;
  assign n11594 = ~controllable_BtoR_REQ1 & ~n11593;
  assign n11595 = ~n7344 & ~n11594;
  assign n11596 = ~controllable_BtoR_REQ0 & ~n11595;
  assign n11597 = ~controllable_BtoR_REQ0 & ~n11596;
  assign n11598 = ~i_RtoB_ACK0 & ~n11597;
  assign n11599 = ~n11519 & ~n11598;
  assign n11600 = ~controllable_DEQ & ~n11599;
  assign n11601 = ~n11592 & ~n11600;
  assign n11602 = i_FULL & ~n11601;
  assign n11603 = ~i_RtoB_ACK1 & ~n11536;
  assign n11604 = ~controllable_BtoR_REQ1 & ~n11603;
  assign n11605 = ~n11538 & ~n11604;
  assign n11606 = ~controllable_BtoR_REQ0 & ~n11605;
  assign n11607 = ~controllable_BtoR_REQ0 & ~n11606;
  assign n11608 = ~i_RtoB_ACK0 & ~n11607;
  assign n11609 = ~i_RtoB_ACK0 & ~n11608;
  assign n11610 = controllable_DEQ & ~n11609;
  assign n11611 = ~controllable_DEQ & ~n11534;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = ~i_FULL & ~n11612;
  assign n11614 = ~n11602 & ~n11613;
  assign n11615 = ~i_nEMPTY & ~n11614;
  assign n11616 = ~n11579 & ~n11615;
  assign n11617 = ~controllable_BtoS_ACK0 & ~n11616;
  assign n11618 = ~n11504 & ~n11617;
  assign n11619 = n4465 & ~n11618;
  assign n11620 = ~n7599 & ~n11617;
  assign n11621 = ~n4465 & ~n11620;
  assign n11622 = ~n11619 & ~n11621;
  assign n11623 = i_StoB_REQ10 & ~n11622;
  assign n11624 = ~i_StoB_REQ14 & ~n7880;
  assign n11625 = controllable_BtoS_ACK14 & ~n11624;
  assign n11626 = i_StoB_REQ14 & ~n8454;
  assign n11627 = ~n7880 & ~n11626;
  assign n11628 = ~controllable_BtoS_ACK14 & ~n11627;
  assign n11629 = ~n11625 & ~n11628;
  assign n11630 = controllable_ENQ & ~n11629;
  assign n11631 = controllable_ENQ & ~n11630;
  assign n11632 = i_RtoB_ACK1 & ~n11631;
  assign n11633 = ~n7887 & ~n7897;
  assign n11634 = controllable_BtoS_ACK14 & ~n11633;
  assign n11635 = i_StoB_REQ14 & ~n7910;
  assign n11636 = ~n7897 & ~n11635;
  assign n11637 = ~controllable_BtoS_ACK14 & ~n11636;
  assign n11638 = ~n11634 & ~n11637;
  assign n11639 = controllable_ENQ & ~n11638;
  assign n11640 = controllable_ENQ & ~n11639;
  assign n11641 = ~i_RtoB_ACK1 & ~n11640;
  assign n11642 = ~n11632 & ~n11641;
  assign n11643 = controllable_BtoR_REQ1 & ~n11642;
  assign n11644 = ~n7690 & ~n7911;
  assign n11645 = controllable_BtoS_ACK14 & ~n11644;
  assign n11646 = ~controllable_BtoS_ACK14 & ~n7910;
  assign n11647 = ~n11645 & ~n11646;
  assign n11648 = controllable_ENQ & ~n11647;
  assign n11649 = controllable_ENQ & ~n11648;
  assign n11650 = ~controllable_BtoR_REQ1 & ~n11649;
  assign n11651 = ~n11643 & ~n11650;
  assign n11652 = ~controllable_BtoR_REQ0 & ~n11651;
  assign n11653 = ~controllable_BtoR_REQ0 & ~n11652;
  assign n11654 = i_RtoB_ACK0 & ~n11653;
  assign n11655 = ~controllable_ENQ & ~n11629;
  assign n11656 = ~n11402 & ~n11655;
  assign n11657 = i_RtoB_ACK1 & ~n11656;
  assign n11658 = ~controllable_ENQ & ~n11638;
  assign n11659 = ~n11402 & ~n11658;
  assign n11660 = ~i_RtoB_ACK1 & ~n11659;
  assign n11661 = ~n11657 & ~n11660;
  assign n11662 = controllable_BtoR_REQ1 & ~n11661;
  assign n11663 = i_RtoB_ACK1 & ~n11649;
  assign n11664 = ~controllable_ENQ & ~n11647;
  assign n11665 = ~n11402 & ~n11664;
  assign n11666 = ~i_RtoB_ACK1 & ~n11665;
  assign n11667 = ~n11663 & ~n11666;
  assign n11668 = ~controllable_BtoR_REQ1 & ~n11667;
  assign n11669 = ~n11662 & ~n11668;
  assign n11670 = ~controllable_BtoR_REQ0 & ~n11669;
  assign n11671 = ~controllable_BtoR_REQ0 & ~n11670;
  assign n11672 = ~i_RtoB_ACK0 & ~n11671;
  assign n11673 = ~n11654 & ~n11672;
  assign n11674 = controllable_DEQ & ~n11673;
  assign n11675 = i_RtoB_ACK1 & ~n11629;
  assign n11676 = ~i_RtoB_ACK1 & ~n11638;
  assign n11677 = ~n11675 & ~n11676;
  assign n11678 = controllable_BtoR_REQ1 & ~n11677;
  assign n11679 = ~controllable_BtoR_REQ1 & ~n11647;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~controllable_BtoR_REQ0 & ~n11680;
  assign n11682 = ~controllable_BtoR_REQ0 & ~n11681;
  assign n11683 = i_RtoB_ACK0 & ~n11682;
  assign n11684 = i_RtoB_ACK1 & ~n11647;
  assign n11685 = ~n11429 & ~n11684;
  assign n11686 = ~controllable_BtoR_REQ1 & ~n11685;
  assign n11687 = ~n11427 & ~n11686;
  assign n11688 = ~controllable_BtoR_REQ0 & ~n11687;
  assign n11689 = ~controllable_BtoR_REQ0 & ~n11688;
  assign n11690 = ~i_RtoB_ACK0 & ~n11689;
  assign n11691 = ~n11683 & ~n11690;
  assign n11692 = ~controllable_DEQ & ~n11691;
  assign n11693 = ~n11674 & ~n11692;
  assign n11694 = i_FULL & ~n11693;
  assign n11695 = ~n11648 & ~n11655;
  assign n11696 = i_RtoB_ACK1 & ~n11695;
  assign n11697 = ~n11648 & ~n11658;
  assign n11698 = ~i_RtoB_ACK1 & ~n11697;
  assign n11699 = ~n11696 & ~n11698;
  assign n11700 = controllable_BtoR_REQ1 & ~n11699;
  assign n11701 = ~i_RtoB_ACK1 & ~n11647;
  assign n11702 = ~n11663 & ~n11701;
  assign n11703 = ~controllable_BtoR_REQ1 & ~n11702;
  assign n11704 = ~n11700 & ~n11703;
  assign n11705 = ~controllable_BtoR_REQ0 & ~n11704;
  assign n11706 = ~controllable_BtoR_REQ0 & ~n11705;
  assign n11707 = ~i_RtoB_ACK0 & ~n11706;
  assign n11708 = ~n11654 & ~n11707;
  assign n11709 = controllable_DEQ & ~n11708;
  assign n11710 = controllable_BtoR_REQ1 & ~n11665;
  assign n11711 = ~n11666 & ~n11684;
  assign n11712 = ~controllable_BtoR_REQ1 & ~n11711;
  assign n11713 = ~n11710 & ~n11712;
  assign n11714 = ~controllable_BtoR_REQ0 & ~n11713;
  assign n11715 = ~controllable_BtoR_REQ0 & ~n11714;
  assign n11716 = ~i_RtoB_ACK0 & ~n11715;
  assign n11717 = ~n11683 & ~n11716;
  assign n11718 = ~controllable_DEQ & ~n11717;
  assign n11719 = ~n11709 & ~n11718;
  assign n11720 = ~i_FULL & ~n11719;
  assign n11721 = ~n11694 & ~n11720;
  assign n11722 = i_nEMPTY & ~n11721;
  assign n11723 = ~controllable_ENQ & ~n11655;
  assign n11724 = i_RtoB_ACK1 & ~n11723;
  assign n11725 = ~controllable_ENQ & ~n11658;
  assign n11726 = ~i_RtoB_ACK1 & ~n11725;
  assign n11727 = ~n11724 & ~n11726;
  assign n11728 = controllable_BtoR_REQ1 & ~n11727;
  assign n11729 = ~controllable_ENQ & ~n11664;
  assign n11730 = ~i_RtoB_ACK1 & ~n11729;
  assign n11731 = ~i_RtoB_ACK1 & ~n11730;
  assign n11732 = ~controllable_BtoR_REQ1 & ~n11731;
  assign n11733 = ~n11728 & ~n11732;
  assign n11734 = ~controllable_BtoR_REQ0 & ~n11733;
  assign n11735 = ~controllable_BtoR_REQ0 & ~n11734;
  assign n11736 = ~i_RtoB_ACK0 & ~n11735;
  assign n11737 = ~i_RtoB_ACK0 & ~n11736;
  assign n11738 = controllable_DEQ & ~n11737;
  assign n11739 = ~n11479 & ~n11663;
  assign n11740 = ~controllable_BtoR_REQ1 & ~n11739;
  assign n11741 = ~n11478 & ~n11740;
  assign n11742 = ~controllable_BtoR_REQ0 & ~n11741;
  assign n11743 = ~controllable_BtoR_REQ0 & ~n11742;
  assign n11744 = ~i_RtoB_ACK0 & ~n11743;
  assign n11745 = ~n11654 & ~n11744;
  assign n11746 = ~controllable_DEQ & ~n11745;
  assign n11747 = ~n11738 & ~n11746;
  assign n11748 = i_FULL & ~n11747;
  assign n11749 = ~i_RtoB_ACK1 & ~n11701;
  assign n11750 = ~controllable_BtoR_REQ1 & ~n11749;
  assign n11751 = ~n11678 & ~n11750;
  assign n11752 = ~controllable_BtoR_REQ0 & ~n11751;
  assign n11753 = ~controllable_BtoR_REQ0 & ~n11752;
  assign n11754 = ~i_RtoB_ACK0 & ~n11753;
  assign n11755 = ~i_RtoB_ACK0 & ~n11754;
  assign n11756 = controllable_DEQ & ~n11755;
  assign n11757 = ~n11660 & ~n11663;
  assign n11758 = ~controllable_BtoR_REQ1 & ~n11757;
  assign n11759 = ~n11662 & ~n11758;
  assign n11760 = ~controllable_BtoR_REQ0 & ~n11759;
  assign n11761 = ~controllable_BtoR_REQ0 & ~n11760;
  assign n11762 = ~i_RtoB_ACK0 & ~n11761;
  assign n11763 = ~n11654 & ~n11762;
  assign n11764 = ~controllable_DEQ & ~n11763;
  assign n11765 = ~n11756 & ~n11764;
  assign n11766 = ~i_FULL & ~n11765;
  assign n11767 = ~n11748 & ~n11766;
  assign n11768 = ~i_nEMPTY & ~n11767;
  assign n11769 = ~n11722 & ~n11768;
  assign n11770 = controllable_BtoS_ACK0 & ~n11769;
  assign n11771 = ~i_StoB_REQ14 & ~n8051;
  assign n11772 = controllable_BtoS_ACK14 & ~n11771;
  assign n11773 = i_StoB_REQ14 & ~n7187;
  assign n11774 = ~n8051 & ~n11773;
  assign n11775 = ~controllable_BtoS_ACK14 & ~n11774;
  assign n11776 = ~n11772 & ~n11775;
  assign n11777 = controllable_ENQ & ~n11776;
  assign n11778 = controllable_ENQ & ~n11777;
  assign n11779 = i_RtoB_ACK1 & ~n11778;
  assign n11780 = ~n7197 & ~n8066;
  assign n11781 = controllable_BtoS_ACK14 & ~n11780;
  assign n11782 = i_StoB_REQ14 & ~n7223;
  assign n11783 = ~n8066 & ~n11782;
  assign n11784 = ~controllable_BtoS_ACK14 & ~n11783;
  assign n11785 = ~n11781 & ~n11784;
  assign n11786 = controllable_ENQ & ~n11785;
  assign n11787 = controllable_ENQ & ~n11786;
  assign n11788 = ~i_RtoB_ACK1 & ~n11787;
  assign n11789 = ~n11779 & ~n11788;
  assign n11790 = controllable_BtoR_REQ1 & ~n11789;
  assign n11791 = ~n5322 & ~n8078;
  assign n11792 = controllable_BtoS_ACK14 & ~n11791;
  assign n11793 = ~controllable_BtoS_ACK14 & ~n7223;
  assign n11794 = ~n11792 & ~n11793;
  assign n11795 = controllable_ENQ & ~n11794;
  assign n11796 = controllable_ENQ & ~n11795;
  assign n11797 = ~controllable_BtoR_REQ1 & ~n11796;
  assign n11798 = ~n11790 & ~n11797;
  assign n11799 = ~controllable_BtoR_REQ0 & ~n11798;
  assign n11800 = ~controllable_BtoR_REQ0 & ~n11799;
  assign n11801 = i_RtoB_ACK0 & ~n11800;
  assign n11802 = ~controllable_ENQ & ~n11776;
  assign n11803 = ~n7256 & ~n11802;
  assign n11804 = i_RtoB_ACK1 & ~n11803;
  assign n11805 = ~controllable_ENQ & ~n11785;
  assign n11806 = ~n7256 & ~n11805;
  assign n11807 = ~i_RtoB_ACK1 & ~n11806;
  assign n11808 = ~n11804 & ~n11807;
  assign n11809 = controllable_BtoR_REQ1 & ~n11808;
  assign n11810 = i_RtoB_ACK1 & ~n11796;
  assign n11811 = ~controllable_ENQ & ~n11794;
  assign n11812 = ~n7256 & ~n11811;
  assign n11813 = ~i_RtoB_ACK1 & ~n11812;
  assign n11814 = ~n11810 & ~n11813;
  assign n11815 = ~controllable_BtoR_REQ1 & ~n11814;
  assign n11816 = ~n11809 & ~n11815;
  assign n11817 = ~controllable_BtoR_REQ0 & ~n11816;
  assign n11818 = ~controllable_BtoR_REQ0 & ~n11817;
  assign n11819 = ~i_RtoB_ACK0 & ~n11818;
  assign n11820 = ~n11801 & ~n11819;
  assign n11821 = controllable_DEQ & ~n11820;
  assign n11822 = i_RtoB_ACK1 & ~n11776;
  assign n11823 = ~i_RtoB_ACK1 & ~n11785;
  assign n11824 = ~n11822 & ~n11823;
  assign n11825 = controllable_BtoR_REQ1 & ~n11824;
  assign n11826 = ~controllable_BtoR_REQ1 & ~n11794;
  assign n11827 = ~n11825 & ~n11826;
  assign n11828 = ~controllable_BtoR_REQ0 & ~n11827;
  assign n11829 = ~controllable_BtoR_REQ0 & ~n11828;
  assign n11830 = i_RtoB_ACK0 & ~n11829;
  assign n11831 = i_RtoB_ACK1 & ~n11794;
  assign n11832 = ~n7288 & ~n11831;
  assign n11833 = ~controllable_BtoR_REQ1 & ~n11832;
  assign n11834 = ~n7286 & ~n11833;
  assign n11835 = ~controllable_BtoR_REQ0 & ~n11834;
  assign n11836 = ~controllable_BtoR_REQ0 & ~n11835;
  assign n11837 = ~i_RtoB_ACK0 & ~n11836;
  assign n11838 = ~n11830 & ~n11837;
  assign n11839 = ~controllable_DEQ & ~n11838;
  assign n11840 = ~n11821 & ~n11839;
  assign n11841 = i_FULL & ~n11840;
  assign n11842 = ~n11795 & ~n11802;
  assign n11843 = i_RtoB_ACK1 & ~n11842;
  assign n11844 = ~n11795 & ~n11805;
  assign n11845 = ~i_RtoB_ACK1 & ~n11844;
  assign n11846 = ~n11843 & ~n11845;
  assign n11847 = controllable_BtoR_REQ1 & ~n11846;
  assign n11848 = ~i_RtoB_ACK1 & ~n11794;
  assign n11849 = ~n11810 & ~n11848;
  assign n11850 = ~controllable_BtoR_REQ1 & ~n11849;
  assign n11851 = ~n11847 & ~n11850;
  assign n11852 = ~controllable_BtoR_REQ0 & ~n11851;
  assign n11853 = ~controllable_BtoR_REQ0 & ~n11852;
  assign n11854 = ~i_RtoB_ACK0 & ~n11853;
  assign n11855 = ~n11801 & ~n11854;
  assign n11856 = controllable_DEQ & ~n11855;
  assign n11857 = controllable_BtoR_REQ1 & ~n11812;
  assign n11858 = ~n11813 & ~n11831;
  assign n11859 = ~controllable_BtoR_REQ1 & ~n11858;
  assign n11860 = ~n11857 & ~n11859;
  assign n11861 = ~controllable_BtoR_REQ0 & ~n11860;
  assign n11862 = ~controllable_BtoR_REQ0 & ~n11861;
  assign n11863 = ~i_RtoB_ACK0 & ~n11862;
  assign n11864 = ~n11830 & ~n11863;
  assign n11865 = ~controllable_DEQ & ~n11864;
  assign n11866 = ~n11856 & ~n11865;
  assign n11867 = ~i_FULL & ~n11866;
  assign n11868 = ~n11841 & ~n11867;
  assign n11869 = i_nEMPTY & ~n11868;
  assign n11870 = ~controllable_ENQ & ~n11802;
  assign n11871 = i_RtoB_ACK1 & ~n11870;
  assign n11872 = ~controllable_ENQ & ~n11805;
  assign n11873 = ~i_RtoB_ACK1 & ~n11872;
  assign n11874 = ~n11871 & ~n11873;
  assign n11875 = controllable_BtoR_REQ1 & ~n11874;
  assign n11876 = ~controllable_ENQ & ~n11811;
  assign n11877 = ~i_RtoB_ACK1 & ~n11876;
  assign n11878 = ~i_RtoB_ACK1 & ~n11877;
  assign n11879 = ~controllable_BtoR_REQ1 & ~n11878;
  assign n11880 = ~n11875 & ~n11879;
  assign n11881 = ~controllable_BtoR_REQ0 & ~n11880;
  assign n11882 = ~controllable_BtoR_REQ0 & ~n11881;
  assign n11883 = ~i_RtoB_ACK0 & ~n11882;
  assign n11884 = ~i_RtoB_ACK0 & ~n11883;
  assign n11885 = controllable_DEQ & ~n11884;
  assign n11886 = ~n7345 & ~n11810;
  assign n11887 = ~controllable_BtoR_REQ1 & ~n11886;
  assign n11888 = ~n7344 & ~n11887;
  assign n11889 = ~controllable_BtoR_REQ0 & ~n11888;
  assign n11890 = ~controllable_BtoR_REQ0 & ~n11889;
  assign n11891 = ~i_RtoB_ACK0 & ~n11890;
  assign n11892 = ~n11801 & ~n11891;
  assign n11893 = ~controllable_DEQ & ~n11892;
  assign n11894 = ~n11885 & ~n11893;
  assign n11895 = i_FULL & ~n11894;
  assign n11896 = ~i_RtoB_ACK1 & ~n11848;
  assign n11897 = ~controllable_BtoR_REQ1 & ~n11896;
  assign n11898 = ~n11825 & ~n11897;
  assign n11899 = ~controllable_BtoR_REQ0 & ~n11898;
  assign n11900 = ~controllable_BtoR_REQ0 & ~n11899;
  assign n11901 = ~i_RtoB_ACK0 & ~n11900;
  assign n11902 = ~i_RtoB_ACK0 & ~n11901;
  assign n11903 = controllable_DEQ & ~n11902;
  assign n11904 = ~n11807 & ~n11810;
  assign n11905 = ~controllable_BtoR_REQ1 & ~n11904;
  assign n11906 = ~n11809 & ~n11905;
  assign n11907 = ~controllable_BtoR_REQ0 & ~n11906;
  assign n11908 = ~controllable_BtoR_REQ0 & ~n11907;
  assign n11909 = ~i_RtoB_ACK0 & ~n11908;
  assign n11910 = ~n11801 & ~n11909;
  assign n11911 = ~controllable_DEQ & ~n11910;
  assign n11912 = ~n11903 & ~n11911;
  assign n11913 = ~i_FULL & ~n11912;
  assign n11914 = ~n11895 & ~n11913;
  assign n11915 = ~i_nEMPTY & ~n11914;
  assign n11916 = ~n11869 & ~n11915;
  assign n11917 = ~controllable_BtoS_ACK0 & ~n11916;
  assign n11918 = ~n11770 & ~n11917;
  assign n11919 = n4465 & ~n11918;
  assign n11920 = ~n7379 & ~n11919;
  assign n11921 = ~i_StoB_REQ10 & ~n11920;
  assign n11922 = ~n11623 & ~n11921;
  assign n11923 = ~controllable_BtoS_ACK10 & ~n11922;
  assign n11924 = ~n11382 & ~n11923;
  assign n11925 = n4464 & ~n11924;
  assign n11926 = ~n7878 & ~n11380;
  assign n11927 = controllable_BtoS_ACK10 & ~n11926;
  assign n11928 = ~n7909 & ~n11386;
  assign n11929 = controllable_ENQ & ~n11928;
  assign n11930 = controllable_ENQ & ~n11929;
  assign n11931 = ~i_RtoB_ACK1 & ~n11930;
  assign n11932 = ~n5237 & ~n11931;
  assign n11933 = controllable_BtoR_REQ1 & ~n11932;
  assign n11934 = ~controllable_BtoR_REQ1 & ~n11930;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = ~controllable_BtoR_REQ0 & ~n11935;
  assign n11937 = ~controllable_BtoR_REQ0 & ~n11936;
  assign n11938 = i_RtoB_ACK0 & ~n11937;
  assign n11939 = ~n5271 & ~n7926;
  assign n11940 = i_RtoB_ACK1 & ~n11939;
  assign n11941 = ~controllable_ENQ & ~n11928;
  assign n11942 = ~n7926 & ~n11941;
  assign n11943 = ~i_RtoB_ACK1 & ~n11942;
  assign n11944 = ~n11940 & ~n11943;
  assign n11945 = controllable_BtoR_REQ1 & ~n11944;
  assign n11946 = i_RtoB_ACK1 & ~n11930;
  assign n11947 = ~n11943 & ~n11946;
  assign n11948 = ~controllable_BtoR_REQ1 & ~n11947;
  assign n11949 = ~n11945 & ~n11948;
  assign n11950 = ~controllable_BtoR_REQ0 & ~n11949;
  assign n11951 = ~controllable_BtoR_REQ0 & ~n11950;
  assign n11952 = ~i_RtoB_ACK0 & ~n11951;
  assign n11953 = ~n11938 & ~n11952;
  assign n11954 = controllable_DEQ & ~n11953;
  assign n11955 = ~i_RtoB_ACK1 & ~n11928;
  assign n11956 = ~n7563 & ~n11955;
  assign n11957 = controllable_BtoR_REQ1 & ~n11956;
  assign n11958 = ~controllable_BtoR_REQ1 & ~n11928;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = ~controllable_BtoR_REQ0 & ~n11959;
  assign n11961 = ~controllable_BtoR_REQ0 & ~n11960;
  assign n11962 = i_RtoB_ACK0 & ~n11961;
  assign n11963 = i_RtoB_ACK1 & ~n11928;
  assign n11964 = ~n7958 & ~n11963;
  assign n11965 = ~controllable_BtoR_REQ1 & ~n11964;
  assign n11966 = ~n7956 & ~n11965;
  assign n11967 = ~controllable_BtoR_REQ0 & ~n11966;
  assign n11968 = ~controllable_BtoR_REQ0 & ~n11967;
  assign n11969 = ~i_RtoB_ACK0 & ~n11968;
  assign n11970 = ~n11962 & ~n11969;
  assign n11971 = ~controllable_DEQ & ~n11970;
  assign n11972 = ~n11954 & ~n11971;
  assign n11973 = i_FULL & ~n11972;
  assign n11974 = ~n5271 & ~n11929;
  assign n11975 = i_RtoB_ACK1 & ~n11974;
  assign n11976 = ~n11955 & ~n11975;
  assign n11977 = controllable_BtoR_REQ1 & ~n11976;
  assign n11978 = ~n11946 & ~n11955;
  assign n11979 = ~controllable_BtoR_REQ1 & ~n11978;
  assign n11980 = ~n11977 & ~n11979;
  assign n11981 = ~controllable_BtoR_REQ0 & ~n11980;
  assign n11982 = ~controllable_BtoR_REQ0 & ~n11981;
  assign n11983 = ~i_RtoB_ACK0 & ~n11982;
  assign n11984 = ~n11938 & ~n11983;
  assign n11985 = controllable_DEQ & ~n11984;
  assign n11986 = controllable_BtoR_REQ1 & ~n11942;
  assign n11987 = ~n11943 & ~n11963;
  assign n11988 = ~controllable_BtoR_REQ1 & ~n11987;
  assign n11989 = ~n11986 & ~n11988;
  assign n11990 = ~controllable_BtoR_REQ0 & ~n11989;
  assign n11991 = ~controllable_BtoR_REQ0 & ~n11990;
  assign n11992 = ~i_RtoB_ACK0 & ~n11991;
  assign n11993 = ~n11962 & ~n11992;
  assign n11994 = ~controllable_DEQ & ~n11993;
  assign n11995 = ~n11985 & ~n11994;
  assign n11996 = ~i_FULL & ~n11995;
  assign n11997 = ~n11973 & ~n11996;
  assign n11998 = i_nEMPTY & ~n11997;
  assign n11999 = ~controllable_ENQ & ~n11941;
  assign n12000 = ~i_RtoB_ACK1 & ~n11999;
  assign n12001 = ~n7574 & ~n12000;
  assign n12002 = controllable_BtoR_REQ1 & ~n12001;
  assign n12003 = ~i_RtoB_ACK1 & ~n12000;
  assign n12004 = ~controllable_BtoR_REQ1 & ~n12003;
  assign n12005 = ~n12002 & ~n12004;
  assign n12006 = ~controllable_BtoR_REQ0 & ~n12005;
  assign n12007 = ~controllable_BtoR_REQ0 & ~n12006;
  assign n12008 = ~i_RtoB_ACK0 & ~n12007;
  assign n12009 = ~i_RtoB_ACK0 & ~n12008;
  assign n12010 = controllable_DEQ & ~n12009;
  assign n12011 = ~n8015 & ~n11946;
  assign n12012 = ~controllable_BtoR_REQ1 & ~n12011;
  assign n12013 = ~n8014 & ~n12012;
  assign n12014 = ~controllable_BtoR_REQ0 & ~n12013;
  assign n12015 = ~controllable_BtoR_REQ0 & ~n12014;
  assign n12016 = ~i_RtoB_ACK0 & ~n12015;
  assign n12017 = ~n11938 & ~n12016;
  assign n12018 = ~controllable_DEQ & ~n12017;
  assign n12019 = ~n12010 & ~n12018;
  assign n12020 = i_FULL & ~n12019;
  assign n12021 = ~i_RtoB_ACK1 & ~n11955;
  assign n12022 = ~controllable_BtoR_REQ1 & ~n12021;
  assign n12023 = ~n11957 & ~n12022;
  assign n12024 = ~controllable_BtoR_REQ0 & ~n12023;
  assign n12025 = ~controllable_BtoR_REQ0 & ~n12024;
  assign n12026 = ~i_RtoB_ACK0 & ~n12025;
  assign n12027 = ~i_RtoB_ACK0 & ~n12026;
  assign n12028 = controllable_DEQ & ~n12027;
  assign n12029 = ~controllable_DEQ & ~n11953;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = ~i_FULL & ~n12030;
  assign n12032 = ~n12020 & ~n12031;
  assign n12033 = ~i_nEMPTY & ~n12032;
  assign n12034 = ~n11998 & ~n12033;
  assign n12035 = controllable_BtoS_ACK0 & ~n12034;
  assign n12036 = ~n8077 & ~n11508;
  assign n12037 = controllable_ENQ & ~n12036;
  assign n12038 = controllable_ENQ & ~n12037;
  assign n12039 = ~i_RtoB_ACK1 & ~n12038;
  assign n12040 = ~n8861 & ~n12039;
  assign n12041 = controllable_BtoR_REQ1 & ~n12040;
  assign n12042 = ~controllable_BtoR_REQ1 & ~n12038;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = ~controllable_BtoR_REQ0 & ~n12043;
  assign n12045 = ~controllable_BtoR_REQ0 & ~n12044;
  assign n12046 = i_RtoB_ACK0 & ~n12045;
  assign n12047 = ~n8090 & ~n8864;
  assign n12048 = i_RtoB_ACK1 & ~n12047;
  assign n12049 = ~controllable_ENQ & ~n12036;
  assign n12050 = ~n8090 & ~n12049;
  assign n12051 = ~i_RtoB_ACK1 & ~n12050;
  assign n12052 = ~n12048 & ~n12051;
  assign n12053 = controllable_BtoR_REQ1 & ~n12052;
  assign n12054 = i_RtoB_ACK1 & ~n12038;
  assign n12055 = ~n12051 & ~n12054;
  assign n12056 = ~controllable_BtoR_REQ1 & ~n12055;
  assign n12057 = ~n12053 & ~n12056;
  assign n12058 = ~controllable_BtoR_REQ0 & ~n12057;
  assign n12059 = ~controllable_BtoR_REQ0 & ~n12058;
  assign n12060 = ~i_RtoB_ACK0 & ~n12059;
  assign n12061 = ~n12046 & ~n12060;
  assign n12062 = controllable_DEQ & ~n12061;
  assign n12063 = ~i_RtoB_ACK1 & ~n12036;
  assign n12064 = ~n8883 & ~n12063;
  assign n12065 = controllable_BtoR_REQ1 & ~n12064;
  assign n12066 = ~controllable_BtoR_REQ1 & ~n12036;
  assign n12067 = ~n12065 & ~n12066;
  assign n12068 = ~controllable_BtoR_REQ0 & ~n12067;
  assign n12069 = ~controllable_BtoR_REQ0 & ~n12068;
  assign n12070 = i_RtoB_ACK0 & ~n12069;
  assign n12071 = i_RtoB_ACK1 & ~n12036;
  assign n12072 = ~n8122 & ~n12071;
  assign n12073 = ~controllable_BtoR_REQ1 & ~n12072;
  assign n12074 = ~n8120 & ~n12073;
  assign n12075 = ~controllable_BtoR_REQ0 & ~n12074;
  assign n12076 = ~controllable_BtoR_REQ0 & ~n12075;
  assign n12077 = ~i_RtoB_ACK0 & ~n12076;
  assign n12078 = ~n12070 & ~n12077;
  assign n12079 = ~controllable_DEQ & ~n12078;
  assign n12080 = ~n12062 & ~n12079;
  assign n12081 = i_FULL & ~n12080;
  assign n12082 = ~n8864 & ~n12037;
  assign n12083 = i_RtoB_ACK1 & ~n12082;
  assign n12084 = ~n12063 & ~n12083;
  assign n12085 = controllable_BtoR_REQ1 & ~n12084;
  assign n12086 = ~n12054 & ~n12063;
  assign n12087 = ~controllable_BtoR_REQ1 & ~n12086;
  assign n12088 = ~n12085 & ~n12087;
  assign n12089 = ~controllable_BtoR_REQ0 & ~n12088;
  assign n12090 = ~controllable_BtoR_REQ0 & ~n12089;
  assign n12091 = ~i_RtoB_ACK0 & ~n12090;
  assign n12092 = ~n12046 & ~n12091;
  assign n12093 = controllable_DEQ & ~n12092;
  assign n12094 = controllable_BtoR_REQ1 & ~n12050;
  assign n12095 = ~n12051 & ~n12071;
  assign n12096 = ~controllable_BtoR_REQ1 & ~n12095;
  assign n12097 = ~n12094 & ~n12096;
  assign n12098 = ~controllable_BtoR_REQ0 & ~n12097;
  assign n12099 = ~controllable_BtoR_REQ0 & ~n12098;
  assign n12100 = ~i_RtoB_ACK0 & ~n12099;
  assign n12101 = ~n12070 & ~n12100;
  assign n12102 = ~controllable_DEQ & ~n12101;
  assign n12103 = ~n12093 & ~n12102;
  assign n12104 = ~i_FULL & ~n12103;
  assign n12105 = ~n12081 & ~n12104;
  assign n12106 = i_nEMPTY & ~n12105;
  assign n12107 = ~controllable_ENQ & ~n12049;
  assign n12108 = ~i_RtoB_ACK1 & ~n12107;
  assign n12109 = ~n11580 & ~n12108;
  assign n12110 = controllable_BtoR_REQ1 & ~n12109;
  assign n12111 = ~i_RtoB_ACK1 & ~n12108;
  assign n12112 = ~controllable_BtoR_REQ1 & ~n12111;
  assign n12113 = ~n12110 & ~n12112;
  assign n12114 = ~controllable_BtoR_REQ0 & ~n12113;
  assign n12115 = ~controllable_BtoR_REQ0 & ~n12114;
  assign n12116 = ~i_RtoB_ACK0 & ~n12115;
  assign n12117 = ~i_RtoB_ACK0 & ~n12116;
  assign n12118 = controllable_DEQ & ~n12117;
  assign n12119 = ~n8179 & ~n12054;
  assign n12120 = ~controllable_BtoR_REQ1 & ~n12119;
  assign n12121 = ~n8178 & ~n12120;
  assign n12122 = ~controllable_BtoR_REQ0 & ~n12121;
  assign n12123 = ~controllable_BtoR_REQ0 & ~n12122;
  assign n12124 = ~i_RtoB_ACK0 & ~n12123;
  assign n12125 = ~n12046 & ~n12124;
  assign n12126 = ~controllable_DEQ & ~n12125;
  assign n12127 = ~n12118 & ~n12126;
  assign n12128 = i_FULL & ~n12127;
  assign n12129 = ~i_RtoB_ACK1 & ~n12063;
  assign n12130 = ~controllable_BtoR_REQ1 & ~n12129;
  assign n12131 = ~n12065 & ~n12130;
  assign n12132 = ~controllable_BtoR_REQ0 & ~n12131;
  assign n12133 = ~controllable_BtoR_REQ0 & ~n12132;
  assign n12134 = ~i_RtoB_ACK0 & ~n12133;
  assign n12135 = ~i_RtoB_ACK0 & ~n12134;
  assign n12136 = controllable_DEQ & ~n12135;
  assign n12137 = ~controllable_DEQ & ~n12061;
  assign n12138 = ~n12136 & ~n12137;
  assign n12139 = ~i_FULL & ~n12138;
  assign n12140 = ~n12128 & ~n12139;
  assign n12141 = ~i_nEMPTY & ~n12140;
  assign n12142 = ~n12106 & ~n12141;
  assign n12143 = ~controllable_BtoS_ACK0 & ~n12142;
  assign n12144 = ~n12035 & ~n12143;
  assign n12145 = n4465 & ~n12144;
  assign n12146 = ~n8666 & ~n12143;
  assign n12147 = ~n4465 & ~n12146;
  assign n12148 = ~n12145 & ~n12147;
  assign n12149 = i_StoB_REQ10 & ~n12148;
  assign n12150 = ~n8451 & ~n12149;
  assign n12151 = ~controllable_BtoS_ACK10 & ~n12150;
  assign n12152 = ~n11927 & ~n12151;
  assign n12153 = ~n4464 & ~n12152;
  assign n12154 = ~n11925 & ~n12153;
  assign n12155 = n4463 & ~n12154;
  assign n12156 = ~i_StoB_REQ14 & ~n10453;
  assign n12157 = ~i_StoB_REQ14 & ~n12156;
  assign n12158 = controllable_BtoS_ACK14 & ~n12157;
  assign n12159 = ~n5216 & ~n12156;
  assign n12160 = ~controllable_BtoS_ACK14 & ~n12159;
  assign n12161 = ~n12158 & ~n12160;
  assign n12162 = controllable_ENQ & ~n12161;
  assign n12163 = controllable_ENQ & ~n12162;
  assign n12164 = ~i_RtoB_ACK1 & ~n12163;
  assign n12165 = ~n11150 & ~n12164;
  assign n12166 = ~controllable_BtoR_REQ1 & ~n12165;
  assign n12167 = ~n11138 & ~n12166;
  assign n12168 = ~controllable_BtoR_REQ0 & ~n12167;
  assign n12169 = ~controllable_BtoR_REQ0 & ~n12168;
  assign n12170 = i_RtoB_ACK0 & ~n12169;
  assign n12171 = ~n5237 & ~n11153;
  assign n12172 = controllable_BtoR_REQ1 & ~n12171;
  assign n12173 = ~controllable_ENQ & ~n12161;
  assign n12174 = ~n5230 & ~n12173;
  assign n12175 = ~i_RtoB_ACK1 & ~n12174;
  assign n12176 = ~n11150 & ~n12175;
  assign n12177 = ~controllable_BtoR_REQ1 & ~n12176;
  assign n12178 = ~n12172 & ~n12177;
  assign n12179 = ~controllable_BtoR_REQ0 & ~n12178;
  assign n12180 = ~controllable_BtoR_REQ0 & ~n12179;
  assign n12181 = ~i_RtoB_ACK0 & ~n12180;
  assign n12182 = ~n12170 & ~n12181;
  assign n12183 = controllable_DEQ & ~n12182;
  assign n12184 = i_RtoB_ACK1 & ~n11142;
  assign n12185 = ~i_RtoB_ACK1 & ~n12161;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~controllable_BtoR_REQ1 & ~n12186;
  assign n12188 = ~n11167 & ~n12187;
  assign n12189 = ~controllable_BtoR_REQ0 & ~n12188;
  assign n12190 = ~controllable_BtoR_REQ0 & ~n12189;
  assign n12191 = i_RtoB_ACK0 & ~n12190;
  assign n12192 = ~n7563 & ~n11156;
  assign n12193 = controllable_BtoR_REQ1 & ~n12192;
  assign n12194 = ~n5243 & ~n12184;
  assign n12195 = ~controllable_BtoR_REQ1 & ~n12194;
  assign n12196 = ~n12193 & ~n12195;
  assign n12197 = ~controllable_BtoR_REQ0 & ~n12196;
  assign n12198 = ~controllable_BtoR_REQ0 & ~n12197;
  assign n12199 = ~i_RtoB_ACK0 & ~n12198;
  assign n12200 = ~n12191 & ~n12199;
  assign n12201 = ~controllable_DEQ & ~n12200;
  assign n12202 = ~n12183 & ~n12201;
  assign n12203 = i_nEMPTY & ~n12202;
  assign n12204 = ~controllable_ENQ & ~n12173;
  assign n12205 = ~i_RtoB_ACK1 & ~n12204;
  assign n12206 = ~i_RtoB_ACK1 & ~n12205;
  assign n12207 = ~controllable_BtoR_REQ1 & ~n12206;
  assign n12208 = ~n11183 & ~n12207;
  assign n12209 = ~controllable_BtoR_REQ0 & ~n12208;
  assign n12210 = ~controllable_BtoR_REQ0 & ~n12209;
  assign n12211 = ~i_RtoB_ACK0 & ~n12210;
  assign n12212 = ~i_RtoB_ACK0 & ~n12211;
  assign n12213 = controllable_DEQ & ~n12212;
  assign n12214 = ~i_RtoB_ACK1 & ~n11144;
  assign n12215 = ~n5237 & ~n12214;
  assign n12216 = controllable_BtoR_REQ1 & ~n12215;
  assign n12217 = ~n8755 & ~n11150;
  assign n12218 = ~controllable_BtoR_REQ1 & ~n12217;
  assign n12219 = ~n12216 & ~n12218;
  assign n12220 = ~controllable_BtoR_REQ0 & ~n12219;
  assign n12221 = ~controllable_BtoR_REQ0 & ~n12220;
  assign n12222 = ~i_RtoB_ACK0 & ~n12221;
  assign n12223 = ~n12170 & ~n12222;
  assign n12224 = ~controllable_DEQ & ~n12223;
  assign n12225 = ~n12213 & ~n12224;
  assign n12226 = i_FULL & ~n12225;
  assign n12227 = ~i_RtoB_ACK1 & ~n12185;
  assign n12228 = ~controllable_BtoR_REQ1 & ~n12227;
  assign n12229 = ~n11167 & ~n12228;
  assign n12230 = ~controllable_BtoR_REQ0 & ~n12229;
  assign n12231 = ~controllable_BtoR_REQ0 & ~n12230;
  assign n12232 = ~i_RtoB_ACK0 & ~n12231;
  assign n12233 = ~i_RtoB_ACK0 & ~n12232;
  assign n12234 = controllable_DEQ & ~n12233;
  assign n12235 = ~n5240 & ~n11150;
  assign n12236 = ~controllable_BtoR_REQ1 & ~n12235;
  assign n12237 = ~n12172 & ~n12236;
  assign n12238 = ~controllable_BtoR_REQ0 & ~n12237;
  assign n12239 = ~controllable_BtoR_REQ0 & ~n12238;
  assign n12240 = ~i_RtoB_ACK0 & ~n12239;
  assign n12241 = ~n12170 & ~n12240;
  assign n12242 = ~controllable_DEQ & ~n12241;
  assign n12243 = ~n12234 & ~n12242;
  assign n12244 = ~i_FULL & ~n12243;
  assign n12245 = ~n12226 & ~n12244;
  assign n12246 = ~i_nEMPTY & ~n12245;
  assign n12247 = ~n12203 & ~n12246;
  assign n12248 = controllable_BtoS_ACK0 & ~n12247;
  assign n12249 = ~i_StoB_REQ14 & ~n10583;
  assign n12250 = ~i_StoB_REQ14 & ~n12249;
  assign n12251 = controllable_BtoS_ACK14 & ~n12250;
  assign n12252 = ~n8048 & ~n12249;
  assign n12253 = ~controllable_BtoS_ACK14 & ~n12252;
  assign n12254 = ~n12251 & ~n12253;
  assign n12255 = controllable_ENQ & ~n12254;
  assign n12256 = controllable_ENQ & ~n12255;
  assign n12257 = ~i_RtoB_ACK1 & ~n12256;
  assign n12258 = ~n5343 & ~n12257;
  assign n12259 = ~controllable_BtoR_REQ1 & ~n12258;
  assign n12260 = ~n5330 & ~n12259;
  assign n12261 = ~controllable_BtoR_REQ0 & ~n12260;
  assign n12262 = ~controllable_BtoR_REQ0 & ~n12261;
  assign n12263 = i_RtoB_ACK0 & ~n12262;
  assign n12264 = ~controllable_ENQ & ~n12254;
  assign n12265 = ~n8852 & ~n12264;
  assign n12266 = ~i_RtoB_ACK1 & ~n12265;
  assign n12267 = ~n5343 & ~n12266;
  assign n12268 = ~controllable_BtoR_REQ1 & ~n12267;
  assign n12269 = ~n8972 & ~n12268;
  assign n12270 = ~controllable_BtoR_REQ0 & ~n12269;
  assign n12271 = ~controllable_BtoR_REQ0 & ~n12270;
  assign n12272 = ~i_RtoB_ACK0 & ~n12271;
  assign n12273 = ~n12263 & ~n12272;
  assign n12274 = controllable_DEQ & ~n12273;
  assign n12275 = ~i_RtoB_ACK1 & ~n12254;
  assign n12276 = ~n8983 & ~n12275;
  assign n12277 = ~controllable_BtoR_REQ1 & ~n12276;
  assign n12278 = ~n5360 & ~n12277;
  assign n12279 = ~controllable_BtoR_REQ0 & ~n12278;
  assign n12280 = ~controllable_BtoR_REQ0 & ~n12279;
  assign n12281 = i_RtoB_ACK0 & ~n12280;
  assign n12282 = ~n8985 & ~n8991;
  assign n12283 = ~controllable_BtoR_REQ0 & ~n12282;
  assign n12284 = ~controllable_BtoR_REQ0 & ~n12283;
  assign n12285 = ~i_RtoB_ACK0 & ~n12284;
  assign n12286 = ~n12281 & ~n12285;
  assign n12287 = ~controllable_DEQ & ~n12286;
  assign n12288 = ~n12274 & ~n12287;
  assign n12289 = i_nEMPTY & ~n12288;
  assign n12290 = ~controllable_ENQ & ~n12264;
  assign n12291 = ~i_RtoB_ACK1 & ~n12290;
  assign n12292 = ~i_RtoB_ACK1 & ~n12291;
  assign n12293 = ~controllable_BtoR_REQ1 & ~n12292;
  assign n12294 = ~n5376 & ~n12293;
  assign n12295 = ~controllable_BtoR_REQ0 & ~n12294;
  assign n12296 = ~controllable_BtoR_REQ0 & ~n12295;
  assign n12297 = ~i_RtoB_ACK0 & ~n12296;
  assign n12298 = ~i_RtoB_ACK0 & ~n12297;
  assign n12299 = controllable_DEQ & ~n12298;
  assign n12300 = ~n8966 & ~n9028;
  assign n12301 = ~controllable_BtoR_REQ0 & ~n12300;
  assign n12302 = ~controllable_BtoR_REQ0 & ~n12301;
  assign n12303 = ~i_RtoB_ACK0 & ~n12302;
  assign n12304 = ~n12263 & ~n12303;
  assign n12305 = ~controllable_DEQ & ~n12304;
  assign n12306 = ~n12299 & ~n12305;
  assign n12307 = i_FULL & ~n12306;
  assign n12308 = ~i_RtoB_ACK1 & ~n12275;
  assign n12309 = ~controllable_BtoR_REQ1 & ~n12308;
  assign n12310 = ~n5360 & ~n12309;
  assign n12311 = ~controllable_BtoR_REQ0 & ~n12310;
  assign n12312 = ~controllable_BtoR_REQ0 & ~n12311;
  assign n12313 = ~i_RtoB_ACK0 & ~n12312;
  assign n12314 = ~i_RtoB_ACK0 & ~n12313;
  assign n12315 = controllable_DEQ & ~n12314;
  assign n12316 = ~n8852 & ~n8946;
  assign n12317 = ~i_RtoB_ACK1 & ~n12316;
  assign n12318 = ~n5343 & ~n12317;
  assign n12319 = ~controllable_BtoR_REQ1 & ~n12318;
  assign n12320 = ~n8972 & ~n12319;
  assign n12321 = ~controllable_BtoR_REQ0 & ~n12320;
  assign n12322 = ~controllable_BtoR_REQ0 & ~n12321;
  assign n12323 = ~i_RtoB_ACK0 & ~n12322;
  assign n12324 = ~n12263 & ~n12323;
  assign n12325 = ~controllable_DEQ & ~n12324;
  assign n12326 = ~n12315 & ~n12325;
  assign n12327 = ~i_FULL & ~n12326;
  assign n12328 = ~n12307 & ~n12327;
  assign n12329 = ~i_nEMPTY & ~n12328;
  assign n12330 = ~n12289 & ~n12329;
  assign n12331 = ~controllable_BtoS_ACK0 & ~n12330;
  assign n12332 = ~n12248 & ~n12331;
  assign n12333 = n4465 & ~n12332;
  assign n12334 = ~n8989 & ~n12285;
  assign n12335 = ~controllable_DEQ & ~n12334;
  assign n12336 = ~n9007 & ~n12335;
  assign n12337 = i_nEMPTY & ~n12336;
  assign n12338 = ~n8970 & ~n12303;
  assign n12339 = ~controllable_DEQ & ~n12338;
  assign n12340 = ~n9025 & ~n12339;
  assign n12341 = i_FULL & ~n12340;
  assign n12342 = ~n8970 & ~n12323;
  assign n12343 = ~controllable_DEQ & ~n12342;
  assign n12344 = ~n9042 & ~n12343;
  assign n12345 = ~i_FULL & ~n12344;
  assign n12346 = ~n12341 & ~n12345;
  assign n12347 = ~i_nEMPTY & ~n12346;
  assign n12348 = ~n12337 & ~n12347;
  assign n12349 = ~controllable_BtoS_ACK0 & ~n12348;
  assign n12350 = ~n5307 & ~n12349;
  assign n12351 = ~n4465 & ~n12350;
  assign n12352 = ~n12333 & ~n12351;
  assign n12353 = i_StoB_REQ10 & ~n12352;
  assign n12354 = ~n11380 & ~n12353;
  assign n12355 = controllable_BtoS_ACK10 & ~n12354;
  assign n12356 = ~n9836 & ~n11410;
  assign n12357 = ~controllable_BtoR_REQ1 & ~n12356;
  assign n12358 = ~n11392 & ~n12357;
  assign n12359 = ~controllable_BtoR_REQ0 & ~n12358;
  assign n12360 = ~controllable_BtoR_REQ0 & ~n12359;
  assign n12361 = i_RtoB_ACK0 & ~n12360;
  assign n12362 = ~n10149 & ~n11407;
  assign n12363 = controllable_BtoR_REQ1 & ~n12362;
  assign n12364 = ~i_StoB_REQ14 & ~n10472;
  assign n12365 = ~n7690 & ~n12364;
  assign n12366 = controllable_BtoS_ACK14 & ~n12365;
  assign n12367 = ~n10473 & ~n12366;
  assign n12368 = controllable_ENQ & ~n12367;
  assign n12369 = ~n9545 & ~n12368;
  assign n12370 = ~i_RtoB_ACK1 & ~n12369;
  assign n12371 = ~n11410 & ~n12370;
  assign n12372 = ~controllable_BtoR_REQ1 & ~n12371;
  assign n12373 = ~n12363 & ~n12372;
  assign n12374 = ~controllable_BtoR_REQ0 & ~n12373;
  assign n12375 = ~controllable_BtoR_REQ0 & ~n12374;
  assign n12376 = ~i_RtoB_ACK0 & ~n12375;
  assign n12377 = ~n12361 & ~n12376;
  assign n12378 = controllable_DEQ & ~n12377;
  assign n12379 = ~n9813 & ~n11428;
  assign n12380 = ~controllable_BtoR_REQ1 & ~n12379;
  assign n12381 = ~n11421 & ~n12380;
  assign n12382 = ~controllable_BtoR_REQ0 & ~n12381;
  assign n12383 = ~controllable_BtoR_REQ0 & ~n12382;
  assign n12384 = i_RtoB_ACK0 & ~n12383;
  assign n12385 = ~n9517 & ~n11429;
  assign n12386 = controllable_BtoR_REQ1 & ~n12385;
  assign n12387 = ~i_RtoB_ACK1 & ~n12367;
  assign n12388 = ~n11428 & ~n12387;
  assign n12389 = ~controllable_BtoR_REQ1 & ~n12388;
  assign n12390 = ~n12386 & ~n12389;
  assign n12391 = ~controllable_BtoR_REQ0 & ~n12390;
  assign n12392 = ~controllable_BtoR_REQ0 & ~n12391;
  assign n12393 = ~i_RtoB_ACK0 & ~n12392;
  assign n12394 = ~n12384 & ~n12393;
  assign n12395 = ~controllable_DEQ & ~n12394;
  assign n12396 = ~n12378 & ~n12395;
  assign n12397 = i_FULL & ~n12396;
  assign n12398 = ~n10149 & ~n11419;
  assign n12399 = controllable_BtoR_REQ1 & ~n12398;
  assign n12400 = ~n9813 & ~n11410;
  assign n12401 = ~controllable_BtoR_REQ1 & ~n12400;
  assign n12402 = ~n12399 & ~n12401;
  assign n12403 = ~controllable_BtoR_REQ0 & ~n12402;
  assign n12404 = ~controllable_BtoR_REQ0 & ~n12403;
  assign n12405 = ~i_RtoB_ACK0 & ~n12404;
  assign n12406 = ~n12361 & ~n12405;
  assign n12407 = controllable_DEQ & ~n12406;
  assign n12408 = ~n9517 & ~n11407;
  assign n12409 = controllable_BtoR_REQ1 & ~n12408;
  assign n12410 = ~n11428 & ~n12370;
  assign n12411 = ~controllable_BtoR_REQ1 & ~n12410;
  assign n12412 = ~n12409 & ~n12411;
  assign n12413 = ~controllable_BtoR_REQ0 & ~n12412;
  assign n12414 = ~controllable_BtoR_REQ0 & ~n12413;
  assign n12415 = ~i_RtoB_ACK0 & ~n12414;
  assign n12416 = ~n12384 & ~n12415;
  assign n12417 = ~controllable_DEQ & ~n12416;
  assign n12418 = ~n12407 & ~n12417;
  assign n12419 = ~i_FULL & ~n12418;
  assign n12420 = ~n12397 & ~n12419;
  assign n12421 = i_nEMPTY & ~n12420;
  assign n12422 = ~n10049 & ~n11468;
  assign n12423 = ~controllable_BtoR_REQ0 & ~n12422;
  assign n12424 = ~controllable_BtoR_REQ0 & ~n12423;
  assign n12425 = ~i_RtoB_ACK0 & ~n12424;
  assign n12426 = ~i_RtoB_ACK0 & ~n12425;
  assign n12427 = controllable_DEQ & ~n12426;
  assign n12428 = ~n9571 & ~n11479;
  assign n12429 = controllable_BtoR_REQ1 & ~n12428;
  assign n12430 = controllable_ENQ & ~n12368;
  assign n12431 = ~i_RtoB_ACK1 & ~n12430;
  assign n12432 = ~n11410 & ~n12431;
  assign n12433 = ~controllable_BtoR_REQ1 & ~n12432;
  assign n12434 = ~n12429 & ~n12433;
  assign n12435 = ~controllable_BtoR_REQ0 & ~n12434;
  assign n12436 = ~controllable_BtoR_REQ0 & ~n12435;
  assign n12437 = ~i_RtoB_ACK0 & ~n12436;
  assign n12438 = ~n12361 & ~n12437;
  assign n12439 = ~controllable_DEQ & ~n12438;
  assign n12440 = ~n12427 & ~n12439;
  assign n12441 = i_FULL & ~n12440;
  assign n12442 = ~n10061 & ~n11421;
  assign n12443 = ~controllable_BtoR_REQ0 & ~n12442;
  assign n12444 = ~controllable_BtoR_REQ0 & ~n12443;
  assign n12445 = ~i_RtoB_ACK0 & ~n12444;
  assign n12446 = ~i_RtoB_ACK0 & ~n12445;
  assign n12447 = controllable_DEQ & ~n12446;
  assign n12448 = ~controllable_DEQ & ~n12377;
  assign n12449 = ~n12447 & ~n12448;
  assign n12450 = ~i_FULL & ~n12449;
  assign n12451 = ~n12441 & ~n12450;
  assign n12452 = ~i_nEMPTY & ~n12451;
  assign n12453 = ~n12421 & ~n12452;
  assign n12454 = controllable_BtoS_ACK0 & ~n12453;
  assign n12455 = ~n9871 & ~n11527;
  assign n12456 = ~controllable_BtoR_REQ1 & ~n12455;
  assign n12457 = ~n11514 & ~n12456;
  assign n12458 = ~controllable_BtoR_REQ0 & ~n12457;
  assign n12459 = ~controllable_BtoR_REQ0 & ~n12458;
  assign n12460 = i_RtoB_ACK0 & ~n12459;
  assign n12461 = ~n8864 & ~n9635;
  assign n12462 = i_RtoB_ACK1 & ~n12461;
  assign n12463 = ~n11524 & ~n12462;
  assign n12464 = controllable_BtoR_REQ1 & ~n12463;
  assign n12465 = ~n9895 & ~n11527;
  assign n12466 = ~controllable_BtoR_REQ1 & ~n12465;
  assign n12467 = ~n12464 & ~n12466;
  assign n12468 = ~controllable_BtoR_REQ0 & ~n12467;
  assign n12469 = ~controllable_BtoR_REQ0 & ~n12468;
  assign n12470 = ~i_RtoB_ACK0 & ~n12469;
  assign n12471 = ~n12460 & ~n12470;
  assign n12472 = controllable_DEQ & ~n12471;
  assign n12473 = ~n9904 & ~n11544;
  assign n12474 = ~controllable_BtoR_REQ1 & ~n12473;
  assign n12475 = ~n11538 & ~n12474;
  assign n12476 = ~controllable_BtoR_REQ0 & ~n12475;
  assign n12477 = ~controllable_BtoR_REQ0 & ~n12476;
  assign n12478 = i_RtoB_ACK0 & ~n12477;
  assign n12479 = ~n9913 & ~n11544;
  assign n12480 = ~controllable_BtoR_REQ1 & ~n12479;
  assign n12481 = ~n9912 & ~n12480;
  assign n12482 = ~controllable_BtoR_REQ0 & ~n12481;
  assign n12483 = ~controllable_BtoR_REQ0 & ~n12482;
  assign n12484 = ~i_RtoB_ACK0 & ~n12483;
  assign n12485 = ~n12478 & ~n12484;
  assign n12486 = ~controllable_DEQ & ~n12485;
  assign n12487 = ~n12472 & ~n12486;
  assign n12488 = i_FULL & ~n12487;
  assign n12489 = ~n11536 & ~n12462;
  assign n12490 = controllable_BtoR_REQ1 & ~n12489;
  assign n12491 = ~n9904 & ~n11527;
  assign n12492 = ~controllable_BtoR_REQ1 & ~n12491;
  assign n12493 = ~n12490 & ~n12492;
  assign n12494 = ~controllable_BtoR_REQ0 & ~n12493;
  assign n12495 = ~controllable_BtoR_REQ0 & ~n12494;
  assign n12496 = ~i_RtoB_ACK0 & ~n12495;
  assign n12497 = ~n12460 & ~n12496;
  assign n12498 = controllable_DEQ & ~n12497;
  assign n12499 = ~n9664 & ~n11524;
  assign n12500 = controllable_BtoR_REQ1 & ~n12499;
  assign n12501 = ~n9895 & ~n11544;
  assign n12502 = ~controllable_BtoR_REQ1 & ~n12501;
  assign n12503 = ~n12500 & ~n12502;
  assign n12504 = ~controllable_BtoR_REQ0 & ~n12503;
  assign n12505 = ~controllable_BtoR_REQ0 & ~n12504;
  assign n12506 = ~i_RtoB_ACK0 & ~n12505;
  assign n12507 = ~n12478 & ~n12506;
  assign n12508 = ~controllable_DEQ & ~n12507;
  assign n12509 = ~n12498 & ~n12508;
  assign n12510 = ~i_FULL & ~n12509;
  assign n12511 = ~n12488 & ~n12510;
  assign n12512 = i_nEMPTY & ~n12511;
  assign n12513 = ~n9951 & ~n11584;
  assign n12514 = ~controllable_BtoR_REQ0 & ~n12513;
  assign n12515 = ~controllable_BtoR_REQ0 & ~n12514;
  assign n12516 = ~i_RtoB_ACK0 & ~n12515;
  assign n12517 = ~i_RtoB_ACK0 & ~n12516;
  assign n12518 = controllable_DEQ & ~n12517;
  assign n12519 = ~n9961 & ~n11527;
  assign n12520 = ~controllable_BtoR_REQ1 & ~n12519;
  assign n12521 = ~n9959 & ~n12520;
  assign n12522 = ~controllable_BtoR_REQ0 & ~n12521;
  assign n12523 = ~controllable_BtoR_REQ0 & ~n12522;
  assign n12524 = ~i_RtoB_ACK0 & ~n12523;
  assign n12525 = ~n12460 & ~n12524;
  assign n12526 = ~controllable_DEQ & ~n12525;
  assign n12527 = ~n12518 & ~n12526;
  assign n12528 = i_FULL & ~n12527;
  assign n12529 = ~n9973 & ~n11538;
  assign n12530 = ~controllable_BtoR_REQ0 & ~n12529;
  assign n12531 = ~controllable_BtoR_REQ0 & ~n12530;
  assign n12532 = ~i_RtoB_ACK0 & ~n12531;
  assign n12533 = ~i_RtoB_ACK0 & ~n12532;
  assign n12534 = controllable_DEQ & ~n12533;
  assign n12535 = ~controllable_DEQ & ~n12471;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = ~i_FULL & ~n12536;
  assign n12538 = ~n12528 & ~n12537;
  assign n12539 = ~i_nEMPTY & ~n12538;
  assign n12540 = ~n12512 & ~n12539;
  assign n12541 = ~controllable_BtoS_ACK0 & ~n12540;
  assign n12542 = ~n12454 & ~n12541;
  assign n12543 = n4465 & ~n12542;
  assign n12544 = ~n10190 & ~n12541;
  assign n12545 = ~n4465 & ~n12544;
  assign n12546 = ~n12543 & ~n12545;
  assign n12547 = i_StoB_REQ10 & ~n12546;
  assign n12548 = ~n9836 & ~n11663;
  assign n12549 = ~controllable_BtoR_REQ1 & ~n12548;
  assign n12550 = ~n11643 & ~n12549;
  assign n12551 = ~controllable_BtoR_REQ0 & ~n12550;
  assign n12552 = ~controllable_BtoR_REQ0 & ~n12551;
  assign n12553 = i_RtoB_ACK0 & ~n12552;
  assign n12554 = ~n9302 & ~n11655;
  assign n12555 = i_RtoB_ACK1 & ~n12554;
  assign n12556 = ~n11660 & ~n12555;
  assign n12557 = controllable_BtoR_REQ1 & ~n12556;
  assign n12558 = ~n11663 & ~n12370;
  assign n12559 = ~controllable_BtoR_REQ1 & ~n12558;
  assign n12560 = ~n12557 & ~n12559;
  assign n12561 = ~controllable_BtoR_REQ0 & ~n12560;
  assign n12562 = ~controllable_BtoR_REQ0 & ~n12561;
  assign n12563 = ~i_RtoB_ACK0 & ~n12562;
  assign n12564 = ~n12553 & ~n12563;
  assign n12565 = controllable_DEQ & ~n12564;
  assign n12566 = ~n9813 & ~n11684;
  assign n12567 = ~controllable_BtoR_REQ1 & ~n12566;
  assign n12568 = ~n11678 & ~n12567;
  assign n12569 = ~controllable_BtoR_REQ0 & ~n12568;
  assign n12570 = ~controllable_BtoR_REQ0 & ~n12569;
  assign n12571 = i_RtoB_ACK0 & ~n12570;
  assign n12572 = ~n11684 & ~n12387;
  assign n12573 = ~controllable_BtoR_REQ1 & ~n12572;
  assign n12574 = ~n12386 & ~n12573;
  assign n12575 = ~controllable_BtoR_REQ0 & ~n12574;
  assign n12576 = ~controllable_BtoR_REQ0 & ~n12575;
  assign n12577 = ~i_RtoB_ACK0 & ~n12576;
  assign n12578 = ~n12571 & ~n12577;
  assign n12579 = ~controllable_DEQ & ~n12578;
  assign n12580 = ~n12565 & ~n12579;
  assign n12581 = i_FULL & ~n12580;
  assign n12582 = ~n11698 & ~n12555;
  assign n12583 = controllable_BtoR_REQ1 & ~n12582;
  assign n12584 = ~n9813 & ~n11663;
  assign n12585 = ~controllable_BtoR_REQ1 & ~n12584;
  assign n12586 = ~n12583 & ~n12585;
  assign n12587 = ~controllable_BtoR_REQ0 & ~n12586;
  assign n12588 = ~controllable_BtoR_REQ0 & ~n12587;
  assign n12589 = ~i_RtoB_ACK0 & ~n12588;
  assign n12590 = ~n12553 & ~n12589;
  assign n12591 = controllable_DEQ & ~n12590;
  assign n12592 = ~n9517 & ~n11666;
  assign n12593 = controllable_BtoR_REQ1 & ~n12592;
  assign n12594 = ~n11684 & ~n12370;
  assign n12595 = ~controllable_BtoR_REQ1 & ~n12594;
  assign n12596 = ~n12593 & ~n12595;
  assign n12597 = ~controllable_BtoR_REQ0 & ~n12596;
  assign n12598 = ~controllable_BtoR_REQ0 & ~n12597;
  assign n12599 = ~i_RtoB_ACK0 & ~n12598;
  assign n12600 = ~n12571 & ~n12599;
  assign n12601 = ~controllable_DEQ & ~n12600;
  assign n12602 = ~n12591 & ~n12601;
  assign n12603 = ~i_FULL & ~n12602;
  assign n12604 = ~n12581 & ~n12603;
  assign n12605 = i_nEMPTY & ~n12604;
  assign n12606 = ~n10049 & ~n11728;
  assign n12607 = ~controllable_BtoR_REQ0 & ~n12606;
  assign n12608 = ~controllable_BtoR_REQ0 & ~n12607;
  assign n12609 = ~i_RtoB_ACK0 & ~n12608;
  assign n12610 = ~i_RtoB_ACK0 & ~n12609;
  assign n12611 = controllable_DEQ & ~n12610;
  assign n12612 = ~n11663 & ~n12431;
  assign n12613 = ~controllable_BtoR_REQ1 & ~n12612;
  assign n12614 = ~n12429 & ~n12613;
  assign n12615 = ~controllable_BtoR_REQ0 & ~n12614;
  assign n12616 = ~controllable_BtoR_REQ0 & ~n12615;
  assign n12617 = ~i_RtoB_ACK0 & ~n12616;
  assign n12618 = ~n12553 & ~n12617;
  assign n12619 = ~controllable_DEQ & ~n12618;
  assign n12620 = ~n12611 & ~n12619;
  assign n12621 = i_FULL & ~n12620;
  assign n12622 = ~n10061 & ~n11678;
  assign n12623 = ~controllable_BtoR_REQ0 & ~n12622;
  assign n12624 = ~controllable_BtoR_REQ0 & ~n12623;
  assign n12625 = ~i_RtoB_ACK0 & ~n12624;
  assign n12626 = ~i_RtoB_ACK0 & ~n12625;
  assign n12627 = controllable_DEQ & ~n12626;
  assign n12628 = ~n9597 & ~n12368;
  assign n12629 = ~i_RtoB_ACK1 & ~n12628;
  assign n12630 = ~n11663 & ~n12629;
  assign n12631 = ~controllable_BtoR_REQ1 & ~n12630;
  assign n12632 = ~n12557 & ~n12631;
  assign n12633 = ~controllable_BtoR_REQ0 & ~n12632;
  assign n12634 = ~controllable_BtoR_REQ0 & ~n12633;
  assign n12635 = ~i_RtoB_ACK0 & ~n12634;
  assign n12636 = ~n12553 & ~n12635;
  assign n12637 = ~controllable_DEQ & ~n12636;
  assign n12638 = ~n12627 & ~n12637;
  assign n12639 = ~i_FULL & ~n12638;
  assign n12640 = ~n12621 & ~n12639;
  assign n12641 = ~i_nEMPTY & ~n12640;
  assign n12642 = ~n12605 & ~n12641;
  assign n12643 = controllable_BtoS_ACK0 & ~n12642;
  assign n12644 = ~n9871 & ~n11810;
  assign n12645 = ~controllable_BtoR_REQ1 & ~n12644;
  assign n12646 = ~n11790 & ~n12645;
  assign n12647 = ~controllable_BtoR_REQ0 & ~n12646;
  assign n12648 = ~controllable_BtoR_REQ0 & ~n12647;
  assign n12649 = i_RtoB_ACK0 & ~n12648;
  assign n12650 = ~n9635 & ~n11802;
  assign n12651 = i_RtoB_ACK1 & ~n12650;
  assign n12652 = ~n11807 & ~n12651;
  assign n12653 = controllable_BtoR_REQ1 & ~n12652;
  assign n12654 = ~n9895 & ~n11810;
  assign n12655 = ~controllable_BtoR_REQ1 & ~n12654;
  assign n12656 = ~n12653 & ~n12655;
  assign n12657 = ~controllable_BtoR_REQ0 & ~n12656;
  assign n12658 = ~controllable_BtoR_REQ0 & ~n12657;
  assign n12659 = ~i_RtoB_ACK0 & ~n12658;
  assign n12660 = ~n12649 & ~n12659;
  assign n12661 = controllable_DEQ & ~n12660;
  assign n12662 = ~n9904 & ~n11831;
  assign n12663 = ~controllable_BtoR_REQ1 & ~n12662;
  assign n12664 = ~n11825 & ~n12663;
  assign n12665 = ~controllable_BtoR_REQ0 & ~n12664;
  assign n12666 = ~controllable_BtoR_REQ0 & ~n12665;
  assign n12667 = i_RtoB_ACK0 & ~n12666;
  assign n12668 = ~n9913 & ~n11831;
  assign n12669 = ~controllable_BtoR_REQ1 & ~n12668;
  assign n12670 = ~n9912 & ~n12669;
  assign n12671 = ~controllable_BtoR_REQ0 & ~n12670;
  assign n12672 = ~controllable_BtoR_REQ0 & ~n12671;
  assign n12673 = ~i_RtoB_ACK0 & ~n12672;
  assign n12674 = ~n12667 & ~n12673;
  assign n12675 = ~controllable_DEQ & ~n12674;
  assign n12676 = ~n12661 & ~n12675;
  assign n12677 = i_FULL & ~n12676;
  assign n12678 = ~n11845 & ~n12651;
  assign n12679 = controllable_BtoR_REQ1 & ~n12678;
  assign n12680 = ~n9904 & ~n11810;
  assign n12681 = ~controllable_BtoR_REQ1 & ~n12680;
  assign n12682 = ~n12679 & ~n12681;
  assign n12683 = ~controllable_BtoR_REQ0 & ~n12682;
  assign n12684 = ~controllable_BtoR_REQ0 & ~n12683;
  assign n12685 = ~i_RtoB_ACK0 & ~n12684;
  assign n12686 = ~n12649 & ~n12685;
  assign n12687 = controllable_DEQ & ~n12686;
  assign n12688 = ~n9664 & ~n11813;
  assign n12689 = controllable_BtoR_REQ1 & ~n12688;
  assign n12690 = ~n9895 & ~n11831;
  assign n12691 = ~controllable_BtoR_REQ1 & ~n12690;
  assign n12692 = ~n12689 & ~n12691;
  assign n12693 = ~controllable_BtoR_REQ0 & ~n12692;
  assign n12694 = ~controllable_BtoR_REQ0 & ~n12693;
  assign n12695 = ~i_RtoB_ACK0 & ~n12694;
  assign n12696 = ~n12667 & ~n12695;
  assign n12697 = ~controllable_DEQ & ~n12696;
  assign n12698 = ~n12687 & ~n12697;
  assign n12699 = ~i_FULL & ~n12698;
  assign n12700 = ~n12677 & ~n12699;
  assign n12701 = i_nEMPTY & ~n12700;
  assign n12702 = ~n9951 & ~n11875;
  assign n12703 = ~controllable_BtoR_REQ0 & ~n12702;
  assign n12704 = ~controllable_BtoR_REQ0 & ~n12703;
  assign n12705 = ~i_RtoB_ACK0 & ~n12704;
  assign n12706 = ~i_RtoB_ACK0 & ~n12705;
  assign n12707 = controllable_DEQ & ~n12706;
  assign n12708 = ~n9961 & ~n11810;
  assign n12709 = ~controllable_BtoR_REQ1 & ~n12708;
  assign n12710 = ~n9959 & ~n12709;
  assign n12711 = ~controllable_BtoR_REQ0 & ~n12710;
  assign n12712 = ~controllable_BtoR_REQ0 & ~n12711;
  assign n12713 = ~i_RtoB_ACK0 & ~n12712;
  assign n12714 = ~n12649 & ~n12713;
  assign n12715 = ~controllable_DEQ & ~n12714;
  assign n12716 = ~n12707 & ~n12715;
  assign n12717 = i_FULL & ~n12716;
  assign n12718 = ~n9973 & ~n11825;
  assign n12719 = ~controllable_BtoR_REQ0 & ~n12718;
  assign n12720 = ~controllable_BtoR_REQ0 & ~n12719;
  assign n12721 = ~i_RtoB_ACK0 & ~n12720;
  assign n12722 = ~i_RtoB_ACK0 & ~n12721;
  assign n12723 = controllable_DEQ & ~n12722;
  assign n12724 = ~n9981 & ~n11810;
  assign n12725 = ~controllable_BtoR_REQ1 & ~n12724;
  assign n12726 = ~n12653 & ~n12725;
  assign n12727 = ~controllable_BtoR_REQ0 & ~n12726;
  assign n12728 = ~controllable_BtoR_REQ0 & ~n12727;
  assign n12729 = ~i_RtoB_ACK0 & ~n12728;
  assign n12730 = ~n12649 & ~n12729;
  assign n12731 = ~controllable_DEQ & ~n12730;
  assign n12732 = ~n12723 & ~n12731;
  assign n12733 = ~i_FULL & ~n12732;
  assign n12734 = ~n12717 & ~n12733;
  assign n12735 = ~i_nEMPTY & ~n12734;
  assign n12736 = ~n12701 & ~n12735;
  assign n12737 = ~controllable_BtoS_ACK0 & ~n12736;
  assign n12738 = ~n12643 & ~n12737;
  assign n12739 = n4465 & ~n12738;
  assign n12740 = ~n7081 & ~n9838;
  assign n12741 = ~controllable_BtoR_REQ0 & ~n12740;
  assign n12742 = ~controllable_BtoR_REQ0 & ~n12741;
  assign n12743 = i_RtoB_ACK0 & ~n12742;
  assign n12744 = ~n9791 & ~n10153;
  assign n12745 = ~controllable_BtoR_REQ0 & ~n12744;
  assign n12746 = ~controllable_BtoR_REQ0 & ~n12745;
  assign n12747 = ~i_RtoB_ACK0 & ~n12746;
  assign n12748 = ~n12743 & ~n12747;
  assign n12749 = controllable_DEQ & ~n12748;
  assign n12750 = ~n7114 & ~n9815;
  assign n12751 = ~controllable_BtoR_REQ0 & ~n12750;
  assign n12752 = ~controllable_BtoR_REQ0 & ~n12751;
  assign n12753 = i_RtoB_ACK0 & ~n12752;
  assign n12754 = ~n9819 & ~n12753;
  assign n12755 = ~controllable_DEQ & ~n12754;
  assign n12756 = ~n12749 & ~n12755;
  assign n12757 = i_nEMPTY & ~n12756;
  assign n12758 = ~n7131 & ~n10049;
  assign n12759 = ~controllable_BtoR_REQ0 & ~n12758;
  assign n12760 = ~controllable_BtoR_REQ0 & ~n12759;
  assign n12761 = ~i_RtoB_ACK0 & ~n12760;
  assign n12762 = ~i_RtoB_ACK0 & ~n12761;
  assign n12763 = controllable_DEQ & ~n12762;
  assign n12764 = ~n9842 & ~n12743;
  assign n12765 = ~controllable_DEQ & ~n12764;
  assign n12766 = ~n12763 & ~n12765;
  assign n12767 = i_FULL & ~n12766;
  assign n12768 = ~n7114 & ~n10061;
  assign n12769 = ~controllable_BtoR_REQ0 & ~n12768;
  assign n12770 = ~controllable_BtoR_REQ0 & ~n12769;
  assign n12771 = ~i_RtoB_ACK0 & ~n12770;
  assign n12772 = ~i_RtoB_ACK0 & ~n12771;
  assign n12773 = controllable_DEQ & ~n12772;
  assign n12774 = ~n9862 & ~n12743;
  assign n12775 = ~controllable_DEQ & ~n12774;
  assign n12776 = ~n12773 & ~n12775;
  assign n12777 = ~i_FULL & ~n12776;
  assign n12778 = ~n12767 & ~n12777;
  assign n12779 = ~i_nEMPTY & ~n12778;
  assign n12780 = ~n12757 & ~n12779;
  assign n12781 = controllable_BtoS_ACK0 & ~n12780;
  assign n12782 = ~n9995 & ~n12781;
  assign n12783 = ~n4465 & ~n12782;
  assign n12784 = ~n12739 & ~n12783;
  assign n12785 = ~i_StoB_REQ10 & ~n12784;
  assign n12786 = ~n12547 & ~n12785;
  assign n12787 = ~controllable_BtoS_ACK10 & ~n12786;
  assign n12788 = ~n12355 & ~n12787;
  assign n12789 = n4464 & ~n12788;
  assign n12790 = ~n10278 & ~n10284;
  assign n12791 = ~controllable_BtoR_REQ0 & ~n12790;
  assign n12792 = ~controllable_BtoR_REQ0 & ~n12791;
  assign n12793 = ~i_RtoB_ACK0 & ~n12792;
  assign n12794 = ~n10282 & ~n12793;
  assign n12795 = ~controllable_DEQ & ~n12794;
  assign n12796 = ~n10300 & ~n12795;
  assign n12797 = i_nEMPTY & ~n12796;
  assign n12798 = ~n10259 & ~n10321;
  assign n12799 = ~controllable_BtoR_REQ0 & ~n12798;
  assign n12800 = ~controllable_BtoR_REQ0 & ~n12799;
  assign n12801 = ~i_RtoB_ACK0 & ~n12800;
  assign n12802 = ~n10263 & ~n12801;
  assign n12803 = ~controllable_DEQ & ~n12802;
  assign n12804 = ~n10318 & ~n12803;
  assign n12805 = i_FULL & ~n12804;
  assign n12806 = ~n5240 & ~n7710;
  assign n12807 = ~controllable_BtoR_REQ1 & ~n12806;
  assign n12808 = ~n10265 & ~n12807;
  assign n12809 = ~controllable_BtoR_REQ0 & ~n12808;
  assign n12810 = ~controllable_BtoR_REQ0 & ~n12809;
  assign n12811 = ~i_RtoB_ACK0 & ~n12810;
  assign n12812 = ~n10263 & ~n12811;
  assign n12813 = ~controllable_DEQ & ~n12812;
  assign n12814 = ~n10335 & ~n12813;
  assign n12815 = ~i_FULL & ~n12814;
  assign n12816 = ~n12805 & ~n12815;
  assign n12817 = ~i_nEMPTY & ~n12816;
  assign n12818 = ~n12797 & ~n12817;
  assign n12819 = controllable_BtoS_ACK0 & ~n12818;
  assign n12820 = ~n10372 & ~n10378;
  assign n12821 = ~controllable_BtoR_REQ0 & ~n12820;
  assign n12822 = ~controllable_BtoR_REQ0 & ~n12821;
  assign n12823 = ~i_RtoB_ACK0 & ~n12822;
  assign n12824 = ~n10376 & ~n12823;
  assign n12825 = ~controllable_DEQ & ~n12824;
  assign n12826 = ~n10394 & ~n12825;
  assign n12827 = i_nEMPTY & ~n12826;
  assign n12828 = ~n10353 & ~n10415;
  assign n12829 = ~controllable_BtoR_REQ0 & ~n12828;
  assign n12830 = ~controllable_BtoR_REQ0 & ~n12829;
  assign n12831 = ~i_RtoB_ACK0 & ~n12830;
  assign n12832 = ~n10357 & ~n12831;
  assign n12833 = ~controllable_DEQ & ~n12832;
  assign n12834 = ~n10412 & ~n12833;
  assign n12835 = i_FULL & ~n12834;
  assign n12836 = ~n7802 & ~n12317;
  assign n12837 = ~controllable_BtoR_REQ1 & ~n12836;
  assign n12838 = ~n10359 & ~n12837;
  assign n12839 = ~controllable_BtoR_REQ0 & ~n12838;
  assign n12840 = ~controllable_BtoR_REQ0 & ~n12839;
  assign n12841 = ~i_RtoB_ACK0 & ~n12840;
  assign n12842 = ~n10357 & ~n12841;
  assign n12843 = ~controllable_DEQ & ~n12842;
  assign n12844 = ~n10429 & ~n12843;
  assign n12845 = ~i_FULL & ~n12844;
  assign n12846 = ~n12835 & ~n12845;
  assign n12847 = ~i_nEMPTY & ~n12846;
  assign n12848 = ~n12827 & ~n12847;
  assign n12849 = ~controllable_BtoS_ACK0 & ~n12848;
  assign n12850 = ~n12819 & ~n12849;
  assign n12851 = n4465 & ~n12850;
  assign n12852 = ~n5307 & ~n12849;
  assign n12853 = ~n4465 & ~n12852;
  assign n12854 = ~n12851 & ~n12853;
  assign n12855 = i_StoB_REQ10 & ~n12854;
  assign n12856 = ~n11380 & ~n12855;
  assign n12857 = controllable_BtoS_ACK10 & ~n12856;
  assign n12858 = ~n9836 & ~n11946;
  assign n12859 = ~controllable_BtoR_REQ1 & ~n12858;
  assign n12860 = ~n11933 & ~n12859;
  assign n12861 = ~controllable_BtoR_REQ0 & ~n12860;
  assign n12862 = ~controllable_BtoR_REQ0 & ~n12861;
  assign n12863 = i_RtoB_ACK0 & ~n12862;
  assign n12864 = ~n10149 & ~n11943;
  assign n12865 = controllable_BtoR_REQ1 & ~n12864;
  assign n12866 = ~n10522 & ~n11946;
  assign n12867 = ~controllable_BtoR_REQ1 & ~n12866;
  assign n12868 = ~n12865 & ~n12867;
  assign n12869 = ~controllable_BtoR_REQ0 & ~n12868;
  assign n12870 = ~controllable_BtoR_REQ0 & ~n12869;
  assign n12871 = ~i_RtoB_ACK0 & ~n12870;
  assign n12872 = ~n12863 & ~n12871;
  assign n12873 = controllable_DEQ & ~n12872;
  assign n12874 = ~n9813 & ~n11963;
  assign n12875 = ~controllable_BtoR_REQ1 & ~n12874;
  assign n12876 = ~n11957 & ~n12875;
  assign n12877 = ~controllable_BtoR_REQ0 & ~n12876;
  assign n12878 = ~controllable_BtoR_REQ0 & ~n12877;
  assign n12879 = i_RtoB_ACK0 & ~n12878;
  assign n12880 = ~n10496 & ~n11963;
  assign n12881 = ~controllable_BtoR_REQ1 & ~n12880;
  assign n12882 = ~n10495 & ~n12881;
  assign n12883 = ~controllable_BtoR_REQ0 & ~n12882;
  assign n12884 = ~controllable_BtoR_REQ0 & ~n12883;
  assign n12885 = ~i_RtoB_ACK0 & ~n12884;
  assign n12886 = ~n12879 & ~n12885;
  assign n12887 = ~controllable_DEQ & ~n12886;
  assign n12888 = ~n12873 & ~n12887;
  assign n12889 = i_FULL & ~n12888;
  assign n12890 = ~n10149 & ~n11955;
  assign n12891 = controllable_BtoR_REQ1 & ~n12890;
  assign n12892 = ~n9813 & ~n11946;
  assign n12893 = ~controllable_BtoR_REQ1 & ~n12892;
  assign n12894 = ~n12891 & ~n12893;
  assign n12895 = ~controllable_BtoR_REQ0 & ~n12894;
  assign n12896 = ~controllable_BtoR_REQ0 & ~n12895;
  assign n12897 = ~i_RtoB_ACK0 & ~n12896;
  assign n12898 = ~n12863 & ~n12897;
  assign n12899 = controllable_DEQ & ~n12898;
  assign n12900 = ~n9517 & ~n11943;
  assign n12901 = controllable_BtoR_REQ1 & ~n12900;
  assign n12902 = ~n10522 & ~n11963;
  assign n12903 = ~controllable_BtoR_REQ1 & ~n12902;
  assign n12904 = ~n12901 & ~n12903;
  assign n12905 = ~controllable_BtoR_REQ0 & ~n12904;
  assign n12906 = ~controllable_BtoR_REQ0 & ~n12905;
  assign n12907 = ~i_RtoB_ACK0 & ~n12906;
  assign n12908 = ~n12879 & ~n12907;
  assign n12909 = ~controllable_DEQ & ~n12908;
  assign n12910 = ~n12899 & ~n12909;
  assign n12911 = ~i_FULL & ~n12910;
  assign n12912 = ~n12889 & ~n12911;
  assign n12913 = i_nEMPTY & ~n12912;
  assign n12914 = ~n10049 & ~n12002;
  assign n12915 = ~controllable_BtoR_REQ0 & ~n12914;
  assign n12916 = ~controllable_BtoR_REQ0 & ~n12915;
  assign n12917 = ~i_RtoB_ACK0 & ~n12916;
  assign n12918 = ~i_RtoB_ACK0 & ~n12917;
  assign n12919 = controllable_DEQ & ~n12918;
  assign n12920 = ~n10548 & ~n11946;
  assign n12921 = ~controllable_BtoR_REQ1 & ~n12920;
  assign n12922 = ~n10546 & ~n12921;
  assign n12923 = ~controllable_BtoR_REQ0 & ~n12922;
  assign n12924 = ~controllable_BtoR_REQ0 & ~n12923;
  assign n12925 = ~i_RtoB_ACK0 & ~n12924;
  assign n12926 = ~n12863 & ~n12925;
  assign n12927 = ~controllable_DEQ & ~n12926;
  assign n12928 = ~n12919 & ~n12927;
  assign n12929 = i_FULL & ~n12928;
  assign n12930 = ~n10061 & ~n11957;
  assign n12931 = ~controllable_BtoR_REQ0 & ~n12930;
  assign n12932 = ~controllable_BtoR_REQ0 & ~n12931;
  assign n12933 = ~i_RtoB_ACK0 & ~n12932;
  assign n12934 = ~i_RtoB_ACK0 & ~n12933;
  assign n12935 = controllable_DEQ & ~n12934;
  assign n12936 = ~controllable_DEQ & ~n12872;
  assign n12937 = ~n12935 & ~n12936;
  assign n12938 = ~i_FULL & ~n12937;
  assign n12939 = ~n12929 & ~n12938;
  assign n12940 = ~i_nEMPTY & ~n12939;
  assign n12941 = ~n12913 & ~n12940;
  assign n12942 = controllable_BtoS_ACK0 & ~n12941;
  assign n12943 = ~n9871 & ~n12054;
  assign n12944 = ~controllable_BtoR_REQ1 & ~n12943;
  assign n12945 = ~n12041 & ~n12944;
  assign n12946 = ~controllable_BtoR_REQ0 & ~n12945;
  assign n12947 = ~controllable_BtoR_REQ0 & ~n12946;
  assign n12948 = i_RtoB_ACK0 & ~n12947;
  assign n12949 = ~n12051 & ~n12462;
  assign n12950 = controllable_BtoR_REQ1 & ~n12949;
  assign n12951 = ~n10649 & ~n12054;
  assign n12952 = ~controllable_BtoR_REQ1 & ~n12951;
  assign n12953 = ~n12950 & ~n12952;
  assign n12954 = ~controllable_BtoR_REQ0 & ~n12953;
  assign n12955 = ~controllable_BtoR_REQ0 & ~n12954;
  assign n12956 = ~i_RtoB_ACK0 & ~n12955;
  assign n12957 = ~n12948 & ~n12956;
  assign n12958 = controllable_DEQ & ~n12957;
  assign n12959 = ~n9904 & ~n12071;
  assign n12960 = ~controllable_BtoR_REQ1 & ~n12959;
  assign n12961 = ~n12065 & ~n12960;
  assign n12962 = ~controllable_BtoR_REQ0 & ~n12961;
  assign n12963 = ~controllable_BtoR_REQ0 & ~n12962;
  assign n12964 = i_RtoB_ACK0 & ~n12963;
  assign n12965 = ~n10623 & ~n12071;
  assign n12966 = ~controllable_BtoR_REQ1 & ~n12965;
  assign n12967 = ~n10622 & ~n12966;
  assign n12968 = ~controllable_BtoR_REQ0 & ~n12967;
  assign n12969 = ~controllable_BtoR_REQ0 & ~n12968;
  assign n12970 = ~i_RtoB_ACK0 & ~n12969;
  assign n12971 = ~n12964 & ~n12970;
  assign n12972 = ~controllable_DEQ & ~n12971;
  assign n12973 = ~n12958 & ~n12972;
  assign n12974 = i_FULL & ~n12973;
  assign n12975 = ~n12063 & ~n12462;
  assign n12976 = controllable_BtoR_REQ1 & ~n12975;
  assign n12977 = ~n9904 & ~n12054;
  assign n12978 = ~controllable_BtoR_REQ1 & ~n12977;
  assign n12979 = ~n12976 & ~n12978;
  assign n12980 = ~controllable_BtoR_REQ0 & ~n12979;
  assign n12981 = ~controllable_BtoR_REQ0 & ~n12980;
  assign n12982 = ~i_RtoB_ACK0 & ~n12981;
  assign n12983 = ~n12948 & ~n12982;
  assign n12984 = controllable_DEQ & ~n12983;
  assign n12985 = ~n9664 & ~n12051;
  assign n12986 = controllable_BtoR_REQ1 & ~n12985;
  assign n12987 = ~n10649 & ~n12071;
  assign n12988 = ~controllable_BtoR_REQ1 & ~n12987;
  assign n12989 = ~n12986 & ~n12988;
  assign n12990 = ~controllable_BtoR_REQ0 & ~n12989;
  assign n12991 = ~controllable_BtoR_REQ0 & ~n12990;
  assign n12992 = ~i_RtoB_ACK0 & ~n12991;
  assign n12993 = ~n12964 & ~n12992;
  assign n12994 = ~controllable_DEQ & ~n12993;
  assign n12995 = ~n12984 & ~n12994;
  assign n12996 = ~i_FULL & ~n12995;
  assign n12997 = ~n12974 & ~n12996;
  assign n12998 = i_nEMPTY & ~n12997;
  assign n12999 = ~n9951 & ~n12110;
  assign n13000 = ~controllable_BtoR_REQ0 & ~n12999;
  assign n13001 = ~controllable_BtoR_REQ0 & ~n13000;
  assign n13002 = ~i_RtoB_ACK0 & ~n13001;
  assign n13003 = ~i_RtoB_ACK0 & ~n13002;
  assign n13004 = controllable_DEQ & ~n13003;
  assign n13005 = ~n10675 & ~n12054;
  assign n13006 = ~controllable_BtoR_REQ1 & ~n13005;
  assign n13007 = ~n10673 & ~n13006;
  assign n13008 = ~controllable_BtoR_REQ0 & ~n13007;
  assign n13009 = ~controllable_BtoR_REQ0 & ~n13008;
  assign n13010 = ~i_RtoB_ACK0 & ~n13009;
  assign n13011 = ~n12948 & ~n13010;
  assign n13012 = ~controllable_DEQ & ~n13011;
  assign n13013 = ~n13004 & ~n13012;
  assign n13014 = i_FULL & ~n13013;
  assign n13015 = ~n9973 & ~n12065;
  assign n13016 = ~controllable_BtoR_REQ0 & ~n13015;
  assign n13017 = ~controllable_BtoR_REQ0 & ~n13016;
  assign n13018 = ~i_RtoB_ACK0 & ~n13017;
  assign n13019 = ~i_RtoB_ACK0 & ~n13018;
  assign n13020 = controllable_DEQ & ~n13019;
  assign n13021 = ~controllable_DEQ & ~n12957;
  assign n13022 = ~n13020 & ~n13021;
  assign n13023 = ~i_FULL & ~n13022;
  assign n13024 = ~n13014 & ~n13023;
  assign n13025 = ~i_nEMPTY & ~n13024;
  assign n13026 = ~n12998 & ~n13025;
  assign n13027 = ~controllable_BtoS_ACK0 & ~n13026;
  assign n13028 = ~n12942 & ~n13027;
  assign n13029 = n4465 & ~n13028;
  assign n13030 = ~n11059 & ~n13027;
  assign n13031 = ~n4465 & ~n13030;
  assign n13032 = ~n13029 & ~n13031;
  assign n13033 = i_StoB_REQ10 & ~n13032;
  assign n13034 = ~n7905 & ~n10882;
  assign n13035 = ~controllable_BtoR_REQ0 & ~n13034;
  assign n13036 = ~controllable_BtoR_REQ0 & ~n13035;
  assign n13037 = i_RtoB_ACK0 & ~n13036;
  assign n13038 = ~n10470 & ~n10892;
  assign n13039 = ~controllable_BtoR_REQ0 & ~n13038;
  assign n13040 = ~controllable_BtoR_REQ0 & ~n13039;
  assign n13041 = ~i_RtoB_ACK0 & ~n13040;
  assign n13042 = ~n13037 & ~n13041;
  assign n13043 = controllable_DEQ & ~n13042;
  assign n13044 = ~n7950 & ~n10900;
  assign n13045 = ~controllable_BtoR_REQ0 & ~n13044;
  assign n13046 = ~controllable_BtoR_REQ0 & ~n13045;
  assign n13047 = i_RtoB_ACK0 & ~n13046;
  assign n13048 = ~n10502 & ~n13047;
  assign n13049 = ~controllable_DEQ & ~n13048;
  assign n13050 = ~n13043 & ~n13049;
  assign n13051 = i_FULL & ~n13050;
  assign n13052 = ~n10508 & ~n10912;
  assign n13053 = ~controllable_BtoR_REQ0 & ~n13052;
  assign n13054 = ~controllable_BtoR_REQ0 & ~n13053;
  assign n13055 = ~i_RtoB_ACK0 & ~n13054;
  assign n13056 = ~n13037 & ~n13055;
  assign n13057 = controllable_DEQ & ~n13056;
  assign n13058 = ~n10528 & ~n13047;
  assign n13059 = ~controllable_DEQ & ~n13058;
  assign n13060 = ~n13057 & ~n13059;
  assign n13061 = ~i_FULL & ~n13060;
  assign n13062 = ~n13051 & ~n13061;
  assign n13063 = i_nEMPTY & ~n13062;
  assign n13064 = ~n8002 & ~n10049;
  assign n13065 = ~controllable_BtoR_REQ0 & ~n13064;
  assign n13066 = ~controllable_BtoR_REQ0 & ~n13065;
  assign n13067 = ~i_RtoB_ACK0 & ~n13066;
  assign n13068 = ~i_RtoB_ACK0 & ~n13067;
  assign n13069 = controllable_DEQ & ~n13068;
  assign n13070 = ~n10554 & ~n13037;
  assign n13071 = ~controllable_DEQ & ~n13070;
  assign n13072 = ~n13069 & ~n13071;
  assign n13073 = i_FULL & ~n13072;
  assign n13074 = ~n7950 & ~n10061;
  assign n13075 = ~controllable_BtoR_REQ0 & ~n13074;
  assign n13076 = ~controllable_BtoR_REQ0 & ~n13075;
  assign n13077 = ~i_RtoB_ACK0 & ~n13076;
  assign n13078 = ~i_RtoB_ACK0 & ~n13077;
  assign n13079 = controllable_DEQ & ~n13078;
  assign n13080 = ~n10574 & ~n13037;
  assign n13081 = ~controllable_DEQ & ~n13080;
  assign n13082 = ~n13079 & ~n13081;
  assign n13083 = ~i_FULL & ~n13082;
  assign n13084 = ~n13073 & ~n13083;
  assign n13085 = ~i_nEMPTY & ~n13084;
  assign n13086 = ~n13063 & ~n13085;
  assign n13087 = controllable_BtoS_ACK0 & ~n13086;
  assign n13088 = ~n8074 & ~n10949;
  assign n13089 = ~controllable_BtoR_REQ0 & ~n13088;
  assign n13090 = ~controllable_BtoR_REQ0 & ~n13089;
  assign n13091 = i_RtoB_ACK0 & ~n13090;
  assign n13092 = ~n10600 & ~n10959;
  assign n13093 = ~controllable_BtoR_REQ0 & ~n13092;
  assign n13094 = ~controllable_BtoR_REQ0 & ~n13093;
  assign n13095 = ~i_RtoB_ACK0 & ~n13094;
  assign n13096 = ~n13091 & ~n13095;
  assign n13097 = controllable_DEQ & ~n13096;
  assign n13098 = ~n8114 & ~n10967;
  assign n13099 = ~controllable_BtoR_REQ0 & ~n13098;
  assign n13100 = ~controllable_BtoR_REQ0 & ~n13099;
  assign n13101 = i_RtoB_ACK0 & ~n13100;
  assign n13102 = ~n10629 & ~n13101;
  assign n13103 = ~controllable_DEQ & ~n13102;
  assign n13104 = ~n13097 & ~n13103;
  assign n13105 = i_FULL & ~n13104;
  assign n13106 = ~n10635 & ~n10979;
  assign n13107 = ~controllable_BtoR_REQ0 & ~n13106;
  assign n13108 = ~controllable_BtoR_REQ0 & ~n13107;
  assign n13109 = ~i_RtoB_ACK0 & ~n13108;
  assign n13110 = ~n13091 & ~n13109;
  assign n13111 = controllable_DEQ & ~n13110;
  assign n13112 = ~n10655 & ~n13101;
  assign n13113 = ~controllable_DEQ & ~n13112;
  assign n13114 = ~n13111 & ~n13113;
  assign n13115 = ~i_FULL & ~n13114;
  assign n13116 = ~n13105 & ~n13115;
  assign n13117 = i_nEMPTY & ~n13116;
  assign n13118 = ~n8166 & ~n9951;
  assign n13119 = ~controllable_BtoR_REQ0 & ~n13118;
  assign n13120 = ~controllable_BtoR_REQ0 & ~n13119;
  assign n13121 = ~i_RtoB_ACK0 & ~n13120;
  assign n13122 = ~i_RtoB_ACK0 & ~n13121;
  assign n13123 = controllable_DEQ & ~n13122;
  assign n13124 = ~n10681 & ~n13091;
  assign n13125 = ~controllable_DEQ & ~n13124;
  assign n13126 = ~n13123 & ~n13125;
  assign n13127 = i_FULL & ~n13126;
  assign n13128 = ~n8114 & ~n9973;
  assign n13129 = ~controllable_BtoR_REQ0 & ~n13128;
  assign n13130 = ~controllable_BtoR_REQ0 & ~n13129;
  assign n13131 = ~i_RtoB_ACK0 & ~n13130;
  assign n13132 = ~i_RtoB_ACK0 & ~n13131;
  assign n13133 = controllable_DEQ & ~n13132;
  assign n13134 = ~n10701 & ~n13091;
  assign n13135 = ~controllable_DEQ & ~n13134;
  assign n13136 = ~n13133 & ~n13135;
  assign n13137 = ~i_FULL & ~n13136;
  assign n13138 = ~n13127 & ~n13137;
  assign n13139 = ~i_nEMPTY & ~n13138;
  assign n13140 = ~n13117 & ~n13139;
  assign n13141 = ~controllable_BtoS_ACK0 & ~n13140;
  assign n13142 = ~n13087 & ~n13141;
  assign n13143 = n4465 & ~n13142;
  assign n13144 = ~n10876 & ~n13143;
  assign n13145 = ~i_StoB_REQ10 & ~n13144;
  assign n13146 = ~n13033 & ~n13145;
  assign n13147 = ~controllable_BtoS_ACK10 & ~n13146;
  assign n13148 = ~n12857 & ~n13147;
  assign n13149 = ~n4464 & ~n13148;
  assign n13150 = ~n12789 & ~n13149;
  assign n13151 = ~n4463 & ~n13150;
  assign n13152 = ~n12155 & ~n13151;
  assign n13153 = ~n4462 & ~n13152;
  assign n13154 = ~n11130 & ~n13153;
  assign n13155 = n4461 & ~n13154;
  assign n13156 = ~n5040 & ~n8763;
  assign n13157 = ~controllable_BtoR_REQ0 & ~n13156;
  assign n13158 = ~controllable_BtoR_REQ0 & ~n13157;
  assign n13159 = ~i_RtoB_ACK0 & ~n13158;
  assign n13160 = ~n5031 & ~n13159;
  assign n13161 = controllable_DEQ & ~n13160;
  assign n13162 = ~n5054 & ~n8786;
  assign n13163 = ~controllable_DEQ & ~n13162;
  assign n13164 = ~n13161 & ~n13163;
  assign n13165 = i_nEMPTY & ~n13164;
  assign n13166 = ~n5031 & ~n8823;
  assign n13167 = ~controllable_DEQ & ~n13166;
  assign n13168 = ~n5076 & ~n13167;
  assign n13169 = i_FULL & ~n13168;
  assign n13170 = ~controllable_BtoR_REQ1 & ~n5036;
  assign n13171 = ~n8763 & ~n13170;
  assign n13172 = ~controllable_BtoR_REQ0 & ~n13171;
  assign n13173 = ~controllable_BtoR_REQ0 & ~n13172;
  assign n13174 = ~i_RtoB_ACK0 & ~n13173;
  assign n13175 = ~n5031 & ~n13174;
  assign n13176 = ~controllable_DEQ & ~n13175;
  assign n13177 = ~n5091 & ~n13176;
  assign n13178 = ~i_FULL & ~n13177;
  assign n13179 = ~n13169 & ~n13178;
  assign n13180 = ~i_nEMPTY & ~n13179;
  assign n13181 = ~n13165 & ~n13180;
  assign n13182 = controllable_BtoS_ACK0 & ~n13181;
  assign n13183 = ~n5137 & ~n8863;
  assign n13184 = ~controllable_BtoR_REQ0 & ~n13183;
  assign n13185 = ~controllable_BtoR_REQ0 & ~n13184;
  assign n13186 = ~i_RtoB_ACK0 & ~n13185;
  assign n13187 = ~n5128 & ~n13186;
  assign n13188 = controllable_DEQ & ~n13187;
  assign n13189 = ~n5151 & ~n8889;
  assign n13190 = ~controllable_DEQ & ~n13189;
  assign n13191 = ~n13188 & ~n13190;
  assign n13192 = i_nEMPTY & ~n13191;
  assign n13193 = ~n5128 & ~n8930;
  assign n13194 = ~controllable_DEQ & ~n13193;
  assign n13195 = ~n5173 & ~n13194;
  assign n13196 = i_FULL & ~n13195;
  assign n13197 = ~controllable_BtoR_REQ1 & ~n5133;
  assign n13198 = ~n8863 & ~n13197;
  assign n13199 = ~controllable_BtoR_REQ0 & ~n13198;
  assign n13200 = ~controllable_BtoR_REQ0 & ~n13199;
  assign n13201 = ~i_RtoB_ACK0 & ~n13200;
  assign n13202 = ~n5128 & ~n13201;
  assign n13203 = ~controllable_DEQ & ~n13202;
  assign n13204 = ~n5188 & ~n13203;
  assign n13205 = ~i_FULL & ~n13204;
  assign n13206 = ~n13196 & ~n13205;
  assign n13207 = ~i_nEMPTY & ~n13206;
  assign n13208 = ~n13192 & ~n13207;
  assign n13209 = ~controllable_BtoS_ACK0 & ~n13208;
  assign n13210 = ~n13182 & ~n13209;
  assign n13211 = n4465 & ~n13210;
  assign n13212 = ~n5351 & ~n8972;
  assign n13213 = ~controllable_BtoR_REQ0 & ~n13212;
  assign n13214 = ~controllable_BtoR_REQ0 & ~n13213;
  assign n13215 = ~i_RtoB_ACK0 & ~n13214;
  assign n13216 = ~n5342 & ~n13215;
  assign n13217 = controllable_DEQ & ~n13216;
  assign n13218 = ~n5365 & ~n8995;
  assign n13219 = ~controllable_DEQ & ~n13218;
  assign n13220 = ~n13217 & ~n13219;
  assign n13221 = i_nEMPTY & ~n13220;
  assign n13222 = ~n5342 & ~n9032;
  assign n13223 = ~controllable_DEQ & ~n13222;
  assign n13224 = ~n5387 & ~n13223;
  assign n13225 = i_FULL & ~n13224;
  assign n13226 = ~controllable_BtoR_REQ1 & ~n5347;
  assign n13227 = ~n8972 & ~n13226;
  assign n13228 = ~controllable_BtoR_REQ0 & ~n13227;
  assign n13229 = ~controllable_BtoR_REQ0 & ~n13228;
  assign n13230 = ~i_RtoB_ACK0 & ~n13229;
  assign n13231 = ~n5342 & ~n13230;
  assign n13232 = ~controllable_DEQ & ~n13231;
  assign n13233 = ~n5402 & ~n13232;
  assign n13234 = ~i_FULL & ~n13233;
  assign n13235 = ~n13225 & ~n13234;
  assign n13236 = ~i_nEMPTY & ~n13235;
  assign n13237 = ~n13221 & ~n13236;
  assign n13238 = ~controllable_BtoS_ACK0 & ~n13237;
  assign n13239 = ~n5307 & ~n13238;
  assign n13240 = ~n4465 & ~n13239;
  assign n13241 = ~n13211 & ~n13240;
  assign n13242 = i_StoB_REQ10 & ~n13241;
  assign n13243 = ~n6765 & ~n9291;
  assign n13244 = i_RtoB_ACK1 & ~n13243;
  assign n13245 = ~n6770 & ~n13244;
  assign n13246 = controllable_BtoR_REQ1 & ~n13245;
  assign n13247 = ~n6778 & ~n13246;
  assign n13248 = ~controllable_BtoR_REQ0 & ~n13247;
  assign n13249 = ~controllable_BtoR_REQ0 & ~n13248;
  assign n13250 = ~i_RtoB_ACK0 & ~n13249;
  assign n13251 = ~n6585 & ~n13250;
  assign n13252 = controllable_DEQ & ~n13251;
  assign n13253 = i_RtoB_ACK1 & ~n9290;
  assign n13254 = ~n6796 & ~n13253;
  assign n13255 = controllable_BtoR_REQ1 & ~n13254;
  assign n13256 = ~n6798 & ~n13255;
  assign n13257 = ~controllable_BtoR_REQ0 & ~n13256;
  assign n13258 = ~controllable_BtoR_REQ0 & ~n13257;
  assign n13259 = ~i_RtoB_ACK0 & ~n13258;
  assign n13260 = ~n6793 & ~n13259;
  assign n13261 = ~controllable_DEQ & ~n13260;
  assign n13262 = ~n13252 & ~n13261;
  assign n13263 = i_FULL & ~n13262;
  assign n13264 = ~n6810 & ~n13244;
  assign n13265 = controllable_BtoR_REQ1 & ~n13264;
  assign n13266 = ~n6815 & ~n13265;
  assign n13267 = ~controllable_BtoR_REQ0 & ~n13266;
  assign n13268 = ~controllable_BtoR_REQ0 & ~n13267;
  assign n13269 = ~i_RtoB_ACK0 & ~n13268;
  assign n13270 = ~n6585 & ~n13269;
  assign n13271 = controllable_DEQ & ~n13270;
  assign n13272 = ~n6776 & ~n13253;
  assign n13273 = controllable_BtoR_REQ1 & ~n13272;
  assign n13274 = ~n6824 & ~n13273;
  assign n13275 = ~controllable_BtoR_REQ0 & ~n13274;
  assign n13276 = ~controllable_BtoR_REQ0 & ~n13275;
  assign n13277 = ~i_RtoB_ACK0 & ~n13276;
  assign n13278 = ~n6793 & ~n13277;
  assign n13279 = ~controllable_DEQ & ~n13278;
  assign n13280 = ~n13271 & ~n13279;
  assign n13281 = ~i_FULL & ~n13280;
  assign n13282 = ~n13263 & ~n13281;
  assign n13283 = i_nEMPTY & ~n13282;
  assign n13284 = i_RtoB_ACK1 & ~n9292;
  assign n13285 = ~n6853 & ~n13284;
  assign n13286 = controllable_BtoR_REQ1 & ~n13285;
  assign n13287 = ~n6855 & ~n13286;
  assign n13288 = ~controllable_BtoR_REQ0 & ~n13287;
  assign n13289 = ~controllable_BtoR_REQ0 & ~n13288;
  assign n13290 = ~i_RtoB_ACK0 & ~n13289;
  assign n13291 = ~n6585 & ~n13290;
  assign n13292 = ~controllable_DEQ & ~n13291;
  assign n13293 = ~n6850 & ~n13292;
  assign n13294 = i_FULL & ~n13293;
  assign n13295 = ~n6873 & ~n13246;
  assign n13296 = ~controllable_BtoR_REQ0 & ~n13295;
  assign n13297 = ~controllable_BtoR_REQ0 & ~n13296;
  assign n13298 = ~i_RtoB_ACK0 & ~n13297;
  assign n13299 = ~n6585 & ~n13298;
  assign n13300 = ~controllable_DEQ & ~n13299;
  assign n13301 = ~n6871 & ~n13300;
  assign n13302 = ~i_FULL & ~n13301;
  assign n13303 = ~n13294 & ~n13302;
  assign n13304 = ~i_nEMPTY & ~n13303;
  assign n13305 = ~n13283 & ~n13304;
  assign n13306 = controllable_BtoS_ACK0 & ~n13305;
  assign n13307 = ~n6931 & ~n9622;
  assign n13308 = i_RtoB_ACK1 & ~n13307;
  assign n13309 = ~n6936 & ~n13308;
  assign n13310 = controllable_BtoR_REQ1 & ~n13309;
  assign n13311 = ~n6944 & ~n13310;
  assign n13312 = ~controllable_BtoR_REQ0 & ~n13311;
  assign n13313 = ~controllable_BtoR_REQ0 & ~n13312;
  assign n13314 = ~i_RtoB_ACK0 & ~n13313;
  assign n13315 = ~n6924 & ~n13314;
  assign n13316 = controllable_DEQ & ~n13315;
  assign n13317 = i_RtoB_ACK1 & ~n9621;
  assign n13318 = ~n6962 & ~n13317;
  assign n13319 = controllable_BtoR_REQ1 & ~n13318;
  assign n13320 = ~n6964 & ~n13319;
  assign n13321 = ~controllable_BtoR_REQ0 & ~n13320;
  assign n13322 = ~controllable_BtoR_REQ0 & ~n13321;
  assign n13323 = ~i_RtoB_ACK0 & ~n13322;
  assign n13324 = ~n6959 & ~n13323;
  assign n13325 = ~controllable_DEQ & ~n13324;
  assign n13326 = ~n13316 & ~n13325;
  assign n13327 = i_FULL & ~n13326;
  assign n13328 = ~n6976 & ~n13308;
  assign n13329 = controllable_BtoR_REQ1 & ~n13328;
  assign n13330 = ~n6981 & ~n13329;
  assign n13331 = ~controllable_BtoR_REQ0 & ~n13330;
  assign n13332 = ~controllable_BtoR_REQ0 & ~n13331;
  assign n13333 = ~i_RtoB_ACK0 & ~n13332;
  assign n13334 = ~n6924 & ~n13333;
  assign n13335 = controllable_DEQ & ~n13334;
  assign n13336 = ~n6942 & ~n13317;
  assign n13337 = controllable_BtoR_REQ1 & ~n13336;
  assign n13338 = ~n6990 & ~n13337;
  assign n13339 = ~controllable_BtoR_REQ0 & ~n13338;
  assign n13340 = ~controllable_BtoR_REQ0 & ~n13339;
  assign n13341 = ~i_RtoB_ACK0 & ~n13340;
  assign n13342 = ~n6959 & ~n13341;
  assign n13343 = ~controllable_DEQ & ~n13342;
  assign n13344 = ~n13335 & ~n13343;
  assign n13345 = ~i_FULL & ~n13344;
  assign n13346 = ~n13327 & ~n13345;
  assign n13347 = i_nEMPTY & ~n13346;
  assign n13348 = i_RtoB_ACK1 & ~n9623;
  assign n13349 = ~n7019 & ~n13348;
  assign n13350 = controllable_BtoR_REQ1 & ~n13349;
  assign n13351 = ~n7021 & ~n13350;
  assign n13352 = ~controllable_BtoR_REQ0 & ~n13351;
  assign n13353 = ~controllable_BtoR_REQ0 & ~n13352;
  assign n13354 = ~i_RtoB_ACK0 & ~n13353;
  assign n13355 = ~n6924 & ~n13354;
  assign n13356 = ~controllable_DEQ & ~n13355;
  assign n13357 = ~n7016 & ~n13356;
  assign n13358 = i_FULL & ~n13357;
  assign n13359 = ~n7039 & ~n13310;
  assign n13360 = ~controllable_BtoR_REQ0 & ~n13359;
  assign n13361 = ~controllable_BtoR_REQ0 & ~n13360;
  assign n13362 = ~i_RtoB_ACK0 & ~n13361;
  assign n13363 = ~n6924 & ~n13362;
  assign n13364 = ~controllable_DEQ & ~n13363;
  assign n13365 = ~n7037 & ~n13364;
  assign n13366 = ~i_FULL & ~n13365;
  assign n13367 = ~n13358 & ~n13366;
  assign n13368 = ~i_nEMPTY & ~n13367;
  assign n13369 = ~n13347 & ~n13368;
  assign n13370 = ~controllable_BtoS_ACK0 & ~n13369;
  assign n13371 = ~n13306 & ~n13370;
  assign n13372 = n4465 & ~n13371;
  assign n13373 = ~n5238 & ~n9779;
  assign n13374 = i_RtoB_ACK1 & ~n13373;
  assign n13375 = ~n7098 & ~n13374;
  assign n13376 = controllable_BtoR_REQ1 & ~n13375;
  assign n13377 = ~n7104 & ~n13376;
  assign n13378 = ~controllable_BtoR_REQ0 & ~n13377;
  assign n13379 = ~controllable_BtoR_REQ0 & ~n13378;
  assign n13380 = ~i_RtoB_ACK0 & ~n13379;
  assign n13381 = ~n7093 & ~n13380;
  assign n13382 = controllable_DEQ & ~n13381;
  assign n13383 = i_RtoB_ACK1 & ~n9778;
  assign n13384 = ~n7102 & ~n13383;
  assign n13385 = controllable_BtoR_REQ1 & ~n13384;
  assign n13386 = ~n7115 & ~n13385;
  assign n13387 = ~controllable_BtoR_REQ0 & ~n13386;
  assign n13388 = ~controllable_BtoR_REQ0 & ~n13387;
  assign n13389 = ~i_RtoB_ACK0 & ~n13388;
  assign n13390 = ~n7119 & ~n13389;
  assign n13391 = ~controllable_DEQ & ~n13390;
  assign n13392 = ~n13382 & ~n13391;
  assign n13393 = i_nEMPTY & ~n13392;
  assign n13394 = i_RtoB_ACK1 & ~n9780;
  assign n13395 = ~n7546 & ~n13394;
  assign n13396 = controllable_BtoR_REQ1 & ~n13395;
  assign n13397 = ~n7089 & ~n13396;
  assign n13398 = ~controllable_BtoR_REQ0 & ~n13397;
  assign n13399 = ~controllable_BtoR_REQ0 & ~n13398;
  assign n13400 = ~i_RtoB_ACK0 & ~n13399;
  assign n13401 = ~n7093 & ~n13400;
  assign n13402 = ~controllable_DEQ & ~n13401;
  assign n13403 = ~n7142 & ~n13402;
  assign n13404 = i_FULL & ~n13403;
  assign n13405 = ~n7159 & ~n13376;
  assign n13406 = ~controllable_BtoR_REQ0 & ~n13405;
  assign n13407 = ~controllable_BtoR_REQ0 & ~n13406;
  assign n13408 = ~i_RtoB_ACK0 & ~n13407;
  assign n13409 = ~n7093 & ~n13408;
  assign n13410 = ~controllable_DEQ & ~n13409;
  assign n13411 = ~n7157 & ~n13410;
  assign n13412 = ~i_FULL & ~n13411;
  assign n13413 = ~n13404 & ~n13412;
  assign n13414 = ~i_nEMPTY & ~n13413;
  assign n13415 = ~n13393 & ~n13414;
  assign n13416 = controllable_BtoS_ACK0 & ~n13415;
  assign n13417 = ~n7270 & ~n9881;
  assign n13418 = ~controllable_BtoR_REQ0 & ~n13417;
  assign n13419 = ~controllable_BtoR_REQ0 & ~n13418;
  assign n13420 = ~i_RtoB_ACK0 & ~n13419;
  assign n13421 = ~n7246 & ~n13420;
  assign n13422 = controllable_DEQ & ~n13421;
  assign n13423 = ~n7290 & ~n9912;
  assign n13424 = ~controllable_BtoR_REQ0 & ~n13423;
  assign n13425 = ~controllable_BtoR_REQ0 & ~n13424;
  assign n13426 = ~i_RtoB_ACK0 & ~n13425;
  assign n13427 = ~n7285 & ~n13426;
  assign n13428 = ~controllable_DEQ & ~n13427;
  assign n13429 = ~n13422 & ~n13428;
  assign n13430 = i_FULL & ~n13429;
  assign n13431 = ~n7307 & ~n9925;
  assign n13432 = ~controllable_BtoR_REQ0 & ~n13431;
  assign n13433 = ~controllable_BtoR_REQ0 & ~n13432;
  assign n13434 = ~i_RtoB_ACK0 & ~n13433;
  assign n13435 = ~n7246 & ~n13434;
  assign n13436 = controllable_DEQ & ~n13435;
  assign n13437 = ~n7316 & ~n9935;
  assign n13438 = ~controllable_BtoR_REQ0 & ~n13437;
  assign n13439 = ~controllable_BtoR_REQ0 & ~n13438;
  assign n13440 = ~i_RtoB_ACK0 & ~n13439;
  assign n13441 = ~n7285 & ~n13440;
  assign n13442 = ~controllable_DEQ & ~n13441;
  assign n13443 = ~n13436 & ~n13442;
  assign n13444 = ~i_FULL & ~n13443;
  assign n13445 = ~n13430 & ~n13444;
  assign n13446 = i_nEMPTY & ~n13445;
  assign n13447 = ~n7347 & ~n9959;
  assign n13448 = ~controllable_BtoR_REQ0 & ~n13447;
  assign n13449 = ~controllable_BtoR_REQ0 & ~n13448;
  assign n13450 = ~i_RtoB_ACK0 & ~n13449;
  assign n13451 = ~n7246 & ~n13450;
  assign n13452 = ~controllable_DEQ & ~n13451;
  assign n13453 = ~n7342 & ~n13452;
  assign n13454 = i_FULL & ~n13453;
  assign n13455 = ~n7365 & ~n9881;
  assign n13456 = ~controllable_BtoR_REQ0 & ~n13455;
  assign n13457 = ~controllable_BtoR_REQ0 & ~n13456;
  assign n13458 = ~i_RtoB_ACK0 & ~n13457;
  assign n13459 = ~n7246 & ~n13458;
  assign n13460 = ~controllable_DEQ & ~n13459;
  assign n13461 = ~n7363 & ~n13460;
  assign n13462 = ~i_FULL & ~n13461;
  assign n13463 = ~n13454 & ~n13462;
  assign n13464 = ~i_nEMPTY & ~n13463;
  assign n13465 = ~n13446 & ~n13464;
  assign n13466 = ~controllable_BtoS_ACK0 & ~n13465;
  assign n13467 = ~n13416 & ~n13466;
  assign n13468 = ~n4465 & ~n13467;
  assign n13469 = ~n13372 & ~n13468;
  assign n13470 = ~i_StoB_REQ10 & ~n13469;
  assign n13471 = ~n13242 & ~n13470;
  assign n13472 = controllable_BtoS_ACK10 & ~n13471;
  assign n13473 = ~n6778 & ~n10011;
  assign n13474 = ~controllable_BtoR_REQ0 & ~n13473;
  assign n13475 = ~controllable_BtoR_REQ0 & ~n13474;
  assign n13476 = ~i_RtoB_ACK0 & ~n13475;
  assign n13477 = ~n7398 & ~n13476;
  assign n13478 = controllable_DEQ & ~n13477;
  assign n13479 = ~n6798 & ~n9519;
  assign n13480 = ~controllable_BtoR_REQ0 & ~n13479;
  assign n13481 = ~controllable_BtoR_REQ0 & ~n13480;
  assign n13482 = ~i_RtoB_ACK0 & ~n13481;
  assign n13483 = ~n7416 & ~n13482;
  assign n13484 = ~controllable_DEQ & ~n13483;
  assign n13485 = ~n13478 & ~n13484;
  assign n13486 = i_FULL & ~n13485;
  assign n13487 = ~n6815 & ~n10031;
  assign n13488 = ~controllable_BtoR_REQ0 & ~n13487;
  assign n13489 = ~controllable_BtoR_REQ0 & ~n13488;
  assign n13490 = ~i_RtoB_ACK0 & ~n13489;
  assign n13491 = ~n7398 & ~n13490;
  assign n13492 = controllable_DEQ & ~n13491;
  assign n13493 = ~n6824 & ~n9544;
  assign n13494 = ~controllable_BtoR_REQ0 & ~n13493;
  assign n13495 = ~controllable_BtoR_REQ0 & ~n13494;
  assign n13496 = ~i_RtoB_ACK0 & ~n13495;
  assign n13497 = ~n7416 & ~n13496;
  assign n13498 = ~controllable_DEQ & ~n13497;
  assign n13499 = ~n13492 & ~n13498;
  assign n13500 = ~i_FULL & ~n13499;
  assign n13501 = ~n13486 & ~n13500;
  assign n13502 = i_nEMPTY & ~n13501;
  assign n13503 = ~n6855 & ~n9573;
  assign n13504 = ~controllable_BtoR_REQ0 & ~n13503;
  assign n13505 = ~controllable_BtoR_REQ0 & ~n13504;
  assign n13506 = ~i_RtoB_ACK0 & ~n13505;
  assign n13507 = ~n7398 & ~n13506;
  assign n13508 = ~controllable_DEQ & ~n13507;
  assign n13509 = ~n7446 & ~n13508;
  assign n13510 = i_FULL & ~n13509;
  assign n13511 = ~controllable_DEQ & ~n13477;
  assign n13512 = ~n7456 & ~n13511;
  assign n13513 = ~i_FULL & ~n13512;
  assign n13514 = ~n13510 & ~n13513;
  assign n13515 = ~i_nEMPTY & ~n13514;
  assign n13516 = ~n13502 & ~n13515;
  assign n13517 = controllable_BtoS_ACK0 & ~n13516;
  assign n13518 = ~n6944 & ~n10084;
  assign n13519 = ~controllable_BtoR_REQ0 & ~n13518;
  assign n13520 = ~controllable_BtoR_REQ0 & ~n13519;
  assign n13521 = ~i_RtoB_ACK0 & ~n13520;
  assign n13522 = ~n7478 & ~n13521;
  assign n13523 = controllable_DEQ & ~n13522;
  assign n13524 = ~n6964 & ~n9666;
  assign n13525 = ~controllable_BtoR_REQ0 & ~n13524;
  assign n13526 = ~controllable_BtoR_REQ0 & ~n13525;
  assign n13527 = ~i_RtoB_ACK0 & ~n13526;
  assign n13528 = ~n7496 & ~n13527;
  assign n13529 = ~controllable_DEQ & ~n13528;
  assign n13530 = ~n13523 & ~n13529;
  assign n13531 = i_FULL & ~n13530;
  assign n13532 = ~n6981 & ~n10104;
  assign n13533 = ~controllable_BtoR_REQ0 & ~n13532;
  assign n13534 = ~controllable_BtoR_REQ0 & ~n13533;
  assign n13535 = ~i_RtoB_ACK0 & ~n13534;
  assign n13536 = ~n7478 & ~n13535;
  assign n13537 = controllable_DEQ & ~n13536;
  assign n13538 = ~n6990 & ~n9691;
  assign n13539 = ~controllable_BtoR_REQ0 & ~n13538;
  assign n13540 = ~controllable_BtoR_REQ0 & ~n13539;
  assign n13541 = ~i_RtoB_ACK0 & ~n13540;
  assign n13542 = ~n7496 & ~n13541;
  assign n13543 = ~controllable_DEQ & ~n13542;
  assign n13544 = ~n13537 & ~n13543;
  assign n13545 = ~i_FULL & ~n13544;
  assign n13546 = ~n13531 & ~n13545;
  assign n13547 = i_nEMPTY & ~n13546;
  assign n13548 = ~n7021 & ~n9720;
  assign n13549 = ~controllable_BtoR_REQ0 & ~n13548;
  assign n13550 = ~controllable_BtoR_REQ0 & ~n13549;
  assign n13551 = ~i_RtoB_ACK0 & ~n13550;
  assign n13552 = ~n7478 & ~n13551;
  assign n13553 = ~controllable_DEQ & ~n13552;
  assign n13554 = ~n7526 & ~n13553;
  assign n13555 = i_FULL & ~n13554;
  assign n13556 = ~controllable_DEQ & ~n13522;
  assign n13557 = ~n7536 & ~n13556;
  assign n13558 = ~i_FULL & ~n13557;
  assign n13559 = ~n13555 & ~n13558;
  assign n13560 = ~i_nEMPTY & ~n13559;
  assign n13561 = ~n13547 & ~n13560;
  assign n13562 = ~controllable_BtoS_ACK0 & ~n13561;
  assign n13563 = ~n13517 & ~n13562;
  assign n13564 = n4465 & ~n13563;
  assign n13565 = ~n7104 & ~n10151;
  assign n13566 = ~controllable_BtoR_REQ0 & ~n13565;
  assign n13567 = ~controllable_BtoR_REQ0 & ~n13566;
  assign n13568 = ~i_RtoB_ACK0 & ~n13567;
  assign n13569 = ~n7552 & ~n13568;
  assign n13570 = controllable_DEQ & ~n13569;
  assign n13571 = ~n7115 & ~n9812;
  assign n13572 = ~controllable_BtoR_REQ0 & ~n13571;
  assign n13573 = ~controllable_BtoR_REQ0 & ~n13572;
  assign n13574 = ~i_RtoB_ACK0 & ~n13573;
  assign n13575 = ~n7569 & ~n13574;
  assign n13576 = ~controllable_DEQ & ~n13575;
  assign n13577 = ~n13570 & ~n13576;
  assign n13578 = i_nEMPTY & ~n13577;
  assign n13579 = ~n7089 & ~n9835;
  assign n13580 = ~controllable_BtoR_REQ0 & ~n13579;
  assign n13581 = ~controllable_BtoR_REQ0 & ~n13580;
  assign n13582 = ~i_RtoB_ACK0 & ~n13581;
  assign n13583 = ~n7552 & ~n13582;
  assign n13584 = ~controllable_DEQ & ~n13583;
  assign n13585 = ~n7582 & ~n13584;
  assign n13586 = i_FULL & ~n13585;
  assign n13587 = ~controllable_DEQ & ~n13569;
  assign n13588 = ~n7592 & ~n13587;
  assign n13589 = ~i_FULL & ~n13588;
  assign n13590 = ~n13586 & ~n13589;
  assign n13591 = ~i_nEMPTY & ~n13590;
  assign n13592 = ~n13578 & ~n13591;
  assign n13593 = controllable_BtoS_ACK0 & ~n13592;
  assign n13594 = ~n7270 & ~n10198;
  assign n13595 = ~controllable_BtoR_REQ0 & ~n13594;
  assign n13596 = ~controllable_BtoR_REQ0 & ~n13595;
  assign n13597 = ~i_RtoB_ACK0 & ~n13596;
  assign n13598 = ~n7614 & ~n13597;
  assign n13599 = controllable_DEQ & ~n13598;
  assign n13600 = ~n7632 & ~n13426;
  assign n13601 = ~controllable_DEQ & ~n13600;
  assign n13602 = ~n13599 & ~n13601;
  assign n13603 = i_FULL & ~n13602;
  assign n13604 = ~n7307 & ~n10214;
  assign n13605 = ~controllable_BtoR_REQ0 & ~n13604;
  assign n13606 = ~controllable_BtoR_REQ0 & ~n13605;
  assign n13607 = ~i_RtoB_ACK0 & ~n13606;
  assign n13608 = ~n7614 & ~n13607;
  assign n13609 = controllable_DEQ & ~n13608;
  assign n13610 = ~n7632 & ~n13440;
  assign n13611 = ~controllable_DEQ & ~n13610;
  assign n13612 = ~n13609 & ~n13611;
  assign n13613 = ~i_FULL & ~n13612;
  assign n13614 = ~n13603 & ~n13613;
  assign n13615 = i_nEMPTY & ~n13614;
  assign n13616 = ~n7614 & ~n13450;
  assign n13617 = ~controllable_DEQ & ~n13616;
  assign n13618 = ~n7662 & ~n13617;
  assign n13619 = i_FULL & ~n13618;
  assign n13620 = ~controllable_DEQ & ~n13598;
  assign n13621 = ~n7672 & ~n13620;
  assign n13622 = ~i_FULL & ~n13621;
  assign n13623 = ~n13619 & ~n13622;
  assign n13624 = ~i_nEMPTY & ~n13623;
  assign n13625 = ~n13615 & ~n13624;
  assign n13626 = ~controllable_BtoS_ACK0 & ~n13625;
  assign n13627 = ~n13593 & ~n13626;
  assign n13628 = ~n4465 & ~n13627;
  assign n13629 = ~n13564 & ~n13628;
  assign n13630 = i_StoB_REQ10 & ~n13629;
  assign n13631 = ~n13470 & ~n13630;
  assign n13632 = ~controllable_BtoS_ACK10 & ~n13631;
  assign n13633 = ~n13472 & ~n13632;
  assign n13634 = n4464 & ~n13633;
  assign n13635 = ~n7718 & ~n10265;
  assign n13636 = ~controllable_BtoR_REQ0 & ~n13635;
  assign n13637 = ~controllable_BtoR_REQ0 & ~n13636;
  assign n13638 = ~i_RtoB_ACK0 & ~n13637;
  assign n13639 = ~n7709 & ~n13638;
  assign n13640 = controllable_DEQ & ~n13639;
  assign n13641 = ~n7732 & ~n10288;
  assign n13642 = ~controllable_DEQ & ~n13641;
  assign n13643 = ~n13640 & ~n13642;
  assign n13644 = i_nEMPTY & ~n13643;
  assign n13645 = ~n7709 & ~n10325;
  assign n13646 = ~controllable_DEQ & ~n13645;
  assign n13647 = ~n7754 & ~n13646;
  assign n13648 = i_FULL & ~n13647;
  assign n13649 = ~controllable_BtoR_REQ1 & ~n7714;
  assign n13650 = ~n10265 & ~n13649;
  assign n13651 = ~controllable_BtoR_REQ0 & ~n13650;
  assign n13652 = ~controllable_BtoR_REQ0 & ~n13651;
  assign n13653 = ~i_RtoB_ACK0 & ~n13652;
  assign n13654 = ~n7709 & ~n13653;
  assign n13655 = ~controllable_DEQ & ~n13654;
  assign n13656 = ~n7769 & ~n13655;
  assign n13657 = ~i_FULL & ~n13656;
  assign n13658 = ~n13648 & ~n13657;
  assign n13659 = ~i_nEMPTY & ~n13658;
  assign n13660 = ~n13644 & ~n13659;
  assign n13661 = controllable_BtoS_ACK0 & ~n13660;
  assign n13662 = ~n7810 & ~n10359;
  assign n13663 = ~controllable_BtoR_REQ0 & ~n13662;
  assign n13664 = ~controllable_BtoR_REQ0 & ~n13663;
  assign n13665 = ~i_RtoB_ACK0 & ~n13664;
  assign n13666 = ~n7801 & ~n13665;
  assign n13667 = controllable_DEQ & ~n13666;
  assign n13668 = ~n7824 & ~n10382;
  assign n13669 = ~controllable_DEQ & ~n13668;
  assign n13670 = ~n13667 & ~n13669;
  assign n13671 = i_nEMPTY & ~n13670;
  assign n13672 = ~n7801 & ~n10419;
  assign n13673 = ~controllable_DEQ & ~n13672;
  assign n13674 = ~n7846 & ~n13673;
  assign n13675 = i_FULL & ~n13674;
  assign n13676 = ~controllable_BtoR_REQ1 & ~n7806;
  assign n13677 = ~n10359 & ~n13676;
  assign n13678 = ~controllable_BtoR_REQ0 & ~n13677;
  assign n13679 = ~controllable_BtoR_REQ0 & ~n13678;
  assign n13680 = ~i_RtoB_ACK0 & ~n13679;
  assign n13681 = ~n7801 & ~n13680;
  assign n13682 = ~controllable_DEQ & ~n13681;
  assign n13683 = ~n7861 & ~n13682;
  assign n13684 = ~i_FULL & ~n13683;
  assign n13685 = ~n13675 & ~n13684;
  assign n13686 = ~i_nEMPTY & ~n13685;
  assign n13687 = ~n13671 & ~n13686;
  assign n13688 = ~controllable_BtoS_ACK0 & ~n13687;
  assign n13689 = ~n13661 & ~n13688;
  assign n13690 = n4465 & ~n13689;
  assign n13691 = ~n5307 & ~n13688;
  assign n13692 = ~n4465 & ~n13691;
  assign n13693 = ~n13690 & ~n13692;
  assign n13694 = i_StoB_REQ10 & ~n13693;
  assign n13695 = ~n7927 & ~n10458;
  assign n13696 = i_RtoB_ACK1 & ~n13695;
  assign n13697 = ~n7932 & ~n13696;
  assign n13698 = controllable_BtoR_REQ1 & ~n13697;
  assign n13699 = ~n7940 & ~n13698;
  assign n13700 = ~controllable_BtoR_REQ0 & ~n13699;
  assign n13701 = ~controllable_BtoR_REQ0 & ~n13700;
  assign n13702 = ~i_RtoB_ACK0 & ~n13701;
  assign n13703 = ~n7921 & ~n13702;
  assign n13704 = controllable_DEQ & ~n13703;
  assign n13705 = i_RtoB_ACK1 & ~n10457;
  assign n13706 = ~n7958 & ~n13705;
  assign n13707 = controllable_BtoR_REQ1 & ~n13706;
  assign n13708 = ~n7960 & ~n13707;
  assign n13709 = ~controllable_BtoR_REQ0 & ~n13708;
  assign n13710 = ~controllable_BtoR_REQ0 & ~n13709;
  assign n13711 = ~i_RtoB_ACK0 & ~n13710;
  assign n13712 = ~n7955 & ~n13711;
  assign n13713 = ~controllable_DEQ & ~n13712;
  assign n13714 = ~n13704 & ~n13713;
  assign n13715 = i_FULL & ~n13714;
  assign n13716 = ~n7972 & ~n13696;
  assign n13717 = controllable_BtoR_REQ1 & ~n13716;
  assign n13718 = ~n7977 & ~n13717;
  assign n13719 = ~controllable_BtoR_REQ0 & ~n13718;
  assign n13720 = ~controllable_BtoR_REQ0 & ~n13719;
  assign n13721 = ~i_RtoB_ACK0 & ~n13720;
  assign n13722 = ~n7921 & ~n13721;
  assign n13723 = controllable_DEQ & ~n13722;
  assign n13724 = ~n7938 & ~n13705;
  assign n13725 = controllable_BtoR_REQ1 & ~n13724;
  assign n13726 = ~n7986 & ~n13725;
  assign n13727 = ~controllable_BtoR_REQ0 & ~n13726;
  assign n13728 = ~controllable_BtoR_REQ0 & ~n13727;
  assign n13729 = ~i_RtoB_ACK0 & ~n13728;
  assign n13730 = ~n7955 & ~n13729;
  assign n13731 = ~controllable_DEQ & ~n13730;
  assign n13732 = ~n13723 & ~n13731;
  assign n13733 = ~i_FULL & ~n13732;
  assign n13734 = ~n13715 & ~n13733;
  assign n13735 = i_nEMPTY & ~n13734;
  assign n13736 = i_RtoB_ACK1 & ~n10459;
  assign n13737 = ~n8015 & ~n13736;
  assign n13738 = controllable_BtoR_REQ1 & ~n13737;
  assign n13739 = ~n8017 & ~n13738;
  assign n13740 = ~controllable_BtoR_REQ0 & ~n13739;
  assign n13741 = ~controllable_BtoR_REQ0 & ~n13740;
  assign n13742 = ~i_RtoB_ACK0 & ~n13741;
  assign n13743 = ~n7921 & ~n13742;
  assign n13744 = ~controllable_DEQ & ~n13743;
  assign n13745 = ~n8012 & ~n13744;
  assign n13746 = i_FULL & ~n13745;
  assign n13747 = ~n8035 & ~n13698;
  assign n13748 = ~controllable_BtoR_REQ0 & ~n13747;
  assign n13749 = ~controllable_BtoR_REQ0 & ~n13748;
  assign n13750 = ~i_RtoB_ACK0 & ~n13749;
  assign n13751 = ~n7921 & ~n13750;
  assign n13752 = ~controllable_DEQ & ~n13751;
  assign n13753 = ~n8033 & ~n13752;
  assign n13754 = ~i_FULL & ~n13753;
  assign n13755 = ~n13746 & ~n13754;
  assign n13756 = ~i_nEMPTY & ~n13755;
  assign n13757 = ~n13735 & ~n13756;
  assign n13758 = controllable_BtoS_ACK0 & ~n13757;
  assign n13759 = ~n8091 & ~n10588;
  assign n13760 = i_RtoB_ACK1 & ~n13759;
  assign n13761 = ~n8096 & ~n13760;
  assign n13762 = controllable_BtoR_REQ1 & ~n13761;
  assign n13763 = ~n8104 & ~n13762;
  assign n13764 = ~controllable_BtoR_REQ0 & ~n13763;
  assign n13765 = ~controllable_BtoR_REQ0 & ~n13764;
  assign n13766 = ~i_RtoB_ACK0 & ~n13765;
  assign n13767 = ~n8088 & ~n13766;
  assign n13768 = controllable_DEQ & ~n13767;
  assign n13769 = i_RtoB_ACK1 & ~n10587;
  assign n13770 = ~n8122 & ~n13769;
  assign n13771 = controllable_BtoR_REQ1 & ~n13770;
  assign n13772 = ~n8124 & ~n13771;
  assign n13773 = ~controllable_BtoR_REQ0 & ~n13772;
  assign n13774 = ~controllable_BtoR_REQ0 & ~n13773;
  assign n13775 = ~i_RtoB_ACK0 & ~n13774;
  assign n13776 = ~n8119 & ~n13775;
  assign n13777 = ~controllable_DEQ & ~n13776;
  assign n13778 = ~n13768 & ~n13777;
  assign n13779 = i_FULL & ~n13778;
  assign n13780 = ~n8136 & ~n13760;
  assign n13781 = controllable_BtoR_REQ1 & ~n13780;
  assign n13782 = ~n8141 & ~n13781;
  assign n13783 = ~controllable_BtoR_REQ0 & ~n13782;
  assign n13784 = ~controllable_BtoR_REQ0 & ~n13783;
  assign n13785 = ~i_RtoB_ACK0 & ~n13784;
  assign n13786 = ~n8088 & ~n13785;
  assign n13787 = controllable_DEQ & ~n13786;
  assign n13788 = ~n8102 & ~n13769;
  assign n13789 = controllable_BtoR_REQ1 & ~n13788;
  assign n13790 = ~n8150 & ~n13789;
  assign n13791 = ~controllable_BtoR_REQ0 & ~n13790;
  assign n13792 = ~controllable_BtoR_REQ0 & ~n13791;
  assign n13793 = ~i_RtoB_ACK0 & ~n13792;
  assign n13794 = ~n8119 & ~n13793;
  assign n13795 = ~controllable_DEQ & ~n13794;
  assign n13796 = ~n13787 & ~n13795;
  assign n13797 = ~i_FULL & ~n13796;
  assign n13798 = ~n13779 & ~n13797;
  assign n13799 = i_nEMPTY & ~n13798;
  assign n13800 = i_RtoB_ACK1 & ~n10589;
  assign n13801 = ~n8179 & ~n13800;
  assign n13802 = controllable_BtoR_REQ1 & ~n13801;
  assign n13803 = ~n8181 & ~n13802;
  assign n13804 = ~controllable_BtoR_REQ0 & ~n13803;
  assign n13805 = ~controllable_BtoR_REQ0 & ~n13804;
  assign n13806 = ~i_RtoB_ACK0 & ~n13805;
  assign n13807 = ~n8088 & ~n13806;
  assign n13808 = ~controllable_DEQ & ~n13807;
  assign n13809 = ~n8176 & ~n13808;
  assign n13810 = i_FULL & ~n13809;
  assign n13811 = ~n8199 & ~n13762;
  assign n13812 = ~controllable_BtoR_REQ0 & ~n13811;
  assign n13813 = ~controllable_BtoR_REQ0 & ~n13812;
  assign n13814 = ~i_RtoB_ACK0 & ~n13813;
  assign n13815 = ~n8088 & ~n13814;
  assign n13816 = ~controllable_DEQ & ~n13815;
  assign n13817 = ~n8197 & ~n13816;
  assign n13818 = ~i_FULL & ~n13817;
  assign n13819 = ~n13810 & ~n13818;
  assign n13820 = ~i_nEMPTY & ~n13819;
  assign n13821 = ~n13799 & ~n13820;
  assign n13822 = ~controllable_BtoS_ACK0 & ~n13821;
  assign n13823 = ~n13758 & ~n13822;
  assign n13824 = n4465 & ~n13823;
  assign n13825 = ~n8242 & ~n10719;
  assign n13826 = ~controllable_BtoR_REQ0 & ~n13825;
  assign n13827 = ~controllable_BtoR_REQ0 & ~n13826;
  assign n13828 = ~i_RtoB_ACK0 & ~n13827;
  assign n13829 = ~n8231 & ~n13828;
  assign n13830 = controllable_DEQ & ~n13829;
  assign n13831 = ~n8252 & ~n10736;
  assign n13832 = ~controllable_BtoR_REQ0 & ~n13831;
  assign n13833 = ~controllable_BtoR_REQ0 & ~n13832;
  assign n13834 = ~i_RtoB_ACK0 & ~n13833;
  assign n13835 = ~n8256 & ~n13834;
  assign n13836 = ~controllable_DEQ & ~n13835;
  assign n13837 = ~n13830 & ~n13836;
  assign n13838 = i_nEMPTY & ~n13837;
  assign n13839 = ~n8227 & ~n10752;
  assign n13840 = ~controllable_BtoR_REQ0 & ~n13839;
  assign n13841 = ~controllable_BtoR_REQ0 & ~n13840;
  assign n13842 = ~i_RtoB_ACK0 & ~n13841;
  assign n13843 = ~n8231 & ~n13842;
  assign n13844 = ~controllable_DEQ & ~n13843;
  assign n13845 = ~n8278 & ~n13844;
  assign n13846 = i_FULL & ~n13845;
  assign n13847 = ~n8295 & ~n10719;
  assign n13848 = ~controllable_BtoR_REQ0 & ~n13847;
  assign n13849 = ~controllable_BtoR_REQ0 & ~n13848;
  assign n13850 = ~i_RtoB_ACK0 & ~n13849;
  assign n13851 = ~n8231 & ~n13850;
  assign n13852 = ~controllable_DEQ & ~n13851;
  assign n13853 = ~n8293 & ~n13852;
  assign n13854 = ~i_FULL & ~n13853;
  assign n13855 = ~n13846 & ~n13854;
  assign n13856 = ~i_nEMPTY & ~n13855;
  assign n13857 = ~n13838 & ~n13856;
  assign n13858 = controllable_BtoS_ACK0 & ~n13857;
  assign n13859 = ~n8345 & ~n10790;
  assign n13860 = ~controllable_BtoR_REQ0 & ~n13859;
  assign n13861 = ~controllable_BtoR_REQ0 & ~n13860;
  assign n13862 = ~i_RtoB_ACK0 & ~n13861;
  assign n13863 = ~n8331 & ~n13862;
  assign n13864 = controllable_DEQ & ~n13863;
  assign n13865 = ~n8363 & ~n10622;
  assign n13866 = ~controllable_BtoR_REQ0 & ~n13865;
  assign n13867 = ~controllable_BtoR_REQ0 & ~n13866;
  assign n13868 = ~i_RtoB_ACK0 & ~n13867;
  assign n13869 = ~n8360 & ~n13868;
  assign n13870 = ~controllable_DEQ & ~n13869;
  assign n13871 = ~n13864 & ~n13870;
  assign n13872 = i_FULL & ~n13871;
  assign n13873 = ~n8380 & ~n10816;
  assign n13874 = ~controllable_BtoR_REQ0 & ~n13873;
  assign n13875 = ~controllable_BtoR_REQ0 & ~n13874;
  assign n13876 = ~i_RtoB_ACK0 & ~n13875;
  assign n13877 = ~n8331 & ~n13876;
  assign n13878 = controllable_DEQ & ~n13877;
  assign n13879 = ~n8389 & ~n10826;
  assign n13880 = ~controllable_BtoR_REQ0 & ~n13879;
  assign n13881 = ~controllable_BtoR_REQ0 & ~n13880;
  assign n13882 = ~i_RtoB_ACK0 & ~n13881;
  assign n13883 = ~n8360 & ~n13882;
  assign n13884 = ~controllable_DEQ & ~n13883;
  assign n13885 = ~n13878 & ~n13884;
  assign n13886 = ~i_FULL & ~n13885;
  assign n13887 = ~n13872 & ~n13886;
  assign n13888 = i_nEMPTY & ~n13887;
  assign n13889 = ~n8417 & ~n10673;
  assign n13890 = ~controllable_BtoR_REQ0 & ~n13889;
  assign n13891 = ~controllable_BtoR_REQ0 & ~n13890;
  assign n13892 = ~i_RtoB_ACK0 & ~n13891;
  assign n13893 = ~n8331 & ~n13892;
  assign n13894 = ~controllable_DEQ & ~n13893;
  assign n13895 = ~n8415 & ~n13894;
  assign n13896 = i_FULL & ~n13895;
  assign n13897 = ~n8435 & ~n10790;
  assign n13898 = ~controllable_BtoR_REQ0 & ~n13897;
  assign n13899 = ~controllable_BtoR_REQ0 & ~n13898;
  assign n13900 = ~i_RtoB_ACK0 & ~n13899;
  assign n13901 = ~n8331 & ~n13900;
  assign n13902 = ~controllable_DEQ & ~n13901;
  assign n13903 = ~n8433 & ~n13902;
  assign n13904 = ~i_FULL & ~n13903;
  assign n13905 = ~n13896 & ~n13904;
  assign n13906 = ~i_nEMPTY & ~n13905;
  assign n13907 = ~n13888 & ~n13906;
  assign n13908 = ~controllable_BtoS_ACK0 & ~n13907;
  assign n13909 = ~n13858 & ~n13908;
  assign n13910 = ~n4465 & ~n13909;
  assign n13911 = ~n13824 & ~n13910;
  assign n13912 = ~i_StoB_REQ10 & ~n13911;
  assign n13913 = ~n13694 & ~n13912;
  assign n13914 = controllable_BtoS_ACK10 & ~n13913;
  assign n13915 = ~n7940 & ~n10890;
  assign n13916 = ~controllable_BtoR_REQ0 & ~n13915;
  assign n13917 = ~controllable_BtoR_REQ0 & ~n13916;
  assign n13918 = ~i_RtoB_ACK0 & ~n13917;
  assign n13919 = ~n8468 & ~n13918;
  assign n13920 = controllable_DEQ & ~n13919;
  assign n13921 = ~n7960 & ~n10495;
  assign n13922 = ~controllable_BtoR_REQ0 & ~n13921;
  assign n13923 = ~controllable_BtoR_REQ0 & ~n13922;
  assign n13924 = ~i_RtoB_ACK0 & ~n13923;
  assign n13925 = ~n8486 & ~n13924;
  assign n13926 = ~controllable_DEQ & ~n13925;
  assign n13927 = ~n13920 & ~n13926;
  assign n13928 = i_FULL & ~n13927;
  assign n13929 = ~n7977 & ~n10910;
  assign n13930 = ~controllable_BtoR_REQ0 & ~n13929;
  assign n13931 = ~controllable_BtoR_REQ0 & ~n13930;
  assign n13932 = ~i_RtoB_ACK0 & ~n13931;
  assign n13933 = ~n8468 & ~n13932;
  assign n13934 = controllable_DEQ & ~n13933;
  assign n13935 = ~n7986 & ~n10520;
  assign n13936 = ~controllable_BtoR_REQ0 & ~n13935;
  assign n13937 = ~controllable_BtoR_REQ0 & ~n13936;
  assign n13938 = ~i_RtoB_ACK0 & ~n13937;
  assign n13939 = ~n8486 & ~n13938;
  assign n13940 = ~controllable_DEQ & ~n13939;
  assign n13941 = ~n13934 & ~n13940;
  assign n13942 = ~i_FULL & ~n13941;
  assign n13943 = ~n13928 & ~n13942;
  assign n13944 = i_nEMPTY & ~n13943;
  assign n13945 = ~n8017 & ~n10546;
  assign n13946 = ~controllable_BtoR_REQ0 & ~n13945;
  assign n13947 = ~controllable_BtoR_REQ0 & ~n13946;
  assign n13948 = ~i_RtoB_ACK0 & ~n13947;
  assign n13949 = ~n8468 & ~n13948;
  assign n13950 = ~controllable_DEQ & ~n13949;
  assign n13951 = ~n8516 & ~n13950;
  assign n13952 = i_FULL & ~n13951;
  assign n13953 = ~controllable_DEQ & ~n13919;
  assign n13954 = ~n8526 & ~n13953;
  assign n13955 = ~i_FULL & ~n13954;
  assign n13956 = ~n13952 & ~n13955;
  assign n13957 = ~i_nEMPTY & ~n13956;
  assign n13958 = ~n13944 & ~n13957;
  assign n13959 = controllable_BtoS_ACK0 & ~n13958;
  assign n13960 = ~n8104 & ~n10957;
  assign n13961 = ~controllable_BtoR_REQ0 & ~n13960;
  assign n13962 = ~controllable_BtoR_REQ0 & ~n13961;
  assign n13963 = ~i_RtoB_ACK0 & ~n13962;
  assign n13964 = ~n8547 & ~n13963;
  assign n13965 = controllable_DEQ & ~n13964;
  assign n13966 = ~n8124 & ~n10622;
  assign n13967 = ~controllable_BtoR_REQ0 & ~n13966;
  assign n13968 = ~controllable_BtoR_REQ0 & ~n13967;
  assign n13969 = ~i_RtoB_ACK0 & ~n13968;
  assign n13970 = ~n8565 & ~n13969;
  assign n13971 = ~controllable_DEQ & ~n13970;
  assign n13972 = ~n13965 & ~n13971;
  assign n13973 = i_FULL & ~n13972;
  assign n13974 = ~n8141 & ~n10977;
  assign n13975 = ~controllable_BtoR_REQ0 & ~n13974;
  assign n13976 = ~controllable_BtoR_REQ0 & ~n13975;
  assign n13977 = ~i_RtoB_ACK0 & ~n13976;
  assign n13978 = ~n8547 & ~n13977;
  assign n13979 = controllable_DEQ & ~n13978;
  assign n13980 = ~n8150 & ~n10647;
  assign n13981 = ~controllable_BtoR_REQ0 & ~n13980;
  assign n13982 = ~controllable_BtoR_REQ0 & ~n13981;
  assign n13983 = ~i_RtoB_ACK0 & ~n13982;
  assign n13984 = ~n8565 & ~n13983;
  assign n13985 = ~controllable_DEQ & ~n13984;
  assign n13986 = ~n13979 & ~n13985;
  assign n13987 = ~i_FULL & ~n13986;
  assign n13988 = ~n13973 & ~n13987;
  assign n13989 = i_nEMPTY & ~n13988;
  assign n13990 = ~n8181 & ~n10673;
  assign n13991 = ~controllable_BtoR_REQ0 & ~n13990;
  assign n13992 = ~controllable_BtoR_REQ0 & ~n13991;
  assign n13993 = ~i_RtoB_ACK0 & ~n13992;
  assign n13994 = ~n8547 & ~n13993;
  assign n13995 = ~controllable_DEQ & ~n13994;
  assign n13996 = ~n8595 & ~n13995;
  assign n13997 = i_FULL & ~n13996;
  assign n13998 = ~controllable_DEQ & ~n13964;
  assign n13999 = ~n8605 & ~n13998;
  assign n14000 = ~i_FULL & ~n13999;
  assign n14001 = ~n13997 & ~n14000;
  assign n14002 = ~i_nEMPTY & ~n14001;
  assign n14003 = ~n13989 & ~n14002;
  assign n14004 = ~controllable_BtoS_ACK0 & ~n14003;
  assign n14005 = ~n13959 & ~n14004;
  assign n14006 = n4465 & ~n14005;
  assign n14007 = ~n8242 & ~n11022;
  assign n14008 = ~controllable_BtoR_REQ0 & ~n14007;
  assign n14009 = ~controllable_BtoR_REQ0 & ~n14008;
  assign n14010 = ~i_RtoB_ACK0 & ~n14009;
  assign n14011 = ~n8621 & ~n14010;
  assign n14012 = controllable_DEQ & ~n14011;
  assign n14013 = ~n8637 & ~n13834;
  assign n14014 = ~controllable_DEQ & ~n14013;
  assign n14015 = ~n14012 & ~n14014;
  assign n14016 = i_nEMPTY & ~n14015;
  assign n14017 = ~n8621 & ~n13842;
  assign n14018 = ~controllable_DEQ & ~n14017;
  assign n14019 = ~n8649 & ~n14018;
  assign n14020 = i_FULL & ~n14019;
  assign n14021 = ~controllable_DEQ & ~n14011;
  assign n14022 = ~n8659 & ~n14021;
  assign n14023 = ~i_FULL & ~n14022;
  assign n14024 = ~n14020 & ~n14023;
  assign n14025 = ~i_nEMPTY & ~n14024;
  assign n14026 = ~n14016 & ~n14025;
  assign n14027 = controllable_BtoS_ACK0 & ~n14026;
  assign n14028 = ~n8345 & ~n11067;
  assign n14029 = ~controllable_BtoR_REQ0 & ~n14028;
  assign n14030 = ~controllable_BtoR_REQ0 & ~n14029;
  assign n14031 = ~i_RtoB_ACK0 & ~n14030;
  assign n14032 = ~n8679 & ~n14031;
  assign n14033 = controllable_DEQ & ~n14032;
  assign n14034 = ~n8697 & ~n13868;
  assign n14035 = ~controllable_DEQ & ~n14034;
  assign n14036 = ~n14033 & ~n14035;
  assign n14037 = i_FULL & ~n14036;
  assign n14038 = ~n8380 & ~n11083;
  assign n14039 = ~controllable_BtoR_REQ0 & ~n14038;
  assign n14040 = ~controllable_BtoR_REQ0 & ~n14039;
  assign n14041 = ~i_RtoB_ACK0 & ~n14040;
  assign n14042 = ~n8679 & ~n14041;
  assign n14043 = controllable_DEQ & ~n14042;
  assign n14044 = ~n8697 & ~n13882;
  assign n14045 = ~controllable_DEQ & ~n14044;
  assign n14046 = ~n14043 & ~n14045;
  assign n14047 = ~i_FULL & ~n14046;
  assign n14048 = ~n14037 & ~n14047;
  assign n14049 = i_nEMPTY & ~n14048;
  assign n14050 = ~n8679 & ~n13892;
  assign n14051 = ~controllable_DEQ & ~n14050;
  assign n14052 = ~n8727 & ~n14051;
  assign n14053 = i_FULL & ~n14052;
  assign n14054 = ~controllable_DEQ & ~n14032;
  assign n14055 = ~n8737 & ~n14054;
  assign n14056 = ~i_FULL & ~n14055;
  assign n14057 = ~n14053 & ~n14056;
  assign n14058 = ~i_nEMPTY & ~n14057;
  assign n14059 = ~n14049 & ~n14058;
  assign n14060 = ~controllable_BtoS_ACK0 & ~n14059;
  assign n14061 = ~n14027 & ~n14060;
  assign n14062 = ~n4465 & ~n14061;
  assign n14063 = ~n14006 & ~n14062;
  assign n14064 = i_StoB_REQ10 & ~n14063;
  assign n14065 = ~n13912 & ~n14064;
  assign n14066 = ~controllable_BtoS_ACK10 & ~n14065;
  assign n14067 = ~n13914 & ~n14066;
  assign n14068 = ~n4464 & ~n14067;
  assign n14069 = ~n13634 & ~n14068;
  assign n14070 = n4463 & ~n14069;
  assign n14071 = ~n11128 & ~n14070;
  assign n14072 = n4462 & ~n14071;
  assign n14073 = i_RtoB_ACK1 & ~n12163;
  assign n14074 = ~n11153 & ~n14073;
  assign n14075 = controllable_BtoR_REQ1 & ~n14074;
  assign n14076 = ~n11158 & ~n14075;
  assign n14077 = ~controllable_BtoR_REQ0 & ~n14076;
  assign n14078 = ~controllable_BtoR_REQ0 & ~n14077;
  assign n14079 = ~i_RtoB_ACK0 & ~n14078;
  assign n14080 = ~n11149 & ~n14079;
  assign n14081 = controllable_DEQ & ~n14080;
  assign n14082 = i_RtoB_ACK1 & ~n12161;
  assign n14083 = ~n11156 & ~n14082;
  assign n14084 = controllable_BtoR_REQ1 & ~n14083;
  assign n14085 = ~n11168 & ~n14084;
  assign n14086 = ~controllable_BtoR_REQ0 & ~n14085;
  assign n14087 = ~controllable_BtoR_REQ0 & ~n14086;
  assign n14088 = ~i_RtoB_ACK0 & ~n14087;
  assign n14089 = ~n11172 & ~n14088;
  assign n14090 = ~controllable_DEQ & ~n14089;
  assign n14091 = ~n14081 & ~n14090;
  assign n14092 = i_nEMPTY & ~n14091;
  assign n14093 = ~n12214 & ~n14073;
  assign n14094 = controllable_BtoR_REQ1 & ~n14093;
  assign n14095 = ~n11145 & ~n14094;
  assign n14096 = ~controllable_BtoR_REQ0 & ~n14095;
  assign n14097 = ~controllable_BtoR_REQ0 & ~n14096;
  assign n14098 = ~i_RtoB_ACK0 & ~n14097;
  assign n14099 = ~n11149 & ~n14098;
  assign n14100 = ~controllable_DEQ & ~n14099;
  assign n14101 = ~n11194 & ~n14100;
  assign n14102 = i_FULL & ~n14101;
  assign n14103 = ~controllable_BtoR_REQ1 & ~n11154;
  assign n14104 = ~n14075 & ~n14103;
  assign n14105 = ~controllable_BtoR_REQ0 & ~n14104;
  assign n14106 = ~controllable_BtoR_REQ0 & ~n14105;
  assign n14107 = ~i_RtoB_ACK0 & ~n14106;
  assign n14108 = ~n11149 & ~n14107;
  assign n14109 = ~controllable_DEQ & ~n14108;
  assign n14110 = ~n11209 & ~n14109;
  assign n14111 = ~i_FULL & ~n14110;
  assign n14112 = ~n14102 & ~n14111;
  assign n14113 = ~i_nEMPTY & ~n14112;
  assign n14114 = ~n14092 & ~n14113;
  assign n14115 = controllable_BtoS_ACK0 & ~n14114;
  assign n14116 = i_RtoB_ACK1 & ~n12256;
  assign n14117 = ~n5346 & ~n14116;
  assign n14118 = controllable_BtoR_REQ1 & ~n14117;
  assign n14119 = ~n5351 & ~n14118;
  assign n14120 = ~controllable_BtoR_REQ0 & ~n14119;
  assign n14121 = ~controllable_BtoR_REQ0 & ~n14120;
  assign n14122 = ~i_RtoB_ACK0 & ~n14121;
  assign n14123 = ~n5342 & ~n14122;
  assign n14124 = controllable_DEQ & ~n14123;
  assign n14125 = i_RtoB_ACK1 & ~n12254;
  assign n14126 = ~n5349 & ~n14125;
  assign n14127 = controllable_BtoR_REQ1 & ~n14126;
  assign n14128 = ~n5361 & ~n14127;
  assign n14129 = ~controllable_BtoR_REQ0 & ~n14128;
  assign n14130 = ~controllable_BtoR_REQ0 & ~n14129;
  assign n14131 = ~i_RtoB_ACK0 & ~n14130;
  assign n14132 = ~n5365 & ~n14131;
  assign n14133 = ~controllable_DEQ & ~n14132;
  assign n14134 = ~n14124 & ~n14133;
  assign n14135 = i_nEMPTY & ~n14134;
  assign n14136 = ~n9026 & ~n14116;
  assign n14137 = controllable_BtoR_REQ1 & ~n14136;
  assign n14138 = ~n5338 & ~n14137;
  assign n14139 = ~controllable_BtoR_REQ0 & ~n14138;
  assign n14140 = ~controllable_BtoR_REQ0 & ~n14139;
  assign n14141 = ~i_RtoB_ACK0 & ~n14140;
  assign n14142 = ~n5342 & ~n14141;
  assign n14143 = ~controllable_DEQ & ~n14142;
  assign n14144 = ~n5387 & ~n14143;
  assign n14145 = i_FULL & ~n14144;
  assign n14146 = ~n13226 & ~n14118;
  assign n14147 = ~controllable_BtoR_REQ0 & ~n14146;
  assign n14148 = ~controllable_BtoR_REQ0 & ~n14147;
  assign n14149 = ~i_RtoB_ACK0 & ~n14148;
  assign n14150 = ~n5342 & ~n14149;
  assign n14151 = ~controllable_DEQ & ~n14150;
  assign n14152 = ~n5402 & ~n14151;
  assign n14153 = ~i_FULL & ~n14152;
  assign n14154 = ~n14145 & ~n14153;
  assign n14155 = ~i_nEMPTY & ~n14154;
  assign n14156 = ~n14135 & ~n14155;
  assign n14157 = ~controllable_BtoS_ACK0 & ~n14156;
  assign n14158 = ~n14115 & ~n14157;
  assign n14159 = n4465 & ~n14158;
  assign n14160 = ~n13240 & ~n14159;
  assign n14161 = i_StoB_REQ10 & ~n14160;
  assign n14162 = ~n11380 & ~n14161;
  assign n14163 = controllable_BtoS_ACK10 & ~n14162;
  assign n14164 = ~n11412 & ~n12363;
  assign n14165 = ~controllable_BtoR_REQ0 & ~n14164;
  assign n14166 = ~controllable_BtoR_REQ0 & ~n14165;
  assign n14167 = ~i_RtoB_ACK0 & ~n14166;
  assign n14168 = ~n11397 & ~n14167;
  assign n14169 = controllable_DEQ & ~n14168;
  assign n14170 = ~n11431 & ~n12386;
  assign n14171 = ~controllable_BtoR_REQ0 & ~n14170;
  assign n14172 = ~controllable_BtoR_REQ0 & ~n14171;
  assign n14173 = ~i_RtoB_ACK0 & ~n14172;
  assign n14174 = ~n11426 & ~n14173;
  assign n14175 = ~controllable_DEQ & ~n14174;
  assign n14176 = ~n14169 & ~n14175;
  assign n14177 = i_FULL & ~n14176;
  assign n14178 = ~n11445 & ~n12399;
  assign n14179 = ~controllable_BtoR_REQ0 & ~n14178;
  assign n14180 = ~controllable_BtoR_REQ0 & ~n14179;
  assign n14181 = ~i_RtoB_ACK0 & ~n14180;
  assign n14182 = ~n11397 & ~n14181;
  assign n14183 = controllable_DEQ & ~n14182;
  assign n14184 = ~n11454 & ~n12409;
  assign n14185 = ~controllable_BtoR_REQ0 & ~n14184;
  assign n14186 = ~controllable_BtoR_REQ0 & ~n14185;
  assign n14187 = ~i_RtoB_ACK0 & ~n14186;
  assign n14188 = ~n11426 & ~n14187;
  assign n14189 = ~controllable_DEQ & ~n14188;
  assign n14190 = ~n14183 & ~n14189;
  assign n14191 = ~i_FULL & ~n14190;
  assign n14192 = ~n14177 & ~n14191;
  assign n14193 = i_nEMPTY & ~n14192;
  assign n14194 = ~n11481 & ~n12429;
  assign n14195 = ~controllable_BtoR_REQ0 & ~n14194;
  assign n14196 = ~controllable_BtoR_REQ0 & ~n14195;
  assign n14197 = ~i_RtoB_ACK0 & ~n14196;
  assign n14198 = ~n11397 & ~n14197;
  assign n14199 = ~controllable_DEQ & ~n14198;
  assign n14200 = ~n11476 & ~n14199;
  assign n14201 = i_FULL & ~n14200;
  assign n14202 = ~controllable_DEQ & ~n14168;
  assign n14203 = ~n11497 & ~n14202;
  assign n14204 = ~i_FULL & ~n14203;
  assign n14205 = ~n14201 & ~n14204;
  assign n14206 = ~i_nEMPTY & ~n14205;
  assign n14207 = ~n14193 & ~n14206;
  assign n14208 = controllable_BtoS_ACK0 & ~n14207;
  assign n14209 = ~n11529 & ~n12464;
  assign n14210 = ~controllable_BtoR_REQ0 & ~n14209;
  assign n14211 = ~controllable_BtoR_REQ0 & ~n14210;
  assign n14212 = ~i_RtoB_ACK0 & ~n14211;
  assign n14213 = ~n11519 & ~n14212;
  assign n14214 = controllable_DEQ & ~n14213;
  assign n14215 = ~n9912 & ~n11546;
  assign n14216 = ~controllable_BtoR_REQ0 & ~n14215;
  assign n14217 = ~controllable_BtoR_REQ0 & ~n14216;
  assign n14218 = ~i_RtoB_ACK0 & ~n14217;
  assign n14219 = ~n11543 & ~n14218;
  assign n14220 = ~controllable_DEQ & ~n14219;
  assign n14221 = ~n14214 & ~n14220;
  assign n14222 = i_FULL & ~n14221;
  assign n14223 = ~n11560 & ~n12490;
  assign n14224 = ~controllable_BtoR_REQ0 & ~n14223;
  assign n14225 = ~controllable_BtoR_REQ0 & ~n14224;
  assign n14226 = ~i_RtoB_ACK0 & ~n14225;
  assign n14227 = ~n11519 & ~n14226;
  assign n14228 = controllable_DEQ & ~n14227;
  assign n14229 = ~n11569 & ~n12500;
  assign n14230 = ~controllable_BtoR_REQ0 & ~n14229;
  assign n14231 = ~controllable_BtoR_REQ0 & ~n14230;
  assign n14232 = ~i_RtoB_ACK0 & ~n14231;
  assign n14233 = ~n11543 & ~n14232;
  assign n14234 = ~controllable_DEQ & ~n14233;
  assign n14235 = ~n14228 & ~n14234;
  assign n14236 = ~i_FULL & ~n14235;
  assign n14237 = ~n14222 & ~n14236;
  assign n14238 = i_nEMPTY & ~n14237;
  assign n14239 = ~n9959 & ~n11594;
  assign n14240 = ~controllable_BtoR_REQ0 & ~n14239;
  assign n14241 = ~controllable_BtoR_REQ0 & ~n14240;
  assign n14242 = ~i_RtoB_ACK0 & ~n14241;
  assign n14243 = ~n11519 & ~n14242;
  assign n14244 = ~controllable_DEQ & ~n14243;
  assign n14245 = ~n11592 & ~n14244;
  assign n14246 = i_FULL & ~n14245;
  assign n14247 = ~controllable_DEQ & ~n14213;
  assign n14248 = ~n11610 & ~n14247;
  assign n14249 = ~i_FULL & ~n14248;
  assign n14250 = ~n14246 & ~n14249;
  assign n14251 = ~i_nEMPTY & ~n14250;
  assign n14252 = ~n14238 & ~n14251;
  assign n14253 = ~controllable_BtoS_ACK0 & ~n14252;
  assign n14254 = ~n14208 & ~n14253;
  assign n14255 = n4465 & ~n14254;
  assign n14256 = ~n13593 & ~n14253;
  assign n14257 = ~n4465 & ~n14256;
  assign n14258 = ~n14255 & ~n14257;
  assign n14259 = i_StoB_REQ10 & ~n14258;
  assign n14260 = ~n11668 & ~n12557;
  assign n14261 = ~controllable_BtoR_REQ0 & ~n14260;
  assign n14262 = ~controllable_BtoR_REQ0 & ~n14261;
  assign n14263 = ~i_RtoB_ACK0 & ~n14262;
  assign n14264 = ~n11654 & ~n14263;
  assign n14265 = controllable_DEQ & ~n14264;
  assign n14266 = ~n11686 & ~n12386;
  assign n14267 = ~controllable_BtoR_REQ0 & ~n14266;
  assign n14268 = ~controllable_BtoR_REQ0 & ~n14267;
  assign n14269 = ~i_RtoB_ACK0 & ~n14268;
  assign n14270 = ~n11683 & ~n14269;
  assign n14271 = ~controllable_DEQ & ~n14270;
  assign n14272 = ~n14265 & ~n14271;
  assign n14273 = i_FULL & ~n14272;
  assign n14274 = ~n11703 & ~n12583;
  assign n14275 = ~controllable_BtoR_REQ0 & ~n14274;
  assign n14276 = ~controllable_BtoR_REQ0 & ~n14275;
  assign n14277 = ~i_RtoB_ACK0 & ~n14276;
  assign n14278 = ~n11654 & ~n14277;
  assign n14279 = controllable_DEQ & ~n14278;
  assign n14280 = ~n11712 & ~n12593;
  assign n14281 = ~controllable_BtoR_REQ0 & ~n14280;
  assign n14282 = ~controllable_BtoR_REQ0 & ~n14281;
  assign n14283 = ~i_RtoB_ACK0 & ~n14282;
  assign n14284 = ~n11683 & ~n14283;
  assign n14285 = ~controllable_DEQ & ~n14284;
  assign n14286 = ~n14279 & ~n14285;
  assign n14287 = ~i_FULL & ~n14286;
  assign n14288 = ~n14273 & ~n14287;
  assign n14289 = i_nEMPTY & ~n14288;
  assign n14290 = ~n11740 & ~n12429;
  assign n14291 = ~controllable_BtoR_REQ0 & ~n14290;
  assign n14292 = ~controllable_BtoR_REQ0 & ~n14291;
  assign n14293 = ~i_RtoB_ACK0 & ~n14292;
  assign n14294 = ~n11654 & ~n14293;
  assign n14295 = ~controllable_DEQ & ~n14294;
  assign n14296 = ~n11738 & ~n14295;
  assign n14297 = i_FULL & ~n14296;
  assign n14298 = ~n11758 & ~n12557;
  assign n14299 = ~controllable_BtoR_REQ0 & ~n14298;
  assign n14300 = ~controllable_BtoR_REQ0 & ~n14299;
  assign n14301 = ~i_RtoB_ACK0 & ~n14300;
  assign n14302 = ~n11654 & ~n14301;
  assign n14303 = ~controllable_DEQ & ~n14302;
  assign n14304 = ~n11756 & ~n14303;
  assign n14305 = ~i_FULL & ~n14304;
  assign n14306 = ~n14297 & ~n14305;
  assign n14307 = ~i_nEMPTY & ~n14306;
  assign n14308 = ~n14289 & ~n14307;
  assign n14309 = controllable_BtoS_ACK0 & ~n14308;
  assign n14310 = ~n11815 & ~n12653;
  assign n14311 = ~controllable_BtoR_REQ0 & ~n14310;
  assign n14312 = ~controllable_BtoR_REQ0 & ~n14311;
  assign n14313 = ~i_RtoB_ACK0 & ~n14312;
  assign n14314 = ~n11801 & ~n14313;
  assign n14315 = controllable_DEQ & ~n14314;
  assign n14316 = ~n9912 & ~n11833;
  assign n14317 = ~controllable_BtoR_REQ0 & ~n14316;
  assign n14318 = ~controllable_BtoR_REQ0 & ~n14317;
  assign n14319 = ~i_RtoB_ACK0 & ~n14318;
  assign n14320 = ~n11830 & ~n14319;
  assign n14321 = ~controllable_DEQ & ~n14320;
  assign n14322 = ~n14315 & ~n14321;
  assign n14323 = i_FULL & ~n14322;
  assign n14324 = ~n11850 & ~n12679;
  assign n14325 = ~controllable_BtoR_REQ0 & ~n14324;
  assign n14326 = ~controllable_BtoR_REQ0 & ~n14325;
  assign n14327 = ~i_RtoB_ACK0 & ~n14326;
  assign n14328 = ~n11801 & ~n14327;
  assign n14329 = controllable_DEQ & ~n14328;
  assign n14330 = ~n11859 & ~n12689;
  assign n14331 = ~controllable_BtoR_REQ0 & ~n14330;
  assign n14332 = ~controllable_BtoR_REQ0 & ~n14331;
  assign n14333 = ~i_RtoB_ACK0 & ~n14332;
  assign n14334 = ~n11830 & ~n14333;
  assign n14335 = ~controllable_DEQ & ~n14334;
  assign n14336 = ~n14329 & ~n14335;
  assign n14337 = ~i_FULL & ~n14336;
  assign n14338 = ~n14323 & ~n14337;
  assign n14339 = i_nEMPTY & ~n14338;
  assign n14340 = ~n9959 & ~n11887;
  assign n14341 = ~controllable_BtoR_REQ0 & ~n14340;
  assign n14342 = ~controllable_BtoR_REQ0 & ~n14341;
  assign n14343 = ~i_RtoB_ACK0 & ~n14342;
  assign n14344 = ~n11801 & ~n14343;
  assign n14345 = ~controllable_DEQ & ~n14344;
  assign n14346 = ~n11885 & ~n14345;
  assign n14347 = i_FULL & ~n14346;
  assign n14348 = ~n11905 & ~n12653;
  assign n14349 = ~controllable_BtoR_REQ0 & ~n14348;
  assign n14350 = ~controllable_BtoR_REQ0 & ~n14349;
  assign n14351 = ~i_RtoB_ACK0 & ~n14350;
  assign n14352 = ~n11801 & ~n14351;
  assign n14353 = ~controllable_DEQ & ~n14352;
  assign n14354 = ~n11903 & ~n14353;
  assign n14355 = ~i_FULL & ~n14354;
  assign n14356 = ~n14347 & ~n14355;
  assign n14357 = ~i_nEMPTY & ~n14356;
  assign n14358 = ~n14339 & ~n14357;
  assign n14359 = ~controllable_BtoS_ACK0 & ~n14358;
  assign n14360 = ~n14309 & ~n14359;
  assign n14361 = n4465 & ~n14360;
  assign n14362 = ~n7104 & ~n9791;
  assign n14363 = ~controllable_BtoR_REQ0 & ~n14362;
  assign n14364 = ~controllable_BtoR_REQ0 & ~n14363;
  assign n14365 = ~i_RtoB_ACK0 & ~n14364;
  assign n14366 = ~n7093 & ~n14365;
  assign n14367 = controllable_DEQ & ~n14366;
  assign n14368 = ~n7119 & ~n13574;
  assign n14369 = ~controllable_DEQ & ~n14368;
  assign n14370 = ~n14367 & ~n14369;
  assign n14371 = i_nEMPTY & ~n14370;
  assign n14372 = ~n7093 & ~n13582;
  assign n14373 = ~controllable_DEQ & ~n14372;
  assign n14374 = ~n7142 & ~n14373;
  assign n14375 = i_FULL & ~n14374;
  assign n14376 = ~n7159 & ~n9791;
  assign n14377 = ~controllable_BtoR_REQ0 & ~n14376;
  assign n14378 = ~controllable_BtoR_REQ0 & ~n14377;
  assign n14379 = ~i_RtoB_ACK0 & ~n14378;
  assign n14380 = ~n7093 & ~n14379;
  assign n14381 = ~controllable_DEQ & ~n14380;
  assign n14382 = ~n7157 & ~n14381;
  assign n14383 = ~i_FULL & ~n14382;
  assign n14384 = ~n14375 & ~n14383;
  assign n14385 = ~i_nEMPTY & ~n14384;
  assign n14386 = ~n14371 & ~n14385;
  assign n14387 = controllable_BtoS_ACK0 & ~n14386;
  assign n14388 = ~n13466 & ~n14387;
  assign n14389 = ~n4465 & ~n14388;
  assign n14390 = ~n14361 & ~n14389;
  assign n14391 = ~i_StoB_REQ10 & ~n14390;
  assign n14392 = ~n14259 & ~n14391;
  assign n14393 = ~controllable_BtoS_ACK10 & ~n14392;
  assign n14394 = ~n14163 & ~n14393;
  assign n14395 = n4464 & ~n14394;
  assign n14396 = ~n11380 & ~n13694;
  assign n14397 = controllable_BtoS_ACK10 & ~n14396;
  assign n14398 = ~n11948 & ~n12865;
  assign n14399 = ~controllable_BtoR_REQ0 & ~n14398;
  assign n14400 = ~controllable_BtoR_REQ0 & ~n14399;
  assign n14401 = ~i_RtoB_ACK0 & ~n14400;
  assign n14402 = ~n11938 & ~n14401;
  assign n14403 = controllable_DEQ & ~n14402;
  assign n14404 = ~n10495 & ~n11965;
  assign n14405 = ~controllable_BtoR_REQ0 & ~n14404;
  assign n14406 = ~controllable_BtoR_REQ0 & ~n14405;
  assign n14407 = ~i_RtoB_ACK0 & ~n14406;
  assign n14408 = ~n11962 & ~n14407;
  assign n14409 = ~controllable_DEQ & ~n14408;
  assign n14410 = ~n14403 & ~n14409;
  assign n14411 = i_FULL & ~n14410;
  assign n14412 = ~n11979 & ~n12891;
  assign n14413 = ~controllable_BtoR_REQ0 & ~n14412;
  assign n14414 = ~controllable_BtoR_REQ0 & ~n14413;
  assign n14415 = ~i_RtoB_ACK0 & ~n14414;
  assign n14416 = ~n11938 & ~n14415;
  assign n14417 = controllable_DEQ & ~n14416;
  assign n14418 = ~n11988 & ~n12901;
  assign n14419 = ~controllable_BtoR_REQ0 & ~n14418;
  assign n14420 = ~controllable_BtoR_REQ0 & ~n14419;
  assign n14421 = ~i_RtoB_ACK0 & ~n14420;
  assign n14422 = ~n11962 & ~n14421;
  assign n14423 = ~controllable_DEQ & ~n14422;
  assign n14424 = ~n14417 & ~n14423;
  assign n14425 = ~i_FULL & ~n14424;
  assign n14426 = ~n14411 & ~n14425;
  assign n14427 = i_nEMPTY & ~n14426;
  assign n14428 = ~n10546 & ~n12012;
  assign n14429 = ~controllable_BtoR_REQ0 & ~n14428;
  assign n14430 = ~controllable_BtoR_REQ0 & ~n14429;
  assign n14431 = ~i_RtoB_ACK0 & ~n14430;
  assign n14432 = ~n11938 & ~n14431;
  assign n14433 = ~controllable_DEQ & ~n14432;
  assign n14434 = ~n12010 & ~n14433;
  assign n14435 = i_FULL & ~n14434;
  assign n14436 = ~controllable_DEQ & ~n14402;
  assign n14437 = ~n12028 & ~n14436;
  assign n14438 = ~i_FULL & ~n14437;
  assign n14439 = ~n14435 & ~n14438;
  assign n14440 = ~i_nEMPTY & ~n14439;
  assign n14441 = ~n14427 & ~n14440;
  assign n14442 = controllable_BtoS_ACK0 & ~n14441;
  assign n14443 = ~n12056 & ~n12950;
  assign n14444 = ~controllable_BtoR_REQ0 & ~n14443;
  assign n14445 = ~controllable_BtoR_REQ0 & ~n14444;
  assign n14446 = ~i_RtoB_ACK0 & ~n14445;
  assign n14447 = ~n12046 & ~n14446;
  assign n14448 = controllable_DEQ & ~n14447;
  assign n14449 = ~n10622 & ~n12073;
  assign n14450 = ~controllable_BtoR_REQ0 & ~n14449;
  assign n14451 = ~controllable_BtoR_REQ0 & ~n14450;
  assign n14452 = ~i_RtoB_ACK0 & ~n14451;
  assign n14453 = ~n12070 & ~n14452;
  assign n14454 = ~controllable_DEQ & ~n14453;
  assign n14455 = ~n14448 & ~n14454;
  assign n14456 = i_FULL & ~n14455;
  assign n14457 = ~n12087 & ~n12976;
  assign n14458 = ~controllable_BtoR_REQ0 & ~n14457;
  assign n14459 = ~controllable_BtoR_REQ0 & ~n14458;
  assign n14460 = ~i_RtoB_ACK0 & ~n14459;
  assign n14461 = ~n12046 & ~n14460;
  assign n14462 = controllable_DEQ & ~n14461;
  assign n14463 = ~n12096 & ~n12986;
  assign n14464 = ~controllable_BtoR_REQ0 & ~n14463;
  assign n14465 = ~controllable_BtoR_REQ0 & ~n14464;
  assign n14466 = ~i_RtoB_ACK0 & ~n14465;
  assign n14467 = ~n12070 & ~n14466;
  assign n14468 = ~controllable_DEQ & ~n14467;
  assign n14469 = ~n14462 & ~n14468;
  assign n14470 = ~i_FULL & ~n14469;
  assign n14471 = ~n14456 & ~n14470;
  assign n14472 = i_nEMPTY & ~n14471;
  assign n14473 = ~n10673 & ~n12120;
  assign n14474 = ~controllable_BtoR_REQ0 & ~n14473;
  assign n14475 = ~controllable_BtoR_REQ0 & ~n14474;
  assign n14476 = ~i_RtoB_ACK0 & ~n14475;
  assign n14477 = ~n12046 & ~n14476;
  assign n14478 = ~controllable_DEQ & ~n14477;
  assign n14479 = ~n12118 & ~n14478;
  assign n14480 = i_FULL & ~n14479;
  assign n14481 = ~controllable_DEQ & ~n14447;
  assign n14482 = ~n12136 & ~n14481;
  assign n14483 = ~i_FULL & ~n14482;
  assign n14484 = ~n14480 & ~n14483;
  assign n14485 = ~i_nEMPTY & ~n14484;
  assign n14486 = ~n14472 & ~n14485;
  assign n14487 = ~controllable_BtoS_ACK0 & ~n14486;
  assign n14488 = ~n14442 & ~n14487;
  assign n14489 = n4465 & ~n14488;
  assign n14490 = ~n14027 & ~n14487;
  assign n14491 = ~n4465 & ~n14490;
  assign n14492 = ~n14489 & ~n14491;
  assign n14493 = i_StoB_REQ10 & ~n14492;
  assign n14494 = ~n7940 & ~n10470;
  assign n14495 = ~controllable_BtoR_REQ0 & ~n14494;
  assign n14496 = ~controllable_BtoR_REQ0 & ~n14495;
  assign n14497 = ~i_RtoB_ACK0 & ~n14496;
  assign n14498 = ~n7921 & ~n14497;
  assign n14499 = controllable_DEQ & ~n14498;
  assign n14500 = ~n7955 & ~n13924;
  assign n14501 = ~controllable_DEQ & ~n14500;
  assign n14502 = ~n14499 & ~n14501;
  assign n14503 = i_FULL & ~n14502;
  assign n14504 = ~n7977 & ~n10508;
  assign n14505 = ~controllable_BtoR_REQ0 & ~n14504;
  assign n14506 = ~controllable_BtoR_REQ0 & ~n14505;
  assign n14507 = ~i_RtoB_ACK0 & ~n14506;
  assign n14508 = ~n7921 & ~n14507;
  assign n14509 = controllable_DEQ & ~n14508;
  assign n14510 = ~n7955 & ~n13938;
  assign n14511 = ~controllable_DEQ & ~n14510;
  assign n14512 = ~n14509 & ~n14511;
  assign n14513 = ~i_FULL & ~n14512;
  assign n14514 = ~n14503 & ~n14513;
  assign n14515 = i_nEMPTY & ~n14514;
  assign n14516 = ~n7921 & ~n13948;
  assign n14517 = ~controllable_DEQ & ~n14516;
  assign n14518 = ~n8012 & ~n14517;
  assign n14519 = i_FULL & ~n14518;
  assign n14520 = ~n8035 & ~n10470;
  assign n14521 = ~controllable_BtoR_REQ0 & ~n14520;
  assign n14522 = ~controllable_BtoR_REQ0 & ~n14521;
  assign n14523 = ~i_RtoB_ACK0 & ~n14522;
  assign n14524 = ~n7921 & ~n14523;
  assign n14525 = ~controllable_DEQ & ~n14524;
  assign n14526 = ~n8033 & ~n14525;
  assign n14527 = ~i_FULL & ~n14526;
  assign n14528 = ~n14519 & ~n14527;
  assign n14529 = ~i_nEMPTY & ~n14528;
  assign n14530 = ~n14515 & ~n14529;
  assign n14531 = controllable_BtoS_ACK0 & ~n14530;
  assign n14532 = ~n8104 & ~n10600;
  assign n14533 = ~controllable_BtoR_REQ0 & ~n14532;
  assign n14534 = ~controllable_BtoR_REQ0 & ~n14533;
  assign n14535 = ~i_RtoB_ACK0 & ~n14534;
  assign n14536 = ~n8088 & ~n14535;
  assign n14537 = controllable_DEQ & ~n14536;
  assign n14538 = ~n8119 & ~n13969;
  assign n14539 = ~controllable_DEQ & ~n14538;
  assign n14540 = ~n14537 & ~n14539;
  assign n14541 = i_FULL & ~n14540;
  assign n14542 = ~n8141 & ~n10635;
  assign n14543 = ~controllable_BtoR_REQ0 & ~n14542;
  assign n14544 = ~controllable_BtoR_REQ0 & ~n14543;
  assign n14545 = ~i_RtoB_ACK0 & ~n14544;
  assign n14546 = ~n8088 & ~n14545;
  assign n14547 = controllable_DEQ & ~n14546;
  assign n14548 = ~n8119 & ~n13983;
  assign n14549 = ~controllable_DEQ & ~n14548;
  assign n14550 = ~n14547 & ~n14549;
  assign n14551 = ~i_FULL & ~n14550;
  assign n14552 = ~n14541 & ~n14551;
  assign n14553 = i_nEMPTY & ~n14552;
  assign n14554 = ~n8088 & ~n13993;
  assign n14555 = ~controllable_DEQ & ~n14554;
  assign n14556 = ~n8176 & ~n14555;
  assign n14557 = i_FULL & ~n14556;
  assign n14558 = ~n8199 & ~n10600;
  assign n14559 = ~controllable_BtoR_REQ0 & ~n14558;
  assign n14560 = ~controllable_BtoR_REQ0 & ~n14559;
  assign n14561 = ~i_RtoB_ACK0 & ~n14560;
  assign n14562 = ~n8088 & ~n14561;
  assign n14563 = ~controllable_DEQ & ~n14562;
  assign n14564 = ~n8197 & ~n14563;
  assign n14565 = ~i_FULL & ~n14564;
  assign n14566 = ~n14557 & ~n14565;
  assign n14567 = ~i_nEMPTY & ~n14566;
  assign n14568 = ~n14553 & ~n14567;
  assign n14569 = ~controllable_BtoS_ACK0 & ~n14568;
  assign n14570 = ~n14531 & ~n14569;
  assign n14571 = n4465 & ~n14570;
  assign n14572 = ~n13910 & ~n14571;
  assign n14573 = ~i_StoB_REQ10 & ~n14572;
  assign n14574 = ~n14493 & ~n14573;
  assign n14575 = ~controllable_BtoS_ACK10 & ~n14574;
  assign n14576 = ~n14397 & ~n14575;
  assign n14577 = ~n4464 & ~n14576;
  assign n14578 = ~n14395 & ~n14577;
  assign n14579 = n4463 & ~n14578;
  assign n14580 = ~n13151 & ~n14579;
  assign n14581 = ~n4462 & ~n14580;
  assign n14582 = ~n14072 & ~n14581;
  assign n14583 = ~n4461 & ~n14582;
  assign n14584 = ~n13155 & ~n14583;
  assign n14585 = ~n4459 & ~n14584;
  assign n14586 = ~i_RtoB_ACK1 & ~n8817;
  assign n14587 = ~controllable_BtoR_REQ1 & ~n14586;
  assign n14588 = ~controllable_BtoR_REQ1 & ~n14587;
  assign n14589 = controllable_BtoR_REQ0 & ~n14588;
  assign n14590 = ~controllable_BtoR_REQ1 & ~n5027;
  assign n14591 = ~controllable_BtoR_REQ0 & ~n14590;
  assign n14592 = ~n14589 & ~n14591;
  assign n14593 = i_RtoB_ACK0 & ~n14592;
  assign n14594 = i_RtoB_ACK1 & ~n5016;
  assign n14595 = ~n5035 & ~n14594;
  assign n14596 = ~controllable_BtoR_REQ1 & ~n14595;
  assign n14597 = ~controllable_BtoR_REQ1 & ~n14596;
  assign n14598 = controllable_BtoR_REQ0 & ~n14597;
  assign n14599 = ~controllable_BtoR_REQ1 & ~n5040;
  assign n14600 = ~controllable_BtoR_REQ0 & ~n14599;
  assign n14601 = ~n14598 & ~n14600;
  assign n14602 = ~i_RtoB_ACK0 & ~n14601;
  assign n14603 = ~n14593 & ~n14602;
  assign n14604 = controllable_DEQ & ~n14603;
  assign n14605 = ~controllable_BtoR_REQ1 & ~n5085;
  assign n14606 = controllable_BtoR_REQ0 & ~n14605;
  assign n14607 = ~controllable_BtoR_REQ1 & ~n5050;
  assign n14608 = ~controllable_BtoR_REQ0 & ~n14607;
  assign n14609 = ~n14606 & ~n14608;
  assign n14610 = i_RtoB_ACK0 & ~n14609;
  assign n14611 = i_RtoB_ACK1 & ~n5014;
  assign n14612 = ~n5038 & ~n14611;
  assign n14613 = ~controllable_BtoR_REQ1 & ~n14612;
  assign n14614 = ~controllable_BtoR_REQ1 & ~n14613;
  assign n14615 = controllable_BtoR_REQ0 & ~n14614;
  assign n14616 = ~n14608 & ~n14615;
  assign n14617 = ~i_RtoB_ACK0 & ~n14616;
  assign n14618 = ~n14610 & ~n14617;
  assign n14619 = ~controllable_DEQ & ~n14618;
  assign n14620 = ~n14604 & ~n14619;
  assign n14621 = i_nEMPTY & ~n14620;
  assign n14622 = ~controllable_BtoR_REQ1 & ~n5064;
  assign n14623 = ~controllable_BtoR_REQ1 & ~n14622;
  assign n14624 = controllable_BtoR_REQ0 & ~n14623;
  assign n14625 = ~controllable_BtoR_REQ1 & ~n5070;
  assign n14626 = ~controllable_BtoR_REQ0 & ~n14625;
  assign n14627 = ~n14624 & ~n14626;
  assign n14628 = ~i_RtoB_ACK0 & ~n14627;
  assign n14629 = ~i_RtoB_ACK0 & ~n14628;
  assign n14630 = controllable_DEQ & ~n14629;
  assign n14631 = ~n8817 & ~n14594;
  assign n14632 = ~controllable_BtoR_REQ1 & ~n14631;
  assign n14633 = ~controllable_BtoR_REQ1 & ~n14632;
  assign n14634 = controllable_BtoR_REQ0 & ~n14633;
  assign n14635 = ~n14591 & ~n14634;
  assign n14636 = ~i_RtoB_ACK0 & ~n14635;
  assign n14637 = ~n14593 & ~n14636;
  assign n14638 = ~controllable_DEQ & ~n14637;
  assign n14639 = ~n14630 & ~n14638;
  assign n14640 = i_FULL & ~n14639;
  assign n14641 = ~controllable_BtoR_REQ1 & ~n5048;
  assign n14642 = ~controllable_BtoR_REQ1 & ~n14641;
  assign n14643 = controllable_BtoR_REQ0 & ~n14642;
  assign n14644 = ~controllable_BtoR_REQ0 & ~n14605;
  assign n14645 = ~n14643 & ~n14644;
  assign n14646 = ~i_RtoB_ACK0 & ~n14645;
  assign n14647 = ~i_RtoB_ACK0 & ~n14646;
  assign n14648 = controllable_DEQ & ~n14647;
  assign n14649 = ~controllable_BtoR_REQ1 & ~n13170;
  assign n14650 = ~controllable_BtoR_REQ0 & ~n14649;
  assign n14651 = ~n14598 & ~n14650;
  assign n14652 = ~i_RtoB_ACK0 & ~n14651;
  assign n14653 = ~n14593 & ~n14652;
  assign n14654 = ~controllable_DEQ & ~n14653;
  assign n14655 = ~n14648 & ~n14654;
  assign n14656 = ~i_FULL & ~n14655;
  assign n14657 = ~n14640 & ~n14656;
  assign n14658 = ~i_nEMPTY & ~n14657;
  assign n14659 = ~n14621 & ~n14658;
  assign n14660 = controllable_BtoS_ACK0 & ~n14659;
  assign n14661 = ~i_RtoB_ACK1 & ~n8924;
  assign n14662 = ~controllable_BtoR_REQ1 & ~n14661;
  assign n14663 = ~controllable_BtoR_REQ1 & ~n14662;
  assign n14664 = controllable_BtoR_REQ0 & ~n14663;
  assign n14665 = ~controllable_BtoR_REQ1 & ~n5124;
  assign n14666 = ~controllable_BtoR_REQ0 & ~n14665;
  assign n14667 = ~n14664 & ~n14666;
  assign n14668 = i_RtoB_ACK0 & ~n14667;
  assign n14669 = i_RtoB_ACK1 & ~n5113;
  assign n14670 = ~n5132 & ~n14669;
  assign n14671 = ~controllable_BtoR_REQ1 & ~n14670;
  assign n14672 = ~controllable_BtoR_REQ1 & ~n14671;
  assign n14673 = controllable_BtoR_REQ0 & ~n14672;
  assign n14674 = ~controllable_BtoR_REQ1 & ~n5137;
  assign n14675 = ~controllable_BtoR_REQ0 & ~n14674;
  assign n14676 = ~n14673 & ~n14675;
  assign n14677 = ~i_RtoB_ACK0 & ~n14676;
  assign n14678 = ~n14668 & ~n14677;
  assign n14679 = controllable_DEQ & ~n14678;
  assign n14680 = ~controllable_BtoR_REQ1 & ~n5182;
  assign n14681 = controllable_BtoR_REQ0 & ~n14680;
  assign n14682 = ~controllable_BtoR_REQ1 & ~n5147;
  assign n14683 = ~controllable_BtoR_REQ0 & ~n14682;
  assign n14684 = ~n14681 & ~n14683;
  assign n14685 = i_RtoB_ACK0 & ~n14684;
  assign n14686 = i_RtoB_ACK1 & ~n5111;
  assign n14687 = ~n5135 & ~n14686;
  assign n14688 = ~controllable_BtoR_REQ1 & ~n14687;
  assign n14689 = ~controllable_BtoR_REQ1 & ~n14688;
  assign n14690 = controllable_BtoR_REQ0 & ~n14689;
  assign n14691 = ~n14683 & ~n14690;
  assign n14692 = ~i_RtoB_ACK0 & ~n14691;
  assign n14693 = ~n14685 & ~n14692;
  assign n14694 = ~controllable_DEQ & ~n14693;
  assign n14695 = ~n14679 & ~n14694;
  assign n14696 = i_nEMPTY & ~n14695;
  assign n14697 = ~controllable_BtoR_REQ1 & ~n5161;
  assign n14698 = ~controllable_BtoR_REQ1 & ~n14697;
  assign n14699 = controllable_BtoR_REQ0 & ~n14698;
  assign n14700 = ~controllable_BtoR_REQ1 & ~n5167;
  assign n14701 = ~controllable_BtoR_REQ0 & ~n14700;
  assign n14702 = ~n14699 & ~n14701;
  assign n14703 = ~i_RtoB_ACK0 & ~n14702;
  assign n14704 = ~i_RtoB_ACK0 & ~n14703;
  assign n14705 = controllable_DEQ & ~n14704;
  assign n14706 = ~n8924 & ~n14669;
  assign n14707 = ~controllable_BtoR_REQ1 & ~n14706;
  assign n14708 = ~controllable_BtoR_REQ1 & ~n14707;
  assign n14709 = controllable_BtoR_REQ0 & ~n14708;
  assign n14710 = ~n14666 & ~n14709;
  assign n14711 = ~i_RtoB_ACK0 & ~n14710;
  assign n14712 = ~n14668 & ~n14711;
  assign n14713 = ~controllable_DEQ & ~n14712;
  assign n14714 = ~n14705 & ~n14713;
  assign n14715 = i_FULL & ~n14714;
  assign n14716 = ~controllable_BtoR_REQ1 & ~n5145;
  assign n14717 = ~controllable_BtoR_REQ1 & ~n14716;
  assign n14718 = controllable_BtoR_REQ0 & ~n14717;
  assign n14719 = ~controllable_BtoR_REQ0 & ~n14680;
  assign n14720 = ~n14718 & ~n14719;
  assign n14721 = ~i_RtoB_ACK0 & ~n14720;
  assign n14722 = ~i_RtoB_ACK0 & ~n14721;
  assign n14723 = controllable_DEQ & ~n14722;
  assign n14724 = ~controllable_BtoR_REQ1 & ~n13197;
  assign n14725 = ~controllable_BtoR_REQ0 & ~n14724;
  assign n14726 = ~n14673 & ~n14725;
  assign n14727 = ~i_RtoB_ACK0 & ~n14726;
  assign n14728 = ~n14668 & ~n14727;
  assign n14729 = ~controllable_DEQ & ~n14728;
  assign n14730 = ~n14723 & ~n14729;
  assign n14731 = ~i_FULL & ~n14730;
  assign n14732 = ~n14715 & ~n14731;
  assign n14733 = ~i_nEMPTY & ~n14732;
  assign n14734 = ~n14696 & ~n14733;
  assign n14735 = ~controllable_BtoS_ACK0 & ~n14734;
  assign n14736 = ~n14660 & ~n14735;
  assign n14737 = n4465 & ~n14736;
  assign n14738 = ~i_RtoB_ACK1 & ~n8755;
  assign n14739 = ~controllable_BtoR_REQ1 & ~n14738;
  assign n14740 = ~controllable_BtoR_REQ1 & ~n14739;
  assign n14741 = controllable_BtoR_REQ0 & ~n14740;
  assign n14742 = ~controllable_BtoR_REQ1 & ~n5232;
  assign n14743 = ~controllable_BtoR_REQ0 & ~n14742;
  assign n14744 = ~n14741 & ~n14743;
  assign n14745 = i_RtoB_ACK0 & ~n14744;
  assign n14746 = ~n5240 & ~n7054;
  assign n14747 = ~controllable_BtoR_REQ1 & ~n14746;
  assign n14748 = ~controllable_BtoR_REQ1 & ~n14747;
  assign n14749 = controllable_BtoR_REQ0 & ~n14748;
  assign n14750 = ~controllable_BtoR_REQ1 & ~n5245;
  assign n14751 = ~controllable_BtoR_REQ0 & ~n14750;
  assign n14752 = ~n14749 & ~n14751;
  assign n14753 = ~i_RtoB_ACK0 & ~n14752;
  assign n14754 = ~n14745 & ~n14753;
  assign n14755 = controllable_DEQ & ~n14754;
  assign n14756 = ~controllable_BtoR_REQ1 & ~n5290;
  assign n14757 = controllable_BtoR_REQ0 & ~n14756;
  assign n14758 = ~controllable_BtoR_REQ1 & ~n5255;
  assign n14759 = ~controllable_BtoR_REQ0 & ~n14758;
  assign n14760 = ~n14757 & ~n14759;
  assign n14761 = i_RtoB_ACK0 & ~n14760;
  assign n14762 = ~n5243 & ~n7111;
  assign n14763 = ~controllable_BtoR_REQ1 & ~n14762;
  assign n14764 = ~controllable_BtoR_REQ1 & ~n14763;
  assign n14765 = controllable_BtoR_REQ0 & ~n14764;
  assign n14766 = ~n14759 & ~n14765;
  assign n14767 = ~i_RtoB_ACK0 & ~n14766;
  assign n14768 = ~n14761 & ~n14767;
  assign n14769 = ~controllable_DEQ & ~n14768;
  assign n14770 = ~n14755 & ~n14769;
  assign n14771 = i_nEMPTY & ~n14770;
  assign n14772 = ~controllable_BtoR_REQ1 & ~n5269;
  assign n14773 = ~controllable_BtoR_REQ1 & ~n14772;
  assign n14774 = controllable_BtoR_REQ0 & ~n14773;
  assign n14775 = ~controllable_BtoR_REQ1 & ~n5275;
  assign n14776 = ~controllable_BtoR_REQ0 & ~n14775;
  assign n14777 = ~n14774 & ~n14776;
  assign n14778 = ~i_RtoB_ACK0 & ~n14777;
  assign n14779 = ~i_RtoB_ACK0 & ~n14778;
  assign n14780 = controllable_DEQ & ~n14779;
  assign n14781 = ~n7054 & ~n8755;
  assign n14782 = ~controllable_BtoR_REQ1 & ~n14781;
  assign n14783 = ~controllable_BtoR_REQ1 & ~n14782;
  assign n14784 = controllable_BtoR_REQ0 & ~n14783;
  assign n14785 = ~n14743 & ~n14784;
  assign n14786 = ~i_RtoB_ACK0 & ~n14785;
  assign n14787 = ~n14745 & ~n14786;
  assign n14788 = ~controllable_DEQ & ~n14787;
  assign n14789 = ~n14780 & ~n14788;
  assign n14790 = i_FULL & ~n14789;
  assign n14791 = ~controllable_BtoR_REQ1 & ~n5253;
  assign n14792 = ~controllable_BtoR_REQ1 & ~n14791;
  assign n14793 = controllable_BtoR_REQ0 & ~n14792;
  assign n14794 = ~controllable_BtoR_REQ0 & ~n14756;
  assign n14795 = ~n14793 & ~n14794;
  assign n14796 = ~i_RtoB_ACK0 & ~n14795;
  assign n14797 = ~i_RtoB_ACK0 & ~n14796;
  assign n14798 = controllable_DEQ & ~n14797;
  assign n14799 = ~controllable_BtoR_REQ1 & ~n5241;
  assign n14800 = ~controllable_BtoR_REQ1 & ~n14799;
  assign n14801 = ~controllable_BtoR_REQ0 & ~n14800;
  assign n14802 = ~n14749 & ~n14801;
  assign n14803 = ~i_RtoB_ACK0 & ~n14802;
  assign n14804 = ~n14745 & ~n14803;
  assign n14805 = ~controllable_DEQ & ~n14804;
  assign n14806 = ~n14798 & ~n14805;
  assign n14807 = ~i_FULL & ~n14806;
  assign n14808 = ~n14790 & ~n14807;
  assign n14809 = ~i_nEMPTY & ~n14808;
  assign n14810 = ~n14771 & ~n14809;
  assign n14811 = controllable_BtoS_ACK0 & ~n14810;
  assign n14812 = ~i_RtoB_ACK1 & ~n9026;
  assign n14813 = ~controllable_BtoR_REQ1 & ~n14812;
  assign n14814 = ~controllable_BtoR_REQ1 & ~n14813;
  assign n14815 = controllable_BtoR_REQ0 & ~n14814;
  assign n14816 = ~controllable_BtoR_REQ1 & ~n5338;
  assign n14817 = ~controllable_BtoR_REQ0 & ~n14816;
  assign n14818 = ~n14815 & ~n14817;
  assign n14819 = i_RtoB_ACK0 & ~n14818;
  assign n14820 = i_RtoB_ACK1 & ~n5327;
  assign n14821 = ~n5346 & ~n14820;
  assign n14822 = ~controllable_BtoR_REQ1 & ~n14821;
  assign n14823 = ~controllable_BtoR_REQ1 & ~n14822;
  assign n14824 = controllable_BtoR_REQ0 & ~n14823;
  assign n14825 = ~controllable_BtoR_REQ1 & ~n5351;
  assign n14826 = ~controllable_BtoR_REQ0 & ~n14825;
  assign n14827 = ~n14824 & ~n14826;
  assign n14828 = ~i_RtoB_ACK0 & ~n14827;
  assign n14829 = ~n14819 & ~n14828;
  assign n14830 = controllable_DEQ & ~n14829;
  assign n14831 = ~controllable_BtoR_REQ1 & ~n5396;
  assign n14832 = controllable_BtoR_REQ0 & ~n14831;
  assign n14833 = ~controllable_BtoR_REQ1 & ~n5361;
  assign n14834 = ~controllable_BtoR_REQ0 & ~n14833;
  assign n14835 = ~n14832 & ~n14834;
  assign n14836 = i_RtoB_ACK0 & ~n14835;
  assign n14837 = i_RtoB_ACK1 & ~n5325;
  assign n14838 = ~n5349 & ~n14837;
  assign n14839 = ~controllable_BtoR_REQ1 & ~n14838;
  assign n14840 = ~controllable_BtoR_REQ1 & ~n14839;
  assign n14841 = controllable_BtoR_REQ0 & ~n14840;
  assign n14842 = ~n14834 & ~n14841;
  assign n14843 = ~i_RtoB_ACK0 & ~n14842;
  assign n14844 = ~n14836 & ~n14843;
  assign n14845 = ~controllable_DEQ & ~n14844;
  assign n14846 = ~n14830 & ~n14845;
  assign n14847 = i_nEMPTY & ~n14846;
  assign n14848 = ~controllable_BtoR_REQ1 & ~n5375;
  assign n14849 = ~controllable_BtoR_REQ1 & ~n14848;
  assign n14850 = controllable_BtoR_REQ0 & ~n14849;
  assign n14851 = ~controllable_BtoR_REQ1 & ~n5381;
  assign n14852 = ~controllable_BtoR_REQ0 & ~n14851;
  assign n14853 = ~n14850 & ~n14852;
  assign n14854 = ~i_RtoB_ACK0 & ~n14853;
  assign n14855 = ~i_RtoB_ACK0 & ~n14854;
  assign n14856 = controllable_DEQ & ~n14855;
  assign n14857 = ~n9026 & ~n14820;
  assign n14858 = ~controllable_BtoR_REQ1 & ~n14857;
  assign n14859 = ~controllable_BtoR_REQ1 & ~n14858;
  assign n14860 = controllable_BtoR_REQ0 & ~n14859;
  assign n14861 = ~n14817 & ~n14860;
  assign n14862 = ~i_RtoB_ACK0 & ~n14861;
  assign n14863 = ~n14819 & ~n14862;
  assign n14864 = ~controllable_DEQ & ~n14863;
  assign n14865 = ~n14856 & ~n14864;
  assign n14866 = i_FULL & ~n14865;
  assign n14867 = ~controllable_BtoR_REQ1 & ~n5359;
  assign n14868 = ~controllable_BtoR_REQ1 & ~n14867;
  assign n14869 = controllable_BtoR_REQ0 & ~n14868;
  assign n14870 = ~controllable_BtoR_REQ0 & ~n14831;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = ~i_RtoB_ACK0 & ~n14871;
  assign n14873 = ~i_RtoB_ACK0 & ~n14872;
  assign n14874 = controllable_DEQ & ~n14873;
  assign n14875 = ~controllable_BtoR_REQ1 & ~n13226;
  assign n14876 = ~controllable_BtoR_REQ0 & ~n14875;
  assign n14877 = ~n14824 & ~n14876;
  assign n14878 = ~i_RtoB_ACK0 & ~n14877;
  assign n14879 = ~n14819 & ~n14878;
  assign n14880 = ~controllable_DEQ & ~n14879;
  assign n14881 = ~n14874 & ~n14880;
  assign n14882 = ~i_FULL & ~n14881;
  assign n14883 = ~n14866 & ~n14882;
  assign n14884 = ~i_nEMPTY & ~n14883;
  assign n14885 = ~n14847 & ~n14884;
  assign n14886 = ~controllable_BtoS_ACK0 & ~n14885;
  assign n14887 = ~n14811 & ~n14886;
  assign n14888 = ~n4465 & ~n14887;
  assign n14889 = ~n14737 & ~n14888;
  assign n14890 = i_StoB_REQ10 & ~n14889;
  assign n14891 = ~i_RtoB_ACK1 & ~n6766;
  assign n14892 = ~n5859 & ~n14891;
  assign n14893 = ~controllable_BtoR_REQ1 & ~n14892;
  assign n14894 = ~controllable_BtoR_REQ1 & ~n14893;
  assign n14895 = controllable_BtoR_REQ0 & ~n14894;
  assign n14896 = ~controllable_BtoR_REQ1 & ~n6581;
  assign n14897 = ~controllable_BtoR_REQ0 & ~n14896;
  assign n14898 = ~n14895 & ~n14897;
  assign n14899 = i_RtoB_ACK0 & ~n14898;
  assign n14900 = i_RtoB_ACK1 & ~n6570;
  assign n14901 = ~n6770 & ~n14900;
  assign n14902 = ~controllable_BtoR_REQ1 & ~n14901;
  assign n14903 = ~controllable_BtoR_REQ1 & ~n14902;
  assign n14904 = controllable_BtoR_REQ0 & ~n14903;
  assign n14905 = ~controllable_BtoR_REQ1 & ~n6778;
  assign n14906 = ~controllable_BtoR_REQ0 & ~n14905;
  assign n14907 = ~n14904 & ~n14906;
  assign n14908 = ~i_RtoB_ACK0 & ~n14907;
  assign n14909 = ~n14899 & ~n14908;
  assign n14910 = controllable_DEQ & ~n14909;
  assign n14911 = ~n6785 & ~n6796;
  assign n14912 = ~controllable_BtoR_REQ1 & ~n14911;
  assign n14913 = ~controllable_BtoR_REQ1 & ~n14912;
  assign n14914 = controllable_BtoR_REQ0 & ~n14913;
  assign n14915 = ~controllable_BtoR_REQ1 & ~n6789;
  assign n14916 = ~controllable_BtoR_REQ0 & ~n14915;
  assign n14917 = ~n14914 & ~n14916;
  assign n14918 = i_RtoB_ACK0 & ~n14917;
  assign n14919 = i_RtoB_ACK1 & ~n6568;
  assign n14920 = ~n6796 & ~n14919;
  assign n14921 = ~controllable_BtoR_REQ1 & ~n14920;
  assign n14922 = ~controllable_BtoR_REQ1 & ~n14921;
  assign n14923 = controllable_BtoR_REQ0 & ~n14922;
  assign n14924 = ~controllable_BtoR_REQ1 & ~n6798;
  assign n14925 = ~controllable_BtoR_REQ0 & ~n14924;
  assign n14926 = ~n14923 & ~n14925;
  assign n14927 = ~i_RtoB_ACK0 & ~n14926;
  assign n14928 = ~n14918 & ~n14927;
  assign n14929 = ~controllable_DEQ & ~n14928;
  assign n14930 = ~n14910 & ~n14929;
  assign n14931 = i_FULL & ~n14930;
  assign n14932 = ~i_RtoB_ACK1 & ~n6807;
  assign n14933 = ~n5859 & ~n14932;
  assign n14934 = ~controllable_BtoR_REQ1 & ~n14933;
  assign n14935 = ~controllable_BtoR_REQ1 & ~n14934;
  assign n14936 = controllable_BtoR_REQ0 & ~n14935;
  assign n14937 = ~n14897 & ~n14936;
  assign n14938 = i_RtoB_ACK0 & ~n14937;
  assign n14939 = ~n6810 & ~n14900;
  assign n14940 = ~controllable_BtoR_REQ1 & ~n14939;
  assign n14941 = ~controllable_BtoR_REQ1 & ~n14940;
  assign n14942 = controllable_BtoR_REQ0 & ~n14941;
  assign n14943 = ~controllable_BtoR_REQ1 & ~n6815;
  assign n14944 = ~controllable_BtoR_REQ0 & ~n14943;
  assign n14945 = ~n14942 & ~n14944;
  assign n14946 = ~i_RtoB_ACK0 & ~n14945;
  assign n14947 = ~n14938 & ~n14946;
  assign n14948 = controllable_DEQ & ~n14947;
  assign n14949 = ~n6776 & ~n6785;
  assign n14950 = ~controllable_BtoR_REQ1 & ~n14949;
  assign n14951 = ~controllable_BtoR_REQ1 & ~n14950;
  assign n14952 = controllable_BtoR_REQ0 & ~n14951;
  assign n14953 = ~n14916 & ~n14952;
  assign n14954 = i_RtoB_ACK0 & ~n14953;
  assign n14955 = ~n6776 & ~n14919;
  assign n14956 = ~controllable_BtoR_REQ1 & ~n14955;
  assign n14957 = ~controllable_BtoR_REQ1 & ~n14956;
  assign n14958 = controllable_BtoR_REQ0 & ~n14957;
  assign n14959 = ~controllable_BtoR_REQ1 & ~n6824;
  assign n14960 = ~controllable_BtoR_REQ0 & ~n14959;
  assign n14961 = ~n14958 & ~n14960;
  assign n14962 = ~i_RtoB_ACK0 & ~n14961;
  assign n14963 = ~n14954 & ~n14962;
  assign n14964 = ~controllable_DEQ & ~n14963;
  assign n14965 = ~n14948 & ~n14964;
  assign n14966 = ~i_FULL & ~n14965;
  assign n14967 = ~n14931 & ~n14966;
  assign n14968 = i_nEMPTY & ~n14967;
  assign n14969 = ~i_RtoB_ACK1 & ~n6835;
  assign n14970 = ~i_RtoB_ACK1 & ~n14969;
  assign n14971 = ~controllable_BtoR_REQ1 & ~n14970;
  assign n14972 = ~controllable_BtoR_REQ1 & ~n14971;
  assign n14973 = controllable_BtoR_REQ0 & ~n14972;
  assign n14974 = controllable_BtoR_REQ0 & ~n14973;
  assign n14975 = i_RtoB_ACK0 & ~n14974;
  assign n14976 = ~i_RtoB_ACK1 & ~n6838;
  assign n14977 = ~controllable_BtoR_REQ1 & ~n14976;
  assign n14978 = ~controllable_BtoR_REQ1 & ~n14977;
  assign n14979 = controllable_BtoR_REQ0 & ~n14978;
  assign n14980 = ~controllable_BtoR_REQ1 & ~n6844;
  assign n14981 = ~controllable_BtoR_REQ0 & ~n14980;
  assign n14982 = ~n14979 & ~n14981;
  assign n14983 = ~i_RtoB_ACK0 & ~n14982;
  assign n14984 = ~n14975 & ~n14983;
  assign n14985 = controllable_DEQ & ~n14984;
  assign n14986 = ~n5859 & ~n6853;
  assign n14987 = ~controllable_BtoR_REQ1 & ~n14986;
  assign n14988 = ~controllable_BtoR_REQ1 & ~n14987;
  assign n14989 = controllable_BtoR_REQ0 & ~n14988;
  assign n14990 = ~n14897 & ~n14989;
  assign n14991 = i_RtoB_ACK0 & ~n14990;
  assign n14992 = ~n6853 & ~n14900;
  assign n14993 = ~controllable_BtoR_REQ1 & ~n14992;
  assign n14994 = ~controllable_BtoR_REQ1 & ~n14993;
  assign n14995 = controllable_BtoR_REQ0 & ~n14994;
  assign n14996 = ~controllable_BtoR_REQ1 & ~n6855;
  assign n14997 = ~controllable_BtoR_REQ0 & ~n14996;
  assign n14998 = ~n14995 & ~n14997;
  assign n14999 = ~i_RtoB_ACK0 & ~n14998;
  assign n15000 = ~n14991 & ~n14999;
  assign n15001 = ~controllable_DEQ & ~n15000;
  assign n15002 = ~n14985 & ~n15001;
  assign n15003 = i_FULL & ~n15002;
  assign n15004 = ~i_RtoB_ACK1 & ~n5856;
  assign n15005 = ~i_RtoB_ACK1 & ~n15004;
  assign n15006 = ~controllable_BtoR_REQ1 & ~n15005;
  assign n15007 = ~controllable_BtoR_REQ1 & ~n15006;
  assign n15008 = controllable_BtoR_REQ0 & ~n15007;
  assign n15009 = controllable_BtoR_REQ0 & ~n15008;
  assign n15010 = i_RtoB_ACK0 & ~n15009;
  assign n15011 = ~i_RtoB_ACK1 & ~n6786;
  assign n15012 = ~controllable_BtoR_REQ1 & ~n15011;
  assign n15013 = ~controllable_BtoR_REQ1 & ~n15012;
  assign n15014 = controllable_BtoR_REQ0 & ~n15013;
  assign n15015 = ~controllable_BtoR_REQ1 & ~n6865;
  assign n15016 = ~controllable_BtoR_REQ0 & ~n15015;
  assign n15017 = ~n15014 & ~n15016;
  assign n15018 = ~i_RtoB_ACK0 & ~n15017;
  assign n15019 = ~n15010 & ~n15018;
  assign n15020 = controllable_DEQ & ~n15019;
  assign n15021 = ~controllable_BtoR_REQ1 & ~n6873;
  assign n15022 = ~controllable_BtoR_REQ0 & ~n15021;
  assign n15023 = ~n14904 & ~n15022;
  assign n15024 = ~i_RtoB_ACK0 & ~n15023;
  assign n15025 = ~n14899 & ~n15024;
  assign n15026 = ~controllable_DEQ & ~n15025;
  assign n15027 = ~n15020 & ~n15026;
  assign n15028 = ~i_FULL & ~n15027;
  assign n15029 = ~n15003 & ~n15028;
  assign n15030 = ~i_nEMPTY & ~n15029;
  assign n15031 = ~n14968 & ~n15030;
  assign n15032 = controllable_BtoS_ACK0 & ~n15031;
  assign n15033 = ~i_RtoB_ACK1 & ~n6932;
  assign n15034 = ~n6897 & ~n15033;
  assign n15035 = ~controllable_BtoR_REQ1 & ~n15034;
  assign n15036 = ~controllable_BtoR_REQ1 & ~n15035;
  assign n15037 = controllable_BtoR_REQ0 & ~n15036;
  assign n15038 = ~controllable_BtoR_REQ1 & ~n6920;
  assign n15039 = ~controllable_BtoR_REQ0 & ~n15038;
  assign n15040 = ~n15037 & ~n15039;
  assign n15041 = i_RtoB_ACK0 & ~n15040;
  assign n15042 = i_RtoB_ACK1 & ~n6909;
  assign n15043 = ~n6936 & ~n15042;
  assign n15044 = ~controllable_BtoR_REQ1 & ~n15043;
  assign n15045 = ~controllable_BtoR_REQ1 & ~n15044;
  assign n15046 = controllable_BtoR_REQ0 & ~n15045;
  assign n15047 = ~controllable_BtoR_REQ1 & ~n6944;
  assign n15048 = ~controllable_BtoR_REQ0 & ~n15047;
  assign n15049 = ~n15046 & ~n15048;
  assign n15050 = ~i_RtoB_ACK0 & ~n15049;
  assign n15051 = ~n15041 & ~n15050;
  assign n15052 = controllable_DEQ & ~n15051;
  assign n15053 = ~n6951 & ~n6962;
  assign n15054 = ~controllable_BtoR_REQ1 & ~n15053;
  assign n15055 = ~controllable_BtoR_REQ1 & ~n15054;
  assign n15056 = controllable_BtoR_REQ0 & ~n15055;
  assign n15057 = ~controllable_BtoR_REQ1 & ~n6955;
  assign n15058 = ~controllable_BtoR_REQ0 & ~n15057;
  assign n15059 = ~n15056 & ~n15058;
  assign n15060 = i_RtoB_ACK0 & ~n15059;
  assign n15061 = i_RtoB_ACK1 & ~n6907;
  assign n15062 = ~n6962 & ~n15061;
  assign n15063 = ~controllable_BtoR_REQ1 & ~n15062;
  assign n15064 = ~controllable_BtoR_REQ1 & ~n15063;
  assign n15065 = controllable_BtoR_REQ0 & ~n15064;
  assign n15066 = ~controllable_BtoR_REQ1 & ~n6964;
  assign n15067 = ~controllable_BtoR_REQ0 & ~n15066;
  assign n15068 = ~n15065 & ~n15067;
  assign n15069 = ~i_RtoB_ACK0 & ~n15068;
  assign n15070 = ~n15060 & ~n15069;
  assign n15071 = ~controllable_DEQ & ~n15070;
  assign n15072 = ~n15052 & ~n15071;
  assign n15073 = i_FULL & ~n15072;
  assign n15074 = ~i_RtoB_ACK1 & ~n6973;
  assign n15075 = ~n6897 & ~n15074;
  assign n15076 = ~controllable_BtoR_REQ1 & ~n15075;
  assign n15077 = ~controllable_BtoR_REQ1 & ~n15076;
  assign n15078 = controllable_BtoR_REQ0 & ~n15077;
  assign n15079 = ~n15039 & ~n15078;
  assign n15080 = i_RtoB_ACK0 & ~n15079;
  assign n15081 = ~n6976 & ~n15042;
  assign n15082 = ~controllable_BtoR_REQ1 & ~n15081;
  assign n15083 = ~controllable_BtoR_REQ1 & ~n15082;
  assign n15084 = controllable_BtoR_REQ0 & ~n15083;
  assign n15085 = ~controllable_BtoR_REQ1 & ~n6981;
  assign n15086 = ~controllable_BtoR_REQ0 & ~n15085;
  assign n15087 = ~n15084 & ~n15086;
  assign n15088 = ~i_RtoB_ACK0 & ~n15087;
  assign n15089 = ~n15080 & ~n15088;
  assign n15090 = controllable_DEQ & ~n15089;
  assign n15091 = ~n6942 & ~n6951;
  assign n15092 = ~controllable_BtoR_REQ1 & ~n15091;
  assign n15093 = ~controllable_BtoR_REQ1 & ~n15092;
  assign n15094 = controllable_BtoR_REQ0 & ~n15093;
  assign n15095 = ~n15058 & ~n15094;
  assign n15096 = i_RtoB_ACK0 & ~n15095;
  assign n15097 = ~n6942 & ~n15061;
  assign n15098 = ~controllable_BtoR_REQ1 & ~n15097;
  assign n15099 = ~controllable_BtoR_REQ1 & ~n15098;
  assign n15100 = controllable_BtoR_REQ0 & ~n15099;
  assign n15101 = ~controllable_BtoR_REQ1 & ~n6990;
  assign n15102 = ~controllable_BtoR_REQ0 & ~n15101;
  assign n15103 = ~n15100 & ~n15102;
  assign n15104 = ~i_RtoB_ACK0 & ~n15103;
  assign n15105 = ~n15096 & ~n15104;
  assign n15106 = ~controllable_DEQ & ~n15105;
  assign n15107 = ~n15090 & ~n15106;
  assign n15108 = ~i_FULL & ~n15107;
  assign n15109 = ~n15073 & ~n15108;
  assign n15110 = i_nEMPTY & ~n15109;
  assign n15111 = ~i_RtoB_ACK1 & ~n7001;
  assign n15112 = ~i_RtoB_ACK1 & ~n15111;
  assign n15113 = ~controllable_BtoR_REQ1 & ~n15112;
  assign n15114 = ~controllable_BtoR_REQ1 & ~n15113;
  assign n15115 = controllable_BtoR_REQ0 & ~n15114;
  assign n15116 = controllable_BtoR_REQ0 & ~n15115;
  assign n15117 = i_RtoB_ACK0 & ~n15116;
  assign n15118 = ~i_RtoB_ACK1 & ~n7004;
  assign n15119 = ~controllable_BtoR_REQ1 & ~n15118;
  assign n15120 = ~controllable_BtoR_REQ1 & ~n15119;
  assign n15121 = controllable_BtoR_REQ0 & ~n15120;
  assign n15122 = ~controllable_BtoR_REQ1 & ~n7010;
  assign n15123 = ~controllable_BtoR_REQ0 & ~n15122;
  assign n15124 = ~n15121 & ~n15123;
  assign n15125 = ~i_RtoB_ACK0 & ~n15124;
  assign n15126 = ~n15117 & ~n15125;
  assign n15127 = controllable_DEQ & ~n15126;
  assign n15128 = ~n6897 & ~n7019;
  assign n15129 = ~controllable_BtoR_REQ1 & ~n15128;
  assign n15130 = ~controllable_BtoR_REQ1 & ~n15129;
  assign n15131 = controllable_BtoR_REQ0 & ~n15130;
  assign n15132 = ~n15039 & ~n15131;
  assign n15133 = i_RtoB_ACK0 & ~n15132;
  assign n15134 = ~n7019 & ~n15042;
  assign n15135 = ~controllable_BtoR_REQ1 & ~n15134;
  assign n15136 = ~controllable_BtoR_REQ1 & ~n15135;
  assign n15137 = controllable_BtoR_REQ0 & ~n15136;
  assign n15138 = ~controllable_BtoR_REQ1 & ~n7021;
  assign n15139 = ~controllable_BtoR_REQ0 & ~n15138;
  assign n15140 = ~n15137 & ~n15139;
  assign n15141 = ~i_RtoB_ACK0 & ~n15140;
  assign n15142 = ~n15133 & ~n15141;
  assign n15143 = ~controllable_DEQ & ~n15142;
  assign n15144 = ~n15127 & ~n15143;
  assign n15145 = i_FULL & ~n15144;
  assign n15146 = ~i_RtoB_ACK1 & ~n6894;
  assign n15147 = ~i_RtoB_ACK1 & ~n15146;
  assign n15148 = ~controllable_BtoR_REQ1 & ~n15147;
  assign n15149 = ~controllable_BtoR_REQ1 & ~n15148;
  assign n15150 = controllable_BtoR_REQ0 & ~n15149;
  assign n15151 = controllable_BtoR_REQ0 & ~n15150;
  assign n15152 = i_RtoB_ACK0 & ~n15151;
  assign n15153 = ~i_RtoB_ACK1 & ~n6952;
  assign n15154 = ~controllable_BtoR_REQ1 & ~n15153;
  assign n15155 = ~controllable_BtoR_REQ1 & ~n15154;
  assign n15156 = controllable_BtoR_REQ0 & ~n15155;
  assign n15157 = ~controllable_BtoR_REQ1 & ~n7031;
  assign n15158 = ~controllable_BtoR_REQ0 & ~n15157;
  assign n15159 = ~n15156 & ~n15158;
  assign n15160 = ~i_RtoB_ACK0 & ~n15159;
  assign n15161 = ~n15152 & ~n15160;
  assign n15162 = controllable_DEQ & ~n15161;
  assign n15163 = ~controllable_BtoR_REQ1 & ~n7039;
  assign n15164 = ~controllable_BtoR_REQ0 & ~n15163;
  assign n15165 = ~n15046 & ~n15164;
  assign n15166 = ~i_RtoB_ACK0 & ~n15165;
  assign n15167 = ~n15041 & ~n15166;
  assign n15168 = ~controllable_DEQ & ~n15167;
  assign n15169 = ~n15162 & ~n15168;
  assign n15170 = ~i_FULL & ~n15169;
  assign n15171 = ~n15145 & ~n15170;
  assign n15172 = ~i_nEMPTY & ~n15171;
  assign n15173 = ~n15110 & ~n15172;
  assign n15174 = ~controllable_BtoS_ACK0 & ~n15173;
  assign n15175 = ~n15032 & ~n15174;
  assign n15176 = n4465 & ~n15175;
  assign n15177 = ~i_RtoB_ACK1 & ~n7094;
  assign n15178 = ~n7054 & ~n15177;
  assign n15179 = ~controllable_BtoR_REQ1 & ~n15178;
  assign n15180 = ~controllable_BtoR_REQ1 & ~n15179;
  assign n15181 = controllable_BtoR_REQ0 & ~n15180;
  assign n15182 = ~controllable_BtoR_REQ1 & ~n7089;
  assign n15183 = ~controllable_BtoR_REQ0 & ~n15182;
  assign n15184 = ~n15181 & ~n15183;
  assign n15185 = i_RtoB_ACK0 & ~n15184;
  assign n15186 = i_RtoB_ACK1 & ~n7078;
  assign n15187 = ~n7098 & ~n15186;
  assign n15188 = ~controllable_BtoR_REQ1 & ~n15187;
  assign n15189 = ~controllable_BtoR_REQ1 & ~n15188;
  assign n15190 = controllable_BtoR_REQ0 & ~n15189;
  assign n15191 = ~controllable_BtoR_REQ1 & ~n7104;
  assign n15192 = ~controllable_BtoR_REQ0 & ~n15191;
  assign n15193 = ~n15190 & ~n15192;
  assign n15194 = ~i_RtoB_ACK0 & ~n15193;
  assign n15195 = ~n15185 & ~n15194;
  assign n15196 = controllable_DEQ & ~n15195;
  assign n15197 = ~n7102 & ~n7111;
  assign n15198 = ~controllable_BtoR_REQ1 & ~n15197;
  assign n15199 = ~controllable_BtoR_REQ1 & ~n15198;
  assign n15200 = controllable_BtoR_REQ0 & ~n15199;
  assign n15201 = ~controllable_BtoR_REQ1 & ~n7115;
  assign n15202 = ~controllable_BtoR_REQ0 & ~n15201;
  assign n15203 = ~n15200 & ~n15202;
  assign n15204 = i_RtoB_ACK0 & ~n15203;
  assign n15205 = i_RtoB_ACK1 & ~n7076;
  assign n15206 = ~n7102 & ~n15205;
  assign n15207 = ~controllable_BtoR_REQ1 & ~n15206;
  assign n15208 = ~controllable_BtoR_REQ1 & ~n15207;
  assign n15209 = controllable_BtoR_REQ0 & ~n15208;
  assign n15210 = ~n15202 & ~n15209;
  assign n15211 = ~i_RtoB_ACK0 & ~n15210;
  assign n15212 = ~n15204 & ~n15211;
  assign n15213 = ~controllable_DEQ & ~n15212;
  assign n15214 = ~n15196 & ~n15213;
  assign n15215 = i_nEMPTY & ~n15214;
  assign n15216 = controllable_BtoR_REQ0 & ~n14774;
  assign n15217 = i_RtoB_ACK0 & ~n15216;
  assign n15218 = ~i_RtoB_ACK1 & ~n7129;
  assign n15219 = ~controllable_BtoR_REQ1 & ~n15218;
  assign n15220 = ~controllable_BtoR_REQ1 & ~n15219;
  assign n15221 = controllable_BtoR_REQ0 & ~n15220;
  assign n15222 = ~controllable_BtoR_REQ1 & ~n7136;
  assign n15223 = ~controllable_BtoR_REQ0 & ~n15222;
  assign n15224 = ~n15221 & ~n15223;
  assign n15225 = ~i_RtoB_ACK0 & ~n15224;
  assign n15226 = ~n15217 & ~n15225;
  assign n15227 = controllable_DEQ & ~n15226;
  assign n15228 = ~n7054 & ~n7546;
  assign n15229 = ~controllable_BtoR_REQ1 & ~n15228;
  assign n15230 = ~controllable_BtoR_REQ1 & ~n15229;
  assign n15231 = controllable_BtoR_REQ0 & ~n15230;
  assign n15232 = ~n15183 & ~n15231;
  assign n15233 = i_RtoB_ACK0 & ~n15232;
  assign n15234 = ~n7546 & ~n15186;
  assign n15235 = ~controllable_BtoR_REQ1 & ~n15234;
  assign n15236 = ~controllable_BtoR_REQ1 & ~n15235;
  assign n15237 = controllable_BtoR_REQ0 & ~n15236;
  assign n15238 = ~n15183 & ~n15237;
  assign n15239 = ~i_RtoB_ACK0 & ~n15238;
  assign n15240 = ~n15233 & ~n15239;
  assign n15241 = ~controllable_DEQ & ~n15240;
  assign n15242 = ~n15227 & ~n15241;
  assign n15243 = i_FULL & ~n15242;
  assign n15244 = controllable_BtoR_REQ0 & ~n14793;
  assign n15245 = i_RtoB_ACK0 & ~n15244;
  assign n15246 = ~i_RtoB_ACK1 & ~n7112;
  assign n15247 = ~controllable_BtoR_REQ1 & ~n15246;
  assign n15248 = ~controllable_BtoR_REQ1 & ~n15247;
  assign n15249 = controllable_BtoR_REQ0 & ~n15248;
  assign n15250 = ~controllable_BtoR_REQ1 & ~n7151;
  assign n15251 = ~controllable_BtoR_REQ0 & ~n15250;
  assign n15252 = ~n15249 & ~n15251;
  assign n15253 = ~i_RtoB_ACK0 & ~n15252;
  assign n15254 = ~n15245 & ~n15253;
  assign n15255 = controllable_DEQ & ~n15254;
  assign n15256 = ~controllable_BtoR_REQ1 & ~n7159;
  assign n15257 = ~controllable_BtoR_REQ0 & ~n15256;
  assign n15258 = ~n15190 & ~n15257;
  assign n15259 = ~i_RtoB_ACK0 & ~n15258;
  assign n15260 = ~n15185 & ~n15259;
  assign n15261 = ~controllable_DEQ & ~n15260;
  assign n15262 = ~n15255 & ~n15261;
  assign n15263 = ~i_FULL & ~n15262;
  assign n15264 = ~n15243 & ~n15263;
  assign n15265 = ~i_nEMPTY & ~n15264;
  assign n15266 = ~n15215 & ~n15265;
  assign n15267 = controllable_BtoS_ACK0 & ~n15266;
  assign n15268 = ~i_RtoB_ACK1 & ~n7258;
  assign n15269 = ~n7196 & ~n15268;
  assign n15270 = ~controllable_BtoR_REQ1 & ~n15269;
  assign n15271 = ~controllable_BtoR_REQ1 & ~n15270;
  assign n15272 = controllable_BtoR_REQ0 & ~n15271;
  assign n15273 = ~controllable_BtoR_REQ1 & ~n7242;
  assign n15274 = ~controllable_BtoR_REQ0 & ~n15273;
  assign n15275 = ~n15272 & ~n15274;
  assign n15276 = i_RtoB_ACK0 & ~n15275;
  assign n15277 = i_RtoB_ACK1 & ~n7231;
  assign n15278 = ~n7262 & ~n15277;
  assign n15279 = ~controllable_BtoR_REQ1 & ~n15278;
  assign n15280 = ~controllable_BtoR_REQ1 & ~n15279;
  assign n15281 = controllable_BtoR_REQ0 & ~n15280;
  assign n15282 = ~controllable_BtoR_REQ1 & ~n7270;
  assign n15283 = ~controllable_BtoR_REQ0 & ~n15282;
  assign n15284 = ~n15281 & ~n15283;
  assign n15285 = ~i_RtoB_ACK0 & ~n15284;
  assign n15286 = ~n15276 & ~n15285;
  assign n15287 = controllable_DEQ & ~n15286;
  assign n15288 = ~n7277 & ~n7288;
  assign n15289 = ~controllable_BtoR_REQ1 & ~n15288;
  assign n15290 = ~controllable_BtoR_REQ1 & ~n15289;
  assign n15291 = controllable_BtoR_REQ0 & ~n15290;
  assign n15292 = ~controllable_BtoR_REQ1 & ~n7281;
  assign n15293 = ~controllable_BtoR_REQ0 & ~n15292;
  assign n15294 = ~n15291 & ~n15293;
  assign n15295 = i_RtoB_ACK0 & ~n15294;
  assign n15296 = i_RtoB_ACK1 & ~n7229;
  assign n15297 = ~n7288 & ~n15296;
  assign n15298 = ~controllable_BtoR_REQ1 & ~n15297;
  assign n15299 = ~controllable_BtoR_REQ1 & ~n15298;
  assign n15300 = controllable_BtoR_REQ0 & ~n15299;
  assign n15301 = ~controllable_BtoR_REQ1 & ~n7290;
  assign n15302 = ~controllable_BtoR_REQ0 & ~n15301;
  assign n15303 = ~n15300 & ~n15302;
  assign n15304 = ~i_RtoB_ACK0 & ~n15303;
  assign n15305 = ~n15295 & ~n15304;
  assign n15306 = ~controllable_DEQ & ~n15305;
  assign n15307 = ~n15287 & ~n15306;
  assign n15308 = i_FULL & ~n15307;
  assign n15309 = ~i_RtoB_ACK1 & ~n7299;
  assign n15310 = ~n7196 & ~n15309;
  assign n15311 = ~controllable_BtoR_REQ1 & ~n15310;
  assign n15312 = ~controllable_BtoR_REQ1 & ~n15311;
  assign n15313 = controllable_BtoR_REQ0 & ~n15312;
  assign n15314 = ~n15274 & ~n15313;
  assign n15315 = i_RtoB_ACK0 & ~n15314;
  assign n15316 = ~n7302 & ~n15277;
  assign n15317 = ~controllable_BtoR_REQ1 & ~n15316;
  assign n15318 = ~controllable_BtoR_REQ1 & ~n15317;
  assign n15319 = controllable_BtoR_REQ0 & ~n15318;
  assign n15320 = ~controllable_BtoR_REQ1 & ~n7307;
  assign n15321 = ~controllable_BtoR_REQ0 & ~n15320;
  assign n15322 = ~n15319 & ~n15321;
  assign n15323 = ~i_RtoB_ACK0 & ~n15322;
  assign n15324 = ~n15315 & ~n15323;
  assign n15325 = controllable_DEQ & ~n15324;
  assign n15326 = ~n7268 & ~n7277;
  assign n15327 = ~controllable_BtoR_REQ1 & ~n15326;
  assign n15328 = ~controllable_BtoR_REQ1 & ~n15327;
  assign n15329 = controllable_BtoR_REQ0 & ~n15328;
  assign n15330 = ~n15293 & ~n15329;
  assign n15331 = i_RtoB_ACK0 & ~n15330;
  assign n15332 = ~n7268 & ~n15296;
  assign n15333 = ~controllable_BtoR_REQ1 & ~n15332;
  assign n15334 = ~controllable_BtoR_REQ1 & ~n15333;
  assign n15335 = controllable_BtoR_REQ0 & ~n15334;
  assign n15336 = ~controllable_BtoR_REQ1 & ~n7316;
  assign n15337 = ~controllable_BtoR_REQ0 & ~n15336;
  assign n15338 = ~n15335 & ~n15337;
  assign n15339 = ~i_RtoB_ACK0 & ~n15338;
  assign n15340 = ~n15331 & ~n15339;
  assign n15341 = ~controllable_DEQ & ~n15340;
  assign n15342 = ~n15325 & ~n15341;
  assign n15343 = ~i_FULL & ~n15342;
  assign n15344 = ~n15308 & ~n15343;
  assign n15345 = i_nEMPTY & ~n15344;
  assign n15346 = ~i_RtoB_ACK1 & ~n7327;
  assign n15347 = ~i_RtoB_ACK1 & ~n15346;
  assign n15348 = ~controllable_BtoR_REQ1 & ~n15347;
  assign n15349 = ~controllable_BtoR_REQ1 & ~n15348;
  assign n15350 = controllable_BtoR_REQ0 & ~n15349;
  assign n15351 = controllable_BtoR_REQ0 & ~n15350;
  assign n15352 = i_RtoB_ACK0 & ~n15351;
  assign n15353 = ~i_RtoB_ACK1 & ~n7330;
  assign n15354 = ~controllable_BtoR_REQ1 & ~n15353;
  assign n15355 = ~controllable_BtoR_REQ1 & ~n15354;
  assign n15356 = controllable_BtoR_REQ0 & ~n15355;
  assign n15357 = ~controllable_BtoR_REQ1 & ~n7336;
  assign n15358 = ~controllable_BtoR_REQ0 & ~n15357;
  assign n15359 = ~n15356 & ~n15358;
  assign n15360 = ~i_RtoB_ACK0 & ~n15359;
  assign n15361 = ~n15352 & ~n15360;
  assign n15362 = controllable_DEQ & ~n15361;
  assign n15363 = ~n7196 & ~n7345;
  assign n15364 = ~controllable_BtoR_REQ1 & ~n15363;
  assign n15365 = ~controllable_BtoR_REQ1 & ~n15364;
  assign n15366 = controllable_BtoR_REQ0 & ~n15365;
  assign n15367 = ~n15274 & ~n15366;
  assign n15368 = i_RtoB_ACK0 & ~n15367;
  assign n15369 = ~n7345 & ~n15277;
  assign n15370 = ~controllable_BtoR_REQ1 & ~n15369;
  assign n15371 = ~controllable_BtoR_REQ1 & ~n15370;
  assign n15372 = controllable_BtoR_REQ0 & ~n15371;
  assign n15373 = ~controllable_BtoR_REQ1 & ~n7347;
  assign n15374 = ~controllable_BtoR_REQ0 & ~n15373;
  assign n15375 = ~n15372 & ~n15374;
  assign n15376 = ~i_RtoB_ACK0 & ~n15375;
  assign n15377 = ~n15368 & ~n15376;
  assign n15378 = ~controllable_DEQ & ~n15377;
  assign n15379 = ~n15362 & ~n15378;
  assign n15380 = i_FULL & ~n15379;
  assign n15381 = ~i_RtoB_ACK1 & ~n7193;
  assign n15382 = ~i_RtoB_ACK1 & ~n15381;
  assign n15383 = ~controllable_BtoR_REQ1 & ~n15382;
  assign n15384 = ~controllable_BtoR_REQ1 & ~n15383;
  assign n15385 = controllable_BtoR_REQ0 & ~n15384;
  assign n15386 = controllable_BtoR_REQ0 & ~n15385;
  assign n15387 = i_RtoB_ACK0 & ~n15386;
  assign n15388 = ~i_RtoB_ACK1 & ~n7278;
  assign n15389 = ~controllable_BtoR_REQ1 & ~n15388;
  assign n15390 = ~controllable_BtoR_REQ1 & ~n15389;
  assign n15391 = controllable_BtoR_REQ0 & ~n15390;
  assign n15392 = ~controllable_BtoR_REQ1 & ~n7357;
  assign n15393 = ~controllable_BtoR_REQ0 & ~n15392;
  assign n15394 = ~n15391 & ~n15393;
  assign n15395 = ~i_RtoB_ACK0 & ~n15394;
  assign n15396 = ~n15387 & ~n15395;
  assign n15397 = controllable_DEQ & ~n15396;
  assign n15398 = ~controllable_BtoR_REQ1 & ~n7365;
  assign n15399 = ~controllable_BtoR_REQ0 & ~n15398;
  assign n15400 = ~n15281 & ~n15399;
  assign n15401 = ~i_RtoB_ACK0 & ~n15400;
  assign n15402 = ~n15276 & ~n15401;
  assign n15403 = ~controllable_DEQ & ~n15402;
  assign n15404 = ~n15397 & ~n15403;
  assign n15405 = ~i_FULL & ~n15404;
  assign n15406 = ~n15380 & ~n15405;
  assign n15407 = ~i_nEMPTY & ~n15406;
  assign n15408 = ~n15345 & ~n15407;
  assign n15409 = ~controllable_BtoS_ACK0 & ~n15408;
  assign n15410 = ~n15267 & ~n15409;
  assign n15411 = ~n4465 & ~n15410;
  assign n15412 = ~n15176 & ~n15411;
  assign n15413 = ~i_StoB_REQ10 & ~n15412;
  assign n15414 = ~n14890 & ~n15413;
  assign n15415 = controllable_BtoS_ACK10 & ~n15414;
  assign n15416 = ~i_RtoB_ACK1 & ~n7400;
  assign n15417 = ~n7391 & ~n15416;
  assign n15418 = ~controllable_BtoR_REQ1 & ~n15417;
  assign n15419 = ~controllable_BtoR_REQ1 & ~n15418;
  assign n15420 = controllable_BtoR_REQ0 & ~n15419;
  assign n15421 = ~n14897 & ~n15420;
  assign n15422 = i_RtoB_ACK0 & ~n15421;
  assign n15423 = ~i_RtoB_ACK0 & ~n14905;
  assign n15424 = ~n15422 & ~n15423;
  assign n15425 = controllable_DEQ & ~n15424;
  assign n15426 = ~n6796 & ~n7410;
  assign n15427 = ~controllable_BtoR_REQ1 & ~n15426;
  assign n15428 = ~controllable_BtoR_REQ1 & ~n15427;
  assign n15429 = controllable_BtoR_REQ0 & ~n15428;
  assign n15430 = ~n14916 & ~n15429;
  assign n15431 = i_RtoB_ACK0 & ~n15430;
  assign n15432 = ~i_RtoB_ACK0 & ~n14924;
  assign n15433 = ~n15431 & ~n15432;
  assign n15434 = ~controllable_DEQ & ~n15433;
  assign n15435 = ~n15425 & ~n15434;
  assign n15436 = i_FULL & ~n15435;
  assign n15437 = ~i_RtoB_ACK1 & ~n7421;
  assign n15438 = ~n7391 & ~n15437;
  assign n15439 = ~controllable_BtoR_REQ1 & ~n15438;
  assign n15440 = ~controllable_BtoR_REQ1 & ~n15439;
  assign n15441 = controllable_BtoR_REQ0 & ~n15440;
  assign n15442 = ~n14897 & ~n15441;
  assign n15443 = i_RtoB_ACK0 & ~n15442;
  assign n15444 = ~i_RtoB_ACK0 & ~n14943;
  assign n15445 = ~n15443 & ~n15444;
  assign n15446 = controllable_DEQ & ~n15445;
  assign n15447 = ~n6776 & ~n7410;
  assign n15448 = ~controllable_BtoR_REQ1 & ~n15447;
  assign n15449 = ~controllable_BtoR_REQ1 & ~n15448;
  assign n15450 = controllable_BtoR_REQ0 & ~n15449;
  assign n15451 = ~n14916 & ~n15450;
  assign n15452 = i_RtoB_ACK0 & ~n15451;
  assign n15453 = ~i_RtoB_ACK0 & ~n14959;
  assign n15454 = ~n15452 & ~n15453;
  assign n15455 = ~controllable_DEQ & ~n15454;
  assign n15456 = ~n15446 & ~n15455;
  assign n15457 = ~i_FULL & ~n15456;
  assign n15458 = ~n15436 & ~n15457;
  assign n15459 = i_nEMPTY & ~n15458;
  assign n15460 = ~i_RtoB_ACK1 & ~n7437;
  assign n15461 = ~i_RtoB_ACK1 & ~n15460;
  assign n15462 = ~controllable_BtoR_REQ1 & ~n15461;
  assign n15463 = ~controllable_BtoR_REQ1 & ~n15462;
  assign n15464 = controllable_BtoR_REQ0 & ~n15463;
  assign n15465 = controllable_BtoR_REQ0 & ~n15464;
  assign n15466 = i_RtoB_ACK0 & ~n15465;
  assign n15467 = ~i_RtoB_ACK0 & ~n14980;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = controllable_DEQ & ~n15468;
  assign n15470 = ~n6853 & ~n7391;
  assign n15471 = ~controllable_BtoR_REQ1 & ~n15470;
  assign n15472 = ~controllable_BtoR_REQ1 & ~n15471;
  assign n15473 = controllable_BtoR_REQ0 & ~n15472;
  assign n15474 = ~n14897 & ~n15473;
  assign n15475 = i_RtoB_ACK0 & ~n15474;
  assign n15476 = ~i_RtoB_ACK0 & ~n14996;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = ~controllable_DEQ & ~n15477;
  assign n15479 = ~n15469 & ~n15478;
  assign n15480 = i_FULL & ~n15479;
  assign n15481 = ~i_RtoB_ACK1 & ~n7388;
  assign n15482 = ~i_RtoB_ACK1 & ~n15481;
  assign n15483 = ~controllable_BtoR_REQ1 & ~n15482;
  assign n15484 = ~controllable_BtoR_REQ1 & ~n15483;
  assign n15485 = controllable_BtoR_REQ0 & ~n15484;
  assign n15486 = controllable_BtoR_REQ0 & ~n15485;
  assign n15487 = i_RtoB_ACK0 & ~n15486;
  assign n15488 = ~i_RtoB_ACK0 & ~n15015;
  assign n15489 = ~n15487 & ~n15488;
  assign n15490 = controllable_DEQ & ~n15489;
  assign n15491 = ~controllable_DEQ & ~n15424;
  assign n15492 = ~n15490 & ~n15491;
  assign n15493 = ~i_FULL & ~n15492;
  assign n15494 = ~n15480 & ~n15493;
  assign n15495 = ~i_nEMPTY & ~n15494;
  assign n15496 = ~n15459 & ~n15495;
  assign n15497 = controllable_BtoS_ACK0 & ~n15496;
  assign n15498 = ~i_RtoB_ACK1 & ~n7480;
  assign n15499 = ~n7471 & ~n15498;
  assign n15500 = ~controllable_BtoR_REQ1 & ~n15499;
  assign n15501 = ~controllable_BtoR_REQ1 & ~n15500;
  assign n15502 = controllable_BtoR_REQ0 & ~n15501;
  assign n15503 = ~n15039 & ~n15502;
  assign n15504 = i_RtoB_ACK0 & ~n15503;
  assign n15505 = ~i_RtoB_ACK0 & ~n15047;
  assign n15506 = ~n15504 & ~n15505;
  assign n15507 = controllable_DEQ & ~n15506;
  assign n15508 = ~n6962 & ~n7490;
  assign n15509 = ~controllable_BtoR_REQ1 & ~n15508;
  assign n15510 = ~controllable_BtoR_REQ1 & ~n15509;
  assign n15511 = controllable_BtoR_REQ0 & ~n15510;
  assign n15512 = ~n15058 & ~n15511;
  assign n15513 = i_RtoB_ACK0 & ~n15512;
  assign n15514 = ~i_RtoB_ACK0 & ~n15066;
  assign n15515 = ~n15513 & ~n15514;
  assign n15516 = ~controllable_DEQ & ~n15515;
  assign n15517 = ~n15507 & ~n15516;
  assign n15518 = i_FULL & ~n15517;
  assign n15519 = ~i_RtoB_ACK1 & ~n7501;
  assign n15520 = ~n7471 & ~n15519;
  assign n15521 = ~controllable_BtoR_REQ1 & ~n15520;
  assign n15522 = ~controllable_BtoR_REQ1 & ~n15521;
  assign n15523 = controllable_BtoR_REQ0 & ~n15522;
  assign n15524 = ~n15039 & ~n15523;
  assign n15525 = i_RtoB_ACK0 & ~n15524;
  assign n15526 = ~i_RtoB_ACK0 & ~n15085;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = controllable_DEQ & ~n15527;
  assign n15529 = ~n6942 & ~n7490;
  assign n15530 = ~controllable_BtoR_REQ1 & ~n15529;
  assign n15531 = ~controllable_BtoR_REQ1 & ~n15530;
  assign n15532 = controllable_BtoR_REQ0 & ~n15531;
  assign n15533 = ~n15058 & ~n15532;
  assign n15534 = i_RtoB_ACK0 & ~n15533;
  assign n15535 = ~i_RtoB_ACK0 & ~n15101;
  assign n15536 = ~n15534 & ~n15535;
  assign n15537 = ~controllable_DEQ & ~n15536;
  assign n15538 = ~n15528 & ~n15537;
  assign n15539 = ~i_FULL & ~n15538;
  assign n15540 = ~n15518 & ~n15539;
  assign n15541 = i_nEMPTY & ~n15540;
  assign n15542 = ~i_RtoB_ACK1 & ~n7517;
  assign n15543 = ~i_RtoB_ACK1 & ~n15542;
  assign n15544 = ~controllable_BtoR_REQ1 & ~n15543;
  assign n15545 = ~controllable_BtoR_REQ1 & ~n15544;
  assign n15546 = controllable_BtoR_REQ0 & ~n15545;
  assign n15547 = controllable_BtoR_REQ0 & ~n15546;
  assign n15548 = i_RtoB_ACK0 & ~n15547;
  assign n15549 = ~i_RtoB_ACK0 & ~n15122;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = controllable_DEQ & ~n15550;
  assign n15552 = ~n7019 & ~n7471;
  assign n15553 = ~controllable_BtoR_REQ1 & ~n15552;
  assign n15554 = ~controllable_BtoR_REQ1 & ~n15553;
  assign n15555 = controllable_BtoR_REQ0 & ~n15554;
  assign n15556 = ~n15039 & ~n15555;
  assign n15557 = i_RtoB_ACK0 & ~n15556;
  assign n15558 = ~i_RtoB_ACK0 & ~n15138;
  assign n15559 = ~n15557 & ~n15558;
  assign n15560 = ~controllable_DEQ & ~n15559;
  assign n15561 = ~n15551 & ~n15560;
  assign n15562 = i_FULL & ~n15561;
  assign n15563 = ~i_RtoB_ACK1 & ~n7468;
  assign n15564 = ~i_RtoB_ACK1 & ~n15563;
  assign n15565 = ~controllable_BtoR_REQ1 & ~n15564;
  assign n15566 = ~controllable_BtoR_REQ1 & ~n15565;
  assign n15567 = controllable_BtoR_REQ0 & ~n15566;
  assign n15568 = controllable_BtoR_REQ0 & ~n15567;
  assign n15569 = i_RtoB_ACK0 & ~n15568;
  assign n15570 = ~i_RtoB_ACK0 & ~n15157;
  assign n15571 = ~n15569 & ~n15570;
  assign n15572 = controllable_DEQ & ~n15571;
  assign n15573 = ~controllable_DEQ & ~n15506;
  assign n15574 = ~n15572 & ~n15573;
  assign n15575 = ~i_FULL & ~n15574;
  assign n15576 = ~n15562 & ~n15575;
  assign n15577 = ~i_nEMPTY & ~n15576;
  assign n15578 = ~n15541 & ~n15577;
  assign n15579 = ~controllable_BtoS_ACK0 & ~n15578;
  assign n15580 = ~n15497 & ~n15579;
  assign n15581 = n4465 & ~n15580;
  assign n15582 = ~i_RtoB_ACK1 & ~n7553;
  assign n15583 = ~n5237 & ~n15582;
  assign n15584 = ~controllable_BtoR_REQ1 & ~n15583;
  assign n15585 = ~controllable_BtoR_REQ1 & ~n15584;
  assign n15586 = controllable_BtoR_REQ0 & ~n15585;
  assign n15587 = ~n15183 & ~n15586;
  assign n15588 = i_RtoB_ACK0 & ~n15587;
  assign n15589 = ~i_RtoB_ACK0 & ~n15191;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = controllable_DEQ & ~n15590;
  assign n15592 = ~controllable_BtoR_REQ1 & ~n7564;
  assign n15593 = ~controllable_BtoR_REQ1 & ~n15592;
  assign n15594 = controllable_BtoR_REQ0 & ~n15593;
  assign n15595 = ~n15202 & ~n15594;
  assign n15596 = i_RtoB_ACK0 & ~n15595;
  assign n15597 = ~i_RtoB_ACK0 & ~n15201;
  assign n15598 = ~n15596 & ~n15597;
  assign n15599 = ~controllable_DEQ & ~n15598;
  assign n15600 = ~n15591 & ~n15599;
  assign n15601 = i_nEMPTY & ~n15600;
  assign n15602 = controllable_BtoR_REQ0 & ~n14775;
  assign n15603 = controllable_BtoR_REQ0 & ~n15602;
  assign n15604 = i_RtoB_ACK0 & ~n15603;
  assign n15605 = ~i_RtoB_ACK0 & ~n15222;
  assign n15606 = ~n15604 & ~n15605;
  assign n15607 = controllable_DEQ & ~n15606;
  assign n15608 = ~controllable_BtoR_REQ1 & ~n7547;
  assign n15609 = ~controllable_BtoR_REQ1 & ~n15608;
  assign n15610 = controllable_BtoR_REQ0 & ~n15609;
  assign n15611 = ~n15183 & ~n15610;
  assign n15612 = i_RtoB_ACK0 & ~n15611;
  assign n15613 = ~i_RtoB_ACK0 & ~n15182;
  assign n15614 = ~n15612 & ~n15613;
  assign n15615 = ~controllable_DEQ & ~n15614;
  assign n15616 = ~n15607 & ~n15615;
  assign n15617 = i_FULL & ~n15616;
  assign n15618 = controllable_BtoR_REQ0 & ~n14757;
  assign n15619 = i_RtoB_ACK0 & ~n15618;
  assign n15620 = ~i_RtoB_ACK0 & ~n15250;
  assign n15621 = ~n15619 & ~n15620;
  assign n15622 = controllable_DEQ & ~n15621;
  assign n15623 = ~controllable_DEQ & ~n15590;
  assign n15624 = ~n15622 & ~n15623;
  assign n15625 = ~i_FULL & ~n15624;
  assign n15626 = ~n15617 & ~n15625;
  assign n15627 = ~i_nEMPTY & ~n15626;
  assign n15628 = ~n15601 & ~n15627;
  assign n15629 = controllable_BtoS_ACK0 & ~n15628;
  assign n15630 = ~i_RtoB_ACK1 & ~n7616;
  assign n15631 = ~n7607 & ~n15630;
  assign n15632 = ~controllable_BtoR_REQ1 & ~n15631;
  assign n15633 = ~controllable_BtoR_REQ1 & ~n15632;
  assign n15634 = controllable_BtoR_REQ0 & ~n15633;
  assign n15635 = ~n15274 & ~n15634;
  assign n15636 = i_RtoB_ACK0 & ~n15635;
  assign n15637 = ~i_RtoB_ACK0 & ~n15282;
  assign n15638 = ~n15636 & ~n15637;
  assign n15639 = controllable_DEQ & ~n15638;
  assign n15640 = ~n7288 & ~n7626;
  assign n15641 = ~controllable_BtoR_REQ1 & ~n15640;
  assign n15642 = ~controllable_BtoR_REQ1 & ~n15641;
  assign n15643 = controllable_BtoR_REQ0 & ~n15642;
  assign n15644 = ~n15293 & ~n15643;
  assign n15645 = i_RtoB_ACK0 & ~n15644;
  assign n15646 = ~i_RtoB_ACK0 & ~n15301;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = ~controllable_DEQ & ~n15647;
  assign n15649 = ~n15639 & ~n15648;
  assign n15650 = i_FULL & ~n15649;
  assign n15651 = ~i_RtoB_ACK1 & ~n7637;
  assign n15652 = ~n7607 & ~n15651;
  assign n15653 = ~controllable_BtoR_REQ1 & ~n15652;
  assign n15654 = ~controllable_BtoR_REQ1 & ~n15653;
  assign n15655 = controllable_BtoR_REQ0 & ~n15654;
  assign n15656 = ~n15274 & ~n15655;
  assign n15657 = i_RtoB_ACK0 & ~n15656;
  assign n15658 = ~i_RtoB_ACK0 & ~n15320;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = controllable_DEQ & ~n15659;
  assign n15661 = ~n7268 & ~n7626;
  assign n15662 = ~controllable_BtoR_REQ1 & ~n15661;
  assign n15663 = ~controllable_BtoR_REQ1 & ~n15662;
  assign n15664 = controllable_BtoR_REQ0 & ~n15663;
  assign n15665 = ~n15293 & ~n15664;
  assign n15666 = i_RtoB_ACK0 & ~n15665;
  assign n15667 = ~i_RtoB_ACK0 & ~n15336;
  assign n15668 = ~n15666 & ~n15667;
  assign n15669 = ~controllable_DEQ & ~n15668;
  assign n15670 = ~n15660 & ~n15669;
  assign n15671 = ~i_FULL & ~n15670;
  assign n15672 = ~n15650 & ~n15671;
  assign n15673 = i_nEMPTY & ~n15672;
  assign n15674 = ~i_RtoB_ACK1 & ~n7653;
  assign n15675 = ~i_RtoB_ACK1 & ~n15674;
  assign n15676 = ~controllable_BtoR_REQ1 & ~n15675;
  assign n15677 = ~controllable_BtoR_REQ1 & ~n15676;
  assign n15678 = controllable_BtoR_REQ0 & ~n15677;
  assign n15679 = controllable_BtoR_REQ0 & ~n15678;
  assign n15680 = i_RtoB_ACK0 & ~n15679;
  assign n15681 = ~i_RtoB_ACK0 & ~n15357;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = controllable_DEQ & ~n15682;
  assign n15684 = ~n7345 & ~n7607;
  assign n15685 = ~controllable_BtoR_REQ1 & ~n15684;
  assign n15686 = ~controllable_BtoR_REQ1 & ~n15685;
  assign n15687 = controllable_BtoR_REQ0 & ~n15686;
  assign n15688 = ~n15274 & ~n15687;
  assign n15689 = i_RtoB_ACK0 & ~n15688;
  assign n15690 = ~i_RtoB_ACK0 & ~n15373;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = ~controllable_DEQ & ~n15691;
  assign n15693 = ~n15683 & ~n15692;
  assign n15694 = i_FULL & ~n15693;
  assign n15695 = ~i_RtoB_ACK1 & ~n7604;
  assign n15696 = ~i_RtoB_ACK1 & ~n15695;
  assign n15697 = ~controllable_BtoR_REQ1 & ~n15696;
  assign n15698 = ~controllable_BtoR_REQ1 & ~n15697;
  assign n15699 = controllable_BtoR_REQ0 & ~n15698;
  assign n15700 = controllable_BtoR_REQ0 & ~n15699;
  assign n15701 = i_RtoB_ACK0 & ~n15700;
  assign n15702 = ~i_RtoB_ACK0 & ~n15392;
  assign n15703 = ~n15701 & ~n15702;
  assign n15704 = controllable_DEQ & ~n15703;
  assign n15705 = ~controllable_DEQ & ~n15638;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = ~i_FULL & ~n15706;
  assign n15708 = ~n15694 & ~n15707;
  assign n15709 = ~i_nEMPTY & ~n15708;
  assign n15710 = ~n15673 & ~n15709;
  assign n15711 = ~controllable_BtoS_ACK0 & ~n15710;
  assign n15712 = ~n15629 & ~n15711;
  assign n15713 = ~n4465 & ~n15712;
  assign n15714 = ~n15581 & ~n15713;
  assign n15715 = i_StoB_REQ10 & ~n15714;
  assign n15716 = ~n15413 & ~n15715;
  assign n15717 = ~controllable_BtoS_ACK10 & ~n15716;
  assign n15718 = ~n15415 & ~n15717;
  assign n15719 = n4464 & ~n15718;
  assign n15720 = ~i_RtoB_ACK1 & ~n10319;
  assign n15721 = ~controllable_BtoR_REQ1 & ~n15720;
  assign n15722 = ~controllable_BtoR_REQ1 & ~n15721;
  assign n15723 = controllable_BtoR_REQ0 & ~n15722;
  assign n15724 = ~controllable_BtoR_REQ1 & ~n7705;
  assign n15725 = ~controllable_BtoR_REQ0 & ~n15724;
  assign n15726 = ~n15723 & ~n15725;
  assign n15727 = i_RtoB_ACK0 & ~n15726;
  assign n15728 = i_RtoB_ACK1 & ~n7697;
  assign n15729 = ~n7713 & ~n15728;
  assign n15730 = ~controllable_BtoR_REQ1 & ~n15729;
  assign n15731 = ~controllable_BtoR_REQ1 & ~n15730;
  assign n15732 = controllable_BtoR_REQ0 & ~n15731;
  assign n15733 = ~controllable_BtoR_REQ1 & ~n7718;
  assign n15734 = ~controllable_BtoR_REQ0 & ~n15733;
  assign n15735 = ~n15732 & ~n15734;
  assign n15736 = ~i_RtoB_ACK0 & ~n15735;
  assign n15737 = ~n15727 & ~n15736;
  assign n15738 = controllable_DEQ & ~n15737;
  assign n15739 = ~controllable_BtoR_REQ1 & ~n7763;
  assign n15740 = controllable_BtoR_REQ0 & ~n15739;
  assign n15741 = ~controllable_BtoR_REQ1 & ~n7728;
  assign n15742 = ~controllable_BtoR_REQ0 & ~n15741;
  assign n15743 = ~n15740 & ~n15742;
  assign n15744 = i_RtoB_ACK0 & ~n15743;
  assign n15745 = i_RtoB_ACK1 & ~n7695;
  assign n15746 = ~n7716 & ~n15745;
  assign n15747 = ~controllable_BtoR_REQ1 & ~n15746;
  assign n15748 = ~controllable_BtoR_REQ1 & ~n15747;
  assign n15749 = controllable_BtoR_REQ0 & ~n15748;
  assign n15750 = ~n15742 & ~n15749;
  assign n15751 = ~i_RtoB_ACK0 & ~n15750;
  assign n15752 = ~n15744 & ~n15751;
  assign n15753 = ~controllable_DEQ & ~n15752;
  assign n15754 = ~n15738 & ~n15753;
  assign n15755 = i_nEMPTY & ~n15754;
  assign n15756 = ~controllable_BtoR_REQ1 & ~n7742;
  assign n15757 = ~controllable_BtoR_REQ1 & ~n15756;
  assign n15758 = controllable_BtoR_REQ0 & ~n15757;
  assign n15759 = ~controllable_BtoR_REQ1 & ~n7748;
  assign n15760 = ~controllable_BtoR_REQ0 & ~n15759;
  assign n15761 = ~n15758 & ~n15760;
  assign n15762 = ~i_RtoB_ACK0 & ~n15761;
  assign n15763 = ~i_RtoB_ACK0 & ~n15762;
  assign n15764 = controllable_DEQ & ~n15763;
  assign n15765 = ~n10319 & ~n15728;
  assign n15766 = ~controllable_BtoR_REQ1 & ~n15765;
  assign n15767 = ~controllable_BtoR_REQ1 & ~n15766;
  assign n15768 = controllable_BtoR_REQ0 & ~n15767;
  assign n15769 = ~n15725 & ~n15768;
  assign n15770 = ~i_RtoB_ACK0 & ~n15769;
  assign n15771 = ~n15727 & ~n15770;
  assign n15772 = ~controllable_DEQ & ~n15771;
  assign n15773 = ~n15764 & ~n15772;
  assign n15774 = i_FULL & ~n15773;
  assign n15775 = ~controllable_BtoR_REQ1 & ~n7726;
  assign n15776 = ~controllable_BtoR_REQ1 & ~n15775;
  assign n15777 = controllable_BtoR_REQ0 & ~n15776;
  assign n15778 = ~controllable_BtoR_REQ0 & ~n15739;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = ~i_RtoB_ACK0 & ~n15779;
  assign n15781 = ~i_RtoB_ACK0 & ~n15780;
  assign n15782 = controllable_DEQ & ~n15781;
  assign n15783 = ~controllable_BtoR_REQ1 & ~n13649;
  assign n15784 = ~controllable_BtoR_REQ0 & ~n15783;
  assign n15785 = ~n15732 & ~n15784;
  assign n15786 = ~i_RtoB_ACK0 & ~n15785;
  assign n15787 = ~n15727 & ~n15786;
  assign n15788 = ~controllable_DEQ & ~n15787;
  assign n15789 = ~n15782 & ~n15788;
  assign n15790 = ~i_FULL & ~n15789;
  assign n15791 = ~n15774 & ~n15790;
  assign n15792 = ~i_nEMPTY & ~n15791;
  assign n15793 = ~n15755 & ~n15792;
  assign n15794 = controllable_BtoS_ACK0 & ~n15793;
  assign n15795 = ~i_RtoB_ACK1 & ~n10413;
  assign n15796 = ~controllable_BtoR_REQ1 & ~n15795;
  assign n15797 = ~controllable_BtoR_REQ1 & ~n15796;
  assign n15798 = controllable_BtoR_REQ0 & ~n15797;
  assign n15799 = ~controllable_BtoR_REQ1 & ~n7797;
  assign n15800 = ~controllable_BtoR_REQ0 & ~n15799;
  assign n15801 = ~n15798 & ~n15800;
  assign n15802 = i_RtoB_ACK0 & ~n15801;
  assign n15803 = i_RtoB_ACK1 & ~n7787;
  assign n15804 = ~n7805 & ~n15803;
  assign n15805 = ~controllable_BtoR_REQ1 & ~n15804;
  assign n15806 = ~controllable_BtoR_REQ1 & ~n15805;
  assign n15807 = controllable_BtoR_REQ0 & ~n15806;
  assign n15808 = ~controllable_BtoR_REQ1 & ~n7810;
  assign n15809 = ~controllable_BtoR_REQ0 & ~n15808;
  assign n15810 = ~n15807 & ~n15809;
  assign n15811 = ~i_RtoB_ACK0 & ~n15810;
  assign n15812 = ~n15802 & ~n15811;
  assign n15813 = controllable_DEQ & ~n15812;
  assign n15814 = ~controllable_BtoR_REQ1 & ~n7855;
  assign n15815 = controllable_BtoR_REQ0 & ~n15814;
  assign n15816 = ~controllable_BtoR_REQ1 & ~n7820;
  assign n15817 = ~controllable_BtoR_REQ0 & ~n15816;
  assign n15818 = ~n15815 & ~n15817;
  assign n15819 = i_RtoB_ACK0 & ~n15818;
  assign n15820 = i_RtoB_ACK1 & ~n7785;
  assign n15821 = ~n7808 & ~n15820;
  assign n15822 = ~controllable_BtoR_REQ1 & ~n15821;
  assign n15823 = ~controllable_BtoR_REQ1 & ~n15822;
  assign n15824 = controllable_BtoR_REQ0 & ~n15823;
  assign n15825 = ~n15817 & ~n15824;
  assign n15826 = ~i_RtoB_ACK0 & ~n15825;
  assign n15827 = ~n15819 & ~n15826;
  assign n15828 = ~controllable_DEQ & ~n15827;
  assign n15829 = ~n15813 & ~n15828;
  assign n15830 = i_nEMPTY & ~n15829;
  assign n15831 = ~controllable_BtoR_REQ1 & ~n7834;
  assign n15832 = ~controllable_BtoR_REQ1 & ~n15831;
  assign n15833 = controllable_BtoR_REQ0 & ~n15832;
  assign n15834 = ~controllable_BtoR_REQ1 & ~n7840;
  assign n15835 = ~controllable_BtoR_REQ0 & ~n15834;
  assign n15836 = ~n15833 & ~n15835;
  assign n15837 = ~i_RtoB_ACK0 & ~n15836;
  assign n15838 = ~i_RtoB_ACK0 & ~n15837;
  assign n15839 = controllable_DEQ & ~n15838;
  assign n15840 = ~n10413 & ~n15803;
  assign n15841 = ~controllable_BtoR_REQ1 & ~n15840;
  assign n15842 = ~controllable_BtoR_REQ1 & ~n15841;
  assign n15843 = controllable_BtoR_REQ0 & ~n15842;
  assign n15844 = ~n15800 & ~n15843;
  assign n15845 = ~i_RtoB_ACK0 & ~n15844;
  assign n15846 = ~n15802 & ~n15845;
  assign n15847 = ~controllable_DEQ & ~n15846;
  assign n15848 = ~n15839 & ~n15847;
  assign n15849 = i_FULL & ~n15848;
  assign n15850 = ~controllable_BtoR_REQ1 & ~n7818;
  assign n15851 = ~controllable_BtoR_REQ1 & ~n15850;
  assign n15852 = controllable_BtoR_REQ0 & ~n15851;
  assign n15853 = ~controllable_BtoR_REQ0 & ~n15814;
  assign n15854 = ~n15852 & ~n15853;
  assign n15855 = ~i_RtoB_ACK0 & ~n15854;
  assign n15856 = ~i_RtoB_ACK0 & ~n15855;
  assign n15857 = controllable_DEQ & ~n15856;
  assign n15858 = ~controllable_BtoR_REQ1 & ~n13676;
  assign n15859 = ~controllable_BtoR_REQ0 & ~n15858;
  assign n15860 = ~n15807 & ~n15859;
  assign n15861 = ~i_RtoB_ACK0 & ~n15860;
  assign n15862 = ~n15802 & ~n15861;
  assign n15863 = ~controllable_DEQ & ~n15862;
  assign n15864 = ~n15857 & ~n15863;
  assign n15865 = ~i_FULL & ~n15864;
  assign n15866 = ~n15849 & ~n15865;
  assign n15867 = ~i_nEMPTY & ~n15866;
  assign n15868 = ~n15830 & ~n15867;
  assign n15869 = ~controllable_BtoS_ACK0 & ~n15868;
  assign n15870 = ~n15794 & ~n15869;
  assign n15871 = n4465 & ~n15870;
  assign n15872 = ~n14811 & ~n15869;
  assign n15873 = ~n4465 & ~n15872;
  assign n15874 = ~n15871 & ~n15873;
  assign n15875 = i_StoB_REQ10 & ~n15874;
  assign n15876 = ~i_RtoB_ACK1 & ~n7928;
  assign n15877 = ~n7886 & ~n15876;
  assign n15878 = ~controllable_BtoR_REQ1 & ~n15877;
  assign n15879 = ~controllable_BtoR_REQ1 & ~n15878;
  assign n15880 = controllable_BtoR_REQ0 & ~n15879;
  assign n15881 = ~controllable_BtoR_REQ1 & ~n7917;
  assign n15882 = ~controllable_BtoR_REQ0 & ~n15881;
  assign n15883 = ~n15880 & ~n15882;
  assign n15884 = i_RtoB_ACK0 & ~n15883;
  assign n15885 = i_RtoB_ACK1 & ~n7902;
  assign n15886 = ~n7932 & ~n15885;
  assign n15887 = ~controllable_BtoR_REQ1 & ~n15886;
  assign n15888 = ~controllable_BtoR_REQ1 & ~n15887;
  assign n15889 = controllable_BtoR_REQ0 & ~n15888;
  assign n15890 = ~controllable_BtoR_REQ1 & ~n7940;
  assign n15891 = ~controllable_BtoR_REQ0 & ~n15890;
  assign n15892 = ~n15889 & ~n15891;
  assign n15893 = ~i_RtoB_ACK0 & ~n15892;
  assign n15894 = ~n15884 & ~n15893;
  assign n15895 = controllable_DEQ & ~n15894;
  assign n15896 = ~n7947 & ~n7958;
  assign n15897 = ~controllable_BtoR_REQ1 & ~n15896;
  assign n15898 = ~controllable_BtoR_REQ1 & ~n15897;
  assign n15899 = controllable_BtoR_REQ0 & ~n15898;
  assign n15900 = ~controllable_BtoR_REQ1 & ~n7951;
  assign n15901 = ~controllable_BtoR_REQ0 & ~n15900;
  assign n15902 = ~n15899 & ~n15901;
  assign n15903 = i_RtoB_ACK0 & ~n15902;
  assign n15904 = i_RtoB_ACK1 & ~n7900;
  assign n15905 = ~n7958 & ~n15904;
  assign n15906 = ~controllable_BtoR_REQ1 & ~n15905;
  assign n15907 = ~controllable_BtoR_REQ1 & ~n15906;
  assign n15908 = controllable_BtoR_REQ0 & ~n15907;
  assign n15909 = ~controllable_BtoR_REQ1 & ~n7960;
  assign n15910 = ~controllable_BtoR_REQ0 & ~n15909;
  assign n15911 = ~n15908 & ~n15910;
  assign n15912 = ~i_RtoB_ACK0 & ~n15911;
  assign n15913 = ~n15903 & ~n15912;
  assign n15914 = ~controllable_DEQ & ~n15913;
  assign n15915 = ~n15895 & ~n15914;
  assign n15916 = i_FULL & ~n15915;
  assign n15917 = ~i_RtoB_ACK1 & ~n7969;
  assign n15918 = ~n7886 & ~n15917;
  assign n15919 = ~controllable_BtoR_REQ1 & ~n15918;
  assign n15920 = ~controllable_BtoR_REQ1 & ~n15919;
  assign n15921 = controllable_BtoR_REQ0 & ~n15920;
  assign n15922 = ~n15882 & ~n15921;
  assign n15923 = i_RtoB_ACK0 & ~n15922;
  assign n15924 = ~n7972 & ~n15885;
  assign n15925 = ~controllable_BtoR_REQ1 & ~n15924;
  assign n15926 = ~controllable_BtoR_REQ1 & ~n15925;
  assign n15927 = controllable_BtoR_REQ0 & ~n15926;
  assign n15928 = ~controllable_BtoR_REQ1 & ~n7977;
  assign n15929 = ~controllable_BtoR_REQ0 & ~n15928;
  assign n15930 = ~n15927 & ~n15929;
  assign n15931 = ~i_RtoB_ACK0 & ~n15930;
  assign n15932 = ~n15923 & ~n15931;
  assign n15933 = controllable_DEQ & ~n15932;
  assign n15934 = ~n7938 & ~n7947;
  assign n15935 = ~controllable_BtoR_REQ1 & ~n15934;
  assign n15936 = ~controllable_BtoR_REQ1 & ~n15935;
  assign n15937 = controllable_BtoR_REQ0 & ~n15936;
  assign n15938 = ~n15901 & ~n15937;
  assign n15939 = i_RtoB_ACK0 & ~n15938;
  assign n15940 = ~n7938 & ~n15904;
  assign n15941 = ~controllable_BtoR_REQ1 & ~n15940;
  assign n15942 = ~controllable_BtoR_REQ1 & ~n15941;
  assign n15943 = controllable_BtoR_REQ0 & ~n15942;
  assign n15944 = ~controllable_BtoR_REQ1 & ~n7986;
  assign n15945 = ~controllable_BtoR_REQ0 & ~n15944;
  assign n15946 = ~n15943 & ~n15945;
  assign n15947 = ~i_RtoB_ACK0 & ~n15946;
  assign n15948 = ~n15939 & ~n15947;
  assign n15949 = ~controllable_DEQ & ~n15948;
  assign n15950 = ~n15933 & ~n15949;
  assign n15951 = ~i_FULL & ~n15950;
  assign n15952 = ~n15916 & ~n15951;
  assign n15953 = i_nEMPTY & ~n15952;
  assign n15954 = ~i_RtoB_ACK1 & ~n7997;
  assign n15955 = ~i_RtoB_ACK1 & ~n15954;
  assign n15956 = ~controllable_BtoR_REQ1 & ~n15955;
  assign n15957 = ~controllable_BtoR_REQ1 & ~n15956;
  assign n15958 = controllable_BtoR_REQ0 & ~n15957;
  assign n15959 = controllable_BtoR_REQ0 & ~n15958;
  assign n15960 = i_RtoB_ACK0 & ~n15959;
  assign n15961 = ~i_RtoB_ACK1 & ~n8000;
  assign n15962 = ~controllable_BtoR_REQ1 & ~n15961;
  assign n15963 = ~controllable_BtoR_REQ1 & ~n15962;
  assign n15964 = controllable_BtoR_REQ0 & ~n15963;
  assign n15965 = ~controllable_BtoR_REQ1 & ~n8006;
  assign n15966 = ~controllable_BtoR_REQ0 & ~n15965;
  assign n15967 = ~n15964 & ~n15966;
  assign n15968 = ~i_RtoB_ACK0 & ~n15967;
  assign n15969 = ~n15960 & ~n15968;
  assign n15970 = controllable_DEQ & ~n15969;
  assign n15971 = ~n7886 & ~n8015;
  assign n15972 = ~controllable_BtoR_REQ1 & ~n15971;
  assign n15973 = ~controllable_BtoR_REQ1 & ~n15972;
  assign n15974 = controllable_BtoR_REQ0 & ~n15973;
  assign n15975 = ~n15882 & ~n15974;
  assign n15976 = i_RtoB_ACK0 & ~n15975;
  assign n15977 = ~n8015 & ~n15885;
  assign n15978 = ~controllable_BtoR_REQ1 & ~n15977;
  assign n15979 = ~controllable_BtoR_REQ1 & ~n15978;
  assign n15980 = controllable_BtoR_REQ0 & ~n15979;
  assign n15981 = ~controllable_BtoR_REQ1 & ~n8017;
  assign n15982 = ~controllable_BtoR_REQ0 & ~n15981;
  assign n15983 = ~n15980 & ~n15982;
  assign n15984 = ~i_RtoB_ACK0 & ~n15983;
  assign n15985 = ~n15976 & ~n15984;
  assign n15986 = ~controllable_DEQ & ~n15985;
  assign n15987 = ~n15970 & ~n15986;
  assign n15988 = i_FULL & ~n15987;
  assign n15989 = ~i_RtoB_ACK1 & ~n7883;
  assign n15990 = ~i_RtoB_ACK1 & ~n15989;
  assign n15991 = ~controllable_BtoR_REQ1 & ~n15990;
  assign n15992 = ~controllable_BtoR_REQ1 & ~n15991;
  assign n15993 = controllable_BtoR_REQ0 & ~n15992;
  assign n15994 = controllable_BtoR_REQ0 & ~n15993;
  assign n15995 = i_RtoB_ACK0 & ~n15994;
  assign n15996 = ~i_RtoB_ACK1 & ~n7948;
  assign n15997 = ~controllable_BtoR_REQ1 & ~n15996;
  assign n15998 = ~controllable_BtoR_REQ1 & ~n15997;
  assign n15999 = controllable_BtoR_REQ0 & ~n15998;
  assign n16000 = ~controllable_BtoR_REQ1 & ~n8027;
  assign n16001 = ~controllable_BtoR_REQ0 & ~n16000;
  assign n16002 = ~n15999 & ~n16001;
  assign n16003 = ~i_RtoB_ACK0 & ~n16002;
  assign n16004 = ~n15995 & ~n16003;
  assign n16005 = controllable_DEQ & ~n16004;
  assign n16006 = ~controllable_BtoR_REQ1 & ~n8035;
  assign n16007 = ~controllable_BtoR_REQ0 & ~n16006;
  assign n16008 = ~n15889 & ~n16007;
  assign n16009 = ~i_RtoB_ACK0 & ~n16008;
  assign n16010 = ~n15884 & ~n16009;
  assign n16011 = ~controllable_DEQ & ~n16010;
  assign n16012 = ~n16005 & ~n16011;
  assign n16013 = ~i_FULL & ~n16012;
  assign n16014 = ~n15988 & ~n16013;
  assign n16015 = ~i_nEMPTY & ~n16014;
  assign n16016 = ~n15953 & ~n16015;
  assign n16017 = controllable_BtoS_ACK0 & ~n16016;
  assign n16018 = ~i_RtoB_ACK1 & ~n8092;
  assign n16019 = ~n8057 & ~n16018;
  assign n16020 = ~controllable_BtoR_REQ1 & ~n16019;
  assign n16021 = ~controllable_BtoR_REQ1 & ~n16020;
  assign n16022 = controllable_BtoR_REQ0 & ~n16021;
  assign n16023 = ~controllable_BtoR_REQ1 & ~n8084;
  assign n16024 = ~controllable_BtoR_REQ0 & ~n16023;
  assign n16025 = ~n16022 & ~n16024;
  assign n16026 = i_RtoB_ACK0 & ~n16025;
  assign n16027 = i_RtoB_ACK1 & ~n8071;
  assign n16028 = ~n8096 & ~n16027;
  assign n16029 = ~controllable_BtoR_REQ1 & ~n16028;
  assign n16030 = ~controllable_BtoR_REQ1 & ~n16029;
  assign n16031 = controllable_BtoR_REQ0 & ~n16030;
  assign n16032 = ~controllable_BtoR_REQ1 & ~n8104;
  assign n16033 = ~controllable_BtoR_REQ0 & ~n16032;
  assign n16034 = ~n16031 & ~n16033;
  assign n16035 = ~i_RtoB_ACK0 & ~n16034;
  assign n16036 = ~n16026 & ~n16035;
  assign n16037 = controllable_DEQ & ~n16036;
  assign n16038 = ~n8111 & ~n8122;
  assign n16039 = ~controllable_BtoR_REQ1 & ~n16038;
  assign n16040 = ~controllable_BtoR_REQ1 & ~n16039;
  assign n16041 = controllable_BtoR_REQ0 & ~n16040;
  assign n16042 = ~controllable_BtoR_REQ1 & ~n8115;
  assign n16043 = ~controllable_BtoR_REQ0 & ~n16042;
  assign n16044 = ~n16041 & ~n16043;
  assign n16045 = i_RtoB_ACK0 & ~n16044;
  assign n16046 = i_RtoB_ACK1 & ~n8069;
  assign n16047 = ~n8122 & ~n16046;
  assign n16048 = ~controllable_BtoR_REQ1 & ~n16047;
  assign n16049 = ~controllable_BtoR_REQ1 & ~n16048;
  assign n16050 = controllable_BtoR_REQ0 & ~n16049;
  assign n16051 = ~controllable_BtoR_REQ1 & ~n8124;
  assign n16052 = ~controllable_BtoR_REQ0 & ~n16051;
  assign n16053 = ~n16050 & ~n16052;
  assign n16054 = ~i_RtoB_ACK0 & ~n16053;
  assign n16055 = ~n16045 & ~n16054;
  assign n16056 = ~controllable_DEQ & ~n16055;
  assign n16057 = ~n16037 & ~n16056;
  assign n16058 = i_FULL & ~n16057;
  assign n16059 = ~i_RtoB_ACK1 & ~n8133;
  assign n16060 = ~n8057 & ~n16059;
  assign n16061 = ~controllable_BtoR_REQ1 & ~n16060;
  assign n16062 = ~controllable_BtoR_REQ1 & ~n16061;
  assign n16063 = controllable_BtoR_REQ0 & ~n16062;
  assign n16064 = ~n16024 & ~n16063;
  assign n16065 = i_RtoB_ACK0 & ~n16064;
  assign n16066 = ~n8136 & ~n16027;
  assign n16067 = ~controllable_BtoR_REQ1 & ~n16066;
  assign n16068 = ~controllable_BtoR_REQ1 & ~n16067;
  assign n16069 = controllable_BtoR_REQ0 & ~n16068;
  assign n16070 = ~controllable_BtoR_REQ1 & ~n8141;
  assign n16071 = ~controllable_BtoR_REQ0 & ~n16070;
  assign n16072 = ~n16069 & ~n16071;
  assign n16073 = ~i_RtoB_ACK0 & ~n16072;
  assign n16074 = ~n16065 & ~n16073;
  assign n16075 = controllable_DEQ & ~n16074;
  assign n16076 = ~n8102 & ~n8111;
  assign n16077 = ~controllable_BtoR_REQ1 & ~n16076;
  assign n16078 = ~controllable_BtoR_REQ1 & ~n16077;
  assign n16079 = controllable_BtoR_REQ0 & ~n16078;
  assign n16080 = ~n16043 & ~n16079;
  assign n16081 = i_RtoB_ACK0 & ~n16080;
  assign n16082 = ~n8102 & ~n16046;
  assign n16083 = ~controllable_BtoR_REQ1 & ~n16082;
  assign n16084 = ~controllable_BtoR_REQ1 & ~n16083;
  assign n16085 = controllable_BtoR_REQ0 & ~n16084;
  assign n16086 = ~controllable_BtoR_REQ1 & ~n8150;
  assign n16087 = ~controllable_BtoR_REQ0 & ~n16086;
  assign n16088 = ~n16085 & ~n16087;
  assign n16089 = ~i_RtoB_ACK0 & ~n16088;
  assign n16090 = ~n16081 & ~n16089;
  assign n16091 = ~controllable_DEQ & ~n16090;
  assign n16092 = ~n16075 & ~n16091;
  assign n16093 = ~i_FULL & ~n16092;
  assign n16094 = ~n16058 & ~n16093;
  assign n16095 = i_nEMPTY & ~n16094;
  assign n16096 = ~i_RtoB_ACK1 & ~n8161;
  assign n16097 = ~i_RtoB_ACK1 & ~n16096;
  assign n16098 = ~controllable_BtoR_REQ1 & ~n16097;
  assign n16099 = ~controllable_BtoR_REQ1 & ~n16098;
  assign n16100 = controllable_BtoR_REQ0 & ~n16099;
  assign n16101 = controllable_BtoR_REQ0 & ~n16100;
  assign n16102 = i_RtoB_ACK0 & ~n16101;
  assign n16103 = ~i_RtoB_ACK1 & ~n8164;
  assign n16104 = ~controllable_BtoR_REQ1 & ~n16103;
  assign n16105 = ~controllable_BtoR_REQ1 & ~n16104;
  assign n16106 = controllable_BtoR_REQ0 & ~n16105;
  assign n16107 = ~controllable_BtoR_REQ1 & ~n8170;
  assign n16108 = ~controllable_BtoR_REQ0 & ~n16107;
  assign n16109 = ~n16106 & ~n16108;
  assign n16110 = ~i_RtoB_ACK0 & ~n16109;
  assign n16111 = ~n16102 & ~n16110;
  assign n16112 = controllable_DEQ & ~n16111;
  assign n16113 = ~n8057 & ~n8179;
  assign n16114 = ~controllable_BtoR_REQ1 & ~n16113;
  assign n16115 = ~controllable_BtoR_REQ1 & ~n16114;
  assign n16116 = controllable_BtoR_REQ0 & ~n16115;
  assign n16117 = ~n16024 & ~n16116;
  assign n16118 = i_RtoB_ACK0 & ~n16117;
  assign n16119 = ~n8179 & ~n16027;
  assign n16120 = ~controllable_BtoR_REQ1 & ~n16119;
  assign n16121 = ~controllable_BtoR_REQ1 & ~n16120;
  assign n16122 = controllable_BtoR_REQ0 & ~n16121;
  assign n16123 = ~controllable_BtoR_REQ1 & ~n8181;
  assign n16124 = ~controllable_BtoR_REQ0 & ~n16123;
  assign n16125 = ~n16122 & ~n16124;
  assign n16126 = ~i_RtoB_ACK0 & ~n16125;
  assign n16127 = ~n16118 & ~n16126;
  assign n16128 = ~controllable_DEQ & ~n16127;
  assign n16129 = ~n16112 & ~n16128;
  assign n16130 = i_FULL & ~n16129;
  assign n16131 = ~i_RtoB_ACK1 & ~n8054;
  assign n16132 = ~i_RtoB_ACK1 & ~n16131;
  assign n16133 = ~controllable_BtoR_REQ1 & ~n16132;
  assign n16134 = ~controllable_BtoR_REQ1 & ~n16133;
  assign n16135 = controllable_BtoR_REQ0 & ~n16134;
  assign n16136 = controllable_BtoR_REQ0 & ~n16135;
  assign n16137 = i_RtoB_ACK0 & ~n16136;
  assign n16138 = ~i_RtoB_ACK1 & ~n8112;
  assign n16139 = ~controllable_BtoR_REQ1 & ~n16138;
  assign n16140 = ~controllable_BtoR_REQ1 & ~n16139;
  assign n16141 = controllable_BtoR_REQ0 & ~n16140;
  assign n16142 = ~controllable_BtoR_REQ1 & ~n8191;
  assign n16143 = ~controllable_BtoR_REQ0 & ~n16142;
  assign n16144 = ~n16141 & ~n16143;
  assign n16145 = ~i_RtoB_ACK0 & ~n16144;
  assign n16146 = ~n16137 & ~n16145;
  assign n16147 = controllable_DEQ & ~n16146;
  assign n16148 = ~controllable_BtoR_REQ1 & ~n8199;
  assign n16149 = ~controllable_BtoR_REQ0 & ~n16148;
  assign n16150 = ~n16031 & ~n16149;
  assign n16151 = ~i_RtoB_ACK0 & ~n16150;
  assign n16152 = ~n16026 & ~n16151;
  assign n16153 = ~controllable_DEQ & ~n16152;
  assign n16154 = ~n16147 & ~n16153;
  assign n16155 = ~i_FULL & ~n16154;
  assign n16156 = ~n16130 & ~n16155;
  assign n16157 = ~i_nEMPTY & ~n16156;
  assign n16158 = ~n16095 & ~n16157;
  assign n16159 = ~controllable_BtoS_ACK0 & ~n16158;
  assign n16160 = ~n16017 & ~n16159;
  assign n16161 = n4465 & ~n16160;
  assign n16162 = ~i_RtoB_ACK1 & ~n8232;
  assign n16163 = ~n7054 & ~n16162;
  assign n16164 = ~controllable_BtoR_REQ1 & ~n16163;
  assign n16165 = ~controllable_BtoR_REQ1 & ~n16164;
  assign n16166 = controllable_BtoR_REQ0 & ~n16165;
  assign n16167 = ~controllable_BtoR_REQ1 & ~n8227;
  assign n16168 = ~controllable_BtoR_REQ0 & ~n16167;
  assign n16169 = ~n16166 & ~n16168;
  assign n16170 = i_RtoB_ACK0 & ~n16169;
  assign n16171 = i_RtoB_ACK1 & ~n8218;
  assign n16172 = ~n8236 & ~n16171;
  assign n16173 = ~controllable_BtoR_REQ1 & ~n16172;
  assign n16174 = ~controllable_BtoR_REQ1 & ~n16173;
  assign n16175 = controllable_BtoR_REQ0 & ~n16174;
  assign n16176 = ~controllable_BtoR_REQ1 & ~n8242;
  assign n16177 = ~controllable_BtoR_REQ0 & ~n16176;
  assign n16178 = ~n16175 & ~n16177;
  assign n16179 = ~i_RtoB_ACK0 & ~n16178;
  assign n16180 = ~n16170 & ~n16179;
  assign n16181 = controllable_DEQ & ~n16180;
  assign n16182 = ~n7111 & ~n8240;
  assign n16183 = ~controllable_BtoR_REQ1 & ~n16182;
  assign n16184 = ~controllable_BtoR_REQ1 & ~n16183;
  assign n16185 = controllable_BtoR_REQ0 & ~n16184;
  assign n16186 = ~controllable_BtoR_REQ1 & ~n8252;
  assign n16187 = ~controllable_BtoR_REQ0 & ~n16186;
  assign n16188 = ~n16185 & ~n16187;
  assign n16189 = i_RtoB_ACK0 & ~n16188;
  assign n16190 = i_RtoB_ACK1 & ~n8216;
  assign n16191 = ~n8240 & ~n16190;
  assign n16192 = ~controllable_BtoR_REQ1 & ~n16191;
  assign n16193 = ~controllable_BtoR_REQ1 & ~n16192;
  assign n16194 = controllable_BtoR_REQ0 & ~n16193;
  assign n16195 = ~n16187 & ~n16194;
  assign n16196 = ~i_RtoB_ACK0 & ~n16195;
  assign n16197 = ~n16189 & ~n16196;
  assign n16198 = ~controllable_DEQ & ~n16197;
  assign n16199 = ~n16181 & ~n16198;
  assign n16200 = i_nEMPTY & ~n16199;
  assign n16201 = ~i_RtoB_ACK1 & ~n8265;
  assign n16202 = ~controllable_BtoR_REQ1 & ~n16201;
  assign n16203 = ~controllable_BtoR_REQ1 & ~n16202;
  assign n16204 = controllable_BtoR_REQ0 & ~n16203;
  assign n16205 = ~controllable_BtoR_REQ1 & ~n8272;
  assign n16206 = ~controllable_BtoR_REQ0 & ~n16205;
  assign n16207 = ~n16204 & ~n16206;
  assign n16208 = ~i_RtoB_ACK0 & ~n16207;
  assign n16209 = ~n15217 & ~n16208;
  assign n16210 = controllable_DEQ & ~n16209;
  assign n16211 = ~n7054 & ~n8615;
  assign n16212 = ~controllable_BtoR_REQ1 & ~n16211;
  assign n16213 = ~controllable_BtoR_REQ1 & ~n16212;
  assign n16214 = controllable_BtoR_REQ0 & ~n16213;
  assign n16215 = ~n16168 & ~n16214;
  assign n16216 = i_RtoB_ACK0 & ~n16215;
  assign n16217 = ~n8615 & ~n16171;
  assign n16218 = ~controllable_BtoR_REQ1 & ~n16217;
  assign n16219 = ~controllable_BtoR_REQ1 & ~n16218;
  assign n16220 = controllable_BtoR_REQ0 & ~n16219;
  assign n16221 = ~n16168 & ~n16220;
  assign n16222 = ~i_RtoB_ACK0 & ~n16221;
  assign n16223 = ~n16216 & ~n16222;
  assign n16224 = ~controllable_DEQ & ~n16223;
  assign n16225 = ~n16210 & ~n16224;
  assign n16226 = i_FULL & ~n16225;
  assign n16227 = ~i_RtoB_ACK1 & ~n8249;
  assign n16228 = ~controllable_BtoR_REQ1 & ~n16227;
  assign n16229 = ~controllable_BtoR_REQ1 & ~n16228;
  assign n16230 = controllable_BtoR_REQ0 & ~n16229;
  assign n16231 = ~controllable_BtoR_REQ1 & ~n8287;
  assign n16232 = ~controllable_BtoR_REQ0 & ~n16231;
  assign n16233 = ~n16230 & ~n16232;
  assign n16234 = ~i_RtoB_ACK0 & ~n16233;
  assign n16235 = ~n15245 & ~n16234;
  assign n16236 = controllable_DEQ & ~n16235;
  assign n16237 = ~controllable_BtoR_REQ1 & ~n8295;
  assign n16238 = ~controllable_BtoR_REQ0 & ~n16237;
  assign n16239 = ~n16175 & ~n16238;
  assign n16240 = ~i_RtoB_ACK0 & ~n16239;
  assign n16241 = ~n16170 & ~n16240;
  assign n16242 = ~controllable_DEQ & ~n16241;
  assign n16243 = ~n16236 & ~n16242;
  assign n16244 = ~i_FULL & ~n16243;
  assign n16245 = ~n16226 & ~n16244;
  assign n16246 = ~i_nEMPTY & ~n16245;
  assign n16247 = ~n16200 & ~n16246;
  assign n16248 = controllable_BtoS_ACK0 & ~n16247;
  assign n16249 = ~i_RtoB_ACK1 & ~n8333;
  assign n16250 = ~n8313 & ~n16249;
  assign n16251 = ~controllable_BtoR_REQ1 & ~n16250;
  assign n16252 = ~controllable_BtoR_REQ1 & ~n16251;
  assign n16253 = controllable_BtoR_REQ0 & ~n16252;
  assign n16254 = ~controllable_BtoR_REQ1 & ~n8327;
  assign n16255 = ~controllable_BtoR_REQ0 & ~n16254;
  assign n16256 = ~n16253 & ~n16255;
  assign n16257 = i_RtoB_ACK0 & ~n16256;
  assign n16258 = i_RtoB_ACK1 & ~n8318;
  assign n16259 = ~n8337 & ~n16258;
  assign n16260 = ~controllable_BtoR_REQ1 & ~n16259;
  assign n16261 = ~controllable_BtoR_REQ1 & ~n16260;
  assign n16262 = controllable_BtoR_REQ0 & ~n16261;
  assign n16263 = ~controllable_BtoR_REQ1 & ~n8345;
  assign n16264 = ~controllable_BtoR_REQ0 & ~n16263;
  assign n16265 = ~n16262 & ~n16264;
  assign n16266 = ~i_RtoB_ACK0 & ~n16265;
  assign n16267 = ~n16257 & ~n16266;
  assign n16268 = controllable_DEQ & ~n16267;
  assign n16269 = ~n8122 & ~n8352;
  assign n16270 = ~controllable_BtoR_REQ1 & ~n16269;
  assign n16271 = ~controllable_BtoR_REQ1 & ~n16270;
  assign n16272 = controllable_BtoR_REQ0 & ~n16271;
  assign n16273 = ~controllable_BtoR_REQ1 & ~n8356;
  assign n16274 = ~controllable_BtoR_REQ0 & ~n16273;
  assign n16275 = ~n16272 & ~n16274;
  assign n16276 = i_RtoB_ACK0 & ~n16275;
  assign n16277 = i_RtoB_ACK1 & ~n8316;
  assign n16278 = ~n8122 & ~n16277;
  assign n16279 = ~controllable_BtoR_REQ1 & ~n16278;
  assign n16280 = ~controllable_BtoR_REQ1 & ~n16279;
  assign n16281 = controllable_BtoR_REQ0 & ~n16280;
  assign n16282 = ~controllable_BtoR_REQ1 & ~n8363;
  assign n16283 = ~controllable_BtoR_REQ0 & ~n16282;
  assign n16284 = ~n16281 & ~n16283;
  assign n16285 = ~i_RtoB_ACK0 & ~n16284;
  assign n16286 = ~n16276 & ~n16285;
  assign n16287 = ~controllable_DEQ & ~n16286;
  assign n16288 = ~n16268 & ~n16287;
  assign n16289 = i_FULL & ~n16288;
  assign n16290 = ~i_RtoB_ACK1 & ~n8372;
  assign n16291 = ~n8313 & ~n16290;
  assign n16292 = ~controllable_BtoR_REQ1 & ~n16291;
  assign n16293 = ~controllable_BtoR_REQ1 & ~n16292;
  assign n16294 = controllable_BtoR_REQ0 & ~n16293;
  assign n16295 = ~n16255 & ~n16294;
  assign n16296 = i_RtoB_ACK0 & ~n16295;
  assign n16297 = ~n8375 & ~n16258;
  assign n16298 = ~controllable_BtoR_REQ1 & ~n16297;
  assign n16299 = ~controllable_BtoR_REQ1 & ~n16298;
  assign n16300 = controllable_BtoR_REQ0 & ~n16299;
  assign n16301 = ~controllable_BtoR_REQ1 & ~n8380;
  assign n16302 = ~controllable_BtoR_REQ0 & ~n16301;
  assign n16303 = ~n16300 & ~n16302;
  assign n16304 = ~i_RtoB_ACK0 & ~n16303;
  assign n16305 = ~n16296 & ~n16304;
  assign n16306 = controllable_DEQ & ~n16305;
  assign n16307 = ~n8343 & ~n8352;
  assign n16308 = ~controllable_BtoR_REQ1 & ~n16307;
  assign n16309 = ~controllable_BtoR_REQ1 & ~n16308;
  assign n16310 = controllable_BtoR_REQ0 & ~n16309;
  assign n16311 = ~n16274 & ~n16310;
  assign n16312 = i_RtoB_ACK0 & ~n16311;
  assign n16313 = ~n8343 & ~n16277;
  assign n16314 = ~controllable_BtoR_REQ1 & ~n16313;
  assign n16315 = ~controllable_BtoR_REQ1 & ~n16314;
  assign n16316 = controllable_BtoR_REQ0 & ~n16315;
  assign n16317 = ~controllable_BtoR_REQ1 & ~n8389;
  assign n16318 = ~controllable_BtoR_REQ0 & ~n16317;
  assign n16319 = ~n16316 & ~n16318;
  assign n16320 = ~i_RtoB_ACK0 & ~n16319;
  assign n16321 = ~n16312 & ~n16320;
  assign n16322 = ~controllable_DEQ & ~n16321;
  assign n16323 = ~n16306 & ~n16322;
  assign n16324 = ~i_FULL & ~n16323;
  assign n16325 = ~n16289 & ~n16324;
  assign n16326 = i_nEMPTY & ~n16325;
  assign n16327 = ~i_RtoB_ACK1 & ~n8400;
  assign n16328 = ~i_RtoB_ACK1 & ~n16327;
  assign n16329 = ~controllable_BtoR_REQ1 & ~n16328;
  assign n16330 = ~controllable_BtoR_REQ1 & ~n16329;
  assign n16331 = controllable_BtoR_REQ0 & ~n16330;
  assign n16332 = controllable_BtoR_REQ0 & ~n16331;
  assign n16333 = i_RtoB_ACK0 & ~n16332;
  assign n16334 = ~i_RtoB_ACK1 & ~n8403;
  assign n16335 = ~controllable_BtoR_REQ1 & ~n16334;
  assign n16336 = ~controllable_BtoR_REQ1 & ~n16335;
  assign n16337 = controllable_BtoR_REQ0 & ~n16336;
  assign n16338 = ~controllable_BtoR_REQ1 & ~n8409;
  assign n16339 = ~controllable_BtoR_REQ0 & ~n16338;
  assign n16340 = ~n16337 & ~n16339;
  assign n16341 = ~i_RtoB_ACK0 & ~n16340;
  assign n16342 = ~n16333 & ~n16341;
  assign n16343 = controllable_DEQ & ~n16342;
  assign n16344 = ~n8179 & ~n8313;
  assign n16345 = ~controllable_BtoR_REQ1 & ~n16344;
  assign n16346 = ~controllable_BtoR_REQ1 & ~n16345;
  assign n16347 = controllable_BtoR_REQ0 & ~n16346;
  assign n16348 = ~n16255 & ~n16347;
  assign n16349 = i_RtoB_ACK0 & ~n16348;
  assign n16350 = ~n8179 & ~n16258;
  assign n16351 = ~controllable_BtoR_REQ1 & ~n16350;
  assign n16352 = ~controllable_BtoR_REQ1 & ~n16351;
  assign n16353 = controllable_BtoR_REQ0 & ~n16352;
  assign n16354 = ~controllable_BtoR_REQ1 & ~n8417;
  assign n16355 = ~controllable_BtoR_REQ0 & ~n16354;
  assign n16356 = ~n16353 & ~n16355;
  assign n16357 = ~i_RtoB_ACK0 & ~n16356;
  assign n16358 = ~n16349 & ~n16357;
  assign n16359 = ~controllable_DEQ & ~n16358;
  assign n16360 = ~n16343 & ~n16359;
  assign n16361 = i_FULL & ~n16360;
  assign n16362 = ~i_RtoB_ACK1 & ~n8310;
  assign n16363 = ~i_RtoB_ACK1 & ~n16362;
  assign n16364 = ~controllable_BtoR_REQ1 & ~n16363;
  assign n16365 = ~controllable_BtoR_REQ1 & ~n16364;
  assign n16366 = controllable_BtoR_REQ0 & ~n16365;
  assign n16367 = controllable_BtoR_REQ0 & ~n16366;
  assign n16368 = i_RtoB_ACK0 & ~n16367;
  assign n16369 = ~i_RtoB_ACK1 & ~n8353;
  assign n16370 = ~controllable_BtoR_REQ1 & ~n16369;
  assign n16371 = ~controllable_BtoR_REQ1 & ~n16370;
  assign n16372 = controllable_BtoR_REQ0 & ~n16371;
  assign n16373 = ~controllable_BtoR_REQ1 & ~n8427;
  assign n16374 = ~controllable_BtoR_REQ0 & ~n16373;
  assign n16375 = ~n16372 & ~n16374;
  assign n16376 = ~i_RtoB_ACK0 & ~n16375;
  assign n16377 = ~n16368 & ~n16376;
  assign n16378 = controllable_DEQ & ~n16377;
  assign n16379 = ~controllable_BtoR_REQ1 & ~n8435;
  assign n16380 = ~controllable_BtoR_REQ0 & ~n16379;
  assign n16381 = ~n16262 & ~n16380;
  assign n16382 = ~i_RtoB_ACK0 & ~n16381;
  assign n16383 = ~n16257 & ~n16382;
  assign n16384 = ~controllable_DEQ & ~n16383;
  assign n16385 = ~n16378 & ~n16384;
  assign n16386 = ~i_FULL & ~n16385;
  assign n16387 = ~n16361 & ~n16386;
  assign n16388 = ~i_nEMPTY & ~n16387;
  assign n16389 = ~n16326 & ~n16388;
  assign n16390 = ~controllable_BtoS_ACK0 & ~n16389;
  assign n16391 = ~n16248 & ~n16390;
  assign n16392 = ~n4465 & ~n16391;
  assign n16393 = ~n16161 & ~n16392;
  assign n16394 = ~i_StoB_REQ10 & ~n16393;
  assign n16395 = ~n15875 & ~n16394;
  assign n16396 = controllable_BtoS_ACK10 & ~n16395;
  assign n16397 = ~i_RtoB_ACK1 & ~n8470;
  assign n16398 = ~n8461 & ~n16397;
  assign n16399 = ~controllable_BtoR_REQ1 & ~n16398;
  assign n16400 = ~controllable_BtoR_REQ1 & ~n16399;
  assign n16401 = controllable_BtoR_REQ0 & ~n16400;
  assign n16402 = ~n15882 & ~n16401;
  assign n16403 = i_RtoB_ACK0 & ~n16402;
  assign n16404 = ~i_RtoB_ACK0 & ~n15890;
  assign n16405 = ~n16403 & ~n16404;
  assign n16406 = controllable_DEQ & ~n16405;
  assign n16407 = ~n7958 & ~n8480;
  assign n16408 = ~controllable_BtoR_REQ1 & ~n16407;
  assign n16409 = ~controllable_BtoR_REQ1 & ~n16408;
  assign n16410 = controllable_BtoR_REQ0 & ~n16409;
  assign n16411 = ~n15901 & ~n16410;
  assign n16412 = i_RtoB_ACK0 & ~n16411;
  assign n16413 = ~i_RtoB_ACK0 & ~n15909;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = ~controllable_DEQ & ~n16414;
  assign n16416 = ~n16406 & ~n16415;
  assign n16417 = i_FULL & ~n16416;
  assign n16418 = ~i_RtoB_ACK1 & ~n8491;
  assign n16419 = ~n8461 & ~n16418;
  assign n16420 = ~controllable_BtoR_REQ1 & ~n16419;
  assign n16421 = ~controllable_BtoR_REQ1 & ~n16420;
  assign n16422 = controllable_BtoR_REQ0 & ~n16421;
  assign n16423 = ~n15882 & ~n16422;
  assign n16424 = i_RtoB_ACK0 & ~n16423;
  assign n16425 = ~i_RtoB_ACK0 & ~n15928;
  assign n16426 = ~n16424 & ~n16425;
  assign n16427 = controllable_DEQ & ~n16426;
  assign n16428 = ~n7938 & ~n8480;
  assign n16429 = ~controllable_BtoR_REQ1 & ~n16428;
  assign n16430 = ~controllable_BtoR_REQ1 & ~n16429;
  assign n16431 = controllable_BtoR_REQ0 & ~n16430;
  assign n16432 = ~n15901 & ~n16431;
  assign n16433 = i_RtoB_ACK0 & ~n16432;
  assign n16434 = ~i_RtoB_ACK0 & ~n15944;
  assign n16435 = ~n16433 & ~n16434;
  assign n16436 = ~controllable_DEQ & ~n16435;
  assign n16437 = ~n16427 & ~n16436;
  assign n16438 = ~i_FULL & ~n16437;
  assign n16439 = ~n16417 & ~n16438;
  assign n16440 = i_nEMPTY & ~n16439;
  assign n16441 = ~i_RtoB_ACK1 & ~n8507;
  assign n16442 = ~i_RtoB_ACK1 & ~n16441;
  assign n16443 = ~controllable_BtoR_REQ1 & ~n16442;
  assign n16444 = ~controllable_BtoR_REQ1 & ~n16443;
  assign n16445 = controllable_BtoR_REQ0 & ~n16444;
  assign n16446 = controllable_BtoR_REQ0 & ~n16445;
  assign n16447 = i_RtoB_ACK0 & ~n16446;
  assign n16448 = ~i_RtoB_ACK0 & ~n15965;
  assign n16449 = ~n16447 & ~n16448;
  assign n16450 = controllable_DEQ & ~n16449;
  assign n16451 = ~n8015 & ~n8461;
  assign n16452 = ~controllable_BtoR_REQ1 & ~n16451;
  assign n16453 = ~controllable_BtoR_REQ1 & ~n16452;
  assign n16454 = controllable_BtoR_REQ0 & ~n16453;
  assign n16455 = ~n15882 & ~n16454;
  assign n16456 = i_RtoB_ACK0 & ~n16455;
  assign n16457 = ~i_RtoB_ACK0 & ~n15981;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = ~controllable_DEQ & ~n16458;
  assign n16460 = ~n16450 & ~n16459;
  assign n16461 = i_FULL & ~n16460;
  assign n16462 = ~i_RtoB_ACK1 & ~n8458;
  assign n16463 = ~i_RtoB_ACK1 & ~n16462;
  assign n16464 = ~controllable_BtoR_REQ1 & ~n16463;
  assign n16465 = ~controllable_BtoR_REQ1 & ~n16464;
  assign n16466 = controllable_BtoR_REQ0 & ~n16465;
  assign n16467 = controllable_BtoR_REQ0 & ~n16466;
  assign n16468 = i_RtoB_ACK0 & ~n16467;
  assign n16469 = ~i_RtoB_ACK0 & ~n16000;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = controllable_DEQ & ~n16470;
  assign n16472 = ~controllable_DEQ & ~n16405;
  assign n16473 = ~n16471 & ~n16472;
  assign n16474 = ~i_FULL & ~n16473;
  assign n16475 = ~n16461 & ~n16474;
  assign n16476 = ~i_nEMPTY & ~n16475;
  assign n16477 = ~n16440 & ~n16476;
  assign n16478 = controllable_BtoS_ACK0 & ~n16477;
  assign n16479 = ~i_RtoB_ACK1 & ~n8549;
  assign n16480 = ~n8540 & ~n16479;
  assign n16481 = ~controllable_BtoR_REQ1 & ~n16480;
  assign n16482 = ~controllable_BtoR_REQ1 & ~n16481;
  assign n16483 = controllable_BtoR_REQ0 & ~n16482;
  assign n16484 = ~n16024 & ~n16483;
  assign n16485 = i_RtoB_ACK0 & ~n16484;
  assign n16486 = ~i_RtoB_ACK0 & ~n16032;
  assign n16487 = ~n16485 & ~n16486;
  assign n16488 = controllable_DEQ & ~n16487;
  assign n16489 = ~n8122 & ~n8559;
  assign n16490 = ~controllable_BtoR_REQ1 & ~n16489;
  assign n16491 = ~controllable_BtoR_REQ1 & ~n16490;
  assign n16492 = controllable_BtoR_REQ0 & ~n16491;
  assign n16493 = ~n16043 & ~n16492;
  assign n16494 = i_RtoB_ACK0 & ~n16493;
  assign n16495 = ~i_RtoB_ACK0 & ~n16051;
  assign n16496 = ~n16494 & ~n16495;
  assign n16497 = ~controllable_DEQ & ~n16496;
  assign n16498 = ~n16488 & ~n16497;
  assign n16499 = i_FULL & ~n16498;
  assign n16500 = ~i_RtoB_ACK1 & ~n8570;
  assign n16501 = ~n8540 & ~n16500;
  assign n16502 = ~controllable_BtoR_REQ1 & ~n16501;
  assign n16503 = ~controllable_BtoR_REQ1 & ~n16502;
  assign n16504 = controllable_BtoR_REQ0 & ~n16503;
  assign n16505 = ~n16024 & ~n16504;
  assign n16506 = i_RtoB_ACK0 & ~n16505;
  assign n16507 = ~i_RtoB_ACK0 & ~n16070;
  assign n16508 = ~n16506 & ~n16507;
  assign n16509 = controllable_DEQ & ~n16508;
  assign n16510 = ~n8102 & ~n8559;
  assign n16511 = ~controllable_BtoR_REQ1 & ~n16510;
  assign n16512 = ~controllable_BtoR_REQ1 & ~n16511;
  assign n16513 = controllable_BtoR_REQ0 & ~n16512;
  assign n16514 = ~n16043 & ~n16513;
  assign n16515 = i_RtoB_ACK0 & ~n16514;
  assign n16516 = ~i_RtoB_ACK0 & ~n16086;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = ~controllable_DEQ & ~n16517;
  assign n16519 = ~n16509 & ~n16518;
  assign n16520 = ~i_FULL & ~n16519;
  assign n16521 = ~n16499 & ~n16520;
  assign n16522 = i_nEMPTY & ~n16521;
  assign n16523 = ~i_RtoB_ACK1 & ~n8586;
  assign n16524 = ~i_RtoB_ACK1 & ~n16523;
  assign n16525 = ~controllable_BtoR_REQ1 & ~n16524;
  assign n16526 = ~controllable_BtoR_REQ1 & ~n16525;
  assign n16527 = controllable_BtoR_REQ0 & ~n16526;
  assign n16528 = controllable_BtoR_REQ0 & ~n16527;
  assign n16529 = i_RtoB_ACK0 & ~n16528;
  assign n16530 = ~i_RtoB_ACK0 & ~n16107;
  assign n16531 = ~n16529 & ~n16530;
  assign n16532 = controllable_DEQ & ~n16531;
  assign n16533 = ~n8179 & ~n8540;
  assign n16534 = ~controllable_BtoR_REQ1 & ~n16533;
  assign n16535 = ~controllable_BtoR_REQ1 & ~n16534;
  assign n16536 = controllable_BtoR_REQ0 & ~n16535;
  assign n16537 = ~n16024 & ~n16536;
  assign n16538 = i_RtoB_ACK0 & ~n16537;
  assign n16539 = ~i_RtoB_ACK0 & ~n16123;
  assign n16540 = ~n16538 & ~n16539;
  assign n16541 = ~controllable_DEQ & ~n16540;
  assign n16542 = ~n16532 & ~n16541;
  assign n16543 = i_FULL & ~n16542;
  assign n16544 = ~i_RtoB_ACK1 & ~n8537;
  assign n16545 = ~i_RtoB_ACK1 & ~n16544;
  assign n16546 = ~controllable_BtoR_REQ1 & ~n16545;
  assign n16547 = ~controllable_BtoR_REQ1 & ~n16546;
  assign n16548 = controllable_BtoR_REQ0 & ~n16547;
  assign n16549 = controllable_BtoR_REQ0 & ~n16548;
  assign n16550 = i_RtoB_ACK0 & ~n16549;
  assign n16551 = ~i_RtoB_ACK0 & ~n16142;
  assign n16552 = ~n16550 & ~n16551;
  assign n16553 = controllable_DEQ & ~n16552;
  assign n16554 = ~controllable_DEQ & ~n16487;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = ~i_FULL & ~n16555;
  assign n16557 = ~n16543 & ~n16556;
  assign n16558 = ~i_nEMPTY & ~n16557;
  assign n16559 = ~n16522 & ~n16558;
  assign n16560 = ~controllable_BtoS_ACK0 & ~n16559;
  assign n16561 = ~n16478 & ~n16560;
  assign n16562 = n4465 & ~n16561;
  assign n16563 = ~i_RtoB_ACK1 & ~n8622;
  assign n16564 = ~n5237 & ~n16563;
  assign n16565 = ~controllable_BtoR_REQ1 & ~n16564;
  assign n16566 = ~controllable_BtoR_REQ1 & ~n16565;
  assign n16567 = controllable_BtoR_REQ0 & ~n16566;
  assign n16568 = ~n16168 & ~n16567;
  assign n16569 = i_RtoB_ACK0 & ~n16568;
  assign n16570 = ~i_RtoB_ACK0 & ~n16176;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = controllable_DEQ & ~n16571;
  assign n16573 = ~controllable_BtoR_REQ1 & ~n8632;
  assign n16574 = ~controllable_BtoR_REQ1 & ~n16573;
  assign n16575 = controllable_BtoR_REQ0 & ~n16574;
  assign n16576 = ~n16187 & ~n16575;
  assign n16577 = i_RtoB_ACK0 & ~n16576;
  assign n16578 = ~i_RtoB_ACK0 & ~n16186;
  assign n16579 = ~n16577 & ~n16578;
  assign n16580 = ~controllable_DEQ & ~n16579;
  assign n16581 = ~n16572 & ~n16580;
  assign n16582 = i_nEMPTY & ~n16581;
  assign n16583 = ~i_RtoB_ACK0 & ~n16205;
  assign n16584 = ~n15604 & ~n16583;
  assign n16585 = controllable_DEQ & ~n16584;
  assign n16586 = ~controllable_BtoR_REQ1 & ~n8616;
  assign n16587 = ~controllable_BtoR_REQ1 & ~n16586;
  assign n16588 = controllable_BtoR_REQ0 & ~n16587;
  assign n16589 = ~n16168 & ~n16588;
  assign n16590 = i_RtoB_ACK0 & ~n16589;
  assign n16591 = ~i_RtoB_ACK0 & ~n16167;
  assign n16592 = ~n16590 & ~n16591;
  assign n16593 = ~controllable_DEQ & ~n16592;
  assign n16594 = ~n16585 & ~n16593;
  assign n16595 = i_FULL & ~n16594;
  assign n16596 = ~i_RtoB_ACK0 & ~n16231;
  assign n16597 = ~n15619 & ~n16596;
  assign n16598 = controllable_DEQ & ~n16597;
  assign n16599 = ~controllable_DEQ & ~n16571;
  assign n16600 = ~n16598 & ~n16599;
  assign n16601 = ~i_FULL & ~n16600;
  assign n16602 = ~n16595 & ~n16601;
  assign n16603 = ~i_nEMPTY & ~n16602;
  assign n16604 = ~n16582 & ~n16603;
  assign n16605 = controllable_BtoS_ACK0 & ~n16604;
  assign n16606 = ~i_RtoB_ACK1 & ~n8681;
  assign n16607 = ~n8672 & ~n16606;
  assign n16608 = ~controllable_BtoR_REQ1 & ~n16607;
  assign n16609 = ~controllable_BtoR_REQ1 & ~n16608;
  assign n16610 = controllable_BtoR_REQ0 & ~n16609;
  assign n16611 = ~n16255 & ~n16610;
  assign n16612 = i_RtoB_ACK0 & ~n16611;
  assign n16613 = ~i_RtoB_ACK0 & ~n16263;
  assign n16614 = ~n16612 & ~n16613;
  assign n16615 = controllable_DEQ & ~n16614;
  assign n16616 = ~n8122 & ~n8691;
  assign n16617 = ~controllable_BtoR_REQ1 & ~n16616;
  assign n16618 = ~controllable_BtoR_REQ1 & ~n16617;
  assign n16619 = controllable_BtoR_REQ0 & ~n16618;
  assign n16620 = ~n16274 & ~n16619;
  assign n16621 = i_RtoB_ACK0 & ~n16620;
  assign n16622 = ~i_RtoB_ACK0 & ~n16282;
  assign n16623 = ~n16621 & ~n16622;
  assign n16624 = ~controllable_DEQ & ~n16623;
  assign n16625 = ~n16615 & ~n16624;
  assign n16626 = i_FULL & ~n16625;
  assign n16627 = ~i_RtoB_ACK1 & ~n8702;
  assign n16628 = ~n8672 & ~n16627;
  assign n16629 = ~controllable_BtoR_REQ1 & ~n16628;
  assign n16630 = ~controllable_BtoR_REQ1 & ~n16629;
  assign n16631 = controllable_BtoR_REQ0 & ~n16630;
  assign n16632 = ~n16255 & ~n16631;
  assign n16633 = i_RtoB_ACK0 & ~n16632;
  assign n16634 = ~i_RtoB_ACK0 & ~n16301;
  assign n16635 = ~n16633 & ~n16634;
  assign n16636 = controllable_DEQ & ~n16635;
  assign n16637 = ~n8343 & ~n8691;
  assign n16638 = ~controllable_BtoR_REQ1 & ~n16637;
  assign n16639 = ~controllable_BtoR_REQ1 & ~n16638;
  assign n16640 = controllable_BtoR_REQ0 & ~n16639;
  assign n16641 = ~n16274 & ~n16640;
  assign n16642 = i_RtoB_ACK0 & ~n16641;
  assign n16643 = ~i_RtoB_ACK0 & ~n16317;
  assign n16644 = ~n16642 & ~n16643;
  assign n16645 = ~controllable_DEQ & ~n16644;
  assign n16646 = ~n16636 & ~n16645;
  assign n16647 = ~i_FULL & ~n16646;
  assign n16648 = ~n16626 & ~n16647;
  assign n16649 = i_nEMPTY & ~n16648;
  assign n16650 = ~i_RtoB_ACK1 & ~n8718;
  assign n16651 = ~i_RtoB_ACK1 & ~n16650;
  assign n16652 = ~controllable_BtoR_REQ1 & ~n16651;
  assign n16653 = ~controllable_BtoR_REQ1 & ~n16652;
  assign n16654 = controllable_BtoR_REQ0 & ~n16653;
  assign n16655 = controllable_BtoR_REQ0 & ~n16654;
  assign n16656 = i_RtoB_ACK0 & ~n16655;
  assign n16657 = ~i_RtoB_ACK0 & ~n16338;
  assign n16658 = ~n16656 & ~n16657;
  assign n16659 = controllable_DEQ & ~n16658;
  assign n16660 = ~n8179 & ~n8672;
  assign n16661 = ~controllable_BtoR_REQ1 & ~n16660;
  assign n16662 = ~controllable_BtoR_REQ1 & ~n16661;
  assign n16663 = controllable_BtoR_REQ0 & ~n16662;
  assign n16664 = ~n16255 & ~n16663;
  assign n16665 = i_RtoB_ACK0 & ~n16664;
  assign n16666 = ~i_RtoB_ACK0 & ~n16354;
  assign n16667 = ~n16665 & ~n16666;
  assign n16668 = ~controllable_DEQ & ~n16667;
  assign n16669 = ~n16659 & ~n16668;
  assign n16670 = i_FULL & ~n16669;
  assign n16671 = ~i_RtoB_ACK1 & ~n8669;
  assign n16672 = ~i_RtoB_ACK1 & ~n16671;
  assign n16673 = ~controllable_BtoR_REQ1 & ~n16672;
  assign n16674 = ~controllable_BtoR_REQ1 & ~n16673;
  assign n16675 = controllable_BtoR_REQ0 & ~n16674;
  assign n16676 = controllable_BtoR_REQ0 & ~n16675;
  assign n16677 = i_RtoB_ACK0 & ~n16676;
  assign n16678 = ~i_RtoB_ACK0 & ~n16373;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = controllable_DEQ & ~n16679;
  assign n16681 = ~controllable_DEQ & ~n16614;
  assign n16682 = ~n16680 & ~n16681;
  assign n16683 = ~i_FULL & ~n16682;
  assign n16684 = ~n16670 & ~n16683;
  assign n16685 = ~i_nEMPTY & ~n16684;
  assign n16686 = ~n16649 & ~n16685;
  assign n16687 = ~controllable_BtoS_ACK0 & ~n16686;
  assign n16688 = ~n16605 & ~n16687;
  assign n16689 = ~n4465 & ~n16688;
  assign n16690 = ~n16562 & ~n16689;
  assign n16691 = i_StoB_REQ10 & ~n16690;
  assign n16692 = ~n16394 & ~n16691;
  assign n16693 = ~controllable_BtoS_ACK10 & ~n16692;
  assign n16694 = ~n16396 & ~n16693;
  assign n16695 = ~n4464 & ~n16694;
  assign n16696 = ~n15719 & ~n16695;
  assign n16697 = n4463 & ~n16696;
  assign n16698 = ~n14591 & ~n14741;
  assign n16699 = i_RtoB_ACK0 & ~n16698;
  assign n16700 = ~n14602 & ~n16699;
  assign n16701 = controllable_DEQ & ~n16700;
  assign n16702 = ~n14608 & ~n14757;
  assign n16703 = i_RtoB_ACK0 & ~n16702;
  assign n16704 = ~n14617 & ~n16703;
  assign n16705 = ~controllable_DEQ & ~n16704;
  assign n16706 = ~n16701 & ~n16705;
  assign n16707 = i_nEMPTY & ~n16706;
  assign n16708 = ~n14636 & ~n16699;
  assign n16709 = ~controllable_DEQ & ~n16708;
  assign n16710 = ~n14630 & ~n16709;
  assign n16711 = i_FULL & ~n16710;
  assign n16712 = ~n14652 & ~n16699;
  assign n16713 = ~controllable_DEQ & ~n16712;
  assign n16714 = ~n14648 & ~n16713;
  assign n16715 = ~i_FULL & ~n16714;
  assign n16716 = ~n16711 & ~n16715;
  assign n16717 = ~i_nEMPTY & ~n16716;
  assign n16718 = ~n16707 & ~n16717;
  assign n16719 = controllable_BtoS_ACK0 & ~n16718;
  assign n16720 = ~i_RtoB_ACK1 & ~n8854;
  assign n16721 = ~controllable_BtoR_REQ1 & ~n16720;
  assign n16722 = ~controllable_BtoR_REQ1 & ~n16721;
  assign n16723 = controllable_BtoR_REQ0 & ~n16722;
  assign n16724 = ~n14666 & ~n16723;
  assign n16725 = i_RtoB_ACK0 & ~n16724;
  assign n16726 = ~n14677 & ~n16725;
  assign n16727 = controllable_DEQ & ~n16726;
  assign n16728 = ~controllable_BtoR_REQ1 & ~n8936;
  assign n16729 = controllable_BtoR_REQ0 & ~n16728;
  assign n16730 = ~n14683 & ~n16729;
  assign n16731 = i_RtoB_ACK0 & ~n16730;
  assign n16732 = ~n14692 & ~n16731;
  assign n16733 = ~controllable_DEQ & ~n16732;
  assign n16734 = ~n16727 & ~n16733;
  assign n16735 = i_nEMPTY & ~n16734;
  assign n16736 = ~n14711 & ~n16725;
  assign n16737 = ~controllable_DEQ & ~n16736;
  assign n16738 = ~n14705 & ~n16737;
  assign n16739 = i_FULL & ~n16738;
  assign n16740 = ~n14727 & ~n16725;
  assign n16741 = ~controllable_DEQ & ~n16740;
  assign n16742 = ~n14723 & ~n16741;
  assign n16743 = ~i_FULL & ~n16742;
  assign n16744 = ~n16739 & ~n16743;
  assign n16745 = ~i_nEMPTY & ~n16744;
  assign n16746 = ~n16735 & ~n16745;
  assign n16747 = ~controllable_BtoS_ACK0 & ~n16746;
  assign n16748 = ~n16719 & ~n16747;
  assign n16749 = n4465 & ~n16748;
  assign n16750 = ~n14817 & ~n16723;
  assign n16751 = i_RtoB_ACK0 & ~n16750;
  assign n16752 = ~n14828 & ~n16751;
  assign n16753 = controllable_DEQ & ~n16752;
  assign n16754 = ~n14834 & ~n16729;
  assign n16755 = i_RtoB_ACK0 & ~n16754;
  assign n16756 = ~n14843 & ~n16755;
  assign n16757 = ~controllable_DEQ & ~n16756;
  assign n16758 = ~n16753 & ~n16757;
  assign n16759 = i_nEMPTY & ~n16758;
  assign n16760 = ~n14862 & ~n16751;
  assign n16761 = ~controllable_DEQ & ~n16760;
  assign n16762 = ~n14856 & ~n16761;
  assign n16763 = i_FULL & ~n16762;
  assign n16764 = ~n14878 & ~n16751;
  assign n16765 = ~controllable_DEQ & ~n16764;
  assign n16766 = ~n14874 & ~n16765;
  assign n16767 = ~i_FULL & ~n16766;
  assign n16768 = ~n16763 & ~n16767;
  assign n16769 = ~i_nEMPTY & ~n16768;
  assign n16770 = ~n16759 & ~n16769;
  assign n16771 = ~controllable_BtoS_ACK0 & ~n16770;
  assign n16772 = ~n14811 & ~n16771;
  assign n16773 = ~n4465 & ~n16772;
  assign n16774 = ~n16749 & ~n16773;
  assign n16775 = i_StoB_REQ10 & ~n16774;
  assign n16776 = ~i_RtoB_ACK1 & ~n13243;
  assign n16777 = ~n5859 & ~n16776;
  assign n16778 = ~controllable_BtoR_REQ1 & ~n16777;
  assign n16779 = ~controllable_BtoR_REQ1 & ~n16778;
  assign n16780 = controllable_BtoR_REQ0 & ~n16779;
  assign n16781 = ~n14897 & ~n16780;
  assign n16782 = i_RtoB_ACK0 & ~n16781;
  assign n16783 = ~n14908 & ~n16782;
  assign n16784 = controllable_DEQ & ~n16783;
  assign n16785 = ~n6785 & ~n9510;
  assign n16786 = ~controllable_BtoR_REQ1 & ~n16785;
  assign n16787 = ~controllable_BtoR_REQ1 & ~n16786;
  assign n16788 = controllable_BtoR_REQ0 & ~n16787;
  assign n16789 = ~n14916 & ~n16788;
  assign n16790 = i_RtoB_ACK0 & ~n16789;
  assign n16791 = ~n14927 & ~n16790;
  assign n16792 = ~controllable_DEQ & ~n16791;
  assign n16793 = ~n16784 & ~n16792;
  assign n16794 = i_FULL & ~n16793;
  assign n16795 = ~n14946 & ~n16782;
  assign n16796 = controllable_DEQ & ~n16795;
  assign n16797 = ~n14962 & ~n16790;
  assign n16798 = ~controllable_DEQ & ~n16797;
  assign n16799 = ~n16796 & ~n16798;
  assign n16800 = ~i_FULL & ~n16799;
  assign n16801 = ~n16794 & ~n16800;
  assign n16802 = i_nEMPTY & ~n16801;
  assign n16803 = ~n5859 & ~n9293;
  assign n16804 = ~controllable_BtoR_REQ1 & ~n16803;
  assign n16805 = ~controllable_BtoR_REQ1 & ~n16804;
  assign n16806 = controllable_BtoR_REQ0 & ~n16805;
  assign n16807 = ~n14897 & ~n16806;
  assign n16808 = i_RtoB_ACK0 & ~n16807;
  assign n16809 = ~n14999 & ~n16808;
  assign n16810 = ~controllable_DEQ & ~n16809;
  assign n16811 = ~n14985 & ~n16810;
  assign n16812 = i_FULL & ~n16811;
  assign n16813 = ~n15024 & ~n16782;
  assign n16814 = ~controllable_DEQ & ~n16813;
  assign n16815 = ~n15020 & ~n16814;
  assign n16816 = ~i_FULL & ~n16815;
  assign n16817 = ~n16812 & ~n16816;
  assign n16818 = ~i_nEMPTY & ~n16817;
  assign n16819 = ~n16802 & ~n16818;
  assign n16820 = controllable_BtoS_ACK0 & ~n16819;
  assign n16821 = ~i_RtoB_ACK1 & ~n13307;
  assign n16822 = ~n6897 & ~n16821;
  assign n16823 = ~controllable_BtoR_REQ1 & ~n16822;
  assign n16824 = ~controllable_BtoR_REQ1 & ~n16823;
  assign n16825 = controllable_BtoR_REQ0 & ~n16824;
  assign n16826 = ~n15039 & ~n16825;
  assign n16827 = i_RtoB_ACK0 & ~n16826;
  assign n16828 = ~n15050 & ~n16827;
  assign n16829 = controllable_DEQ & ~n16828;
  assign n16830 = ~n6951 & ~n9657;
  assign n16831 = ~controllable_BtoR_REQ1 & ~n16830;
  assign n16832 = ~controllable_BtoR_REQ1 & ~n16831;
  assign n16833 = controllable_BtoR_REQ0 & ~n16832;
  assign n16834 = ~n15058 & ~n16833;
  assign n16835 = i_RtoB_ACK0 & ~n16834;
  assign n16836 = ~n15069 & ~n16835;
  assign n16837 = ~controllable_DEQ & ~n16836;
  assign n16838 = ~n16829 & ~n16837;
  assign n16839 = i_FULL & ~n16838;
  assign n16840 = ~n15088 & ~n16827;
  assign n16841 = controllable_DEQ & ~n16840;
  assign n16842 = ~n15104 & ~n16835;
  assign n16843 = ~controllable_DEQ & ~n16842;
  assign n16844 = ~n16841 & ~n16843;
  assign n16845 = ~i_FULL & ~n16844;
  assign n16846 = ~n16839 & ~n16845;
  assign n16847 = i_nEMPTY & ~n16846;
  assign n16848 = ~n6897 & ~n9624;
  assign n16849 = ~controllable_BtoR_REQ1 & ~n16848;
  assign n16850 = ~controllable_BtoR_REQ1 & ~n16849;
  assign n16851 = controllable_BtoR_REQ0 & ~n16850;
  assign n16852 = ~n15039 & ~n16851;
  assign n16853 = i_RtoB_ACK0 & ~n16852;
  assign n16854 = ~n15141 & ~n16853;
  assign n16855 = ~controllable_DEQ & ~n16854;
  assign n16856 = ~n15127 & ~n16855;
  assign n16857 = i_FULL & ~n16856;
  assign n16858 = ~n15166 & ~n16827;
  assign n16859 = ~controllable_DEQ & ~n16858;
  assign n16860 = ~n15162 & ~n16859;
  assign n16861 = ~i_FULL & ~n16860;
  assign n16862 = ~n16857 & ~n16861;
  assign n16863 = ~i_nEMPTY & ~n16862;
  assign n16864 = ~n16847 & ~n16863;
  assign n16865 = ~controllable_BtoS_ACK0 & ~n16864;
  assign n16866 = ~n16820 & ~n16865;
  assign n16867 = n4465 & ~n16866;
  assign n16868 = ~i_RtoB_ACK1 & ~n13373;
  assign n16869 = ~n7054 & ~n16868;
  assign n16870 = ~controllable_BtoR_REQ1 & ~n16869;
  assign n16871 = ~controllable_BtoR_REQ1 & ~n16870;
  assign n16872 = controllable_BtoR_REQ0 & ~n16871;
  assign n16873 = ~n15183 & ~n16872;
  assign n16874 = i_RtoB_ACK0 & ~n16873;
  assign n16875 = ~n15194 & ~n16874;
  assign n16876 = controllable_DEQ & ~n16875;
  assign n16877 = ~n7111 & ~n9804;
  assign n16878 = ~controllable_BtoR_REQ1 & ~n16877;
  assign n16879 = ~controllable_BtoR_REQ1 & ~n16878;
  assign n16880 = controllable_BtoR_REQ0 & ~n16879;
  assign n16881 = ~n15202 & ~n16880;
  assign n16882 = i_RtoB_ACK0 & ~n16881;
  assign n16883 = ~n15211 & ~n16882;
  assign n16884 = ~controllable_DEQ & ~n16883;
  assign n16885 = ~n16876 & ~n16884;
  assign n16886 = i_nEMPTY & ~n16885;
  assign n16887 = ~n7054 & ~n9781;
  assign n16888 = ~controllable_BtoR_REQ1 & ~n16887;
  assign n16889 = ~controllable_BtoR_REQ1 & ~n16888;
  assign n16890 = controllable_BtoR_REQ0 & ~n16889;
  assign n16891 = ~n15183 & ~n16890;
  assign n16892 = i_RtoB_ACK0 & ~n16891;
  assign n16893 = ~n15239 & ~n16892;
  assign n16894 = ~controllable_DEQ & ~n16893;
  assign n16895 = ~n15227 & ~n16894;
  assign n16896 = i_FULL & ~n16895;
  assign n16897 = ~n15259 & ~n16874;
  assign n16898 = ~controllable_DEQ & ~n16897;
  assign n16899 = ~n15255 & ~n16898;
  assign n16900 = ~i_FULL & ~n16899;
  assign n16901 = ~n16896 & ~n16900;
  assign n16902 = ~i_nEMPTY & ~n16901;
  assign n16903 = ~n16886 & ~n16902;
  assign n16904 = controllable_BtoS_ACK0 & ~n16903;
  assign n16905 = ~i_RtoB_ACK1 & ~n9878;
  assign n16906 = ~n7196 & ~n16905;
  assign n16907 = ~controllable_BtoR_REQ1 & ~n16906;
  assign n16908 = ~controllable_BtoR_REQ1 & ~n16907;
  assign n16909 = controllable_BtoR_REQ0 & ~n16908;
  assign n16910 = ~n15274 & ~n16909;
  assign n16911 = i_RtoB_ACK0 & ~n16910;
  assign n16912 = ~n15285 & ~n16911;
  assign n16913 = controllable_DEQ & ~n16912;
  assign n16914 = ~n7277 & ~n9904;
  assign n16915 = ~controllable_BtoR_REQ1 & ~n16914;
  assign n16916 = ~controllable_BtoR_REQ1 & ~n16915;
  assign n16917 = controllable_BtoR_REQ0 & ~n16916;
  assign n16918 = ~n15293 & ~n16917;
  assign n16919 = i_RtoB_ACK0 & ~n16918;
  assign n16920 = ~n15304 & ~n16919;
  assign n16921 = ~controllable_DEQ & ~n16920;
  assign n16922 = ~n16913 & ~n16921;
  assign n16923 = i_FULL & ~n16922;
  assign n16924 = ~n15323 & ~n16911;
  assign n16925 = controllable_DEQ & ~n16924;
  assign n16926 = ~n15339 & ~n16919;
  assign n16927 = ~controllable_DEQ & ~n16926;
  assign n16928 = ~n16925 & ~n16927;
  assign n16929 = ~i_FULL & ~n16928;
  assign n16930 = ~n16923 & ~n16929;
  assign n16931 = i_nEMPTY & ~n16930;
  assign n16932 = ~n7196 & ~n9871;
  assign n16933 = ~controllable_BtoR_REQ1 & ~n16932;
  assign n16934 = ~controllable_BtoR_REQ1 & ~n16933;
  assign n16935 = controllable_BtoR_REQ0 & ~n16934;
  assign n16936 = ~n15274 & ~n16935;
  assign n16937 = i_RtoB_ACK0 & ~n16936;
  assign n16938 = ~n15376 & ~n16937;
  assign n16939 = ~controllable_DEQ & ~n16938;
  assign n16940 = ~n15362 & ~n16939;
  assign n16941 = i_FULL & ~n16940;
  assign n16942 = ~n15401 & ~n16911;
  assign n16943 = ~controllable_DEQ & ~n16942;
  assign n16944 = ~n15397 & ~n16943;
  assign n16945 = ~i_FULL & ~n16944;
  assign n16946 = ~n16941 & ~n16945;
  assign n16947 = ~i_nEMPTY & ~n16946;
  assign n16948 = ~n16931 & ~n16947;
  assign n16949 = ~controllable_BtoS_ACK0 & ~n16948;
  assign n16950 = ~n16904 & ~n16949;
  assign n16951 = ~n4465 & ~n16950;
  assign n16952 = ~n16867 & ~n16951;
  assign n16953 = ~i_StoB_REQ10 & ~n16952;
  assign n16954 = ~n16775 & ~n16953;
  assign n16955 = controllable_BtoS_ACK10 & ~n16954;
  assign n16956 = ~i_RtoB_ACK1 & ~n10008;
  assign n16957 = ~n7391 & ~n16956;
  assign n16958 = ~controllable_BtoR_REQ1 & ~n16957;
  assign n16959 = ~controllable_BtoR_REQ1 & ~n16958;
  assign n16960 = controllable_BtoR_REQ0 & ~n16959;
  assign n16961 = ~n14897 & ~n16960;
  assign n16962 = i_RtoB_ACK0 & ~n16961;
  assign n16963 = ~n15423 & ~n16962;
  assign n16964 = controllable_DEQ & ~n16963;
  assign n16965 = ~n7410 & ~n9813;
  assign n16966 = ~controllable_BtoR_REQ1 & ~n16965;
  assign n16967 = ~controllable_BtoR_REQ1 & ~n16966;
  assign n16968 = controllable_BtoR_REQ0 & ~n16967;
  assign n16969 = ~n14916 & ~n16968;
  assign n16970 = i_RtoB_ACK0 & ~n16969;
  assign n16971 = ~n15432 & ~n16970;
  assign n16972 = ~controllable_DEQ & ~n16971;
  assign n16973 = ~n16964 & ~n16972;
  assign n16974 = i_FULL & ~n16973;
  assign n16975 = ~n15444 & ~n16962;
  assign n16976 = controllable_DEQ & ~n16975;
  assign n16977 = ~n15453 & ~n16970;
  assign n16978 = ~controllable_DEQ & ~n16977;
  assign n16979 = ~n16976 & ~n16978;
  assign n16980 = ~i_FULL & ~n16979;
  assign n16981 = ~n16974 & ~n16980;
  assign n16982 = i_nEMPTY & ~n16981;
  assign n16983 = ~n7391 & ~n9836;
  assign n16984 = ~controllable_BtoR_REQ1 & ~n16983;
  assign n16985 = ~controllable_BtoR_REQ1 & ~n16984;
  assign n16986 = controllable_BtoR_REQ0 & ~n16985;
  assign n16987 = ~n14897 & ~n16986;
  assign n16988 = i_RtoB_ACK0 & ~n16987;
  assign n16989 = ~n15476 & ~n16988;
  assign n16990 = ~controllable_DEQ & ~n16989;
  assign n16991 = ~n15469 & ~n16990;
  assign n16992 = i_FULL & ~n16991;
  assign n16993 = ~controllable_DEQ & ~n16963;
  assign n16994 = ~n15490 & ~n16993;
  assign n16995 = ~i_FULL & ~n16994;
  assign n16996 = ~n16992 & ~n16995;
  assign n16997 = ~i_nEMPTY & ~n16996;
  assign n16998 = ~n16982 & ~n16997;
  assign n16999 = controllable_BtoS_ACK0 & ~n16998;
  assign n17000 = ~i_RtoB_ACK1 & ~n10081;
  assign n17001 = ~n7471 & ~n17000;
  assign n17002 = ~controllable_BtoR_REQ1 & ~n17001;
  assign n17003 = ~controllable_BtoR_REQ1 & ~n17002;
  assign n17004 = controllable_BtoR_REQ0 & ~n17003;
  assign n17005 = ~n15039 & ~n17004;
  assign n17006 = i_RtoB_ACK0 & ~n17005;
  assign n17007 = ~n15505 & ~n17006;
  assign n17008 = controllable_DEQ & ~n17007;
  assign n17009 = ~n7490 & ~n9904;
  assign n17010 = ~controllable_BtoR_REQ1 & ~n17009;
  assign n17011 = ~controllable_BtoR_REQ1 & ~n17010;
  assign n17012 = controllable_BtoR_REQ0 & ~n17011;
  assign n17013 = ~n15058 & ~n17012;
  assign n17014 = i_RtoB_ACK0 & ~n17013;
  assign n17015 = ~n15514 & ~n17014;
  assign n17016 = ~controllable_DEQ & ~n17015;
  assign n17017 = ~n17008 & ~n17016;
  assign n17018 = i_FULL & ~n17017;
  assign n17019 = ~n15526 & ~n17006;
  assign n17020 = controllable_DEQ & ~n17019;
  assign n17021 = ~n15535 & ~n17014;
  assign n17022 = ~controllable_DEQ & ~n17021;
  assign n17023 = ~n17020 & ~n17022;
  assign n17024 = ~i_FULL & ~n17023;
  assign n17025 = ~n17018 & ~n17024;
  assign n17026 = i_nEMPTY & ~n17025;
  assign n17027 = ~n7471 & ~n9871;
  assign n17028 = ~controllable_BtoR_REQ1 & ~n17027;
  assign n17029 = ~controllable_BtoR_REQ1 & ~n17028;
  assign n17030 = controllable_BtoR_REQ0 & ~n17029;
  assign n17031 = ~n15039 & ~n17030;
  assign n17032 = i_RtoB_ACK0 & ~n17031;
  assign n17033 = ~n15558 & ~n17032;
  assign n17034 = ~controllable_DEQ & ~n17033;
  assign n17035 = ~n15551 & ~n17034;
  assign n17036 = i_FULL & ~n17035;
  assign n17037 = ~controllable_DEQ & ~n17007;
  assign n17038 = ~n15572 & ~n17037;
  assign n17039 = ~i_FULL & ~n17038;
  assign n17040 = ~n17036 & ~n17039;
  assign n17041 = ~i_nEMPTY & ~n17040;
  assign n17042 = ~n17026 & ~n17041;
  assign n17043 = ~controllable_BtoS_ACK0 & ~n17042;
  assign n17044 = ~n16999 & ~n17043;
  assign n17045 = n4465 & ~n17044;
  assign n17046 = ~i_RtoB_ACK1 & ~n10148;
  assign n17047 = ~n5237 & ~n17046;
  assign n17048 = ~controllable_BtoR_REQ1 & ~n17047;
  assign n17049 = ~controllable_BtoR_REQ1 & ~n17048;
  assign n17050 = controllable_BtoR_REQ0 & ~n17049;
  assign n17051 = ~n15183 & ~n17050;
  assign n17052 = i_RtoB_ACK0 & ~n17051;
  assign n17053 = ~n15589 & ~n17052;
  assign n17054 = controllable_DEQ & ~n17053;
  assign n17055 = ~n7563 & ~n9813;
  assign n17056 = ~controllable_BtoR_REQ1 & ~n17055;
  assign n17057 = ~controllable_BtoR_REQ1 & ~n17056;
  assign n17058 = controllable_BtoR_REQ0 & ~n17057;
  assign n17059 = ~n15202 & ~n17058;
  assign n17060 = i_RtoB_ACK0 & ~n17059;
  assign n17061 = ~n15597 & ~n17060;
  assign n17062 = ~controllable_DEQ & ~n17061;
  assign n17063 = ~n17054 & ~n17062;
  assign n17064 = i_nEMPTY & ~n17063;
  assign n17065 = ~n5237 & ~n9836;
  assign n17066 = ~controllable_BtoR_REQ1 & ~n17065;
  assign n17067 = ~controllable_BtoR_REQ1 & ~n17066;
  assign n17068 = controllable_BtoR_REQ0 & ~n17067;
  assign n17069 = ~n15183 & ~n17068;
  assign n17070 = i_RtoB_ACK0 & ~n17069;
  assign n17071 = ~n15613 & ~n17070;
  assign n17072 = ~controllable_DEQ & ~n17071;
  assign n17073 = ~n15607 & ~n17072;
  assign n17074 = i_FULL & ~n17073;
  assign n17075 = ~controllable_DEQ & ~n17053;
  assign n17076 = ~n15622 & ~n17075;
  assign n17077 = ~i_FULL & ~n17076;
  assign n17078 = ~n17074 & ~n17077;
  assign n17079 = ~i_nEMPTY & ~n17078;
  assign n17080 = ~n17064 & ~n17079;
  assign n17081 = controllable_BtoS_ACK0 & ~n17080;
  assign n17082 = ~i_RtoB_ACK1 & ~n10195;
  assign n17083 = ~n7607 & ~n17082;
  assign n17084 = ~controllable_BtoR_REQ1 & ~n17083;
  assign n17085 = ~controllable_BtoR_REQ1 & ~n17084;
  assign n17086 = controllable_BtoR_REQ0 & ~n17085;
  assign n17087 = ~n15274 & ~n17086;
  assign n17088 = i_RtoB_ACK0 & ~n17087;
  assign n17089 = ~n15637 & ~n17088;
  assign n17090 = controllable_DEQ & ~n17089;
  assign n17091 = ~n7626 & ~n9904;
  assign n17092 = ~controllable_BtoR_REQ1 & ~n17091;
  assign n17093 = ~controllable_BtoR_REQ1 & ~n17092;
  assign n17094 = controllable_BtoR_REQ0 & ~n17093;
  assign n17095 = ~n15293 & ~n17094;
  assign n17096 = i_RtoB_ACK0 & ~n17095;
  assign n17097 = ~n15646 & ~n17096;
  assign n17098 = ~controllable_DEQ & ~n17097;
  assign n17099 = ~n17090 & ~n17098;
  assign n17100 = i_FULL & ~n17099;
  assign n17101 = ~n15658 & ~n17088;
  assign n17102 = controllable_DEQ & ~n17101;
  assign n17103 = ~n15667 & ~n17096;
  assign n17104 = ~controllable_DEQ & ~n17103;
  assign n17105 = ~n17102 & ~n17104;
  assign n17106 = ~i_FULL & ~n17105;
  assign n17107 = ~n17100 & ~n17106;
  assign n17108 = i_nEMPTY & ~n17107;
  assign n17109 = ~n7607 & ~n9871;
  assign n17110 = ~controllable_BtoR_REQ1 & ~n17109;
  assign n17111 = ~controllable_BtoR_REQ1 & ~n17110;
  assign n17112 = controllable_BtoR_REQ0 & ~n17111;
  assign n17113 = ~n15274 & ~n17112;
  assign n17114 = i_RtoB_ACK0 & ~n17113;
  assign n17115 = ~n15690 & ~n17114;
  assign n17116 = ~controllable_DEQ & ~n17115;
  assign n17117 = ~n15683 & ~n17116;
  assign n17118 = i_FULL & ~n17117;
  assign n17119 = ~controllable_DEQ & ~n17089;
  assign n17120 = ~n15704 & ~n17119;
  assign n17121 = ~i_FULL & ~n17120;
  assign n17122 = ~n17118 & ~n17121;
  assign n17123 = ~i_nEMPTY & ~n17122;
  assign n17124 = ~n17108 & ~n17123;
  assign n17125 = ~controllable_BtoS_ACK0 & ~n17124;
  assign n17126 = ~n17081 & ~n17125;
  assign n17127 = ~n4465 & ~n17126;
  assign n17128 = ~n17045 & ~n17127;
  assign n17129 = i_StoB_REQ10 & ~n17128;
  assign n17130 = ~n16953 & ~n17129;
  assign n17131 = ~controllable_BtoS_ACK10 & ~n17130;
  assign n17132 = ~n16955 & ~n17131;
  assign n17133 = n4464 & ~n17132;
  assign n17134 = ~n14741 & ~n15725;
  assign n17135 = i_RtoB_ACK0 & ~n17134;
  assign n17136 = ~n15736 & ~n17135;
  assign n17137 = controllable_DEQ & ~n17136;
  assign n17138 = ~n14757 & ~n15742;
  assign n17139 = i_RtoB_ACK0 & ~n17138;
  assign n17140 = ~n15751 & ~n17139;
  assign n17141 = ~controllable_DEQ & ~n17140;
  assign n17142 = ~n17137 & ~n17141;
  assign n17143 = i_nEMPTY & ~n17142;
  assign n17144 = ~n15770 & ~n17135;
  assign n17145 = ~controllable_DEQ & ~n17144;
  assign n17146 = ~n15764 & ~n17145;
  assign n17147 = i_FULL & ~n17146;
  assign n17148 = ~n15786 & ~n17135;
  assign n17149 = ~controllable_DEQ & ~n17148;
  assign n17150 = ~n15782 & ~n17149;
  assign n17151 = ~i_FULL & ~n17150;
  assign n17152 = ~n17147 & ~n17151;
  assign n17153 = ~i_nEMPTY & ~n17152;
  assign n17154 = ~n17143 & ~n17153;
  assign n17155 = controllable_BtoS_ACK0 & ~n17154;
  assign n17156 = ~n15800 & ~n16723;
  assign n17157 = i_RtoB_ACK0 & ~n17156;
  assign n17158 = ~n15811 & ~n17157;
  assign n17159 = controllable_DEQ & ~n17158;
  assign n17160 = ~n15817 & ~n16729;
  assign n17161 = i_RtoB_ACK0 & ~n17160;
  assign n17162 = ~n15826 & ~n17161;
  assign n17163 = ~controllable_DEQ & ~n17162;
  assign n17164 = ~n17159 & ~n17163;
  assign n17165 = i_nEMPTY & ~n17164;
  assign n17166 = ~n15845 & ~n17157;
  assign n17167 = ~controllable_DEQ & ~n17166;
  assign n17168 = ~n15839 & ~n17167;
  assign n17169 = i_FULL & ~n17168;
  assign n17170 = ~n15861 & ~n17157;
  assign n17171 = ~controllable_DEQ & ~n17170;
  assign n17172 = ~n15857 & ~n17171;
  assign n17173 = ~i_FULL & ~n17172;
  assign n17174 = ~n17169 & ~n17173;
  assign n17175 = ~i_nEMPTY & ~n17174;
  assign n17176 = ~n17165 & ~n17175;
  assign n17177 = ~controllable_BtoS_ACK0 & ~n17176;
  assign n17178 = ~n17155 & ~n17177;
  assign n17179 = n4465 & ~n17178;
  assign n17180 = ~n14811 & ~n17177;
  assign n17181 = ~n4465 & ~n17180;
  assign n17182 = ~n17179 & ~n17181;
  assign n17183 = i_StoB_REQ10 & ~n17182;
  assign n17184 = ~i_RtoB_ACK1 & ~n13695;
  assign n17185 = ~n7886 & ~n17184;
  assign n17186 = ~controllable_BtoR_REQ1 & ~n17185;
  assign n17187 = ~controllable_BtoR_REQ1 & ~n17186;
  assign n17188 = controllable_BtoR_REQ0 & ~n17187;
  assign n17189 = ~n15882 & ~n17188;
  assign n17190 = i_RtoB_ACK0 & ~n17189;
  assign n17191 = ~n15893 & ~n17190;
  assign n17192 = controllable_DEQ & ~n17191;
  assign n17193 = ~n7947 & ~n10487;
  assign n17194 = ~controllable_BtoR_REQ1 & ~n17193;
  assign n17195 = ~controllable_BtoR_REQ1 & ~n17194;
  assign n17196 = controllable_BtoR_REQ0 & ~n17195;
  assign n17197 = ~n15901 & ~n17196;
  assign n17198 = i_RtoB_ACK0 & ~n17197;
  assign n17199 = ~n15912 & ~n17198;
  assign n17200 = ~controllable_DEQ & ~n17199;
  assign n17201 = ~n17192 & ~n17200;
  assign n17202 = i_FULL & ~n17201;
  assign n17203 = ~n15931 & ~n17190;
  assign n17204 = controllable_DEQ & ~n17203;
  assign n17205 = ~n15947 & ~n17198;
  assign n17206 = ~controllable_DEQ & ~n17205;
  assign n17207 = ~n17204 & ~n17206;
  assign n17208 = ~i_FULL & ~n17207;
  assign n17209 = ~n17202 & ~n17208;
  assign n17210 = i_nEMPTY & ~n17209;
  assign n17211 = ~n7886 & ~n10460;
  assign n17212 = ~controllable_BtoR_REQ1 & ~n17211;
  assign n17213 = ~controllable_BtoR_REQ1 & ~n17212;
  assign n17214 = controllable_BtoR_REQ0 & ~n17213;
  assign n17215 = ~n15882 & ~n17214;
  assign n17216 = i_RtoB_ACK0 & ~n17215;
  assign n17217 = ~n15984 & ~n17216;
  assign n17218 = ~controllable_DEQ & ~n17217;
  assign n17219 = ~n15970 & ~n17218;
  assign n17220 = i_FULL & ~n17219;
  assign n17221 = ~n16009 & ~n17190;
  assign n17222 = ~controllable_DEQ & ~n17221;
  assign n17223 = ~n16005 & ~n17222;
  assign n17224 = ~i_FULL & ~n17223;
  assign n17225 = ~n17220 & ~n17224;
  assign n17226 = ~i_nEMPTY & ~n17225;
  assign n17227 = ~n17210 & ~n17226;
  assign n17228 = controllable_BtoS_ACK0 & ~n17227;
  assign n17229 = ~i_RtoB_ACK1 & ~n13759;
  assign n17230 = ~n8057 & ~n17229;
  assign n17231 = ~controllable_BtoR_REQ1 & ~n17230;
  assign n17232 = ~controllable_BtoR_REQ1 & ~n17231;
  assign n17233 = controllable_BtoR_REQ0 & ~n17232;
  assign n17234 = ~n16024 & ~n17233;
  assign n17235 = i_RtoB_ACK0 & ~n17234;
  assign n17236 = ~n16035 & ~n17235;
  assign n17237 = controllable_DEQ & ~n17236;
  assign n17238 = ~n8111 & ~n10614;
  assign n17239 = ~controllable_BtoR_REQ1 & ~n17238;
  assign n17240 = ~controllable_BtoR_REQ1 & ~n17239;
  assign n17241 = controllable_BtoR_REQ0 & ~n17240;
  assign n17242 = ~n16043 & ~n17241;
  assign n17243 = i_RtoB_ACK0 & ~n17242;
  assign n17244 = ~n16054 & ~n17243;
  assign n17245 = ~controllable_DEQ & ~n17244;
  assign n17246 = ~n17237 & ~n17245;
  assign n17247 = i_FULL & ~n17246;
  assign n17248 = ~n16073 & ~n17235;
  assign n17249 = controllable_DEQ & ~n17248;
  assign n17250 = ~n16089 & ~n17243;
  assign n17251 = ~controllable_DEQ & ~n17250;
  assign n17252 = ~n17249 & ~n17251;
  assign n17253 = ~i_FULL & ~n17252;
  assign n17254 = ~n17247 & ~n17253;
  assign n17255 = i_nEMPTY & ~n17254;
  assign n17256 = ~n8057 & ~n10590;
  assign n17257 = ~controllable_BtoR_REQ1 & ~n17256;
  assign n17258 = ~controllable_BtoR_REQ1 & ~n17257;
  assign n17259 = controllable_BtoR_REQ0 & ~n17258;
  assign n17260 = ~n16024 & ~n17259;
  assign n17261 = i_RtoB_ACK0 & ~n17260;
  assign n17262 = ~n16126 & ~n17261;
  assign n17263 = ~controllable_DEQ & ~n17262;
  assign n17264 = ~n16112 & ~n17263;
  assign n17265 = i_FULL & ~n17264;
  assign n17266 = ~n16151 & ~n17235;
  assign n17267 = ~controllable_DEQ & ~n17266;
  assign n17268 = ~n16147 & ~n17267;
  assign n17269 = ~i_FULL & ~n17268;
  assign n17270 = ~n17265 & ~n17269;
  assign n17271 = ~i_nEMPTY & ~n17270;
  assign n17272 = ~n17255 & ~n17271;
  assign n17273 = ~controllable_BtoS_ACK0 & ~n17272;
  assign n17274 = ~n17228 & ~n17273;
  assign n17275 = n4465 & ~n17274;
  assign n17276 = ~i_RtoB_ACK1 & ~n9788;
  assign n17277 = ~n7054 & ~n17276;
  assign n17278 = ~controllable_BtoR_REQ1 & ~n17277;
  assign n17279 = ~controllable_BtoR_REQ1 & ~n17278;
  assign n17280 = controllable_BtoR_REQ0 & ~n17279;
  assign n17281 = ~n16168 & ~n17280;
  assign n17282 = i_RtoB_ACK0 & ~n17281;
  assign n17283 = ~n16179 & ~n17282;
  assign n17284 = controllable_DEQ & ~n17283;
  assign n17285 = ~n7111 & ~n9813;
  assign n17286 = ~controllable_BtoR_REQ1 & ~n17285;
  assign n17287 = ~controllable_BtoR_REQ1 & ~n17286;
  assign n17288 = controllable_BtoR_REQ0 & ~n17287;
  assign n17289 = ~n16187 & ~n17288;
  assign n17290 = i_RtoB_ACK0 & ~n17289;
  assign n17291 = ~n16196 & ~n17290;
  assign n17292 = ~controllable_DEQ & ~n17291;
  assign n17293 = ~n17284 & ~n17292;
  assign n17294 = i_nEMPTY & ~n17293;
  assign n17295 = ~n7054 & ~n9836;
  assign n17296 = ~controllable_BtoR_REQ1 & ~n17295;
  assign n17297 = ~controllable_BtoR_REQ1 & ~n17296;
  assign n17298 = controllable_BtoR_REQ0 & ~n17297;
  assign n17299 = ~n16168 & ~n17298;
  assign n17300 = i_RtoB_ACK0 & ~n17299;
  assign n17301 = ~n16222 & ~n17300;
  assign n17302 = ~controllable_DEQ & ~n17301;
  assign n17303 = ~n16210 & ~n17302;
  assign n17304 = i_FULL & ~n17303;
  assign n17305 = ~n16240 & ~n17282;
  assign n17306 = ~controllable_DEQ & ~n17305;
  assign n17307 = ~n16236 & ~n17306;
  assign n17308 = ~i_FULL & ~n17307;
  assign n17309 = ~n17304 & ~n17308;
  assign n17310 = ~i_nEMPTY & ~n17309;
  assign n17311 = ~n17294 & ~n17310;
  assign n17312 = controllable_BtoS_ACK0 & ~n17311;
  assign n17313 = ~i_RtoB_ACK1 & ~n10787;
  assign n17314 = ~n8313 & ~n17313;
  assign n17315 = ~controllable_BtoR_REQ1 & ~n17314;
  assign n17316 = ~controllable_BtoR_REQ1 & ~n17315;
  assign n17317 = controllable_BtoR_REQ0 & ~n17316;
  assign n17318 = ~n16255 & ~n17317;
  assign n17319 = i_RtoB_ACK0 & ~n17318;
  assign n17320 = ~n16266 & ~n17319;
  assign n17321 = controllable_DEQ & ~n17320;
  assign n17322 = ~n8352 & ~n9904;
  assign n17323 = ~controllable_BtoR_REQ1 & ~n17322;
  assign n17324 = ~controllable_BtoR_REQ1 & ~n17323;
  assign n17325 = controllable_BtoR_REQ0 & ~n17324;
  assign n17326 = ~n16274 & ~n17325;
  assign n17327 = i_RtoB_ACK0 & ~n17326;
  assign n17328 = ~n16285 & ~n17327;
  assign n17329 = ~controllable_DEQ & ~n17328;
  assign n17330 = ~n17321 & ~n17329;
  assign n17331 = i_FULL & ~n17330;
  assign n17332 = ~n16304 & ~n17319;
  assign n17333 = controllable_DEQ & ~n17332;
  assign n17334 = ~n16320 & ~n17327;
  assign n17335 = ~controllable_DEQ & ~n17334;
  assign n17336 = ~n17333 & ~n17335;
  assign n17337 = ~i_FULL & ~n17336;
  assign n17338 = ~n17331 & ~n17337;
  assign n17339 = i_nEMPTY & ~n17338;
  assign n17340 = ~n8313 & ~n9871;
  assign n17341 = ~controllable_BtoR_REQ1 & ~n17340;
  assign n17342 = ~controllable_BtoR_REQ1 & ~n17341;
  assign n17343 = controllable_BtoR_REQ0 & ~n17342;
  assign n17344 = ~n16255 & ~n17343;
  assign n17345 = i_RtoB_ACK0 & ~n17344;
  assign n17346 = ~n16357 & ~n17345;
  assign n17347 = ~controllable_DEQ & ~n17346;
  assign n17348 = ~n16343 & ~n17347;
  assign n17349 = i_FULL & ~n17348;
  assign n17350 = ~n16382 & ~n17319;
  assign n17351 = ~controllable_DEQ & ~n17350;
  assign n17352 = ~n16378 & ~n17351;
  assign n17353 = ~i_FULL & ~n17352;
  assign n17354 = ~n17349 & ~n17353;
  assign n17355 = ~i_nEMPTY & ~n17354;
  assign n17356 = ~n17339 & ~n17355;
  assign n17357 = ~controllable_BtoS_ACK0 & ~n17356;
  assign n17358 = ~n17312 & ~n17357;
  assign n17359 = ~n4465 & ~n17358;
  assign n17360 = ~n17275 & ~n17359;
  assign n17361 = ~i_StoB_REQ10 & ~n17360;
  assign n17362 = ~n17183 & ~n17361;
  assign n17363 = controllable_BtoS_ACK10 & ~n17362;
  assign n17364 = ~i_RtoB_ACK1 & ~n10887;
  assign n17365 = ~n8461 & ~n17364;
  assign n17366 = ~controllable_BtoR_REQ1 & ~n17365;
  assign n17367 = ~controllable_BtoR_REQ1 & ~n17366;
  assign n17368 = controllable_BtoR_REQ0 & ~n17367;
  assign n17369 = ~n15882 & ~n17368;
  assign n17370 = i_RtoB_ACK0 & ~n17369;
  assign n17371 = ~n16404 & ~n17370;
  assign n17372 = controllable_DEQ & ~n17371;
  assign n17373 = ~n8480 & ~n9813;
  assign n17374 = ~controllable_BtoR_REQ1 & ~n17373;
  assign n17375 = ~controllable_BtoR_REQ1 & ~n17374;
  assign n17376 = controllable_BtoR_REQ0 & ~n17375;
  assign n17377 = ~n15901 & ~n17376;
  assign n17378 = i_RtoB_ACK0 & ~n17377;
  assign n17379 = ~n16413 & ~n17378;
  assign n17380 = ~controllable_DEQ & ~n17379;
  assign n17381 = ~n17372 & ~n17380;
  assign n17382 = i_FULL & ~n17381;
  assign n17383 = ~n16425 & ~n17370;
  assign n17384 = controllable_DEQ & ~n17383;
  assign n17385 = ~n16434 & ~n17378;
  assign n17386 = ~controllable_DEQ & ~n17385;
  assign n17387 = ~n17384 & ~n17386;
  assign n17388 = ~i_FULL & ~n17387;
  assign n17389 = ~n17382 & ~n17388;
  assign n17390 = i_nEMPTY & ~n17389;
  assign n17391 = ~n8461 & ~n9836;
  assign n17392 = ~controllable_BtoR_REQ1 & ~n17391;
  assign n17393 = ~controllable_BtoR_REQ1 & ~n17392;
  assign n17394 = controllable_BtoR_REQ0 & ~n17393;
  assign n17395 = ~n15882 & ~n17394;
  assign n17396 = i_RtoB_ACK0 & ~n17395;
  assign n17397 = ~n16457 & ~n17396;
  assign n17398 = ~controllable_DEQ & ~n17397;
  assign n17399 = ~n16450 & ~n17398;
  assign n17400 = i_FULL & ~n17399;
  assign n17401 = ~controllable_DEQ & ~n17371;
  assign n17402 = ~n16471 & ~n17401;
  assign n17403 = ~i_FULL & ~n17402;
  assign n17404 = ~n17400 & ~n17403;
  assign n17405 = ~i_nEMPTY & ~n17404;
  assign n17406 = ~n17390 & ~n17405;
  assign n17407 = controllable_BtoS_ACK0 & ~n17406;
  assign n17408 = ~i_RtoB_ACK1 & ~n10954;
  assign n17409 = ~n8540 & ~n17408;
  assign n17410 = ~controllable_BtoR_REQ1 & ~n17409;
  assign n17411 = ~controllable_BtoR_REQ1 & ~n17410;
  assign n17412 = controllable_BtoR_REQ0 & ~n17411;
  assign n17413 = ~n16024 & ~n17412;
  assign n17414 = i_RtoB_ACK0 & ~n17413;
  assign n17415 = ~n16486 & ~n17414;
  assign n17416 = controllable_DEQ & ~n17415;
  assign n17417 = ~n8559 & ~n9904;
  assign n17418 = ~controllable_BtoR_REQ1 & ~n17417;
  assign n17419 = ~controllable_BtoR_REQ1 & ~n17418;
  assign n17420 = controllable_BtoR_REQ0 & ~n17419;
  assign n17421 = ~n16043 & ~n17420;
  assign n17422 = i_RtoB_ACK0 & ~n17421;
  assign n17423 = ~n16495 & ~n17422;
  assign n17424 = ~controllable_DEQ & ~n17423;
  assign n17425 = ~n17416 & ~n17424;
  assign n17426 = i_FULL & ~n17425;
  assign n17427 = ~n16507 & ~n17414;
  assign n17428 = controllable_DEQ & ~n17427;
  assign n17429 = ~n16516 & ~n17422;
  assign n17430 = ~controllable_DEQ & ~n17429;
  assign n17431 = ~n17428 & ~n17430;
  assign n17432 = ~i_FULL & ~n17431;
  assign n17433 = ~n17426 & ~n17432;
  assign n17434 = i_nEMPTY & ~n17433;
  assign n17435 = ~n8540 & ~n9871;
  assign n17436 = ~controllable_BtoR_REQ1 & ~n17435;
  assign n17437 = ~controllable_BtoR_REQ1 & ~n17436;
  assign n17438 = controllable_BtoR_REQ0 & ~n17437;
  assign n17439 = ~n16024 & ~n17438;
  assign n17440 = i_RtoB_ACK0 & ~n17439;
  assign n17441 = ~n16539 & ~n17440;
  assign n17442 = ~controllable_DEQ & ~n17441;
  assign n17443 = ~n16532 & ~n17442;
  assign n17444 = i_FULL & ~n17443;
  assign n17445 = ~controllable_DEQ & ~n17415;
  assign n17446 = ~n16553 & ~n17445;
  assign n17447 = ~i_FULL & ~n17446;
  assign n17448 = ~n17444 & ~n17447;
  assign n17449 = ~i_nEMPTY & ~n17448;
  assign n17450 = ~n17434 & ~n17449;
  assign n17451 = ~controllable_BtoS_ACK0 & ~n17450;
  assign n17452 = ~n17407 & ~n17451;
  assign n17453 = n4465 & ~n17452;
  assign n17454 = ~n16168 & ~n17050;
  assign n17455 = i_RtoB_ACK0 & ~n17454;
  assign n17456 = ~n16570 & ~n17455;
  assign n17457 = controllable_DEQ & ~n17456;
  assign n17458 = ~n16187 & ~n17058;
  assign n17459 = i_RtoB_ACK0 & ~n17458;
  assign n17460 = ~n16578 & ~n17459;
  assign n17461 = ~controllable_DEQ & ~n17460;
  assign n17462 = ~n17457 & ~n17461;
  assign n17463 = i_nEMPTY & ~n17462;
  assign n17464 = ~n16168 & ~n17068;
  assign n17465 = i_RtoB_ACK0 & ~n17464;
  assign n17466 = ~n16591 & ~n17465;
  assign n17467 = ~controllable_DEQ & ~n17466;
  assign n17468 = ~n16585 & ~n17467;
  assign n17469 = i_FULL & ~n17468;
  assign n17470 = ~controllable_DEQ & ~n17456;
  assign n17471 = ~n16598 & ~n17470;
  assign n17472 = ~i_FULL & ~n17471;
  assign n17473 = ~n17469 & ~n17472;
  assign n17474 = ~i_nEMPTY & ~n17473;
  assign n17475 = ~n17463 & ~n17474;
  assign n17476 = controllable_BtoS_ACK0 & ~n17475;
  assign n17477 = ~i_RtoB_ACK1 & ~n11064;
  assign n17478 = ~n8672 & ~n17477;
  assign n17479 = ~controllable_BtoR_REQ1 & ~n17478;
  assign n17480 = ~controllable_BtoR_REQ1 & ~n17479;
  assign n17481 = controllable_BtoR_REQ0 & ~n17480;
  assign n17482 = ~n16255 & ~n17481;
  assign n17483 = i_RtoB_ACK0 & ~n17482;
  assign n17484 = ~n16613 & ~n17483;
  assign n17485 = controllable_DEQ & ~n17484;
  assign n17486 = ~n8691 & ~n9904;
  assign n17487 = ~controllable_BtoR_REQ1 & ~n17486;
  assign n17488 = ~controllable_BtoR_REQ1 & ~n17487;
  assign n17489 = controllable_BtoR_REQ0 & ~n17488;
  assign n17490 = ~n16274 & ~n17489;
  assign n17491 = i_RtoB_ACK0 & ~n17490;
  assign n17492 = ~n16622 & ~n17491;
  assign n17493 = ~controllable_DEQ & ~n17492;
  assign n17494 = ~n17485 & ~n17493;
  assign n17495 = i_FULL & ~n17494;
  assign n17496 = ~n16634 & ~n17483;
  assign n17497 = controllable_DEQ & ~n17496;
  assign n17498 = ~n16643 & ~n17491;
  assign n17499 = ~controllable_DEQ & ~n17498;
  assign n17500 = ~n17497 & ~n17499;
  assign n17501 = ~i_FULL & ~n17500;
  assign n17502 = ~n17495 & ~n17501;
  assign n17503 = i_nEMPTY & ~n17502;
  assign n17504 = ~n8672 & ~n9871;
  assign n17505 = ~controllable_BtoR_REQ1 & ~n17504;
  assign n17506 = ~controllable_BtoR_REQ1 & ~n17505;
  assign n17507 = controllable_BtoR_REQ0 & ~n17506;
  assign n17508 = ~n16255 & ~n17507;
  assign n17509 = i_RtoB_ACK0 & ~n17508;
  assign n17510 = ~n16666 & ~n17509;
  assign n17511 = ~controllable_DEQ & ~n17510;
  assign n17512 = ~n16659 & ~n17511;
  assign n17513 = i_FULL & ~n17512;
  assign n17514 = ~controllable_DEQ & ~n17484;
  assign n17515 = ~n16680 & ~n17514;
  assign n17516 = ~i_FULL & ~n17515;
  assign n17517 = ~n17513 & ~n17516;
  assign n17518 = ~i_nEMPTY & ~n17517;
  assign n17519 = ~n17503 & ~n17518;
  assign n17520 = ~controllable_BtoS_ACK0 & ~n17519;
  assign n17521 = ~n17476 & ~n17520;
  assign n17522 = ~n4465 & ~n17521;
  assign n17523 = ~n17453 & ~n17522;
  assign n17524 = i_StoB_REQ10 & ~n17523;
  assign n17525 = ~n17361 & ~n17524;
  assign n17526 = ~controllable_BtoS_ACK10 & ~n17525;
  assign n17527 = ~n17363 & ~n17526;
  assign n17528 = ~n4464 & ~n17527;
  assign n17529 = ~n17133 & ~n17528;
  assign n17530 = ~n4463 & ~n17529;
  assign n17531 = ~n16697 & ~n17530;
  assign n17532 = n4462 & ~n17531;
  assign n17533 = ~i_RtoB_ACK1 & ~n12214;
  assign n17534 = ~controllable_BtoR_REQ1 & ~n17533;
  assign n17535 = ~controllable_BtoR_REQ1 & ~n17534;
  assign n17536 = controllable_BtoR_REQ0 & ~n17535;
  assign n17537 = ~controllable_BtoR_REQ1 & ~n11145;
  assign n17538 = ~controllable_BtoR_REQ0 & ~n17537;
  assign n17539 = ~n17536 & ~n17538;
  assign n17540 = i_RtoB_ACK0 & ~n17539;
  assign n17541 = i_RtoB_ACK1 & ~n11135;
  assign n17542 = ~n11153 & ~n17541;
  assign n17543 = ~controllable_BtoR_REQ1 & ~n17542;
  assign n17544 = ~controllable_BtoR_REQ1 & ~n17543;
  assign n17545 = controllable_BtoR_REQ0 & ~n17544;
  assign n17546 = ~controllable_BtoR_REQ1 & ~n11158;
  assign n17547 = ~controllable_BtoR_REQ0 & ~n17546;
  assign n17548 = ~n17545 & ~n17547;
  assign n17549 = ~i_RtoB_ACK0 & ~n17548;
  assign n17550 = ~n17540 & ~n17549;
  assign n17551 = controllable_DEQ & ~n17550;
  assign n17552 = ~controllable_BtoR_REQ1 & ~n11203;
  assign n17553 = controllable_BtoR_REQ0 & ~n17552;
  assign n17554 = ~controllable_BtoR_REQ1 & ~n11168;
  assign n17555 = ~controllable_BtoR_REQ0 & ~n17554;
  assign n17556 = ~n17553 & ~n17555;
  assign n17557 = i_RtoB_ACK0 & ~n17556;
  assign n17558 = i_RtoB_ACK1 & ~n11133;
  assign n17559 = ~n11156 & ~n17558;
  assign n17560 = ~controllable_BtoR_REQ1 & ~n17559;
  assign n17561 = ~controllable_BtoR_REQ1 & ~n17560;
  assign n17562 = controllable_BtoR_REQ0 & ~n17561;
  assign n17563 = ~n17555 & ~n17562;
  assign n17564 = ~i_RtoB_ACK0 & ~n17563;
  assign n17565 = ~n17557 & ~n17564;
  assign n17566 = ~controllable_DEQ & ~n17565;
  assign n17567 = ~n17551 & ~n17566;
  assign n17568 = i_nEMPTY & ~n17567;
  assign n17569 = ~controllable_BtoR_REQ1 & ~n11182;
  assign n17570 = ~controllable_BtoR_REQ1 & ~n17569;
  assign n17571 = controllable_BtoR_REQ0 & ~n17570;
  assign n17572 = ~controllable_BtoR_REQ1 & ~n11188;
  assign n17573 = ~controllable_BtoR_REQ0 & ~n17572;
  assign n17574 = ~n17571 & ~n17573;
  assign n17575 = ~i_RtoB_ACK0 & ~n17574;
  assign n17576 = ~i_RtoB_ACK0 & ~n17575;
  assign n17577 = controllable_DEQ & ~n17576;
  assign n17578 = ~n12214 & ~n17541;
  assign n17579 = ~controllable_BtoR_REQ1 & ~n17578;
  assign n17580 = ~controllable_BtoR_REQ1 & ~n17579;
  assign n17581 = controllable_BtoR_REQ0 & ~n17580;
  assign n17582 = ~n17538 & ~n17581;
  assign n17583 = ~i_RtoB_ACK0 & ~n17582;
  assign n17584 = ~n17540 & ~n17583;
  assign n17585 = ~controllable_DEQ & ~n17584;
  assign n17586 = ~n17577 & ~n17585;
  assign n17587 = i_FULL & ~n17586;
  assign n17588 = ~controllable_BtoR_REQ1 & ~n11166;
  assign n17589 = ~controllable_BtoR_REQ1 & ~n17588;
  assign n17590 = controllable_BtoR_REQ0 & ~n17589;
  assign n17591 = ~controllable_BtoR_REQ0 & ~n17552;
  assign n17592 = ~n17590 & ~n17591;
  assign n17593 = ~i_RtoB_ACK0 & ~n17592;
  assign n17594 = ~i_RtoB_ACK0 & ~n17593;
  assign n17595 = controllable_DEQ & ~n17594;
  assign n17596 = ~controllable_BtoR_REQ1 & ~n14103;
  assign n17597 = ~controllable_BtoR_REQ0 & ~n17596;
  assign n17598 = ~n17545 & ~n17597;
  assign n17599 = ~i_RtoB_ACK0 & ~n17598;
  assign n17600 = ~n17540 & ~n17599;
  assign n17601 = ~controllable_DEQ & ~n17600;
  assign n17602 = ~n17595 & ~n17601;
  assign n17603 = ~i_FULL & ~n17602;
  assign n17604 = ~n17587 & ~n17603;
  assign n17605 = ~i_nEMPTY & ~n17604;
  assign n17606 = ~n17568 & ~n17605;
  assign n17607 = controllable_BtoS_ACK0 & ~n17606;
  assign n17608 = ~n14886 & ~n17607;
  assign n17609 = n4465 & ~n17608;
  assign n17610 = ~n14888 & ~n17609;
  assign n17611 = i_StoB_REQ10 & ~n17610;
  assign n17612 = ~controllable_BtoR_REQ1 & ~n11230;
  assign n17613 = ~controllable_BtoR_REQ0 & ~n17612;
  assign n17614 = ~n17280 & ~n17613;
  assign n17615 = i_RtoB_ACK0 & ~n17614;
  assign n17616 = i_RtoB_ACK1 & ~n11226;
  assign n17617 = ~n9856 & ~n17616;
  assign n17618 = ~controllable_BtoR_REQ1 & ~n17617;
  assign n17619 = ~controllable_BtoR_REQ1 & ~n17618;
  assign n17620 = controllable_BtoR_REQ0 & ~n17619;
  assign n17621 = ~controllable_BtoR_REQ1 & ~n11238;
  assign n17622 = ~controllable_BtoR_REQ0 & ~n17621;
  assign n17623 = ~n17620 & ~n17622;
  assign n17624 = ~i_RtoB_ACK0 & ~n17623;
  assign n17625 = ~n17615 & ~n17624;
  assign n17626 = controllable_DEQ & ~n17625;
  assign n17627 = ~controllable_BtoR_REQ1 & ~n11248;
  assign n17628 = ~controllable_BtoR_REQ0 & ~n17627;
  assign n17629 = ~n17288 & ~n17628;
  assign n17630 = i_RtoB_ACK0 & ~n17629;
  assign n17631 = i_RtoB_ACK1 & ~n9596;
  assign n17632 = ~n9813 & ~n17631;
  assign n17633 = ~controllable_BtoR_REQ1 & ~n17632;
  assign n17634 = ~controllable_BtoR_REQ1 & ~n17633;
  assign n17635 = controllable_BtoR_REQ0 & ~n17634;
  assign n17636 = ~n17628 & ~n17635;
  assign n17637 = ~i_RtoB_ACK0 & ~n17636;
  assign n17638 = ~n17630 & ~n17637;
  assign n17639 = ~controllable_DEQ & ~n17638;
  assign n17640 = ~n17626 & ~n17639;
  assign n17641 = i_nEMPTY & ~n17640;
  assign n17642 = ~i_RtoB_ACK1 & ~n11261;
  assign n17643 = ~controllable_BtoR_REQ1 & ~n17642;
  assign n17644 = ~controllable_BtoR_REQ1 & ~n17643;
  assign n17645 = controllable_BtoR_REQ0 & ~n17644;
  assign n17646 = ~controllable_BtoR_REQ1 & ~n10049;
  assign n17647 = ~controllable_BtoR_REQ0 & ~n17646;
  assign n17648 = ~n17645 & ~n17647;
  assign n17649 = ~i_RtoB_ACK0 & ~n17648;
  assign n17650 = ~n15217 & ~n17649;
  assign n17651 = controllable_DEQ & ~n17650;
  assign n17652 = ~n17298 & ~n17613;
  assign n17653 = i_RtoB_ACK0 & ~n17652;
  assign n17654 = ~n9836 & ~n17616;
  assign n17655 = ~controllable_BtoR_REQ1 & ~n17654;
  assign n17656 = ~controllable_BtoR_REQ1 & ~n17655;
  assign n17657 = controllable_BtoR_REQ0 & ~n17656;
  assign n17658 = ~n17613 & ~n17657;
  assign n17659 = ~i_RtoB_ACK0 & ~n17658;
  assign n17660 = ~n17653 & ~n17659;
  assign n17661 = ~controllable_DEQ & ~n17660;
  assign n17662 = ~n17651 & ~n17661;
  assign n17663 = i_FULL & ~n17662;
  assign n17664 = ~i_RtoB_ACK1 & ~n11245;
  assign n17665 = ~controllable_BtoR_REQ1 & ~n17664;
  assign n17666 = ~controllable_BtoR_REQ1 & ~n17665;
  assign n17667 = controllable_BtoR_REQ0 & ~n17666;
  assign n17668 = ~controllable_BtoR_REQ1 & ~n10061;
  assign n17669 = ~controllable_BtoR_REQ0 & ~n17668;
  assign n17670 = ~n17667 & ~n17669;
  assign n17671 = ~i_RtoB_ACK0 & ~n17670;
  assign n17672 = ~n15245 & ~n17671;
  assign n17673 = controllable_DEQ & ~n17672;
  assign n17674 = ~controllable_BtoR_REQ1 & ~n11284;
  assign n17675 = ~controllable_BtoR_REQ0 & ~n17674;
  assign n17676 = ~n17620 & ~n17675;
  assign n17677 = ~i_RtoB_ACK0 & ~n17676;
  assign n17678 = ~n17615 & ~n17677;
  assign n17679 = ~controllable_DEQ & ~n17678;
  assign n17680 = ~n17673 & ~n17679;
  assign n17681 = ~i_FULL & ~n17680;
  assign n17682 = ~n17663 & ~n17681;
  assign n17683 = ~i_nEMPTY & ~n17682;
  assign n17684 = ~n17641 & ~n17683;
  assign n17685 = controllable_BtoS_ACK0 & ~n17684;
  assign n17686 = ~i_RtoB_ACK1 & ~n11310;
  assign n17687 = ~n11299 & ~n17686;
  assign n17688 = ~controllable_BtoR_REQ1 & ~n17687;
  assign n17689 = ~controllable_BtoR_REQ1 & ~n17688;
  assign n17690 = controllable_BtoR_REQ0 & ~n17689;
  assign n17691 = ~controllable_BtoR_REQ1 & ~n11305;
  assign n17692 = ~controllable_BtoR_REQ0 & ~n17691;
  assign n17693 = ~n17690 & ~n17692;
  assign n17694 = i_RtoB_ACK0 & ~n17693;
  assign n17695 = i_RtoB_ACK1 & ~n11301;
  assign n17696 = ~n11313 & ~n17695;
  assign n17697 = ~controllable_BtoR_REQ1 & ~n17696;
  assign n17698 = ~controllable_BtoR_REQ1 & ~n17697;
  assign n17699 = controllable_BtoR_REQ0 & ~n17698;
  assign n17700 = ~controllable_BtoR_REQ1 & ~n11317;
  assign n17701 = ~controllable_BtoR_REQ0 & ~n17700;
  assign n17702 = ~n17699 & ~n17701;
  assign n17703 = ~i_RtoB_ACK0 & ~n17702;
  assign n17704 = ~n17694 & ~n17703;
  assign n17705 = controllable_DEQ & ~n17704;
  assign n17706 = ~n9904 & ~n11324;
  assign n17707 = ~controllable_BtoR_REQ1 & ~n17706;
  assign n17708 = ~controllable_BtoR_REQ1 & ~n17707;
  assign n17709 = controllable_BtoR_REQ0 & ~n17708;
  assign n17710 = ~controllable_BtoR_REQ1 & ~n11328;
  assign n17711 = ~controllable_BtoR_REQ0 & ~n17710;
  assign n17712 = ~n17709 & ~n17711;
  assign n17713 = i_RtoB_ACK0 & ~n17712;
  assign n17714 = i_RtoB_ACK1 & ~n9746;
  assign n17715 = ~n9904 & ~n17714;
  assign n17716 = ~controllable_BtoR_REQ1 & ~n17715;
  assign n17717 = ~controllable_BtoR_REQ1 & ~n17716;
  assign n17718 = controllable_BtoR_REQ0 & ~n17717;
  assign n17719 = ~n17711 & ~n17718;
  assign n17720 = ~i_RtoB_ACK0 & ~n17719;
  assign n17721 = ~n17713 & ~n17720;
  assign n17722 = ~controllable_DEQ & ~n17721;
  assign n17723 = ~n17705 & ~n17722;
  assign n17724 = i_nEMPTY & ~n17723;
  assign n17725 = ~i_RtoB_ACK1 & ~n11340;
  assign n17726 = ~i_RtoB_ACK1 & ~n17725;
  assign n17727 = ~controllable_BtoR_REQ1 & ~n17726;
  assign n17728 = ~controllable_BtoR_REQ1 & ~n17727;
  assign n17729 = controllable_BtoR_REQ0 & ~n17728;
  assign n17730 = controllable_BtoR_REQ0 & ~n17729;
  assign n17731 = i_RtoB_ACK0 & ~n17730;
  assign n17732 = ~i_RtoB_ACK1 & ~n11343;
  assign n17733 = ~controllable_BtoR_REQ1 & ~n17732;
  assign n17734 = ~controllable_BtoR_REQ1 & ~n17733;
  assign n17735 = controllable_BtoR_REQ0 & ~n17734;
  assign n17736 = ~controllable_BtoR_REQ1 & ~n9951;
  assign n17737 = ~controllable_BtoR_REQ0 & ~n17736;
  assign n17738 = ~n17735 & ~n17737;
  assign n17739 = ~i_RtoB_ACK0 & ~n17738;
  assign n17740 = ~n17731 & ~n17739;
  assign n17741 = controllable_DEQ & ~n17740;
  assign n17742 = ~n9871 & ~n11299;
  assign n17743 = ~controllable_BtoR_REQ1 & ~n17742;
  assign n17744 = ~controllable_BtoR_REQ1 & ~n17743;
  assign n17745 = controllable_BtoR_REQ0 & ~n17744;
  assign n17746 = ~n17692 & ~n17745;
  assign n17747 = i_RtoB_ACK0 & ~n17746;
  assign n17748 = ~n9871 & ~n17695;
  assign n17749 = ~controllable_BtoR_REQ1 & ~n17748;
  assign n17750 = ~controllable_BtoR_REQ1 & ~n17749;
  assign n17751 = controllable_BtoR_REQ0 & ~n17750;
  assign n17752 = ~n17692 & ~n17751;
  assign n17753 = ~i_RtoB_ACK0 & ~n17752;
  assign n17754 = ~n17747 & ~n17753;
  assign n17755 = ~controllable_DEQ & ~n17754;
  assign n17756 = ~n17741 & ~n17755;
  assign n17757 = i_FULL & ~n17756;
  assign n17758 = ~i_RtoB_ACK1 & ~n8945;
  assign n17759 = ~i_RtoB_ACK1 & ~n17758;
  assign n17760 = ~controllable_BtoR_REQ1 & ~n17759;
  assign n17761 = ~controllable_BtoR_REQ1 & ~n17760;
  assign n17762 = controllable_BtoR_REQ0 & ~n17761;
  assign n17763 = controllable_BtoR_REQ0 & ~n17762;
  assign n17764 = i_RtoB_ACK0 & ~n17763;
  assign n17765 = ~i_RtoB_ACK1 & ~n11325;
  assign n17766 = ~controllable_BtoR_REQ1 & ~n17765;
  assign n17767 = ~controllable_BtoR_REQ1 & ~n17766;
  assign n17768 = controllable_BtoR_REQ0 & ~n17767;
  assign n17769 = ~controllable_BtoR_REQ1 & ~n9973;
  assign n17770 = ~controllable_BtoR_REQ0 & ~n17769;
  assign n17771 = ~n17768 & ~n17770;
  assign n17772 = ~i_RtoB_ACK0 & ~n17771;
  assign n17773 = ~n17764 & ~n17772;
  assign n17774 = controllable_DEQ & ~n17773;
  assign n17775 = ~controllable_BtoR_REQ1 & ~n11366;
  assign n17776 = ~controllable_BtoR_REQ0 & ~n17775;
  assign n17777 = ~n17699 & ~n17776;
  assign n17778 = ~i_RtoB_ACK0 & ~n17777;
  assign n17779 = ~n17694 & ~n17778;
  assign n17780 = ~controllable_DEQ & ~n17779;
  assign n17781 = ~n17774 & ~n17780;
  assign n17782 = ~i_FULL & ~n17781;
  assign n17783 = ~n17757 & ~n17782;
  assign n17784 = ~i_nEMPTY & ~n17783;
  assign n17785 = ~n17724 & ~n17784;
  assign n17786 = ~controllable_BtoS_ACK0 & ~n17785;
  assign n17787 = ~n17685 & ~n17786;
  assign n17788 = ~i_StoB_REQ10 & ~n17787;
  assign n17789 = ~n17611 & ~n17788;
  assign n17790 = controllable_BtoS_ACK10 & ~n17789;
  assign n17791 = ~i_RtoB_ACK1 & ~n11403;
  assign n17792 = ~n5237 & ~n17791;
  assign n17793 = ~controllable_BtoR_REQ1 & ~n17792;
  assign n17794 = ~controllable_BtoR_REQ1 & ~n17793;
  assign n17795 = controllable_BtoR_REQ0 & ~n17794;
  assign n17796 = ~controllable_BtoR_REQ1 & ~n11393;
  assign n17797 = ~controllable_BtoR_REQ0 & ~n17796;
  assign n17798 = ~n17795 & ~n17797;
  assign n17799 = i_RtoB_ACK0 & ~n17798;
  assign n17800 = ~controllable_BtoR_REQ1 & ~n11412;
  assign n17801 = ~i_RtoB_ACK0 & ~n17800;
  assign n17802 = ~n17799 & ~n17801;
  assign n17803 = controllable_DEQ & ~n17802;
  assign n17804 = ~n7563 & ~n11429;
  assign n17805 = ~controllable_BtoR_REQ1 & ~n17804;
  assign n17806 = ~controllable_BtoR_REQ1 & ~n17805;
  assign n17807 = controllable_BtoR_REQ0 & ~n17806;
  assign n17808 = ~controllable_BtoR_REQ1 & ~n11422;
  assign n17809 = ~controllable_BtoR_REQ0 & ~n17808;
  assign n17810 = ~n17807 & ~n17809;
  assign n17811 = i_RtoB_ACK0 & ~n17810;
  assign n17812 = ~controllable_BtoR_REQ1 & ~n11431;
  assign n17813 = ~i_RtoB_ACK0 & ~n17812;
  assign n17814 = ~n17811 & ~n17813;
  assign n17815 = ~controllable_DEQ & ~n17814;
  assign n17816 = ~n17803 & ~n17815;
  assign n17817 = i_FULL & ~n17816;
  assign n17818 = ~i_RtoB_ACK1 & ~n11440;
  assign n17819 = ~n5237 & ~n17818;
  assign n17820 = ~controllable_BtoR_REQ1 & ~n17819;
  assign n17821 = ~controllable_BtoR_REQ1 & ~n17820;
  assign n17822 = controllable_BtoR_REQ0 & ~n17821;
  assign n17823 = ~n17797 & ~n17822;
  assign n17824 = i_RtoB_ACK0 & ~n17823;
  assign n17825 = ~controllable_BtoR_REQ1 & ~n11445;
  assign n17826 = ~i_RtoB_ACK0 & ~n17825;
  assign n17827 = ~n17824 & ~n17826;
  assign n17828 = controllable_DEQ & ~n17827;
  assign n17829 = ~n7563 & ~n11407;
  assign n17830 = ~controllable_BtoR_REQ1 & ~n17829;
  assign n17831 = ~controllable_BtoR_REQ1 & ~n17830;
  assign n17832 = controllable_BtoR_REQ0 & ~n17831;
  assign n17833 = ~n17809 & ~n17832;
  assign n17834 = i_RtoB_ACK0 & ~n17833;
  assign n17835 = ~controllable_BtoR_REQ1 & ~n11454;
  assign n17836 = ~i_RtoB_ACK0 & ~n17835;
  assign n17837 = ~n17834 & ~n17836;
  assign n17838 = ~controllable_DEQ & ~n17837;
  assign n17839 = ~n17828 & ~n17838;
  assign n17840 = ~i_FULL & ~n17839;
  assign n17841 = ~n17817 & ~n17840;
  assign n17842 = i_nEMPTY & ~n17841;
  assign n17843 = ~controllable_BtoR_REQ1 & ~n11470;
  assign n17844 = ~i_RtoB_ACK0 & ~n17843;
  assign n17845 = ~n15604 & ~n17844;
  assign n17846 = controllable_DEQ & ~n17845;
  assign n17847 = ~n5237 & ~n11479;
  assign n17848 = ~controllable_BtoR_REQ1 & ~n17847;
  assign n17849 = ~controllable_BtoR_REQ1 & ~n17848;
  assign n17850 = controllable_BtoR_REQ0 & ~n17849;
  assign n17851 = ~n17797 & ~n17850;
  assign n17852 = i_RtoB_ACK0 & ~n17851;
  assign n17853 = ~controllable_BtoR_REQ1 & ~n11481;
  assign n17854 = ~i_RtoB_ACK0 & ~n17853;
  assign n17855 = ~n17852 & ~n17854;
  assign n17856 = ~controllable_DEQ & ~n17855;
  assign n17857 = ~n17846 & ~n17856;
  assign n17858 = i_FULL & ~n17857;
  assign n17859 = ~controllable_BtoR_REQ1 & ~n11491;
  assign n17860 = ~i_RtoB_ACK0 & ~n17859;
  assign n17861 = ~n15619 & ~n17860;
  assign n17862 = controllable_DEQ & ~n17861;
  assign n17863 = ~controllable_DEQ & ~n17802;
  assign n17864 = ~n17862 & ~n17863;
  assign n17865 = ~i_FULL & ~n17864;
  assign n17866 = ~n17858 & ~n17865;
  assign n17867 = ~i_nEMPTY & ~n17866;
  assign n17868 = ~n17842 & ~n17867;
  assign n17869 = controllable_BtoS_ACK0 & ~n17868;
  assign n17870 = ~i_RtoB_ACK1 & ~n11520;
  assign n17871 = ~n8861 & ~n17870;
  assign n17872 = ~controllable_BtoR_REQ1 & ~n17871;
  assign n17873 = ~controllable_BtoR_REQ1 & ~n17872;
  assign n17874 = controllable_BtoR_REQ0 & ~n17873;
  assign n17875 = ~controllable_BtoR_REQ1 & ~n11515;
  assign n17876 = ~controllable_BtoR_REQ0 & ~n17875;
  assign n17877 = ~n17874 & ~n17876;
  assign n17878 = i_RtoB_ACK0 & ~n17877;
  assign n17879 = ~controllable_BtoR_REQ1 & ~n11529;
  assign n17880 = ~i_RtoB_ACK0 & ~n17879;
  assign n17881 = ~n17878 & ~n17880;
  assign n17882 = controllable_DEQ & ~n17881;
  assign n17883 = ~n7288 & ~n8883;
  assign n17884 = ~controllable_BtoR_REQ1 & ~n17883;
  assign n17885 = ~controllable_BtoR_REQ1 & ~n17884;
  assign n17886 = controllable_BtoR_REQ0 & ~n17885;
  assign n17887 = ~controllable_BtoR_REQ1 & ~n11539;
  assign n17888 = ~controllable_BtoR_REQ0 & ~n17887;
  assign n17889 = ~n17886 & ~n17888;
  assign n17890 = i_RtoB_ACK0 & ~n17889;
  assign n17891 = ~controllable_BtoR_REQ1 & ~n11546;
  assign n17892 = ~i_RtoB_ACK0 & ~n17891;
  assign n17893 = ~n17890 & ~n17892;
  assign n17894 = ~controllable_DEQ & ~n17893;
  assign n17895 = ~n17882 & ~n17894;
  assign n17896 = i_FULL & ~n17895;
  assign n17897 = ~i_RtoB_ACK1 & ~n11555;
  assign n17898 = ~n8861 & ~n17897;
  assign n17899 = ~controllable_BtoR_REQ1 & ~n17898;
  assign n17900 = ~controllable_BtoR_REQ1 & ~n17899;
  assign n17901 = controllable_BtoR_REQ0 & ~n17900;
  assign n17902 = ~n17876 & ~n17901;
  assign n17903 = i_RtoB_ACK0 & ~n17902;
  assign n17904 = ~controllable_BtoR_REQ1 & ~n11560;
  assign n17905 = ~i_RtoB_ACK0 & ~n17904;
  assign n17906 = ~n17903 & ~n17905;
  assign n17907 = controllable_DEQ & ~n17906;
  assign n17908 = ~n8883 & ~n11524;
  assign n17909 = ~controllable_BtoR_REQ1 & ~n17908;
  assign n17910 = ~controllable_BtoR_REQ1 & ~n17909;
  assign n17911 = controllable_BtoR_REQ0 & ~n17910;
  assign n17912 = ~n17888 & ~n17911;
  assign n17913 = i_RtoB_ACK0 & ~n17912;
  assign n17914 = ~controllable_BtoR_REQ1 & ~n11569;
  assign n17915 = ~i_RtoB_ACK0 & ~n17914;
  assign n17916 = ~n17913 & ~n17915;
  assign n17917 = ~controllable_DEQ & ~n17916;
  assign n17918 = ~n17907 & ~n17917;
  assign n17919 = ~i_FULL & ~n17918;
  assign n17920 = ~n17896 & ~n17919;
  assign n17921 = i_nEMPTY & ~n17920;
  assign n17922 = ~controllable_BtoR_REQ1 & ~n8917;
  assign n17923 = controllable_BtoR_REQ0 & ~n17922;
  assign n17924 = controllable_BtoR_REQ0 & ~n17923;
  assign n17925 = i_RtoB_ACK0 & ~n17924;
  assign n17926 = ~controllable_BtoR_REQ1 & ~n11586;
  assign n17927 = ~i_RtoB_ACK0 & ~n17926;
  assign n17928 = ~n17925 & ~n17927;
  assign n17929 = controllable_DEQ & ~n17928;
  assign n17930 = ~n7345 & ~n8861;
  assign n17931 = ~controllable_BtoR_REQ1 & ~n17930;
  assign n17932 = ~controllable_BtoR_REQ1 & ~n17931;
  assign n17933 = controllable_BtoR_REQ0 & ~n17932;
  assign n17934 = ~n17876 & ~n17933;
  assign n17935 = i_RtoB_ACK0 & ~n17934;
  assign n17936 = ~controllable_BtoR_REQ1 & ~n11594;
  assign n17937 = ~i_RtoB_ACK0 & ~n17936;
  assign n17938 = ~n17935 & ~n17937;
  assign n17939 = ~controllable_DEQ & ~n17938;
  assign n17940 = ~n17929 & ~n17939;
  assign n17941 = i_FULL & ~n17940;
  assign n17942 = controllable_BtoR_REQ0 & ~n16729;
  assign n17943 = i_RtoB_ACK0 & ~n17942;
  assign n17944 = ~controllable_BtoR_REQ1 & ~n11604;
  assign n17945 = ~i_RtoB_ACK0 & ~n17944;
  assign n17946 = ~n17943 & ~n17945;
  assign n17947 = controllable_DEQ & ~n17946;
  assign n17948 = ~controllable_DEQ & ~n17881;
  assign n17949 = ~n17947 & ~n17948;
  assign n17950 = ~i_FULL & ~n17949;
  assign n17951 = ~n17941 & ~n17950;
  assign n17952 = ~i_nEMPTY & ~n17951;
  assign n17953 = ~n17921 & ~n17952;
  assign n17954 = ~controllable_BtoS_ACK0 & ~n17953;
  assign n17955 = ~n17869 & ~n17954;
  assign n17956 = n4465 & ~n17955;
  assign n17957 = ~n15629 & ~n17954;
  assign n17958 = ~n4465 & ~n17957;
  assign n17959 = ~n17956 & ~n17958;
  assign n17960 = i_StoB_REQ10 & ~n17959;
  assign n17961 = ~i_RtoB_ACK1 & ~n11656;
  assign n17962 = ~n11632 & ~n17961;
  assign n17963 = ~controllable_BtoR_REQ1 & ~n17962;
  assign n17964 = ~controllable_BtoR_REQ1 & ~n17963;
  assign n17965 = controllable_BtoR_REQ0 & ~n17964;
  assign n17966 = ~controllable_BtoR_REQ1 & ~n11650;
  assign n17967 = ~controllable_BtoR_REQ0 & ~n17966;
  assign n17968 = ~n17965 & ~n17967;
  assign n17969 = i_RtoB_ACK0 & ~n17968;
  assign n17970 = i_RtoB_ACK1 & ~n11640;
  assign n17971 = ~n11660 & ~n17970;
  assign n17972 = ~controllable_BtoR_REQ1 & ~n17971;
  assign n17973 = ~controllable_BtoR_REQ1 & ~n17972;
  assign n17974 = controllable_BtoR_REQ0 & ~n17973;
  assign n17975 = ~controllable_BtoR_REQ1 & ~n11668;
  assign n17976 = ~controllable_BtoR_REQ0 & ~n17975;
  assign n17977 = ~n17974 & ~n17976;
  assign n17978 = ~i_RtoB_ACK0 & ~n17977;
  assign n17979 = ~n17969 & ~n17978;
  assign n17980 = controllable_DEQ & ~n17979;
  assign n17981 = ~n11429 & ~n11675;
  assign n17982 = ~controllable_BtoR_REQ1 & ~n17981;
  assign n17983 = ~controllable_BtoR_REQ1 & ~n17982;
  assign n17984 = controllable_BtoR_REQ0 & ~n17983;
  assign n17985 = ~controllable_BtoR_REQ1 & ~n11679;
  assign n17986 = ~controllable_BtoR_REQ0 & ~n17985;
  assign n17987 = ~n17984 & ~n17986;
  assign n17988 = i_RtoB_ACK0 & ~n17987;
  assign n17989 = i_RtoB_ACK1 & ~n11638;
  assign n17990 = ~n11429 & ~n17989;
  assign n17991 = ~controllable_BtoR_REQ1 & ~n17990;
  assign n17992 = ~controllable_BtoR_REQ1 & ~n17991;
  assign n17993 = controllable_BtoR_REQ0 & ~n17992;
  assign n17994 = ~controllable_BtoR_REQ1 & ~n11686;
  assign n17995 = ~controllable_BtoR_REQ0 & ~n17994;
  assign n17996 = ~n17993 & ~n17995;
  assign n17997 = ~i_RtoB_ACK0 & ~n17996;
  assign n17998 = ~n17988 & ~n17997;
  assign n17999 = ~controllable_DEQ & ~n17998;
  assign n18000 = ~n17980 & ~n17999;
  assign n18001 = i_FULL & ~n18000;
  assign n18002 = ~i_RtoB_ACK1 & ~n11695;
  assign n18003 = ~n11632 & ~n18002;
  assign n18004 = ~controllable_BtoR_REQ1 & ~n18003;
  assign n18005 = ~controllable_BtoR_REQ1 & ~n18004;
  assign n18006 = controllable_BtoR_REQ0 & ~n18005;
  assign n18007 = ~n17967 & ~n18006;
  assign n18008 = i_RtoB_ACK0 & ~n18007;
  assign n18009 = ~n11698 & ~n17970;
  assign n18010 = ~controllable_BtoR_REQ1 & ~n18009;
  assign n18011 = ~controllable_BtoR_REQ1 & ~n18010;
  assign n18012 = controllable_BtoR_REQ0 & ~n18011;
  assign n18013 = ~controllable_BtoR_REQ1 & ~n11703;
  assign n18014 = ~controllable_BtoR_REQ0 & ~n18013;
  assign n18015 = ~n18012 & ~n18014;
  assign n18016 = ~i_RtoB_ACK0 & ~n18015;
  assign n18017 = ~n18008 & ~n18016;
  assign n18018 = controllable_DEQ & ~n18017;
  assign n18019 = ~n11666 & ~n11675;
  assign n18020 = ~controllable_BtoR_REQ1 & ~n18019;
  assign n18021 = ~controllable_BtoR_REQ1 & ~n18020;
  assign n18022 = controllable_BtoR_REQ0 & ~n18021;
  assign n18023 = ~n17986 & ~n18022;
  assign n18024 = i_RtoB_ACK0 & ~n18023;
  assign n18025 = ~n11666 & ~n17989;
  assign n18026 = ~controllable_BtoR_REQ1 & ~n18025;
  assign n18027 = ~controllable_BtoR_REQ1 & ~n18026;
  assign n18028 = controllable_BtoR_REQ0 & ~n18027;
  assign n18029 = ~controllable_BtoR_REQ1 & ~n11712;
  assign n18030 = ~controllable_BtoR_REQ0 & ~n18029;
  assign n18031 = ~n18028 & ~n18030;
  assign n18032 = ~i_RtoB_ACK0 & ~n18031;
  assign n18033 = ~n18024 & ~n18032;
  assign n18034 = ~controllable_DEQ & ~n18033;
  assign n18035 = ~n18018 & ~n18034;
  assign n18036 = ~i_FULL & ~n18035;
  assign n18037 = ~n18001 & ~n18036;
  assign n18038 = i_nEMPTY & ~n18037;
  assign n18039 = ~i_RtoB_ACK1 & ~n11723;
  assign n18040 = ~i_RtoB_ACK1 & ~n18039;
  assign n18041 = ~controllable_BtoR_REQ1 & ~n18040;
  assign n18042 = ~controllable_BtoR_REQ1 & ~n18041;
  assign n18043 = controllable_BtoR_REQ0 & ~n18042;
  assign n18044 = controllable_BtoR_REQ0 & ~n18043;
  assign n18045 = i_RtoB_ACK0 & ~n18044;
  assign n18046 = ~i_RtoB_ACK1 & ~n11726;
  assign n18047 = ~controllable_BtoR_REQ1 & ~n18046;
  assign n18048 = ~controllable_BtoR_REQ1 & ~n18047;
  assign n18049 = controllable_BtoR_REQ0 & ~n18048;
  assign n18050 = ~controllable_BtoR_REQ1 & ~n11732;
  assign n18051 = ~controllable_BtoR_REQ0 & ~n18050;
  assign n18052 = ~n18049 & ~n18051;
  assign n18053 = ~i_RtoB_ACK0 & ~n18052;
  assign n18054 = ~n18045 & ~n18053;
  assign n18055 = controllable_DEQ & ~n18054;
  assign n18056 = ~n11479 & ~n11632;
  assign n18057 = ~controllable_BtoR_REQ1 & ~n18056;
  assign n18058 = ~controllable_BtoR_REQ1 & ~n18057;
  assign n18059 = controllable_BtoR_REQ0 & ~n18058;
  assign n18060 = ~n17967 & ~n18059;
  assign n18061 = i_RtoB_ACK0 & ~n18060;
  assign n18062 = ~n11479 & ~n17970;
  assign n18063 = ~controllable_BtoR_REQ1 & ~n18062;
  assign n18064 = ~controllable_BtoR_REQ1 & ~n18063;
  assign n18065 = controllable_BtoR_REQ0 & ~n18064;
  assign n18066 = ~controllable_BtoR_REQ1 & ~n11740;
  assign n18067 = ~controllable_BtoR_REQ0 & ~n18066;
  assign n18068 = ~n18065 & ~n18067;
  assign n18069 = ~i_RtoB_ACK0 & ~n18068;
  assign n18070 = ~n18061 & ~n18069;
  assign n18071 = ~controllable_DEQ & ~n18070;
  assign n18072 = ~n18055 & ~n18071;
  assign n18073 = i_FULL & ~n18072;
  assign n18074 = ~i_RtoB_ACK1 & ~n11629;
  assign n18075 = ~i_RtoB_ACK1 & ~n18074;
  assign n18076 = ~controllable_BtoR_REQ1 & ~n18075;
  assign n18077 = ~controllable_BtoR_REQ1 & ~n18076;
  assign n18078 = controllable_BtoR_REQ0 & ~n18077;
  assign n18079 = controllable_BtoR_REQ0 & ~n18078;
  assign n18080 = i_RtoB_ACK0 & ~n18079;
  assign n18081 = ~i_RtoB_ACK1 & ~n11676;
  assign n18082 = ~controllable_BtoR_REQ1 & ~n18081;
  assign n18083 = ~controllable_BtoR_REQ1 & ~n18082;
  assign n18084 = controllable_BtoR_REQ0 & ~n18083;
  assign n18085 = ~controllable_BtoR_REQ1 & ~n11750;
  assign n18086 = ~controllable_BtoR_REQ0 & ~n18085;
  assign n18087 = ~n18084 & ~n18086;
  assign n18088 = ~i_RtoB_ACK0 & ~n18087;
  assign n18089 = ~n18080 & ~n18088;
  assign n18090 = controllable_DEQ & ~n18089;
  assign n18091 = ~controllable_BtoR_REQ1 & ~n11758;
  assign n18092 = ~controllable_BtoR_REQ0 & ~n18091;
  assign n18093 = ~n17974 & ~n18092;
  assign n18094 = ~i_RtoB_ACK0 & ~n18093;
  assign n18095 = ~n17969 & ~n18094;
  assign n18096 = ~controllable_DEQ & ~n18095;
  assign n18097 = ~n18090 & ~n18096;
  assign n18098 = ~i_FULL & ~n18097;
  assign n18099 = ~n18073 & ~n18098;
  assign n18100 = ~i_nEMPTY & ~n18099;
  assign n18101 = ~n18038 & ~n18100;
  assign n18102 = controllable_BtoS_ACK0 & ~n18101;
  assign n18103 = ~i_RtoB_ACK1 & ~n11803;
  assign n18104 = ~n11779 & ~n18103;
  assign n18105 = ~controllable_BtoR_REQ1 & ~n18104;
  assign n18106 = ~controllable_BtoR_REQ1 & ~n18105;
  assign n18107 = controllable_BtoR_REQ0 & ~n18106;
  assign n18108 = ~controllable_BtoR_REQ1 & ~n11797;
  assign n18109 = ~controllable_BtoR_REQ0 & ~n18108;
  assign n18110 = ~n18107 & ~n18109;
  assign n18111 = i_RtoB_ACK0 & ~n18110;
  assign n18112 = i_RtoB_ACK1 & ~n11787;
  assign n18113 = ~n11807 & ~n18112;
  assign n18114 = ~controllable_BtoR_REQ1 & ~n18113;
  assign n18115 = ~controllable_BtoR_REQ1 & ~n18114;
  assign n18116 = controllable_BtoR_REQ0 & ~n18115;
  assign n18117 = ~controllable_BtoR_REQ1 & ~n11815;
  assign n18118 = ~controllable_BtoR_REQ0 & ~n18117;
  assign n18119 = ~n18116 & ~n18118;
  assign n18120 = ~i_RtoB_ACK0 & ~n18119;
  assign n18121 = ~n18111 & ~n18120;
  assign n18122 = controllable_DEQ & ~n18121;
  assign n18123 = ~n7288 & ~n11822;
  assign n18124 = ~controllable_BtoR_REQ1 & ~n18123;
  assign n18125 = ~controllable_BtoR_REQ1 & ~n18124;
  assign n18126 = controllable_BtoR_REQ0 & ~n18125;
  assign n18127 = ~controllable_BtoR_REQ1 & ~n11826;
  assign n18128 = ~controllable_BtoR_REQ0 & ~n18127;
  assign n18129 = ~n18126 & ~n18128;
  assign n18130 = i_RtoB_ACK0 & ~n18129;
  assign n18131 = i_RtoB_ACK1 & ~n11785;
  assign n18132 = ~n7288 & ~n18131;
  assign n18133 = ~controllable_BtoR_REQ1 & ~n18132;
  assign n18134 = ~controllable_BtoR_REQ1 & ~n18133;
  assign n18135 = controllable_BtoR_REQ0 & ~n18134;
  assign n18136 = ~controllable_BtoR_REQ1 & ~n11833;
  assign n18137 = ~controllable_BtoR_REQ0 & ~n18136;
  assign n18138 = ~n18135 & ~n18137;
  assign n18139 = ~i_RtoB_ACK0 & ~n18138;
  assign n18140 = ~n18130 & ~n18139;
  assign n18141 = ~controllable_DEQ & ~n18140;
  assign n18142 = ~n18122 & ~n18141;
  assign n18143 = i_FULL & ~n18142;
  assign n18144 = ~i_RtoB_ACK1 & ~n11842;
  assign n18145 = ~n11779 & ~n18144;
  assign n18146 = ~controllable_BtoR_REQ1 & ~n18145;
  assign n18147 = ~controllable_BtoR_REQ1 & ~n18146;
  assign n18148 = controllable_BtoR_REQ0 & ~n18147;
  assign n18149 = ~n18109 & ~n18148;
  assign n18150 = i_RtoB_ACK0 & ~n18149;
  assign n18151 = ~n11845 & ~n18112;
  assign n18152 = ~controllable_BtoR_REQ1 & ~n18151;
  assign n18153 = ~controllable_BtoR_REQ1 & ~n18152;
  assign n18154 = controllable_BtoR_REQ0 & ~n18153;
  assign n18155 = ~controllable_BtoR_REQ1 & ~n11850;
  assign n18156 = ~controllable_BtoR_REQ0 & ~n18155;
  assign n18157 = ~n18154 & ~n18156;
  assign n18158 = ~i_RtoB_ACK0 & ~n18157;
  assign n18159 = ~n18150 & ~n18158;
  assign n18160 = controllable_DEQ & ~n18159;
  assign n18161 = ~n11813 & ~n11822;
  assign n18162 = ~controllable_BtoR_REQ1 & ~n18161;
  assign n18163 = ~controllable_BtoR_REQ1 & ~n18162;
  assign n18164 = controllable_BtoR_REQ0 & ~n18163;
  assign n18165 = ~n18128 & ~n18164;
  assign n18166 = i_RtoB_ACK0 & ~n18165;
  assign n18167 = ~n11813 & ~n18131;
  assign n18168 = ~controllable_BtoR_REQ1 & ~n18167;
  assign n18169 = ~controllable_BtoR_REQ1 & ~n18168;
  assign n18170 = controllable_BtoR_REQ0 & ~n18169;
  assign n18171 = ~controllable_BtoR_REQ1 & ~n11859;
  assign n18172 = ~controllable_BtoR_REQ0 & ~n18171;
  assign n18173 = ~n18170 & ~n18172;
  assign n18174 = ~i_RtoB_ACK0 & ~n18173;
  assign n18175 = ~n18166 & ~n18174;
  assign n18176 = ~controllable_DEQ & ~n18175;
  assign n18177 = ~n18160 & ~n18176;
  assign n18178 = ~i_FULL & ~n18177;
  assign n18179 = ~n18143 & ~n18178;
  assign n18180 = i_nEMPTY & ~n18179;
  assign n18181 = ~i_RtoB_ACK1 & ~n11870;
  assign n18182 = ~i_RtoB_ACK1 & ~n18181;
  assign n18183 = ~controllable_BtoR_REQ1 & ~n18182;
  assign n18184 = ~controllable_BtoR_REQ1 & ~n18183;
  assign n18185 = controllable_BtoR_REQ0 & ~n18184;
  assign n18186 = controllable_BtoR_REQ0 & ~n18185;
  assign n18187 = i_RtoB_ACK0 & ~n18186;
  assign n18188 = ~i_RtoB_ACK1 & ~n11873;
  assign n18189 = ~controllable_BtoR_REQ1 & ~n18188;
  assign n18190 = ~controllable_BtoR_REQ1 & ~n18189;
  assign n18191 = controllable_BtoR_REQ0 & ~n18190;
  assign n18192 = ~controllable_BtoR_REQ1 & ~n11879;
  assign n18193 = ~controllable_BtoR_REQ0 & ~n18192;
  assign n18194 = ~n18191 & ~n18193;
  assign n18195 = ~i_RtoB_ACK0 & ~n18194;
  assign n18196 = ~n18187 & ~n18195;
  assign n18197 = controllable_DEQ & ~n18196;
  assign n18198 = ~n7345 & ~n11779;
  assign n18199 = ~controllable_BtoR_REQ1 & ~n18198;
  assign n18200 = ~controllable_BtoR_REQ1 & ~n18199;
  assign n18201 = controllable_BtoR_REQ0 & ~n18200;
  assign n18202 = ~n18109 & ~n18201;
  assign n18203 = i_RtoB_ACK0 & ~n18202;
  assign n18204 = ~n7345 & ~n18112;
  assign n18205 = ~controllable_BtoR_REQ1 & ~n18204;
  assign n18206 = ~controllable_BtoR_REQ1 & ~n18205;
  assign n18207 = controllable_BtoR_REQ0 & ~n18206;
  assign n18208 = ~controllable_BtoR_REQ1 & ~n11887;
  assign n18209 = ~controllable_BtoR_REQ0 & ~n18208;
  assign n18210 = ~n18207 & ~n18209;
  assign n18211 = ~i_RtoB_ACK0 & ~n18210;
  assign n18212 = ~n18203 & ~n18211;
  assign n18213 = ~controllable_DEQ & ~n18212;
  assign n18214 = ~n18197 & ~n18213;
  assign n18215 = i_FULL & ~n18214;
  assign n18216 = ~i_RtoB_ACK1 & ~n11776;
  assign n18217 = ~i_RtoB_ACK1 & ~n18216;
  assign n18218 = ~controllable_BtoR_REQ1 & ~n18217;
  assign n18219 = ~controllable_BtoR_REQ1 & ~n18218;
  assign n18220 = controllable_BtoR_REQ0 & ~n18219;
  assign n18221 = controllable_BtoR_REQ0 & ~n18220;
  assign n18222 = i_RtoB_ACK0 & ~n18221;
  assign n18223 = ~i_RtoB_ACK1 & ~n11823;
  assign n18224 = ~controllable_BtoR_REQ1 & ~n18223;
  assign n18225 = ~controllable_BtoR_REQ1 & ~n18224;
  assign n18226 = controllable_BtoR_REQ0 & ~n18225;
  assign n18227 = ~controllable_BtoR_REQ1 & ~n11897;
  assign n18228 = ~controllable_BtoR_REQ0 & ~n18227;
  assign n18229 = ~n18226 & ~n18228;
  assign n18230 = ~i_RtoB_ACK0 & ~n18229;
  assign n18231 = ~n18222 & ~n18230;
  assign n18232 = controllable_DEQ & ~n18231;
  assign n18233 = ~controllable_BtoR_REQ1 & ~n11905;
  assign n18234 = ~controllable_BtoR_REQ0 & ~n18233;
  assign n18235 = ~n18116 & ~n18234;
  assign n18236 = ~i_RtoB_ACK0 & ~n18235;
  assign n18237 = ~n18111 & ~n18236;
  assign n18238 = ~controllable_DEQ & ~n18237;
  assign n18239 = ~n18232 & ~n18238;
  assign n18240 = ~i_FULL & ~n18239;
  assign n18241 = ~n18215 & ~n18240;
  assign n18242 = ~i_nEMPTY & ~n18241;
  assign n18243 = ~n18180 & ~n18242;
  assign n18244 = ~controllable_BtoS_ACK0 & ~n18243;
  assign n18245 = ~n18102 & ~n18244;
  assign n18246 = n4465 & ~n18245;
  assign n18247 = ~n15411 & ~n18246;
  assign n18248 = ~i_StoB_REQ10 & ~n18247;
  assign n18249 = ~n17960 & ~n18248;
  assign n18250 = ~controllable_BtoS_ACK10 & ~n18249;
  assign n18251 = ~n17790 & ~n18250;
  assign n18252 = n4464 & ~n18251;
  assign n18253 = ~n15875 & ~n17788;
  assign n18254 = controllable_BtoS_ACK10 & ~n18253;
  assign n18255 = ~i_RtoB_ACK1 & ~n11939;
  assign n18256 = ~n5237 & ~n18255;
  assign n18257 = ~controllable_BtoR_REQ1 & ~n18256;
  assign n18258 = ~controllable_BtoR_REQ1 & ~n18257;
  assign n18259 = controllable_BtoR_REQ0 & ~n18258;
  assign n18260 = ~controllable_BtoR_REQ1 & ~n11934;
  assign n18261 = ~controllable_BtoR_REQ0 & ~n18260;
  assign n18262 = ~n18259 & ~n18261;
  assign n18263 = i_RtoB_ACK0 & ~n18262;
  assign n18264 = ~controllable_BtoR_REQ1 & ~n11948;
  assign n18265 = ~i_RtoB_ACK0 & ~n18264;
  assign n18266 = ~n18263 & ~n18265;
  assign n18267 = controllable_DEQ & ~n18266;
  assign n18268 = ~n7563 & ~n7958;
  assign n18269 = ~controllable_BtoR_REQ1 & ~n18268;
  assign n18270 = ~controllable_BtoR_REQ1 & ~n18269;
  assign n18271 = controllable_BtoR_REQ0 & ~n18270;
  assign n18272 = ~controllable_BtoR_REQ1 & ~n11958;
  assign n18273 = ~controllable_BtoR_REQ0 & ~n18272;
  assign n18274 = ~n18271 & ~n18273;
  assign n18275 = i_RtoB_ACK0 & ~n18274;
  assign n18276 = ~controllable_BtoR_REQ1 & ~n11965;
  assign n18277 = ~i_RtoB_ACK0 & ~n18276;
  assign n18278 = ~n18275 & ~n18277;
  assign n18279 = ~controllable_DEQ & ~n18278;
  assign n18280 = ~n18267 & ~n18279;
  assign n18281 = i_FULL & ~n18280;
  assign n18282 = ~i_RtoB_ACK1 & ~n11974;
  assign n18283 = ~n5237 & ~n18282;
  assign n18284 = ~controllable_BtoR_REQ1 & ~n18283;
  assign n18285 = ~controllable_BtoR_REQ1 & ~n18284;
  assign n18286 = controllable_BtoR_REQ0 & ~n18285;
  assign n18287 = ~n18261 & ~n18286;
  assign n18288 = i_RtoB_ACK0 & ~n18287;
  assign n18289 = ~controllable_BtoR_REQ1 & ~n11979;
  assign n18290 = ~i_RtoB_ACK0 & ~n18289;
  assign n18291 = ~n18288 & ~n18290;
  assign n18292 = controllable_DEQ & ~n18291;
  assign n18293 = ~n7563 & ~n11943;
  assign n18294 = ~controllable_BtoR_REQ1 & ~n18293;
  assign n18295 = ~controllable_BtoR_REQ1 & ~n18294;
  assign n18296 = controllable_BtoR_REQ0 & ~n18295;
  assign n18297 = ~n18273 & ~n18296;
  assign n18298 = i_RtoB_ACK0 & ~n18297;
  assign n18299 = ~controllable_BtoR_REQ1 & ~n11988;
  assign n18300 = ~i_RtoB_ACK0 & ~n18299;
  assign n18301 = ~n18298 & ~n18300;
  assign n18302 = ~controllable_DEQ & ~n18301;
  assign n18303 = ~n18292 & ~n18302;
  assign n18304 = ~i_FULL & ~n18303;
  assign n18305 = ~n18281 & ~n18304;
  assign n18306 = i_nEMPTY & ~n18305;
  assign n18307 = ~controllable_BtoR_REQ1 & ~n12004;
  assign n18308 = ~i_RtoB_ACK0 & ~n18307;
  assign n18309 = ~n15604 & ~n18308;
  assign n18310 = controllable_DEQ & ~n18309;
  assign n18311 = ~n5237 & ~n8015;
  assign n18312 = ~controllable_BtoR_REQ1 & ~n18311;
  assign n18313 = ~controllable_BtoR_REQ1 & ~n18312;
  assign n18314 = controllable_BtoR_REQ0 & ~n18313;
  assign n18315 = ~n18261 & ~n18314;
  assign n18316 = i_RtoB_ACK0 & ~n18315;
  assign n18317 = ~controllable_BtoR_REQ1 & ~n12012;
  assign n18318 = ~i_RtoB_ACK0 & ~n18317;
  assign n18319 = ~n18316 & ~n18318;
  assign n18320 = ~controllable_DEQ & ~n18319;
  assign n18321 = ~n18310 & ~n18320;
  assign n18322 = i_FULL & ~n18321;
  assign n18323 = ~controllable_BtoR_REQ1 & ~n12022;
  assign n18324 = ~i_RtoB_ACK0 & ~n18323;
  assign n18325 = ~n15619 & ~n18324;
  assign n18326 = controllable_DEQ & ~n18325;
  assign n18327 = ~controllable_DEQ & ~n18266;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = ~i_FULL & ~n18328;
  assign n18330 = ~n18322 & ~n18329;
  assign n18331 = ~i_nEMPTY & ~n18330;
  assign n18332 = ~n18306 & ~n18331;
  assign n18333 = controllable_BtoS_ACK0 & ~n18332;
  assign n18334 = ~i_RtoB_ACK1 & ~n12047;
  assign n18335 = ~n8861 & ~n18334;
  assign n18336 = ~controllable_BtoR_REQ1 & ~n18335;
  assign n18337 = ~controllable_BtoR_REQ1 & ~n18336;
  assign n18338 = controllable_BtoR_REQ0 & ~n18337;
  assign n18339 = ~controllable_BtoR_REQ1 & ~n12042;
  assign n18340 = ~controllable_BtoR_REQ0 & ~n18339;
  assign n18341 = ~n18338 & ~n18340;
  assign n18342 = i_RtoB_ACK0 & ~n18341;
  assign n18343 = ~controllable_BtoR_REQ1 & ~n12056;
  assign n18344 = ~i_RtoB_ACK0 & ~n18343;
  assign n18345 = ~n18342 & ~n18344;
  assign n18346 = controllable_DEQ & ~n18345;
  assign n18347 = ~n8122 & ~n8883;
  assign n18348 = ~controllable_BtoR_REQ1 & ~n18347;
  assign n18349 = ~controllable_BtoR_REQ1 & ~n18348;
  assign n18350 = controllable_BtoR_REQ0 & ~n18349;
  assign n18351 = ~controllable_BtoR_REQ1 & ~n12066;
  assign n18352 = ~controllable_BtoR_REQ0 & ~n18351;
  assign n18353 = ~n18350 & ~n18352;
  assign n18354 = i_RtoB_ACK0 & ~n18353;
  assign n18355 = ~controllable_BtoR_REQ1 & ~n12073;
  assign n18356 = ~i_RtoB_ACK0 & ~n18355;
  assign n18357 = ~n18354 & ~n18356;
  assign n18358 = ~controllable_DEQ & ~n18357;
  assign n18359 = ~n18346 & ~n18358;
  assign n18360 = i_FULL & ~n18359;
  assign n18361 = ~i_RtoB_ACK1 & ~n12082;
  assign n18362 = ~n8861 & ~n18361;
  assign n18363 = ~controllable_BtoR_REQ1 & ~n18362;
  assign n18364 = ~controllable_BtoR_REQ1 & ~n18363;
  assign n18365 = controllable_BtoR_REQ0 & ~n18364;
  assign n18366 = ~n18340 & ~n18365;
  assign n18367 = i_RtoB_ACK0 & ~n18366;
  assign n18368 = ~controllable_BtoR_REQ1 & ~n12087;
  assign n18369 = ~i_RtoB_ACK0 & ~n18368;
  assign n18370 = ~n18367 & ~n18369;
  assign n18371 = controllable_DEQ & ~n18370;
  assign n18372 = ~n8883 & ~n12051;
  assign n18373 = ~controllable_BtoR_REQ1 & ~n18372;
  assign n18374 = ~controllable_BtoR_REQ1 & ~n18373;
  assign n18375 = controllable_BtoR_REQ0 & ~n18374;
  assign n18376 = ~n18352 & ~n18375;
  assign n18377 = i_RtoB_ACK0 & ~n18376;
  assign n18378 = ~controllable_BtoR_REQ1 & ~n12096;
  assign n18379 = ~i_RtoB_ACK0 & ~n18378;
  assign n18380 = ~n18377 & ~n18379;
  assign n18381 = ~controllable_DEQ & ~n18380;
  assign n18382 = ~n18371 & ~n18381;
  assign n18383 = ~i_FULL & ~n18382;
  assign n18384 = ~n18360 & ~n18383;
  assign n18385 = i_nEMPTY & ~n18384;
  assign n18386 = ~controllable_BtoR_REQ1 & ~n12112;
  assign n18387 = ~i_RtoB_ACK0 & ~n18386;
  assign n18388 = ~n17925 & ~n18387;
  assign n18389 = controllable_DEQ & ~n18388;
  assign n18390 = ~n8179 & ~n8861;
  assign n18391 = ~controllable_BtoR_REQ1 & ~n18390;
  assign n18392 = ~controllable_BtoR_REQ1 & ~n18391;
  assign n18393 = controllable_BtoR_REQ0 & ~n18392;
  assign n18394 = ~n18340 & ~n18393;
  assign n18395 = i_RtoB_ACK0 & ~n18394;
  assign n18396 = ~controllable_BtoR_REQ1 & ~n12120;
  assign n18397 = ~i_RtoB_ACK0 & ~n18396;
  assign n18398 = ~n18395 & ~n18397;
  assign n18399 = ~controllable_DEQ & ~n18398;
  assign n18400 = ~n18389 & ~n18399;
  assign n18401 = i_FULL & ~n18400;
  assign n18402 = ~controllable_BtoR_REQ1 & ~n12130;
  assign n18403 = ~i_RtoB_ACK0 & ~n18402;
  assign n18404 = ~n17943 & ~n18403;
  assign n18405 = controllable_DEQ & ~n18404;
  assign n18406 = ~controllable_DEQ & ~n18345;
  assign n18407 = ~n18405 & ~n18406;
  assign n18408 = ~i_FULL & ~n18407;
  assign n18409 = ~n18401 & ~n18408;
  assign n18410 = ~i_nEMPTY & ~n18409;
  assign n18411 = ~n18385 & ~n18410;
  assign n18412 = ~controllable_BtoS_ACK0 & ~n18411;
  assign n18413 = ~n18333 & ~n18412;
  assign n18414 = n4465 & ~n18413;
  assign n18415 = ~n16605 & ~n18412;
  assign n18416 = ~n4465 & ~n18415;
  assign n18417 = ~n18414 & ~n18416;
  assign n18418 = i_StoB_REQ10 & ~n18417;
  assign n18419 = ~n16394 & ~n18418;
  assign n18420 = ~controllable_BtoS_ACK10 & ~n18419;
  assign n18421 = ~n18254 & ~n18420;
  assign n18422 = ~n4464 & ~n18421;
  assign n18423 = ~n18252 & ~n18422;
  assign n18424 = n4463 & ~n18423;
  assign n18425 = ~i_RtoB_ACK1 & ~n12164;
  assign n18426 = ~controllable_BtoR_REQ1 & ~n18425;
  assign n18427 = ~controllable_BtoR_REQ1 & ~n18426;
  assign n18428 = controllable_BtoR_REQ0 & ~n18427;
  assign n18429 = ~n17538 & ~n18428;
  assign n18430 = i_RtoB_ACK0 & ~n18429;
  assign n18431 = ~n17549 & ~n18430;
  assign n18432 = controllable_DEQ & ~n18431;
  assign n18433 = ~controllable_BtoR_REQ1 & ~n12228;
  assign n18434 = controllable_BtoR_REQ0 & ~n18433;
  assign n18435 = ~n17555 & ~n18434;
  assign n18436 = i_RtoB_ACK0 & ~n18435;
  assign n18437 = ~n17564 & ~n18436;
  assign n18438 = ~controllable_DEQ & ~n18437;
  assign n18439 = ~n18432 & ~n18438;
  assign n18440 = i_nEMPTY & ~n18439;
  assign n18441 = ~n17583 & ~n18430;
  assign n18442 = ~controllable_DEQ & ~n18441;
  assign n18443 = ~n17577 & ~n18442;
  assign n18444 = i_FULL & ~n18443;
  assign n18445 = ~n17599 & ~n18430;
  assign n18446 = ~controllable_DEQ & ~n18445;
  assign n18447 = ~n17595 & ~n18446;
  assign n18448 = ~i_FULL & ~n18447;
  assign n18449 = ~n18444 & ~n18448;
  assign n18450 = ~i_nEMPTY & ~n18449;
  assign n18451 = ~n18440 & ~n18450;
  assign n18452 = controllable_BtoS_ACK0 & ~n18451;
  assign n18453 = ~i_RtoB_ACK1 & ~n12257;
  assign n18454 = ~controllable_BtoR_REQ1 & ~n18453;
  assign n18455 = ~controllable_BtoR_REQ1 & ~n18454;
  assign n18456 = controllable_BtoR_REQ0 & ~n18455;
  assign n18457 = ~n14817 & ~n18456;
  assign n18458 = i_RtoB_ACK0 & ~n18457;
  assign n18459 = ~n14828 & ~n18458;
  assign n18460 = controllable_DEQ & ~n18459;
  assign n18461 = ~controllable_BtoR_REQ1 & ~n12309;
  assign n18462 = controllable_BtoR_REQ0 & ~n18461;
  assign n18463 = ~n14834 & ~n18462;
  assign n18464 = i_RtoB_ACK0 & ~n18463;
  assign n18465 = ~n14843 & ~n18464;
  assign n18466 = ~controllable_DEQ & ~n18465;
  assign n18467 = ~n18460 & ~n18466;
  assign n18468 = i_nEMPTY & ~n18467;
  assign n18469 = ~n14862 & ~n18458;
  assign n18470 = ~controllable_DEQ & ~n18469;
  assign n18471 = ~n14856 & ~n18470;
  assign n18472 = i_FULL & ~n18471;
  assign n18473 = ~n14878 & ~n18458;
  assign n18474 = ~controllable_DEQ & ~n18473;
  assign n18475 = ~n14874 & ~n18474;
  assign n18476 = ~i_FULL & ~n18475;
  assign n18477 = ~n18472 & ~n18476;
  assign n18478 = ~i_nEMPTY & ~n18477;
  assign n18479 = ~n18468 & ~n18478;
  assign n18480 = ~controllable_BtoS_ACK0 & ~n18479;
  assign n18481 = ~n18452 & ~n18480;
  assign n18482 = n4465 & ~n18481;
  assign n18483 = ~n16773 & ~n18482;
  assign n18484 = i_StoB_REQ10 & ~n18483;
  assign n18485 = ~n17788 & ~n18484;
  assign n18486 = controllable_BtoS_ACK10 & ~n18485;
  assign n18487 = ~n17050 & ~n17797;
  assign n18488 = i_RtoB_ACK0 & ~n18487;
  assign n18489 = ~n17801 & ~n18488;
  assign n18490 = controllable_DEQ & ~n18489;
  assign n18491 = ~n17058 & ~n17809;
  assign n18492 = i_RtoB_ACK0 & ~n18491;
  assign n18493 = ~n17813 & ~n18492;
  assign n18494 = ~controllable_DEQ & ~n18493;
  assign n18495 = ~n18490 & ~n18494;
  assign n18496 = i_FULL & ~n18495;
  assign n18497 = ~n17826 & ~n18488;
  assign n18498 = controllable_DEQ & ~n18497;
  assign n18499 = ~n17836 & ~n18492;
  assign n18500 = ~controllable_DEQ & ~n18499;
  assign n18501 = ~n18498 & ~n18500;
  assign n18502 = ~i_FULL & ~n18501;
  assign n18503 = ~n18496 & ~n18502;
  assign n18504 = i_nEMPTY & ~n18503;
  assign n18505 = ~n17068 & ~n17797;
  assign n18506 = i_RtoB_ACK0 & ~n18505;
  assign n18507 = ~n17854 & ~n18506;
  assign n18508 = ~controllable_DEQ & ~n18507;
  assign n18509 = ~n17846 & ~n18508;
  assign n18510 = i_FULL & ~n18509;
  assign n18511 = ~controllable_DEQ & ~n18489;
  assign n18512 = ~n17862 & ~n18511;
  assign n18513 = ~i_FULL & ~n18512;
  assign n18514 = ~n18510 & ~n18513;
  assign n18515 = ~i_nEMPTY & ~n18514;
  assign n18516 = ~n18504 & ~n18515;
  assign n18517 = controllable_BtoS_ACK0 & ~n18516;
  assign n18518 = ~i_RtoB_ACK1 & ~n12461;
  assign n18519 = ~n8861 & ~n18518;
  assign n18520 = ~controllable_BtoR_REQ1 & ~n18519;
  assign n18521 = ~controllable_BtoR_REQ1 & ~n18520;
  assign n18522 = controllable_BtoR_REQ0 & ~n18521;
  assign n18523 = ~n17876 & ~n18522;
  assign n18524 = i_RtoB_ACK0 & ~n18523;
  assign n18525 = ~n17880 & ~n18524;
  assign n18526 = controllable_DEQ & ~n18525;
  assign n18527 = ~n8883 & ~n9904;
  assign n18528 = ~controllable_BtoR_REQ1 & ~n18527;
  assign n18529 = ~controllable_BtoR_REQ1 & ~n18528;
  assign n18530 = controllable_BtoR_REQ0 & ~n18529;
  assign n18531 = ~n17888 & ~n18530;
  assign n18532 = i_RtoB_ACK0 & ~n18531;
  assign n18533 = ~n17892 & ~n18532;
  assign n18534 = ~controllable_DEQ & ~n18533;
  assign n18535 = ~n18526 & ~n18534;
  assign n18536 = i_FULL & ~n18535;
  assign n18537 = ~n17905 & ~n18524;
  assign n18538 = controllable_DEQ & ~n18537;
  assign n18539 = ~n17915 & ~n18532;
  assign n18540 = ~controllable_DEQ & ~n18539;
  assign n18541 = ~n18538 & ~n18540;
  assign n18542 = ~i_FULL & ~n18541;
  assign n18543 = ~n18536 & ~n18542;
  assign n18544 = i_nEMPTY & ~n18543;
  assign n18545 = ~n8861 & ~n9871;
  assign n18546 = ~controllable_BtoR_REQ1 & ~n18545;
  assign n18547 = ~controllable_BtoR_REQ1 & ~n18546;
  assign n18548 = controllable_BtoR_REQ0 & ~n18547;
  assign n18549 = ~n17876 & ~n18548;
  assign n18550 = i_RtoB_ACK0 & ~n18549;
  assign n18551 = ~n17937 & ~n18550;
  assign n18552 = ~controllable_DEQ & ~n18551;
  assign n18553 = ~n17929 & ~n18552;
  assign n18554 = i_FULL & ~n18553;
  assign n18555 = ~controllable_DEQ & ~n18525;
  assign n18556 = ~n17947 & ~n18555;
  assign n18557 = ~i_FULL & ~n18556;
  assign n18558 = ~n18554 & ~n18557;
  assign n18559 = ~i_nEMPTY & ~n18558;
  assign n18560 = ~n18544 & ~n18559;
  assign n18561 = ~controllable_BtoS_ACK0 & ~n18560;
  assign n18562 = ~n18517 & ~n18561;
  assign n18563 = n4465 & ~n18562;
  assign n18564 = ~n17081 & ~n18561;
  assign n18565 = ~n4465 & ~n18564;
  assign n18566 = ~n18563 & ~n18565;
  assign n18567 = i_StoB_REQ10 & ~n18566;
  assign n18568 = ~i_RtoB_ACK1 & ~n12554;
  assign n18569 = ~n11632 & ~n18568;
  assign n18570 = ~controllable_BtoR_REQ1 & ~n18569;
  assign n18571 = ~controllable_BtoR_REQ1 & ~n18570;
  assign n18572 = controllable_BtoR_REQ0 & ~n18571;
  assign n18573 = ~n17967 & ~n18572;
  assign n18574 = i_RtoB_ACK0 & ~n18573;
  assign n18575 = ~n17978 & ~n18574;
  assign n18576 = controllable_DEQ & ~n18575;
  assign n18577 = ~n9813 & ~n11675;
  assign n18578 = ~controllable_BtoR_REQ1 & ~n18577;
  assign n18579 = ~controllable_BtoR_REQ1 & ~n18578;
  assign n18580 = controllable_BtoR_REQ0 & ~n18579;
  assign n18581 = ~n17986 & ~n18580;
  assign n18582 = i_RtoB_ACK0 & ~n18581;
  assign n18583 = ~n17997 & ~n18582;
  assign n18584 = ~controllable_DEQ & ~n18583;
  assign n18585 = ~n18576 & ~n18584;
  assign n18586 = i_FULL & ~n18585;
  assign n18587 = ~n18016 & ~n18574;
  assign n18588 = controllable_DEQ & ~n18587;
  assign n18589 = ~n18032 & ~n18582;
  assign n18590 = ~controllable_DEQ & ~n18589;
  assign n18591 = ~n18588 & ~n18590;
  assign n18592 = ~i_FULL & ~n18591;
  assign n18593 = ~n18586 & ~n18592;
  assign n18594 = i_nEMPTY & ~n18593;
  assign n18595 = ~n9836 & ~n11632;
  assign n18596 = ~controllable_BtoR_REQ1 & ~n18595;
  assign n18597 = ~controllable_BtoR_REQ1 & ~n18596;
  assign n18598 = controllable_BtoR_REQ0 & ~n18597;
  assign n18599 = ~n17967 & ~n18598;
  assign n18600 = i_RtoB_ACK0 & ~n18599;
  assign n18601 = ~n18069 & ~n18600;
  assign n18602 = ~controllable_DEQ & ~n18601;
  assign n18603 = ~n18055 & ~n18602;
  assign n18604 = i_FULL & ~n18603;
  assign n18605 = ~n18094 & ~n18574;
  assign n18606 = ~controllable_DEQ & ~n18605;
  assign n18607 = ~n18090 & ~n18606;
  assign n18608 = ~i_FULL & ~n18607;
  assign n18609 = ~n18604 & ~n18608;
  assign n18610 = ~i_nEMPTY & ~n18609;
  assign n18611 = ~n18594 & ~n18610;
  assign n18612 = controllable_BtoS_ACK0 & ~n18611;
  assign n18613 = ~i_RtoB_ACK1 & ~n12650;
  assign n18614 = ~n11779 & ~n18613;
  assign n18615 = ~controllable_BtoR_REQ1 & ~n18614;
  assign n18616 = ~controllable_BtoR_REQ1 & ~n18615;
  assign n18617 = controllable_BtoR_REQ0 & ~n18616;
  assign n18618 = ~n18109 & ~n18617;
  assign n18619 = i_RtoB_ACK0 & ~n18618;
  assign n18620 = ~n18120 & ~n18619;
  assign n18621 = controllable_DEQ & ~n18620;
  assign n18622 = ~n9904 & ~n11822;
  assign n18623 = ~controllable_BtoR_REQ1 & ~n18622;
  assign n18624 = ~controllable_BtoR_REQ1 & ~n18623;
  assign n18625 = controllable_BtoR_REQ0 & ~n18624;
  assign n18626 = ~n18128 & ~n18625;
  assign n18627 = i_RtoB_ACK0 & ~n18626;
  assign n18628 = ~n18139 & ~n18627;
  assign n18629 = ~controllable_DEQ & ~n18628;
  assign n18630 = ~n18621 & ~n18629;
  assign n18631 = i_FULL & ~n18630;
  assign n18632 = ~n18158 & ~n18619;
  assign n18633 = controllable_DEQ & ~n18632;
  assign n18634 = ~n18174 & ~n18627;
  assign n18635 = ~controllable_DEQ & ~n18634;
  assign n18636 = ~n18633 & ~n18635;
  assign n18637 = ~i_FULL & ~n18636;
  assign n18638 = ~n18631 & ~n18637;
  assign n18639 = i_nEMPTY & ~n18638;
  assign n18640 = ~n9871 & ~n11779;
  assign n18641 = ~controllable_BtoR_REQ1 & ~n18640;
  assign n18642 = ~controllable_BtoR_REQ1 & ~n18641;
  assign n18643 = controllable_BtoR_REQ0 & ~n18642;
  assign n18644 = ~n18109 & ~n18643;
  assign n18645 = i_RtoB_ACK0 & ~n18644;
  assign n18646 = ~n18211 & ~n18645;
  assign n18647 = ~controllable_DEQ & ~n18646;
  assign n18648 = ~n18197 & ~n18647;
  assign n18649 = i_FULL & ~n18648;
  assign n18650 = ~n18236 & ~n18619;
  assign n18651 = ~controllable_DEQ & ~n18650;
  assign n18652 = ~n18232 & ~n18651;
  assign n18653 = ~i_FULL & ~n18652;
  assign n18654 = ~n18649 & ~n18653;
  assign n18655 = ~i_nEMPTY & ~n18654;
  assign n18656 = ~n18639 & ~n18655;
  assign n18657 = ~controllable_BtoS_ACK0 & ~n18656;
  assign n18658 = ~n18612 & ~n18657;
  assign n18659 = n4465 & ~n18658;
  assign n18660 = ~n15183 & ~n17280;
  assign n18661 = i_RtoB_ACK0 & ~n18660;
  assign n18662 = ~n15194 & ~n18661;
  assign n18663 = controllable_DEQ & ~n18662;
  assign n18664 = ~n15202 & ~n17288;
  assign n18665 = i_RtoB_ACK0 & ~n18664;
  assign n18666 = ~n15211 & ~n18665;
  assign n18667 = ~controllable_DEQ & ~n18666;
  assign n18668 = ~n18663 & ~n18667;
  assign n18669 = i_nEMPTY & ~n18668;
  assign n18670 = ~n15183 & ~n17298;
  assign n18671 = i_RtoB_ACK0 & ~n18670;
  assign n18672 = ~n15239 & ~n18671;
  assign n18673 = ~controllable_DEQ & ~n18672;
  assign n18674 = ~n15227 & ~n18673;
  assign n18675 = i_FULL & ~n18674;
  assign n18676 = ~n15259 & ~n18661;
  assign n18677 = ~controllable_DEQ & ~n18676;
  assign n18678 = ~n15255 & ~n18677;
  assign n18679 = ~i_FULL & ~n18678;
  assign n18680 = ~n18675 & ~n18679;
  assign n18681 = ~i_nEMPTY & ~n18680;
  assign n18682 = ~n18669 & ~n18681;
  assign n18683 = controllable_BtoS_ACK0 & ~n18682;
  assign n18684 = ~n16949 & ~n18683;
  assign n18685 = ~n4465 & ~n18684;
  assign n18686 = ~n18659 & ~n18685;
  assign n18687 = ~i_StoB_REQ10 & ~n18686;
  assign n18688 = ~n18567 & ~n18687;
  assign n18689 = ~controllable_BtoS_ACK10 & ~n18688;
  assign n18690 = ~n18486 & ~n18689;
  assign n18691 = n4464 & ~n18690;
  assign n18692 = ~n17183 & ~n17788;
  assign n18693 = controllable_BtoS_ACK10 & ~n18692;
  assign n18694 = ~n17050 & ~n18261;
  assign n18695 = i_RtoB_ACK0 & ~n18694;
  assign n18696 = ~n18265 & ~n18695;
  assign n18697 = controllable_DEQ & ~n18696;
  assign n18698 = ~n17058 & ~n18273;
  assign n18699 = i_RtoB_ACK0 & ~n18698;
  assign n18700 = ~n18277 & ~n18699;
  assign n18701 = ~controllable_DEQ & ~n18700;
  assign n18702 = ~n18697 & ~n18701;
  assign n18703 = i_FULL & ~n18702;
  assign n18704 = ~n18290 & ~n18695;
  assign n18705 = controllable_DEQ & ~n18704;
  assign n18706 = ~n18300 & ~n18699;
  assign n18707 = ~controllable_DEQ & ~n18706;
  assign n18708 = ~n18705 & ~n18707;
  assign n18709 = ~i_FULL & ~n18708;
  assign n18710 = ~n18703 & ~n18709;
  assign n18711 = i_nEMPTY & ~n18710;
  assign n18712 = ~n17068 & ~n18261;
  assign n18713 = i_RtoB_ACK0 & ~n18712;
  assign n18714 = ~n18318 & ~n18713;
  assign n18715 = ~controllable_DEQ & ~n18714;
  assign n18716 = ~n18310 & ~n18715;
  assign n18717 = i_FULL & ~n18716;
  assign n18718 = ~controllable_DEQ & ~n18696;
  assign n18719 = ~n18326 & ~n18718;
  assign n18720 = ~i_FULL & ~n18719;
  assign n18721 = ~n18717 & ~n18720;
  assign n18722 = ~i_nEMPTY & ~n18721;
  assign n18723 = ~n18711 & ~n18722;
  assign n18724 = controllable_BtoS_ACK0 & ~n18723;
  assign n18725 = ~n18340 & ~n18522;
  assign n18726 = i_RtoB_ACK0 & ~n18725;
  assign n18727 = ~n18344 & ~n18726;
  assign n18728 = controllable_DEQ & ~n18727;
  assign n18729 = ~n18352 & ~n18530;
  assign n18730 = i_RtoB_ACK0 & ~n18729;
  assign n18731 = ~n18356 & ~n18730;
  assign n18732 = ~controllable_DEQ & ~n18731;
  assign n18733 = ~n18728 & ~n18732;
  assign n18734 = i_FULL & ~n18733;
  assign n18735 = ~n18369 & ~n18726;
  assign n18736 = controllable_DEQ & ~n18735;
  assign n18737 = ~n18379 & ~n18730;
  assign n18738 = ~controllable_DEQ & ~n18737;
  assign n18739 = ~n18736 & ~n18738;
  assign n18740 = ~i_FULL & ~n18739;
  assign n18741 = ~n18734 & ~n18740;
  assign n18742 = i_nEMPTY & ~n18741;
  assign n18743 = ~n18340 & ~n18548;
  assign n18744 = i_RtoB_ACK0 & ~n18743;
  assign n18745 = ~n18397 & ~n18744;
  assign n18746 = ~controllable_DEQ & ~n18745;
  assign n18747 = ~n18389 & ~n18746;
  assign n18748 = i_FULL & ~n18747;
  assign n18749 = ~controllable_DEQ & ~n18727;
  assign n18750 = ~n18405 & ~n18749;
  assign n18751 = ~i_FULL & ~n18750;
  assign n18752 = ~n18748 & ~n18751;
  assign n18753 = ~i_nEMPTY & ~n18752;
  assign n18754 = ~n18742 & ~n18753;
  assign n18755 = ~controllable_BtoS_ACK0 & ~n18754;
  assign n18756 = ~n18724 & ~n18755;
  assign n18757 = n4465 & ~n18756;
  assign n18758 = ~n17476 & ~n18755;
  assign n18759 = ~n4465 & ~n18758;
  assign n18760 = ~n18757 & ~n18759;
  assign n18761 = i_StoB_REQ10 & ~n18760;
  assign n18762 = ~i_RtoB_ACK1 & ~n10467;
  assign n18763 = ~n7886 & ~n18762;
  assign n18764 = ~controllable_BtoR_REQ1 & ~n18763;
  assign n18765 = ~controllable_BtoR_REQ1 & ~n18764;
  assign n18766 = controllable_BtoR_REQ0 & ~n18765;
  assign n18767 = ~n15882 & ~n18766;
  assign n18768 = i_RtoB_ACK0 & ~n18767;
  assign n18769 = ~n15893 & ~n18768;
  assign n18770 = controllable_DEQ & ~n18769;
  assign n18771 = ~n7947 & ~n9813;
  assign n18772 = ~controllable_BtoR_REQ1 & ~n18771;
  assign n18773 = ~controllable_BtoR_REQ1 & ~n18772;
  assign n18774 = controllable_BtoR_REQ0 & ~n18773;
  assign n18775 = ~n15901 & ~n18774;
  assign n18776 = i_RtoB_ACK0 & ~n18775;
  assign n18777 = ~n15912 & ~n18776;
  assign n18778 = ~controllable_DEQ & ~n18777;
  assign n18779 = ~n18770 & ~n18778;
  assign n18780 = i_FULL & ~n18779;
  assign n18781 = ~n15931 & ~n18768;
  assign n18782 = controllable_DEQ & ~n18781;
  assign n18783 = ~n15947 & ~n18776;
  assign n18784 = ~controllable_DEQ & ~n18783;
  assign n18785 = ~n18782 & ~n18784;
  assign n18786 = ~i_FULL & ~n18785;
  assign n18787 = ~n18780 & ~n18786;
  assign n18788 = i_nEMPTY & ~n18787;
  assign n18789 = ~n7886 & ~n9836;
  assign n18790 = ~controllable_BtoR_REQ1 & ~n18789;
  assign n18791 = ~controllable_BtoR_REQ1 & ~n18790;
  assign n18792 = controllable_BtoR_REQ0 & ~n18791;
  assign n18793 = ~n15882 & ~n18792;
  assign n18794 = i_RtoB_ACK0 & ~n18793;
  assign n18795 = ~n15984 & ~n18794;
  assign n18796 = ~controllable_DEQ & ~n18795;
  assign n18797 = ~n15970 & ~n18796;
  assign n18798 = i_FULL & ~n18797;
  assign n18799 = ~n16009 & ~n18768;
  assign n18800 = ~controllable_DEQ & ~n18799;
  assign n18801 = ~n16005 & ~n18800;
  assign n18802 = ~i_FULL & ~n18801;
  assign n18803 = ~n18798 & ~n18802;
  assign n18804 = ~i_nEMPTY & ~n18803;
  assign n18805 = ~n18788 & ~n18804;
  assign n18806 = controllable_BtoS_ACK0 & ~n18805;
  assign n18807 = ~i_RtoB_ACK1 & ~n10597;
  assign n18808 = ~n8057 & ~n18807;
  assign n18809 = ~controllable_BtoR_REQ1 & ~n18808;
  assign n18810 = ~controllable_BtoR_REQ1 & ~n18809;
  assign n18811 = controllable_BtoR_REQ0 & ~n18810;
  assign n18812 = ~n16024 & ~n18811;
  assign n18813 = i_RtoB_ACK0 & ~n18812;
  assign n18814 = ~n16035 & ~n18813;
  assign n18815 = controllable_DEQ & ~n18814;
  assign n18816 = ~n8111 & ~n9904;
  assign n18817 = ~controllable_BtoR_REQ1 & ~n18816;
  assign n18818 = ~controllable_BtoR_REQ1 & ~n18817;
  assign n18819 = controllable_BtoR_REQ0 & ~n18818;
  assign n18820 = ~n16043 & ~n18819;
  assign n18821 = i_RtoB_ACK0 & ~n18820;
  assign n18822 = ~n16054 & ~n18821;
  assign n18823 = ~controllable_DEQ & ~n18822;
  assign n18824 = ~n18815 & ~n18823;
  assign n18825 = i_FULL & ~n18824;
  assign n18826 = ~n16073 & ~n18813;
  assign n18827 = controllable_DEQ & ~n18826;
  assign n18828 = ~n16089 & ~n18821;
  assign n18829 = ~controllable_DEQ & ~n18828;
  assign n18830 = ~n18827 & ~n18829;
  assign n18831 = ~i_FULL & ~n18830;
  assign n18832 = ~n18825 & ~n18831;
  assign n18833 = i_nEMPTY & ~n18832;
  assign n18834 = ~n8057 & ~n9871;
  assign n18835 = ~controllable_BtoR_REQ1 & ~n18834;
  assign n18836 = ~controllable_BtoR_REQ1 & ~n18835;
  assign n18837 = controllable_BtoR_REQ0 & ~n18836;
  assign n18838 = ~n16024 & ~n18837;
  assign n18839 = i_RtoB_ACK0 & ~n18838;
  assign n18840 = ~n16126 & ~n18839;
  assign n18841 = ~controllable_DEQ & ~n18840;
  assign n18842 = ~n16112 & ~n18841;
  assign n18843 = i_FULL & ~n18842;
  assign n18844 = ~n16151 & ~n18813;
  assign n18845 = ~controllable_DEQ & ~n18844;
  assign n18846 = ~n16147 & ~n18845;
  assign n18847 = ~i_FULL & ~n18846;
  assign n18848 = ~n18843 & ~n18847;
  assign n18849 = ~i_nEMPTY & ~n18848;
  assign n18850 = ~n18833 & ~n18849;
  assign n18851 = ~controllable_BtoS_ACK0 & ~n18850;
  assign n18852 = ~n18806 & ~n18851;
  assign n18853 = n4465 & ~n18852;
  assign n18854 = ~n17359 & ~n18853;
  assign n18855 = ~i_StoB_REQ10 & ~n18854;
  assign n18856 = ~n18761 & ~n18855;
  assign n18857 = ~controllable_BtoS_ACK10 & ~n18856;
  assign n18858 = ~n18693 & ~n18857;
  assign n18859 = ~n4464 & ~n18858;
  assign n18860 = ~n18691 & ~n18859;
  assign n18861 = ~n4463 & ~n18860;
  assign n18862 = ~n18424 & ~n18861;
  assign n18863 = ~n4462 & ~n18862;
  assign n18864 = ~n17532 & ~n18863;
  assign n18865 = n4461 & ~n18864;
  assign n18866 = ~n5237 & ~n8765;
  assign n18867 = ~controllable_BtoR_REQ1 & ~n18866;
  assign n18868 = ~controllable_BtoR_REQ1 & ~n18867;
  assign n18869 = ~controllable_BtoR_REQ0 & ~n18868;
  assign n18870 = ~n14598 & ~n18869;
  assign n18871 = ~i_RtoB_ACK0 & ~n18870;
  assign n18872 = ~n16699 & ~n18871;
  assign n18873 = controllable_DEQ & ~n18872;
  assign n18874 = ~controllable_BtoR_REQ1 & ~n8781;
  assign n18875 = ~controllable_BtoR_REQ1 & ~n18874;
  assign n18876 = ~controllable_BtoR_REQ0 & ~n18875;
  assign n18877 = ~n14615 & ~n18876;
  assign n18878 = ~i_RtoB_ACK0 & ~n18877;
  assign n18879 = ~n16703 & ~n18878;
  assign n18880 = ~controllable_DEQ & ~n18879;
  assign n18881 = ~n18873 & ~n18880;
  assign n18882 = i_FULL & ~n18881;
  assign n18883 = ~n14598 & ~n14751;
  assign n18884 = ~i_RtoB_ACK0 & ~n18883;
  assign n18885 = ~n16699 & ~n18884;
  assign n18886 = controllable_DEQ & ~n18885;
  assign n18887 = ~n7563 & ~n8765;
  assign n18888 = ~controllable_BtoR_REQ1 & ~n18887;
  assign n18889 = ~controllable_BtoR_REQ1 & ~n18888;
  assign n18890 = ~controllable_BtoR_REQ0 & ~n18889;
  assign n18891 = ~n14615 & ~n18890;
  assign n18892 = ~i_RtoB_ACK0 & ~n18891;
  assign n18893 = ~n16703 & ~n18892;
  assign n18894 = ~controllable_DEQ & ~n18893;
  assign n18895 = ~n18886 & ~n18894;
  assign n18896 = ~i_FULL & ~n18895;
  assign n18897 = ~n18882 & ~n18896;
  assign n18898 = i_nEMPTY & ~n18897;
  assign n18899 = ~n14624 & ~n14776;
  assign n18900 = ~i_RtoB_ACK0 & ~n18899;
  assign n18901 = ~i_RtoB_ACK0 & ~n18900;
  assign n18902 = controllable_DEQ & ~n18901;
  assign n18903 = ~controllable_BtoR_REQ1 & ~n8818;
  assign n18904 = ~controllable_BtoR_REQ1 & ~n18903;
  assign n18905 = ~controllable_BtoR_REQ0 & ~n18904;
  assign n18906 = ~n14634 & ~n18905;
  assign n18907 = ~i_RtoB_ACK0 & ~n18906;
  assign n18908 = ~n16699 & ~n18907;
  assign n18909 = ~controllable_DEQ & ~n18908;
  assign n18910 = ~n18902 & ~n18909;
  assign n18911 = i_FULL & ~n18910;
  assign n18912 = ~n14643 & ~n14794;
  assign n18913 = ~i_RtoB_ACK0 & ~n18912;
  assign n18914 = ~i_RtoB_ACK0 & ~n18913;
  assign n18915 = controllable_DEQ & ~n18914;
  assign n18916 = ~n5237 & ~n8835;
  assign n18917 = ~controllable_BtoR_REQ1 & ~n18916;
  assign n18918 = ~controllable_BtoR_REQ1 & ~n18917;
  assign n18919 = ~controllable_BtoR_REQ0 & ~n18918;
  assign n18920 = ~n14598 & ~n18919;
  assign n18921 = ~i_RtoB_ACK0 & ~n18920;
  assign n18922 = ~n16699 & ~n18921;
  assign n18923 = ~controllable_DEQ & ~n18922;
  assign n18924 = ~n18915 & ~n18923;
  assign n18925 = ~i_FULL & ~n18924;
  assign n18926 = ~n18911 & ~n18925;
  assign n18927 = ~i_nEMPTY & ~n18926;
  assign n18928 = ~n18898 & ~n18927;
  assign n18929 = controllable_BtoS_ACK0 & ~n18928;
  assign n18930 = ~n8861 & ~n8866;
  assign n18931 = ~controllable_BtoR_REQ1 & ~n18930;
  assign n18932 = ~controllable_BtoR_REQ1 & ~n18931;
  assign n18933 = ~controllable_BtoR_REQ0 & ~n18932;
  assign n18934 = ~n14673 & ~n18933;
  assign n18935 = ~i_RtoB_ACK0 & ~n18934;
  assign n18936 = ~n16725 & ~n18935;
  assign n18937 = controllable_DEQ & ~n18936;
  assign n18938 = ~controllable_BtoR_REQ1 & ~n8884;
  assign n18939 = ~controllable_BtoR_REQ1 & ~n18938;
  assign n18940 = ~controllable_BtoR_REQ0 & ~n18939;
  assign n18941 = ~n14690 & ~n18940;
  assign n18942 = ~i_RtoB_ACK0 & ~n18941;
  assign n18943 = ~n16731 & ~n18942;
  assign n18944 = ~controllable_DEQ & ~n18943;
  assign n18945 = ~n18937 & ~n18944;
  assign n18946 = i_FULL & ~n18945;
  assign n18947 = ~n8861 & ~n8876;
  assign n18948 = ~controllable_BtoR_REQ1 & ~n18947;
  assign n18949 = ~controllable_BtoR_REQ1 & ~n18948;
  assign n18950 = ~controllable_BtoR_REQ0 & ~n18949;
  assign n18951 = ~n14673 & ~n18950;
  assign n18952 = ~i_RtoB_ACK0 & ~n18951;
  assign n18953 = ~n16725 & ~n18952;
  assign n18954 = controllable_DEQ & ~n18953;
  assign n18955 = ~n8866 & ~n8883;
  assign n18956 = ~controllable_BtoR_REQ1 & ~n18955;
  assign n18957 = ~controllable_BtoR_REQ1 & ~n18956;
  assign n18958 = ~controllable_BtoR_REQ0 & ~n18957;
  assign n18959 = ~n14690 & ~n18958;
  assign n18960 = ~i_RtoB_ACK0 & ~n18959;
  assign n18961 = ~n16731 & ~n18960;
  assign n18962 = ~controllable_DEQ & ~n18961;
  assign n18963 = ~n18954 & ~n18962;
  assign n18964 = ~i_FULL & ~n18963;
  assign n18965 = ~n18946 & ~n18964;
  assign n18966 = i_nEMPTY & ~n18965;
  assign n18967 = ~controllable_BtoR_REQ0 & ~n17922;
  assign n18968 = ~n14699 & ~n18967;
  assign n18969 = ~i_RtoB_ACK0 & ~n18968;
  assign n18970 = ~i_RtoB_ACK0 & ~n18969;
  assign n18971 = controllable_DEQ & ~n18970;
  assign n18972 = ~controllable_BtoR_REQ1 & ~n8925;
  assign n18973 = ~controllable_BtoR_REQ1 & ~n18972;
  assign n18974 = ~controllable_BtoR_REQ0 & ~n18973;
  assign n18975 = ~n14709 & ~n18974;
  assign n18976 = ~i_RtoB_ACK0 & ~n18975;
  assign n18977 = ~n16725 & ~n18976;
  assign n18978 = ~controllable_DEQ & ~n18977;
  assign n18979 = ~n18971 & ~n18978;
  assign n18980 = i_FULL & ~n18979;
  assign n18981 = ~controllable_BtoR_REQ0 & ~n16728;
  assign n18982 = ~n14718 & ~n18981;
  assign n18983 = ~i_RtoB_ACK0 & ~n18982;
  assign n18984 = ~i_RtoB_ACK0 & ~n18983;
  assign n18985 = controllable_DEQ & ~n18984;
  assign n18986 = ~n8861 & ~n8948;
  assign n18987 = ~controllable_BtoR_REQ1 & ~n18986;
  assign n18988 = ~controllable_BtoR_REQ1 & ~n18987;
  assign n18989 = ~controllable_BtoR_REQ0 & ~n18988;
  assign n18990 = ~n14673 & ~n18989;
  assign n18991 = ~i_RtoB_ACK0 & ~n18990;
  assign n18992 = ~n16725 & ~n18991;
  assign n18993 = ~controllable_DEQ & ~n18992;
  assign n18994 = ~n18985 & ~n18993;
  assign n18995 = ~i_FULL & ~n18994;
  assign n18996 = ~n18980 & ~n18995;
  assign n18997 = ~i_nEMPTY & ~n18996;
  assign n18998 = ~n18966 & ~n18997;
  assign n18999 = ~controllable_BtoS_ACK0 & ~n18998;
  assign n19000 = ~n18929 & ~n18999;
  assign n19001 = n4465 & ~n19000;
  assign n19002 = ~n8861 & ~n8974;
  assign n19003 = ~controllable_BtoR_REQ1 & ~n19002;
  assign n19004 = ~controllable_BtoR_REQ1 & ~n19003;
  assign n19005 = ~controllable_BtoR_REQ0 & ~n19004;
  assign n19006 = ~n14824 & ~n19005;
  assign n19007 = ~i_RtoB_ACK0 & ~n19006;
  assign n19008 = ~n16751 & ~n19007;
  assign n19009 = controllable_DEQ & ~n19008;
  assign n19010 = ~controllable_BtoR_REQ1 & ~n8990;
  assign n19011 = ~controllable_BtoR_REQ1 & ~n19010;
  assign n19012 = ~controllable_BtoR_REQ0 & ~n19011;
  assign n19013 = ~n14841 & ~n19012;
  assign n19014 = ~i_RtoB_ACK0 & ~n19013;
  assign n19015 = ~n16755 & ~n19014;
  assign n19016 = ~controllable_DEQ & ~n19015;
  assign n19017 = ~n19009 & ~n19016;
  assign n19018 = i_FULL & ~n19017;
  assign n19019 = ~n14824 & ~n18950;
  assign n19020 = ~i_RtoB_ACK0 & ~n19019;
  assign n19021 = ~n16751 & ~n19020;
  assign n19022 = controllable_DEQ & ~n19021;
  assign n19023 = ~n8883 & ~n8974;
  assign n19024 = ~controllable_BtoR_REQ1 & ~n19023;
  assign n19025 = ~controllable_BtoR_REQ1 & ~n19024;
  assign n19026 = ~controllable_BtoR_REQ0 & ~n19025;
  assign n19027 = ~n14841 & ~n19026;
  assign n19028 = ~i_RtoB_ACK0 & ~n19027;
  assign n19029 = ~n16755 & ~n19028;
  assign n19030 = ~controllable_DEQ & ~n19029;
  assign n19031 = ~n19022 & ~n19030;
  assign n19032 = ~i_FULL & ~n19031;
  assign n19033 = ~n19018 & ~n19032;
  assign n19034 = i_nEMPTY & ~n19033;
  assign n19035 = ~n14850 & ~n18967;
  assign n19036 = ~i_RtoB_ACK0 & ~n19035;
  assign n19037 = ~i_RtoB_ACK0 & ~n19036;
  assign n19038 = controllable_DEQ & ~n19037;
  assign n19039 = ~controllable_BtoR_REQ1 & ~n9027;
  assign n19040 = ~controllable_BtoR_REQ1 & ~n19039;
  assign n19041 = ~controllable_BtoR_REQ0 & ~n19040;
  assign n19042 = ~n14860 & ~n19041;
  assign n19043 = ~i_RtoB_ACK0 & ~n19042;
  assign n19044 = ~n16751 & ~n19043;
  assign n19045 = ~controllable_DEQ & ~n19044;
  assign n19046 = ~n19038 & ~n19045;
  assign n19047 = i_FULL & ~n19046;
  assign n19048 = ~n14869 & ~n18981;
  assign n19049 = ~i_RtoB_ACK0 & ~n19048;
  assign n19050 = ~i_RtoB_ACK0 & ~n19049;
  assign n19051 = controllable_DEQ & ~n19050;
  assign n19052 = ~n8861 & ~n9044;
  assign n19053 = ~controllable_BtoR_REQ1 & ~n19052;
  assign n19054 = ~controllable_BtoR_REQ1 & ~n19053;
  assign n19055 = ~controllable_BtoR_REQ0 & ~n19054;
  assign n19056 = ~n14824 & ~n19055;
  assign n19057 = ~i_RtoB_ACK0 & ~n19056;
  assign n19058 = ~n16751 & ~n19057;
  assign n19059 = ~controllable_DEQ & ~n19058;
  assign n19060 = ~n19051 & ~n19059;
  assign n19061 = ~i_FULL & ~n19060;
  assign n19062 = ~n19047 & ~n19061;
  assign n19063 = ~i_nEMPTY & ~n19062;
  assign n19064 = ~n19034 & ~n19063;
  assign n19065 = ~controllable_BtoS_ACK0 & ~n19064;
  assign n19066 = ~n14811 & ~n19065;
  assign n19067 = ~n4465 & ~n19066;
  assign n19068 = ~n19001 & ~n19067;
  assign n19069 = i_StoB_REQ10 & ~n19068;
  assign n19070 = ~i_RtoB_ACK1 & ~n9303;
  assign n19071 = ~n5859 & ~n19070;
  assign n19072 = ~controllable_BtoR_REQ1 & ~n19071;
  assign n19073 = ~controllable_BtoR_REQ1 & ~n19072;
  assign n19074 = controllable_BtoR_REQ0 & ~n19073;
  assign n19075 = ~n14897 & ~n19074;
  assign n19076 = i_RtoB_ACK0 & ~n19075;
  assign n19077 = ~n9501 & ~n13284;
  assign n19078 = ~controllable_BtoR_REQ1 & ~n19077;
  assign n19079 = ~controllable_BtoR_REQ1 & ~n19078;
  assign n19080 = ~controllable_BtoR_REQ0 & ~n19079;
  assign n19081 = ~n14904 & ~n19080;
  assign n19082 = ~i_RtoB_ACK0 & ~n19081;
  assign n19083 = ~n19076 & ~n19082;
  assign n19084 = controllable_DEQ & ~n19083;
  assign n19085 = ~n6785 & ~n9813;
  assign n19086 = ~controllable_BtoR_REQ1 & ~n19085;
  assign n19087 = ~controllable_BtoR_REQ1 & ~n19086;
  assign n19088 = controllable_BtoR_REQ0 & ~n19087;
  assign n19089 = ~n14916 & ~n19088;
  assign n19090 = i_RtoB_ACK0 & ~n19089;
  assign n19091 = ~n9520 & ~n13253;
  assign n19092 = ~controllable_BtoR_REQ1 & ~n19091;
  assign n19093 = ~controllable_BtoR_REQ1 & ~n19092;
  assign n19094 = ~controllable_BtoR_REQ0 & ~n19093;
  assign n19095 = ~n14923 & ~n19094;
  assign n19096 = ~i_RtoB_ACK0 & ~n19095;
  assign n19097 = ~n19090 & ~n19096;
  assign n19098 = ~controllable_DEQ & ~n19097;
  assign n19099 = ~n19084 & ~n19098;
  assign n19100 = i_FULL & ~n19099;
  assign n19101 = ~n9534 & ~n13284;
  assign n19102 = ~controllable_BtoR_REQ1 & ~n19101;
  assign n19103 = ~controllable_BtoR_REQ1 & ~n19102;
  assign n19104 = ~controllable_BtoR_REQ0 & ~n19103;
  assign n19105 = ~n14942 & ~n19104;
  assign n19106 = ~i_RtoB_ACK0 & ~n19105;
  assign n19107 = ~n19076 & ~n19106;
  assign n19108 = controllable_DEQ & ~n19107;
  assign n19109 = ~n9547 & ~n13253;
  assign n19110 = ~controllable_BtoR_REQ1 & ~n19109;
  assign n19111 = ~controllable_BtoR_REQ1 & ~n19110;
  assign n19112 = ~controllable_BtoR_REQ0 & ~n19111;
  assign n19113 = ~n14958 & ~n19112;
  assign n19114 = ~i_RtoB_ACK0 & ~n19113;
  assign n19115 = ~n19090 & ~n19114;
  assign n19116 = ~controllable_DEQ & ~n19115;
  assign n19117 = ~n19108 & ~n19116;
  assign n19118 = ~i_FULL & ~n19117;
  assign n19119 = ~n19100 & ~n19118;
  assign n19120 = i_nEMPTY & ~n19119;
  assign n19121 = ~controllable_BtoR_REQ1 & ~n9563;
  assign n19122 = ~controllable_BtoR_REQ0 & ~n19121;
  assign n19123 = ~n14979 & ~n19122;
  assign n19124 = ~i_RtoB_ACK0 & ~n19123;
  assign n19125 = ~n14975 & ~n19124;
  assign n19126 = controllable_DEQ & ~n19125;
  assign n19127 = ~n5859 & ~n9836;
  assign n19128 = ~controllable_BtoR_REQ1 & ~n19127;
  assign n19129 = ~controllable_BtoR_REQ1 & ~n19128;
  assign n19130 = controllable_BtoR_REQ0 & ~n19129;
  assign n19131 = ~n14897 & ~n19130;
  assign n19132 = i_RtoB_ACK0 & ~n19131;
  assign n19133 = ~n9575 & ~n13284;
  assign n19134 = ~controllable_BtoR_REQ1 & ~n19133;
  assign n19135 = ~controllable_BtoR_REQ1 & ~n19134;
  assign n19136 = ~controllable_BtoR_REQ0 & ~n19135;
  assign n19137 = ~n14995 & ~n19136;
  assign n19138 = ~i_RtoB_ACK0 & ~n19137;
  assign n19139 = ~n19132 & ~n19138;
  assign n19140 = ~controllable_DEQ & ~n19139;
  assign n19141 = ~n19126 & ~n19140;
  assign n19142 = i_FULL & ~n19141;
  assign n19143 = ~controllable_BtoR_REQ1 & ~n9587;
  assign n19144 = ~controllable_BtoR_REQ0 & ~n19143;
  assign n19145 = ~n15014 & ~n19144;
  assign n19146 = ~i_RtoB_ACK0 & ~n19145;
  assign n19147 = ~n15010 & ~n19146;
  assign n19148 = controllable_DEQ & ~n19147;
  assign n19149 = ~n9599 & ~n13284;
  assign n19150 = ~controllable_BtoR_REQ1 & ~n19149;
  assign n19151 = ~controllable_BtoR_REQ1 & ~n19150;
  assign n19152 = ~controllable_BtoR_REQ0 & ~n19151;
  assign n19153 = ~n14904 & ~n19152;
  assign n19154 = ~i_RtoB_ACK0 & ~n19153;
  assign n19155 = ~n19076 & ~n19154;
  assign n19156 = ~controllable_DEQ & ~n19155;
  assign n19157 = ~n19148 & ~n19156;
  assign n19158 = ~i_FULL & ~n19157;
  assign n19159 = ~n19142 & ~n19158;
  assign n19160 = ~i_nEMPTY & ~n19159;
  assign n19161 = ~n19120 & ~n19160;
  assign n19162 = controllable_BtoS_ACK0 & ~n19161;
  assign n19163 = ~i_RtoB_ACK1 & ~n9636;
  assign n19164 = ~n6897 & ~n19163;
  assign n19165 = ~controllable_BtoR_REQ1 & ~n19164;
  assign n19166 = ~controllable_BtoR_REQ1 & ~n19165;
  assign n19167 = controllable_BtoR_REQ0 & ~n19166;
  assign n19168 = ~n15039 & ~n19167;
  assign n19169 = i_RtoB_ACK0 & ~n19168;
  assign n19170 = ~n9648 & ~n13348;
  assign n19171 = ~controllable_BtoR_REQ1 & ~n19170;
  assign n19172 = ~controllable_BtoR_REQ1 & ~n19171;
  assign n19173 = ~controllable_BtoR_REQ0 & ~n19172;
  assign n19174 = ~n15046 & ~n19173;
  assign n19175 = ~i_RtoB_ACK0 & ~n19174;
  assign n19176 = ~n19169 & ~n19175;
  assign n19177 = controllable_DEQ & ~n19176;
  assign n19178 = ~n6951 & ~n9904;
  assign n19179 = ~controllable_BtoR_REQ1 & ~n19178;
  assign n19180 = ~controllable_BtoR_REQ1 & ~n19179;
  assign n19181 = controllable_BtoR_REQ0 & ~n19180;
  assign n19182 = ~n15058 & ~n19181;
  assign n19183 = i_RtoB_ACK0 & ~n19182;
  assign n19184 = ~n9667 & ~n13317;
  assign n19185 = ~controllable_BtoR_REQ1 & ~n19184;
  assign n19186 = ~controllable_BtoR_REQ1 & ~n19185;
  assign n19187 = ~controllable_BtoR_REQ0 & ~n19186;
  assign n19188 = ~n15065 & ~n19187;
  assign n19189 = ~i_RtoB_ACK0 & ~n19188;
  assign n19190 = ~n19183 & ~n19189;
  assign n19191 = ~controllable_DEQ & ~n19190;
  assign n19192 = ~n19177 & ~n19191;
  assign n19193 = i_FULL & ~n19192;
  assign n19194 = ~n9681 & ~n13348;
  assign n19195 = ~controllable_BtoR_REQ1 & ~n19194;
  assign n19196 = ~controllable_BtoR_REQ1 & ~n19195;
  assign n19197 = ~controllable_BtoR_REQ0 & ~n19196;
  assign n19198 = ~n15084 & ~n19197;
  assign n19199 = ~i_RtoB_ACK0 & ~n19198;
  assign n19200 = ~n19169 & ~n19199;
  assign n19201 = controllable_DEQ & ~n19200;
  assign n19202 = ~n9694 & ~n13317;
  assign n19203 = ~controllable_BtoR_REQ1 & ~n19202;
  assign n19204 = ~controllable_BtoR_REQ1 & ~n19203;
  assign n19205 = ~controllable_BtoR_REQ0 & ~n19204;
  assign n19206 = ~n15100 & ~n19205;
  assign n19207 = ~i_RtoB_ACK0 & ~n19206;
  assign n19208 = ~n19183 & ~n19207;
  assign n19209 = ~controllable_DEQ & ~n19208;
  assign n19210 = ~n19201 & ~n19209;
  assign n19211 = ~i_FULL & ~n19210;
  assign n19212 = ~n19193 & ~n19211;
  assign n19213 = i_nEMPTY & ~n19212;
  assign n19214 = ~controllable_BtoR_REQ1 & ~n9710;
  assign n19215 = ~controllable_BtoR_REQ0 & ~n19214;
  assign n19216 = ~n15121 & ~n19215;
  assign n19217 = ~i_RtoB_ACK0 & ~n19216;
  assign n19218 = ~n15117 & ~n19217;
  assign n19219 = controllable_DEQ & ~n19218;
  assign n19220 = ~n6897 & ~n9871;
  assign n19221 = ~controllable_BtoR_REQ1 & ~n19220;
  assign n19222 = ~controllable_BtoR_REQ1 & ~n19221;
  assign n19223 = controllable_BtoR_REQ0 & ~n19222;
  assign n19224 = ~n15039 & ~n19223;
  assign n19225 = i_RtoB_ACK0 & ~n19224;
  assign n19226 = ~n9722 & ~n13348;
  assign n19227 = ~controllable_BtoR_REQ1 & ~n19226;
  assign n19228 = ~controllable_BtoR_REQ1 & ~n19227;
  assign n19229 = ~controllable_BtoR_REQ0 & ~n19228;
  assign n19230 = ~n15137 & ~n19229;
  assign n19231 = ~i_RtoB_ACK0 & ~n19230;
  assign n19232 = ~n19225 & ~n19231;
  assign n19233 = ~controllable_DEQ & ~n19232;
  assign n19234 = ~n19219 & ~n19233;
  assign n19235 = i_FULL & ~n19234;
  assign n19236 = ~controllable_BtoR_REQ1 & ~n9734;
  assign n19237 = ~controllable_BtoR_REQ0 & ~n19236;
  assign n19238 = ~n15156 & ~n19237;
  assign n19239 = ~i_RtoB_ACK0 & ~n19238;
  assign n19240 = ~n15152 & ~n19239;
  assign n19241 = controllable_DEQ & ~n19240;
  assign n19242 = ~n9749 & ~n13348;
  assign n19243 = ~controllable_BtoR_REQ1 & ~n19242;
  assign n19244 = ~controllable_BtoR_REQ1 & ~n19243;
  assign n19245 = ~controllable_BtoR_REQ0 & ~n19244;
  assign n19246 = ~n15046 & ~n19245;
  assign n19247 = ~i_RtoB_ACK0 & ~n19246;
  assign n19248 = ~n19169 & ~n19247;
  assign n19249 = ~controllable_DEQ & ~n19248;
  assign n19250 = ~n19241 & ~n19249;
  assign n19251 = ~i_FULL & ~n19250;
  assign n19252 = ~n19235 & ~n19251;
  assign n19253 = ~i_nEMPTY & ~n19252;
  assign n19254 = ~n19213 & ~n19253;
  assign n19255 = ~controllable_BtoS_ACK0 & ~n19254;
  assign n19256 = ~n19162 & ~n19255;
  assign n19257 = n4465 & ~n19256;
  assign n19258 = ~n9794 & ~n13394;
  assign n19259 = ~controllable_BtoR_REQ1 & ~n19258;
  assign n19260 = ~controllable_BtoR_REQ1 & ~n19259;
  assign n19261 = ~controllable_BtoR_REQ0 & ~n19260;
  assign n19262 = ~n15190 & ~n19261;
  assign n19263 = ~i_RtoB_ACK0 & ~n19262;
  assign n19264 = ~n18661 & ~n19263;
  assign n19265 = controllable_DEQ & ~n19264;
  assign n19266 = ~n9813 & ~n13383;
  assign n19267 = ~controllable_BtoR_REQ1 & ~n19266;
  assign n19268 = ~controllable_BtoR_REQ1 & ~n19267;
  assign n19269 = ~controllable_BtoR_REQ0 & ~n19268;
  assign n19270 = ~n15209 & ~n19269;
  assign n19271 = ~i_RtoB_ACK0 & ~n19270;
  assign n19272 = ~n18665 & ~n19271;
  assign n19273 = ~controllable_DEQ & ~n19272;
  assign n19274 = ~n19265 & ~n19273;
  assign n19275 = i_nEMPTY & ~n19274;
  assign n19276 = ~controllable_BtoR_REQ1 & ~n9827;
  assign n19277 = ~controllable_BtoR_REQ0 & ~n19276;
  assign n19278 = ~n15221 & ~n19277;
  assign n19279 = ~i_RtoB_ACK0 & ~n19278;
  assign n19280 = ~n15217 & ~n19279;
  assign n19281 = controllable_DEQ & ~n19280;
  assign n19282 = ~n9836 & ~n13394;
  assign n19283 = ~controllable_BtoR_REQ1 & ~n19282;
  assign n19284 = ~controllable_BtoR_REQ1 & ~n19283;
  assign n19285 = ~controllable_BtoR_REQ0 & ~n19284;
  assign n19286 = ~n15237 & ~n19285;
  assign n19287 = ~i_RtoB_ACK0 & ~n19286;
  assign n19288 = ~n18671 & ~n19287;
  assign n19289 = ~controllable_DEQ & ~n19288;
  assign n19290 = ~n19281 & ~n19289;
  assign n19291 = i_FULL & ~n19290;
  assign n19292 = ~controllable_BtoR_REQ1 & ~n9848;
  assign n19293 = ~controllable_BtoR_REQ0 & ~n19292;
  assign n19294 = ~n15249 & ~n19293;
  assign n19295 = ~i_RtoB_ACK0 & ~n19294;
  assign n19296 = ~n15245 & ~n19295;
  assign n19297 = controllable_DEQ & ~n19296;
  assign n19298 = ~n9856 & ~n13394;
  assign n19299 = ~controllable_BtoR_REQ1 & ~n19298;
  assign n19300 = ~controllable_BtoR_REQ1 & ~n19299;
  assign n19301 = ~controllable_BtoR_REQ0 & ~n19300;
  assign n19302 = ~n15190 & ~n19301;
  assign n19303 = ~i_RtoB_ACK0 & ~n19302;
  assign n19304 = ~n18661 & ~n19303;
  assign n19305 = ~controllable_DEQ & ~n19304;
  assign n19306 = ~n19297 & ~n19305;
  assign n19307 = ~i_FULL & ~n19306;
  assign n19308 = ~n19291 & ~n19307;
  assign n19309 = ~i_nEMPTY & ~n19308;
  assign n19310 = ~n19275 & ~n19309;
  assign n19311 = controllable_BtoS_ACK0 & ~n19310;
  assign n19312 = ~n9718 & ~n9895;
  assign n19313 = ~controllable_BtoR_REQ1 & ~n19312;
  assign n19314 = ~controllable_BtoR_REQ1 & ~n19313;
  assign n19315 = ~controllable_BtoR_REQ0 & ~n19314;
  assign n19316 = ~n15281 & ~n19315;
  assign n19317 = ~i_RtoB_ACK0 & ~n19316;
  assign n19318 = ~n16911 & ~n19317;
  assign n19319 = controllable_DEQ & ~n19318;
  assign n19320 = ~n9664 & ~n9913;
  assign n19321 = ~controllable_BtoR_REQ1 & ~n19320;
  assign n19322 = ~controllable_BtoR_REQ1 & ~n19321;
  assign n19323 = ~controllable_BtoR_REQ0 & ~n19322;
  assign n19324 = ~n15300 & ~n19323;
  assign n19325 = ~i_RtoB_ACK0 & ~n19324;
  assign n19326 = ~n16919 & ~n19325;
  assign n19327 = ~controllable_DEQ & ~n19326;
  assign n19328 = ~n19319 & ~n19327;
  assign n19329 = i_FULL & ~n19328;
  assign n19330 = ~n15319 & ~n17701;
  assign n19331 = ~i_RtoB_ACK0 & ~n19330;
  assign n19332 = ~n16911 & ~n19331;
  assign n19333 = controllable_DEQ & ~n19332;
  assign n19334 = ~n9664 & ~n9895;
  assign n19335 = ~controllable_BtoR_REQ1 & ~n19334;
  assign n19336 = ~controllable_BtoR_REQ1 & ~n19335;
  assign n19337 = ~controllable_BtoR_REQ0 & ~n19336;
  assign n19338 = ~n15335 & ~n19337;
  assign n19339 = ~i_RtoB_ACK0 & ~n19338;
  assign n19340 = ~n16919 & ~n19339;
  assign n19341 = ~controllable_DEQ & ~n19340;
  assign n19342 = ~n19333 & ~n19341;
  assign n19343 = ~i_FULL & ~n19342;
  assign n19344 = ~n19329 & ~n19343;
  assign n19345 = i_nEMPTY & ~n19344;
  assign n19346 = ~n15356 & ~n17737;
  assign n19347 = ~i_RtoB_ACK0 & ~n19346;
  assign n19348 = ~n15352 & ~n19347;
  assign n19349 = controllable_DEQ & ~n19348;
  assign n19350 = ~n9718 & ~n9961;
  assign n19351 = ~controllable_BtoR_REQ1 & ~n19350;
  assign n19352 = ~controllable_BtoR_REQ1 & ~n19351;
  assign n19353 = ~controllable_BtoR_REQ0 & ~n19352;
  assign n19354 = ~n15372 & ~n19353;
  assign n19355 = ~i_RtoB_ACK0 & ~n19354;
  assign n19356 = ~n16937 & ~n19355;
  assign n19357 = ~controllable_DEQ & ~n19356;
  assign n19358 = ~n19349 & ~n19357;
  assign n19359 = i_FULL & ~n19358;
  assign n19360 = ~n15391 & ~n17770;
  assign n19361 = ~i_RtoB_ACK0 & ~n19360;
  assign n19362 = ~n15387 & ~n19361;
  assign n19363 = controllable_DEQ & ~n19362;
  assign n19364 = ~n9718 & ~n9981;
  assign n19365 = ~controllable_BtoR_REQ1 & ~n19364;
  assign n19366 = ~controllable_BtoR_REQ1 & ~n19365;
  assign n19367 = ~controllable_BtoR_REQ0 & ~n19366;
  assign n19368 = ~n15281 & ~n19367;
  assign n19369 = ~i_RtoB_ACK0 & ~n19368;
  assign n19370 = ~n16911 & ~n19369;
  assign n19371 = ~controllable_DEQ & ~n19370;
  assign n19372 = ~n19363 & ~n19371;
  assign n19373 = ~i_FULL & ~n19372;
  assign n19374 = ~n19359 & ~n19373;
  assign n19375 = ~i_nEMPTY & ~n19374;
  assign n19376 = ~n19345 & ~n19375;
  assign n19377 = ~controllable_BtoS_ACK0 & ~n19376;
  assign n19378 = ~n19311 & ~n19377;
  assign n19379 = ~n4465 & ~n19378;
  assign n19380 = ~n19257 & ~n19379;
  assign n19381 = ~i_StoB_REQ10 & ~n19380;
  assign n19382 = ~n19069 & ~n19381;
  assign n19383 = controllable_BtoS_ACK10 & ~n19382;
  assign n19384 = controllable_BtoR_REQ0 & ~n14905;
  assign n19385 = ~n9547 & ~n9571;
  assign n19386 = ~controllable_BtoR_REQ1 & ~n19385;
  assign n19387 = ~controllable_BtoR_REQ1 & ~n19386;
  assign n19388 = ~controllable_BtoR_REQ0 & ~n19387;
  assign n19389 = ~n19384 & ~n19388;
  assign n19390 = ~i_RtoB_ACK0 & ~n19389;
  assign n19391 = ~n16962 & ~n19390;
  assign n19392 = controllable_DEQ & ~n19391;
  assign n19393 = controllable_BtoR_REQ0 & ~n14924;
  assign n19394 = ~n9517 & ~n9520;
  assign n19395 = ~controllable_BtoR_REQ1 & ~n19394;
  assign n19396 = ~controllable_BtoR_REQ1 & ~n19395;
  assign n19397 = ~controllable_BtoR_REQ0 & ~n19396;
  assign n19398 = ~n19393 & ~n19397;
  assign n19399 = ~i_RtoB_ACK0 & ~n19398;
  assign n19400 = ~n16970 & ~n19399;
  assign n19401 = ~controllable_DEQ & ~n19400;
  assign n19402 = ~n19392 & ~n19401;
  assign n19403 = i_FULL & ~n19402;
  assign n19404 = controllable_BtoR_REQ0 & ~n14943;
  assign n19405 = ~n17622 & ~n19404;
  assign n19406 = ~i_RtoB_ACK0 & ~n19405;
  assign n19407 = ~n16962 & ~n19406;
  assign n19408 = controllable_DEQ & ~n19407;
  assign n19409 = controllable_BtoR_REQ0 & ~n14959;
  assign n19410 = ~n9517 & ~n9547;
  assign n19411 = ~controllable_BtoR_REQ1 & ~n19410;
  assign n19412 = ~controllable_BtoR_REQ1 & ~n19411;
  assign n19413 = ~controllable_BtoR_REQ0 & ~n19412;
  assign n19414 = ~n19409 & ~n19413;
  assign n19415 = ~i_RtoB_ACK0 & ~n19414;
  assign n19416 = ~n16970 & ~n19415;
  assign n19417 = ~controllable_DEQ & ~n19416;
  assign n19418 = ~n19408 & ~n19417;
  assign n19419 = ~i_FULL & ~n19418;
  assign n19420 = ~n19403 & ~n19419;
  assign n19421 = i_nEMPTY & ~n19420;
  assign n19422 = controllable_BtoR_REQ0 & ~n14980;
  assign n19423 = ~n17647 & ~n19422;
  assign n19424 = ~i_RtoB_ACK0 & ~n19423;
  assign n19425 = ~n15466 & ~n19424;
  assign n19426 = controllable_DEQ & ~n19425;
  assign n19427 = controllable_BtoR_REQ0 & ~n14996;
  assign n19428 = ~n9571 & ~n9575;
  assign n19429 = ~controllable_BtoR_REQ1 & ~n19428;
  assign n19430 = ~controllable_BtoR_REQ1 & ~n19429;
  assign n19431 = ~controllable_BtoR_REQ0 & ~n19430;
  assign n19432 = ~n19427 & ~n19431;
  assign n19433 = ~i_RtoB_ACK0 & ~n19432;
  assign n19434 = ~n16988 & ~n19433;
  assign n19435 = ~controllable_DEQ & ~n19434;
  assign n19436 = ~n19426 & ~n19435;
  assign n19437 = i_FULL & ~n19436;
  assign n19438 = controllable_BtoR_REQ0 & ~n15015;
  assign n19439 = ~n17669 & ~n19438;
  assign n19440 = ~i_RtoB_ACK0 & ~n19439;
  assign n19441 = ~n15487 & ~n19440;
  assign n19442 = controllable_DEQ & ~n19441;
  assign n19443 = ~controllable_DEQ & ~n19391;
  assign n19444 = ~n19442 & ~n19443;
  assign n19445 = ~i_FULL & ~n19444;
  assign n19446 = ~n19437 & ~n19445;
  assign n19447 = ~i_nEMPTY & ~n19446;
  assign n19448 = ~n19421 & ~n19447;
  assign n19449 = controllable_BtoS_ACK0 & ~n19448;
  assign n19450 = controllable_BtoR_REQ0 & ~n15047;
  assign n19451 = ~n9694 & ~n9718;
  assign n19452 = ~controllable_BtoR_REQ1 & ~n19451;
  assign n19453 = ~controllable_BtoR_REQ1 & ~n19452;
  assign n19454 = ~controllable_BtoR_REQ0 & ~n19453;
  assign n19455 = ~n19450 & ~n19454;
  assign n19456 = ~i_RtoB_ACK0 & ~n19455;
  assign n19457 = ~n17006 & ~n19456;
  assign n19458 = controllable_DEQ & ~n19457;
  assign n19459 = controllable_BtoR_REQ0 & ~n15066;
  assign n19460 = ~n9664 & ~n9667;
  assign n19461 = ~controllable_BtoR_REQ1 & ~n19460;
  assign n19462 = ~controllable_BtoR_REQ1 & ~n19461;
  assign n19463 = ~controllable_BtoR_REQ0 & ~n19462;
  assign n19464 = ~n19459 & ~n19463;
  assign n19465 = ~i_RtoB_ACK0 & ~n19464;
  assign n19466 = ~n17014 & ~n19465;
  assign n19467 = ~controllable_DEQ & ~n19466;
  assign n19468 = ~n19458 & ~n19467;
  assign n19469 = i_FULL & ~n19468;
  assign n19470 = controllable_BtoR_REQ0 & ~n15085;
  assign n19471 = ~n17701 & ~n19470;
  assign n19472 = ~i_RtoB_ACK0 & ~n19471;
  assign n19473 = ~n17006 & ~n19472;
  assign n19474 = controllable_DEQ & ~n19473;
  assign n19475 = controllable_BtoR_REQ0 & ~n15101;
  assign n19476 = ~n9664 & ~n9694;
  assign n19477 = ~controllable_BtoR_REQ1 & ~n19476;
  assign n19478 = ~controllable_BtoR_REQ1 & ~n19477;
  assign n19479 = ~controllable_BtoR_REQ0 & ~n19478;
  assign n19480 = ~n19475 & ~n19479;
  assign n19481 = ~i_RtoB_ACK0 & ~n19480;
  assign n19482 = ~n17014 & ~n19481;
  assign n19483 = ~controllable_DEQ & ~n19482;
  assign n19484 = ~n19474 & ~n19483;
  assign n19485 = ~i_FULL & ~n19484;
  assign n19486 = ~n19469 & ~n19485;
  assign n19487 = i_nEMPTY & ~n19486;
  assign n19488 = controllable_BtoR_REQ0 & ~n15122;
  assign n19489 = ~n17737 & ~n19488;
  assign n19490 = ~i_RtoB_ACK0 & ~n19489;
  assign n19491 = ~n15548 & ~n19490;
  assign n19492 = controllable_DEQ & ~n19491;
  assign n19493 = controllable_BtoR_REQ0 & ~n15138;
  assign n19494 = ~n9718 & ~n9722;
  assign n19495 = ~controllable_BtoR_REQ1 & ~n19494;
  assign n19496 = ~controllable_BtoR_REQ1 & ~n19495;
  assign n19497 = ~controllable_BtoR_REQ0 & ~n19496;
  assign n19498 = ~n19493 & ~n19497;
  assign n19499 = ~i_RtoB_ACK0 & ~n19498;
  assign n19500 = ~n17032 & ~n19499;
  assign n19501 = ~controllable_DEQ & ~n19500;
  assign n19502 = ~n19492 & ~n19501;
  assign n19503 = i_FULL & ~n19502;
  assign n19504 = controllable_BtoR_REQ0 & ~n15157;
  assign n19505 = ~n17770 & ~n19504;
  assign n19506 = ~i_RtoB_ACK0 & ~n19505;
  assign n19507 = ~n15569 & ~n19506;
  assign n19508 = controllable_DEQ & ~n19507;
  assign n19509 = ~controllable_DEQ & ~n19457;
  assign n19510 = ~n19508 & ~n19509;
  assign n19511 = ~i_FULL & ~n19510;
  assign n19512 = ~n19503 & ~n19511;
  assign n19513 = ~i_nEMPTY & ~n19512;
  assign n19514 = ~n19487 & ~n19513;
  assign n19515 = ~controllable_BtoS_ACK0 & ~n19514;
  assign n19516 = ~n19449 & ~n19515;
  assign n19517 = n4465 & ~n19516;
  assign n19518 = controllable_BtoR_REQ0 & ~n15191;
  assign n19519 = ~n17622 & ~n19518;
  assign n19520 = ~i_RtoB_ACK0 & ~n19519;
  assign n19521 = ~n17052 & ~n19520;
  assign n19522 = controllable_DEQ & ~n19521;
  assign n19523 = controllable_BtoR_REQ0 & ~n15201;
  assign n19524 = ~n17628 & ~n19523;
  assign n19525 = ~i_RtoB_ACK0 & ~n19524;
  assign n19526 = ~n17060 & ~n19525;
  assign n19527 = ~controllable_DEQ & ~n19526;
  assign n19528 = ~n19522 & ~n19527;
  assign n19529 = i_nEMPTY & ~n19528;
  assign n19530 = controllable_BtoR_REQ0 & ~n15222;
  assign n19531 = ~n17647 & ~n19530;
  assign n19532 = ~i_RtoB_ACK0 & ~n19531;
  assign n19533 = ~n15604 & ~n19532;
  assign n19534 = controllable_DEQ & ~n19533;
  assign n19535 = controllable_BtoR_REQ0 & ~n15182;
  assign n19536 = ~n17613 & ~n19535;
  assign n19537 = ~i_RtoB_ACK0 & ~n19536;
  assign n19538 = ~n17070 & ~n19537;
  assign n19539 = ~controllable_DEQ & ~n19538;
  assign n19540 = ~n19534 & ~n19539;
  assign n19541 = i_FULL & ~n19540;
  assign n19542 = controllable_BtoR_REQ0 & ~n15250;
  assign n19543 = ~n17669 & ~n19542;
  assign n19544 = ~i_RtoB_ACK0 & ~n19543;
  assign n19545 = ~n15619 & ~n19544;
  assign n19546 = controllable_DEQ & ~n19545;
  assign n19547 = ~controllable_DEQ & ~n19521;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = ~i_FULL & ~n19548;
  assign n19550 = ~n19541 & ~n19549;
  assign n19551 = ~i_nEMPTY & ~n19550;
  assign n19552 = ~n19529 & ~n19551;
  assign n19553 = controllable_BtoS_ACK0 & ~n19552;
  assign n19554 = controllable_BtoR_REQ0 & ~n15282;
  assign n19555 = ~n19315 & ~n19554;
  assign n19556 = ~i_RtoB_ACK0 & ~n19555;
  assign n19557 = ~n17088 & ~n19556;
  assign n19558 = controllable_DEQ & ~n19557;
  assign n19559 = controllable_BtoR_REQ0 & ~n15301;
  assign n19560 = ~n19323 & ~n19559;
  assign n19561 = ~i_RtoB_ACK0 & ~n19560;
  assign n19562 = ~n17096 & ~n19561;
  assign n19563 = ~controllable_DEQ & ~n19562;
  assign n19564 = ~n19558 & ~n19563;
  assign n19565 = i_FULL & ~n19564;
  assign n19566 = controllable_BtoR_REQ0 & ~n15320;
  assign n19567 = ~n17701 & ~n19566;
  assign n19568 = ~i_RtoB_ACK0 & ~n19567;
  assign n19569 = ~n17088 & ~n19568;
  assign n19570 = controllable_DEQ & ~n19569;
  assign n19571 = controllable_BtoR_REQ0 & ~n15336;
  assign n19572 = ~n19337 & ~n19571;
  assign n19573 = ~i_RtoB_ACK0 & ~n19572;
  assign n19574 = ~n17096 & ~n19573;
  assign n19575 = ~controllable_DEQ & ~n19574;
  assign n19576 = ~n19570 & ~n19575;
  assign n19577 = ~i_FULL & ~n19576;
  assign n19578 = ~n19565 & ~n19577;
  assign n19579 = i_nEMPTY & ~n19578;
  assign n19580 = controllable_BtoR_REQ0 & ~n15357;
  assign n19581 = ~n17737 & ~n19580;
  assign n19582 = ~i_RtoB_ACK0 & ~n19581;
  assign n19583 = ~n15680 & ~n19582;
  assign n19584 = controllable_DEQ & ~n19583;
  assign n19585 = controllable_BtoR_REQ0 & ~n15373;
  assign n19586 = ~n19353 & ~n19585;
  assign n19587 = ~i_RtoB_ACK0 & ~n19586;
  assign n19588 = ~n17114 & ~n19587;
  assign n19589 = ~controllable_DEQ & ~n19588;
  assign n19590 = ~n19584 & ~n19589;
  assign n19591 = i_FULL & ~n19590;
  assign n19592 = controllable_BtoR_REQ0 & ~n15392;
  assign n19593 = ~n17770 & ~n19592;
  assign n19594 = ~i_RtoB_ACK0 & ~n19593;
  assign n19595 = ~n15701 & ~n19594;
  assign n19596 = controllable_DEQ & ~n19595;
  assign n19597 = ~controllable_DEQ & ~n19557;
  assign n19598 = ~n19596 & ~n19597;
  assign n19599 = ~i_FULL & ~n19598;
  assign n19600 = ~n19591 & ~n19599;
  assign n19601 = ~i_nEMPTY & ~n19600;
  assign n19602 = ~n19579 & ~n19601;
  assign n19603 = ~controllable_BtoS_ACK0 & ~n19602;
  assign n19604 = ~n19553 & ~n19603;
  assign n19605 = ~n4465 & ~n19604;
  assign n19606 = ~n19517 & ~n19605;
  assign n19607 = i_StoB_REQ10 & ~n19606;
  assign n19608 = ~n19381 & ~n19607;
  assign n19609 = ~controllable_BtoS_ACK10 & ~n19608;
  assign n19610 = ~n19383 & ~n19609;
  assign n19611 = n4464 & ~n19610;
  assign n19612 = ~n5237 & ~n10267;
  assign n19613 = ~controllable_BtoR_REQ1 & ~n19612;
  assign n19614 = ~controllable_BtoR_REQ1 & ~n19613;
  assign n19615 = ~controllable_BtoR_REQ0 & ~n19614;
  assign n19616 = ~n15732 & ~n19615;
  assign n19617 = ~i_RtoB_ACK0 & ~n19616;
  assign n19618 = ~n17135 & ~n19617;
  assign n19619 = controllable_DEQ & ~n19618;
  assign n19620 = ~controllable_BtoR_REQ1 & ~n10283;
  assign n19621 = ~controllable_BtoR_REQ1 & ~n19620;
  assign n19622 = ~controllable_BtoR_REQ0 & ~n19621;
  assign n19623 = ~n15749 & ~n19622;
  assign n19624 = ~i_RtoB_ACK0 & ~n19623;
  assign n19625 = ~n17139 & ~n19624;
  assign n19626 = ~controllable_DEQ & ~n19625;
  assign n19627 = ~n19619 & ~n19626;
  assign n19628 = i_FULL & ~n19627;
  assign n19629 = ~n14751 & ~n15732;
  assign n19630 = ~i_RtoB_ACK0 & ~n19629;
  assign n19631 = ~n17135 & ~n19630;
  assign n19632 = controllable_DEQ & ~n19631;
  assign n19633 = ~n7563 & ~n10267;
  assign n19634 = ~controllable_BtoR_REQ1 & ~n19633;
  assign n19635 = ~controllable_BtoR_REQ1 & ~n19634;
  assign n19636 = ~controllable_BtoR_REQ0 & ~n19635;
  assign n19637 = ~n15749 & ~n19636;
  assign n19638 = ~i_RtoB_ACK0 & ~n19637;
  assign n19639 = ~n17139 & ~n19638;
  assign n19640 = ~controllable_DEQ & ~n19639;
  assign n19641 = ~n19632 & ~n19640;
  assign n19642 = ~i_FULL & ~n19641;
  assign n19643 = ~n19628 & ~n19642;
  assign n19644 = i_nEMPTY & ~n19643;
  assign n19645 = ~n14776 & ~n15758;
  assign n19646 = ~i_RtoB_ACK0 & ~n19645;
  assign n19647 = ~i_RtoB_ACK0 & ~n19646;
  assign n19648 = controllable_DEQ & ~n19647;
  assign n19649 = ~controllable_BtoR_REQ1 & ~n10320;
  assign n19650 = ~controllable_BtoR_REQ1 & ~n19649;
  assign n19651 = ~controllable_BtoR_REQ0 & ~n19650;
  assign n19652 = ~n15768 & ~n19651;
  assign n19653 = ~i_RtoB_ACK0 & ~n19652;
  assign n19654 = ~n17135 & ~n19653;
  assign n19655 = ~controllable_DEQ & ~n19654;
  assign n19656 = ~n19648 & ~n19655;
  assign n19657 = i_FULL & ~n19656;
  assign n19658 = ~n14794 & ~n15777;
  assign n19659 = ~i_RtoB_ACK0 & ~n19658;
  assign n19660 = ~i_RtoB_ACK0 & ~n19659;
  assign n19661 = controllable_DEQ & ~n19660;
  assign n19662 = ~n5237 & ~n10337;
  assign n19663 = ~controllable_BtoR_REQ1 & ~n19662;
  assign n19664 = ~controllable_BtoR_REQ1 & ~n19663;
  assign n19665 = ~controllable_BtoR_REQ0 & ~n19664;
  assign n19666 = ~n15732 & ~n19665;
  assign n19667 = ~i_RtoB_ACK0 & ~n19666;
  assign n19668 = ~n17135 & ~n19667;
  assign n19669 = ~controllable_DEQ & ~n19668;
  assign n19670 = ~n19661 & ~n19669;
  assign n19671 = ~i_FULL & ~n19670;
  assign n19672 = ~n19657 & ~n19671;
  assign n19673 = ~i_nEMPTY & ~n19672;
  assign n19674 = ~n19644 & ~n19673;
  assign n19675 = controllable_BtoS_ACK0 & ~n19674;
  assign n19676 = ~n8861 & ~n10361;
  assign n19677 = ~controllable_BtoR_REQ1 & ~n19676;
  assign n19678 = ~controllable_BtoR_REQ1 & ~n19677;
  assign n19679 = ~controllable_BtoR_REQ0 & ~n19678;
  assign n19680 = ~n15807 & ~n19679;
  assign n19681 = ~i_RtoB_ACK0 & ~n19680;
  assign n19682 = ~n17157 & ~n19681;
  assign n19683 = controllable_DEQ & ~n19682;
  assign n19684 = ~controllable_BtoR_REQ1 & ~n10377;
  assign n19685 = ~controllable_BtoR_REQ1 & ~n19684;
  assign n19686 = ~controllable_BtoR_REQ0 & ~n19685;
  assign n19687 = ~n15824 & ~n19686;
  assign n19688 = ~i_RtoB_ACK0 & ~n19687;
  assign n19689 = ~n17161 & ~n19688;
  assign n19690 = ~controllable_DEQ & ~n19689;
  assign n19691 = ~n19683 & ~n19690;
  assign n19692 = i_FULL & ~n19691;
  assign n19693 = ~n15807 & ~n18950;
  assign n19694 = ~i_RtoB_ACK0 & ~n19693;
  assign n19695 = ~n17157 & ~n19694;
  assign n19696 = controllable_DEQ & ~n19695;
  assign n19697 = ~n8883 & ~n10361;
  assign n19698 = ~controllable_BtoR_REQ1 & ~n19697;
  assign n19699 = ~controllable_BtoR_REQ1 & ~n19698;
  assign n19700 = ~controllable_BtoR_REQ0 & ~n19699;
  assign n19701 = ~n15824 & ~n19700;
  assign n19702 = ~i_RtoB_ACK0 & ~n19701;
  assign n19703 = ~n17161 & ~n19702;
  assign n19704 = ~controllable_DEQ & ~n19703;
  assign n19705 = ~n19696 & ~n19704;
  assign n19706 = ~i_FULL & ~n19705;
  assign n19707 = ~n19692 & ~n19706;
  assign n19708 = i_nEMPTY & ~n19707;
  assign n19709 = ~n15833 & ~n18967;
  assign n19710 = ~i_RtoB_ACK0 & ~n19709;
  assign n19711 = ~i_RtoB_ACK0 & ~n19710;
  assign n19712 = controllable_DEQ & ~n19711;
  assign n19713 = ~controllable_BtoR_REQ1 & ~n10414;
  assign n19714 = ~controllable_BtoR_REQ1 & ~n19713;
  assign n19715 = ~controllable_BtoR_REQ0 & ~n19714;
  assign n19716 = ~n15843 & ~n19715;
  assign n19717 = ~i_RtoB_ACK0 & ~n19716;
  assign n19718 = ~n17157 & ~n19717;
  assign n19719 = ~controllable_DEQ & ~n19718;
  assign n19720 = ~n19712 & ~n19719;
  assign n19721 = i_FULL & ~n19720;
  assign n19722 = ~n15852 & ~n18981;
  assign n19723 = ~i_RtoB_ACK0 & ~n19722;
  assign n19724 = ~i_RtoB_ACK0 & ~n19723;
  assign n19725 = controllable_DEQ & ~n19724;
  assign n19726 = ~n8861 & ~n10431;
  assign n19727 = ~controllable_BtoR_REQ1 & ~n19726;
  assign n19728 = ~controllable_BtoR_REQ1 & ~n19727;
  assign n19729 = ~controllable_BtoR_REQ0 & ~n19728;
  assign n19730 = ~n15807 & ~n19729;
  assign n19731 = ~i_RtoB_ACK0 & ~n19730;
  assign n19732 = ~n17157 & ~n19731;
  assign n19733 = ~controllable_DEQ & ~n19732;
  assign n19734 = ~n19725 & ~n19733;
  assign n19735 = ~i_FULL & ~n19734;
  assign n19736 = ~n19721 & ~n19735;
  assign n19737 = ~i_nEMPTY & ~n19736;
  assign n19738 = ~n19708 & ~n19737;
  assign n19739 = ~controllable_BtoS_ACK0 & ~n19738;
  assign n19740 = ~n19675 & ~n19739;
  assign n19741 = n4465 & ~n19740;
  assign n19742 = ~n14811 & ~n19739;
  assign n19743 = ~n4465 & ~n19742;
  assign n19744 = ~n19741 & ~n19743;
  assign n19745 = i_StoB_REQ10 & ~n19744;
  assign n19746 = ~n10478 & ~n13736;
  assign n19747 = ~controllable_BtoR_REQ1 & ~n19746;
  assign n19748 = ~controllable_BtoR_REQ1 & ~n19747;
  assign n19749 = ~controllable_BtoR_REQ0 & ~n19748;
  assign n19750 = ~n15889 & ~n19749;
  assign n19751 = ~i_RtoB_ACK0 & ~n19750;
  assign n19752 = ~n18768 & ~n19751;
  assign n19753 = controllable_DEQ & ~n19752;
  assign n19754 = ~n10496 & ~n13705;
  assign n19755 = ~controllable_BtoR_REQ1 & ~n19754;
  assign n19756 = ~controllable_BtoR_REQ1 & ~n19755;
  assign n19757 = ~controllable_BtoR_REQ0 & ~n19756;
  assign n19758 = ~n15908 & ~n19757;
  assign n19759 = ~i_RtoB_ACK0 & ~n19758;
  assign n19760 = ~n18776 & ~n19759;
  assign n19761 = ~controllable_DEQ & ~n19760;
  assign n19762 = ~n19753 & ~n19761;
  assign n19763 = i_FULL & ~n19762;
  assign n19764 = ~n10510 & ~n13736;
  assign n19765 = ~controllable_BtoR_REQ1 & ~n19764;
  assign n19766 = ~controllable_BtoR_REQ1 & ~n19765;
  assign n19767 = ~controllable_BtoR_REQ0 & ~n19766;
  assign n19768 = ~n15927 & ~n19767;
  assign n19769 = ~i_RtoB_ACK0 & ~n19768;
  assign n19770 = ~n18768 & ~n19769;
  assign n19771 = controllable_DEQ & ~n19770;
  assign n19772 = ~n10522 & ~n13705;
  assign n19773 = ~controllable_BtoR_REQ1 & ~n19772;
  assign n19774 = ~controllable_BtoR_REQ1 & ~n19773;
  assign n19775 = ~controllable_BtoR_REQ0 & ~n19774;
  assign n19776 = ~n15943 & ~n19775;
  assign n19777 = ~i_RtoB_ACK0 & ~n19776;
  assign n19778 = ~n18776 & ~n19777;
  assign n19779 = ~controllable_DEQ & ~n19778;
  assign n19780 = ~n19771 & ~n19779;
  assign n19781 = ~i_FULL & ~n19780;
  assign n19782 = ~n19763 & ~n19781;
  assign n19783 = i_nEMPTY & ~n19782;
  assign n19784 = ~controllable_BtoR_REQ1 & ~n10538;
  assign n19785 = ~controllable_BtoR_REQ0 & ~n19784;
  assign n19786 = ~n15964 & ~n19785;
  assign n19787 = ~i_RtoB_ACK0 & ~n19786;
  assign n19788 = ~n15960 & ~n19787;
  assign n19789 = controllable_DEQ & ~n19788;
  assign n19790 = ~n10548 & ~n13736;
  assign n19791 = ~controllable_BtoR_REQ1 & ~n19790;
  assign n19792 = ~controllable_BtoR_REQ1 & ~n19791;
  assign n19793 = ~controllable_BtoR_REQ0 & ~n19792;
  assign n19794 = ~n15980 & ~n19793;
  assign n19795 = ~i_RtoB_ACK0 & ~n19794;
  assign n19796 = ~n18794 & ~n19795;
  assign n19797 = ~controllable_DEQ & ~n19796;
  assign n19798 = ~n19789 & ~n19797;
  assign n19799 = i_FULL & ~n19798;
  assign n19800 = ~controllable_BtoR_REQ1 & ~n10560;
  assign n19801 = ~controllable_BtoR_REQ0 & ~n19800;
  assign n19802 = ~n15999 & ~n19801;
  assign n19803 = ~i_RtoB_ACK0 & ~n19802;
  assign n19804 = ~n15995 & ~n19803;
  assign n19805 = controllable_DEQ & ~n19804;
  assign n19806 = ~n10568 & ~n13736;
  assign n19807 = ~controllable_BtoR_REQ1 & ~n19806;
  assign n19808 = ~controllable_BtoR_REQ1 & ~n19807;
  assign n19809 = ~controllable_BtoR_REQ0 & ~n19808;
  assign n19810 = ~n15889 & ~n19809;
  assign n19811 = ~i_RtoB_ACK0 & ~n19810;
  assign n19812 = ~n18768 & ~n19811;
  assign n19813 = ~controllable_DEQ & ~n19812;
  assign n19814 = ~n19805 & ~n19813;
  assign n19815 = ~i_FULL & ~n19814;
  assign n19816 = ~n19799 & ~n19815;
  assign n19817 = ~i_nEMPTY & ~n19816;
  assign n19818 = ~n19783 & ~n19817;
  assign n19819 = controllable_BtoS_ACK0 & ~n19818;
  assign n19820 = ~n10605 & ~n13800;
  assign n19821 = ~controllable_BtoR_REQ1 & ~n19820;
  assign n19822 = ~controllable_BtoR_REQ1 & ~n19821;
  assign n19823 = ~controllable_BtoR_REQ0 & ~n19822;
  assign n19824 = ~n16031 & ~n19823;
  assign n19825 = ~i_RtoB_ACK0 & ~n19824;
  assign n19826 = ~n18813 & ~n19825;
  assign n19827 = controllable_DEQ & ~n19826;
  assign n19828 = ~n10623 & ~n13769;
  assign n19829 = ~controllable_BtoR_REQ1 & ~n19828;
  assign n19830 = ~controllable_BtoR_REQ1 & ~n19829;
  assign n19831 = ~controllable_BtoR_REQ0 & ~n19830;
  assign n19832 = ~n16050 & ~n19831;
  assign n19833 = ~i_RtoB_ACK0 & ~n19832;
  assign n19834 = ~n18821 & ~n19833;
  assign n19835 = ~controllable_DEQ & ~n19834;
  assign n19836 = ~n19827 & ~n19835;
  assign n19837 = i_FULL & ~n19836;
  assign n19838 = ~n10637 & ~n13800;
  assign n19839 = ~controllable_BtoR_REQ1 & ~n19838;
  assign n19840 = ~controllable_BtoR_REQ1 & ~n19839;
  assign n19841 = ~controllable_BtoR_REQ0 & ~n19840;
  assign n19842 = ~n16069 & ~n19841;
  assign n19843 = ~i_RtoB_ACK0 & ~n19842;
  assign n19844 = ~n18813 & ~n19843;
  assign n19845 = controllable_DEQ & ~n19844;
  assign n19846 = ~n10649 & ~n13769;
  assign n19847 = ~controllable_BtoR_REQ1 & ~n19846;
  assign n19848 = ~controllable_BtoR_REQ1 & ~n19847;
  assign n19849 = ~controllable_BtoR_REQ0 & ~n19848;
  assign n19850 = ~n16085 & ~n19849;
  assign n19851 = ~i_RtoB_ACK0 & ~n19850;
  assign n19852 = ~n18821 & ~n19851;
  assign n19853 = ~controllable_DEQ & ~n19852;
  assign n19854 = ~n19845 & ~n19853;
  assign n19855 = ~i_FULL & ~n19854;
  assign n19856 = ~n19837 & ~n19855;
  assign n19857 = i_nEMPTY & ~n19856;
  assign n19858 = ~controllable_BtoR_REQ1 & ~n10665;
  assign n19859 = ~controllable_BtoR_REQ0 & ~n19858;
  assign n19860 = ~n16106 & ~n19859;
  assign n19861 = ~i_RtoB_ACK0 & ~n19860;
  assign n19862 = ~n16102 & ~n19861;
  assign n19863 = controllable_DEQ & ~n19862;
  assign n19864 = ~n10675 & ~n13800;
  assign n19865 = ~controllable_BtoR_REQ1 & ~n19864;
  assign n19866 = ~controllable_BtoR_REQ1 & ~n19865;
  assign n19867 = ~controllable_BtoR_REQ0 & ~n19866;
  assign n19868 = ~n16122 & ~n19867;
  assign n19869 = ~i_RtoB_ACK0 & ~n19868;
  assign n19870 = ~n18839 & ~n19869;
  assign n19871 = ~controllable_DEQ & ~n19870;
  assign n19872 = ~n19863 & ~n19871;
  assign n19873 = i_FULL & ~n19872;
  assign n19874 = ~controllable_BtoR_REQ1 & ~n10687;
  assign n19875 = ~controllable_BtoR_REQ0 & ~n19874;
  assign n19876 = ~n16141 & ~n19875;
  assign n19877 = ~i_RtoB_ACK0 & ~n19876;
  assign n19878 = ~n16137 & ~n19877;
  assign n19879 = controllable_DEQ & ~n19878;
  assign n19880 = ~n10695 & ~n13800;
  assign n19881 = ~controllable_BtoR_REQ1 & ~n19880;
  assign n19882 = ~controllable_BtoR_REQ1 & ~n19881;
  assign n19883 = ~controllable_BtoR_REQ0 & ~n19882;
  assign n19884 = ~n16031 & ~n19883;
  assign n19885 = ~i_RtoB_ACK0 & ~n19884;
  assign n19886 = ~n18813 & ~n19885;
  assign n19887 = ~controllable_DEQ & ~n19886;
  assign n19888 = ~n19879 & ~n19887;
  assign n19889 = ~i_FULL & ~n19888;
  assign n19890 = ~n19873 & ~n19889;
  assign n19891 = ~i_nEMPTY & ~n19890;
  assign n19892 = ~n19857 & ~n19891;
  assign n19893 = ~controllable_BtoS_ACK0 & ~n19892;
  assign n19894 = ~n19819 & ~n19893;
  assign n19895 = n4465 & ~n19894;
  assign n19896 = ~n16175 & ~n17622;
  assign n19897 = ~i_RtoB_ACK0 & ~n19896;
  assign n19898 = ~n17282 & ~n19897;
  assign n19899 = controllable_DEQ & ~n19898;
  assign n19900 = ~n16194 & ~n17628;
  assign n19901 = ~i_RtoB_ACK0 & ~n19900;
  assign n19902 = ~n17290 & ~n19901;
  assign n19903 = ~controllable_DEQ & ~n19902;
  assign n19904 = ~n19899 & ~n19903;
  assign n19905 = i_nEMPTY & ~n19904;
  assign n19906 = ~n16204 & ~n17647;
  assign n19907 = ~i_RtoB_ACK0 & ~n19906;
  assign n19908 = ~n15217 & ~n19907;
  assign n19909 = controllable_DEQ & ~n19908;
  assign n19910 = ~n16220 & ~n17613;
  assign n19911 = ~i_RtoB_ACK0 & ~n19910;
  assign n19912 = ~n17300 & ~n19911;
  assign n19913 = ~controllable_DEQ & ~n19912;
  assign n19914 = ~n19909 & ~n19913;
  assign n19915 = i_FULL & ~n19914;
  assign n19916 = ~n16230 & ~n17669;
  assign n19917 = ~i_RtoB_ACK0 & ~n19916;
  assign n19918 = ~n15245 & ~n19917;
  assign n19919 = controllable_DEQ & ~n19918;
  assign n19920 = ~n16175 & ~n17675;
  assign n19921 = ~i_RtoB_ACK0 & ~n19920;
  assign n19922 = ~n17282 & ~n19921;
  assign n19923 = ~controllable_DEQ & ~n19922;
  assign n19924 = ~n19919 & ~n19923;
  assign n19925 = ~i_FULL & ~n19924;
  assign n19926 = ~n19915 & ~n19925;
  assign n19927 = ~i_nEMPTY & ~n19926;
  assign n19928 = ~n19905 & ~n19927;
  assign n19929 = controllable_BtoS_ACK0 & ~n19928;
  assign n19930 = ~n9718 & ~n10649;
  assign n19931 = ~controllable_BtoR_REQ1 & ~n19930;
  assign n19932 = ~controllable_BtoR_REQ1 & ~n19931;
  assign n19933 = ~controllable_BtoR_REQ0 & ~n19932;
  assign n19934 = ~n16262 & ~n19933;
  assign n19935 = ~i_RtoB_ACK0 & ~n19934;
  assign n19936 = ~n17319 & ~n19935;
  assign n19937 = controllable_DEQ & ~n19936;
  assign n19938 = ~n9664 & ~n10623;
  assign n19939 = ~controllable_BtoR_REQ1 & ~n19938;
  assign n19940 = ~controllable_BtoR_REQ1 & ~n19939;
  assign n19941 = ~controllable_BtoR_REQ0 & ~n19940;
  assign n19942 = ~n16281 & ~n19941;
  assign n19943 = ~i_RtoB_ACK0 & ~n19942;
  assign n19944 = ~n17327 & ~n19943;
  assign n19945 = ~controllable_DEQ & ~n19944;
  assign n19946 = ~n19937 & ~n19945;
  assign n19947 = i_FULL & ~n19946;
  assign n19948 = ~n16300 & ~n17701;
  assign n19949 = ~i_RtoB_ACK0 & ~n19948;
  assign n19950 = ~n17319 & ~n19949;
  assign n19951 = controllable_DEQ & ~n19950;
  assign n19952 = ~n9664 & ~n10649;
  assign n19953 = ~controllable_BtoR_REQ1 & ~n19952;
  assign n19954 = ~controllable_BtoR_REQ1 & ~n19953;
  assign n19955 = ~controllable_BtoR_REQ0 & ~n19954;
  assign n19956 = ~n16316 & ~n19955;
  assign n19957 = ~i_RtoB_ACK0 & ~n19956;
  assign n19958 = ~n17327 & ~n19957;
  assign n19959 = ~controllable_DEQ & ~n19958;
  assign n19960 = ~n19951 & ~n19959;
  assign n19961 = ~i_FULL & ~n19960;
  assign n19962 = ~n19947 & ~n19961;
  assign n19963 = i_nEMPTY & ~n19962;
  assign n19964 = ~n16337 & ~n17737;
  assign n19965 = ~i_RtoB_ACK0 & ~n19964;
  assign n19966 = ~n16333 & ~n19965;
  assign n19967 = controllable_DEQ & ~n19966;
  assign n19968 = ~n9718 & ~n10675;
  assign n19969 = ~controllable_BtoR_REQ1 & ~n19968;
  assign n19970 = ~controllable_BtoR_REQ1 & ~n19969;
  assign n19971 = ~controllable_BtoR_REQ0 & ~n19970;
  assign n19972 = ~n16353 & ~n19971;
  assign n19973 = ~i_RtoB_ACK0 & ~n19972;
  assign n19974 = ~n17345 & ~n19973;
  assign n19975 = ~controllable_DEQ & ~n19974;
  assign n19976 = ~n19967 & ~n19975;
  assign n19977 = i_FULL & ~n19976;
  assign n19978 = ~n16372 & ~n17770;
  assign n19979 = ~i_RtoB_ACK0 & ~n19978;
  assign n19980 = ~n16368 & ~n19979;
  assign n19981 = controllable_DEQ & ~n19980;
  assign n19982 = ~n9718 & ~n10695;
  assign n19983 = ~controllable_BtoR_REQ1 & ~n19982;
  assign n19984 = ~controllable_BtoR_REQ1 & ~n19983;
  assign n19985 = ~controllable_BtoR_REQ0 & ~n19984;
  assign n19986 = ~n16262 & ~n19985;
  assign n19987 = ~i_RtoB_ACK0 & ~n19986;
  assign n19988 = ~n17319 & ~n19987;
  assign n19989 = ~controllable_DEQ & ~n19988;
  assign n19990 = ~n19981 & ~n19989;
  assign n19991 = ~i_FULL & ~n19990;
  assign n19992 = ~n19977 & ~n19991;
  assign n19993 = ~i_nEMPTY & ~n19992;
  assign n19994 = ~n19963 & ~n19993;
  assign n19995 = ~controllable_BtoS_ACK0 & ~n19994;
  assign n19996 = ~n19929 & ~n19995;
  assign n19997 = ~n4465 & ~n19996;
  assign n19998 = ~n19895 & ~n19997;
  assign n19999 = ~i_StoB_REQ10 & ~n19998;
  assign n20000 = ~n19745 & ~n19999;
  assign n20001 = controllable_BtoS_ACK10 & ~n20000;
  assign n20002 = controllable_BtoR_REQ0 & ~n15890;
  assign n20003 = ~n9571 & ~n10522;
  assign n20004 = ~controllable_BtoR_REQ1 & ~n20003;
  assign n20005 = ~controllable_BtoR_REQ1 & ~n20004;
  assign n20006 = ~controllable_BtoR_REQ0 & ~n20005;
  assign n20007 = ~n20002 & ~n20006;
  assign n20008 = ~i_RtoB_ACK0 & ~n20007;
  assign n20009 = ~n17370 & ~n20008;
  assign n20010 = controllable_DEQ & ~n20009;
  assign n20011 = controllable_BtoR_REQ0 & ~n15909;
  assign n20012 = ~n9517 & ~n10496;
  assign n20013 = ~controllable_BtoR_REQ1 & ~n20012;
  assign n20014 = ~controllable_BtoR_REQ1 & ~n20013;
  assign n20015 = ~controllable_BtoR_REQ0 & ~n20014;
  assign n20016 = ~n20011 & ~n20015;
  assign n20017 = ~i_RtoB_ACK0 & ~n20016;
  assign n20018 = ~n17378 & ~n20017;
  assign n20019 = ~controllable_DEQ & ~n20018;
  assign n20020 = ~n20010 & ~n20019;
  assign n20021 = i_FULL & ~n20020;
  assign n20022 = controllable_BtoR_REQ0 & ~n15928;
  assign n20023 = ~n17622 & ~n20022;
  assign n20024 = ~i_RtoB_ACK0 & ~n20023;
  assign n20025 = ~n17370 & ~n20024;
  assign n20026 = controllable_DEQ & ~n20025;
  assign n20027 = controllable_BtoR_REQ0 & ~n15944;
  assign n20028 = ~n9517 & ~n10522;
  assign n20029 = ~controllable_BtoR_REQ1 & ~n20028;
  assign n20030 = ~controllable_BtoR_REQ1 & ~n20029;
  assign n20031 = ~controllable_BtoR_REQ0 & ~n20030;
  assign n20032 = ~n20027 & ~n20031;
  assign n20033 = ~i_RtoB_ACK0 & ~n20032;
  assign n20034 = ~n17378 & ~n20033;
  assign n20035 = ~controllable_DEQ & ~n20034;
  assign n20036 = ~n20026 & ~n20035;
  assign n20037 = ~i_FULL & ~n20036;
  assign n20038 = ~n20021 & ~n20037;
  assign n20039 = i_nEMPTY & ~n20038;
  assign n20040 = controllable_BtoR_REQ0 & ~n15965;
  assign n20041 = ~n17647 & ~n20040;
  assign n20042 = ~i_RtoB_ACK0 & ~n20041;
  assign n20043 = ~n16447 & ~n20042;
  assign n20044 = controllable_DEQ & ~n20043;
  assign n20045 = controllable_BtoR_REQ0 & ~n15981;
  assign n20046 = ~n9571 & ~n10548;
  assign n20047 = ~controllable_BtoR_REQ1 & ~n20046;
  assign n20048 = ~controllable_BtoR_REQ1 & ~n20047;
  assign n20049 = ~controllable_BtoR_REQ0 & ~n20048;
  assign n20050 = ~n20045 & ~n20049;
  assign n20051 = ~i_RtoB_ACK0 & ~n20050;
  assign n20052 = ~n17396 & ~n20051;
  assign n20053 = ~controllable_DEQ & ~n20052;
  assign n20054 = ~n20044 & ~n20053;
  assign n20055 = i_FULL & ~n20054;
  assign n20056 = controllable_BtoR_REQ0 & ~n16000;
  assign n20057 = ~n17669 & ~n20056;
  assign n20058 = ~i_RtoB_ACK0 & ~n20057;
  assign n20059 = ~n16468 & ~n20058;
  assign n20060 = controllable_DEQ & ~n20059;
  assign n20061 = ~controllable_DEQ & ~n20009;
  assign n20062 = ~n20060 & ~n20061;
  assign n20063 = ~i_FULL & ~n20062;
  assign n20064 = ~n20055 & ~n20063;
  assign n20065 = ~i_nEMPTY & ~n20064;
  assign n20066 = ~n20039 & ~n20065;
  assign n20067 = controllable_BtoS_ACK0 & ~n20066;
  assign n20068 = controllable_BtoR_REQ0 & ~n16032;
  assign n20069 = ~n19933 & ~n20068;
  assign n20070 = ~i_RtoB_ACK0 & ~n20069;
  assign n20071 = ~n17414 & ~n20070;
  assign n20072 = controllable_DEQ & ~n20071;
  assign n20073 = controllable_BtoR_REQ0 & ~n16051;
  assign n20074 = ~n19941 & ~n20073;
  assign n20075 = ~i_RtoB_ACK0 & ~n20074;
  assign n20076 = ~n17422 & ~n20075;
  assign n20077 = ~controllable_DEQ & ~n20076;
  assign n20078 = ~n20072 & ~n20077;
  assign n20079 = i_FULL & ~n20078;
  assign n20080 = controllable_BtoR_REQ0 & ~n16070;
  assign n20081 = ~n17701 & ~n20080;
  assign n20082 = ~i_RtoB_ACK0 & ~n20081;
  assign n20083 = ~n17414 & ~n20082;
  assign n20084 = controllable_DEQ & ~n20083;
  assign n20085 = controllable_BtoR_REQ0 & ~n16086;
  assign n20086 = ~n19955 & ~n20085;
  assign n20087 = ~i_RtoB_ACK0 & ~n20086;
  assign n20088 = ~n17422 & ~n20087;
  assign n20089 = ~controllable_DEQ & ~n20088;
  assign n20090 = ~n20084 & ~n20089;
  assign n20091 = ~i_FULL & ~n20090;
  assign n20092 = ~n20079 & ~n20091;
  assign n20093 = i_nEMPTY & ~n20092;
  assign n20094 = controllable_BtoR_REQ0 & ~n16107;
  assign n20095 = ~n17737 & ~n20094;
  assign n20096 = ~i_RtoB_ACK0 & ~n20095;
  assign n20097 = ~n16529 & ~n20096;
  assign n20098 = controllable_DEQ & ~n20097;
  assign n20099 = controllable_BtoR_REQ0 & ~n16123;
  assign n20100 = ~n19971 & ~n20099;
  assign n20101 = ~i_RtoB_ACK0 & ~n20100;
  assign n20102 = ~n17440 & ~n20101;
  assign n20103 = ~controllable_DEQ & ~n20102;
  assign n20104 = ~n20098 & ~n20103;
  assign n20105 = i_FULL & ~n20104;
  assign n20106 = controllable_BtoR_REQ0 & ~n16142;
  assign n20107 = ~n17770 & ~n20106;
  assign n20108 = ~i_RtoB_ACK0 & ~n20107;
  assign n20109 = ~n16550 & ~n20108;
  assign n20110 = controllable_DEQ & ~n20109;
  assign n20111 = ~controllable_DEQ & ~n20071;
  assign n20112 = ~n20110 & ~n20111;
  assign n20113 = ~i_FULL & ~n20112;
  assign n20114 = ~n20105 & ~n20113;
  assign n20115 = ~i_nEMPTY & ~n20114;
  assign n20116 = ~n20093 & ~n20115;
  assign n20117 = ~controllable_BtoS_ACK0 & ~n20116;
  assign n20118 = ~n20067 & ~n20117;
  assign n20119 = n4465 & ~n20118;
  assign n20120 = controllable_BtoR_REQ0 & ~n16176;
  assign n20121 = ~n17622 & ~n20120;
  assign n20122 = ~i_RtoB_ACK0 & ~n20121;
  assign n20123 = ~n17455 & ~n20122;
  assign n20124 = controllable_DEQ & ~n20123;
  assign n20125 = controllable_BtoR_REQ0 & ~n16186;
  assign n20126 = ~n17628 & ~n20125;
  assign n20127 = ~i_RtoB_ACK0 & ~n20126;
  assign n20128 = ~n17459 & ~n20127;
  assign n20129 = ~controllable_DEQ & ~n20128;
  assign n20130 = ~n20124 & ~n20129;
  assign n20131 = i_nEMPTY & ~n20130;
  assign n20132 = controllable_BtoR_REQ0 & ~n16205;
  assign n20133 = ~n17647 & ~n20132;
  assign n20134 = ~i_RtoB_ACK0 & ~n20133;
  assign n20135 = ~n15604 & ~n20134;
  assign n20136 = controllable_DEQ & ~n20135;
  assign n20137 = controllable_BtoR_REQ0 & ~n16167;
  assign n20138 = ~n17613 & ~n20137;
  assign n20139 = ~i_RtoB_ACK0 & ~n20138;
  assign n20140 = ~n17465 & ~n20139;
  assign n20141 = ~controllable_DEQ & ~n20140;
  assign n20142 = ~n20136 & ~n20141;
  assign n20143 = i_FULL & ~n20142;
  assign n20144 = controllable_BtoR_REQ0 & ~n16231;
  assign n20145 = ~n17669 & ~n20144;
  assign n20146 = ~i_RtoB_ACK0 & ~n20145;
  assign n20147 = ~n15619 & ~n20146;
  assign n20148 = controllable_DEQ & ~n20147;
  assign n20149 = ~controllable_DEQ & ~n20123;
  assign n20150 = ~n20148 & ~n20149;
  assign n20151 = ~i_FULL & ~n20150;
  assign n20152 = ~n20143 & ~n20151;
  assign n20153 = ~i_nEMPTY & ~n20152;
  assign n20154 = ~n20131 & ~n20153;
  assign n20155 = controllable_BtoS_ACK0 & ~n20154;
  assign n20156 = controllable_BtoR_REQ0 & ~n16263;
  assign n20157 = ~n19933 & ~n20156;
  assign n20158 = ~i_RtoB_ACK0 & ~n20157;
  assign n20159 = ~n17483 & ~n20158;
  assign n20160 = controllable_DEQ & ~n20159;
  assign n20161 = controllable_BtoR_REQ0 & ~n16282;
  assign n20162 = ~n19941 & ~n20161;
  assign n20163 = ~i_RtoB_ACK0 & ~n20162;
  assign n20164 = ~n17491 & ~n20163;
  assign n20165 = ~controllable_DEQ & ~n20164;
  assign n20166 = ~n20160 & ~n20165;
  assign n20167 = i_FULL & ~n20166;
  assign n20168 = controllable_BtoR_REQ0 & ~n16301;
  assign n20169 = ~n17701 & ~n20168;
  assign n20170 = ~i_RtoB_ACK0 & ~n20169;
  assign n20171 = ~n17483 & ~n20170;
  assign n20172 = controllable_DEQ & ~n20171;
  assign n20173 = controllable_BtoR_REQ0 & ~n16317;
  assign n20174 = ~n19955 & ~n20173;
  assign n20175 = ~i_RtoB_ACK0 & ~n20174;
  assign n20176 = ~n17491 & ~n20175;
  assign n20177 = ~controllable_DEQ & ~n20176;
  assign n20178 = ~n20172 & ~n20177;
  assign n20179 = ~i_FULL & ~n20178;
  assign n20180 = ~n20167 & ~n20179;
  assign n20181 = i_nEMPTY & ~n20180;
  assign n20182 = controllable_BtoR_REQ0 & ~n16338;
  assign n20183 = ~n17737 & ~n20182;
  assign n20184 = ~i_RtoB_ACK0 & ~n20183;
  assign n20185 = ~n16656 & ~n20184;
  assign n20186 = controllable_DEQ & ~n20185;
  assign n20187 = controllable_BtoR_REQ0 & ~n16354;
  assign n20188 = ~n19971 & ~n20187;
  assign n20189 = ~i_RtoB_ACK0 & ~n20188;
  assign n20190 = ~n17509 & ~n20189;
  assign n20191 = ~controllable_DEQ & ~n20190;
  assign n20192 = ~n20186 & ~n20191;
  assign n20193 = i_FULL & ~n20192;
  assign n20194 = controllable_BtoR_REQ0 & ~n16373;
  assign n20195 = ~n17770 & ~n20194;
  assign n20196 = ~i_RtoB_ACK0 & ~n20195;
  assign n20197 = ~n16677 & ~n20196;
  assign n20198 = controllable_DEQ & ~n20197;
  assign n20199 = ~controllable_DEQ & ~n20159;
  assign n20200 = ~n20198 & ~n20199;
  assign n20201 = ~i_FULL & ~n20200;
  assign n20202 = ~n20193 & ~n20201;
  assign n20203 = ~i_nEMPTY & ~n20202;
  assign n20204 = ~n20181 & ~n20203;
  assign n20205 = ~controllable_BtoS_ACK0 & ~n20204;
  assign n20206 = ~n20155 & ~n20205;
  assign n20207 = ~n4465 & ~n20206;
  assign n20208 = ~n20119 & ~n20207;
  assign n20209 = i_StoB_REQ10 & ~n20208;
  assign n20210 = ~n19999 & ~n20209;
  assign n20211 = ~controllable_BtoS_ACK10 & ~n20210;
  assign n20212 = ~n20001 & ~n20211;
  assign n20213 = ~n4464 & ~n20212;
  assign n20214 = ~n19611 & ~n20213;
  assign n20215 = n4462 & ~n20214;
  assign n20216 = ~n14741 & ~n17538;
  assign n20217 = i_RtoB_ACK0 & ~n20216;
  assign n20218 = ~n12175 & ~n14073;
  assign n20219 = ~controllable_BtoR_REQ1 & ~n20218;
  assign n20220 = ~controllable_BtoR_REQ1 & ~n20219;
  assign n20221 = ~controllable_BtoR_REQ0 & ~n20220;
  assign n20222 = ~n17545 & ~n20221;
  assign n20223 = ~i_RtoB_ACK0 & ~n20222;
  assign n20224 = ~n20217 & ~n20223;
  assign n20225 = controllable_DEQ & ~n20224;
  assign n20226 = ~n14757 & ~n17555;
  assign n20227 = i_RtoB_ACK0 & ~n20226;
  assign n20228 = ~n5243 & ~n14082;
  assign n20229 = ~controllable_BtoR_REQ1 & ~n20228;
  assign n20230 = ~controllable_BtoR_REQ1 & ~n20229;
  assign n20231 = ~controllable_BtoR_REQ0 & ~n20230;
  assign n20232 = ~n17562 & ~n20231;
  assign n20233 = ~i_RtoB_ACK0 & ~n20232;
  assign n20234 = ~n20227 & ~n20233;
  assign n20235 = ~controllable_DEQ & ~n20234;
  assign n20236 = ~n20225 & ~n20235;
  assign n20237 = i_nEMPTY & ~n20236;
  assign n20238 = ~controllable_BtoR_REQ1 & ~n12207;
  assign n20239 = ~controllable_BtoR_REQ0 & ~n20238;
  assign n20240 = ~n17571 & ~n20239;
  assign n20241 = ~i_RtoB_ACK0 & ~n20240;
  assign n20242 = ~i_RtoB_ACK0 & ~n20241;
  assign n20243 = controllable_DEQ & ~n20242;
  assign n20244 = ~n8755 & ~n14073;
  assign n20245 = ~controllable_BtoR_REQ1 & ~n20244;
  assign n20246 = ~controllable_BtoR_REQ1 & ~n20245;
  assign n20247 = ~controllable_BtoR_REQ0 & ~n20246;
  assign n20248 = ~n17581 & ~n20247;
  assign n20249 = ~i_RtoB_ACK0 & ~n20248;
  assign n20250 = ~n20217 & ~n20249;
  assign n20251 = ~controllable_DEQ & ~n20250;
  assign n20252 = ~n20243 & ~n20251;
  assign n20253 = i_FULL & ~n20252;
  assign n20254 = ~controllable_BtoR_REQ0 & ~n18433;
  assign n20255 = ~n17590 & ~n20254;
  assign n20256 = ~i_RtoB_ACK0 & ~n20255;
  assign n20257 = ~i_RtoB_ACK0 & ~n20256;
  assign n20258 = controllable_DEQ & ~n20257;
  assign n20259 = ~n5240 & ~n14073;
  assign n20260 = ~controllable_BtoR_REQ1 & ~n20259;
  assign n20261 = ~controllable_BtoR_REQ1 & ~n20260;
  assign n20262 = ~controllable_BtoR_REQ0 & ~n20261;
  assign n20263 = ~n17545 & ~n20262;
  assign n20264 = ~i_RtoB_ACK0 & ~n20263;
  assign n20265 = ~n20217 & ~n20264;
  assign n20266 = ~controllable_DEQ & ~n20265;
  assign n20267 = ~n20258 & ~n20266;
  assign n20268 = ~i_FULL & ~n20267;
  assign n20269 = ~n20253 & ~n20268;
  assign n20270 = ~i_nEMPTY & ~n20269;
  assign n20271 = ~n20237 & ~n20270;
  assign n20272 = controllable_BtoS_ACK0 & ~n20271;
  assign n20273 = ~n12266 & ~n14116;
  assign n20274 = ~controllable_BtoR_REQ1 & ~n20273;
  assign n20275 = ~controllable_BtoR_REQ1 & ~n20274;
  assign n20276 = ~controllable_BtoR_REQ0 & ~n20275;
  assign n20277 = ~n14824 & ~n20276;
  assign n20278 = ~i_RtoB_ACK0 & ~n20277;
  assign n20279 = ~n16751 & ~n20278;
  assign n20280 = controllable_DEQ & ~n20279;
  assign n20281 = ~n8876 & ~n14125;
  assign n20282 = ~controllable_BtoR_REQ1 & ~n20281;
  assign n20283 = ~controllable_BtoR_REQ1 & ~n20282;
  assign n20284 = ~controllable_BtoR_REQ0 & ~n20283;
  assign n20285 = ~n14841 & ~n20284;
  assign n20286 = ~i_RtoB_ACK0 & ~n20285;
  assign n20287 = ~n16755 & ~n20286;
  assign n20288 = ~controllable_DEQ & ~n20287;
  assign n20289 = ~n20280 & ~n20288;
  assign n20290 = i_nEMPTY & ~n20289;
  assign n20291 = ~controllable_BtoR_REQ1 & ~n12293;
  assign n20292 = ~controllable_BtoR_REQ0 & ~n20291;
  assign n20293 = ~n14850 & ~n20292;
  assign n20294 = ~i_RtoB_ACK0 & ~n20293;
  assign n20295 = ~i_RtoB_ACK0 & ~n20294;
  assign n20296 = controllable_DEQ & ~n20295;
  assign n20297 = ~n8854 & ~n14116;
  assign n20298 = ~controllable_BtoR_REQ1 & ~n20297;
  assign n20299 = ~controllable_BtoR_REQ1 & ~n20298;
  assign n20300 = ~controllable_BtoR_REQ0 & ~n20299;
  assign n20301 = ~n14860 & ~n20300;
  assign n20302 = ~i_RtoB_ACK0 & ~n20301;
  assign n20303 = ~n16751 & ~n20302;
  assign n20304 = ~controllable_DEQ & ~n20303;
  assign n20305 = ~n20296 & ~n20304;
  assign n20306 = i_FULL & ~n20305;
  assign n20307 = ~controllable_BtoR_REQ0 & ~n18461;
  assign n20308 = ~n14869 & ~n20307;
  assign n20309 = ~i_RtoB_ACK0 & ~n20308;
  assign n20310 = ~i_RtoB_ACK0 & ~n20309;
  assign n20311 = controllable_DEQ & ~n20310;
  assign n20312 = ~n12317 & ~n14116;
  assign n20313 = ~controllable_BtoR_REQ1 & ~n20312;
  assign n20314 = ~controllable_BtoR_REQ1 & ~n20313;
  assign n20315 = ~controllable_BtoR_REQ0 & ~n20314;
  assign n20316 = ~n14824 & ~n20315;
  assign n20317 = ~i_RtoB_ACK0 & ~n20316;
  assign n20318 = ~n16751 & ~n20317;
  assign n20319 = ~controllable_DEQ & ~n20318;
  assign n20320 = ~n20311 & ~n20319;
  assign n20321 = ~i_FULL & ~n20320;
  assign n20322 = ~n20306 & ~n20321;
  assign n20323 = ~i_nEMPTY & ~n20322;
  assign n20324 = ~n20290 & ~n20323;
  assign n20325 = ~controllable_BtoS_ACK0 & ~n20324;
  assign n20326 = ~n20272 & ~n20325;
  assign n20327 = n4465 & ~n20326;
  assign n20328 = ~controllable_BtoR_REQ1 & ~n8851;
  assign n20329 = ~controllable_BtoR_REQ1 & ~n20328;
  assign n20330 = ~controllable_BtoR_REQ0 & ~n20329;
  assign n20331 = ~n14841 & ~n20330;
  assign n20332 = ~i_RtoB_ACK0 & ~n20331;
  assign n20333 = ~n16755 & ~n20332;
  assign n20334 = ~controllable_DEQ & ~n20333;
  assign n20335 = ~n19022 & ~n20334;
  assign n20336 = i_nEMPTY & ~n20335;
  assign n20337 = ~controllable_BtoR_REQ1 & ~n8853;
  assign n20338 = ~controllable_BtoR_REQ1 & ~n20337;
  assign n20339 = ~controllable_BtoR_REQ0 & ~n20338;
  assign n20340 = ~n14860 & ~n20339;
  assign n20341 = ~i_RtoB_ACK0 & ~n20340;
  assign n20342 = ~n16751 & ~n20341;
  assign n20343 = ~controllable_DEQ & ~n20342;
  assign n20344 = ~n19038 & ~n20343;
  assign n20345 = i_FULL & ~n20344;
  assign n20346 = ~n8861 & ~n12317;
  assign n20347 = ~controllable_BtoR_REQ1 & ~n20346;
  assign n20348 = ~controllable_BtoR_REQ1 & ~n20347;
  assign n20349 = ~controllable_BtoR_REQ0 & ~n20348;
  assign n20350 = ~n14824 & ~n20349;
  assign n20351 = ~i_RtoB_ACK0 & ~n20350;
  assign n20352 = ~n16751 & ~n20351;
  assign n20353 = ~controllable_DEQ & ~n20352;
  assign n20354 = ~n19051 & ~n20353;
  assign n20355 = ~i_FULL & ~n20354;
  assign n20356 = ~n20345 & ~n20355;
  assign n20357 = ~i_nEMPTY & ~n20356;
  assign n20358 = ~n20336 & ~n20357;
  assign n20359 = ~controllable_BtoS_ACK0 & ~n20358;
  assign n20360 = ~n14811 & ~n20359;
  assign n20361 = ~n4465 & ~n20360;
  assign n20362 = ~n20327 & ~n20361;
  assign n20363 = i_StoB_REQ10 & ~n20362;
  assign n20364 = ~n17788 & ~n20363;
  assign n20365 = controllable_BtoS_ACK10 & ~n20364;
  assign n20366 = controllable_BtoR_REQ0 & ~n17800;
  assign n20367 = ~n9571 & ~n12370;
  assign n20368 = ~controllable_BtoR_REQ1 & ~n20367;
  assign n20369 = ~controllable_BtoR_REQ1 & ~n20368;
  assign n20370 = ~controllable_BtoR_REQ0 & ~n20369;
  assign n20371 = ~n20366 & ~n20370;
  assign n20372 = ~i_RtoB_ACK0 & ~n20371;
  assign n20373 = ~n18488 & ~n20372;
  assign n20374 = controllable_DEQ & ~n20373;
  assign n20375 = controllable_BtoR_REQ0 & ~n17812;
  assign n20376 = ~n9517 & ~n12387;
  assign n20377 = ~controllable_BtoR_REQ1 & ~n20376;
  assign n20378 = ~controllable_BtoR_REQ1 & ~n20377;
  assign n20379 = ~controllable_BtoR_REQ0 & ~n20378;
  assign n20380 = ~n20375 & ~n20379;
  assign n20381 = ~i_RtoB_ACK0 & ~n20380;
  assign n20382 = ~n18492 & ~n20381;
  assign n20383 = ~controllable_DEQ & ~n20382;
  assign n20384 = ~n20374 & ~n20383;
  assign n20385 = i_FULL & ~n20384;
  assign n20386 = controllable_BtoR_REQ0 & ~n17825;
  assign n20387 = ~n17622 & ~n20386;
  assign n20388 = ~i_RtoB_ACK0 & ~n20387;
  assign n20389 = ~n18488 & ~n20388;
  assign n20390 = controllable_DEQ & ~n20389;
  assign n20391 = controllable_BtoR_REQ0 & ~n17835;
  assign n20392 = ~n9517 & ~n12370;
  assign n20393 = ~controllable_BtoR_REQ1 & ~n20392;
  assign n20394 = ~controllable_BtoR_REQ1 & ~n20393;
  assign n20395 = ~controllable_BtoR_REQ0 & ~n20394;
  assign n20396 = ~n20391 & ~n20395;
  assign n20397 = ~i_RtoB_ACK0 & ~n20396;
  assign n20398 = ~n18492 & ~n20397;
  assign n20399 = ~controllable_DEQ & ~n20398;
  assign n20400 = ~n20390 & ~n20399;
  assign n20401 = ~i_FULL & ~n20400;
  assign n20402 = ~n20385 & ~n20401;
  assign n20403 = i_nEMPTY & ~n20402;
  assign n20404 = controllable_BtoR_REQ0 & ~n17843;
  assign n20405 = ~n17647 & ~n20404;
  assign n20406 = ~i_RtoB_ACK0 & ~n20405;
  assign n20407 = ~n15604 & ~n20406;
  assign n20408 = controllable_DEQ & ~n20407;
  assign n20409 = controllable_BtoR_REQ0 & ~n17853;
  assign n20410 = ~n9571 & ~n12431;
  assign n20411 = ~controllable_BtoR_REQ1 & ~n20410;
  assign n20412 = ~controllable_BtoR_REQ1 & ~n20411;
  assign n20413 = ~controllable_BtoR_REQ0 & ~n20412;
  assign n20414 = ~n20409 & ~n20413;
  assign n20415 = ~i_RtoB_ACK0 & ~n20414;
  assign n20416 = ~n18506 & ~n20415;
  assign n20417 = ~controllable_DEQ & ~n20416;
  assign n20418 = ~n20408 & ~n20417;
  assign n20419 = i_FULL & ~n20418;
  assign n20420 = controllable_BtoR_REQ0 & ~n17859;
  assign n20421 = ~n17669 & ~n20420;
  assign n20422 = ~i_RtoB_ACK0 & ~n20421;
  assign n20423 = ~n15619 & ~n20422;
  assign n20424 = controllable_DEQ & ~n20423;
  assign n20425 = ~controllable_DEQ & ~n20373;
  assign n20426 = ~n20424 & ~n20425;
  assign n20427 = ~i_FULL & ~n20426;
  assign n20428 = ~n20419 & ~n20427;
  assign n20429 = ~i_nEMPTY & ~n20428;
  assign n20430 = ~n20403 & ~n20429;
  assign n20431 = controllable_BtoS_ACK0 & ~n20430;
  assign n20432 = controllable_BtoR_REQ0 & ~n17879;
  assign n20433 = ~n19315 & ~n20432;
  assign n20434 = ~i_RtoB_ACK0 & ~n20433;
  assign n20435 = ~n18524 & ~n20434;
  assign n20436 = controllable_DEQ & ~n20435;
  assign n20437 = controllable_BtoR_REQ0 & ~n17891;
  assign n20438 = ~n19323 & ~n20437;
  assign n20439 = ~i_RtoB_ACK0 & ~n20438;
  assign n20440 = ~n18532 & ~n20439;
  assign n20441 = ~controllable_DEQ & ~n20440;
  assign n20442 = ~n20436 & ~n20441;
  assign n20443 = i_FULL & ~n20442;
  assign n20444 = controllable_BtoR_REQ0 & ~n17904;
  assign n20445 = ~n17701 & ~n20444;
  assign n20446 = ~i_RtoB_ACK0 & ~n20445;
  assign n20447 = ~n18524 & ~n20446;
  assign n20448 = controllable_DEQ & ~n20447;
  assign n20449 = controllable_BtoR_REQ0 & ~n17914;
  assign n20450 = ~n19337 & ~n20449;
  assign n20451 = ~i_RtoB_ACK0 & ~n20450;
  assign n20452 = ~n18532 & ~n20451;
  assign n20453 = ~controllable_DEQ & ~n20452;
  assign n20454 = ~n20448 & ~n20453;
  assign n20455 = ~i_FULL & ~n20454;
  assign n20456 = ~n20443 & ~n20455;
  assign n20457 = i_nEMPTY & ~n20456;
  assign n20458 = controllable_BtoR_REQ0 & ~n17926;
  assign n20459 = ~n17737 & ~n20458;
  assign n20460 = ~i_RtoB_ACK0 & ~n20459;
  assign n20461 = ~n17925 & ~n20460;
  assign n20462 = controllable_DEQ & ~n20461;
  assign n20463 = controllable_BtoR_REQ0 & ~n17936;
  assign n20464 = ~n19353 & ~n20463;
  assign n20465 = ~i_RtoB_ACK0 & ~n20464;
  assign n20466 = ~n18550 & ~n20465;
  assign n20467 = ~controllable_DEQ & ~n20466;
  assign n20468 = ~n20462 & ~n20467;
  assign n20469 = i_FULL & ~n20468;
  assign n20470 = controllable_BtoR_REQ0 & ~n17944;
  assign n20471 = ~n17770 & ~n20470;
  assign n20472 = ~i_RtoB_ACK0 & ~n20471;
  assign n20473 = ~n17943 & ~n20472;
  assign n20474 = controllable_DEQ & ~n20473;
  assign n20475 = ~controllable_DEQ & ~n20435;
  assign n20476 = ~n20474 & ~n20475;
  assign n20477 = ~i_FULL & ~n20476;
  assign n20478 = ~n20469 & ~n20477;
  assign n20479 = ~i_nEMPTY & ~n20478;
  assign n20480 = ~n20457 & ~n20479;
  assign n20481 = ~controllable_BtoS_ACK0 & ~n20480;
  assign n20482 = ~n20431 & ~n20481;
  assign n20483 = n4465 & ~n20482;
  assign n20484 = ~n19553 & ~n20481;
  assign n20485 = ~n4465 & ~n20484;
  assign n20486 = ~n20483 & ~n20485;
  assign n20487 = i_StoB_REQ10 & ~n20486;
  assign n20488 = ~n17974 & ~n20370;
  assign n20489 = ~i_RtoB_ACK0 & ~n20488;
  assign n20490 = ~n18574 & ~n20489;
  assign n20491 = controllable_DEQ & ~n20490;
  assign n20492 = ~n17993 & ~n20379;
  assign n20493 = ~i_RtoB_ACK0 & ~n20492;
  assign n20494 = ~n18582 & ~n20493;
  assign n20495 = ~controllable_DEQ & ~n20494;
  assign n20496 = ~n20491 & ~n20495;
  assign n20497 = i_FULL & ~n20496;
  assign n20498 = ~n17622 & ~n18012;
  assign n20499 = ~i_RtoB_ACK0 & ~n20498;
  assign n20500 = ~n18574 & ~n20499;
  assign n20501 = controllable_DEQ & ~n20500;
  assign n20502 = ~n18028 & ~n20395;
  assign n20503 = ~i_RtoB_ACK0 & ~n20502;
  assign n20504 = ~n18582 & ~n20503;
  assign n20505 = ~controllable_DEQ & ~n20504;
  assign n20506 = ~n20501 & ~n20505;
  assign n20507 = ~i_FULL & ~n20506;
  assign n20508 = ~n20497 & ~n20507;
  assign n20509 = i_nEMPTY & ~n20508;
  assign n20510 = ~n17647 & ~n18049;
  assign n20511 = ~i_RtoB_ACK0 & ~n20510;
  assign n20512 = ~n18045 & ~n20511;
  assign n20513 = controllable_DEQ & ~n20512;
  assign n20514 = ~n18065 & ~n20413;
  assign n20515 = ~i_RtoB_ACK0 & ~n20514;
  assign n20516 = ~n18600 & ~n20515;
  assign n20517 = ~controllable_DEQ & ~n20516;
  assign n20518 = ~n20513 & ~n20517;
  assign n20519 = i_FULL & ~n20518;
  assign n20520 = ~n17669 & ~n18084;
  assign n20521 = ~i_RtoB_ACK0 & ~n20520;
  assign n20522 = ~n18080 & ~n20521;
  assign n20523 = controllable_DEQ & ~n20522;
  assign n20524 = ~n9571 & ~n12629;
  assign n20525 = ~controllable_BtoR_REQ1 & ~n20524;
  assign n20526 = ~controllable_BtoR_REQ1 & ~n20525;
  assign n20527 = ~controllable_BtoR_REQ0 & ~n20526;
  assign n20528 = ~n17974 & ~n20527;
  assign n20529 = ~i_RtoB_ACK0 & ~n20528;
  assign n20530 = ~n18574 & ~n20529;
  assign n20531 = ~controllable_DEQ & ~n20530;
  assign n20532 = ~n20523 & ~n20531;
  assign n20533 = ~i_FULL & ~n20532;
  assign n20534 = ~n20519 & ~n20533;
  assign n20535 = ~i_nEMPTY & ~n20534;
  assign n20536 = ~n20509 & ~n20535;
  assign n20537 = controllable_BtoS_ACK0 & ~n20536;
  assign n20538 = ~n18116 & ~n19315;
  assign n20539 = ~i_RtoB_ACK0 & ~n20538;
  assign n20540 = ~n18619 & ~n20539;
  assign n20541 = controllable_DEQ & ~n20540;
  assign n20542 = ~n18135 & ~n19323;
  assign n20543 = ~i_RtoB_ACK0 & ~n20542;
  assign n20544 = ~n18627 & ~n20543;
  assign n20545 = ~controllable_DEQ & ~n20544;
  assign n20546 = ~n20541 & ~n20545;
  assign n20547 = i_FULL & ~n20546;
  assign n20548 = ~n17701 & ~n18154;
  assign n20549 = ~i_RtoB_ACK0 & ~n20548;
  assign n20550 = ~n18619 & ~n20549;
  assign n20551 = controllable_DEQ & ~n20550;
  assign n20552 = ~n18170 & ~n19337;
  assign n20553 = ~i_RtoB_ACK0 & ~n20552;
  assign n20554 = ~n18627 & ~n20553;
  assign n20555 = ~controllable_DEQ & ~n20554;
  assign n20556 = ~n20551 & ~n20555;
  assign n20557 = ~i_FULL & ~n20556;
  assign n20558 = ~n20547 & ~n20557;
  assign n20559 = i_nEMPTY & ~n20558;
  assign n20560 = ~n17737 & ~n18191;
  assign n20561 = ~i_RtoB_ACK0 & ~n20560;
  assign n20562 = ~n18187 & ~n20561;
  assign n20563 = controllable_DEQ & ~n20562;
  assign n20564 = ~n18207 & ~n19353;
  assign n20565 = ~i_RtoB_ACK0 & ~n20564;
  assign n20566 = ~n18645 & ~n20565;
  assign n20567 = ~controllable_DEQ & ~n20566;
  assign n20568 = ~n20563 & ~n20567;
  assign n20569 = i_FULL & ~n20568;
  assign n20570 = ~n17770 & ~n18226;
  assign n20571 = ~i_RtoB_ACK0 & ~n20570;
  assign n20572 = ~n18222 & ~n20571;
  assign n20573 = controllable_DEQ & ~n20572;
  assign n20574 = ~n18116 & ~n19367;
  assign n20575 = ~i_RtoB_ACK0 & ~n20574;
  assign n20576 = ~n18619 & ~n20575;
  assign n20577 = ~controllable_DEQ & ~n20576;
  assign n20578 = ~n20573 & ~n20577;
  assign n20579 = ~i_FULL & ~n20578;
  assign n20580 = ~n20569 & ~n20579;
  assign n20581 = ~i_nEMPTY & ~n20580;
  assign n20582 = ~n20559 & ~n20581;
  assign n20583 = ~controllable_BtoS_ACK0 & ~n20582;
  assign n20584 = ~n20537 & ~n20583;
  assign n20585 = n4465 & ~n20584;
  assign n20586 = ~n15190 & ~n17622;
  assign n20587 = ~i_RtoB_ACK0 & ~n20586;
  assign n20588 = ~n18661 & ~n20587;
  assign n20589 = controllable_DEQ & ~n20588;
  assign n20590 = ~n15209 & ~n17628;
  assign n20591 = ~i_RtoB_ACK0 & ~n20590;
  assign n20592 = ~n18665 & ~n20591;
  assign n20593 = ~controllable_DEQ & ~n20592;
  assign n20594 = ~n20589 & ~n20593;
  assign n20595 = i_nEMPTY & ~n20594;
  assign n20596 = ~n15221 & ~n17647;
  assign n20597 = ~i_RtoB_ACK0 & ~n20596;
  assign n20598 = ~n15217 & ~n20597;
  assign n20599 = controllable_DEQ & ~n20598;
  assign n20600 = ~n15237 & ~n17613;
  assign n20601 = ~i_RtoB_ACK0 & ~n20600;
  assign n20602 = ~n18671 & ~n20601;
  assign n20603 = ~controllable_DEQ & ~n20602;
  assign n20604 = ~n20599 & ~n20603;
  assign n20605 = i_FULL & ~n20604;
  assign n20606 = ~n15249 & ~n17669;
  assign n20607 = ~i_RtoB_ACK0 & ~n20606;
  assign n20608 = ~n15245 & ~n20607;
  assign n20609 = controllable_DEQ & ~n20608;
  assign n20610 = ~n15190 & ~n17675;
  assign n20611 = ~i_RtoB_ACK0 & ~n20610;
  assign n20612 = ~n18661 & ~n20611;
  assign n20613 = ~controllable_DEQ & ~n20612;
  assign n20614 = ~n20609 & ~n20613;
  assign n20615 = ~i_FULL & ~n20614;
  assign n20616 = ~n20605 & ~n20615;
  assign n20617 = ~i_nEMPTY & ~n20616;
  assign n20618 = ~n20595 & ~n20617;
  assign n20619 = controllable_BtoS_ACK0 & ~n20618;
  assign n20620 = ~n19377 & ~n20619;
  assign n20621 = ~n4465 & ~n20620;
  assign n20622 = ~n20585 & ~n20621;
  assign n20623 = ~i_StoB_REQ10 & ~n20622;
  assign n20624 = ~n20487 & ~n20623;
  assign n20625 = ~controllable_BtoS_ACK10 & ~n20624;
  assign n20626 = ~n20365 & ~n20625;
  assign n20627 = n4464 & ~n20626;
  assign n20628 = ~n14759 & ~n15749;
  assign n20629 = ~i_RtoB_ACK0 & ~n20628;
  assign n20630 = ~n17139 & ~n20629;
  assign n20631 = ~controllable_DEQ & ~n20630;
  assign n20632 = ~n19632 & ~n20631;
  assign n20633 = i_nEMPTY & ~n20632;
  assign n20634 = ~n14743 & ~n15768;
  assign n20635 = ~i_RtoB_ACK0 & ~n20634;
  assign n20636 = ~n17135 & ~n20635;
  assign n20637 = ~controllable_DEQ & ~n20636;
  assign n20638 = ~n19648 & ~n20637;
  assign n20639 = i_FULL & ~n20638;
  assign n20640 = ~n14801 & ~n15732;
  assign n20641 = ~i_RtoB_ACK0 & ~n20640;
  assign n20642 = ~n17135 & ~n20641;
  assign n20643 = ~controllable_DEQ & ~n20642;
  assign n20644 = ~n19661 & ~n20643;
  assign n20645 = ~i_FULL & ~n20644;
  assign n20646 = ~n20639 & ~n20645;
  assign n20647 = ~i_nEMPTY & ~n20646;
  assign n20648 = ~n20633 & ~n20647;
  assign n20649 = controllable_BtoS_ACK0 & ~n20648;
  assign n20650 = ~n15824 & ~n20330;
  assign n20651 = ~i_RtoB_ACK0 & ~n20650;
  assign n20652 = ~n17161 & ~n20651;
  assign n20653 = ~controllable_DEQ & ~n20652;
  assign n20654 = ~n19696 & ~n20653;
  assign n20655 = i_nEMPTY & ~n20654;
  assign n20656 = ~n15843 & ~n20339;
  assign n20657 = ~i_RtoB_ACK0 & ~n20656;
  assign n20658 = ~n17157 & ~n20657;
  assign n20659 = ~controllable_DEQ & ~n20658;
  assign n20660 = ~n19712 & ~n20659;
  assign n20661 = i_FULL & ~n20660;
  assign n20662 = ~n15807 & ~n20349;
  assign n20663 = ~i_RtoB_ACK0 & ~n20662;
  assign n20664 = ~n17157 & ~n20663;
  assign n20665 = ~controllable_DEQ & ~n20664;
  assign n20666 = ~n19725 & ~n20665;
  assign n20667 = ~i_FULL & ~n20666;
  assign n20668 = ~n20661 & ~n20667;
  assign n20669 = ~i_nEMPTY & ~n20668;
  assign n20670 = ~n20655 & ~n20669;
  assign n20671 = ~controllable_BtoS_ACK0 & ~n20670;
  assign n20672 = ~n20649 & ~n20671;
  assign n20673 = n4465 & ~n20672;
  assign n20674 = ~n14811 & ~n20671;
  assign n20675 = ~n4465 & ~n20674;
  assign n20676 = ~n20673 & ~n20675;
  assign n20677 = i_StoB_REQ10 & ~n20676;
  assign n20678 = ~n17788 & ~n20677;
  assign n20679 = controllable_BtoS_ACK10 & ~n20678;
  assign n20680 = controllable_BtoR_REQ0 & ~n18264;
  assign n20681 = ~n20006 & ~n20680;
  assign n20682 = ~i_RtoB_ACK0 & ~n20681;
  assign n20683 = ~n18695 & ~n20682;
  assign n20684 = controllable_DEQ & ~n20683;
  assign n20685 = controllable_BtoR_REQ0 & ~n18276;
  assign n20686 = ~n20015 & ~n20685;
  assign n20687 = ~i_RtoB_ACK0 & ~n20686;
  assign n20688 = ~n18699 & ~n20687;
  assign n20689 = ~controllable_DEQ & ~n20688;
  assign n20690 = ~n20684 & ~n20689;
  assign n20691 = i_FULL & ~n20690;
  assign n20692 = controllable_BtoR_REQ0 & ~n18289;
  assign n20693 = ~n17622 & ~n20692;
  assign n20694 = ~i_RtoB_ACK0 & ~n20693;
  assign n20695 = ~n18695 & ~n20694;
  assign n20696 = controllable_DEQ & ~n20695;
  assign n20697 = controllable_BtoR_REQ0 & ~n18299;
  assign n20698 = ~n20031 & ~n20697;
  assign n20699 = ~i_RtoB_ACK0 & ~n20698;
  assign n20700 = ~n18699 & ~n20699;
  assign n20701 = ~controllable_DEQ & ~n20700;
  assign n20702 = ~n20696 & ~n20701;
  assign n20703 = ~i_FULL & ~n20702;
  assign n20704 = ~n20691 & ~n20703;
  assign n20705 = i_nEMPTY & ~n20704;
  assign n20706 = controllable_BtoR_REQ0 & ~n18307;
  assign n20707 = ~n17647 & ~n20706;
  assign n20708 = ~i_RtoB_ACK0 & ~n20707;
  assign n20709 = ~n15604 & ~n20708;
  assign n20710 = controllable_DEQ & ~n20709;
  assign n20711 = controllable_BtoR_REQ0 & ~n18317;
  assign n20712 = ~n20049 & ~n20711;
  assign n20713 = ~i_RtoB_ACK0 & ~n20712;
  assign n20714 = ~n18713 & ~n20713;
  assign n20715 = ~controllable_DEQ & ~n20714;
  assign n20716 = ~n20710 & ~n20715;
  assign n20717 = i_FULL & ~n20716;
  assign n20718 = controllable_BtoR_REQ0 & ~n18323;
  assign n20719 = ~n17669 & ~n20718;
  assign n20720 = ~i_RtoB_ACK0 & ~n20719;
  assign n20721 = ~n15619 & ~n20720;
  assign n20722 = controllable_DEQ & ~n20721;
  assign n20723 = ~controllable_DEQ & ~n20683;
  assign n20724 = ~n20722 & ~n20723;
  assign n20725 = ~i_FULL & ~n20724;
  assign n20726 = ~n20717 & ~n20725;
  assign n20727 = ~i_nEMPTY & ~n20726;
  assign n20728 = ~n20705 & ~n20727;
  assign n20729 = controllable_BtoS_ACK0 & ~n20728;
  assign n20730 = controllable_BtoR_REQ0 & ~n18343;
  assign n20731 = ~n19933 & ~n20730;
  assign n20732 = ~i_RtoB_ACK0 & ~n20731;
  assign n20733 = ~n18726 & ~n20732;
  assign n20734 = controllable_DEQ & ~n20733;
  assign n20735 = controllable_BtoR_REQ0 & ~n18355;
  assign n20736 = ~n19941 & ~n20735;
  assign n20737 = ~i_RtoB_ACK0 & ~n20736;
  assign n20738 = ~n18730 & ~n20737;
  assign n20739 = ~controllable_DEQ & ~n20738;
  assign n20740 = ~n20734 & ~n20739;
  assign n20741 = i_FULL & ~n20740;
  assign n20742 = controllable_BtoR_REQ0 & ~n18368;
  assign n20743 = ~n17701 & ~n20742;
  assign n20744 = ~i_RtoB_ACK0 & ~n20743;
  assign n20745 = ~n18726 & ~n20744;
  assign n20746 = controllable_DEQ & ~n20745;
  assign n20747 = controllable_BtoR_REQ0 & ~n18378;
  assign n20748 = ~n19955 & ~n20747;
  assign n20749 = ~i_RtoB_ACK0 & ~n20748;
  assign n20750 = ~n18730 & ~n20749;
  assign n20751 = ~controllable_DEQ & ~n20750;
  assign n20752 = ~n20746 & ~n20751;
  assign n20753 = ~i_FULL & ~n20752;
  assign n20754 = ~n20741 & ~n20753;
  assign n20755 = i_nEMPTY & ~n20754;
  assign n20756 = controllable_BtoR_REQ0 & ~n18386;
  assign n20757 = ~n17737 & ~n20756;
  assign n20758 = ~i_RtoB_ACK0 & ~n20757;
  assign n20759 = ~n17925 & ~n20758;
  assign n20760 = controllable_DEQ & ~n20759;
  assign n20761 = controllable_BtoR_REQ0 & ~n18396;
  assign n20762 = ~n19971 & ~n20761;
  assign n20763 = ~i_RtoB_ACK0 & ~n20762;
  assign n20764 = ~n18744 & ~n20763;
  assign n20765 = ~controllable_DEQ & ~n20764;
  assign n20766 = ~n20760 & ~n20765;
  assign n20767 = i_FULL & ~n20766;
  assign n20768 = controllable_BtoR_REQ0 & ~n18402;
  assign n20769 = ~n17770 & ~n20768;
  assign n20770 = ~i_RtoB_ACK0 & ~n20769;
  assign n20771 = ~n17943 & ~n20770;
  assign n20772 = controllable_DEQ & ~n20771;
  assign n20773 = ~controllable_DEQ & ~n20733;
  assign n20774 = ~n20772 & ~n20773;
  assign n20775 = ~i_FULL & ~n20774;
  assign n20776 = ~n20767 & ~n20775;
  assign n20777 = ~i_nEMPTY & ~n20776;
  assign n20778 = ~n20755 & ~n20777;
  assign n20779 = ~controllable_BtoS_ACK0 & ~n20778;
  assign n20780 = ~n20729 & ~n20779;
  assign n20781 = n4465 & ~n20780;
  assign n20782 = ~n20155 & ~n20779;
  assign n20783 = ~n4465 & ~n20782;
  assign n20784 = ~n20781 & ~n20783;
  assign n20785 = i_StoB_REQ10 & ~n20784;
  assign n20786 = ~n15889 & ~n20006;
  assign n20787 = ~i_RtoB_ACK0 & ~n20786;
  assign n20788 = ~n18768 & ~n20787;
  assign n20789 = controllable_DEQ & ~n20788;
  assign n20790 = ~n15908 & ~n20015;
  assign n20791 = ~i_RtoB_ACK0 & ~n20790;
  assign n20792 = ~n18776 & ~n20791;
  assign n20793 = ~controllable_DEQ & ~n20792;
  assign n20794 = ~n20789 & ~n20793;
  assign n20795 = i_FULL & ~n20794;
  assign n20796 = ~n15927 & ~n17622;
  assign n20797 = ~i_RtoB_ACK0 & ~n20796;
  assign n20798 = ~n18768 & ~n20797;
  assign n20799 = controllable_DEQ & ~n20798;
  assign n20800 = ~n15943 & ~n20031;
  assign n20801 = ~i_RtoB_ACK0 & ~n20800;
  assign n20802 = ~n18776 & ~n20801;
  assign n20803 = ~controllable_DEQ & ~n20802;
  assign n20804 = ~n20799 & ~n20803;
  assign n20805 = ~i_FULL & ~n20804;
  assign n20806 = ~n20795 & ~n20805;
  assign n20807 = i_nEMPTY & ~n20806;
  assign n20808 = ~n15964 & ~n17647;
  assign n20809 = ~i_RtoB_ACK0 & ~n20808;
  assign n20810 = ~n15960 & ~n20809;
  assign n20811 = controllable_DEQ & ~n20810;
  assign n20812 = ~n15980 & ~n20049;
  assign n20813 = ~i_RtoB_ACK0 & ~n20812;
  assign n20814 = ~n18794 & ~n20813;
  assign n20815 = ~controllable_DEQ & ~n20814;
  assign n20816 = ~n20811 & ~n20815;
  assign n20817 = i_FULL & ~n20816;
  assign n20818 = ~n15999 & ~n17669;
  assign n20819 = ~i_RtoB_ACK0 & ~n20818;
  assign n20820 = ~n15995 & ~n20819;
  assign n20821 = controllable_DEQ & ~n20820;
  assign n20822 = ~n9571 & ~n10568;
  assign n20823 = ~controllable_BtoR_REQ1 & ~n20822;
  assign n20824 = ~controllable_BtoR_REQ1 & ~n20823;
  assign n20825 = ~controllable_BtoR_REQ0 & ~n20824;
  assign n20826 = ~n15889 & ~n20825;
  assign n20827 = ~i_RtoB_ACK0 & ~n20826;
  assign n20828 = ~n18768 & ~n20827;
  assign n20829 = ~controllable_DEQ & ~n20828;
  assign n20830 = ~n20821 & ~n20829;
  assign n20831 = ~i_FULL & ~n20830;
  assign n20832 = ~n20817 & ~n20831;
  assign n20833 = ~i_nEMPTY & ~n20832;
  assign n20834 = ~n20807 & ~n20833;
  assign n20835 = controllable_BtoS_ACK0 & ~n20834;
  assign n20836 = ~n16031 & ~n19933;
  assign n20837 = ~i_RtoB_ACK0 & ~n20836;
  assign n20838 = ~n18813 & ~n20837;
  assign n20839 = controllable_DEQ & ~n20838;
  assign n20840 = ~n16050 & ~n19941;
  assign n20841 = ~i_RtoB_ACK0 & ~n20840;
  assign n20842 = ~n18821 & ~n20841;
  assign n20843 = ~controllable_DEQ & ~n20842;
  assign n20844 = ~n20839 & ~n20843;
  assign n20845 = i_FULL & ~n20844;
  assign n20846 = ~n16069 & ~n17701;
  assign n20847 = ~i_RtoB_ACK0 & ~n20846;
  assign n20848 = ~n18813 & ~n20847;
  assign n20849 = controllable_DEQ & ~n20848;
  assign n20850 = ~n16085 & ~n19955;
  assign n20851 = ~i_RtoB_ACK0 & ~n20850;
  assign n20852 = ~n18821 & ~n20851;
  assign n20853 = ~controllable_DEQ & ~n20852;
  assign n20854 = ~n20849 & ~n20853;
  assign n20855 = ~i_FULL & ~n20854;
  assign n20856 = ~n20845 & ~n20855;
  assign n20857 = i_nEMPTY & ~n20856;
  assign n20858 = ~n16106 & ~n17737;
  assign n20859 = ~i_RtoB_ACK0 & ~n20858;
  assign n20860 = ~n16102 & ~n20859;
  assign n20861 = controllable_DEQ & ~n20860;
  assign n20862 = ~n16122 & ~n19971;
  assign n20863 = ~i_RtoB_ACK0 & ~n20862;
  assign n20864 = ~n18839 & ~n20863;
  assign n20865 = ~controllable_DEQ & ~n20864;
  assign n20866 = ~n20861 & ~n20865;
  assign n20867 = i_FULL & ~n20866;
  assign n20868 = ~n16141 & ~n17770;
  assign n20869 = ~i_RtoB_ACK0 & ~n20868;
  assign n20870 = ~n16137 & ~n20869;
  assign n20871 = controllable_DEQ & ~n20870;
  assign n20872 = ~n16031 & ~n19985;
  assign n20873 = ~i_RtoB_ACK0 & ~n20872;
  assign n20874 = ~n18813 & ~n20873;
  assign n20875 = ~controllable_DEQ & ~n20874;
  assign n20876 = ~n20871 & ~n20875;
  assign n20877 = ~i_FULL & ~n20876;
  assign n20878 = ~n20867 & ~n20877;
  assign n20879 = ~i_nEMPTY & ~n20878;
  assign n20880 = ~n20857 & ~n20879;
  assign n20881 = ~controllable_BtoS_ACK0 & ~n20880;
  assign n20882 = ~n20835 & ~n20881;
  assign n20883 = n4465 & ~n20882;
  assign n20884 = ~n19997 & ~n20883;
  assign n20885 = ~i_StoB_REQ10 & ~n20884;
  assign n20886 = ~n20785 & ~n20885;
  assign n20887 = ~controllable_BtoS_ACK10 & ~n20886;
  assign n20888 = ~n20679 & ~n20887;
  assign n20889 = ~n4464 & ~n20888;
  assign n20890 = ~n20627 & ~n20889;
  assign n20891 = ~n4462 & ~n20890;
  assign n20892 = ~n20215 & ~n20891;
  assign n20893 = ~n4461 & ~n20892;
  assign n20894 = ~n18865 & ~n20893;
  assign n20895 = n4459 & ~n20894;
  assign n20896 = ~n14585 & ~n20895;
  assign n20897 = n4455 & ~n20896;
  assign n20898 = ~n5029 & ~n14589;
  assign n20899 = i_RtoB_ACK0 & ~n20898;
  assign n20900 = ~n5042 & ~n14598;
  assign n20901 = ~i_RtoB_ACK0 & ~n20900;
  assign n20902 = ~n20899 & ~n20901;
  assign n20903 = controllable_DEQ & ~n20902;
  assign n20904 = ~n5052 & ~n14606;
  assign n20905 = i_RtoB_ACK0 & ~n20904;
  assign n20906 = ~n5055 & ~n14615;
  assign n20907 = ~i_RtoB_ACK0 & ~n20906;
  assign n20908 = ~n20905 & ~n20907;
  assign n20909 = ~controllable_DEQ & ~n20908;
  assign n20910 = ~n20903 & ~n20909;
  assign n20911 = i_nEMPTY & ~n20910;
  assign n20912 = ~n5072 & ~n14624;
  assign n20913 = ~i_RtoB_ACK0 & ~n20912;
  assign n20914 = ~i_RtoB_ACK0 & ~n20913;
  assign n20915 = controllable_DEQ & ~n20914;
  assign n20916 = ~n5077 & ~n14634;
  assign n20917 = ~i_RtoB_ACK0 & ~n20916;
  assign n20918 = ~n20899 & ~n20917;
  assign n20919 = ~controllable_DEQ & ~n20918;
  assign n20920 = ~n20915 & ~n20919;
  assign n20921 = i_FULL & ~n20920;
  assign n20922 = ~n5087 & ~n14643;
  assign n20923 = ~i_RtoB_ACK0 & ~n20922;
  assign n20924 = ~i_RtoB_ACK0 & ~n20923;
  assign n20925 = controllable_DEQ & ~n20924;
  assign n20926 = ~n5092 & ~n14598;
  assign n20927 = ~i_RtoB_ACK0 & ~n20926;
  assign n20928 = ~n20899 & ~n20927;
  assign n20929 = ~controllable_DEQ & ~n20928;
  assign n20930 = ~n20925 & ~n20929;
  assign n20931 = ~i_FULL & ~n20930;
  assign n20932 = ~n20921 & ~n20931;
  assign n20933 = ~i_nEMPTY & ~n20932;
  assign n20934 = ~n20911 & ~n20933;
  assign n20935 = controllable_BtoS_ACK0 & ~n20934;
  assign n20936 = ~n5126 & ~n14664;
  assign n20937 = i_RtoB_ACK0 & ~n20936;
  assign n20938 = ~n5139 & ~n14673;
  assign n20939 = ~i_RtoB_ACK0 & ~n20938;
  assign n20940 = ~n20937 & ~n20939;
  assign n20941 = controllable_DEQ & ~n20940;
  assign n20942 = ~n5149 & ~n14681;
  assign n20943 = i_RtoB_ACK0 & ~n20942;
  assign n20944 = ~n5152 & ~n14690;
  assign n20945 = ~i_RtoB_ACK0 & ~n20944;
  assign n20946 = ~n20943 & ~n20945;
  assign n20947 = ~controllable_DEQ & ~n20946;
  assign n20948 = ~n20941 & ~n20947;
  assign n20949 = i_nEMPTY & ~n20948;
  assign n20950 = ~n5169 & ~n14699;
  assign n20951 = ~i_RtoB_ACK0 & ~n20950;
  assign n20952 = ~i_RtoB_ACK0 & ~n20951;
  assign n20953 = controllable_DEQ & ~n20952;
  assign n20954 = ~n5174 & ~n14709;
  assign n20955 = ~i_RtoB_ACK0 & ~n20954;
  assign n20956 = ~n20937 & ~n20955;
  assign n20957 = ~controllable_DEQ & ~n20956;
  assign n20958 = ~n20953 & ~n20957;
  assign n20959 = i_FULL & ~n20958;
  assign n20960 = ~n5184 & ~n14718;
  assign n20961 = ~i_RtoB_ACK0 & ~n20960;
  assign n20962 = ~i_RtoB_ACK0 & ~n20961;
  assign n20963 = controllable_DEQ & ~n20962;
  assign n20964 = ~n5189 & ~n14673;
  assign n20965 = ~i_RtoB_ACK0 & ~n20964;
  assign n20966 = ~n20937 & ~n20965;
  assign n20967 = ~controllable_DEQ & ~n20966;
  assign n20968 = ~n20963 & ~n20967;
  assign n20969 = ~i_FULL & ~n20968;
  assign n20970 = ~n20959 & ~n20969;
  assign n20971 = ~i_nEMPTY & ~n20970;
  assign n20972 = ~n20949 & ~n20971;
  assign n20973 = ~controllable_BtoS_ACK0 & ~n20972;
  assign n20974 = ~n20935 & ~n20973;
  assign n20975 = n4465 & ~n20974;
  assign n20976 = ~n5234 & ~n14741;
  assign n20977 = i_RtoB_ACK0 & ~n20976;
  assign n20978 = ~n5247 & ~n14749;
  assign n20979 = ~i_RtoB_ACK0 & ~n20978;
  assign n20980 = ~n20977 & ~n20979;
  assign n20981 = controllable_DEQ & ~n20980;
  assign n20982 = ~n5257 & ~n14757;
  assign n20983 = i_RtoB_ACK0 & ~n20982;
  assign n20984 = ~n5260 & ~n14765;
  assign n20985 = ~i_RtoB_ACK0 & ~n20984;
  assign n20986 = ~n20983 & ~n20985;
  assign n20987 = ~controllable_DEQ & ~n20986;
  assign n20988 = ~n20981 & ~n20987;
  assign n20989 = i_nEMPTY & ~n20988;
  assign n20990 = ~n5277 & ~n14774;
  assign n20991 = ~i_RtoB_ACK0 & ~n20990;
  assign n20992 = ~i_RtoB_ACK0 & ~n20991;
  assign n20993 = controllable_DEQ & ~n20992;
  assign n20994 = ~n5282 & ~n14784;
  assign n20995 = ~i_RtoB_ACK0 & ~n20994;
  assign n20996 = ~n20977 & ~n20995;
  assign n20997 = ~controllable_DEQ & ~n20996;
  assign n20998 = ~n20993 & ~n20997;
  assign n20999 = i_FULL & ~n20998;
  assign n21000 = ~n5292 & ~n14793;
  assign n21001 = ~i_RtoB_ACK0 & ~n21000;
  assign n21002 = ~i_RtoB_ACK0 & ~n21001;
  assign n21003 = controllable_DEQ & ~n21002;
  assign n21004 = ~n5297 & ~n14749;
  assign n21005 = ~i_RtoB_ACK0 & ~n21004;
  assign n21006 = ~n20977 & ~n21005;
  assign n21007 = ~controllable_DEQ & ~n21006;
  assign n21008 = ~n21003 & ~n21007;
  assign n21009 = ~i_FULL & ~n21008;
  assign n21010 = ~n20999 & ~n21009;
  assign n21011 = ~i_nEMPTY & ~n21010;
  assign n21012 = ~n20989 & ~n21011;
  assign n21013 = controllable_BtoS_ACK0 & ~n21012;
  assign n21014 = ~n5340 & ~n14815;
  assign n21015 = i_RtoB_ACK0 & ~n21014;
  assign n21016 = ~n5353 & ~n14824;
  assign n21017 = ~i_RtoB_ACK0 & ~n21016;
  assign n21018 = ~n21015 & ~n21017;
  assign n21019 = controllable_DEQ & ~n21018;
  assign n21020 = ~n5363 & ~n14832;
  assign n21021 = i_RtoB_ACK0 & ~n21020;
  assign n21022 = ~n5366 & ~n14841;
  assign n21023 = ~i_RtoB_ACK0 & ~n21022;
  assign n21024 = ~n21021 & ~n21023;
  assign n21025 = ~controllable_DEQ & ~n21024;
  assign n21026 = ~n21019 & ~n21025;
  assign n21027 = i_nEMPTY & ~n21026;
  assign n21028 = ~n5383 & ~n14850;
  assign n21029 = ~i_RtoB_ACK0 & ~n21028;
  assign n21030 = ~i_RtoB_ACK0 & ~n21029;
  assign n21031 = controllable_DEQ & ~n21030;
  assign n21032 = ~n5388 & ~n14860;
  assign n21033 = ~i_RtoB_ACK0 & ~n21032;
  assign n21034 = ~n21015 & ~n21033;
  assign n21035 = ~controllable_DEQ & ~n21034;
  assign n21036 = ~n21031 & ~n21035;
  assign n21037 = i_FULL & ~n21036;
  assign n21038 = ~n5398 & ~n14869;
  assign n21039 = ~i_RtoB_ACK0 & ~n21038;
  assign n21040 = ~i_RtoB_ACK0 & ~n21039;
  assign n21041 = controllable_DEQ & ~n21040;
  assign n21042 = ~n5403 & ~n14824;
  assign n21043 = ~i_RtoB_ACK0 & ~n21042;
  assign n21044 = ~n21015 & ~n21043;
  assign n21045 = ~controllable_DEQ & ~n21044;
  assign n21046 = ~n21041 & ~n21045;
  assign n21047 = ~i_FULL & ~n21046;
  assign n21048 = ~n21037 & ~n21047;
  assign n21049 = ~i_nEMPTY & ~n21048;
  assign n21050 = ~n21027 & ~n21049;
  assign n21051 = ~controllable_BtoS_ACK0 & ~n21050;
  assign n21052 = ~n21013 & ~n21051;
  assign n21053 = ~n4465 & ~n21052;
  assign n21054 = ~n20975 & ~n21053;
  assign n21055 = i_StoB_REQ10 & ~n21054;
  assign n21056 = ~n6583 & ~n14895;
  assign n21057 = i_RtoB_ACK0 & ~n21056;
  assign n21058 = ~n6780 & ~n14904;
  assign n21059 = ~i_RtoB_ACK0 & ~n21058;
  assign n21060 = ~n21057 & ~n21059;
  assign n21061 = controllable_DEQ & ~n21060;
  assign n21062 = ~n6791 & ~n14914;
  assign n21063 = i_RtoB_ACK0 & ~n21062;
  assign n21064 = ~n6800 & ~n14923;
  assign n21065 = ~i_RtoB_ACK0 & ~n21064;
  assign n21066 = ~n21063 & ~n21065;
  assign n21067 = ~controllable_DEQ & ~n21066;
  assign n21068 = ~n21061 & ~n21067;
  assign n21069 = i_FULL & ~n21068;
  assign n21070 = ~n6583 & ~n14936;
  assign n21071 = i_RtoB_ACK0 & ~n21070;
  assign n21072 = ~n6817 & ~n14942;
  assign n21073 = ~i_RtoB_ACK0 & ~n21072;
  assign n21074 = ~n21071 & ~n21073;
  assign n21075 = controllable_DEQ & ~n21074;
  assign n21076 = ~n6791 & ~n14952;
  assign n21077 = i_RtoB_ACK0 & ~n21076;
  assign n21078 = ~n6826 & ~n14958;
  assign n21079 = ~i_RtoB_ACK0 & ~n21078;
  assign n21080 = ~n21077 & ~n21079;
  assign n21081 = ~controllable_DEQ & ~n21080;
  assign n21082 = ~n21075 & ~n21081;
  assign n21083 = ~i_FULL & ~n21082;
  assign n21084 = ~n21069 & ~n21083;
  assign n21085 = i_nEMPTY & ~n21084;
  assign n21086 = ~n6846 & ~n14979;
  assign n21087 = ~i_RtoB_ACK0 & ~n21086;
  assign n21088 = ~n14975 & ~n21087;
  assign n21089 = controllable_DEQ & ~n21088;
  assign n21090 = ~n6583 & ~n14989;
  assign n21091 = i_RtoB_ACK0 & ~n21090;
  assign n21092 = ~n6857 & ~n14995;
  assign n21093 = ~i_RtoB_ACK0 & ~n21092;
  assign n21094 = ~n21091 & ~n21093;
  assign n21095 = ~controllable_DEQ & ~n21094;
  assign n21096 = ~n21089 & ~n21095;
  assign n21097 = i_FULL & ~n21096;
  assign n21098 = ~n6867 & ~n15014;
  assign n21099 = ~i_RtoB_ACK0 & ~n21098;
  assign n21100 = ~n15010 & ~n21099;
  assign n21101 = controllable_DEQ & ~n21100;
  assign n21102 = ~n6875 & ~n14904;
  assign n21103 = ~i_RtoB_ACK0 & ~n21102;
  assign n21104 = ~n21057 & ~n21103;
  assign n21105 = ~controllable_DEQ & ~n21104;
  assign n21106 = ~n21101 & ~n21105;
  assign n21107 = ~i_FULL & ~n21106;
  assign n21108 = ~n21097 & ~n21107;
  assign n21109 = ~i_nEMPTY & ~n21108;
  assign n21110 = ~n21085 & ~n21109;
  assign n21111 = controllable_BtoS_ACK0 & ~n21110;
  assign n21112 = ~n6922 & ~n15037;
  assign n21113 = i_RtoB_ACK0 & ~n21112;
  assign n21114 = ~n6946 & ~n15046;
  assign n21115 = ~i_RtoB_ACK0 & ~n21114;
  assign n21116 = ~n21113 & ~n21115;
  assign n21117 = controllable_DEQ & ~n21116;
  assign n21118 = ~n6957 & ~n15056;
  assign n21119 = i_RtoB_ACK0 & ~n21118;
  assign n21120 = ~n6966 & ~n15065;
  assign n21121 = ~i_RtoB_ACK0 & ~n21120;
  assign n21122 = ~n21119 & ~n21121;
  assign n21123 = ~controllable_DEQ & ~n21122;
  assign n21124 = ~n21117 & ~n21123;
  assign n21125 = i_FULL & ~n21124;
  assign n21126 = ~n6922 & ~n15078;
  assign n21127 = i_RtoB_ACK0 & ~n21126;
  assign n21128 = ~n6983 & ~n15084;
  assign n21129 = ~i_RtoB_ACK0 & ~n21128;
  assign n21130 = ~n21127 & ~n21129;
  assign n21131 = controllable_DEQ & ~n21130;
  assign n21132 = ~n6957 & ~n15094;
  assign n21133 = i_RtoB_ACK0 & ~n21132;
  assign n21134 = ~n6992 & ~n15100;
  assign n21135 = ~i_RtoB_ACK0 & ~n21134;
  assign n21136 = ~n21133 & ~n21135;
  assign n21137 = ~controllable_DEQ & ~n21136;
  assign n21138 = ~n21131 & ~n21137;
  assign n21139 = ~i_FULL & ~n21138;
  assign n21140 = ~n21125 & ~n21139;
  assign n21141 = i_nEMPTY & ~n21140;
  assign n21142 = ~n7012 & ~n15121;
  assign n21143 = ~i_RtoB_ACK0 & ~n21142;
  assign n21144 = ~n15117 & ~n21143;
  assign n21145 = controllable_DEQ & ~n21144;
  assign n21146 = ~n6922 & ~n15131;
  assign n21147 = i_RtoB_ACK0 & ~n21146;
  assign n21148 = ~n7023 & ~n15137;
  assign n21149 = ~i_RtoB_ACK0 & ~n21148;
  assign n21150 = ~n21147 & ~n21149;
  assign n21151 = ~controllable_DEQ & ~n21150;
  assign n21152 = ~n21145 & ~n21151;
  assign n21153 = i_FULL & ~n21152;
  assign n21154 = ~n7033 & ~n15156;
  assign n21155 = ~i_RtoB_ACK0 & ~n21154;
  assign n21156 = ~n15152 & ~n21155;
  assign n21157 = controllable_DEQ & ~n21156;
  assign n21158 = ~n7041 & ~n15046;
  assign n21159 = ~i_RtoB_ACK0 & ~n21158;
  assign n21160 = ~n21113 & ~n21159;
  assign n21161 = ~controllable_DEQ & ~n21160;
  assign n21162 = ~n21157 & ~n21161;
  assign n21163 = ~i_FULL & ~n21162;
  assign n21164 = ~n21153 & ~n21163;
  assign n21165 = ~i_nEMPTY & ~n21164;
  assign n21166 = ~n21141 & ~n21165;
  assign n21167 = ~controllable_BtoS_ACK0 & ~n21166;
  assign n21168 = ~n21111 & ~n21167;
  assign n21169 = n4465 & ~n21168;
  assign n21170 = ~n7091 & ~n15181;
  assign n21171 = i_RtoB_ACK0 & ~n21170;
  assign n21172 = ~n7106 & ~n15190;
  assign n21173 = ~i_RtoB_ACK0 & ~n21172;
  assign n21174 = ~n21171 & ~n21173;
  assign n21175 = controllable_DEQ & ~n21174;
  assign n21176 = ~n7117 & ~n15200;
  assign n21177 = i_RtoB_ACK0 & ~n21176;
  assign n21178 = ~n7120 & ~n15209;
  assign n21179 = ~i_RtoB_ACK0 & ~n21178;
  assign n21180 = ~n21177 & ~n21179;
  assign n21181 = ~controllable_DEQ & ~n21180;
  assign n21182 = ~n21175 & ~n21181;
  assign n21183 = i_nEMPTY & ~n21182;
  assign n21184 = ~n7138 & ~n15221;
  assign n21185 = ~i_RtoB_ACK0 & ~n21184;
  assign n21186 = ~n15217 & ~n21185;
  assign n21187 = controllable_DEQ & ~n21186;
  assign n21188 = ~n7091 & ~n15231;
  assign n21189 = i_RtoB_ACK0 & ~n21188;
  assign n21190 = ~n7143 & ~n15237;
  assign n21191 = ~i_RtoB_ACK0 & ~n21190;
  assign n21192 = ~n21189 & ~n21191;
  assign n21193 = ~controllable_DEQ & ~n21192;
  assign n21194 = ~n21187 & ~n21193;
  assign n21195 = i_FULL & ~n21194;
  assign n21196 = ~n7153 & ~n15249;
  assign n21197 = ~i_RtoB_ACK0 & ~n21196;
  assign n21198 = ~n15245 & ~n21197;
  assign n21199 = controllable_DEQ & ~n21198;
  assign n21200 = ~n7161 & ~n15190;
  assign n21201 = ~i_RtoB_ACK0 & ~n21200;
  assign n21202 = ~n21171 & ~n21201;
  assign n21203 = ~controllable_DEQ & ~n21202;
  assign n21204 = ~n21199 & ~n21203;
  assign n21205 = ~i_FULL & ~n21204;
  assign n21206 = ~n21195 & ~n21205;
  assign n21207 = ~i_nEMPTY & ~n21206;
  assign n21208 = ~n21183 & ~n21207;
  assign n21209 = controllable_BtoS_ACK0 & ~n21208;
  assign n21210 = ~n7244 & ~n15272;
  assign n21211 = i_RtoB_ACK0 & ~n21210;
  assign n21212 = ~n7272 & ~n15281;
  assign n21213 = ~i_RtoB_ACK0 & ~n21212;
  assign n21214 = ~n21211 & ~n21213;
  assign n21215 = controllable_DEQ & ~n21214;
  assign n21216 = ~n7283 & ~n15291;
  assign n21217 = i_RtoB_ACK0 & ~n21216;
  assign n21218 = ~n7292 & ~n15300;
  assign n21219 = ~i_RtoB_ACK0 & ~n21218;
  assign n21220 = ~n21217 & ~n21219;
  assign n21221 = ~controllable_DEQ & ~n21220;
  assign n21222 = ~n21215 & ~n21221;
  assign n21223 = i_FULL & ~n21222;
  assign n21224 = ~n7244 & ~n15313;
  assign n21225 = i_RtoB_ACK0 & ~n21224;
  assign n21226 = ~n7309 & ~n15319;
  assign n21227 = ~i_RtoB_ACK0 & ~n21226;
  assign n21228 = ~n21225 & ~n21227;
  assign n21229 = controllable_DEQ & ~n21228;
  assign n21230 = ~n7283 & ~n15329;
  assign n21231 = i_RtoB_ACK0 & ~n21230;
  assign n21232 = ~n7318 & ~n15335;
  assign n21233 = ~i_RtoB_ACK0 & ~n21232;
  assign n21234 = ~n21231 & ~n21233;
  assign n21235 = ~controllable_DEQ & ~n21234;
  assign n21236 = ~n21229 & ~n21235;
  assign n21237 = ~i_FULL & ~n21236;
  assign n21238 = ~n21223 & ~n21237;
  assign n21239 = i_nEMPTY & ~n21238;
  assign n21240 = ~n7338 & ~n15356;
  assign n21241 = ~i_RtoB_ACK0 & ~n21240;
  assign n21242 = ~n15352 & ~n21241;
  assign n21243 = controllable_DEQ & ~n21242;
  assign n21244 = ~n7244 & ~n15366;
  assign n21245 = i_RtoB_ACK0 & ~n21244;
  assign n21246 = ~n7349 & ~n15372;
  assign n21247 = ~i_RtoB_ACK0 & ~n21246;
  assign n21248 = ~n21245 & ~n21247;
  assign n21249 = ~controllable_DEQ & ~n21248;
  assign n21250 = ~n21243 & ~n21249;
  assign n21251 = i_FULL & ~n21250;
  assign n21252 = ~n7359 & ~n15391;
  assign n21253 = ~i_RtoB_ACK0 & ~n21252;
  assign n21254 = ~n15387 & ~n21253;
  assign n21255 = controllable_DEQ & ~n21254;
  assign n21256 = ~n7367 & ~n15281;
  assign n21257 = ~i_RtoB_ACK0 & ~n21256;
  assign n21258 = ~n21211 & ~n21257;
  assign n21259 = ~controllable_DEQ & ~n21258;
  assign n21260 = ~n21255 & ~n21259;
  assign n21261 = ~i_FULL & ~n21260;
  assign n21262 = ~n21251 & ~n21261;
  assign n21263 = ~i_nEMPTY & ~n21262;
  assign n21264 = ~n21239 & ~n21263;
  assign n21265 = ~controllable_BtoS_ACK0 & ~n21264;
  assign n21266 = ~n21209 & ~n21265;
  assign n21267 = ~n4465 & ~n21266;
  assign n21268 = ~n21169 & ~n21267;
  assign n21269 = ~i_StoB_REQ10 & ~n21268;
  assign n21270 = ~n21055 & ~n21269;
  assign n21271 = controllable_BtoS_ACK10 & ~n21270;
  assign n21272 = ~n7396 & ~n15420;
  assign n21273 = i_RtoB_ACK0 & ~n21272;
  assign n21274 = ~n7405 & ~n19384;
  assign n21275 = ~i_RtoB_ACK0 & ~n21274;
  assign n21276 = ~n21273 & ~n21275;
  assign n21277 = controllable_DEQ & ~n21276;
  assign n21278 = ~n7414 & ~n15429;
  assign n21279 = i_RtoB_ACK0 & ~n21278;
  assign n21280 = ~n6800 & ~n19393;
  assign n21281 = ~i_RtoB_ACK0 & ~n21280;
  assign n21282 = ~n21279 & ~n21281;
  assign n21283 = ~controllable_DEQ & ~n21282;
  assign n21284 = ~n21277 & ~n21283;
  assign n21285 = i_FULL & ~n21284;
  assign n21286 = ~n7396 & ~n15441;
  assign n21287 = i_RtoB_ACK0 & ~n21286;
  assign n21288 = ~n7426 & ~n19404;
  assign n21289 = ~i_RtoB_ACK0 & ~n21288;
  assign n21290 = ~n21287 & ~n21289;
  assign n21291 = controllable_DEQ & ~n21290;
  assign n21292 = ~n7414 & ~n15450;
  assign n21293 = i_RtoB_ACK0 & ~n21292;
  assign n21294 = ~n6826 & ~n19409;
  assign n21295 = ~i_RtoB_ACK0 & ~n21294;
  assign n21296 = ~n21293 & ~n21295;
  assign n21297 = ~controllable_DEQ & ~n21296;
  assign n21298 = ~n21291 & ~n21297;
  assign n21299 = ~i_FULL & ~n21298;
  assign n21300 = ~n21285 & ~n21299;
  assign n21301 = i_nEMPTY & ~n21300;
  assign n21302 = ~n7442 & ~n19422;
  assign n21303 = ~i_RtoB_ACK0 & ~n21302;
  assign n21304 = ~n15466 & ~n21303;
  assign n21305 = controllable_DEQ & ~n21304;
  assign n21306 = ~n7396 & ~n15473;
  assign n21307 = i_RtoB_ACK0 & ~n21306;
  assign n21308 = ~n6857 & ~n19427;
  assign n21309 = ~i_RtoB_ACK0 & ~n21308;
  assign n21310 = ~n21307 & ~n21309;
  assign n21311 = ~controllable_DEQ & ~n21310;
  assign n21312 = ~n21305 & ~n21311;
  assign n21313 = i_FULL & ~n21312;
  assign n21314 = ~n7452 & ~n19438;
  assign n21315 = ~i_RtoB_ACK0 & ~n21314;
  assign n21316 = ~n15487 & ~n21315;
  assign n21317 = controllable_DEQ & ~n21316;
  assign n21318 = ~controllable_DEQ & ~n21276;
  assign n21319 = ~n21317 & ~n21318;
  assign n21320 = ~i_FULL & ~n21319;
  assign n21321 = ~n21313 & ~n21320;
  assign n21322 = ~i_nEMPTY & ~n21321;
  assign n21323 = ~n21301 & ~n21322;
  assign n21324 = controllable_BtoS_ACK0 & ~n21323;
  assign n21325 = ~n7476 & ~n15502;
  assign n21326 = i_RtoB_ACK0 & ~n21325;
  assign n21327 = ~n7485 & ~n19450;
  assign n21328 = ~i_RtoB_ACK0 & ~n21327;
  assign n21329 = ~n21326 & ~n21328;
  assign n21330 = controllable_DEQ & ~n21329;
  assign n21331 = ~n7494 & ~n15511;
  assign n21332 = i_RtoB_ACK0 & ~n21331;
  assign n21333 = ~n6966 & ~n19459;
  assign n21334 = ~i_RtoB_ACK0 & ~n21333;
  assign n21335 = ~n21332 & ~n21334;
  assign n21336 = ~controllable_DEQ & ~n21335;
  assign n21337 = ~n21330 & ~n21336;
  assign n21338 = i_FULL & ~n21337;
  assign n21339 = ~n7476 & ~n15523;
  assign n21340 = i_RtoB_ACK0 & ~n21339;
  assign n21341 = ~n7506 & ~n19470;
  assign n21342 = ~i_RtoB_ACK0 & ~n21341;
  assign n21343 = ~n21340 & ~n21342;
  assign n21344 = controllable_DEQ & ~n21343;
  assign n21345 = ~n7494 & ~n15532;
  assign n21346 = i_RtoB_ACK0 & ~n21345;
  assign n21347 = ~n6992 & ~n19475;
  assign n21348 = ~i_RtoB_ACK0 & ~n21347;
  assign n21349 = ~n21346 & ~n21348;
  assign n21350 = ~controllable_DEQ & ~n21349;
  assign n21351 = ~n21344 & ~n21350;
  assign n21352 = ~i_FULL & ~n21351;
  assign n21353 = ~n21338 & ~n21352;
  assign n21354 = i_nEMPTY & ~n21353;
  assign n21355 = ~n7522 & ~n19488;
  assign n21356 = ~i_RtoB_ACK0 & ~n21355;
  assign n21357 = ~n15548 & ~n21356;
  assign n21358 = controllable_DEQ & ~n21357;
  assign n21359 = ~n7476 & ~n15555;
  assign n21360 = i_RtoB_ACK0 & ~n21359;
  assign n21361 = ~n7023 & ~n19493;
  assign n21362 = ~i_RtoB_ACK0 & ~n21361;
  assign n21363 = ~n21360 & ~n21362;
  assign n21364 = ~controllable_DEQ & ~n21363;
  assign n21365 = ~n21358 & ~n21364;
  assign n21366 = i_FULL & ~n21365;
  assign n21367 = ~n7532 & ~n19504;
  assign n21368 = ~i_RtoB_ACK0 & ~n21367;
  assign n21369 = ~n15569 & ~n21368;
  assign n21370 = controllable_DEQ & ~n21369;
  assign n21371 = ~controllable_DEQ & ~n21329;
  assign n21372 = ~n21370 & ~n21371;
  assign n21373 = ~i_FULL & ~n21372;
  assign n21374 = ~n21366 & ~n21373;
  assign n21375 = ~i_nEMPTY & ~n21374;
  assign n21376 = ~n21354 & ~n21375;
  assign n21377 = ~controllable_BtoS_ACK0 & ~n21376;
  assign n21378 = ~n21324 & ~n21377;
  assign n21379 = n4465 & ~n21378;
  assign n21380 = ~n7550 & ~n15586;
  assign n21381 = i_RtoB_ACK0 & ~n21380;
  assign n21382 = ~n7558 & ~n19518;
  assign n21383 = ~i_RtoB_ACK0 & ~n21382;
  assign n21384 = ~n21381 & ~n21383;
  assign n21385 = controllable_DEQ & ~n21384;
  assign n21386 = ~n7567 & ~n15594;
  assign n21387 = i_RtoB_ACK0 & ~n21386;
  assign n21388 = ~n7120 & ~n19523;
  assign n21389 = ~i_RtoB_ACK0 & ~n21388;
  assign n21390 = ~n21387 & ~n21389;
  assign n21391 = ~controllable_DEQ & ~n21390;
  assign n21392 = ~n21385 & ~n21391;
  assign n21393 = i_nEMPTY & ~n21392;
  assign n21394 = ~n7578 & ~n19530;
  assign n21395 = ~i_RtoB_ACK0 & ~n21394;
  assign n21396 = ~n15604 & ~n21395;
  assign n21397 = controllable_DEQ & ~n21396;
  assign n21398 = ~n7550 & ~n15610;
  assign n21399 = i_RtoB_ACK0 & ~n21398;
  assign n21400 = ~n7143 & ~n19535;
  assign n21401 = ~i_RtoB_ACK0 & ~n21400;
  assign n21402 = ~n21399 & ~n21401;
  assign n21403 = ~controllable_DEQ & ~n21402;
  assign n21404 = ~n21397 & ~n21403;
  assign n21405 = i_FULL & ~n21404;
  assign n21406 = ~n7588 & ~n19542;
  assign n21407 = ~i_RtoB_ACK0 & ~n21406;
  assign n21408 = ~n15619 & ~n21407;
  assign n21409 = controllable_DEQ & ~n21408;
  assign n21410 = ~controllable_DEQ & ~n21384;
  assign n21411 = ~n21409 & ~n21410;
  assign n21412 = ~i_FULL & ~n21411;
  assign n21413 = ~n21405 & ~n21412;
  assign n21414 = ~i_nEMPTY & ~n21413;
  assign n21415 = ~n21393 & ~n21414;
  assign n21416 = controllable_BtoS_ACK0 & ~n21415;
  assign n21417 = ~n7612 & ~n15634;
  assign n21418 = i_RtoB_ACK0 & ~n21417;
  assign n21419 = ~n7621 & ~n19554;
  assign n21420 = ~i_RtoB_ACK0 & ~n21419;
  assign n21421 = ~n21418 & ~n21420;
  assign n21422 = controllable_DEQ & ~n21421;
  assign n21423 = ~n7630 & ~n15643;
  assign n21424 = i_RtoB_ACK0 & ~n21423;
  assign n21425 = ~n7292 & ~n19559;
  assign n21426 = ~i_RtoB_ACK0 & ~n21425;
  assign n21427 = ~n21424 & ~n21426;
  assign n21428 = ~controllable_DEQ & ~n21427;
  assign n21429 = ~n21422 & ~n21428;
  assign n21430 = i_FULL & ~n21429;
  assign n21431 = ~n7612 & ~n15655;
  assign n21432 = i_RtoB_ACK0 & ~n21431;
  assign n21433 = ~n7642 & ~n19566;
  assign n21434 = ~i_RtoB_ACK0 & ~n21433;
  assign n21435 = ~n21432 & ~n21434;
  assign n21436 = controllable_DEQ & ~n21435;
  assign n21437 = ~n7630 & ~n15664;
  assign n21438 = i_RtoB_ACK0 & ~n21437;
  assign n21439 = ~n7318 & ~n19571;
  assign n21440 = ~i_RtoB_ACK0 & ~n21439;
  assign n21441 = ~n21438 & ~n21440;
  assign n21442 = ~controllable_DEQ & ~n21441;
  assign n21443 = ~n21436 & ~n21442;
  assign n21444 = ~i_FULL & ~n21443;
  assign n21445 = ~n21430 & ~n21444;
  assign n21446 = i_nEMPTY & ~n21445;
  assign n21447 = ~n7658 & ~n19580;
  assign n21448 = ~i_RtoB_ACK0 & ~n21447;
  assign n21449 = ~n15680 & ~n21448;
  assign n21450 = controllable_DEQ & ~n21449;
  assign n21451 = ~n7612 & ~n15687;
  assign n21452 = i_RtoB_ACK0 & ~n21451;
  assign n21453 = ~n7349 & ~n19585;
  assign n21454 = ~i_RtoB_ACK0 & ~n21453;
  assign n21455 = ~n21452 & ~n21454;
  assign n21456 = ~controllable_DEQ & ~n21455;
  assign n21457 = ~n21450 & ~n21456;
  assign n21458 = i_FULL & ~n21457;
  assign n21459 = ~n7668 & ~n19592;
  assign n21460 = ~i_RtoB_ACK0 & ~n21459;
  assign n21461 = ~n15701 & ~n21460;
  assign n21462 = controllable_DEQ & ~n21461;
  assign n21463 = ~controllable_DEQ & ~n21421;
  assign n21464 = ~n21462 & ~n21463;
  assign n21465 = ~i_FULL & ~n21464;
  assign n21466 = ~n21458 & ~n21465;
  assign n21467 = ~i_nEMPTY & ~n21466;
  assign n21468 = ~n21446 & ~n21467;
  assign n21469 = ~controllable_BtoS_ACK0 & ~n21468;
  assign n21470 = ~n21416 & ~n21469;
  assign n21471 = ~n4465 & ~n21470;
  assign n21472 = ~n21379 & ~n21471;
  assign n21473 = i_StoB_REQ10 & ~n21472;
  assign n21474 = ~n21269 & ~n21473;
  assign n21475 = ~controllable_BtoS_ACK10 & ~n21474;
  assign n21476 = ~n21271 & ~n21475;
  assign n21477 = n4464 & ~n21476;
  assign n21478 = ~n7707 & ~n15723;
  assign n21479 = i_RtoB_ACK0 & ~n21478;
  assign n21480 = ~n7720 & ~n15732;
  assign n21481 = ~i_RtoB_ACK0 & ~n21480;
  assign n21482 = ~n21479 & ~n21481;
  assign n21483 = controllable_DEQ & ~n21482;
  assign n21484 = ~n7730 & ~n15740;
  assign n21485 = i_RtoB_ACK0 & ~n21484;
  assign n21486 = ~n7733 & ~n15749;
  assign n21487 = ~i_RtoB_ACK0 & ~n21486;
  assign n21488 = ~n21485 & ~n21487;
  assign n21489 = ~controllable_DEQ & ~n21488;
  assign n21490 = ~n21483 & ~n21489;
  assign n21491 = i_nEMPTY & ~n21490;
  assign n21492 = ~n7750 & ~n15758;
  assign n21493 = ~i_RtoB_ACK0 & ~n21492;
  assign n21494 = ~i_RtoB_ACK0 & ~n21493;
  assign n21495 = controllable_DEQ & ~n21494;
  assign n21496 = ~n7755 & ~n15768;
  assign n21497 = ~i_RtoB_ACK0 & ~n21496;
  assign n21498 = ~n21479 & ~n21497;
  assign n21499 = ~controllable_DEQ & ~n21498;
  assign n21500 = ~n21495 & ~n21499;
  assign n21501 = i_FULL & ~n21500;
  assign n21502 = ~n7765 & ~n15777;
  assign n21503 = ~i_RtoB_ACK0 & ~n21502;
  assign n21504 = ~i_RtoB_ACK0 & ~n21503;
  assign n21505 = controllable_DEQ & ~n21504;
  assign n21506 = ~n7770 & ~n15732;
  assign n21507 = ~i_RtoB_ACK0 & ~n21506;
  assign n21508 = ~n21479 & ~n21507;
  assign n21509 = ~controllable_DEQ & ~n21508;
  assign n21510 = ~n21505 & ~n21509;
  assign n21511 = ~i_FULL & ~n21510;
  assign n21512 = ~n21501 & ~n21511;
  assign n21513 = ~i_nEMPTY & ~n21512;
  assign n21514 = ~n21491 & ~n21513;
  assign n21515 = controllable_BtoS_ACK0 & ~n21514;
  assign n21516 = ~n7799 & ~n15798;
  assign n21517 = i_RtoB_ACK0 & ~n21516;
  assign n21518 = ~n7812 & ~n15807;
  assign n21519 = ~i_RtoB_ACK0 & ~n21518;
  assign n21520 = ~n21517 & ~n21519;
  assign n21521 = controllable_DEQ & ~n21520;
  assign n21522 = ~n7822 & ~n15815;
  assign n21523 = i_RtoB_ACK0 & ~n21522;
  assign n21524 = ~n7825 & ~n15824;
  assign n21525 = ~i_RtoB_ACK0 & ~n21524;
  assign n21526 = ~n21523 & ~n21525;
  assign n21527 = ~controllable_DEQ & ~n21526;
  assign n21528 = ~n21521 & ~n21527;
  assign n21529 = i_nEMPTY & ~n21528;
  assign n21530 = ~n7842 & ~n15833;
  assign n21531 = ~i_RtoB_ACK0 & ~n21530;
  assign n21532 = ~i_RtoB_ACK0 & ~n21531;
  assign n21533 = controllable_DEQ & ~n21532;
  assign n21534 = ~n7847 & ~n15843;
  assign n21535 = ~i_RtoB_ACK0 & ~n21534;
  assign n21536 = ~n21517 & ~n21535;
  assign n21537 = ~controllable_DEQ & ~n21536;
  assign n21538 = ~n21533 & ~n21537;
  assign n21539 = i_FULL & ~n21538;
  assign n21540 = ~n7857 & ~n15852;
  assign n21541 = ~i_RtoB_ACK0 & ~n21540;
  assign n21542 = ~i_RtoB_ACK0 & ~n21541;
  assign n21543 = controllable_DEQ & ~n21542;
  assign n21544 = ~n7862 & ~n15807;
  assign n21545 = ~i_RtoB_ACK0 & ~n21544;
  assign n21546 = ~n21517 & ~n21545;
  assign n21547 = ~controllable_DEQ & ~n21546;
  assign n21548 = ~n21543 & ~n21547;
  assign n21549 = ~i_FULL & ~n21548;
  assign n21550 = ~n21539 & ~n21549;
  assign n21551 = ~i_nEMPTY & ~n21550;
  assign n21552 = ~n21529 & ~n21551;
  assign n21553 = ~controllable_BtoS_ACK0 & ~n21552;
  assign n21554 = ~n21515 & ~n21553;
  assign n21555 = n4465 & ~n21554;
  assign n21556 = ~n21013 & ~n21553;
  assign n21557 = ~n4465 & ~n21556;
  assign n21558 = ~n21555 & ~n21557;
  assign n21559 = i_StoB_REQ10 & ~n21558;
  assign n21560 = ~n7919 & ~n15880;
  assign n21561 = i_RtoB_ACK0 & ~n21560;
  assign n21562 = ~n7942 & ~n15889;
  assign n21563 = ~i_RtoB_ACK0 & ~n21562;
  assign n21564 = ~n21561 & ~n21563;
  assign n21565 = controllable_DEQ & ~n21564;
  assign n21566 = ~n7953 & ~n15899;
  assign n21567 = i_RtoB_ACK0 & ~n21566;
  assign n21568 = ~n7962 & ~n15908;
  assign n21569 = ~i_RtoB_ACK0 & ~n21568;
  assign n21570 = ~n21567 & ~n21569;
  assign n21571 = ~controllable_DEQ & ~n21570;
  assign n21572 = ~n21565 & ~n21571;
  assign n21573 = i_FULL & ~n21572;
  assign n21574 = ~n7919 & ~n15921;
  assign n21575 = i_RtoB_ACK0 & ~n21574;
  assign n21576 = ~n7979 & ~n15927;
  assign n21577 = ~i_RtoB_ACK0 & ~n21576;
  assign n21578 = ~n21575 & ~n21577;
  assign n21579 = controllable_DEQ & ~n21578;
  assign n21580 = ~n7953 & ~n15937;
  assign n21581 = i_RtoB_ACK0 & ~n21580;
  assign n21582 = ~n7988 & ~n15943;
  assign n21583 = ~i_RtoB_ACK0 & ~n21582;
  assign n21584 = ~n21581 & ~n21583;
  assign n21585 = ~controllable_DEQ & ~n21584;
  assign n21586 = ~n21579 & ~n21585;
  assign n21587 = ~i_FULL & ~n21586;
  assign n21588 = ~n21573 & ~n21587;
  assign n21589 = i_nEMPTY & ~n21588;
  assign n21590 = ~n8008 & ~n15964;
  assign n21591 = ~i_RtoB_ACK0 & ~n21590;
  assign n21592 = ~n15960 & ~n21591;
  assign n21593 = controllable_DEQ & ~n21592;
  assign n21594 = ~n7919 & ~n15974;
  assign n21595 = i_RtoB_ACK0 & ~n21594;
  assign n21596 = ~n8019 & ~n15980;
  assign n21597 = ~i_RtoB_ACK0 & ~n21596;
  assign n21598 = ~n21595 & ~n21597;
  assign n21599 = ~controllable_DEQ & ~n21598;
  assign n21600 = ~n21593 & ~n21599;
  assign n21601 = i_FULL & ~n21600;
  assign n21602 = ~n8029 & ~n15999;
  assign n21603 = ~i_RtoB_ACK0 & ~n21602;
  assign n21604 = ~n15995 & ~n21603;
  assign n21605 = controllable_DEQ & ~n21604;
  assign n21606 = ~n8037 & ~n15889;
  assign n21607 = ~i_RtoB_ACK0 & ~n21606;
  assign n21608 = ~n21561 & ~n21607;
  assign n21609 = ~controllable_DEQ & ~n21608;
  assign n21610 = ~n21605 & ~n21609;
  assign n21611 = ~i_FULL & ~n21610;
  assign n21612 = ~n21601 & ~n21611;
  assign n21613 = ~i_nEMPTY & ~n21612;
  assign n21614 = ~n21589 & ~n21613;
  assign n21615 = controllable_BtoS_ACK0 & ~n21614;
  assign n21616 = ~n8086 & ~n16022;
  assign n21617 = i_RtoB_ACK0 & ~n21616;
  assign n21618 = ~n8106 & ~n16031;
  assign n21619 = ~i_RtoB_ACK0 & ~n21618;
  assign n21620 = ~n21617 & ~n21619;
  assign n21621 = controllable_DEQ & ~n21620;
  assign n21622 = ~n8117 & ~n16041;
  assign n21623 = i_RtoB_ACK0 & ~n21622;
  assign n21624 = ~n8126 & ~n16050;
  assign n21625 = ~i_RtoB_ACK0 & ~n21624;
  assign n21626 = ~n21623 & ~n21625;
  assign n21627 = ~controllable_DEQ & ~n21626;
  assign n21628 = ~n21621 & ~n21627;
  assign n21629 = i_FULL & ~n21628;
  assign n21630 = ~n8086 & ~n16063;
  assign n21631 = i_RtoB_ACK0 & ~n21630;
  assign n21632 = ~n8143 & ~n16069;
  assign n21633 = ~i_RtoB_ACK0 & ~n21632;
  assign n21634 = ~n21631 & ~n21633;
  assign n21635 = controllable_DEQ & ~n21634;
  assign n21636 = ~n8117 & ~n16079;
  assign n21637 = i_RtoB_ACK0 & ~n21636;
  assign n21638 = ~n8152 & ~n16085;
  assign n21639 = ~i_RtoB_ACK0 & ~n21638;
  assign n21640 = ~n21637 & ~n21639;
  assign n21641 = ~controllable_DEQ & ~n21640;
  assign n21642 = ~n21635 & ~n21641;
  assign n21643 = ~i_FULL & ~n21642;
  assign n21644 = ~n21629 & ~n21643;
  assign n21645 = i_nEMPTY & ~n21644;
  assign n21646 = ~n8172 & ~n16106;
  assign n21647 = ~i_RtoB_ACK0 & ~n21646;
  assign n21648 = ~n16102 & ~n21647;
  assign n21649 = controllable_DEQ & ~n21648;
  assign n21650 = ~n8086 & ~n16116;
  assign n21651 = i_RtoB_ACK0 & ~n21650;
  assign n21652 = ~n8183 & ~n16122;
  assign n21653 = ~i_RtoB_ACK0 & ~n21652;
  assign n21654 = ~n21651 & ~n21653;
  assign n21655 = ~controllable_DEQ & ~n21654;
  assign n21656 = ~n21649 & ~n21655;
  assign n21657 = i_FULL & ~n21656;
  assign n21658 = ~n8193 & ~n16141;
  assign n21659 = ~i_RtoB_ACK0 & ~n21658;
  assign n21660 = ~n16137 & ~n21659;
  assign n21661 = controllable_DEQ & ~n21660;
  assign n21662 = ~n8201 & ~n16031;
  assign n21663 = ~i_RtoB_ACK0 & ~n21662;
  assign n21664 = ~n21617 & ~n21663;
  assign n21665 = ~controllable_DEQ & ~n21664;
  assign n21666 = ~n21661 & ~n21665;
  assign n21667 = ~i_FULL & ~n21666;
  assign n21668 = ~n21657 & ~n21667;
  assign n21669 = ~i_nEMPTY & ~n21668;
  assign n21670 = ~n21645 & ~n21669;
  assign n21671 = ~controllable_BtoS_ACK0 & ~n21670;
  assign n21672 = ~n21615 & ~n21671;
  assign n21673 = n4465 & ~n21672;
  assign n21674 = ~n8229 & ~n16166;
  assign n21675 = i_RtoB_ACK0 & ~n21674;
  assign n21676 = ~n8244 & ~n16175;
  assign n21677 = ~i_RtoB_ACK0 & ~n21676;
  assign n21678 = ~n21675 & ~n21677;
  assign n21679 = controllable_DEQ & ~n21678;
  assign n21680 = ~n8254 & ~n16185;
  assign n21681 = i_RtoB_ACK0 & ~n21680;
  assign n21682 = ~n8257 & ~n16194;
  assign n21683 = ~i_RtoB_ACK0 & ~n21682;
  assign n21684 = ~n21681 & ~n21683;
  assign n21685 = ~controllable_DEQ & ~n21684;
  assign n21686 = ~n21679 & ~n21685;
  assign n21687 = i_nEMPTY & ~n21686;
  assign n21688 = ~n8274 & ~n16204;
  assign n21689 = ~i_RtoB_ACK0 & ~n21688;
  assign n21690 = ~n15217 & ~n21689;
  assign n21691 = controllable_DEQ & ~n21690;
  assign n21692 = ~n8229 & ~n16214;
  assign n21693 = i_RtoB_ACK0 & ~n21692;
  assign n21694 = ~n8279 & ~n16220;
  assign n21695 = ~i_RtoB_ACK0 & ~n21694;
  assign n21696 = ~n21693 & ~n21695;
  assign n21697 = ~controllable_DEQ & ~n21696;
  assign n21698 = ~n21691 & ~n21697;
  assign n21699 = i_FULL & ~n21698;
  assign n21700 = ~n8289 & ~n16230;
  assign n21701 = ~i_RtoB_ACK0 & ~n21700;
  assign n21702 = ~n15245 & ~n21701;
  assign n21703 = controllable_DEQ & ~n21702;
  assign n21704 = ~n8297 & ~n16175;
  assign n21705 = ~i_RtoB_ACK0 & ~n21704;
  assign n21706 = ~n21675 & ~n21705;
  assign n21707 = ~controllable_DEQ & ~n21706;
  assign n21708 = ~n21703 & ~n21707;
  assign n21709 = ~i_FULL & ~n21708;
  assign n21710 = ~n21699 & ~n21709;
  assign n21711 = ~i_nEMPTY & ~n21710;
  assign n21712 = ~n21687 & ~n21711;
  assign n21713 = controllable_BtoS_ACK0 & ~n21712;
  assign n21714 = ~n8329 & ~n16253;
  assign n21715 = i_RtoB_ACK0 & ~n21714;
  assign n21716 = ~n8347 & ~n16262;
  assign n21717 = ~i_RtoB_ACK0 & ~n21716;
  assign n21718 = ~n21715 & ~n21717;
  assign n21719 = controllable_DEQ & ~n21718;
  assign n21720 = ~n8358 & ~n16272;
  assign n21721 = i_RtoB_ACK0 & ~n21720;
  assign n21722 = ~n8365 & ~n16281;
  assign n21723 = ~i_RtoB_ACK0 & ~n21722;
  assign n21724 = ~n21721 & ~n21723;
  assign n21725 = ~controllable_DEQ & ~n21724;
  assign n21726 = ~n21719 & ~n21725;
  assign n21727 = i_FULL & ~n21726;
  assign n21728 = ~n8329 & ~n16294;
  assign n21729 = i_RtoB_ACK0 & ~n21728;
  assign n21730 = ~n8382 & ~n16300;
  assign n21731 = ~i_RtoB_ACK0 & ~n21730;
  assign n21732 = ~n21729 & ~n21731;
  assign n21733 = controllable_DEQ & ~n21732;
  assign n21734 = ~n8358 & ~n16310;
  assign n21735 = i_RtoB_ACK0 & ~n21734;
  assign n21736 = ~n8391 & ~n16316;
  assign n21737 = ~i_RtoB_ACK0 & ~n21736;
  assign n21738 = ~n21735 & ~n21737;
  assign n21739 = ~controllable_DEQ & ~n21738;
  assign n21740 = ~n21733 & ~n21739;
  assign n21741 = ~i_FULL & ~n21740;
  assign n21742 = ~n21727 & ~n21741;
  assign n21743 = i_nEMPTY & ~n21742;
  assign n21744 = ~n8411 & ~n16337;
  assign n21745 = ~i_RtoB_ACK0 & ~n21744;
  assign n21746 = ~n16333 & ~n21745;
  assign n21747 = controllable_DEQ & ~n21746;
  assign n21748 = ~n8329 & ~n16347;
  assign n21749 = i_RtoB_ACK0 & ~n21748;
  assign n21750 = ~n8419 & ~n16353;
  assign n21751 = ~i_RtoB_ACK0 & ~n21750;
  assign n21752 = ~n21749 & ~n21751;
  assign n21753 = ~controllable_DEQ & ~n21752;
  assign n21754 = ~n21747 & ~n21753;
  assign n21755 = i_FULL & ~n21754;
  assign n21756 = ~n8429 & ~n16372;
  assign n21757 = ~i_RtoB_ACK0 & ~n21756;
  assign n21758 = ~n16368 & ~n21757;
  assign n21759 = controllable_DEQ & ~n21758;
  assign n21760 = ~n8437 & ~n16262;
  assign n21761 = ~i_RtoB_ACK0 & ~n21760;
  assign n21762 = ~n21715 & ~n21761;
  assign n21763 = ~controllable_DEQ & ~n21762;
  assign n21764 = ~n21759 & ~n21763;
  assign n21765 = ~i_FULL & ~n21764;
  assign n21766 = ~n21755 & ~n21765;
  assign n21767 = ~i_nEMPTY & ~n21766;
  assign n21768 = ~n21743 & ~n21767;
  assign n21769 = ~controllable_BtoS_ACK0 & ~n21768;
  assign n21770 = ~n21713 & ~n21769;
  assign n21771 = ~n4465 & ~n21770;
  assign n21772 = ~n21673 & ~n21771;
  assign n21773 = ~i_StoB_REQ10 & ~n21772;
  assign n21774 = ~n21559 & ~n21773;
  assign n21775 = controllable_BtoS_ACK10 & ~n21774;
  assign n21776 = ~n8466 & ~n16401;
  assign n21777 = i_RtoB_ACK0 & ~n21776;
  assign n21778 = ~n8475 & ~n20002;
  assign n21779 = ~i_RtoB_ACK0 & ~n21778;
  assign n21780 = ~n21777 & ~n21779;
  assign n21781 = controllable_DEQ & ~n21780;
  assign n21782 = ~n8484 & ~n16410;
  assign n21783 = i_RtoB_ACK0 & ~n21782;
  assign n21784 = ~n7962 & ~n20011;
  assign n21785 = ~i_RtoB_ACK0 & ~n21784;
  assign n21786 = ~n21783 & ~n21785;
  assign n21787 = ~controllable_DEQ & ~n21786;
  assign n21788 = ~n21781 & ~n21787;
  assign n21789 = i_FULL & ~n21788;
  assign n21790 = ~n8466 & ~n16422;
  assign n21791 = i_RtoB_ACK0 & ~n21790;
  assign n21792 = ~n8496 & ~n20022;
  assign n21793 = ~i_RtoB_ACK0 & ~n21792;
  assign n21794 = ~n21791 & ~n21793;
  assign n21795 = controllable_DEQ & ~n21794;
  assign n21796 = ~n8484 & ~n16431;
  assign n21797 = i_RtoB_ACK0 & ~n21796;
  assign n21798 = ~n7988 & ~n20027;
  assign n21799 = ~i_RtoB_ACK0 & ~n21798;
  assign n21800 = ~n21797 & ~n21799;
  assign n21801 = ~controllable_DEQ & ~n21800;
  assign n21802 = ~n21795 & ~n21801;
  assign n21803 = ~i_FULL & ~n21802;
  assign n21804 = ~n21789 & ~n21803;
  assign n21805 = i_nEMPTY & ~n21804;
  assign n21806 = ~n8512 & ~n20040;
  assign n21807 = ~i_RtoB_ACK0 & ~n21806;
  assign n21808 = ~n16447 & ~n21807;
  assign n21809 = controllable_DEQ & ~n21808;
  assign n21810 = ~n8466 & ~n16454;
  assign n21811 = i_RtoB_ACK0 & ~n21810;
  assign n21812 = ~n8019 & ~n20045;
  assign n21813 = ~i_RtoB_ACK0 & ~n21812;
  assign n21814 = ~n21811 & ~n21813;
  assign n21815 = ~controllable_DEQ & ~n21814;
  assign n21816 = ~n21809 & ~n21815;
  assign n21817 = i_FULL & ~n21816;
  assign n21818 = ~n8522 & ~n20056;
  assign n21819 = ~i_RtoB_ACK0 & ~n21818;
  assign n21820 = ~n16468 & ~n21819;
  assign n21821 = controllable_DEQ & ~n21820;
  assign n21822 = ~controllable_DEQ & ~n21780;
  assign n21823 = ~n21821 & ~n21822;
  assign n21824 = ~i_FULL & ~n21823;
  assign n21825 = ~n21817 & ~n21824;
  assign n21826 = ~i_nEMPTY & ~n21825;
  assign n21827 = ~n21805 & ~n21826;
  assign n21828 = controllable_BtoS_ACK0 & ~n21827;
  assign n21829 = ~n8545 & ~n16483;
  assign n21830 = i_RtoB_ACK0 & ~n21829;
  assign n21831 = ~n8554 & ~n20068;
  assign n21832 = ~i_RtoB_ACK0 & ~n21831;
  assign n21833 = ~n21830 & ~n21832;
  assign n21834 = controllable_DEQ & ~n21833;
  assign n21835 = ~n8563 & ~n16492;
  assign n21836 = i_RtoB_ACK0 & ~n21835;
  assign n21837 = ~n8126 & ~n20073;
  assign n21838 = ~i_RtoB_ACK0 & ~n21837;
  assign n21839 = ~n21836 & ~n21838;
  assign n21840 = ~controllable_DEQ & ~n21839;
  assign n21841 = ~n21834 & ~n21840;
  assign n21842 = i_FULL & ~n21841;
  assign n21843 = ~n8545 & ~n16504;
  assign n21844 = i_RtoB_ACK0 & ~n21843;
  assign n21845 = ~n8575 & ~n20080;
  assign n21846 = ~i_RtoB_ACK0 & ~n21845;
  assign n21847 = ~n21844 & ~n21846;
  assign n21848 = controllable_DEQ & ~n21847;
  assign n21849 = ~n8563 & ~n16513;
  assign n21850 = i_RtoB_ACK0 & ~n21849;
  assign n21851 = ~n8152 & ~n20085;
  assign n21852 = ~i_RtoB_ACK0 & ~n21851;
  assign n21853 = ~n21850 & ~n21852;
  assign n21854 = ~controllable_DEQ & ~n21853;
  assign n21855 = ~n21848 & ~n21854;
  assign n21856 = ~i_FULL & ~n21855;
  assign n21857 = ~n21842 & ~n21856;
  assign n21858 = i_nEMPTY & ~n21857;
  assign n21859 = ~n8591 & ~n20094;
  assign n21860 = ~i_RtoB_ACK0 & ~n21859;
  assign n21861 = ~n16529 & ~n21860;
  assign n21862 = controllable_DEQ & ~n21861;
  assign n21863 = ~n8545 & ~n16536;
  assign n21864 = i_RtoB_ACK0 & ~n21863;
  assign n21865 = ~n8183 & ~n20099;
  assign n21866 = ~i_RtoB_ACK0 & ~n21865;
  assign n21867 = ~n21864 & ~n21866;
  assign n21868 = ~controllable_DEQ & ~n21867;
  assign n21869 = ~n21862 & ~n21868;
  assign n21870 = i_FULL & ~n21869;
  assign n21871 = ~n8601 & ~n20106;
  assign n21872 = ~i_RtoB_ACK0 & ~n21871;
  assign n21873 = ~n16550 & ~n21872;
  assign n21874 = controllable_DEQ & ~n21873;
  assign n21875 = ~controllable_DEQ & ~n21833;
  assign n21876 = ~n21874 & ~n21875;
  assign n21877 = ~i_FULL & ~n21876;
  assign n21878 = ~n21870 & ~n21877;
  assign n21879 = ~i_nEMPTY & ~n21878;
  assign n21880 = ~n21858 & ~n21879;
  assign n21881 = ~controllable_BtoS_ACK0 & ~n21880;
  assign n21882 = ~n21828 & ~n21881;
  assign n21883 = n4465 & ~n21882;
  assign n21884 = ~n8619 & ~n16567;
  assign n21885 = i_RtoB_ACK0 & ~n21884;
  assign n21886 = ~n8627 & ~n20120;
  assign n21887 = ~i_RtoB_ACK0 & ~n21886;
  assign n21888 = ~n21885 & ~n21887;
  assign n21889 = controllable_DEQ & ~n21888;
  assign n21890 = ~n8635 & ~n16575;
  assign n21891 = i_RtoB_ACK0 & ~n21890;
  assign n21892 = ~n8257 & ~n20125;
  assign n21893 = ~i_RtoB_ACK0 & ~n21892;
  assign n21894 = ~n21891 & ~n21893;
  assign n21895 = ~controllable_DEQ & ~n21894;
  assign n21896 = ~n21889 & ~n21895;
  assign n21897 = i_nEMPTY & ~n21896;
  assign n21898 = ~n8645 & ~n20132;
  assign n21899 = ~i_RtoB_ACK0 & ~n21898;
  assign n21900 = ~n15604 & ~n21899;
  assign n21901 = controllable_DEQ & ~n21900;
  assign n21902 = ~n8619 & ~n16588;
  assign n21903 = i_RtoB_ACK0 & ~n21902;
  assign n21904 = ~n8279 & ~n20137;
  assign n21905 = ~i_RtoB_ACK0 & ~n21904;
  assign n21906 = ~n21903 & ~n21905;
  assign n21907 = ~controllable_DEQ & ~n21906;
  assign n21908 = ~n21901 & ~n21907;
  assign n21909 = i_FULL & ~n21908;
  assign n21910 = ~n8655 & ~n20144;
  assign n21911 = ~i_RtoB_ACK0 & ~n21910;
  assign n21912 = ~n15619 & ~n21911;
  assign n21913 = controllable_DEQ & ~n21912;
  assign n21914 = ~controllable_DEQ & ~n21888;
  assign n21915 = ~n21913 & ~n21914;
  assign n21916 = ~i_FULL & ~n21915;
  assign n21917 = ~n21909 & ~n21916;
  assign n21918 = ~i_nEMPTY & ~n21917;
  assign n21919 = ~n21897 & ~n21918;
  assign n21920 = controllable_BtoS_ACK0 & ~n21919;
  assign n21921 = ~n8677 & ~n16610;
  assign n21922 = i_RtoB_ACK0 & ~n21921;
  assign n21923 = ~n8686 & ~n20156;
  assign n21924 = ~i_RtoB_ACK0 & ~n21923;
  assign n21925 = ~n21922 & ~n21924;
  assign n21926 = controllable_DEQ & ~n21925;
  assign n21927 = ~n8695 & ~n16619;
  assign n21928 = i_RtoB_ACK0 & ~n21927;
  assign n21929 = ~n8365 & ~n20161;
  assign n21930 = ~i_RtoB_ACK0 & ~n21929;
  assign n21931 = ~n21928 & ~n21930;
  assign n21932 = ~controllable_DEQ & ~n21931;
  assign n21933 = ~n21926 & ~n21932;
  assign n21934 = i_FULL & ~n21933;
  assign n21935 = ~n8677 & ~n16631;
  assign n21936 = i_RtoB_ACK0 & ~n21935;
  assign n21937 = ~n8707 & ~n20168;
  assign n21938 = ~i_RtoB_ACK0 & ~n21937;
  assign n21939 = ~n21936 & ~n21938;
  assign n21940 = controllable_DEQ & ~n21939;
  assign n21941 = ~n8695 & ~n16640;
  assign n21942 = i_RtoB_ACK0 & ~n21941;
  assign n21943 = ~n8391 & ~n20173;
  assign n21944 = ~i_RtoB_ACK0 & ~n21943;
  assign n21945 = ~n21942 & ~n21944;
  assign n21946 = ~controllable_DEQ & ~n21945;
  assign n21947 = ~n21940 & ~n21946;
  assign n21948 = ~i_FULL & ~n21947;
  assign n21949 = ~n21934 & ~n21948;
  assign n21950 = i_nEMPTY & ~n21949;
  assign n21951 = ~n8723 & ~n20182;
  assign n21952 = ~i_RtoB_ACK0 & ~n21951;
  assign n21953 = ~n16656 & ~n21952;
  assign n21954 = controllable_DEQ & ~n21953;
  assign n21955 = ~n8677 & ~n16663;
  assign n21956 = i_RtoB_ACK0 & ~n21955;
  assign n21957 = ~n8419 & ~n20187;
  assign n21958 = ~i_RtoB_ACK0 & ~n21957;
  assign n21959 = ~n21956 & ~n21958;
  assign n21960 = ~controllable_DEQ & ~n21959;
  assign n21961 = ~n21954 & ~n21960;
  assign n21962 = i_FULL & ~n21961;
  assign n21963 = ~n8733 & ~n20194;
  assign n21964 = ~i_RtoB_ACK0 & ~n21963;
  assign n21965 = ~n16677 & ~n21964;
  assign n21966 = controllable_DEQ & ~n21965;
  assign n21967 = ~controllable_DEQ & ~n21925;
  assign n21968 = ~n21966 & ~n21967;
  assign n21969 = ~i_FULL & ~n21968;
  assign n21970 = ~n21962 & ~n21969;
  assign n21971 = ~i_nEMPTY & ~n21970;
  assign n21972 = ~n21950 & ~n21971;
  assign n21973 = ~controllable_BtoS_ACK0 & ~n21972;
  assign n21974 = ~n21920 & ~n21973;
  assign n21975 = ~n4465 & ~n21974;
  assign n21976 = ~n21883 & ~n21975;
  assign n21977 = i_StoB_REQ10 & ~n21976;
  assign n21978 = ~n21773 & ~n21977;
  assign n21979 = ~controllable_BtoS_ACK10 & ~n21978;
  assign n21980 = ~n21775 & ~n21979;
  assign n21981 = ~n4464 & ~n21980;
  assign n21982 = ~n21477 & ~n21981;
  assign n21983 = n4463 & ~n21982;
  assign n21984 = ~n8759 & ~n14741;
  assign n21985 = i_RtoB_ACK0 & ~n21984;
  assign n21986 = ~n8769 & ~n14598;
  assign n21987 = ~i_RtoB_ACK0 & ~n21986;
  assign n21988 = ~n21985 & ~n21987;
  assign n21989 = controllable_DEQ & ~n21988;
  assign n21990 = ~n8778 & ~n14757;
  assign n21991 = i_RtoB_ACK0 & ~n21990;
  assign n21992 = ~n8784 & ~n14615;
  assign n21993 = ~i_RtoB_ACK0 & ~n21992;
  assign n21994 = ~n21991 & ~n21993;
  assign n21995 = ~controllable_DEQ & ~n21994;
  assign n21996 = ~n21989 & ~n21995;
  assign n21997 = i_FULL & ~n21996;
  assign n21998 = ~n8794 & ~n14598;
  assign n21999 = ~i_RtoB_ACK0 & ~n21998;
  assign n22000 = ~n21985 & ~n21999;
  assign n22001 = controllable_DEQ & ~n22000;
  assign n22002 = ~n8802 & ~n14615;
  assign n22003 = ~i_RtoB_ACK0 & ~n22002;
  assign n22004 = ~n21991 & ~n22003;
  assign n22005 = ~controllable_DEQ & ~n22004;
  assign n22006 = ~n22001 & ~n22005;
  assign n22007 = ~i_FULL & ~n22006;
  assign n22008 = ~n21997 & ~n22007;
  assign n22009 = i_nEMPTY & ~n22008;
  assign n22010 = ~n8812 & ~n14624;
  assign n22011 = ~i_RtoB_ACK0 & ~n22010;
  assign n22012 = ~i_RtoB_ACK0 & ~n22011;
  assign n22013 = controllable_DEQ & ~n22012;
  assign n22014 = ~n8821 & ~n14634;
  assign n22015 = ~i_RtoB_ACK0 & ~n22014;
  assign n22016 = ~n21985 & ~n22015;
  assign n22017 = ~controllable_DEQ & ~n22016;
  assign n22018 = ~n22013 & ~n22017;
  assign n22019 = i_FULL & ~n22018;
  assign n22020 = ~n8829 & ~n14643;
  assign n22021 = ~i_RtoB_ACK0 & ~n22020;
  assign n22022 = ~i_RtoB_ACK0 & ~n22021;
  assign n22023 = controllable_DEQ & ~n22022;
  assign n22024 = ~n8839 & ~n14598;
  assign n22025 = ~i_RtoB_ACK0 & ~n22024;
  assign n22026 = ~n21985 & ~n22025;
  assign n22027 = ~controllable_DEQ & ~n22026;
  assign n22028 = ~n22023 & ~n22027;
  assign n22029 = ~i_FULL & ~n22028;
  assign n22030 = ~n22019 & ~n22029;
  assign n22031 = ~i_nEMPTY & ~n22030;
  assign n22032 = ~n22009 & ~n22031;
  assign n22033 = controllable_BtoS_ACK0 & ~n22032;
  assign n22034 = ~n8858 & ~n16723;
  assign n22035 = i_RtoB_ACK0 & ~n22034;
  assign n22036 = ~n8870 & ~n14673;
  assign n22037 = ~i_RtoB_ACK0 & ~n22036;
  assign n22038 = ~n22035 & ~n22037;
  assign n22039 = controllable_DEQ & ~n22038;
  assign n22040 = ~n8880 & ~n16729;
  assign n22041 = i_RtoB_ACK0 & ~n22040;
  assign n22042 = ~n8887 & ~n14690;
  assign n22043 = ~i_RtoB_ACK0 & ~n22042;
  assign n22044 = ~n22041 & ~n22043;
  assign n22045 = ~controllable_DEQ & ~n22044;
  assign n22046 = ~n22039 & ~n22045;
  assign n22047 = i_FULL & ~n22046;
  assign n22048 = ~n8897 & ~n14673;
  assign n22049 = ~i_RtoB_ACK0 & ~n22048;
  assign n22050 = ~n22035 & ~n22049;
  assign n22051 = controllable_DEQ & ~n22050;
  assign n22052 = ~n8905 & ~n14690;
  assign n22053 = ~i_RtoB_ACK0 & ~n22052;
  assign n22054 = ~n22041 & ~n22053;
  assign n22055 = ~controllable_DEQ & ~n22054;
  assign n22056 = ~n22051 & ~n22055;
  assign n22057 = ~i_FULL & ~n22056;
  assign n22058 = ~n22047 & ~n22057;
  assign n22059 = i_nEMPTY & ~n22058;
  assign n22060 = ~n8919 & ~n14699;
  assign n22061 = ~i_RtoB_ACK0 & ~n22060;
  assign n22062 = ~i_RtoB_ACK0 & ~n22061;
  assign n22063 = controllable_DEQ & ~n22062;
  assign n22064 = ~n8928 & ~n14709;
  assign n22065 = ~i_RtoB_ACK0 & ~n22064;
  assign n22066 = ~n22035 & ~n22065;
  assign n22067 = ~controllable_DEQ & ~n22066;
  assign n22068 = ~n22063 & ~n22067;
  assign n22069 = i_FULL & ~n22068;
  assign n22070 = ~n8938 & ~n14718;
  assign n22071 = ~i_RtoB_ACK0 & ~n22070;
  assign n22072 = ~i_RtoB_ACK0 & ~n22071;
  assign n22073 = controllable_DEQ & ~n22072;
  assign n22074 = ~n8952 & ~n14673;
  assign n22075 = ~i_RtoB_ACK0 & ~n22074;
  assign n22076 = ~n22035 & ~n22075;
  assign n22077 = ~controllable_DEQ & ~n22076;
  assign n22078 = ~n22073 & ~n22077;
  assign n22079 = ~i_FULL & ~n22078;
  assign n22080 = ~n22069 & ~n22079;
  assign n22081 = ~i_nEMPTY & ~n22080;
  assign n22082 = ~n22059 & ~n22081;
  assign n22083 = ~controllable_BtoS_ACK0 & ~n22082;
  assign n22084 = ~n22033 & ~n22083;
  assign n22085 = n4465 & ~n22084;
  assign n22086 = ~n8968 & ~n16723;
  assign n22087 = i_RtoB_ACK0 & ~n22086;
  assign n22088 = ~n8978 & ~n14824;
  assign n22089 = ~i_RtoB_ACK0 & ~n22088;
  assign n22090 = ~n22087 & ~n22089;
  assign n22091 = controllable_DEQ & ~n22090;
  assign n22092 = ~n8987 & ~n16729;
  assign n22093 = i_RtoB_ACK0 & ~n22092;
  assign n22094 = ~n8993 & ~n14841;
  assign n22095 = ~i_RtoB_ACK0 & ~n22094;
  assign n22096 = ~n22093 & ~n22095;
  assign n22097 = ~controllable_DEQ & ~n22096;
  assign n22098 = ~n22091 & ~n22097;
  assign n22099 = i_FULL & ~n22098;
  assign n22100 = ~n9003 & ~n14824;
  assign n22101 = ~i_RtoB_ACK0 & ~n22100;
  assign n22102 = ~n22087 & ~n22101;
  assign n22103 = controllable_DEQ & ~n22102;
  assign n22104 = ~n9011 & ~n14841;
  assign n22105 = ~i_RtoB_ACK0 & ~n22104;
  assign n22106 = ~n22093 & ~n22105;
  assign n22107 = ~controllable_DEQ & ~n22106;
  assign n22108 = ~n22103 & ~n22107;
  assign n22109 = ~i_FULL & ~n22108;
  assign n22110 = ~n22099 & ~n22109;
  assign n22111 = i_nEMPTY & ~n22110;
  assign n22112 = ~n9021 & ~n14850;
  assign n22113 = ~i_RtoB_ACK0 & ~n22112;
  assign n22114 = ~i_RtoB_ACK0 & ~n22113;
  assign n22115 = controllable_DEQ & ~n22114;
  assign n22116 = ~n9030 & ~n14860;
  assign n22117 = ~i_RtoB_ACK0 & ~n22116;
  assign n22118 = ~n22087 & ~n22117;
  assign n22119 = ~controllable_DEQ & ~n22118;
  assign n22120 = ~n22115 & ~n22119;
  assign n22121 = i_FULL & ~n22120;
  assign n22122 = ~n9038 & ~n14869;
  assign n22123 = ~i_RtoB_ACK0 & ~n22122;
  assign n22124 = ~i_RtoB_ACK0 & ~n22123;
  assign n22125 = controllable_DEQ & ~n22124;
  assign n22126 = ~n9048 & ~n14824;
  assign n22127 = ~i_RtoB_ACK0 & ~n22126;
  assign n22128 = ~n22087 & ~n22127;
  assign n22129 = ~controllable_DEQ & ~n22128;
  assign n22130 = ~n22125 & ~n22129;
  assign n22131 = ~i_FULL & ~n22130;
  assign n22132 = ~n22121 & ~n22131;
  assign n22133 = ~i_nEMPTY & ~n22132;
  assign n22134 = ~n22111 & ~n22133;
  assign n22135 = ~controllable_BtoS_ACK0 & ~n22134;
  assign n22136 = ~n21013 & ~n22135;
  assign n22137 = ~n4465 & ~n22136;
  assign n22138 = ~n22085 & ~n22137;
  assign n22139 = i_StoB_REQ10 & ~n22138;
  assign n22140 = ~n9297 & ~n16780;
  assign n22141 = i_RtoB_ACK0 & ~n22140;
  assign n22142 = ~n9505 & ~n14904;
  assign n22143 = ~i_RtoB_ACK0 & ~n22142;
  assign n22144 = ~n22141 & ~n22143;
  assign n22145 = controllable_DEQ & ~n22144;
  assign n22146 = ~n9514 & ~n16788;
  assign n22147 = i_RtoB_ACK0 & ~n22146;
  assign n22148 = ~n9524 & ~n14923;
  assign n22149 = ~i_RtoB_ACK0 & ~n22148;
  assign n22150 = ~n22147 & ~n22149;
  assign n22151 = ~controllable_DEQ & ~n22150;
  assign n22152 = ~n22145 & ~n22151;
  assign n22153 = i_FULL & ~n22152;
  assign n22154 = ~n9538 & ~n14942;
  assign n22155 = ~i_RtoB_ACK0 & ~n22154;
  assign n22156 = ~n22141 & ~n22155;
  assign n22157 = controllable_DEQ & ~n22156;
  assign n22158 = ~n9551 & ~n14958;
  assign n22159 = ~i_RtoB_ACK0 & ~n22158;
  assign n22160 = ~n22147 & ~n22159;
  assign n22161 = ~controllable_DEQ & ~n22160;
  assign n22162 = ~n22157 & ~n22161;
  assign n22163 = ~i_FULL & ~n22162;
  assign n22164 = ~n22153 & ~n22163;
  assign n22165 = i_nEMPTY & ~n22164;
  assign n22166 = ~n9565 & ~n14979;
  assign n22167 = ~i_RtoB_ACK0 & ~n22166;
  assign n22168 = ~n14975 & ~n22167;
  assign n22169 = controllable_DEQ & ~n22168;
  assign n22170 = ~n9297 & ~n16806;
  assign n22171 = i_RtoB_ACK0 & ~n22170;
  assign n22172 = ~n9579 & ~n14995;
  assign n22173 = ~i_RtoB_ACK0 & ~n22172;
  assign n22174 = ~n22171 & ~n22173;
  assign n22175 = ~controllable_DEQ & ~n22174;
  assign n22176 = ~n22169 & ~n22175;
  assign n22177 = i_FULL & ~n22176;
  assign n22178 = ~n9589 & ~n15014;
  assign n22179 = ~i_RtoB_ACK0 & ~n22178;
  assign n22180 = ~n15010 & ~n22179;
  assign n22181 = controllable_DEQ & ~n22180;
  assign n22182 = ~n9603 & ~n14904;
  assign n22183 = ~i_RtoB_ACK0 & ~n22182;
  assign n22184 = ~n22141 & ~n22183;
  assign n22185 = ~controllable_DEQ & ~n22184;
  assign n22186 = ~n22181 & ~n22185;
  assign n22187 = ~i_FULL & ~n22186;
  assign n22188 = ~n22177 & ~n22187;
  assign n22189 = ~i_nEMPTY & ~n22188;
  assign n22190 = ~n22165 & ~n22189;
  assign n22191 = controllable_BtoS_ACK0 & ~n22190;
  assign n22192 = ~n9628 & ~n16825;
  assign n22193 = i_RtoB_ACK0 & ~n22192;
  assign n22194 = ~n9652 & ~n15046;
  assign n22195 = ~i_RtoB_ACK0 & ~n22194;
  assign n22196 = ~n22193 & ~n22195;
  assign n22197 = controllable_DEQ & ~n22196;
  assign n22198 = ~n9661 & ~n16833;
  assign n22199 = i_RtoB_ACK0 & ~n22198;
  assign n22200 = ~n9671 & ~n15065;
  assign n22201 = ~i_RtoB_ACK0 & ~n22200;
  assign n22202 = ~n22199 & ~n22201;
  assign n22203 = ~controllable_DEQ & ~n22202;
  assign n22204 = ~n22197 & ~n22203;
  assign n22205 = i_FULL & ~n22204;
  assign n22206 = ~n9685 & ~n15084;
  assign n22207 = ~i_RtoB_ACK0 & ~n22206;
  assign n22208 = ~n22193 & ~n22207;
  assign n22209 = controllable_DEQ & ~n22208;
  assign n22210 = ~n9698 & ~n15100;
  assign n22211 = ~i_RtoB_ACK0 & ~n22210;
  assign n22212 = ~n22199 & ~n22211;
  assign n22213 = ~controllable_DEQ & ~n22212;
  assign n22214 = ~n22209 & ~n22213;
  assign n22215 = ~i_FULL & ~n22214;
  assign n22216 = ~n22205 & ~n22215;
  assign n22217 = i_nEMPTY & ~n22216;
  assign n22218 = ~n9712 & ~n15121;
  assign n22219 = ~i_RtoB_ACK0 & ~n22218;
  assign n22220 = ~n15117 & ~n22219;
  assign n22221 = controllable_DEQ & ~n22220;
  assign n22222 = ~n9628 & ~n16851;
  assign n22223 = i_RtoB_ACK0 & ~n22222;
  assign n22224 = ~n9726 & ~n15137;
  assign n22225 = ~i_RtoB_ACK0 & ~n22224;
  assign n22226 = ~n22223 & ~n22225;
  assign n22227 = ~controllable_DEQ & ~n22226;
  assign n22228 = ~n22221 & ~n22227;
  assign n22229 = i_FULL & ~n22228;
  assign n22230 = ~n9736 & ~n15156;
  assign n22231 = ~i_RtoB_ACK0 & ~n22230;
  assign n22232 = ~n15152 & ~n22231;
  assign n22233 = controllable_DEQ & ~n22232;
  assign n22234 = ~n9753 & ~n15046;
  assign n22235 = ~i_RtoB_ACK0 & ~n22234;
  assign n22236 = ~n22193 & ~n22235;
  assign n22237 = ~controllable_DEQ & ~n22236;
  assign n22238 = ~n22233 & ~n22237;
  assign n22239 = ~i_FULL & ~n22238;
  assign n22240 = ~n22229 & ~n22239;
  assign n22241 = ~i_nEMPTY & ~n22240;
  assign n22242 = ~n22217 & ~n22241;
  assign n22243 = ~controllable_BtoS_ACK0 & ~n22242;
  assign n22244 = ~n22191 & ~n22243;
  assign n22245 = n4465 & ~n22244;
  assign n22246 = ~n9785 & ~n16872;
  assign n22247 = i_RtoB_ACK0 & ~n22246;
  assign n22248 = ~n9798 & ~n15190;
  assign n22249 = ~i_RtoB_ACK0 & ~n22248;
  assign n22250 = ~n22247 & ~n22249;
  assign n22251 = controllable_DEQ & ~n22250;
  assign n22252 = ~n9808 & ~n16880;
  assign n22253 = i_RtoB_ACK0 & ~n22252;
  assign n22254 = ~n9817 & ~n15209;
  assign n22255 = ~i_RtoB_ACK0 & ~n22254;
  assign n22256 = ~n22253 & ~n22255;
  assign n22257 = ~controllable_DEQ & ~n22256;
  assign n22258 = ~n22251 & ~n22257;
  assign n22259 = i_nEMPTY & ~n22258;
  assign n22260 = ~n9829 & ~n15221;
  assign n22261 = ~i_RtoB_ACK0 & ~n22260;
  assign n22262 = ~n15217 & ~n22261;
  assign n22263 = controllable_DEQ & ~n22262;
  assign n22264 = ~n9785 & ~n16890;
  assign n22265 = i_RtoB_ACK0 & ~n22264;
  assign n22266 = ~n9840 & ~n15237;
  assign n22267 = ~i_RtoB_ACK0 & ~n22266;
  assign n22268 = ~n22265 & ~n22267;
  assign n22269 = ~controllable_DEQ & ~n22268;
  assign n22270 = ~n22263 & ~n22269;
  assign n22271 = i_FULL & ~n22270;
  assign n22272 = ~n9850 & ~n15249;
  assign n22273 = ~i_RtoB_ACK0 & ~n22272;
  assign n22274 = ~n15245 & ~n22273;
  assign n22275 = controllable_DEQ & ~n22274;
  assign n22276 = ~n9860 & ~n15190;
  assign n22277 = ~i_RtoB_ACK0 & ~n22276;
  assign n22278 = ~n22247 & ~n22277;
  assign n22279 = ~controllable_DEQ & ~n22278;
  assign n22280 = ~n22275 & ~n22279;
  assign n22281 = ~i_FULL & ~n22280;
  assign n22282 = ~n22271 & ~n22281;
  assign n22283 = ~i_nEMPTY & ~n22282;
  assign n22284 = ~n22259 & ~n22283;
  assign n22285 = controllable_BtoS_ACK0 & ~n22284;
  assign n22286 = ~n9875 & ~n16909;
  assign n22287 = i_RtoB_ACK0 & ~n22286;
  assign n22288 = ~n9899 & ~n15281;
  assign n22289 = ~i_RtoB_ACK0 & ~n22288;
  assign n22290 = ~n22287 & ~n22289;
  assign n22291 = controllable_DEQ & ~n22290;
  assign n22292 = ~n9908 & ~n16917;
  assign n22293 = i_RtoB_ACK0 & ~n22292;
  assign n22294 = ~n9917 & ~n15300;
  assign n22295 = ~i_RtoB_ACK0 & ~n22294;
  assign n22296 = ~n22293 & ~n22295;
  assign n22297 = ~controllable_DEQ & ~n22296;
  assign n22298 = ~n22291 & ~n22297;
  assign n22299 = i_FULL & ~n22298;
  assign n22300 = ~n9929 & ~n15319;
  assign n22301 = ~i_RtoB_ACK0 & ~n22300;
  assign n22302 = ~n22287 & ~n22301;
  assign n22303 = controllable_DEQ & ~n22302;
  assign n22304 = ~n9939 & ~n15335;
  assign n22305 = ~i_RtoB_ACK0 & ~n22304;
  assign n22306 = ~n22293 & ~n22305;
  assign n22307 = ~controllable_DEQ & ~n22306;
  assign n22308 = ~n22303 & ~n22307;
  assign n22309 = ~i_FULL & ~n22308;
  assign n22310 = ~n22299 & ~n22309;
  assign n22311 = i_nEMPTY & ~n22310;
  assign n22312 = ~n9953 & ~n15356;
  assign n22313 = ~i_RtoB_ACK0 & ~n22312;
  assign n22314 = ~n15352 & ~n22313;
  assign n22315 = controllable_DEQ & ~n22314;
  assign n22316 = ~n9875 & ~n16935;
  assign n22317 = i_RtoB_ACK0 & ~n22316;
  assign n22318 = ~n9965 & ~n15372;
  assign n22319 = ~i_RtoB_ACK0 & ~n22318;
  assign n22320 = ~n22317 & ~n22319;
  assign n22321 = ~controllable_DEQ & ~n22320;
  assign n22322 = ~n22315 & ~n22321;
  assign n22323 = i_FULL & ~n22322;
  assign n22324 = ~n9975 & ~n15391;
  assign n22325 = ~i_RtoB_ACK0 & ~n22324;
  assign n22326 = ~n15387 & ~n22325;
  assign n22327 = controllable_DEQ & ~n22326;
  assign n22328 = ~n9985 & ~n15281;
  assign n22329 = ~i_RtoB_ACK0 & ~n22328;
  assign n22330 = ~n22287 & ~n22329;
  assign n22331 = ~controllable_DEQ & ~n22330;
  assign n22332 = ~n22327 & ~n22331;
  assign n22333 = ~i_FULL & ~n22332;
  assign n22334 = ~n22323 & ~n22333;
  assign n22335 = ~i_nEMPTY & ~n22334;
  assign n22336 = ~n22311 & ~n22335;
  assign n22337 = ~controllable_BtoS_ACK0 & ~n22336;
  assign n22338 = ~n22285 & ~n22337;
  assign n22339 = ~n4465 & ~n22338;
  assign n22340 = ~n22245 & ~n22339;
  assign n22341 = ~i_StoB_REQ10 & ~n22340;
  assign n22342 = ~n22139 & ~n22341;
  assign n22343 = controllable_BtoS_ACK10 & ~n22342;
  assign n22344 = ~n10005 & ~n16960;
  assign n22345 = i_RtoB_ACK0 & ~n22344;
  assign n22346 = ~n10015 & ~n19384;
  assign n22347 = ~i_RtoB_ACK0 & ~n22346;
  assign n22348 = ~n22345 & ~n22347;
  assign n22349 = controllable_DEQ & ~n22348;
  assign n22350 = ~n10023 & ~n16968;
  assign n22351 = i_RtoB_ACK0 & ~n22350;
  assign n22352 = ~n9524 & ~n19393;
  assign n22353 = ~i_RtoB_ACK0 & ~n22352;
  assign n22354 = ~n22351 & ~n22353;
  assign n22355 = ~controllable_DEQ & ~n22354;
  assign n22356 = ~n22349 & ~n22355;
  assign n22357 = i_FULL & ~n22356;
  assign n22358 = ~n10035 & ~n19404;
  assign n22359 = ~i_RtoB_ACK0 & ~n22358;
  assign n22360 = ~n22345 & ~n22359;
  assign n22361 = controllable_DEQ & ~n22360;
  assign n22362 = ~n9551 & ~n19409;
  assign n22363 = ~i_RtoB_ACK0 & ~n22362;
  assign n22364 = ~n22351 & ~n22363;
  assign n22365 = ~controllable_DEQ & ~n22364;
  assign n22366 = ~n22361 & ~n22365;
  assign n22367 = ~i_FULL & ~n22366;
  assign n22368 = ~n22357 & ~n22367;
  assign n22369 = i_nEMPTY & ~n22368;
  assign n22370 = ~n10051 & ~n19422;
  assign n22371 = ~i_RtoB_ACK0 & ~n22370;
  assign n22372 = ~n15466 & ~n22371;
  assign n22373 = controllable_DEQ & ~n22372;
  assign n22374 = ~n10005 & ~n16986;
  assign n22375 = i_RtoB_ACK0 & ~n22374;
  assign n22376 = ~n9579 & ~n19427;
  assign n22377 = ~i_RtoB_ACK0 & ~n22376;
  assign n22378 = ~n22375 & ~n22377;
  assign n22379 = ~controllable_DEQ & ~n22378;
  assign n22380 = ~n22373 & ~n22379;
  assign n22381 = i_FULL & ~n22380;
  assign n22382 = ~n10063 & ~n19438;
  assign n22383 = ~i_RtoB_ACK0 & ~n22382;
  assign n22384 = ~n15487 & ~n22383;
  assign n22385 = controllable_DEQ & ~n22384;
  assign n22386 = ~controllable_DEQ & ~n22348;
  assign n22387 = ~n22385 & ~n22386;
  assign n22388 = ~i_FULL & ~n22387;
  assign n22389 = ~n22381 & ~n22388;
  assign n22390 = ~i_nEMPTY & ~n22389;
  assign n22391 = ~n22369 & ~n22390;
  assign n22392 = controllable_BtoS_ACK0 & ~n22391;
  assign n22393 = ~n10078 & ~n17004;
  assign n22394 = i_RtoB_ACK0 & ~n22393;
  assign n22395 = ~n10088 & ~n19450;
  assign n22396 = ~i_RtoB_ACK0 & ~n22395;
  assign n22397 = ~n22394 & ~n22396;
  assign n22398 = controllable_DEQ & ~n22397;
  assign n22399 = ~n10096 & ~n17012;
  assign n22400 = i_RtoB_ACK0 & ~n22399;
  assign n22401 = ~n9671 & ~n19459;
  assign n22402 = ~i_RtoB_ACK0 & ~n22401;
  assign n22403 = ~n22400 & ~n22402;
  assign n22404 = ~controllable_DEQ & ~n22403;
  assign n22405 = ~n22398 & ~n22404;
  assign n22406 = i_FULL & ~n22405;
  assign n22407 = ~n10108 & ~n19470;
  assign n22408 = ~i_RtoB_ACK0 & ~n22407;
  assign n22409 = ~n22394 & ~n22408;
  assign n22410 = controllable_DEQ & ~n22409;
  assign n22411 = ~n9698 & ~n19475;
  assign n22412 = ~i_RtoB_ACK0 & ~n22411;
  assign n22413 = ~n22400 & ~n22412;
  assign n22414 = ~controllable_DEQ & ~n22413;
  assign n22415 = ~n22410 & ~n22414;
  assign n22416 = ~i_FULL & ~n22415;
  assign n22417 = ~n22406 & ~n22416;
  assign n22418 = i_nEMPTY & ~n22417;
  assign n22419 = ~n10120 & ~n19488;
  assign n22420 = ~i_RtoB_ACK0 & ~n22419;
  assign n22421 = ~n15548 & ~n22420;
  assign n22422 = controllable_DEQ & ~n22421;
  assign n22423 = ~n10078 & ~n17030;
  assign n22424 = i_RtoB_ACK0 & ~n22423;
  assign n22425 = ~n9726 & ~n19493;
  assign n22426 = ~i_RtoB_ACK0 & ~n22425;
  assign n22427 = ~n22424 & ~n22426;
  assign n22428 = ~controllable_DEQ & ~n22427;
  assign n22429 = ~n22422 & ~n22428;
  assign n22430 = i_FULL & ~n22429;
  assign n22431 = ~n10130 & ~n19504;
  assign n22432 = ~i_RtoB_ACK0 & ~n22431;
  assign n22433 = ~n15569 & ~n22432;
  assign n22434 = controllable_DEQ & ~n22433;
  assign n22435 = ~controllable_DEQ & ~n22397;
  assign n22436 = ~n22434 & ~n22435;
  assign n22437 = ~i_FULL & ~n22436;
  assign n22438 = ~n22430 & ~n22437;
  assign n22439 = ~i_nEMPTY & ~n22438;
  assign n22440 = ~n22418 & ~n22439;
  assign n22441 = ~controllable_BtoS_ACK0 & ~n22440;
  assign n22442 = ~n22392 & ~n22441;
  assign n22443 = n4465 & ~n22442;
  assign n22444 = ~n10145 & ~n17050;
  assign n22445 = i_RtoB_ACK0 & ~n22444;
  assign n22446 = ~n10155 & ~n19518;
  assign n22447 = ~i_RtoB_ACK0 & ~n22446;
  assign n22448 = ~n22445 & ~n22447;
  assign n22449 = controllable_DEQ & ~n22448;
  assign n22450 = ~n10161 & ~n17058;
  assign n22451 = i_RtoB_ACK0 & ~n22450;
  assign n22452 = ~n9817 & ~n19523;
  assign n22453 = ~i_RtoB_ACK0 & ~n22452;
  assign n22454 = ~n22451 & ~n22453;
  assign n22455 = ~controllable_DEQ & ~n22454;
  assign n22456 = ~n22449 & ~n22455;
  assign n22457 = i_nEMPTY & ~n22456;
  assign n22458 = ~n10169 & ~n19530;
  assign n22459 = ~i_RtoB_ACK0 & ~n22458;
  assign n22460 = ~n15604 & ~n22459;
  assign n22461 = controllable_DEQ & ~n22460;
  assign n22462 = ~n10145 & ~n17068;
  assign n22463 = i_RtoB_ACK0 & ~n22462;
  assign n22464 = ~n9840 & ~n19535;
  assign n22465 = ~i_RtoB_ACK0 & ~n22464;
  assign n22466 = ~n22463 & ~n22465;
  assign n22467 = ~controllable_DEQ & ~n22466;
  assign n22468 = ~n22461 & ~n22467;
  assign n22469 = i_FULL & ~n22468;
  assign n22470 = ~n10179 & ~n19542;
  assign n22471 = ~i_RtoB_ACK0 & ~n22470;
  assign n22472 = ~n15619 & ~n22471;
  assign n22473 = controllable_DEQ & ~n22472;
  assign n22474 = ~controllable_DEQ & ~n22448;
  assign n22475 = ~n22473 & ~n22474;
  assign n22476 = ~i_FULL & ~n22475;
  assign n22477 = ~n22469 & ~n22476;
  assign n22478 = ~i_nEMPTY & ~n22477;
  assign n22479 = ~n22457 & ~n22478;
  assign n22480 = controllable_BtoS_ACK0 & ~n22479;
  assign n22481 = ~n10192 & ~n17086;
  assign n22482 = i_RtoB_ACK0 & ~n22481;
  assign n22483 = ~n10200 & ~n19554;
  assign n22484 = ~i_RtoB_ACK0 & ~n22483;
  assign n22485 = ~n22482 & ~n22484;
  assign n22486 = controllable_DEQ & ~n22485;
  assign n22487 = ~n10206 & ~n17094;
  assign n22488 = i_RtoB_ACK0 & ~n22487;
  assign n22489 = ~n9917 & ~n19559;
  assign n22490 = ~i_RtoB_ACK0 & ~n22489;
  assign n22491 = ~n22488 & ~n22490;
  assign n22492 = ~controllable_DEQ & ~n22491;
  assign n22493 = ~n22486 & ~n22492;
  assign n22494 = i_FULL & ~n22493;
  assign n22495 = ~n10216 & ~n19566;
  assign n22496 = ~i_RtoB_ACK0 & ~n22495;
  assign n22497 = ~n22482 & ~n22496;
  assign n22498 = controllable_DEQ & ~n22497;
  assign n22499 = ~n9939 & ~n19571;
  assign n22500 = ~i_RtoB_ACK0 & ~n22499;
  assign n22501 = ~n22488 & ~n22500;
  assign n22502 = ~controllable_DEQ & ~n22501;
  assign n22503 = ~n22498 & ~n22502;
  assign n22504 = ~i_FULL & ~n22503;
  assign n22505 = ~n22494 & ~n22504;
  assign n22506 = i_nEMPTY & ~n22505;
  assign n22507 = ~n10228 & ~n19580;
  assign n22508 = ~i_RtoB_ACK0 & ~n22507;
  assign n22509 = ~n15680 & ~n22508;
  assign n22510 = controllable_DEQ & ~n22509;
  assign n22511 = ~n10192 & ~n17112;
  assign n22512 = i_RtoB_ACK0 & ~n22511;
  assign n22513 = ~n9965 & ~n19585;
  assign n22514 = ~i_RtoB_ACK0 & ~n22513;
  assign n22515 = ~n22512 & ~n22514;
  assign n22516 = ~controllable_DEQ & ~n22515;
  assign n22517 = ~n22510 & ~n22516;
  assign n22518 = i_FULL & ~n22517;
  assign n22519 = ~n10238 & ~n19592;
  assign n22520 = ~i_RtoB_ACK0 & ~n22519;
  assign n22521 = ~n15701 & ~n22520;
  assign n22522 = controllable_DEQ & ~n22521;
  assign n22523 = ~controllable_DEQ & ~n22485;
  assign n22524 = ~n22522 & ~n22523;
  assign n22525 = ~i_FULL & ~n22524;
  assign n22526 = ~n22518 & ~n22525;
  assign n22527 = ~i_nEMPTY & ~n22526;
  assign n22528 = ~n22506 & ~n22527;
  assign n22529 = ~controllable_BtoS_ACK0 & ~n22528;
  assign n22530 = ~n22480 & ~n22529;
  assign n22531 = ~n4465 & ~n22530;
  assign n22532 = ~n22443 & ~n22531;
  assign n22533 = i_StoB_REQ10 & ~n22532;
  assign n22534 = ~n22341 & ~n22533;
  assign n22535 = ~controllable_BtoS_ACK10 & ~n22534;
  assign n22536 = ~n22343 & ~n22535;
  assign n22537 = n4464 & ~n22536;
  assign n22538 = ~n10261 & ~n14741;
  assign n22539 = i_RtoB_ACK0 & ~n22538;
  assign n22540 = ~n10271 & ~n15732;
  assign n22541 = ~i_RtoB_ACK0 & ~n22540;
  assign n22542 = ~n22539 & ~n22541;
  assign n22543 = controllable_DEQ & ~n22542;
  assign n22544 = ~n10280 & ~n14757;
  assign n22545 = i_RtoB_ACK0 & ~n22544;
  assign n22546 = ~n10286 & ~n15749;
  assign n22547 = ~i_RtoB_ACK0 & ~n22546;
  assign n22548 = ~n22545 & ~n22547;
  assign n22549 = ~controllable_DEQ & ~n22548;
  assign n22550 = ~n22543 & ~n22549;
  assign n22551 = i_FULL & ~n22550;
  assign n22552 = ~n10296 & ~n15732;
  assign n22553 = ~i_RtoB_ACK0 & ~n22552;
  assign n22554 = ~n22539 & ~n22553;
  assign n22555 = controllable_DEQ & ~n22554;
  assign n22556 = ~n10304 & ~n15749;
  assign n22557 = ~i_RtoB_ACK0 & ~n22556;
  assign n22558 = ~n22545 & ~n22557;
  assign n22559 = ~controllable_DEQ & ~n22558;
  assign n22560 = ~n22555 & ~n22559;
  assign n22561 = ~i_FULL & ~n22560;
  assign n22562 = ~n22551 & ~n22561;
  assign n22563 = i_nEMPTY & ~n22562;
  assign n22564 = ~n10314 & ~n15758;
  assign n22565 = ~i_RtoB_ACK0 & ~n22564;
  assign n22566 = ~i_RtoB_ACK0 & ~n22565;
  assign n22567 = controllable_DEQ & ~n22566;
  assign n22568 = ~n10323 & ~n15768;
  assign n22569 = ~i_RtoB_ACK0 & ~n22568;
  assign n22570 = ~n22539 & ~n22569;
  assign n22571 = ~controllable_DEQ & ~n22570;
  assign n22572 = ~n22567 & ~n22571;
  assign n22573 = i_FULL & ~n22572;
  assign n22574 = ~n10331 & ~n15777;
  assign n22575 = ~i_RtoB_ACK0 & ~n22574;
  assign n22576 = ~i_RtoB_ACK0 & ~n22575;
  assign n22577 = controllable_DEQ & ~n22576;
  assign n22578 = ~n10341 & ~n15732;
  assign n22579 = ~i_RtoB_ACK0 & ~n22578;
  assign n22580 = ~n22539 & ~n22579;
  assign n22581 = ~controllable_DEQ & ~n22580;
  assign n22582 = ~n22577 & ~n22581;
  assign n22583 = ~i_FULL & ~n22582;
  assign n22584 = ~n22573 & ~n22583;
  assign n22585 = ~i_nEMPTY & ~n22584;
  assign n22586 = ~n22563 & ~n22585;
  assign n22587 = controllable_BtoS_ACK0 & ~n22586;
  assign n22588 = ~n10355 & ~n16723;
  assign n22589 = i_RtoB_ACK0 & ~n22588;
  assign n22590 = ~n10365 & ~n15807;
  assign n22591 = ~i_RtoB_ACK0 & ~n22590;
  assign n22592 = ~n22589 & ~n22591;
  assign n22593 = controllable_DEQ & ~n22592;
  assign n22594 = ~n10374 & ~n16729;
  assign n22595 = i_RtoB_ACK0 & ~n22594;
  assign n22596 = ~n10380 & ~n15824;
  assign n22597 = ~i_RtoB_ACK0 & ~n22596;
  assign n22598 = ~n22595 & ~n22597;
  assign n22599 = ~controllable_DEQ & ~n22598;
  assign n22600 = ~n22593 & ~n22599;
  assign n22601 = i_FULL & ~n22600;
  assign n22602 = ~n10390 & ~n15807;
  assign n22603 = ~i_RtoB_ACK0 & ~n22602;
  assign n22604 = ~n22589 & ~n22603;
  assign n22605 = controllable_DEQ & ~n22604;
  assign n22606 = ~n10398 & ~n15824;
  assign n22607 = ~i_RtoB_ACK0 & ~n22606;
  assign n22608 = ~n22595 & ~n22607;
  assign n22609 = ~controllable_DEQ & ~n22608;
  assign n22610 = ~n22605 & ~n22609;
  assign n22611 = ~i_FULL & ~n22610;
  assign n22612 = ~n22601 & ~n22611;
  assign n22613 = i_nEMPTY & ~n22612;
  assign n22614 = ~n10408 & ~n15833;
  assign n22615 = ~i_RtoB_ACK0 & ~n22614;
  assign n22616 = ~i_RtoB_ACK0 & ~n22615;
  assign n22617 = controllable_DEQ & ~n22616;
  assign n22618 = ~n10417 & ~n15843;
  assign n22619 = ~i_RtoB_ACK0 & ~n22618;
  assign n22620 = ~n22589 & ~n22619;
  assign n22621 = ~controllable_DEQ & ~n22620;
  assign n22622 = ~n22617 & ~n22621;
  assign n22623 = i_FULL & ~n22622;
  assign n22624 = ~n10425 & ~n15852;
  assign n22625 = ~i_RtoB_ACK0 & ~n22624;
  assign n22626 = ~i_RtoB_ACK0 & ~n22625;
  assign n22627 = controllable_DEQ & ~n22626;
  assign n22628 = ~n10435 & ~n15807;
  assign n22629 = ~i_RtoB_ACK0 & ~n22628;
  assign n22630 = ~n22589 & ~n22629;
  assign n22631 = ~controllable_DEQ & ~n22630;
  assign n22632 = ~n22627 & ~n22631;
  assign n22633 = ~i_FULL & ~n22632;
  assign n22634 = ~n22623 & ~n22633;
  assign n22635 = ~i_nEMPTY & ~n22634;
  assign n22636 = ~n22613 & ~n22635;
  assign n22637 = ~controllable_BtoS_ACK0 & ~n22636;
  assign n22638 = ~n22587 & ~n22637;
  assign n22639 = n4465 & ~n22638;
  assign n22640 = ~n21013 & ~n22637;
  assign n22641 = ~n4465 & ~n22640;
  assign n22642 = ~n22639 & ~n22641;
  assign n22643 = i_StoB_REQ10 & ~n22642;
  assign n22644 = ~n10464 & ~n17188;
  assign n22645 = i_RtoB_ACK0 & ~n22644;
  assign n22646 = ~n10482 & ~n15889;
  assign n22647 = ~i_RtoB_ACK0 & ~n22646;
  assign n22648 = ~n22645 & ~n22647;
  assign n22649 = controllable_DEQ & ~n22648;
  assign n22650 = ~n10491 & ~n17196;
  assign n22651 = i_RtoB_ACK0 & ~n22650;
  assign n22652 = ~n10500 & ~n15908;
  assign n22653 = ~i_RtoB_ACK0 & ~n22652;
  assign n22654 = ~n22651 & ~n22653;
  assign n22655 = ~controllable_DEQ & ~n22654;
  assign n22656 = ~n22649 & ~n22655;
  assign n22657 = i_FULL & ~n22656;
  assign n22658 = ~n10514 & ~n15927;
  assign n22659 = ~i_RtoB_ACK0 & ~n22658;
  assign n22660 = ~n22645 & ~n22659;
  assign n22661 = controllable_DEQ & ~n22660;
  assign n22662 = ~n10526 & ~n15943;
  assign n22663 = ~i_RtoB_ACK0 & ~n22662;
  assign n22664 = ~n22651 & ~n22663;
  assign n22665 = ~controllable_DEQ & ~n22664;
  assign n22666 = ~n22661 & ~n22665;
  assign n22667 = ~i_FULL & ~n22666;
  assign n22668 = ~n22657 & ~n22667;
  assign n22669 = i_nEMPTY & ~n22668;
  assign n22670 = ~n10540 & ~n15964;
  assign n22671 = ~i_RtoB_ACK0 & ~n22670;
  assign n22672 = ~n15960 & ~n22671;
  assign n22673 = controllable_DEQ & ~n22672;
  assign n22674 = ~n10464 & ~n17214;
  assign n22675 = i_RtoB_ACK0 & ~n22674;
  assign n22676 = ~n10552 & ~n15980;
  assign n22677 = ~i_RtoB_ACK0 & ~n22676;
  assign n22678 = ~n22675 & ~n22677;
  assign n22679 = ~controllable_DEQ & ~n22678;
  assign n22680 = ~n22673 & ~n22679;
  assign n22681 = i_FULL & ~n22680;
  assign n22682 = ~n10562 & ~n15999;
  assign n22683 = ~i_RtoB_ACK0 & ~n22682;
  assign n22684 = ~n15995 & ~n22683;
  assign n22685 = controllable_DEQ & ~n22684;
  assign n22686 = ~n10572 & ~n15889;
  assign n22687 = ~i_RtoB_ACK0 & ~n22686;
  assign n22688 = ~n22645 & ~n22687;
  assign n22689 = ~controllable_DEQ & ~n22688;
  assign n22690 = ~n22685 & ~n22689;
  assign n22691 = ~i_FULL & ~n22690;
  assign n22692 = ~n22681 & ~n22691;
  assign n22693 = ~i_nEMPTY & ~n22692;
  assign n22694 = ~n22669 & ~n22693;
  assign n22695 = controllable_BtoS_ACK0 & ~n22694;
  assign n22696 = ~n10594 & ~n17233;
  assign n22697 = i_RtoB_ACK0 & ~n22696;
  assign n22698 = ~n10609 & ~n16031;
  assign n22699 = ~i_RtoB_ACK0 & ~n22698;
  assign n22700 = ~n22697 & ~n22699;
  assign n22701 = controllable_DEQ & ~n22700;
  assign n22702 = ~n10618 & ~n17241;
  assign n22703 = i_RtoB_ACK0 & ~n22702;
  assign n22704 = ~n10627 & ~n16050;
  assign n22705 = ~i_RtoB_ACK0 & ~n22704;
  assign n22706 = ~n22703 & ~n22705;
  assign n22707 = ~controllable_DEQ & ~n22706;
  assign n22708 = ~n22701 & ~n22707;
  assign n22709 = i_FULL & ~n22708;
  assign n22710 = ~n10641 & ~n16069;
  assign n22711 = ~i_RtoB_ACK0 & ~n22710;
  assign n22712 = ~n22697 & ~n22711;
  assign n22713 = controllable_DEQ & ~n22712;
  assign n22714 = ~n10653 & ~n16085;
  assign n22715 = ~i_RtoB_ACK0 & ~n22714;
  assign n22716 = ~n22703 & ~n22715;
  assign n22717 = ~controllable_DEQ & ~n22716;
  assign n22718 = ~n22713 & ~n22717;
  assign n22719 = ~i_FULL & ~n22718;
  assign n22720 = ~n22709 & ~n22719;
  assign n22721 = i_nEMPTY & ~n22720;
  assign n22722 = ~n10667 & ~n16106;
  assign n22723 = ~i_RtoB_ACK0 & ~n22722;
  assign n22724 = ~n16102 & ~n22723;
  assign n22725 = controllable_DEQ & ~n22724;
  assign n22726 = ~n10594 & ~n17259;
  assign n22727 = i_RtoB_ACK0 & ~n22726;
  assign n22728 = ~n10679 & ~n16122;
  assign n22729 = ~i_RtoB_ACK0 & ~n22728;
  assign n22730 = ~n22727 & ~n22729;
  assign n22731 = ~controllable_DEQ & ~n22730;
  assign n22732 = ~n22725 & ~n22731;
  assign n22733 = i_FULL & ~n22732;
  assign n22734 = ~n10689 & ~n16141;
  assign n22735 = ~i_RtoB_ACK0 & ~n22734;
  assign n22736 = ~n16137 & ~n22735;
  assign n22737 = controllable_DEQ & ~n22736;
  assign n22738 = ~n10699 & ~n16031;
  assign n22739 = ~i_RtoB_ACK0 & ~n22738;
  assign n22740 = ~n22697 & ~n22739;
  assign n22741 = ~controllable_DEQ & ~n22740;
  assign n22742 = ~n22737 & ~n22741;
  assign n22743 = ~i_FULL & ~n22742;
  assign n22744 = ~n22733 & ~n22743;
  assign n22745 = ~i_nEMPTY & ~n22744;
  assign n22746 = ~n22721 & ~n22745;
  assign n22747 = ~controllable_BtoS_ACK0 & ~n22746;
  assign n22748 = ~n22695 & ~n22747;
  assign n22749 = n4465 & ~n22748;
  assign n22750 = ~n10715 & ~n17280;
  assign n22751 = i_RtoB_ACK0 & ~n22750;
  assign n22752 = ~n10723 & ~n16175;
  assign n22753 = ~i_RtoB_ACK0 & ~n22752;
  assign n22754 = ~n22751 & ~n22753;
  assign n22755 = controllable_DEQ & ~n22754;
  assign n22756 = ~n10732 & ~n17288;
  assign n22757 = i_RtoB_ACK0 & ~n22756;
  assign n22758 = ~n10738 & ~n16194;
  assign n22759 = ~i_RtoB_ACK0 & ~n22758;
  assign n22760 = ~n22757 & ~n22759;
  assign n22761 = ~controllable_DEQ & ~n22760;
  assign n22762 = ~n22755 & ~n22761;
  assign n22763 = i_nEMPTY & ~n22762;
  assign n22764 = ~n10746 & ~n16204;
  assign n22765 = ~i_RtoB_ACK0 & ~n22764;
  assign n22766 = ~n15217 & ~n22765;
  assign n22767 = controllable_DEQ & ~n22766;
  assign n22768 = ~n10715 & ~n17298;
  assign n22769 = i_RtoB_ACK0 & ~n22768;
  assign n22770 = ~n10754 & ~n16220;
  assign n22771 = ~i_RtoB_ACK0 & ~n22770;
  assign n22772 = ~n22769 & ~n22771;
  assign n22773 = ~controllable_DEQ & ~n22772;
  assign n22774 = ~n22767 & ~n22773;
  assign n22775 = i_FULL & ~n22774;
  assign n22776 = ~n10762 & ~n16230;
  assign n22777 = ~i_RtoB_ACK0 & ~n22776;
  assign n22778 = ~n15245 & ~n22777;
  assign n22779 = controllable_DEQ & ~n22778;
  assign n22780 = ~n10770 & ~n16175;
  assign n22781 = ~i_RtoB_ACK0 & ~n22780;
  assign n22782 = ~n22751 & ~n22781;
  assign n22783 = ~controllable_DEQ & ~n22782;
  assign n22784 = ~n22779 & ~n22783;
  assign n22785 = ~i_FULL & ~n22784;
  assign n22786 = ~n22775 & ~n22785;
  assign n22787 = ~i_nEMPTY & ~n22786;
  assign n22788 = ~n22763 & ~n22787;
  assign n22789 = controllable_BtoS_ACK0 & ~n22788;
  assign n22790 = ~n10784 & ~n17317;
  assign n22791 = i_RtoB_ACK0 & ~n22790;
  assign n22792 = ~n10794 & ~n16262;
  assign n22793 = ~i_RtoB_ACK0 & ~n22792;
  assign n22794 = ~n22791 & ~n22793;
  assign n22795 = controllable_DEQ & ~n22794;
  assign n22796 = ~n10802 & ~n17325;
  assign n22797 = i_RtoB_ACK0 & ~n22796;
  assign n22798 = ~n10808 & ~n16281;
  assign n22799 = ~i_RtoB_ACK0 & ~n22798;
  assign n22800 = ~n22797 & ~n22799;
  assign n22801 = ~controllable_DEQ & ~n22800;
  assign n22802 = ~n22795 & ~n22801;
  assign n22803 = i_FULL & ~n22802;
  assign n22804 = ~n10820 & ~n16300;
  assign n22805 = ~i_RtoB_ACK0 & ~n22804;
  assign n22806 = ~n22791 & ~n22805;
  assign n22807 = controllable_DEQ & ~n22806;
  assign n22808 = ~n10830 & ~n16316;
  assign n22809 = ~i_RtoB_ACK0 & ~n22808;
  assign n22810 = ~n22797 & ~n22809;
  assign n22811 = ~controllable_DEQ & ~n22810;
  assign n22812 = ~n22807 & ~n22811;
  assign n22813 = ~i_FULL & ~n22812;
  assign n22814 = ~n22803 & ~n22813;
  assign n22815 = i_nEMPTY & ~n22814;
  assign n22816 = ~n10840 & ~n16337;
  assign n22817 = ~i_RtoB_ACK0 & ~n22816;
  assign n22818 = ~n16333 & ~n22817;
  assign n22819 = controllable_DEQ & ~n22818;
  assign n22820 = ~n10784 & ~n17343;
  assign n22821 = i_RtoB_ACK0 & ~n22820;
  assign n22822 = ~n10848 & ~n16353;
  assign n22823 = ~i_RtoB_ACK0 & ~n22822;
  assign n22824 = ~n22821 & ~n22823;
  assign n22825 = ~controllable_DEQ & ~n22824;
  assign n22826 = ~n22819 & ~n22825;
  assign n22827 = i_FULL & ~n22826;
  assign n22828 = ~n10856 & ~n16372;
  assign n22829 = ~i_RtoB_ACK0 & ~n22828;
  assign n22830 = ~n16368 & ~n22829;
  assign n22831 = controllable_DEQ & ~n22830;
  assign n22832 = ~n10864 & ~n16262;
  assign n22833 = ~i_RtoB_ACK0 & ~n22832;
  assign n22834 = ~n22791 & ~n22833;
  assign n22835 = ~controllable_DEQ & ~n22834;
  assign n22836 = ~n22831 & ~n22835;
  assign n22837 = ~i_FULL & ~n22836;
  assign n22838 = ~n22827 & ~n22837;
  assign n22839 = ~i_nEMPTY & ~n22838;
  assign n22840 = ~n22815 & ~n22839;
  assign n22841 = ~controllable_BtoS_ACK0 & ~n22840;
  assign n22842 = ~n22789 & ~n22841;
  assign n22843 = ~n4465 & ~n22842;
  assign n22844 = ~n22749 & ~n22843;
  assign n22845 = ~i_StoB_REQ10 & ~n22844;
  assign n22846 = ~n22643 & ~n22845;
  assign n22847 = controllable_BtoS_ACK10 & ~n22846;
  assign n22848 = ~n10884 & ~n17368;
  assign n22849 = i_RtoB_ACK0 & ~n22848;
  assign n22850 = ~n10894 & ~n20002;
  assign n22851 = ~i_RtoB_ACK0 & ~n22850;
  assign n22852 = ~n22849 & ~n22851;
  assign n22853 = controllable_DEQ & ~n22852;
  assign n22854 = ~n10902 & ~n17376;
  assign n22855 = i_RtoB_ACK0 & ~n22854;
  assign n22856 = ~n10500 & ~n20011;
  assign n22857 = ~i_RtoB_ACK0 & ~n22856;
  assign n22858 = ~n22855 & ~n22857;
  assign n22859 = ~controllable_DEQ & ~n22858;
  assign n22860 = ~n22853 & ~n22859;
  assign n22861 = i_FULL & ~n22860;
  assign n22862 = ~n10914 & ~n20022;
  assign n22863 = ~i_RtoB_ACK0 & ~n22862;
  assign n22864 = ~n22849 & ~n22863;
  assign n22865 = controllable_DEQ & ~n22864;
  assign n22866 = ~n10526 & ~n20027;
  assign n22867 = ~i_RtoB_ACK0 & ~n22866;
  assign n22868 = ~n22855 & ~n22867;
  assign n22869 = ~controllable_DEQ & ~n22868;
  assign n22870 = ~n22865 & ~n22869;
  assign n22871 = ~i_FULL & ~n22870;
  assign n22872 = ~n22861 & ~n22871;
  assign n22873 = i_nEMPTY & ~n22872;
  assign n22874 = ~n10926 & ~n20040;
  assign n22875 = ~i_RtoB_ACK0 & ~n22874;
  assign n22876 = ~n16447 & ~n22875;
  assign n22877 = controllable_DEQ & ~n22876;
  assign n22878 = ~n10884 & ~n17394;
  assign n22879 = i_RtoB_ACK0 & ~n22878;
  assign n22880 = ~n10552 & ~n20045;
  assign n22881 = ~i_RtoB_ACK0 & ~n22880;
  assign n22882 = ~n22879 & ~n22881;
  assign n22883 = ~controllable_DEQ & ~n22882;
  assign n22884 = ~n22877 & ~n22883;
  assign n22885 = i_FULL & ~n22884;
  assign n22886 = ~n10936 & ~n20056;
  assign n22887 = ~i_RtoB_ACK0 & ~n22886;
  assign n22888 = ~n16468 & ~n22887;
  assign n22889 = controllable_DEQ & ~n22888;
  assign n22890 = ~controllable_DEQ & ~n22852;
  assign n22891 = ~n22889 & ~n22890;
  assign n22892 = ~i_FULL & ~n22891;
  assign n22893 = ~n22885 & ~n22892;
  assign n22894 = ~i_nEMPTY & ~n22893;
  assign n22895 = ~n22873 & ~n22894;
  assign n22896 = controllable_BtoS_ACK0 & ~n22895;
  assign n22897 = ~n10951 & ~n17412;
  assign n22898 = i_RtoB_ACK0 & ~n22897;
  assign n22899 = ~n10961 & ~n20068;
  assign n22900 = ~i_RtoB_ACK0 & ~n22899;
  assign n22901 = ~n22898 & ~n22900;
  assign n22902 = controllable_DEQ & ~n22901;
  assign n22903 = ~n10969 & ~n17420;
  assign n22904 = i_RtoB_ACK0 & ~n22903;
  assign n22905 = ~n10627 & ~n20073;
  assign n22906 = ~i_RtoB_ACK0 & ~n22905;
  assign n22907 = ~n22904 & ~n22906;
  assign n22908 = ~controllable_DEQ & ~n22907;
  assign n22909 = ~n22902 & ~n22908;
  assign n22910 = i_FULL & ~n22909;
  assign n22911 = ~n10981 & ~n20080;
  assign n22912 = ~i_RtoB_ACK0 & ~n22911;
  assign n22913 = ~n22898 & ~n22912;
  assign n22914 = controllable_DEQ & ~n22913;
  assign n22915 = ~n10653 & ~n20085;
  assign n22916 = ~i_RtoB_ACK0 & ~n22915;
  assign n22917 = ~n22904 & ~n22916;
  assign n22918 = ~controllable_DEQ & ~n22917;
  assign n22919 = ~n22914 & ~n22918;
  assign n22920 = ~i_FULL & ~n22919;
  assign n22921 = ~n22910 & ~n22920;
  assign n22922 = i_nEMPTY & ~n22921;
  assign n22923 = ~n10993 & ~n20094;
  assign n22924 = ~i_RtoB_ACK0 & ~n22923;
  assign n22925 = ~n16529 & ~n22924;
  assign n22926 = controllable_DEQ & ~n22925;
  assign n22927 = ~n10951 & ~n17438;
  assign n22928 = i_RtoB_ACK0 & ~n22927;
  assign n22929 = ~n10679 & ~n20099;
  assign n22930 = ~i_RtoB_ACK0 & ~n22929;
  assign n22931 = ~n22928 & ~n22930;
  assign n22932 = ~controllable_DEQ & ~n22931;
  assign n22933 = ~n22926 & ~n22932;
  assign n22934 = i_FULL & ~n22933;
  assign n22935 = ~n11003 & ~n20106;
  assign n22936 = ~i_RtoB_ACK0 & ~n22935;
  assign n22937 = ~n16550 & ~n22936;
  assign n22938 = controllable_DEQ & ~n22937;
  assign n22939 = ~controllable_DEQ & ~n22901;
  assign n22940 = ~n22938 & ~n22939;
  assign n22941 = ~i_FULL & ~n22940;
  assign n22942 = ~n22934 & ~n22941;
  assign n22943 = ~i_nEMPTY & ~n22942;
  assign n22944 = ~n22922 & ~n22943;
  assign n22945 = ~controllable_BtoS_ACK0 & ~n22944;
  assign n22946 = ~n22896 & ~n22945;
  assign n22947 = n4465 & ~n22946;
  assign n22948 = ~n11018 & ~n17050;
  assign n22949 = i_RtoB_ACK0 & ~n22948;
  assign n22950 = ~n11024 & ~n20120;
  assign n22951 = ~i_RtoB_ACK0 & ~n22950;
  assign n22952 = ~n22949 & ~n22951;
  assign n22953 = controllable_DEQ & ~n22952;
  assign n22954 = ~n11030 & ~n17058;
  assign n22955 = i_RtoB_ACK0 & ~n22954;
  assign n22956 = ~n10738 & ~n20125;
  assign n22957 = ~i_RtoB_ACK0 & ~n22956;
  assign n22958 = ~n22955 & ~n22957;
  assign n22959 = ~controllable_DEQ & ~n22958;
  assign n22960 = ~n22953 & ~n22959;
  assign n22961 = i_nEMPTY & ~n22960;
  assign n22962 = ~n11038 & ~n20132;
  assign n22963 = ~i_RtoB_ACK0 & ~n22962;
  assign n22964 = ~n15604 & ~n22963;
  assign n22965 = controllable_DEQ & ~n22964;
  assign n22966 = ~n11018 & ~n17068;
  assign n22967 = i_RtoB_ACK0 & ~n22966;
  assign n22968 = ~n10754 & ~n20137;
  assign n22969 = ~i_RtoB_ACK0 & ~n22968;
  assign n22970 = ~n22967 & ~n22969;
  assign n22971 = ~controllable_DEQ & ~n22970;
  assign n22972 = ~n22965 & ~n22971;
  assign n22973 = i_FULL & ~n22972;
  assign n22974 = ~n11048 & ~n20144;
  assign n22975 = ~i_RtoB_ACK0 & ~n22974;
  assign n22976 = ~n15619 & ~n22975;
  assign n22977 = controllable_DEQ & ~n22976;
  assign n22978 = ~controllable_DEQ & ~n22952;
  assign n22979 = ~n22977 & ~n22978;
  assign n22980 = ~i_FULL & ~n22979;
  assign n22981 = ~n22973 & ~n22980;
  assign n22982 = ~i_nEMPTY & ~n22981;
  assign n22983 = ~n22961 & ~n22982;
  assign n22984 = controllable_BtoS_ACK0 & ~n22983;
  assign n22985 = ~n11061 & ~n17481;
  assign n22986 = i_RtoB_ACK0 & ~n22985;
  assign n22987 = ~n11069 & ~n20156;
  assign n22988 = ~i_RtoB_ACK0 & ~n22987;
  assign n22989 = ~n22986 & ~n22988;
  assign n22990 = controllable_DEQ & ~n22989;
  assign n22991 = ~n11075 & ~n17489;
  assign n22992 = i_RtoB_ACK0 & ~n22991;
  assign n22993 = ~n10808 & ~n20161;
  assign n22994 = ~i_RtoB_ACK0 & ~n22993;
  assign n22995 = ~n22992 & ~n22994;
  assign n22996 = ~controllable_DEQ & ~n22995;
  assign n22997 = ~n22990 & ~n22996;
  assign n22998 = i_FULL & ~n22997;
  assign n22999 = ~n11085 & ~n20168;
  assign n23000 = ~i_RtoB_ACK0 & ~n22999;
  assign n23001 = ~n22986 & ~n23000;
  assign n23002 = controllable_DEQ & ~n23001;
  assign n23003 = ~n10830 & ~n20173;
  assign n23004 = ~i_RtoB_ACK0 & ~n23003;
  assign n23005 = ~n22992 & ~n23004;
  assign n23006 = ~controllable_DEQ & ~n23005;
  assign n23007 = ~n23002 & ~n23006;
  assign n23008 = ~i_FULL & ~n23007;
  assign n23009 = ~n22998 & ~n23008;
  assign n23010 = i_nEMPTY & ~n23009;
  assign n23011 = ~n11097 & ~n20182;
  assign n23012 = ~i_RtoB_ACK0 & ~n23011;
  assign n23013 = ~n16656 & ~n23012;
  assign n23014 = controllable_DEQ & ~n23013;
  assign n23015 = ~n11061 & ~n17507;
  assign n23016 = i_RtoB_ACK0 & ~n23015;
  assign n23017 = ~n10848 & ~n20187;
  assign n23018 = ~i_RtoB_ACK0 & ~n23017;
  assign n23019 = ~n23016 & ~n23018;
  assign n23020 = ~controllable_DEQ & ~n23019;
  assign n23021 = ~n23014 & ~n23020;
  assign n23022 = i_FULL & ~n23021;
  assign n23023 = ~n11107 & ~n20194;
  assign n23024 = ~i_RtoB_ACK0 & ~n23023;
  assign n23025 = ~n16677 & ~n23024;
  assign n23026 = controllable_DEQ & ~n23025;
  assign n23027 = ~controllable_DEQ & ~n22989;
  assign n23028 = ~n23026 & ~n23027;
  assign n23029 = ~i_FULL & ~n23028;
  assign n23030 = ~n23022 & ~n23029;
  assign n23031 = ~i_nEMPTY & ~n23030;
  assign n23032 = ~n23010 & ~n23031;
  assign n23033 = ~controllable_BtoS_ACK0 & ~n23032;
  assign n23034 = ~n22984 & ~n23033;
  assign n23035 = ~n4465 & ~n23034;
  assign n23036 = ~n22947 & ~n23035;
  assign n23037 = i_StoB_REQ10 & ~n23036;
  assign n23038 = ~n22845 & ~n23037;
  assign n23039 = ~controllable_BtoS_ACK10 & ~n23038;
  assign n23040 = ~n22847 & ~n23039;
  assign n23041 = ~n4464 & ~n23040;
  assign n23042 = ~n22537 & ~n23041;
  assign n23043 = ~n4463 & ~n23042;
  assign n23044 = ~n21983 & ~n23043;
  assign n23045 = n4462 & ~n23044;
  assign n23046 = ~n11147 & ~n17536;
  assign n23047 = i_RtoB_ACK0 & ~n23046;
  assign n23048 = ~n11160 & ~n17545;
  assign n23049 = ~i_RtoB_ACK0 & ~n23048;
  assign n23050 = ~n23047 & ~n23049;
  assign n23051 = controllable_DEQ & ~n23050;
  assign n23052 = ~n11170 & ~n17553;
  assign n23053 = i_RtoB_ACK0 & ~n23052;
  assign n23054 = ~n11173 & ~n17562;
  assign n23055 = ~i_RtoB_ACK0 & ~n23054;
  assign n23056 = ~n23053 & ~n23055;
  assign n23057 = ~controllable_DEQ & ~n23056;
  assign n23058 = ~n23051 & ~n23057;
  assign n23059 = i_nEMPTY & ~n23058;
  assign n23060 = ~n11190 & ~n17571;
  assign n23061 = ~i_RtoB_ACK0 & ~n23060;
  assign n23062 = ~i_RtoB_ACK0 & ~n23061;
  assign n23063 = controllable_DEQ & ~n23062;
  assign n23064 = ~n11195 & ~n17581;
  assign n23065 = ~i_RtoB_ACK0 & ~n23064;
  assign n23066 = ~n23047 & ~n23065;
  assign n23067 = ~controllable_DEQ & ~n23066;
  assign n23068 = ~n23063 & ~n23067;
  assign n23069 = i_FULL & ~n23068;
  assign n23070 = ~n11205 & ~n17590;
  assign n23071 = ~i_RtoB_ACK0 & ~n23070;
  assign n23072 = ~i_RtoB_ACK0 & ~n23071;
  assign n23073 = controllable_DEQ & ~n23072;
  assign n23074 = ~n11210 & ~n17545;
  assign n23075 = ~i_RtoB_ACK0 & ~n23074;
  assign n23076 = ~n23047 & ~n23075;
  assign n23077 = ~controllable_DEQ & ~n23076;
  assign n23078 = ~n23073 & ~n23077;
  assign n23079 = ~i_FULL & ~n23078;
  assign n23080 = ~n23069 & ~n23079;
  assign n23081 = ~i_nEMPTY & ~n23080;
  assign n23082 = ~n23059 & ~n23081;
  assign n23083 = controllable_BtoS_ACK0 & ~n23082;
  assign n23084 = ~n21051 & ~n23083;
  assign n23085 = n4465 & ~n23084;
  assign n23086 = ~n21053 & ~n23085;
  assign n23087 = i_StoB_REQ10 & ~n23086;
  assign n23088 = ~n11232 & ~n17280;
  assign n23089 = i_RtoB_ACK0 & ~n23088;
  assign n23090 = ~n11240 & ~n17620;
  assign n23091 = ~i_RtoB_ACK0 & ~n23090;
  assign n23092 = ~n23089 & ~n23091;
  assign n23093 = controllable_DEQ & ~n23092;
  assign n23094 = ~n11250 & ~n17288;
  assign n23095 = i_RtoB_ACK0 & ~n23094;
  assign n23096 = ~n11253 & ~n17635;
  assign n23097 = ~i_RtoB_ACK0 & ~n23096;
  assign n23098 = ~n23095 & ~n23097;
  assign n23099 = ~controllable_DEQ & ~n23098;
  assign n23100 = ~n23093 & ~n23099;
  assign n23101 = i_nEMPTY & ~n23100;
  assign n23102 = ~n11265 & ~n17645;
  assign n23103 = ~i_RtoB_ACK0 & ~n23102;
  assign n23104 = ~n15217 & ~n23103;
  assign n23105 = controllable_DEQ & ~n23104;
  assign n23106 = ~n11232 & ~n17298;
  assign n23107 = i_RtoB_ACK0 & ~n23106;
  assign n23108 = ~n11270 & ~n17657;
  assign n23109 = ~i_RtoB_ACK0 & ~n23108;
  assign n23110 = ~n23107 & ~n23109;
  assign n23111 = ~controllable_DEQ & ~n23110;
  assign n23112 = ~n23105 & ~n23111;
  assign n23113 = i_FULL & ~n23112;
  assign n23114 = ~n11278 & ~n17667;
  assign n23115 = ~i_RtoB_ACK0 & ~n23114;
  assign n23116 = ~n15245 & ~n23115;
  assign n23117 = controllable_DEQ & ~n23116;
  assign n23118 = ~n11286 & ~n17620;
  assign n23119 = ~i_RtoB_ACK0 & ~n23118;
  assign n23120 = ~n23089 & ~n23119;
  assign n23121 = ~controllable_DEQ & ~n23120;
  assign n23122 = ~n23117 & ~n23121;
  assign n23123 = ~i_FULL & ~n23122;
  assign n23124 = ~n23113 & ~n23123;
  assign n23125 = ~i_nEMPTY & ~n23124;
  assign n23126 = ~n23101 & ~n23125;
  assign n23127 = controllable_BtoS_ACK0 & ~n23126;
  assign n23128 = ~n11307 & ~n17690;
  assign n23129 = i_RtoB_ACK0 & ~n23128;
  assign n23130 = ~n11319 & ~n17699;
  assign n23131 = ~i_RtoB_ACK0 & ~n23130;
  assign n23132 = ~n23129 & ~n23131;
  assign n23133 = controllable_DEQ & ~n23132;
  assign n23134 = ~n11330 & ~n17709;
  assign n23135 = i_RtoB_ACK0 & ~n23134;
  assign n23136 = ~n11333 & ~n17718;
  assign n23137 = ~i_RtoB_ACK0 & ~n23136;
  assign n23138 = ~n23135 & ~n23137;
  assign n23139 = ~controllable_DEQ & ~n23138;
  assign n23140 = ~n23133 & ~n23139;
  assign n23141 = i_nEMPTY & ~n23140;
  assign n23142 = ~n11347 & ~n17735;
  assign n23143 = ~i_RtoB_ACK0 & ~n23142;
  assign n23144 = ~n17731 & ~n23143;
  assign n23145 = controllable_DEQ & ~n23144;
  assign n23146 = ~n11307 & ~n17745;
  assign n23147 = i_RtoB_ACK0 & ~n23146;
  assign n23148 = ~n11352 & ~n17751;
  assign n23149 = ~i_RtoB_ACK0 & ~n23148;
  assign n23150 = ~n23147 & ~n23149;
  assign n23151 = ~controllable_DEQ & ~n23150;
  assign n23152 = ~n23145 & ~n23151;
  assign n23153 = i_FULL & ~n23152;
  assign n23154 = ~n11360 & ~n17768;
  assign n23155 = ~i_RtoB_ACK0 & ~n23154;
  assign n23156 = ~n17764 & ~n23155;
  assign n23157 = controllable_DEQ & ~n23156;
  assign n23158 = ~n11368 & ~n17699;
  assign n23159 = ~i_RtoB_ACK0 & ~n23158;
  assign n23160 = ~n23129 & ~n23159;
  assign n23161 = ~controllable_DEQ & ~n23160;
  assign n23162 = ~n23157 & ~n23161;
  assign n23163 = ~i_FULL & ~n23162;
  assign n23164 = ~n23153 & ~n23163;
  assign n23165 = ~i_nEMPTY & ~n23164;
  assign n23166 = ~n23141 & ~n23165;
  assign n23167 = ~controllable_BtoS_ACK0 & ~n23166;
  assign n23168 = ~n23127 & ~n23167;
  assign n23169 = ~i_StoB_REQ10 & ~n23168;
  assign n23170 = ~n23087 & ~n23169;
  assign n23171 = controllable_BtoS_ACK10 & ~n23170;
  assign n23172 = ~n11395 & ~n17795;
  assign n23173 = i_RtoB_ACK0 & ~n23172;
  assign n23174 = ~n11414 & ~n20366;
  assign n23175 = ~i_RtoB_ACK0 & ~n23174;
  assign n23176 = ~n23173 & ~n23175;
  assign n23177 = controllable_DEQ & ~n23176;
  assign n23178 = ~n11424 & ~n17807;
  assign n23179 = i_RtoB_ACK0 & ~n23178;
  assign n23180 = ~n11433 & ~n20375;
  assign n23181 = ~i_RtoB_ACK0 & ~n23180;
  assign n23182 = ~n23179 & ~n23181;
  assign n23183 = ~controllable_DEQ & ~n23182;
  assign n23184 = ~n23177 & ~n23183;
  assign n23185 = i_FULL & ~n23184;
  assign n23186 = ~n11395 & ~n17822;
  assign n23187 = i_RtoB_ACK0 & ~n23186;
  assign n23188 = ~n11447 & ~n20386;
  assign n23189 = ~i_RtoB_ACK0 & ~n23188;
  assign n23190 = ~n23187 & ~n23189;
  assign n23191 = controllable_DEQ & ~n23190;
  assign n23192 = ~n11424 & ~n17832;
  assign n23193 = i_RtoB_ACK0 & ~n23192;
  assign n23194 = ~n11456 & ~n20391;
  assign n23195 = ~i_RtoB_ACK0 & ~n23194;
  assign n23196 = ~n23193 & ~n23195;
  assign n23197 = ~controllable_DEQ & ~n23196;
  assign n23198 = ~n23191 & ~n23197;
  assign n23199 = ~i_FULL & ~n23198;
  assign n23200 = ~n23185 & ~n23199;
  assign n23201 = i_nEMPTY & ~n23200;
  assign n23202 = ~n11472 & ~n20404;
  assign n23203 = ~i_RtoB_ACK0 & ~n23202;
  assign n23204 = ~n15604 & ~n23203;
  assign n23205 = controllable_DEQ & ~n23204;
  assign n23206 = ~n11395 & ~n17850;
  assign n23207 = i_RtoB_ACK0 & ~n23206;
  assign n23208 = ~n11483 & ~n20409;
  assign n23209 = ~i_RtoB_ACK0 & ~n23208;
  assign n23210 = ~n23207 & ~n23209;
  assign n23211 = ~controllable_DEQ & ~n23210;
  assign n23212 = ~n23205 & ~n23211;
  assign n23213 = i_FULL & ~n23212;
  assign n23214 = ~n11493 & ~n20420;
  assign n23215 = ~i_RtoB_ACK0 & ~n23214;
  assign n23216 = ~n15619 & ~n23215;
  assign n23217 = controllable_DEQ & ~n23216;
  assign n23218 = ~controllable_DEQ & ~n23176;
  assign n23219 = ~n23217 & ~n23218;
  assign n23220 = ~i_FULL & ~n23219;
  assign n23221 = ~n23213 & ~n23220;
  assign n23222 = ~i_nEMPTY & ~n23221;
  assign n23223 = ~n23201 & ~n23222;
  assign n23224 = controllable_BtoS_ACK0 & ~n23223;
  assign n23225 = ~n11517 & ~n17874;
  assign n23226 = i_RtoB_ACK0 & ~n23225;
  assign n23227 = ~n11531 & ~n20432;
  assign n23228 = ~i_RtoB_ACK0 & ~n23227;
  assign n23229 = ~n23226 & ~n23228;
  assign n23230 = controllable_DEQ & ~n23229;
  assign n23231 = ~n11541 & ~n17886;
  assign n23232 = i_RtoB_ACK0 & ~n23231;
  assign n23233 = ~n11548 & ~n20437;
  assign n23234 = ~i_RtoB_ACK0 & ~n23233;
  assign n23235 = ~n23232 & ~n23234;
  assign n23236 = ~controllable_DEQ & ~n23235;
  assign n23237 = ~n23230 & ~n23236;
  assign n23238 = i_FULL & ~n23237;
  assign n23239 = ~n11517 & ~n17901;
  assign n23240 = i_RtoB_ACK0 & ~n23239;
  assign n23241 = ~n11562 & ~n20444;
  assign n23242 = ~i_RtoB_ACK0 & ~n23241;
  assign n23243 = ~n23240 & ~n23242;
  assign n23244 = controllable_DEQ & ~n23243;
  assign n23245 = ~n11541 & ~n17911;
  assign n23246 = i_RtoB_ACK0 & ~n23245;
  assign n23247 = ~n11571 & ~n20449;
  assign n23248 = ~i_RtoB_ACK0 & ~n23247;
  assign n23249 = ~n23246 & ~n23248;
  assign n23250 = ~controllable_DEQ & ~n23249;
  assign n23251 = ~n23244 & ~n23250;
  assign n23252 = ~i_FULL & ~n23251;
  assign n23253 = ~n23238 & ~n23252;
  assign n23254 = i_nEMPTY & ~n23253;
  assign n23255 = ~n11588 & ~n20458;
  assign n23256 = ~i_RtoB_ACK0 & ~n23255;
  assign n23257 = ~n17925 & ~n23256;
  assign n23258 = controllable_DEQ & ~n23257;
  assign n23259 = ~n11517 & ~n17933;
  assign n23260 = i_RtoB_ACK0 & ~n23259;
  assign n23261 = ~n11596 & ~n20463;
  assign n23262 = ~i_RtoB_ACK0 & ~n23261;
  assign n23263 = ~n23260 & ~n23262;
  assign n23264 = ~controllable_DEQ & ~n23263;
  assign n23265 = ~n23258 & ~n23264;
  assign n23266 = i_FULL & ~n23265;
  assign n23267 = ~n11606 & ~n20470;
  assign n23268 = ~i_RtoB_ACK0 & ~n23267;
  assign n23269 = ~n17943 & ~n23268;
  assign n23270 = controllable_DEQ & ~n23269;
  assign n23271 = ~controllable_DEQ & ~n23229;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = ~i_FULL & ~n23272;
  assign n23274 = ~n23266 & ~n23273;
  assign n23275 = ~i_nEMPTY & ~n23274;
  assign n23276 = ~n23254 & ~n23275;
  assign n23277 = ~controllable_BtoS_ACK0 & ~n23276;
  assign n23278 = ~n23224 & ~n23277;
  assign n23279 = n4465 & ~n23278;
  assign n23280 = ~n21416 & ~n23277;
  assign n23281 = ~n4465 & ~n23280;
  assign n23282 = ~n23279 & ~n23281;
  assign n23283 = i_StoB_REQ10 & ~n23282;
  assign n23284 = ~n11652 & ~n17965;
  assign n23285 = i_RtoB_ACK0 & ~n23284;
  assign n23286 = ~n11670 & ~n17974;
  assign n23287 = ~i_RtoB_ACK0 & ~n23286;
  assign n23288 = ~n23285 & ~n23287;
  assign n23289 = controllable_DEQ & ~n23288;
  assign n23290 = ~n11681 & ~n17984;
  assign n23291 = i_RtoB_ACK0 & ~n23290;
  assign n23292 = ~n11688 & ~n17993;
  assign n23293 = ~i_RtoB_ACK0 & ~n23292;
  assign n23294 = ~n23291 & ~n23293;
  assign n23295 = ~controllable_DEQ & ~n23294;
  assign n23296 = ~n23289 & ~n23295;
  assign n23297 = i_FULL & ~n23296;
  assign n23298 = ~n11652 & ~n18006;
  assign n23299 = i_RtoB_ACK0 & ~n23298;
  assign n23300 = ~n11705 & ~n18012;
  assign n23301 = ~i_RtoB_ACK0 & ~n23300;
  assign n23302 = ~n23299 & ~n23301;
  assign n23303 = controllable_DEQ & ~n23302;
  assign n23304 = ~n11681 & ~n18022;
  assign n23305 = i_RtoB_ACK0 & ~n23304;
  assign n23306 = ~n11714 & ~n18028;
  assign n23307 = ~i_RtoB_ACK0 & ~n23306;
  assign n23308 = ~n23305 & ~n23307;
  assign n23309 = ~controllable_DEQ & ~n23308;
  assign n23310 = ~n23303 & ~n23309;
  assign n23311 = ~i_FULL & ~n23310;
  assign n23312 = ~n23297 & ~n23311;
  assign n23313 = i_nEMPTY & ~n23312;
  assign n23314 = ~n11734 & ~n18049;
  assign n23315 = ~i_RtoB_ACK0 & ~n23314;
  assign n23316 = ~n18045 & ~n23315;
  assign n23317 = controllable_DEQ & ~n23316;
  assign n23318 = ~n11652 & ~n18059;
  assign n23319 = i_RtoB_ACK0 & ~n23318;
  assign n23320 = ~n11742 & ~n18065;
  assign n23321 = ~i_RtoB_ACK0 & ~n23320;
  assign n23322 = ~n23319 & ~n23321;
  assign n23323 = ~controllable_DEQ & ~n23322;
  assign n23324 = ~n23317 & ~n23323;
  assign n23325 = i_FULL & ~n23324;
  assign n23326 = ~n11752 & ~n18084;
  assign n23327 = ~i_RtoB_ACK0 & ~n23326;
  assign n23328 = ~n18080 & ~n23327;
  assign n23329 = controllable_DEQ & ~n23328;
  assign n23330 = ~n11760 & ~n17974;
  assign n23331 = ~i_RtoB_ACK0 & ~n23330;
  assign n23332 = ~n23285 & ~n23331;
  assign n23333 = ~controllable_DEQ & ~n23332;
  assign n23334 = ~n23329 & ~n23333;
  assign n23335 = ~i_FULL & ~n23334;
  assign n23336 = ~n23325 & ~n23335;
  assign n23337 = ~i_nEMPTY & ~n23336;
  assign n23338 = ~n23313 & ~n23337;
  assign n23339 = controllable_BtoS_ACK0 & ~n23338;
  assign n23340 = ~n11799 & ~n18107;
  assign n23341 = i_RtoB_ACK0 & ~n23340;
  assign n23342 = ~n11817 & ~n18116;
  assign n23343 = ~i_RtoB_ACK0 & ~n23342;
  assign n23344 = ~n23341 & ~n23343;
  assign n23345 = controllable_DEQ & ~n23344;
  assign n23346 = ~n11828 & ~n18126;
  assign n23347 = i_RtoB_ACK0 & ~n23346;
  assign n23348 = ~n11835 & ~n18135;
  assign n23349 = ~i_RtoB_ACK0 & ~n23348;
  assign n23350 = ~n23347 & ~n23349;
  assign n23351 = ~controllable_DEQ & ~n23350;
  assign n23352 = ~n23345 & ~n23351;
  assign n23353 = i_FULL & ~n23352;
  assign n23354 = ~n11799 & ~n18148;
  assign n23355 = i_RtoB_ACK0 & ~n23354;
  assign n23356 = ~n11852 & ~n18154;
  assign n23357 = ~i_RtoB_ACK0 & ~n23356;
  assign n23358 = ~n23355 & ~n23357;
  assign n23359 = controllable_DEQ & ~n23358;
  assign n23360 = ~n11828 & ~n18164;
  assign n23361 = i_RtoB_ACK0 & ~n23360;
  assign n23362 = ~n11861 & ~n18170;
  assign n23363 = ~i_RtoB_ACK0 & ~n23362;
  assign n23364 = ~n23361 & ~n23363;
  assign n23365 = ~controllable_DEQ & ~n23364;
  assign n23366 = ~n23359 & ~n23365;
  assign n23367 = ~i_FULL & ~n23366;
  assign n23368 = ~n23353 & ~n23367;
  assign n23369 = i_nEMPTY & ~n23368;
  assign n23370 = ~n11881 & ~n18191;
  assign n23371 = ~i_RtoB_ACK0 & ~n23370;
  assign n23372 = ~n18187 & ~n23371;
  assign n23373 = controllable_DEQ & ~n23372;
  assign n23374 = ~n11799 & ~n18201;
  assign n23375 = i_RtoB_ACK0 & ~n23374;
  assign n23376 = ~n11889 & ~n18207;
  assign n23377 = ~i_RtoB_ACK0 & ~n23376;
  assign n23378 = ~n23375 & ~n23377;
  assign n23379 = ~controllable_DEQ & ~n23378;
  assign n23380 = ~n23373 & ~n23379;
  assign n23381 = i_FULL & ~n23380;
  assign n23382 = ~n11899 & ~n18226;
  assign n23383 = ~i_RtoB_ACK0 & ~n23382;
  assign n23384 = ~n18222 & ~n23383;
  assign n23385 = controllable_DEQ & ~n23384;
  assign n23386 = ~n11907 & ~n18116;
  assign n23387 = ~i_RtoB_ACK0 & ~n23386;
  assign n23388 = ~n23341 & ~n23387;
  assign n23389 = ~controllable_DEQ & ~n23388;
  assign n23390 = ~n23385 & ~n23389;
  assign n23391 = ~i_FULL & ~n23390;
  assign n23392 = ~n23381 & ~n23391;
  assign n23393 = ~i_nEMPTY & ~n23392;
  assign n23394 = ~n23369 & ~n23393;
  assign n23395 = ~controllable_BtoS_ACK0 & ~n23394;
  assign n23396 = ~n23339 & ~n23395;
  assign n23397 = n4465 & ~n23396;
  assign n23398 = ~n21267 & ~n23397;
  assign n23399 = ~i_StoB_REQ10 & ~n23398;
  assign n23400 = ~n23283 & ~n23399;
  assign n23401 = ~controllable_BtoS_ACK10 & ~n23400;
  assign n23402 = ~n23171 & ~n23401;
  assign n23403 = n4464 & ~n23402;
  assign n23404 = ~n21559 & ~n23169;
  assign n23405 = controllable_BtoS_ACK10 & ~n23404;
  assign n23406 = ~n11936 & ~n18259;
  assign n23407 = i_RtoB_ACK0 & ~n23406;
  assign n23408 = ~n11950 & ~n20680;
  assign n23409 = ~i_RtoB_ACK0 & ~n23408;
  assign n23410 = ~n23407 & ~n23409;
  assign n23411 = controllable_DEQ & ~n23410;
  assign n23412 = ~n11960 & ~n18271;
  assign n23413 = i_RtoB_ACK0 & ~n23412;
  assign n23414 = ~n11967 & ~n20685;
  assign n23415 = ~i_RtoB_ACK0 & ~n23414;
  assign n23416 = ~n23413 & ~n23415;
  assign n23417 = ~controllable_DEQ & ~n23416;
  assign n23418 = ~n23411 & ~n23417;
  assign n23419 = i_FULL & ~n23418;
  assign n23420 = ~n11936 & ~n18286;
  assign n23421 = i_RtoB_ACK0 & ~n23420;
  assign n23422 = ~n11981 & ~n20692;
  assign n23423 = ~i_RtoB_ACK0 & ~n23422;
  assign n23424 = ~n23421 & ~n23423;
  assign n23425 = controllable_DEQ & ~n23424;
  assign n23426 = ~n11960 & ~n18296;
  assign n23427 = i_RtoB_ACK0 & ~n23426;
  assign n23428 = ~n11990 & ~n20697;
  assign n23429 = ~i_RtoB_ACK0 & ~n23428;
  assign n23430 = ~n23427 & ~n23429;
  assign n23431 = ~controllable_DEQ & ~n23430;
  assign n23432 = ~n23425 & ~n23431;
  assign n23433 = ~i_FULL & ~n23432;
  assign n23434 = ~n23419 & ~n23433;
  assign n23435 = i_nEMPTY & ~n23434;
  assign n23436 = ~n12006 & ~n20706;
  assign n23437 = ~i_RtoB_ACK0 & ~n23436;
  assign n23438 = ~n15604 & ~n23437;
  assign n23439 = controllable_DEQ & ~n23438;
  assign n23440 = ~n11936 & ~n18314;
  assign n23441 = i_RtoB_ACK0 & ~n23440;
  assign n23442 = ~n12014 & ~n20711;
  assign n23443 = ~i_RtoB_ACK0 & ~n23442;
  assign n23444 = ~n23441 & ~n23443;
  assign n23445 = ~controllable_DEQ & ~n23444;
  assign n23446 = ~n23439 & ~n23445;
  assign n23447 = i_FULL & ~n23446;
  assign n23448 = ~n12024 & ~n20718;
  assign n23449 = ~i_RtoB_ACK0 & ~n23448;
  assign n23450 = ~n15619 & ~n23449;
  assign n23451 = controllable_DEQ & ~n23450;
  assign n23452 = ~controllable_DEQ & ~n23410;
  assign n23453 = ~n23451 & ~n23452;
  assign n23454 = ~i_FULL & ~n23453;
  assign n23455 = ~n23447 & ~n23454;
  assign n23456 = ~i_nEMPTY & ~n23455;
  assign n23457 = ~n23435 & ~n23456;
  assign n23458 = controllable_BtoS_ACK0 & ~n23457;
  assign n23459 = ~n12044 & ~n18338;
  assign n23460 = i_RtoB_ACK0 & ~n23459;
  assign n23461 = ~n12058 & ~n20730;
  assign n23462 = ~i_RtoB_ACK0 & ~n23461;
  assign n23463 = ~n23460 & ~n23462;
  assign n23464 = controllable_DEQ & ~n23463;
  assign n23465 = ~n12068 & ~n18350;
  assign n23466 = i_RtoB_ACK0 & ~n23465;
  assign n23467 = ~n12075 & ~n20735;
  assign n23468 = ~i_RtoB_ACK0 & ~n23467;
  assign n23469 = ~n23466 & ~n23468;
  assign n23470 = ~controllable_DEQ & ~n23469;
  assign n23471 = ~n23464 & ~n23470;
  assign n23472 = i_FULL & ~n23471;
  assign n23473 = ~n12044 & ~n18365;
  assign n23474 = i_RtoB_ACK0 & ~n23473;
  assign n23475 = ~n12089 & ~n20742;
  assign n23476 = ~i_RtoB_ACK0 & ~n23475;
  assign n23477 = ~n23474 & ~n23476;
  assign n23478 = controllable_DEQ & ~n23477;
  assign n23479 = ~n12068 & ~n18375;
  assign n23480 = i_RtoB_ACK0 & ~n23479;
  assign n23481 = ~n12098 & ~n20747;
  assign n23482 = ~i_RtoB_ACK0 & ~n23481;
  assign n23483 = ~n23480 & ~n23482;
  assign n23484 = ~controllable_DEQ & ~n23483;
  assign n23485 = ~n23478 & ~n23484;
  assign n23486 = ~i_FULL & ~n23485;
  assign n23487 = ~n23472 & ~n23486;
  assign n23488 = i_nEMPTY & ~n23487;
  assign n23489 = ~n12114 & ~n20756;
  assign n23490 = ~i_RtoB_ACK0 & ~n23489;
  assign n23491 = ~n17925 & ~n23490;
  assign n23492 = controllable_DEQ & ~n23491;
  assign n23493 = ~n12044 & ~n18393;
  assign n23494 = i_RtoB_ACK0 & ~n23493;
  assign n23495 = ~n12122 & ~n20761;
  assign n23496 = ~i_RtoB_ACK0 & ~n23495;
  assign n23497 = ~n23494 & ~n23496;
  assign n23498 = ~controllable_DEQ & ~n23497;
  assign n23499 = ~n23492 & ~n23498;
  assign n23500 = i_FULL & ~n23499;
  assign n23501 = ~n12132 & ~n20768;
  assign n23502 = ~i_RtoB_ACK0 & ~n23501;
  assign n23503 = ~n17943 & ~n23502;
  assign n23504 = controllable_DEQ & ~n23503;
  assign n23505 = ~controllable_DEQ & ~n23463;
  assign n23506 = ~n23504 & ~n23505;
  assign n23507 = ~i_FULL & ~n23506;
  assign n23508 = ~n23500 & ~n23507;
  assign n23509 = ~i_nEMPTY & ~n23508;
  assign n23510 = ~n23488 & ~n23509;
  assign n23511 = ~controllable_BtoS_ACK0 & ~n23510;
  assign n23512 = ~n23458 & ~n23511;
  assign n23513 = n4465 & ~n23512;
  assign n23514 = ~n21920 & ~n23511;
  assign n23515 = ~n4465 & ~n23514;
  assign n23516 = ~n23513 & ~n23515;
  assign n23517 = i_StoB_REQ10 & ~n23516;
  assign n23518 = ~n21773 & ~n23517;
  assign n23519 = ~controllable_BtoS_ACK10 & ~n23518;
  assign n23520 = ~n23405 & ~n23519;
  assign n23521 = ~n4464 & ~n23520;
  assign n23522 = ~n23403 & ~n23521;
  assign n23523 = n4463 & ~n23522;
  assign n23524 = ~n12168 & ~n18428;
  assign n23525 = i_RtoB_ACK0 & ~n23524;
  assign n23526 = ~n12179 & ~n17545;
  assign n23527 = ~i_RtoB_ACK0 & ~n23526;
  assign n23528 = ~n23525 & ~n23527;
  assign n23529 = controllable_DEQ & ~n23528;
  assign n23530 = ~n12189 & ~n18434;
  assign n23531 = i_RtoB_ACK0 & ~n23530;
  assign n23532 = ~n12197 & ~n17562;
  assign n23533 = ~i_RtoB_ACK0 & ~n23532;
  assign n23534 = ~n23531 & ~n23533;
  assign n23535 = ~controllable_DEQ & ~n23534;
  assign n23536 = ~n23529 & ~n23535;
  assign n23537 = i_nEMPTY & ~n23536;
  assign n23538 = ~n12209 & ~n17571;
  assign n23539 = ~i_RtoB_ACK0 & ~n23538;
  assign n23540 = ~i_RtoB_ACK0 & ~n23539;
  assign n23541 = controllable_DEQ & ~n23540;
  assign n23542 = ~n12220 & ~n17581;
  assign n23543 = ~i_RtoB_ACK0 & ~n23542;
  assign n23544 = ~n23525 & ~n23543;
  assign n23545 = ~controllable_DEQ & ~n23544;
  assign n23546 = ~n23541 & ~n23545;
  assign n23547 = i_FULL & ~n23546;
  assign n23548 = ~n12230 & ~n17590;
  assign n23549 = ~i_RtoB_ACK0 & ~n23548;
  assign n23550 = ~i_RtoB_ACK0 & ~n23549;
  assign n23551 = controllable_DEQ & ~n23550;
  assign n23552 = ~n12238 & ~n17545;
  assign n23553 = ~i_RtoB_ACK0 & ~n23552;
  assign n23554 = ~n23525 & ~n23553;
  assign n23555 = ~controllable_DEQ & ~n23554;
  assign n23556 = ~n23551 & ~n23555;
  assign n23557 = ~i_FULL & ~n23556;
  assign n23558 = ~n23547 & ~n23557;
  assign n23559 = ~i_nEMPTY & ~n23558;
  assign n23560 = ~n23537 & ~n23559;
  assign n23561 = controllable_BtoS_ACK0 & ~n23560;
  assign n23562 = ~n12261 & ~n18456;
  assign n23563 = i_RtoB_ACK0 & ~n23562;
  assign n23564 = ~n12270 & ~n14824;
  assign n23565 = ~i_RtoB_ACK0 & ~n23564;
  assign n23566 = ~n23563 & ~n23565;
  assign n23567 = controllable_DEQ & ~n23566;
  assign n23568 = ~n12279 & ~n18462;
  assign n23569 = i_RtoB_ACK0 & ~n23568;
  assign n23570 = ~n12283 & ~n14841;
  assign n23571 = ~i_RtoB_ACK0 & ~n23570;
  assign n23572 = ~n23569 & ~n23571;
  assign n23573 = ~controllable_DEQ & ~n23572;
  assign n23574 = ~n23567 & ~n23573;
  assign n23575 = i_nEMPTY & ~n23574;
  assign n23576 = ~n12295 & ~n14850;
  assign n23577 = ~i_RtoB_ACK0 & ~n23576;
  assign n23578 = ~i_RtoB_ACK0 & ~n23577;
  assign n23579 = controllable_DEQ & ~n23578;
  assign n23580 = ~n12301 & ~n14860;
  assign n23581 = ~i_RtoB_ACK0 & ~n23580;
  assign n23582 = ~n23563 & ~n23581;
  assign n23583 = ~controllable_DEQ & ~n23582;
  assign n23584 = ~n23579 & ~n23583;
  assign n23585 = i_FULL & ~n23584;
  assign n23586 = ~n12311 & ~n14869;
  assign n23587 = ~i_RtoB_ACK0 & ~n23586;
  assign n23588 = ~i_RtoB_ACK0 & ~n23587;
  assign n23589 = controllable_DEQ & ~n23588;
  assign n23590 = ~n12321 & ~n14824;
  assign n23591 = ~i_RtoB_ACK0 & ~n23590;
  assign n23592 = ~n23563 & ~n23591;
  assign n23593 = ~controllable_DEQ & ~n23592;
  assign n23594 = ~n23589 & ~n23593;
  assign n23595 = ~i_FULL & ~n23594;
  assign n23596 = ~n23585 & ~n23595;
  assign n23597 = ~i_nEMPTY & ~n23596;
  assign n23598 = ~n23575 & ~n23597;
  assign n23599 = ~controllable_BtoS_ACK0 & ~n23598;
  assign n23600 = ~n23561 & ~n23599;
  assign n23601 = n4465 & ~n23600;
  assign n23602 = ~n22093 & ~n23571;
  assign n23603 = ~controllable_DEQ & ~n23602;
  assign n23604 = ~n22103 & ~n23603;
  assign n23605 = i_nEMPTY & ~n23604;
  assign n23606 = ~n22087 & ~n23581;
  assign n23607 = ~controllable_DEQ & ~n23606;
  assign n23608 = ~n22115 & ~n23607;
  assign n23609 = i_FULL & ~n23608;
  assign n23610 = ~n22087 & ~n23591;
  assign n23611 = ~controllable_DEQ & ~n23610;
  assign n23612 = ~n22125 & ~n23611;
  assign n23613 = ~i_FULL & ~n23612;
  assign n23614 = ~n23609 & ~n23613;
  assign n23615 = ~i_nEMPTY & ~n23614;
  assign n23616 = ~n23605 & ~n23615;
  assign n23617 = ~controllable_BtoS_ACK0 & ~n23616;
  assign n23618 = ~n21013 & ~n23617;
  assign n23619 = ~n4465 & ~n23618;
  assign n23620 = ~n23601 & ~n23619;
  assign n23621 = i_StoB_REQ10 & ~n23620;
  assign n23622 = ~n23169 & ~n23621;
  assign n23623 = controllable_BtoS_ACK10 & ~n23622;
  assign n23624 = ~n12359 & ~n17050;
  assign n23625 = i_RtoB_ACK0 & ~n23624;
  assign n23626 = ~n12374 & ~n20366;
  assign n23627 = ~i_RtoB_ACK0 & ~n23626;
  assign n23628 = ~n23625 & ~n23627;
  assign n23629 = controllable_DEQ & ~n23628;
  assign n23630 = ~n12382 & ~n17058;
  assign n23631 = i_RtoB_ACK0 & ~n23630;
  assign n23632 = ~n12391 & ~n20375;
  assign n23633 = ~i_RtoB_ACK0 & ~n23632;
  assign n23634 = ~n23631 & ~n23633;
  assign n23635 = ~controllable_DEQ & ~n23634;
  assign n23636 = ~n23629 & ~n23635;
  assign n23637 = i_FULL & ~n23636;
  assign n23638 = ~n12403 & ~n20386;
  assign n23639 = ~i_RtoB_ACK0 & ~n23638;
  assign n23640 = ~n23625 & ~n23639;
  assign n23641 = controllable_DEQ & ~n23640;
  assign n23642 = ~n12413 & ~n20391;
  assign n23643 = ~i_RtoB_ACK0 & ~n23642;
  assign n23644 = ~n23631 & ~n23643;
  assign n23645 = ~controllable_DEQ & ~n23644;
  assign n23646 = ~n23641 & ~n23645;
  assign n23647 = ~i_FULL & ~n23646;
  assign n23648 = ~n23637 & ~n23647;
  assign n23649 = i_nEMPTY & ~n23648;
  assign n23650 = ~n12423 & ~n20404;
  assign n23651 = ~i_RtoB_ACK0 & ~n23650;
  assign n23652 = ~n15604 & ~n23651;
  assign n23653 = controllable_DEQ & ~n23652;
  assign n23654 = ~n12359 & ~n17068;
  assign n23655 = i_RtoB_ACK0 & ~n23654;
  assign n23656 = ~n12435 & ~n20409;
  assign n23657 = ~i_RtoB_ACK0 & ~n23656;
  assign n23658 = ~n23655 & ~n23657;
  assign n23659 = ~controllable_DEQ & ~n23658;
  assign n23660 = ~n23653 & ~n23659;
  assign n23661 = i_FULL & ~n23660;
  assign n23662 = ~n12443 & ~n20420;
  assign n23663 = ~i_RtoB_ACK0 & ~n23662;
  assign n23664 = ~n15619 & ~n23663;
  assign n23665 = controllable_DEQ & ~n23664;
  assign n23666 = ~controllable_DEQ & ~n23628;
  assign n23667 = ~n23665 & ~n23666;
  assign n23668 = ~i_FULL & ~n23667;
  assign n23669 = ~n23661 & ~n23668;
  assign n23670 = ~i_nEMPTY & ~n23669;
  assign n23671 = ~n23649 & ~n23670;
  assign n23672 = controllable_BtoS_ACK0 & ~n23671;
  assign n23673 = ~n12458 & ~n18522;
  assign n23674 = i_RtoB_ACK0 & ~n23673;
  assign n23675 = ~n12468 & ~n20432;
  assign n23676 = ~i_RtoB_ACK0 & ~n23675;
  assign n23677 = ~n23674 & ~n23676;
  assign n23678 = controllable_DEQ & ~n23677;
  assign n23679 = ~n12476 & ~n18530;
  assign n23680 = i_RtoB_ACK0 & ~n23679;
  assign n23681 = ~n12482 & ~n20437;
  assign n23682 = ~i_RtoB_ACK0 & ~n23681;
  assign n23683 = ~n23680 & ~n23682;
  assign n23684 = ~controllable_DEQ & ~n23683;
  assign n23685 = ~n23678 & ~n23684;
  assign n23686 = i_FULL & ~n23685;
  assign n23687 = ~n12494 & ~n20444;
  assign n23688 = ~i_RtoB_ACK0 & ~n23687;
  assign n23689 = ~n23674 & ~n23688;
  assign n23690 = controllable_DEQ & ~n23689;
  assign n23691 = ~n12504 & ~n20449;
  assign n23692 = ~i_RtoB_ACK0 & ~n23691;
  assign n23693 = ~n23680 & ~n23692;
  assign n23694 = ~controllable_DEQ & ~n23693;
  assign n23695 = ~n23690 & ~n23694;
  assign n23696 = ~i_FULL & ~n23695;
  assign n23697 = ~n23686 & ~n23696;
  assign n23698 = i_nEMPTY & ~n23697;
  assign n23699 = ~n12514 & ~n20458;
  assign n23700 = ~i_RtoB_ACK0 & ~n23699;
  assign n23701 = ~n17925 & ~n23700;
  assign n23702 = controllable_DEQ & ~n23701;
  assign n23703 = ~n12458 & ~n18548;
  assign n23704 = i_RtoB_ACK0 & ~n23703;
  assign n23705 = ~n12522 & ~n20463;
  assign n23706 = ~i_RtoB_ACK0 & ~n23705;
  assign n23707 = ~n23704 & ~n23706;
  assign n23708 = ~controllable_DEQ & ~n23707;
  assign n23709 = ~n23702 & ~n23708;
  assign n23710 = i_FULL & ~n23709;
  assign n23711 = ~n12530 & ~n20470;
  assign n23712 = ~i_RtoB_ACK0 & ~n23711;
  assign n23713 = ~n17943 & ~n23712;
  assign n23714 = controllable_DEQ & ~n23713;
  assign n23715 = ~controllable_DEQ & ~n23677;
  assign n23716 = ~n23714 & ~n23715;
  assign n23717 = ~i_FULL & ~n23716;
  assign n23718 = ~n23710 & ~n23717;
  assign n23719 = ~i_nEMPTY & ~n23718;
  assign n23720 = ~n23698 & ~n23719;
  assign n23721 = ~controllable_BtoS_ACK0 & ~n23720;
  assign n23722 = ~n23672 & ~n23721;
  assign n23723 = n4465 & ~n23722;
  assign n23724 = ~n22480 & ~n23721;
  assign n23725 = ~n4465 & ~n23724;
  assign n23726 = ~n23723 & ~n23725;
  assign n23727 = i_StoB_REQ10 & ~n23726;
  assign n23728 = ~n12551 & ~n18572;
  assign n23729 = i_RtoB_ACK0 & ~n23728;
  assign n23730 = ~n12561 & ~n17974;
  assign n23731 = ~i_RtoB_ACK0 & ~n23730;
  assign n23732 = ~n23729 & ~n23731;
  assign n23733 = controllable_DEQ & ~n23732;
  assign n23734 = ~n12569 & ~n18580;
  assign n23735 = i_RtoB_ACK0 & ~n23734;
  assign n23736 = ~n12575 & ~n17993;
  assign n23737 = ~i_RtoB_ACK0 & ~n23736;
  assign n23738 = ~n23735 & ~n23737;
  assign n23739 = ~controllable_DEQ & ~n23738;
  assign n23740 = ~n23733 & ~n23739;
  assign n23741 = i_FULL & ~n23740;
  assign n23742 = ~n12587 & ~n18012;
  assign n23743 = ~i_RtoB_ACK0 & ~n23742;
  assign n23744 = ~n23729 & ~n23743;
  assign n23745 = controllable_DEQ & ~n23744;
  assign n23746 = ~n12597 & ~n18028;
  assign n23747 = ~i_RtoB_ACK0 & ~n23746;
  assign n23748 = ~n23735 & ~n23747;
  assign n23749 = ~controllable_DEQ & ~n23748;
  assign n23750 = ~n23745 & ~n23749;
  assign n23751 = ~i_FULL & ~n23750;
  assign n23752 = ~n23741 & ~n23751;
  assign n23753 = i_nEMPTY & ~n23752;
  assign n23754 = ~n12607 & ~n18049;
  assign n23755 = ~i_RtoB_ACK0 & ~n23754;
  assign n23756 = ~n18045 & ~n23755;
  assign n23757 = controllable_DEQ & ~n23756;
  assign n23758 = ~n12551 & ~n18598;
  assign n23759 = i_RtoB_ACK0 & ~n23758;
  assign n23760 = ~n12615 & ~n18065;
  assign n23761 = ~i_RtoB_ACK0 & ~n23760;
  assign n23762 = ~n23759 & ~n23761;
  assign n23763 = ~controllable_DEQ & ~n23762;
  assign n23764 = ~n23757 & ~n23763;
  assign n23765 = i_FULL & ~n23764;
  assign n23766 = ~n12623 & ~n18084;
  assign n23767 = ~i_RtoB_ACK0 & ~n23766;
  assign n23768 = ~n18080 & ~n23767;
  assign n23769 = controllable_DEQ & ~n23768;
  assign n23770 = ~n12633 & ~n17974;
  assign n23771 = ~i_RtoB_ACK0 & ~n23770;
  assign n23772 = ~n23729 & ~n23771;
  assign n23773 = ~controllable_DEQ & ~n23772;
  assign n23774 = ~n23769 & ~n23773;
  assign n23775 = ~i_FULL & ~n23774;
  assign n23776 = ~n23765 & ~n23775;
  assign n23777 = ~i_nEMPTY & ~n23776;
  assign n23778 = ~n23753 & ~n23777;
  assign n23779 = controllable_BtoS_ACK0 & ~n23778;
  assign n23780 = ~n12647 & ~n18617;
  assign n23781 = i_RtoB_ACK0 & ~n23780;
  assign n23782 = ~n12657 & ~n18116;
  assign n23783 = ~i_RtoB_ACK0 & ~n23782;
  assign n23784 = ~n23781 & ~n23783;
  assign n23785 = controllable_DEQ & ~n23784;
  assign n23786 = ~n12665 & ~n18625;
  assign n23787 = i_RtoB_ACK0 & ~n23786;
  assign n23788 = ~n12671 & ~n18135;
  assign n23789 = ~i_RtoB_ACK0 & ~n23788;
  assign n23790 = ~n23787 & ~n23789;
  assign n23791 = ~controllable_DEQ & ~n23790;
  assign n23792 = ~n23785 & ~n23791;
  assign n23793 = i_FULL & ~n23792;
  assign n23794 = ~n12683 & ~n18154;
  assign n23795 = ~i_RtoB_ACK0 & ~n23794;
  assign n23796 = ~n23781 & ~n23795;
  assign n23797 = controllable_DEQ & ~n23796;
  assign n23798 = ~n12693 & ~n18170;
  assign n23799 = ~i_RtoB_ACK0 & ~n23798;
  assign n23800 = ~n23787 & ~n23799;
  assign n23801 = ~controllable_DEQ & ~n23800;
  assign n23802 = ~n23797 & ~n23801;
  assign n23803 = ~i_FULL & ~n23802;
  assign n23804 = ~n23793 & ~n23803;
  assign n23805 = i_nEMPTY & ~n23804;
  assign n23806 = ~n12703 & ~n18191;
  assign n23807 = ~i_RtoB_ACK0 & ~n23806;
  assign n23808 = ~n18187 & ~n23807;
  assign n23809 = controllable_DEQ & ~n23808;
  assign n23810 = ~n12647 & ~n18643;
  assign n23811 = i_RtoB_ACK0 & ~n23810;
  assign n23812 = ~n12711 & ~n18207;
  assign n23813 = ~i_RtoB_ACK0 & ~n23812;
  assign n23814 = ~n23811 & ~n23813;
  assign n23815 = ~controllable_DEQ & ~n23814;
  assign n23816 = ~n23809 & ~n23815;
  assign n23817 = i_FULL & ~n23816;
  assign n23818 = ~n12719 & ~n18226;
  assign n23819 = ~i_RtoB_ACK0 & ~n23818;
  assign n23820 = ~n18222 & ~n23819;
  assign n23821 = controllable_DEQ & ~n23820;
  assign n23822 = ~n12727 & ~n18116;
  assign n23823 = ~i_RtoB_ACK0 & ~n23822;
  assign n23824 = ~n23781 & ~n23823;
  assign n23825 = ~controllable_DEQ & ~n23824;
  assign n23826 = ~n23821 & ~n23825;
  assign n23827 = ~i_FULL & ~n23826;
  assign n23828 = ~n23817 & ~n23827;
  assign n23829 = ~i_nEMPTY & ~n23828;
  assign n23830 = ~n23805 & ~n23829;
  assign n23831 = ~controllable_BtoS_ACK0 & ~n23830;
  assign n23832 = ~n23779 & ~n23831;
  assign n23833 = n4465 & ~n23832;
  assign n23834 = ~n12741 & ~n17280;
  assign n23835 = i_RtoB_ACK0 & ~n23834;
  assign n23836 = ~n12745 & ~n15190;
  assign n23837 = ~i_RtoB_ACK0 & ~n23836;
  assign n23838 = ~n23835 & ~n23837;
  assign n23839 = controllable_DEQ & ~n23838;
  assign n23840 = ~n12751 & ~n17288;
  assign n23841 = i_RtoB_ACK0 & ~n23840;
  assign n23842 = ~n22255 & ~n23841;
  assign n23843 = ~controllable_DEQ & ~n23842;
  assign n23844 = ~n23839 & ~n23843;
  assign n23845 = i_nEMPTY & ~n23844;
  assign n23846 = ~n12759 & ~n15221;
  assign n23847 = ~i_RtoB_ACK0 & ~n23846;
  assign n23848 = ~n15217 & ~n23847;
  assign n23849 = controllable_DEQ & ~n23848;
  assign n23850 = ~n12741 & ~n17298;
  assign n23851 = i_RtoB_ACK0 & ~n23850;
  assign n23852 = ~n22267 & ~n23851;
  assign n23853 = ~controllable_DEQ & ~n23852;
  assign n23854 = ~n23849 & ~n23853;
  assign n23855 = i_FULL & ~n23854;
  assign n23856 = ~n12769 & ~n15249;
  assign n23857 = ~i_RtoB_ACK0 & ~n23856;
  assign n23858 = ~n15245 & ~n23857;
  assign n23859 = controllable_DEQ & ~n23858;
  assign n23860 = ~n22277 & ~n23835;
  assign n23861 = ~controllable_DEQ & ~n23860;
  assign n23862 = ~n23859 & ~n23861;
  assign n23863 = ~i_FULL & ~n23862;
  assign n23864 = ~n23855 & ~n23863;
  assign n23865 = ~i_nEMPTY & ~n23864;
  assign n23866 = ~n23845 & ~n23865;
  assign n23867 = controllable_BtoS_ACK0 & ~n23866;
  assign n23868 = ~n22337 & ~n23867;
  assign n23869 = ~n4465 & ~n23868;
  assign n23870 = ~n23833 & ~n23869;
  assign n23871 = ~i_StoB_REQ10 & ~n23870;
  assign n23872 = ~n23727 & ~n23871;
  assign n23873 = ~controllable_BtoS_ACK10 & ~n23872;
  assign n23874 = ~n23623 & ~n23873;
  assign n23875 = n4464 & ~n23874;
  assign n23876 = ~n12791 & ~n15749;
  assign n23877 = ~i_RtoB_ACK0 & ~n23876;
  assign n23878 = ~n22545 & ~n23877;
  assign n23879 = ~controllable_DEQ & ~n23878;
  assign n23880 = ~n22555 & ~n23879;
  assign n23881 = i_nEMPTY & ~n23880;
  assign n23882 = ~n12799 & ~n15768;
  assign n23883 = ~i_RtoB_ACK0 & ~n23882;
  assign n23884 = ~n22539 & ~n23883;
  assign n23885 = ~controllable_DEQ & ~n23884;
  assign n23886 = ~n22567 & ~n23885;
  assign n23887 = i_FULL & ~n23886;
  assign n23888 = ~n12809 & ~n15732;
  assign n23889 = ~i_RtoB_ACK0 & ~n23888;
  assign n23890 = ~n22539 & ~n23889;
  assign n23891 = ~controllable_DEQ & ~n23890;
  assign n23892 = ~n22577 & ~n23891;
  assign n23893 = ~i_FULL & ~n23892;
  assign n23894 = ~n23887 & ~n23893;
  assign n23895 = ~i_nEMPTY & ~n23894;
  assign n23896 = ~n23881 & ~n23895;
  assign n23897 = controllable_BtoS_ACK0 & ~n23896;
  assign n23898 = ~n12821 & ~n15824;
  assign n23899 = ~i_RtoB_ACK0 & ~n23898;
  assign n23900 = ~n22595 & ~n23899;
  assign n23901 = ~controllable_DEQ & ~n23900;
  assign n23902 = ~n22605 & ~n23901;
  assign n23903 = i_nEMPTY & ~n23902;
  assign n23904 = ~n12829 & ~n15843;
  assign n23905 = ~i_RtoB_ACK0 & ~n23904;
  assign n23906 = ~n22589 & ~n23905;
  assign n23907 = ~controllable_DEQ & ~n23906;
  assign n23908 = ~n22617 & ~n23907;
  assign n23909 = i_FULL & ~n23908;
  assign n23910 = ~n12839 & ~n15807;
  assign n23911 = ~i_RtoB_ACK0 & ~n23910;
  assign n23912 = ~n22589 & ~n23911;
  assign n23913 = ~controllable_DEQ & ~n23912;
  assign n23914 = ~n22627 & ~n23913;
  assign n23915 = ~i_FULL & ~n23914;
  assign n23916 = ~n23909 & ~n23915;
  assign n23917 = ~i_nEMPTY & ~n23916;
  assign n23918 = ~n23903 & ~n23917;
  assign n23919 = ~controllable_BtoS_ACK0 & ~n23918;
  assign n23920 = ~n23897 & ~n23919;
  assign n23921 = n4465 & ~n23920;
  assign n23922 = ~n21013 & ~n23919;
  assign n23923 = ~n4465 & ~n23922;
  assign n23924 = ~n23921 & ~n23923;
  assign n23925 = i_StoB_REQ10 & ~n23924;
  assign n23926 = ~n23169 & ~n23925;
  assign n23927 = controllable_BtoS_ACK10 & ~n23926;
  assign n23928 = ~n12861 & ~n17050;
  assign n23929 = i_RtoB_ACK0 & ~n23928;
  assign n23930 = ~n12869 & ~n20680;
  assign n23931 = ~i_RtoB_ACK0 & ~n23930;
  assign n23932 = ~n23929 & ~n23931;
  assign n23933 = controllable_DEQ & ~n23932;
  assign n23934 = ~n12877 & ~n17058;
  assign n23935 = i_RtoB_ACK0 & ~n23934;
  assign n23936 = ~n12883 & ~n20685;
  assign n23937 = ~i_RtoB_ACK0 & ~n23936;
  assign n23938 = ~n23935 & ~n23937;
  assign n23939 = ~controllable_DEQ & ~n23938;
  assign n23940 = ~n23933 & ~n23939;
  assign n23941 = i_FULL & ~n23940;
  assign n23942 = ~n12895 & ~n20692;
  assign n23943 = ~i_RtoB_ACK0 & ~n23942;
  assign n23944 = ~n23929 & ~n23943;
  assign n23945 = controllable_DEQ & ~n23944;
  assign n23946 = ~n12905 & ~n20697;
  assign n23947 = ~i_RtoB_ACK0 & ~n23946;
  assign n23948 = ~n23935 & ~n23947;
  assign n23949 = ~controllable_DEQ & ~n23948;
  assign n23950 = ~n23945 & ~n23949;
  assign n23951 = ~i_FULL & ~n23950;
  assign n23952 = ~n23941 & ~n23951;
  assign n23953 = i_nEMPTY & ~n23952;
  assign n23954 = ~n12915 & ~n20706;
  assign n23955 = ~i_RtoB_ACK0 & ~n23954;
  assign n23956 = ~n15604 & ~n23955;
  assign n23957 = controllable_DEQ & ~n23956;
  assign n23958 = ~n12861 & ~n17068;
  assign n23959 = i_RtoB_ACK0 & ~n23958;
  assign n23960 = ~n12923 & ~n20711;
  assign n23961 = ~i_RtoB_ACK0 & ~n23960;
  assign n23962 = ~n23959 & ~n23961;
  assign n23963 = ~controllable_DEQ & ~n23962;
  assign n23964 = ~n23957 & ~n23963;
  assign n23965 = i_FULL & ~n23964;
  assign n23966 = ~n12931 & ~n20718;
  assign n23967 = ~i_RtoB_ACK0 & ~n23966;
  assign n23968 = ~n15619 & ~n23967;
  assign n23969 = controllable_DEQ & ~n23968;
  assign n23970 = ~controllable_DEQ & ~n23932;
  assign n23971 = ~n23969 & ~n23970;
  assign n23972 = ~i_FULL & ~n23971;
  assign n23973 = ~n23965 & ~n23972;
  assign n23974 = ~i_nEMPTY & ~n23973;
  assign n23975 = ~n23953 & ~n23974;
  assign n23976 = controllable_BtoS_ACK0 & ~n23975;
  assign n23977 = ~n12946 & ~n18522;
  assign n23978 = i_RtoB_ACK0 & ~n23977;
  assign n23979 = ~n12954 & ~n20730;
  assign n23980 = ~i_RtoB_ACK0 & ~n23979;
  assign n23981 = ~n23978 & ~n23980;
  assign n23982 = controllable_DEQ & ~n23981;
  assign n23983 = ~n12962 & ~n18530;
  assign n23984 = i_RtoB_ACK0 & ~n23983;
  assign n23985 = ~n12968 & ~n20735;
  assign n23986 = ~i_RtoB_ACK0 & ~n23985;
  assign n23987 = ~n23984 & ~n23986;
  assign n23988 = ~controllable_DEQ & ~n23987;
  assign n23989 = ~n23982 & ~n23988;
  assign n23990 = i_FULL & ~n23989;
  assign n23991 = ~n12980 & ~n20742;
  assign n23992 = ~i_RtoB_ACK0 & ~n23991;
  assign n23993 = ~n23978 & ~n23992;
  assign n23994 = controllable_DEQ & ~n23993;
  assign n23995 = ~n12990 & ~n20747;
  assign n23996 = ~i_RtoB_ACK0 & ~n23995;
  assign n23997 = ~n23984 & ~n23996;
  assign n23998 = ~controllable_DEQ & ~n23997;
  assign n23999 = ~n23994 & ~n23998;
  assign n24000 = ~i_FULL & ~n23999;
  assign n24001 = ~n23990 & ~n24000;
  assign n24002 = i_nEMPTY & ~n24001;
  assign n24003 = ~n13000 & ~n20756;
  assign n24004 = ~i_RtoB_ACK0 & ~n24003;
  assign n24005 = ~n17925 & ~n24004;
  assign n24006 = controllable_DEQ & ~n24005;
  assign n24007 = ~n12946 & ~n18548;
  assign n24008 = i_RtoB_ACK0 & ~n24007;
  assign n24009 = ~n13008 & ~n20761;
  assign n24010 = ~i_RtoB_ACK0 & ~n24009;
  assign n24011 = ~n24008 & ~n24010;
  assign n24012 = ~controllable_DEQ & ~n24011;
  assign n24013 = ~n24006 & ~n24012;
  assign n24014 = i_FULL & ~n24013;
  assign n24015 = ~n13016 & ~n20768;
  assign n24016 = ~i_RtoB_ACK0 & ~n24015;
  assign n24017 = ~n17943 & ~n24016;
  assign n24018 = controllable_DEQ & ~n24017;
  assign n24019 = ~controllable_DEQ & ~n23981;
  assign n24020 = ~n24018 & ~n24019;
  assign n24021 = ~i_FULL & ~n24020;
  assign n24022 = ~n24014 & ~n24021;
  assign n24023 = ~i_nEMPTY & ~n24022;
  assign n24024 = ~n24002 & ~n24023;
  assign n24025 = ~controllable_BtoS_ACK0 & ~n24024;
  assign n24026 = ~n23976 & ~n24025;
  assign n24027 = n4465 & ~n24026;
  assign n24028 = ~n22984 & ~n24025;
  assign n24029 = ~n4465 & ~n24028;
  assign n24030 = ~n24027 & ~n24029;
  assign n24031 = i_StoB_REQ10 & ~n24030;
  assign n24032 = ~n13035 & ~n18766;
  assign n24033 = i_RtoB_ACK0 & ~n24032;
  assign n24034 = ~n13039 & ~n15889;
  assign n24035 = ~i_RtoB_ACK0 & ~n24034;
  assign n24036 = ~n24033 & ~n24035;
  assign n24037 = controllable_DEQ & ~n24036;
  assign n24038 = ~n13045 & ~n18774;
  assign n24039 = i_RtoB_ACK0 & ~n24038;
  assign n24040 = ~n22653 & ~n24039;
  assign n24041 = ~controllable_DEQ & ~n24040;
  assign n24042 = ~n24037 & ~n24041;
  assign n24043 = i_FULL & ~n24042;
  assign n24044 = ~n13053 & ~n15927;
  assign n24045 = ~i_RtoB_ACK0 & ~n24044;
  assign n24046 = ~n24033 & ~n24045;
  assign n24047 = controllable_DEQ & ~n24046;
  assign n24048 = ~n22663 & ~n24039;
  assign n24049 = ~controllable_DEQ & ~n24048;
  assign n24050 = ~n24047 & ~n24049;
  assign n24051 = ~i_FULL & ~n24050;
  assign n24052 = ~n24043 & ~n24051;
  assign n24053 = i_nEMPTY & ~n24052;
  assign n24054 = ~n13065 & ~n15964;
  assign n24055 = ~i_RtoB_ACK0 & ~n24054;
  assign n24056 = ~n15960 & ~n24055;
  assign n24057 = controllable_DEQ & ~n24056;
  assign n24058 = ~n13035 & ~n18792;
  assign n24059 = i_RtoB_ACK0 & ~n24058;
  assign n24060 = ~n22677 & ~n24059;
  assign n24061 = ~controllable_DEQ & ~n24060;
  assign n24062 = ~n24057 & ~n24061;
  assign n24063 = i_FULL & ~n24062;
  assign n24064 = ~n13075 & ~n15999;
  assign n24065 = ~i_RtoB_ACK0 & ~n24064;
  assign n24066 = ~n15995 & ~n24065;
  assign n24067 = controllable_DEQ & ~n24066;
  assign n24068 = ~n22687 & ~n24033;
  assign n24069 = ~controllable_DEQ & ~n24068;
  assign n24070 = ~n24067 & ~n24069;
  assign n24071 = ~i_FULL & ~n24070;
  assign n24072 = ~n24063 & ~n24071;
  assign n24073 = ~i_nEMPTY & ~n24072;
  assign n24074 = ~n24053 & ~n24073;
  assign n24075 = controllable_BtoS_ACK0 & ~n24074;
  assign n24076 = ~n13089 & ~n18811;
  assign n24077 = i_RtoB_ACK0 & ~n24076;
  assign n24078 = ~n13093 & ~n16031;
  assign n24079 = ~i_RtoB_ACK0 & ~n24078;
  assign n24080 = ~n24077 & ~n24079;
  assign n24081 = controllable_DEQ & ~n24080;
  assign n24082 = ~n13099 & ~n18819;
  assign n24083 = i_RtoB_ACK0 & ~n24082;
  assign n24084 = ~n22705 & ~n24083;
  assign n24085 = ~controllable_DEQ & ~n24084;
  assign n24086 = ~n24081 & ~n24085;
  assign n24087 = i_FULL & ~n24086;
  assign n24088 = ~n13107 & ~n16069;
  assign n24089 = ~i_RtoB_ACK0 & ~n24088;
  assign n24090 = ~n24077 & ~n24089;
  assign n24091 = controllable_DEQ & ~n24090;
  assign n24092 = ~n22715 & ~n24083;
  assign n24093 = ~controllable_DEQ & ~n24092;
  assign n24094 = ~n24091 & ~n24093;
  assign n24095 = ~i_FULL & ~n24094;
  assign n24096 = ~n24087 & ~n24095;
  assign n24097 = i_nEMPTY & ~n24096;
  assign n24098 = ~n13119 & ~n16106;
  assign n24099 = ~i_RtoB_ACK0 & ~n24098;
  assign n24100 = ~n16102 & ~n24099;
  assign n24101 = controllable_DEQ & ~n24100;
  assign n24102 = ~n13089 & ~n18837;
  assign n24103 = i_RtoB_ACK0 & ~n24102;
  assign n24104 = ~n22729 & ~n24103;
  assign n24105 = ~controllable_DEQ & ~n24104;
  assign n24106 = ~n24101 & ~n24105;
  assign n24107 = i_FULL & ~n24106;
  assign n24108 = ~n13129 & ~n16141;
  assign n24109 = ~i_RtoB_ACK0 & ~n24108;
  assign n24110 = ~n16137 & ~n24109;
  assign n24111 = controllable_DEQ & ~n24110;
  assign n24112 = ~n22739 & ~n24077;
  assign n24113 = ~controllable_DEQ & ~n24112;
  assign n24114 = ~n24111 & ~n24113;
  assign n24115 = ~i_FULL & ~n24114;
  assign n24116 = ~n24107 & ~n24115;
  assign n24117 = ~i_nEMPTY & ~n24116;
  assign n24118 = ~n24097 & ~n24117;
  assign n24119 = ~controllable_BtoS_ACK0 & ~n24118;
  assign n24120 = ~n24075 & ~n24119;
  assign n24121 = n4465 & ~n24120;
  assign n24122 = ~n22843 & ~n24121;
  assign n24123 = ~i_StoB_REQ10 & ~n24122;
  assign n24124 = ~n24031 & ~n24123;
  assign n24125 = ~controllable_BtoS_ACK10 & ~n24124;
  assign n24126 = ~n23927 & ~n24125;
  assign n24127 = ~n4464 & ~n24126;
  assign n24128 = ~n23875 & ~n24127;
  assign n24129 = ~n4463 & ~n24128;
  assign n24130 = ~n23523 & ~n24129;
  assign n24131 = ~n4462 & ~n24130;
  assign n24132 = ~n23045 & ~n24131;
  assign n24133 = n4461 & ~n24132;
  assign n24134 = ~n5029 & ~n14741;
  assign n24135 = i_RtoB_ACK0 & ~n24134;
  assign n24136 = ~n13157 & ~n14598;
  assign n24137 = ~i_RtoB_ACK0 & ~n24136;
  assign n24138 = ~n24135 & ~n24137;
  assign n24139 = controllable_DEQ & ~n24138;
  assign n24140 = ~n5052 & ~n14757;
  assign n24141 = i_RtoB_ACK0 & ~n24140;
  assign n24142 = ~n21993 & ~n24141;
  assign n24143 = ~controllable_DEQ & ~n24142;
  assign n24144 = ~n24139 & ~n24143;
  assign n24145 = i_nEMPTY & ~n24144;
  assign n24146 = ~n22015 & ~n24135;
  assign n24147 = ~controllable_DEQ & ~n24146;
  assign n24148 = ~n20915 & ~n24147;
  assign n24149 = i_FULL & ~n24148;
  assign n24150 = ~n13172 & ~n14598;
  assign n24151 = ~i_RtoB_ACK0 & ~n24150;
  assign n24152 = ~n24135 & ~n24151;
  assign n24153 = ~controllable_DEQ & ~n24152;
  assign n24154 = ~n20925 & ~n24153;
  assign n24155 = ~i_FULL & ~n24154;
  assign n24156 = ~n24149 & ~n24155;
  assign n24157 = ~i_nEMPTY & ~n24156;
  assign n24158 = ~n24145 & ~n24157;
  assign n24159 = controllable_BtoS_ACK0 & ~n24158;
  assign n24160 = ~n5126 & ~n16723;
  assign n24161 = i_RtoB_ACK0 & ~n24160;
  assign n24162 = ~n13184 & ~n14673;
  assign n24163 = ~i_RtoB_ACK0 & ~n24162;
  assign n24164 = ~n24161 & ~n24163;
  assign n24165 = controllable_DEQ & ~n24164;
  assign n24166 = ~n5149 & ~n16729;
  assign n24167 = i_RtoB_ACK0 & ~n24166;
  assign n24168 = ~n22043 & ~n24167;
  assign n24169 = ~controllable_DEQ & ~n24168;
  assign n24170 = ~n24165 & ~n24169;
  assign n24171 = i_nEMPTY & ~n24170;
  assign n24172 = ~n22065 & ~n24161;
  assign n24173 = ~controllable_DEQ & ~n24172;
  assign n24174 = ~n20953 & ~n24173;
  assign n24175 = i_FULL & ~n24174;
  assign n24176 = ~n13199 & ~n14673;
  assign n24177 = ~i_RtoB_ACK0 & ~n24176;
  assign n24178 = ~n24161 & ~n24177;
  assign n24179 = ~controllable_DEQ & ~n24178;
  assign n24180 = ~n20963 & ~n24179;
  assign n24181 = ~i_FULL & ~n24180;
  assign n24182 = ~n24175 & ~n24181;
  assign n24183 = ~i_nEMPTY & ~n24182;
  assign n24184 = ~n24171 & ~n24183;
  assign n24185 = ~controllable_BtoS_ACK0 & ~n24184;
  assign n24186 = ~n24159 & ~n24185;
  assign n24187 = n4465 & ~n24186;
  assign n24188 = ~n5340 & ~n16723;
  assign n24189 = i_RtoB_ACK0 & ~n24188;
  assign n24190 = ~n13213 & ~n14824;
  assign n24191 = ~i_RtoB_ACK0 & ~n24190;
  assign n24192 = ~n24189 & ~n24191;
  assign n24193 = controllable_DEQ & ~n24192;
  assign n24194 = ~n5363 & ~n16729;
  assign n24195 = i_RtoB_ACK0 & ~n24194;
  assign n24196 = ~n22095 & ~n24195;
  assign n24197 = ~controllable_DEQ & ~n24196;
  assign n24198 = ~n24193 & ~n24197;
  assign n24199 = i_nEMPTY & ~n24198;
  assign n24200 = ~n22117 & ~n24189;
  assign n24201 = ~controllable_DEQ & ~n24200;
  assign n24202 = ~n21031 & ~n24201;
  assign n24203 = i_FULL & ~n24202;
  assign n24204 = ~n13228 & ~n14824;
  assign n24205 = ~i_RtoB_ACK0 & ~n24204;
  assign n24206 = ~n24189 & ~n24205;
  assign n24207 = ~controllable_DEQ & ~n24206;
  assign n24208 = ~n21041 & ~n24207;
  assign n24209 = ~i_FULL & ~n24208;
  assign n24210 = ~n24203 & ~n24209;
  assign n24211 = ~i_nEMPTY & ~n24210;
  assign n24212 = ~n24199 & ~n24211;
  assign n24213 = ~controllable_BtoS_ACK0 & ~n24212;
  assign n24214 = ~n21013 & ~n24213;
  assign n24215 = ~n4465 & ~n24214;
  assign n24216 = ~n24187 & ~n24215;
  assign n24217 = i_StoB_REQ10 & ~n24216;
  assign n24218 = ~n6583 & ~n19074;
  assign n24219 = i_RtoB_ACK0 & ~n24218;
  assign n24220 = ~n13248 & ~n14904;
  assign n24221 = ~i_RtoB_ACK0 & ~n24220;
  assign n24222 = ~n24219 & ~n24221;
  assign n24223 = controllable_DEQ & ~n24222;
  assign n24224 = ~n6791 & ~n19088;
  assign n24225 = i_RtoB_ACK0 & ~n24224;
  assign n24226 = ~n13257 & ~n14923;
  assign n24227 = ~i_RtoB_ACK0 & ~n24226;
  assign n24228 = ~n24225 & ~n24227;
  assign n24229 = ~controllable_DEQ & ~n24228;
  assign n24230 = ~n24223 & ~n24229;
  assign n24231 = i_FULL & ~n24230;
  assign n24232 = ~n13267 & ~n14942;
  assign n24233 = ~i_RtoB_ACK0 & ~n24232;
  assign n24234 = ~n24219 & ~n24233;
  assign n24235 = controllable_DEQ & ~n24234;
  assign n24236 = ~n13275 & ~n14958;
  assign n24237 = ~i_RtoB_ACK0 & ~n24236;
  assign n24238 = ~n24225 & ~n24237;
  assign n24239 = ~controllable_DEQ & ~n24238;
  assign n24240 = ~n24235 & ~n24239;
  assign n24241 = ~i_FULL & ~n24240;
  assign n24242 = ~n24231 & ~n24241;
  assign n24243 = i_nEMPTY & ~n24242;
  assign n24244 = ~n6583 & ~n19130;
  assign n24245 = i_RtoB_ACK0 & ~n24244;
  assign n24246 = ~n13288 & ~n14995;
  assign n24247 = ~i_RtoB_ACK0 & ~n24246;
  assign n24248 = ~n24245 & ~n24247;
  assign n24249 = ~controllable_DEQ & ~n24248;
  assign n24250 = ~n21089 & ~n24249;
  assign n24251 = i_FULL & ~n24250;
  assign n24252 = ~n13296 & ~n14904;
  assign n24253 = ~i_RtoB_ACK0 & ~n24252;
  assign n24254 = ~n24219 & ~n24253;
  assign n24255 = ~controllable_DEQ & ~n24254;
  assign n24256 = ~n21101 & ~n24255;
  assign n24257 = ~i_FULL & ~n24256;
  assign n24258 = ~n24251 & ~n24257;
  assign n24259 = ~i_nEMPTY & ~n24258;
  assign n24260 = ~n24243 & ~n24259;
  assign n24261 = controllable_BtoS_ACK0 & ~n24260;
  assign n24262 = ~n6922 & ~n19167;
  assign n24263 = i_RtoB_ACK0 & ~n24262;
  assign n24264 = ~n13312 & ~n15046;
  assign n24265 = ~i_RtoB_ACK0 & ~n24264;
  assign n24266 = ~n24263 & ~n24265;
  assign n24267 = controllable_DEQ & ~n24266;
  assign n24268 = ~n6957 & ~n19181;
  assign n24269 = i_RtoB_ACK0 & ~n24268;
  assign n24270 = ~n13321 & ~n15065;
  assign n24271 = ~i_RtoB_ACK0 & ~n24270;
  assign n24272 = ~n24269 & ~n24271;
  assign n24273 = ~controllable_DEQ & ~n24272;
  assign n24274 = ~n24267 & ~n24273;
  assign n24275 = i_FULL & ~n24274;
  assign n24276 = ~n13331 & ~n15084;
  assign n24277 = ~i_RtoB_ACK0 & ~n24276;
  assign n24278 = ~n24263 & ~n24277;
  assign n24279 = controllable_DEQ & ~n24278;
  assign n24280 = ~n13339 & ~n15100;
  assign n24281 = ~i_RtoB_ACK0 & ~n24280;
  assign n24282 = ~n24269 & ~n24281;
  assign n24283 = ~controllable_DEQ & ~n24282;
  assign n24284 = ~n24279 & ~n24283;
  assign n24285 = ~i_FULL & ~n24284;
  assign n24286 = ~n24275 & ~n24285;
  assign n24287 = i_nEMPTY & ~n24286;
  assign n24288 = ~n6922 & ~n19223;
  assign n24289 = i_RtoB_ACK0 & ~n24288;
  assign n24290 = ~n13352 & ~n15137;
  assign n24291 = ~i_RtoB_ACK0 & ~n24290;
  assign n24292 = ~n24289 & ~n24291;
  assign n24293 = ~controllable_DEQ & ~n24292;
  assign n24294 = ~n21145 & ~n24293;
  assign n24295 = i_FULL & ~n24294;
  assign n24296 = ~n13360 & ~n15046;
  assign n24297 = ~i_RtoB_ACK0 & ~n24296;
  assign n24298 = ~n24263 & ~n24297;
  assign n24299 = ~controllable_DEQ & ~n24298;
  assign n24300 = ~n21157 & ~n24299;
  assign n24301 = ~i_FULL & ~n24300;
  assign n24302 = ~n24295 & ~n24301;
  assign n24303 = ~i_nEMPTY & ~n24302;
  assign n24304 = ~n24287 & ~n24303;
  assign n24305 = ~controllable_BtoS_ACK0 & ~n24304;
  assign n24306 = ~n24261 & ~n24305;
  assign n24307 = n4465 & ~n24306;
  assign n24308 = ~n7091 & ~n17280;
  assign n24309 = i_RtoB_ACK0 & ~n24308;
  assign n24310 = ~n13378 & ~n15190;
  assign n24311 = ~i_RtoB_ACK0 & ~n24310;
  assign n24312 = ~n24309 & ~n24311;
  assign n24313 = controllable_DEQ & ~n24312;
  assign n24314 = ~n7117 & ~n17288;
  assign n24315 = i_RtoB_ACK0 & ~n24314;
  assign n24316 = ~n13387 & ~n15209;
  assign n24317 = ~i_RtoB_ACK0 & ~n24316;
  assign n24318 = ~n24315 & ~n24317;
  assign n24319 = ~controllable_DEQ & ~n24318;
  assign n24320 = ~n24313 & ~n24319;
  assign n24321 = i_nEMPTY & ~n24320;
  assign n24322 = ~n7091 & ~n17298;
  assign n24323 = i_RtoB_ACK0 & ~n24322;
  assign n24324 = ~n13398 & ~n15237;
  assign n24325 = ~i_RtoB_ACK0 & ~n24324;
  assign n24326 = ~n24323 & ~n24325;
  assign n24327 = ~controllable_DEQ & ~n24326;
  assign n24328 = ~n21187 & ~n24327;
  assign n24329 = i_FULL & ~n24328;
  assign n24330 = ~n13406 & ~n15190;
  assign n24331 = ~i_RtoB_ACK0 & ~n24330;
  assign n24332 = ~n24309 & ~n24331;
  assign n24333 = ~controllable_DEQ & ~n24332;
  assign n24334 = ~n21199 & ~n24333;
  assign n24335 = ~i_FULL & ~n24334;
  assign n24336 = ~n24329 & ~n24335;
  assign n24337 = ~i_nEMPTY & ~n24336;
  assign n24338 = ~n24321 & ~n24337;
  assign n24339 = controllable_BtoS_ACK0 & ~n24338;
  assign n24340 = ~n7244 & ~n16909;
  assign n24341 = i_RtoB_ACK0 & ~n24340;
  assign n24342 = ~n13418 & ~n15281;
  assign n24343 = ~i_RtoB_ACK0 & ~n24342;
  assign n24344 = ~n24341 & ~n24343;
  assign n24345 = controllable_DEQ & ~n24344;
  assign n24346 = ~n7283 & ~n16917;
  assign n24347 = i_RtoB_ACK0 & ~n24346;
  assign n24348 = ~n13424 & ~n15300;
  assign n24349 = ~i_RtoB_ACK0 & ~n24348;
  assign n24350 = ~n24347 & ~n24349;
  assign n24351 = ~controllable_DEQ & ~n24350;
  assign n24352 = ~n24345 & ~n24351;
  assign n24353 = i_FULL & ~n24352;
  assign n24354 = ~n13432 & ~n15319;
  assign n24355 = ~i_RtoB_ACK0 & ~n24354;
  assign n24356 = ~n24341 & ~n24355;
  assign n24357 = controllable_DEQ & ~n24356;
  assign n24358 = ~n13438 & ~n15335;
  assign n24359 = ~i_RtoB_ACK0 & ~n24358;
  assign n24360 = ~n24347 & ~n24359;
  assign n24361 = ~controllable_DEQ & ~n24360;
  assign n24362 = ~n24357 & ~n24361;
  assign n24363 = ~i_FULL & ~n24362;
  assign n24364 = ~n24353 & ~n24363;
  assign n24365 = i_nEMPTY & ~n24364;
  assign n24366 = ~n7244 & ~n16935;
  assign n24367 = i_RtoB_ACK0 & ~n24366;
  assign n24368 = ~n13448 & ~n15372;
  assign n24369 = ~i_RtoB_ACK0 & ~n24368;
  assign n24370 = ~n24367 & ~n24369;
  assign n24371 = ~controllable_DEQ & ~n24370;
  assign n24372 = ~n21243 & ~n24371;
  assign n24373 = i_FULL & ~n24372;
  assign n24374 = ~n13456 & ~n15281;
  assign n24375 = ~i_RtoB_ACK0 & ~n24374;
  assign n24376 = ~n24341 & ~n24375;
  assign n24377 = ~controllable_DEQ & ~n24376;
  assign n24378 = ~n21255 & ~n24377;
  assign n24379 = ~i_FULL & ~n24378;
  assign n24380 = ~n24373 & ~n24379;
  assign n24381 = ~i_nEMPTY & ~n24380;
  assign n24382 = ~n24365 & ~n24381;
  assign n24383 = ~controllable_BtoS_ACK0 & ~n24382;
  assign n24384 = ~n24339 & ~n24383;
  assign n24385 = ~n4465 & ~n24384;
  assign n24386 = ~n24307 & ~n24385;
  assign n24387 = ~i_StoB_REQ10 & ~n24386;
  assign n24388 = ~n24217 & ~n24387;
  assign n24389 = controllable_BtoS_ACK10 & ~n24388;
  assign n24390 = ~n7396 & ~n16960;
  assign n24391 = i_RtoB_ACK0 & ~n24390;
  assign n24392 = ~n13474 & ~n19384;
  assign n24393 = ~i_RtoB_ACK0 & ~n24392;
  assign n24394 = ~n24391 & ~n24393;
  assign n24395 = controllable_DEQ & ~n24394;
  assign n24396 = ~n7414 & ~n16968;
  assign n24397 = i_RtoB_ACK0 & ~n24396;
  assign n24398 = ~n13480 & ~n19393;
  assign n24399 = ~i_RtoB_ACK0 & ~n24398;
  assign n24400 = ~n24397 & ~n24399;
  assign n24401 = ~controllable_DEQ & ~n24400;
  assign n24402 = ~n24395 & ~n24401;
  assign n24403 = i_FULL & ~n24402;
  assign n24404 = ~n13488 & ~n19404;
  assign n24405 = ~i_RtoB_ACK0 & ~n24404;
  assign n24406 = ~n24391 & ~n24405;
  assign n24407 = controllable_DEQ & ~n24406;
  assign n24408 = ~n13494 & ~n19409;
  assign n24409 = ~i_RtoB_ACK0 & ~n24408;
  assign n24410 = ~n24397 & ~n24409;
  assign n24411 = ~controllable_DEQ & ~n24410;
  assign n24412 = ~n24407 & ~n24411;
  assign n24413 = ~i_FULL & ~n24412;
  assign n24414 = ~n24403 & ~n24413;
  assign n24415 = i_nEMPTY & ~n24414;
  assign n24416 = ~n7396 & ~n16986;
  assign n24417 = i_RtoB_ACK0 & ~n24416;
  assign n24418 = ~n13504 & ~n19427;
  assign n24419 = ~i_RtoB_ACK0 & ~n24418;
  assign n24420 = ~n24417 & ~n24419;
  assign n24421 = ~controllable_DEQ & ~n24420;
  assign n24422 = ~n21305 & ~n24421;
  assign n24423 = i_FULL & ~n24422;
  assign n24424 = ~controllable_DEQ & ~n24394;
  assign n24425 = ~n21317 & ~n24424;
  assign n24426 = ~i_FULL & ~n24425;
  assign n24427 = ~n24423 & ~n24426;
  assign n24428 = ~i_nEMPTY & ~n24427;
  assign n24429 = ~n24415 & ~n24428;
  assign n24430 = controllable_BtoS_ACK0 & ~n24429;
  assign n24431 = ~n7476 & ~n17004;
  assign n24432 = i_RtoB_ACK0 & ~n24431;
  assign n24433 = ~n13519 & ~n19450;
  assign n24434 = ~i_RtoB_ACK0 & ~n24433;
  assign n24435 = ~n24432 & ~n24434;
  assign n24436 = controllable_DEQ & ~n24435;
  assign n24437 = ~n7494 & ~n17012;
  assign n24438 = i_RtoB_ACK0 & ~n24437;
  assign n24439 = ~n13525 & ~n19459;
  assign n24440 = ~i_RtoB_ACK0 & ~n24439;
  assign n24441 = ~n24438 & ~n24440;
  assign n24442 = ~controllable_DEQ & ~n24441;
  assign n24443 = ~n24436 & ~n24442;
  assign n24444 = i_FULL & ~n24443;
  assign n24445 = ~n13533 & ~n19470;
  assign n24446 = ~i_RtoB_ACK0 & ~n24445;
  assign n24447 = ~n24432 & ~n24446;
  assign n24448 = controllable_DEQ & ~n24447;
  assign n24449 = ~n13539 & ~n19475;
  assign n24450 = ~i_RtoB_ACK0 & ~n24449;
  assign n24451 = ~n24438 & ~n24450;
  assign n24452 = ~controllable_DEQ & ~n24451;
  assign n24453 = ~n24448 & ~n24452;
  assign n24454 = ~i_FULL & ~n24453;
  assign n24455 = ~n24444 & ~n24454;
  assign n24456 = i_nEMPTY & ~n24455;
  assign n24457 = ~n7476 & ~n17030;
  assign n24458 = i_RtoB_ACK0 & ~n24457;
  assign n24459 = ~n13549 & ~n19493;
  assign n24460 = ~i_RtoB_ACK0 & ~n24459;
  assign n24461 = ~n24458 & ~n24460;
  assign n24462 = ~controllable_DEQ & ~n24461;
  assign n24463 = ~n21358 & ~n24462;
  assign n24464 = i_FULL & ~n24463;
  assign n24465 = ~controllable_DEQ & ~n24435;
  assign n24466 = ~n21370 & ~n24465;
  assign n24467 = ~i_FULL & ~n24466;
  assign n24468 = ~n24464 & ~n24467;
  assign n24469 = ~i_nEMPTY & ~n24468;
  assign n24470 = ~n24456 & ~n24469;
  assign n24471 = ~controllable_BtoS_ACK0 & ~n24470;
  assign n24472 = ~n24430 & ~n24471;
  assign n24473 = n4465 & ~n24472;
  assign n24474 = ~n7550 & ~n17050;
  assign n24475 = i_RtoB_ACK0 & ~n24474;
  assign n24476 = ~n13566 & ~n19518;
  assign n24477 = ~i_RtoB_ACK0 & ~n24476;
  assign n24478 = ~n24475 & ~n24477;
  assign n24479 = controllable_DEQ & ~n24478;
  assign n24480 = ~n7567 & ~n17058;
  assign n24481 = i_RtoB_ACK0 & ~n24480;
  assign n24482 = ~n13572 & ~n19523;
  assign n24483 = ~i_RtoB_ACK0 & ~n24482;
  assign n24484 = ~n24481 & ~n24483;
  assign n24485 = ~controllable_DEQ & ~n24484;
  assign n24486 = ~n24479 & ~n24485;
  assign n24487 = i_nEMPTY & ~n24486;
  assign n24488 = ~n7550 & ~n17068;
  assign n24489 = i_RtoB_ACK0 & ~n24488;
  assign n24490 = ~n13580 & ~n19535;
  assign n24491 = ~i_RtoB_ACK0 & ~n24490;
  assign n24492 = ~n24489 & ~n24491;
  assign n24493 = ~controllable_DEQ & ~n24492;
  assign n24494 = ~n21397 & ~n24493;
  assign n24495 = i_FULL & ~n24494;
  assign n24496 = ~controllable_DEQ & ~n24478;
  assign n24497 = ~n21409 & ~n24496;
  assign n24498 = ~i_FULL & ~n24497;
  assign n24499 = ~n24495 & ~n24498;
  assign n24500 = ~i_nEMPTY & ~n24499;
  assign n24501 = ~n24487 & ~n24500;
  assign n24502 = controllable_BtoS_ACK0 & ~n24501;
  assign n24503 = ~n7612 & ~n17086;
  assign n24504 = i_RtoB_ACK0 & ~n24503;
  assign n24505 = ~n13595 & ~n19554;
  assign n24506 = ~i_RtoB_ACK0 & ~n24505;
  assign n24507 = ~n24504 & ~n24506;
  assign n24508 = controllable_DEQ & ~n24507;
  assign n24509 = ~n7630 & ~n17094;
  assign n24510 = i_RtoB_ACK0 & ~n24509;
  assign n24511 = ~n13424 & ~n19559;
  assign n24512 = ~i_RtoB_ACK0 & ~n24511;
  assign n24513 = ~n24510 & ~n24512;
  assign n24514 = ~controllable_DEQ & ~n24513;
  assign n24515 = ~n24508 & ~n24514;
  assign n24516 = i_FULL & ~n24515;
  assign n24517 = ~n13605 & ~n19566;
  assign n24518 = ~i_RtoB_ACK0 & ~n24517;
  assign n24519 = ~n24504 & ~n24518;
  assign n24520 = controllable_DEQ & ~n24519;
  assign n24521 = ~n13438 & ~n19571;
  assign n24522 = ~i_RtoB_ACK0 & ~n24521;
  assign n24523 = ~n24510 & ~n24522;
  assign n24524 = ~controllable_DEQ & ~n24523;
  assign n24525 = ~n24520 & ~n24524;
  assign n24526 = ~i_FULL & ~n24525;
  assign n24527 = ~n24516 & ~n24526;
  assign n24528 = i_nEMPTY & ~n24527;
  assign n24529 = ~n7612 & ~n17112;
  assign n24530 = i_RtoB_ACK0 & ~n24529;
  assign n24531 = ~n13448 & ~n19585;
  assign n24532 = ~i_RtoB_ACK0 & ~n24531;
  assign n24533 = ~n24530 & ~n24532;
  assign n24534 = ~controllable_DEQ & ~n24533;
  assign n24535 = ~n21450 & ~n24534;
  assign n24536 = i_FULL & ~n24535;
  assign n24537 = ~controllable_DEQ & ~n24507;
  assign n24538 = ~n21462 & ~n24537;
  assign n24539 = ~i_FULL & ~n24538;
  assign n24540 = ~n24536 & ~n24539;
  assign n24541 = ~i_nEMPTY & ~n24540;
  assign n24542 = ~n24528 & ~n24541;
  assign n24543 = ~controllable_BtoS_ACK0 & ~n24542;
  assign n24544 = ~n24502 & ~n24543;
  assign n24545 = ~n4465 & ~n24544;
  assign n24546 = ~n24473 & ~n24545;
  assign n24547 = i_StoB_REQ10 & ~n24546;
  assign n24548 = ~n24387 & ~n24547;
  assign n24549 = ~controllable_BtoS_ACK10 & ~n24548;
  assign n24550 = ~n24389 & ~n24549;
  assign n24551 = n4464 & ~n24550;
  assign n24552 = ~n7707 & ~n14741;
  assign n24553 = i_RtoB_ACK0 & ~n24552;
  assign n24554 = ~n13636 & ~n15732;
  assign n24555 = ~i_RtoB_ACK0 & ~n24554;
  assign n24556 = ~n24553 & ~n24555;
  assign n24557 = controllable_DEQ & ~n24556;
  assign n24558 = ~n7730 & ~n14757;
  assign n24559 = i_RtoB_ACK0 & ~n24558;
  assign n24560 = ~n22547 & ~n24559;
  assign n24561 = ~controllable_DEQ & ~n24560;
  assign n24562 = ~n24557 & ~n24561;
  assign n24563 = i_nEMPTY & ~n24562;
  assign n24564 = ~n22569 & ~n24553;
  assign n24565 = ~controllable_DEQ & ~n24564;
  assign n24566 = ~n21495 & ~n24565;
  assign n24567 = i_FULL & ~n24566;
  assign n24568 = ~n13651 & ~n15732;
  assign n24569 = ~i_RtoB_ACK0 & ~n24568;
  assign n24570 = ~n24553 & ~n24569;
  assign n24571 = ~controllable_DEQ & ~n24570;
  assign n24572 = ~n21505 & ~n24571;
  assign n24573 = ~i_FULL & ~n24572;
  assign n24574 = ~n24567 & ~n24573;
  assign n24575 = ~i_nEMPTY & ~n24574;
  assign n24576 = ~n24563 & ~n24575;
  assign n24577 = controllable_BtoS_ACK0 & ~n24576;
  assign n24578 = ~n7799 & ~n16723;
  assign n24579 = i_RtoB_ACK0 & ~n24578;
  assign n24580 = ~n13663 & ~n15807;
  assign n24581 = ~i_RtoB_ACK0 & ~n24580;
  assign n24582 = ~n24579 & ~n24581;
  assign n24583 = controllable_DEQ & ~n24582;
  assign n24584 = ~n7822 & ~n16729;
  assign n24585 = i_RtoB_ACK0 & ~n24584;
  assign n24586 = ~n22597 & ~n24585;
  assign n24587 = ~controllable_DEQ & ~n24586;
  assign n24588 = ~n24583 & ~n24587;
  assign n24589 = i_nEMPTY & ~n24588;
  assign n24590 = ~n22619 & ~n24579;
  assign n24591 = ~controllable_DEQ & ~n24590;
  assign n24592 = ~n21533 & ~n24591;
  assign n24593 = i_FULL & ~n24592;
  assign n24594 = ~n13678 & ~n15807;
  assign n24595 = ~i_RtoB_ACK0 & ~n24594;
  assign n24596 = ~n24579 & ~n24595;
  assign n24597 = ~controllable_DEQ & ~n24596;
  assign n24598 = ~n21543 & ~n24597;
  assign n24599 = ~i_FULL & ~n24598;
  assign n24600 = ~n24593 & ~n24599;
  assign n24601 = ~i_nEMPTY & ~n24600;
  assign n24602 = ~n24589 & ~n24601;
  assign n24603 = ~controllable_BtoS_ACK0 & ~n24602;
  assign n24604 = ~n24577 & ~n24603;
  assign n24605 = n4465 & ~n24604;
  assign n24606 = ~n21013 & ~n24603;
  assign n24607 = ~n4465 & ~n24606;
  assign n24608 = ~n24605 & ~n24607;
  assign n24609 = i_StoB_REQ10 & ~n24608;
  assign n24610 = ~n7919 & ~n18766;
  assign n24611 = i_RtoB_ACK0 & ~n24610;
  assign n24612 = ~n13700 & ~n15889;
  assign n24613 = ~i_RtoB_ACK0 & ~n24612;
  assign n24614 = ~n24611 & ~n24613;
  assign n24615 = controllable_DEQ & ~n24614;
  assign n24616 = ~n7953 & ~n18774;
  assign n24617 = i_RtoB_ACK0 & ~n24616;
  assign n24618 = ~n13709 & ~n15908;
  assign n24619 = ~i_RtoB_ACK0 & ~n24618;
  assign n24620 = ~n24617 & ~n24619;
  assign n24621 = ~controllable_DEQ & ~n24620;
  assign n24622 = ~n24615 & ~n24621;
  assign n24623 = i_FULL & ~n24622;
  assign n24624 = ~n13719 & ~n15927;
  assign n24625 = ~i_RtoB_ACK0 & ~n24624;
  assign n24626 = ~n24611 & ~n24625;
  assign n24627 = controllable_DEQ & ~n24626;
  assign n24628 = ~n13727 & ~n15943;
  assign n24629 = ~i_RtoB_ACK0 & ~n24628;
  assign n24630 = ~n24617 & ~n24629;
  assign n24631 = ~controllable_DEQ & ~n24630;
  assign n24632 = ~n24627 & ~n24631;
  assign n24633 = ~i_FULL & ~n24632;
  assign n24634 = ~n24623 & ~n24633;
  assign n24635 = i_nEMPTY & ~n24634;
  assign n24636 = ~n7919 & ~n18792;
  assign n24637 = i_RtoB_ACK0 & ~n24636;
  assign n24638 = ~n13740 & ~n15980;
  assign n24639 = ~i_RtoB_ACK0 & ~n24638;
  assign n24640 = ~n24637 & ~n24639;
  assign n24641 = ~controllable_DEQ & ~n24640;
  assign n24642 = ~n21593 & ~n24641;
  assign n24643 = i_FULL & ~n24642;
  assign n24644 = ~n13748 & ~n15889;
  assign n24645 = ~i_RtoB_ACK0 & ~n24644;
  assign n24646 = ~n24611 & ~n24645;
  assign n24647 = ~controllable_DEQ & ~n24646;
  assign n24648 = ~n21605 & ~n24647;
  assign n24649 = ~i_FULL & ~n24648;
  assign n24650 = ~n24643 & ~n24649;
  assign n24651 = ~i_nEMPTY & ~n24650;
  assign n24652 = ~n24635 & ~n24651;
  assign n24653 = controllable_BtoS_ACK0 & ~n24652;
  assign n24654 = ~n8086 & ~n18811;
  assign n24655 = i_RtoB_ACK0 & ~n24654;
  assign n24656 = ~n13764 & ~n16031;
  assign n24657 = ~i_RtoB_ACK0 & ~n24656;
  assign n24658 = ~n24655 & ~n24657;
  assign n24659 = controllable_DEQ & ~n24658;
  assign n24660 = ~n8117 & ~n18819;
  assign n24661 = i_RtoB_ACK0 & ~n24660;
  assign n24662 = ~n13773 & ~n16050;
  assign n24663 = ~i_RtoB_ACK0 & ~n24662;
  assign n24664 = ~n24661 & ~n24663;
  assign n24665 = ~controllable_DEQ & ~n24664;
  assign n24666 = ~n24659 & ~n24665;
  assign n24667 = i_FULL & ~n24666;
  assign n24668 = ~n13783 & ~n16069;
  assign n24669 = ~i_RtoB_ACK0 & ~n24668;
  assign n24670 = ~n24655 & ~n24669;
  assign n24671 = controllable_DEQ & ~n24670;
  assign n24672 = ~n13791 & ~n16085;
  assign n24673 = ~i_RtoB_ACK0 & ~n24672;
  assign n24674 = ~n24661 & ~n24673;
  assign n24675 = ~controllable_DEQ & ~n24674;
  assign n24676 = ~n24671 & ~n24675;
  assign n24677 = ~i_FULL & ~n24676;
  assign n24678 = ~n24667 & ~n24677;
  assign n24679 = i_nEMPTY & ~n24678;
  assign n24680 = ~n8086 & ~n18837;
  assign n24681 = i_RtoB_ACK0 & ~n24680;
  assign n24682 = ~n13804 & ~n16122;
  assign n24683 = ~i_RtoB_ACK0 & ~n24682;
  assign n24684 = ~n24681 & ~n24683;
  assign n24685 = ~controllable_DEQ & ~n24684;
  assign n24686 = ~n21649 & ~n24685;
  assign n24687 = i_FULL & ~n24686;
  assign n24688 = ~n13812 & ~n16031;
  assign n24689 = ~i_RtoB_ACK0 & ~n24688;
  assign n24690 = ~n24655 & ~n24689;
  assign n24691 = ~controllable_DEQ & ~n24690;
  assign n24692 = ~n21661 & ~n24691;
  assign n24693 = ~i_FULL & ~n24692;
  assign n24694 = ~n24687 & ~n24693;
  assign n24695 = ~i_nEMPTY & ~n24694;
  assign n24696 = ~n24679 & ~n24695;
  assign n24697 = ~controllable_BtoS_ACK0 & ~n24696;
  assign n24698 = ~n24653 & ~n24697;
  assign n24699 = n4465 & ~n24698;
  assign n24700 = ~n8229 & ~n17280;
  assign n24701 = i_RtoB_ACK0 & ~n24700;
  assign n24702 = ~n13826 & ~n16175;
  assign n24703 = ~i_RtoB_ACK0 & ~n24702;
  assign n24704 = ~n24701 & ~n24703;
  assign n24705 = controllable_DEQ & ~n24704;
  assign n24706 = ~n8254 & ~n17288;
  assign n24707 = i_RtoB_ACK0 & ~n24706;
  assign n24708 = ~n13832 & ~n16194;
  assign n24709 = ~i_RtoB_ACK0 & ~n24708;
  assign n24710 = ~n24707 & ~n24709;
  assign n24711 = ~controllable_DEQ & ~n24710;
  assign n24712 = ~n24705 & ~n24711;
  assign n24713 = i_nEMPTY & ~n24712;
  assign n24714 = ~n8229 & ~n17298;
  assign n24715 = i_RtoB_ACK0 & ~n24714;
  assign n24716 = ~n13840 & ~n16220;
  assign n24717 = ~i_RtoB_ACK0 & ~n24716;
  assign n24718 = ~n24715 & ~n24717;
  assign n24719 = ~controllable_DEQ & ~n24718;
  assign n24720 = ~n21691 & ~n24719;
  assign n24721 = i_FULL & ~n24720;
  assign n24722 = ~n13848 & ~n16175;
  assign n24723 = ~i_RtoB_ACK0 & ~n24722;
  assign n24724 = ~n24701 & ~n24723;
  assign n24725 = ~controllable_DEQ & ~n24724;
  assign n24726 = ~n21703 & ~n24725;
  assign n24727 = ~i_FULL & ~n24726;
  assign n24728 = ~n24721 & ~n24727;
  assign n24729 = ~i_nEMPTY & ~n24728;
  assign n24730 = ~n24713 & ~n24729;
  assign n24731 = controllable_BtoS_ACK0 & ~n24730;
  assign n24732 = ~n8329 & ~n17317;
  assign n24733 = i_RtoB_ACK0 & ~n24732;
  assign n24734 = ~n13860 & ~n16262;
  assign n24735 = ~i_RtoB_ACK0 & ~n24734;
  assign n24736 = ~n24733 & ~n24735;
  assign n24737 = controllable_DEQ & ~n24736;
  assign n24738 = ~n8358 & ~n17325;
  assign n24739 = i_RtoB_ACK0 & ~n24738;
  assign n24740 = ~n13866 & ~n16281;
  assign n24741 = ~i_RtoB_ACK0 & ~n24740;
  assign n24742 = ~n24739 & ~n24741;
  assign n24743 = ~controllable_DEQ & ~n24742;
  assign n24744 = ~n24737 & ~n24743;
  assign n24745 = i_FULL & ~n24744;
  assign n24746 = ~n13874 & ~n16300;
  assign n24747 = ~i_RtoB_ACK0 & ~n24746;
  assign n24748 = ~n24733 & ~n24747;
  assign n24749 = controllable_DEQ & ~n24748;
  assign n24750 = ~n13880 & ~n16316;
  assign n24751 = ~i_RtoB_ACK0 & ~n24750;
  assign n24752 = ~n24739 & ~n24751;
  assign n24753 = ~controllable_DEQ & ~n24752;
  assign n24754 = ~n24749 & ~n24753;
  assign n24755 = ~i_FULL & ~n24754;
  assign n24756 = ~n24745 & ~n24755;
  assign n24757 = i_nEMPTY & ~n24756;
  assign n24758 = ~n8329 & ~n17343;
  assign n24759 = i_RtoB_ACK0 & ~n24758;
  assign n24760 = ~n13890 & ~n16353;
  assign n24761 = ~i_RtoB_ACK0 & ~n24760;
  assign n24762 = ~n24759 & ~n24761;
  assign n24763 = ~controllable_DEQ & ~n24762;
  assign n24764 = ~n21747 & ~n24763;
  assign n24765 = i_FULL & ~n24764;
  assign n24766 = ~n13898 & ~n16262;
  assign n24767 = ~i_RtoB_ACK0 & ~n24766;
  assign n24768 = ~n24733 & ~n24767;
  assign n24769 = ~controllable_DEQ & ~n24768;
  assign n24770 = ~n21759 & ~n24769;
  assign n24771 = ~i_FULL & ~n24770;
  assign n24772 = ~n24765 & ~n24771;
  assign n24773 = ~i_nEMPTY & ~n24772;
  assign n24774 = ~n24757 & ~n24773;
  assign n24775 = ~controllable_BtoS_ACK0 & ~n24774;
  assign n24776 = ~n24731 & ~n24775;
  assign n24777 = ~n4465 & ~n24776;
  assign n24778 = ~n24699 & ~n24777;
  assign n24779 = ~i_StoB_REQ10 & ~n24778;
  assign n24780 = ~n24609 & ~n24779;
  assign n24781 = controllable_BtoS_ACK10 & ~n24780;
  assign n24782 = ~n8466 & ~n17368;
  assign n24783 = i_RtoB_ACK0 & ~n24782;
  assign n24784 = ~n13916 & ~n20002;
  assign n24785 = ~i_RtoB_ACK0 & ~n24784;
  assign n24786 = ~n24783 & ~n24785;
  assign n24787 = controllable_DEQ & ~n24786;
  assign n24788 = ~n8484 & ~n17376;
  assign n24789 = i_RtoB_ACK0 & ~n24788;
  assign n24790 = ~n13922 & ~n20011;
  assign n24791 = ~i_RtoB_ACK0 & ~n24790;
  assign n24792 = ~n24789 & ~n24791;
  assign n24793 = ~controllable_DEQ & ~n24792;
  assign n24794 = ~n24787 & ~n24793;
  assign n24795 = i_FULL & ~n24794;
  assign n24796 = ~n13930 & ~n20022;
  assign n24797 = ~i_RtoB_ACK0 & ~n24796;
  assign n24798 = ~n24783 & ~n24797;
  assign n24799 = controllable_DEQ & ~n24798;
  assign n24800 = ~n13936 & ~n20027;
  assign n24801 = ~i_RtoB_ACK0 & ~n24800;
  assign n24802 = ~n24789 & ~n24801;
  assign n24803 = ~controllable_DEQ & ~n24802;
  assign n24804 = ~n24799 & ~n24803;
  assign n24805 = ~i_FULL & ~n24804;
  assign n24806 = ~n24795 & ~n24805;
  assign n24807 = i_nEMPTY & ~n24806;
  assign n24808 = ~n8466 & ~n17394;
  assign n24809 = i_RtoB_ACK0 & ~n24808;
  assign n24810 = ~n13946 & ~n20045;
  assign n24811 = ~i_RtoB_ACK0 & ~n24810;
  assign n24812 = ~n24809 & ~n24811;
  assign n24813 = ~controllable_DEQ & ~n24812;
  assign n24814 = ~n21809 & ~n24813;
  assign n24815 = i_FULL & ~n24814;
  assign n24816 = ~controllable_DEQ & ~n24786;
  assign n24817 = ~n21821 & ~n24816;
  assign n24818 = ~i_FULL & ~n24817;
  assign n24819 = ~n24815 & ~n24818;
  assign n24820 = ~i_nEMPTY & ~n24819;
  assign n24821 = ~n24807 & ~n24820;
  assign n24822 = controllable_BtoS_ACK0 & ~n24821;
  assign n24823 = ~n8545 & ~n17412;
  assign n24824 = i_RtoB_ACK0 & ~n24823;
  assign n24825 = ~n13961 & ~n20068;
  assign n24826 = ~i_RtoB_ACK0 & ~n24825;
  assign n24827 = ~n24824 & ~n24826;
  assign n24828 = controllable_DEQ & ~n24827;
  assign n24829 = ~n8563 & ~n17420;
  assign n24830 = i_RtoB_ACK0 & ~n24829;
  assign n24831 = ~n13967 & ~n20073;
  assign n24832 = ~i_RtoB_ACK0 & ~n24831;
  assign n24833 = ~n24830 & ~n24832;
  assign n24834 = ~controllable_DEQ & ~n24833;
  assign n24835 = ~n24828 & ~n24834;
  assign n24836 = i_FULL & ~n24835;
  assign n24837 = ~n13975 & ~n20080;
  assign n24838 = ~i_RtoB_ACK0 & ~n24837;
  assign n24839 = ~n24824 & ~n24838;
  assign n24840 = controllable_DEQ & ~n24839;
  assign n24841 = ~n13981 & ~n20085;
  assign n24842 = ~i_RtoB_ACK0 & ~n24841;
  assign n24843 = ~n24830 & ~n24842;
  assign n24844 = ~controllable_DEQ & ~n24843;
  assign n24845 = ~n24840 & ~n24844;
  assign n24846 = ~i_FULL & ~n24845;
  assign n24847 = ~n24836 & ~n24846;
  assign n24848 = i_nEMPTY & ~n24847;
  assign n24849 = ~n8545 & ~n17438;
  assign n24850 = i_RtoB_ACK0 & ~n24849;
  assign n24851 = ~n13991 & ~n20099;
  assign n24852 = ~i_RtoB_ACK0 & ~n24851;
  assign n24853 = ~n24850 & ~n24852;
  assign n24854 = ~controllable_DEQ & ~n24853;
  assign n24855 = ~n21862 & ~n24854;
  assign n24856 = i_FULL & ~n24855;
  assign n24857 = ~controllable_DEQ & ~n24827;
  assign n24858 = ~n21874 & ~n24857;
  assign n24859 = ~i_FULL & ~n24858;
  assign n24860 = ~n24856 & ~n24859;
  assign n24861 = ~i_nEMPTY & ~n24860;
  assign n24862 = ~n24848 & ~n24861;
  assign n24863 = ~controllable_BtoS_ACK0 & ~n24862;
  assign n24864 = ~n24822 & ~n24863;
  assign n24865 = n4465 & ~n24864;
  assign n24866 = ~n8619 & ~n17050;
  assign n24867 = i_RtoB_ACK0 & ~n24866;
  assign n24868 = ~n14008 & ~n20120;
  assign n24869 = ~i_RtoB_ACK0 & ~n24868;
  assign n24870 = ~n24867 & ~n24869;
  assign n24871 = controllable_DEQ & ~n24870;
  assign n24872 = ~n8635 & ~n17058;
  assign n24873 = i_RtoB_ACK0 & ~n24872;
  assign n24874 = ~n13832 & ~n20125;
  assign n24875 = ~i_RtoB_ACK0 & ~n24874;
  assign n24876 = ~n24873 & ~n24875;
  assign n24877 = ~controllable_DEQ & ~n24876;
  assign n24878 = ~n24871 & ~n24877;
  assign n24879 = i_nEMPTY & ~n24878;
  assign n24880 = ~n8619 & ~n17068;
  assign n24881 = i_RtoB_ACK0 & ~n24880;
  assign n24882 = ~n13840 & ~n20137;
  assign n24883 = ~i_RtoB_ACK0 & ~n24882;
  assign n24884 = ~n24881 & ~n24883;
  assign n24885 = ~controllable_DEQ & ~n24884;
  assign n24886 = ~n21901 & ~n24885;
  assign n24887 = i_FULL & ~n24886;
  assign n24888 = ~controllable_DEQ & ~n24870;
  assign n24889 = ~n21913 & ~n24888;
  assign n24890 = ~i_FULL & ~n24889;
  assign n24891 = ~n24887 & ~n24890;
  assign n24892 = ~i_nEMPTY & ~n24891;
  assign n24893 = ~n24879 & ~n24892;
  assign n24894 = controllable_BtoS_ACK0 & ~n24893;
  assign n24895 = ~n8677 & ~n17481;
  assign n24896 = i_RtoB_ACK0 & ~n24895;
  assign n24897 = ~n14029 & ~n20156;
  assign n24898 = ~i_RtoB_ACK0 & ~n24897;
  assign n24899 = ~n24896 & ~n24898;
  assign n24900 = controllable_DEQ & ~n24899;
  assign n24901 = ~n8695 & ~n17489;
  assign n24902 = i_RtoB_ACK0 & ~n24901;
  assign n24903 = ~n13866 & ~n20161;
  assign n24904 = ~i_RtoB_ACK0 & ~n24903;
  assign n24905 = ~n24902 & ~n24904;
  assign n24906 = ~controllable_DEQ & ~n24905;
  assign n24907 = ~n24900 & ~n24906;
  assign n24908 = i_FULL & ~n24907;
  assign n24909 = ~n14039 & ~n20168;
  assign n24910 = ~i_RtoB_ACK0 & ~n24909;
  assign n24911 = ~n24896 & ~n24910;
  assign n24912 = controllable_DEQ & ~n24911;
  assign n24913 = ~n13880 & ~n20173;
  assign n24914 = ~i_RtoB_ACK0 & ~n24913;
  assign n24915 = ~n24902 & ~n24914;
  assign n24916 = ~controllable_DEQ & ~n24915;
  assign n24917 = ~n24912 & ~n24916;
  assign n24918 = ~i_FULL & ~n24917;
  assign n24919 = ~n24908 & ~n24918;
  assign n24920 = i_nEMPTY & ~n24919;
  assign n24921 = ~n8677 & ~n17507;
  assign n24922 = i_RtoB_ACK0 & ~n24921;
  assign n24923 = ~n13890 & ~n20187;
  assign n24924 = ~i_RtoB_ACK0 & ~n24923;
  assign n24925 = ~n24922 & ~n24924;
  assign n24926 = ~controllable_DEQ & ~n24925;
  assign n24927 = ~n21954 & ~n24926;
  assign n24928 = i_FULL & ~n24927;
  assign n24929 = ~controllable_DEQ & ~n24899;
  assign n24930 = ~n21966 & ~n24929;
  assign n24931 = ~i_FULL & ~n24930;
  assign n24932 = ~n24928 & ~n24931;
  assign n24933 = ~i_nEMPTY & ~n24932;
  assign n24934 = ~n24920 & ~n24933;
  assign n24935 = ~controllable_BtoS_ACK0 & ~n24934;
  assign n24936 = ~n24894 & ~n24935;
  assign n24937 = ~n4465 & ~n24936;
  assign n24938 = ~n24865 & ~n24937;
  assign n24939 = i_StoB_REQ10 & ~n24938;
  assign n24940 = ~n24779 & ~n24939;
  assign n24941 = ~controllable_BtoS_ACK10 & ~n24940;
  assign n24942 = ~n24781 & ~n24941;
  assign n24943 = ~n4464 & ~n24942;
  assign n24944 = ~n24551 & ~n24943;
  assign n24945 = n4463 & ~n24944;
  assign n24946 = ~n9297 & ~n19074;
  assign n24947 = i_RtoB_ACK0 & ~n24946;
  assign n24948 = ~n22143 & ~n24947;
  assign n24949 = controllable_DEQ & ~n24948;
  assign n24950 = ~n9514 & ~n19088;
  assign n24951 = i_RtoB_ACK0 & ~n24950;
  assign n24952 = ~n22149 & ~n24951;
  assign n24953 = ~controllable_DEQ & ~n24952;
  assign n24954 = ~n24949 & ~n24953;
  assign n24955 = i_FULL & ~n24954;
  assign n24956 = ~n22155 & ~n24947;
  assign n24957 = controllable_DEQ & ~n24956;
  assign n24958 = ~n22159 & ~n24951;
  assign n24959 = ~controllable_DEQ & ~n24958;
  assign n24960 = ~n24957 & ~n24959;
  assign n24961 = ~i_FULL & ~n24960;
  assign n24962 = ~n24955 & ~n24961;
  assign n24963 = i_nEMPTY & ~n24962;
  assign n24964 = ~n9297 & ~n19130;
  assign n24965 = i_RtoB_ACK0 & ~n24964;
  assign n24966 = ~n22173 & ~n24965;
  assign n24967 = ~controllable_DEQ & ~n24966;
  assign n24968 = ~n22169 & ~n24967;
  assign n24969 = i_FULL & ~n24968;
  assign n24970 = ~n22183 & ~n24947;
  assign n24971 = ~controllable_DEQ & ~n24970;
  assign n24972 = ~n22181 & ~n24971;
  assign n24973 = ~i_FULL & ~n24972;
  assign n24974 = ~n24969 & ~n24973;
  assign n24975 = ~i_nEMPTY & ~n24974;
  assign n24976 = ~n24963 & ~n24975;
  assign n24977 = controllable_BtoS_ACK0 & ~n24976;
  assign n24978 = ~n9628 & ~n19167;
  assign n24979 = i_RtoB_ACK0 & ~n24978;
  assign n24980 = ~n22195 & ~n24979;
  assign n24981 = controllable_DEQ & ~n24980;
  assign n24982 = ~n9661 & ~n19181;
  assign n24983 = i_RtoB_ACK0 & ~n24982;
  assign n24984 = ~n22201 & ~n24983;
  assign n24985 = ~controllable_DEQ & ~n24984;
  assign n24986 = ~n24981 & ~n24985;
  assign n24987 = i_FULL & ~n24986;
  assign n24988 = ~n22207 & ~n24979;
  assign n24989 = controllable_DEQ & ~n24988;
  assign n24990 = ~n22211 & ~n24983;
  assign n24991 = ~controllable_DEQ & ~n24990;
  assign n24992 = ~n24989 & ~n24991;
  assign n24993 = ~i_FULL & ~n24992;
  assign n24994 = ~n24987 & ~n24993;
  assign n24995 = i_nEMPTY & ~n24994;
  assign n24996 = ~n9628 & ~n19223;
  assign n24997 = i_RtoB_ACK0 & ~n24996;
  assign n24998 = ~n22225 & ~n24997;
  assign n24999 = ~controllable_DEQ & ~n24998;
  assign n25000 = ~n22221 & ~n24999;
  assign n25001 = i_FULL & ~n25000;
  assign n25002 = ~n22235 & ~n24979;
  assign n25003 = ~controllable_DEQ & ~n25002;
  assign n25004 = ~n22233 & ~n25003;
  assign n25005 = ~i_FULL & ~n25004;
  assign n25006 = ~n25001 & ~n25005;
  assign n25007 = ~i_nEMPTY & ~n25006;
  assign n25008 = ~n24995 & ~n25007;
  assign n25009 = ~controllable_BtoS_ACK0 & ~n25008;
  assign n25010 = ~n24977 & ~n25009;
  assign n25011 = n4465 & ~n25010;
  assign n25012 = ~n9785 & ~n17280;
  assign n25013 = i_RtoB_ACK0 & ~n25012;
  assign n25014 = ~n22249 & ~n25013;
  assign n25015 = controllable_DEQ & ~n25014;
  assign n25016 = ~n9808 & ~n17288;
  assign n25017 = i_RtoB_ACK0 & ~n25016;
  assign n25018 = ~n22255 & ~n25017;
  assign n25019 = ~controllable_DEQ & ~n25018;
  assign n25020 = ~n25015 & ~n25019;
  assign n25021 = i_nEMPTY & ~n25020;
  assign n25022 = ~n9785 & ~n17298;
  assign n25023 = i_RtoB_ACK0 & ~n25022;
  assign n25024 = ~n22267 & ~n25023;
  assign n25025 = ~controllable_DEQ & ~n25024;
  assign n25026 = ~n22263 & ~n25025;
  assign n25027 = i_FULL & ~n25026;
  assign n25028 = ~n22277 & ~n25013;
  assign n25029 = ~controllable_DEQ & ~n25028;
  assign n25030 = ~n22275 & ~n25029;
  assign n25031 = ~i_FULL & ~n25030;
  assign n25032 = ~n25027 & ~n25031;
  assign n25033 = ~i_nEMPTY & ~n25032;
  assign n25034 = ~n25021 & ~n25033;
  assign n25035 = controllable_BtoS_ACK0 & ~n25034;
  assign n25036 = ~n22337 & ~n25035;
  assign n25037 = ~n4465 & ~n25036;
  assign n25038 = ~n25011 & ~n25037;
  assign n25039 = ~i_StoB_REQ10 & ~n25038;
  assign n25040 = ~n22139 & ~n25039;
  assign n25041 = controllable_BtoS_ACK10 & ~n25040;
  assign n25042 = ~n22533 & ~n25039;
  assign n25043 = ~controllable_BtoS_ACK10 & ~n25042;
  assign n25044 = ~n25041 & ~n25043;
  assign n25045 = n4464 & ~n25044;
  assign n25046 = ~n10464 & ~n18766;
  assign n25047 = i_RtoB_ACK0 & ~n25046;
  assign n25048 = ~n22647 & ~n25047;
  assign n25049 = controllable_DEQ & ~n25048;
  assign n25050 = ~n10491 & ~n18774;
  assign n25051 = i_RtoB_ACK0 & ~n25050;
  assign n25052 = ~n22653 & ~n25051;
  assign n25053 = ~controllable_DEQ & ~n25052;
  assign n25054 = ~n25049 & ~n25053;
  assign n25055 = i_FULL & ~n25054;
  assign n25056 = ~n22659 & ~n25047;
  assign n25057 = controllable_DEQ & ~n25056;
  assign n25058 = ~n22663 & ~n25051;
  assign n25059 = ~controllable_DEQ & ~n25058;
  assign n25060 = ~n25057 & ~n25059;
  assign n25061 = ~i_FULL & ~n25060;
  assign n25062 = ~n25055 & ~n25061;
  assign n25063 = i_nEMPTY & ~n25062;
  assign n25064 = ~n10464 & ~n18792;
  assign n25065 = i_RtoB_ACK0 & ~n25064;
  assign n25066 = ~n22677 & ~n25065;
  assign n25067 = ~controllable_DEQ & ~n25066;
  assign n25068 = ~n22673 & ~n25067;
  assign n25069 = i_FULL & ~n25068;
  assign n25070 = ~n22687 & ~n25047;
  assign n25071 = ~controllable_DEQ & ~n25070;
  assign n25072 = ~n22685 & ~n25071;
  assign n25073 = ~i_FULL & ~n25072;
  assign n25074 = ~n25069 & ~n25073;
  assign n25075 = ~i_nEMPTY & ~n25074;
  assign n25076 = ~n25063 & ~n25075;
  assign n25077 = controllable_BtoS_ACK0 & ~n25076;
  assign n25078 = ~n10594 & ~n18811;
  assign n25079 = i_RtoB_ACK0 & ~n25078;
  assign n25080 = ~n22699 & ~n25079;
  assign n25081 = controllable_DEQ & ~n25080;
  assign n25082 = ~n10618 & ~n18819;
  assign n25083 = i_RtoB_ACK0 & ~n25082;
  assign n25084 = ~n22705 & ~n25083;
  assign n25085 = ~controllable_DEQ & ~n25084;
  assign n25086 = ~n25081 & ~n25085;
  assign n25087 = i_FULL & ~n25086;
  assign n25088 = ~n22711 & ~n25079;
  assign n25089 = controllable_DEQ & ~n25088;
  assign n25090 = ~n22715 & ~n25083;
  assign n25091 = ~controllable_DEQ & ~n25090;
  assign n25092 = ~n25089 & ~n25091;
  assign n25093 = ~i_FULL & ~n25092;
  assign n25094 = ~n25087 & ~n25093;
  assign n25095 = i_nEMPTY & ~n25094;
  assign n25096 = ~n10594 & ~n18837;
  assign n25097 = i_RtoB_ACK0 & ~n25096;
  assign n25098 = ~n22729 & ~n25097;
  assign n25099 = ~controllable_DEQ & ~n25098;
  assign n25100 = ~n22725 & ~n25099;
  assign n25101 = i_FULL & ~n25100;
  assign n25102 = ~n22739 & ~n25079;
  assign n25103 = ~controllable_DEQ & ~n25102;
  assign n25104 = ~n22737 & ~n25103;
  assign n25105 = ~i_FULL & ~n25104;
  assign n25106 = ~n25101 & ~n25105;
  assign n25107 = ~i_nEMPTY & ~n25106;
  assign n25108 = ~n25095 & ~n25107;
  assign n25109 = ~controllable_BtoS_ACK0 & ~n25108;
  assign n25110 = ~n25077 & ~n25109;
  assign n25111 = n4465 & ~n25110;
  assign n25112 = ~n22843 & ~n25111;
  assign n25113 = ~i_StoB_REQ10 & ~n25112;
  assign n25114 = ~n22643 & ~n25113;
  assign n25115 = controllable_BtoS_ACK10 & ~n25114;
  assign n25116 = ~n23037 & ~n25113;
  assign n25117 = ~controllable_BtoS_ACK10 & ~n25116;
  assign n25118 = ~n25115 & ~n25117;
  assign n25119 = ~n4464 & ~n25118;
  assign n25120 = ~n25045 & ~n25119;
  assign n25121 = ~n4463 & ~n25120;
  assign n25122 = ~n24945 & ~n25121;
  assign n25123 = n4462 & ~n25122;
  assign n25124 = ~n11147 & ~n14741;
  assign n25125 = i_RtoB_ACK0 & ~n25124;
  assign n25126 = ~n14077 & ~n17545;
  assign n25127 = ~i_RtoB_ACK0 & ~n25126;
  assign n25128 = ~n25125 & ~n25127;
  assign n25129 = controllable_DEQ & ~n25128;
  assign n25130 = ~n11170 & ~n14757;
  assign n25131 = i_RtoB_ACK0 & ~n25130;
  assign n25132 = ~n14086 & ~n17562;
  assign n25133 = ~i_RtoB_ACK0 & ~n25132;
  assign n25134 = ~n25131 & ~n25133;
  assign n25135 = ~controllable_DEQ & ~n25134;
  assign n25136 = ~n25129 & ~n25135;
  assign n25137 = i_nEMPTY & ~n25136;
  assign n25138 = ~n14096 & ~n17581;
  assign n25139 = ~i_RtoB_ACK0 & ~n25138;
  assign n25140 = ~n25125 & ~n25139;
  assign n25141 = ~controllable_DEQ & ~n25140;
  assign n25142 = ~n23063 & ~n25141;
  assign n25143 = i_FULL & ~n25142;
  assign n25144 = ~n14105 & ~n17545;
  assign n25145 = ~i_RtoB_ACK0 & ~n25144;
  assign n25146 = ~n25125 & ~n25145;
  assign n25147 = ~controllable_DEQ & ~n25146;
  assign n25148 = ~n23073 & ~n25147;
  assign n25149 = ~i_FULL & ~n25148;
  assign n25150 = ~n25143 & ~n25149;
  assign n25151 = ~i_nEMPTY & ~n25150;
  assign n25152 = ~n25137 & ~n25151;
  assign n25153 = controllable_BtoS_ACK0 & ~n25152;
  assign n25154 = ~n14120 & ~n14824;
  assign n25155 = ~i_RtoB_ACK0 & ~n25154;
  assign n25156 = ~n24189 & ~n25155;
  assign n25157 = controllable_DEQ & ~n25156;
  assign n25158 = ~n14129 & ~n14841;
  assign n25159 = ~i_RtoB_ACK0 & ~n25158;
  assign n25160 = ~n24195 & ~n25159;
  assign n25161 = ~controllable_DEQ & ~n25160;
  assign n25162 = ~n25157 & ~n25161;
  assign n25163 = i_nEMPTY & ~n25162;
  assign n25164 = ~n14139 & ~n14860;
  assign n25165 = ~i_RtoB_ACK0 & ~n25164;
  assign n25166 = ~n24189 & ~n25165;
  assign n25167 = ~controllable_DEQ & ~n25166;
  assign n25168 = ~n21031 & ~n25167;
  assign n25169 = i_FULL & ~n25168;
  assign n25170 = ~n14147 & ~n14824;
  assign n25171 = ~i_RtoB_ACK0 & ~n25170;
  assign n25172 = ~n24189 & ~n25171;
  assign n25173 = ~controllable_DEQ & ~n25172;
  assign n25174 = ~n21041 & ~n25173;
  assign n25175 = ~i_FULL & ~n25174;
  assign n25176 = ~n25169 & ~n25175;
  assign n25177 = ~i_nEMPTY & ~n25176;
  assign n25178 = ~n25163 & ~n25177;
  assign n25179 = ~controllable_BtoS_ACK0 & ~n25178;
  assign n25180 = ~n25153 & ~n25179;
  assign n25181 = n4465 & ~n25180;
  assign n25182 = ~n24215 & ~n25181;
  assign n25183 = i_StoB_REQ10 & ~n25182;
  assign n25184 = ~n23169 & ~n25183;
  assign n25185 = controllable_BtoS_ACK10 & ~n25184;
  assign n25186 = ~n11395 & ~n17050;
  assign n25187 = i_RtoB_ACK0 & ~n25186;
  assign n25188 = ~n14165 & ~n20366;
  assign n25189 = ~i_RtoB_ACK0 & ~n25188;
  assign n25190 = ~n25187 & ~n25189;
  assign n25191 = controllable_DEQ & ~n25190;
  assign n25192 = ~n11424 & ~n17058;
  assign n25193 = i_RtoB_ACK0 & ~n25192;
  assign n25194 = ~n14171 & ~n20375;
  assign n25195 = ~i_RtoB_ACK0 & ~n25194;
  assign n25196 = ~n25193 & ~n25195;
  assign n25197 = ~controllable_DEQ & ~n25196;
  assign n25198 = ~n25191 & ~n25197;
  assign n25199 = i_FULL & ~n25198;
  assign n25200 = ~n14179 & ~n20386;
  assign n25201 = ~i_RtoB_ACK0 & ~n25200;
  assign n25202 = ~n25187 & ~n25201;
  assign n25203 = controllable_DEQ & ~n25202;
  assign n25204 = ~n14185 & ~n20391;
  assign n25205 = ~i_RtoB_ACK0 & ~n25204;
  assign n25206 = ~n25193 & ~n25205;
  assign n25207 = ~controllable_DEQ & ~n25206;
  assign n25208 = ~n25203 & ~n25207;
  assign n25209 = ~i_FULL & ~n25208;
  assign n25210 = ~n25199 & ~n25209;
  assign n25211 = i_nEMPTY & ~n25210;
  assign n25212 = ~n11395 & ~n17068;
  assign n25213 = i_RtoB_ACK0 & ~n25212;
  assign n25214 = ~n14195 & ~n20409;
  assign n25215 = ~i_RtoB_ACK0 & ~n25214;
  assign n25216 = ~n25213 & ~n25215;
  assign n25217 = ~controllable_DEQ & ~n25216;
  assign n25218 = ~n23205 & ~n25217;
  assign n25219 = i_FULL & ~n25218;
  assign n25220 = ~controllable_DEQ & ~n25190;
  assign n25221 = ~n23217 & ~n25220;
  assign n25222 = ~i_FULL & ~n25221;
  assign n25223 = ~n25219 & ~n25222;
  assign n25224 = ~i_nEMPTY & ~n25223;
  assign n25225 = ~n25211 & ~n25224;
  assign n25226 = controllable_BtoS_ACK0 & ~n25225;
  assign n25227 = ~n11517 & ~n18522;
  assign n25228 = i_RtoB_ACK0 & ~n25227;
  assign n25229 = ~n14210 & ~n20432;
  assign n25230 = ~i_RtoB_ACK0 & ~n25229;
  assign n25231 = ~n25228 & ~n25230;
  assign n25232 = controllable_DEQ & ~n25231;
  assign n25233 = ~n11541 & ~n18530;
  assign n25234 = i_RtoB_ACK0 & ~n25233;
  assign n25235 = ~n14216 & ~n20437;
  assign n25236 = ~i_RtoB_ACK0 & ~n25235;
  assign n25237 = ~n25234 & ~n25236;
  assign n25238 = ~controllable_DEQ & ~n25237;
  assign n25239 = ~n25232 & ~n25238;
  assign n25240 = i_FULL & ~n25239;
  assign n25241 = ~n14224 & ~n20444;
  assign n25242 = ~i_RtoB_ACK0 & ~n25241;
  assign n25243 = ~n25228 & ~n25242;
  assign n25244 = controllable_DEQ & ~n25243;
  assign n25245 = ~n14230 & ~n20449;
  assign n25246 = ~i_RtoB_ACK0 & ~n25245;
  assign n25247 = ~n25234 & ~n25246;
  assign n25248 = ~controllable_DEQ & ~n25247;
  assign n25249 = ~n25244 & ~n25248;
  assign n25250 = ~i_FULL & ~n25249;
  assign n25251 = ~n25240 & ~n25250;
  assign n25252 = i_nEMPTY & ~n25251;
  assign n25253 = ~n11517 & ~n18548;
  assign n25254 = i_RtoB_ACK0 & ~n25253;
  assign n25255 = ~n14240 & ~n20463;
  assign n25256 = ~i_RtoB_ACK0 & ~n25255;
  assign n25257 = ~n25254 & ~n25256;
  assign n25258 = ~controllable_DEQ & ~n25257;
  assign n25259 = ~n23258 & ~n25258;
  assign n25260 = i_FULL & ~n25259;
  assign n25261 = ~controllable_DEQ & ~n25231;
  assign n25262 = ~n23270 & ~n25261;
  assign n25263 = ~i_FULL & ~n25262;
  assign n25264 = ~n25260 & ~n25263;
  assign n25265 = ~i_nEMPTY & ~n25264;
  assign n25266 = ~n25252 & ~n25265;
  assign n25267 = ~controllable_BtoS_ACK0 & ~n25266;
  assign n25268 = ~n25226 & ~n25267;
  assign n25269 = n4465 & ~n25268;
  assign n25270 = ~n24502 & ~n25267;
  assign n25271 = ~n4465 & ~n25270;
  assign n25272 = ~n25269 & ~n25271;
  assign n25273 = i_StoB_REQ10 & ~n25272;
  assign n25274 = ~n11652 & ~n18572;
  assign n25275 = i_RtoB_ACK0 & ~n25274;
  assign n25276 = ~n14261 & ~n17974;
  assign n25277 = ~i_RtoB_ACK0 & ~n25276;
  assign n25278 = ~n25275 & ~n25277;
  assign n25279 = controllable_DEQ & ~n25278;
  assign n25280 = ~n11681 & ~n18580;
  assign n25281 = i_RtoB_ACK0 & ~n25280;
  assign n25282 = ~n14267 & ~n17993;
  assign n25283 = ~i_RtoB_ACK0 & ~n25282;
  assign n25284 = ~n25281 & ~n25283;
  assign n25285 = ~controllable_DEQ & ~n25284;
  assign n25286 = ~n25279 & ~n25285;
  assign n25287 = i_FULL & ~n25286;
  assign n25288 = ~n14275 & ~n18012;
  assign n25289 = ~i_RtoB_ACK0 & ~n25288;
  assign n25290 = ~n25275 & ~n25289;
  assign n25291 = controllable_DEQ & ~n25290;
  assign n25292 = ~n14281 & ~n18028;
  assign n25293 = ~i_RtoB_ACK0 & ~n25292;
  assign n25294 = ~n25281 & ~n25293;
  assign n25295 = ~controllable_DEQ & ~n25294;
  assign n25296 = ~n25291 & ~n25295;
  assign n25297 = ~i_FULL & ~n25296;
  assign n25298 = ~n25287 & ~n25297;
  assign n25299 = i_nEMPTY & ~n25298;
  assign n25300 = ~n11652 & ~n18598;
  assign n25301 = i_RtoB_ACK0 & ~n25300;
  assign n25302 = ~n14291 & ~n18065;
  assign n25303 = ~i_RtoB_ACK0 & ~n25302;
  assign n25304 = ~n25301 & ~n25303;
  assign n25305 = ~controllable_DEQ & ~n25304;
  assign n25306 = ~n23317 & ~n25305;
  assign n25307 = i_FULL & ~n25306;
  assign n25308 = ~n14299 & ~n17974;
  assign n25309 = ~i_RtoB_ACK0 & ~n25308;
  assign n25310 = ~n25275 & ~n25309;
  assign n25311 = ~controllable_DEQ & ~n25310;
  assign n25312 = ~n23329 & ~n25311;
  assign n25313 = ~i_FULL & ~n25312;
  assign n25314 = ~n25307 & ~n25313;
  assign n25315 = ~i_nEMPTY & ~n25314;
  assign n25316 = ~n25299 & ~n25315;
  assign n25317 = controllable_BtoS_ACK0 & ~n25316;
  assign n25318 = ~n11799 & ~n18617;
  assign n25319 = i_RtoB_ACK0 & ~n25318;
  assign n25320 = ~n14311 & ~n18116;
  assign n25321 = ~i_RtoB_ACK0 & ~n25320;
  assign n25322 = ~n25319 & ~n25321;
  assign n25323 = controllable_DEQ & ~n25322;
  assign n25324 = ~n11828 & ~n18625;
  assign n25325 = i_RtoB_ACK0 & ~n25324;
  assign n25326 = ~n14317 & ~n18135;
  assign n25327 = ~i_RtoB_ACK0 & ~n25326;
  assign n25328 = ~n25325 & ~n25327;
  assign n25329 = ~controllable_DEQ & ~n25328;
  assign n25330 = ~n25323 & ~n25329;
  assign n25331 = i_FULL & ~n25330;
  assign n25332 = ~n14325 & ~n18154;
  assign n25333 = ~i_RtoB_ACK0 & ~n25332;
  assign n25334 = ~n25319 & ~n25333;
  assign n25335 = controllable_DEQ & ~n25334;
  assign n25336 = ~n14331 & ~n18170;
  assign n25337 = ~i_RtoB_ACK0 & ~n25336;
  assign n25338 = ~n25325 & ~n25337;
  assign n25339 = ~controllable_DEQ & ~n25338;
  assign n25340 = ~n25335 & ~n25339;
  assign n25341 = ~i_FULL & ~n25340;
  assign n25342 = ~n25331 & ~n25341;
  assign n25343 = i_nEMPTY & ~n25342;
  assign n25344 = ~n11799 & ~n18643;
  assign n25345 = i_RtoB_ACK0 & ~n25344;
  assign n25346 = ~n14341 & ~n18207;
  assign n25347 = ~i_RtoB_ACK0 & ~n25346;
  assign n25348 = ~n25345 & ~n25347;
  assign n25349 = ~controllable_DEQ & ~n25348;
  assign n25350 = ~n23373 & ~n25349;
  assign n25351 = i_FULL & ~n25350;
  assign n25352 = ~n14349 & ~n18116;
  assign n25353 = ~i_RtoB_ACK0 & ~n25352;
  assign n25354 = ~n25319 & ~n25353;
  assign n25355 = ~controllable_DEQ & ~n25354;
  assign n25356 = ~n23385 & ~n25355;
  assign n25357 = ~i_FULL & ~n25356;
  assign n25358 = ~n25351 & ~n25357;
  assign n25359 = ~i_nEMPTY & ~n25358;
  assign n25360 = ~n25343 & ~n25359;
  assign n25361 = ~controllable_BtoS_ACK0 & ~n25360;
  assign n25362 = ~n25317 & ~n25361;
  assign n25363 = n4465 & ~n25362;
  assign n25364 = ~n14363 & ~n15190;
  assign n25365 = ~i_RtoB_ACK0 & ~n25364;
  assign n25366 = ~n24309 & ~n25365;
  assign n25367 = controllable_DEQ & ~n25366;
  assign n25368 = ~n13572 & ~n15209;
  assign n25369 = ~i_RtoB_ACK0 & ~n25368;
  assign n25370 = ~n24315 & ~n25369;
  assign n25371 = ~controllable_DEQ & ~n25370;
  assign n25372 = ~n25367 & ~n25371;
  assign n25373 = i_nEMPTY & ~n25372;
  assign n25374 = ~n13580 & ~n15237;
  assign n25375 = ~i_RtoB_ACK0 & ~n25374;
  assign n25376 = ~n24323 & ~n25375;
  assign n25377 = ~controllable_DEQ & ~n25376;
  assign n25378 = ~n21187 & ~n25377;
  assign n25379 = i_FULL & ~n25378;
  assign n25380 = ~n14377 & ~n15190;
  assign n25381 = ~i_RtoB_ACK0 & ~n25380;
  assign n25382 = ~n24309 & ~n25381;
  assign n25383 = ~controllable_DEQ & ~n25382;
  assign n25384 = ~n21199 & ~n25383;
  assign n25385 = ~i_FULL & ~n25384;
  assign n25386 = ~n25379 & ~n25385;
  assign n25387 = ~i_nEMPTY & ~n25386;
  assign n25388 = ~n25373 & ~n25387;
  assign n25389 = controllable_BtoS_ACK0 & ~n25388;
  assign n25390 = ~n24383 & ~n25389;
  assign n25391 = ~n4465 & ~n25390;
  assign n25392 = ~n25363 & ~n25391;
  assign n25393 = ~i_StoB_REQ10 & ~n25392;
  assign n25394 = ~n25273 & ~n25393;
  assign n25395 = ~controllable_BtoS_ACK10 & ~n25394;
  assign n25396 = ~n25185 & ~n25395;
  assign n25397 = n4464 & ~n25396;
  assign n25398 = ~n23169 & ~n24609;
  assign n25399 = controllable_BtoS_ACK10 & ~n25398;
  assign n25400 = ~n11936 & ~n17050;
  assign n25401 = i_RtoB_ACK0 & ~n25400;
  assign n25402 = ~n14399 & ~n20680;
  assign n25403 = ~i_RtoB_ACK0 & ~n25402;
  assign n25404 = ~n25401 & ~n25403;
  assign n25405 = controllable_DEQ & ~n25404;
  assign n25406 = ~n11960 & ~n17058;
  assign n25407 = i_RtoB_ACK0 & ~n25406;
  assign n25408 = ~n14405 & ~n20685;
  assign n25409 = ~i_RtoB_ACK0 & ~n25408;
  assign n25410 = ~n25407 & ~n25409;
  assign n25411 = ~controllable_DEQ & ~n25410;
  assign n25412 = ~n25405 & ~n25411;
  assign n25413 = i_FULL & ~n25412;
  assign n25414 = ~n14413 & ~n20692;
  assign n25415 = ~i_RtoB_ACK0 & ~n25414;
  assign n25416 = ~n25401 & ~n25415;
  assign n25417 = controllable_DEQ & ~n25416;
  assign n25418 = ~n14419 & ~n20697;
  assign n25419 = ~i_RtoB_ACK0 & ~n25418;
  assign n25420 = ~n25407 & ~n25419;
  assign n25421 = ~controllable_DEQ & ~n25420;
  assign n25422 = ~n25417 & ~n25421;
  assign n25423 = ~i_FULL & ~n25422;
  assign n25424 = ~n25413 & ~n25423;
  assign n25425 = i_nEMPTY & ~n25424;
  assign n25426 = ~n11936 & ~n17068;
  assign n25427 = i_RtoB_ACK0 & ~n25426;
  assign n25428 = ~n14429 & ~n20711;
  assign n25429 = ~i_RtoB_ACK0 & ~n25428;
  assign n25430 = ~n25427 & ~n25429;
  assign n25431 = ~controllable_DEQ & ~n25430;
  assign n25432 = ~n23439 & ~n25431;
  assign n25433 = i_FULL & ~n25432;
  assign n25434 = ~controllable_DEQ & ~n25404;
  assign n25435 = ~n23451 & ~n25434;
  assign n25436 = ~i_FULL & ~n25435;
  assign n25437 = ~n25433 & ~n25436;
  assign n25438 = ~i_nEMPTY & ~n25437;
  assign n25439 = ~n25425 & ~n25438;
  assign n25440 = controllable_BtoS_ACK0 & ~n25439;
  assign n25441 = ~n12044 & ~n18522;
  assign n25442 = i_RtoB_ACK0 & ~n25441;
  assign n25443 = ~n14444 & ~n20730;
  assign n25444 = ~i_RtoB_ACK0 & ~n25443;
  assign n25445 = ~n25442 & ~n25444;
  assign n25446 = controllable_DEQ & ~n25445;
  assign n25447 = ~n12068 & ~n18530;
  assign n25448 = i_RtoB_ACK0 & ~n25447;
  assign n25449 = ~n14450 & ~n20735;
  assign n25450 = ~i_RtoB_ACK0 & ~n25449;
  assign n25451 = ~n25448 & ~n25450;
  assign n25452 = ~controllable_DEQ & ~n25451;
  assign n25453 = ~n25446 & ~n25452;
  assign n25454 = i_FULL & ~n25453;
  assign n25455 = ~n14458 & ~n20742;
  assign n25456 = ~i_RtoB_ACK0 & ~n25455;
  assign n25457 = ~n25442 & ~n25456;
  assign n25458 = controllable_DEQ & ~n25457;
  assign n25459 = ~n14464 & ~n20747;
  assign n25460 = ~i_RtoB_ACK0 & ~n25459;
  assign n25461 = ~n25448 & ~n25460;
  assign n25462 = ~controllable_DEQ & ~n25461;
  assign n25463 = ~n25458 & ~n25462;
  assign n25464 = ~i_FULL & ~n25463;
  assign n25465 = ~n25454 & ~n25464;
  assign n25466 = i_nEMPTY & ~n25465;
  assign n25467 = ~n12044 & ~n18548;
  assign n25468 = i_RtoB_ACK0 & ~n25467;
  assign n25469 = ~n14474 & ~n20761;
  assign n25470 = ~i_RtoB_ACK0 & ~n25469;
  assign n25471 = ~n25468 & ~n25470;
  assign n25472 = ~controllable_DEQ & ~n25471;
  assign n25473 = ~n23492 & ~n25472;
  assign n25474 = i_FULL & ~n25473;
  assign n25475 = ~controllable_DEQ & ~n25445;
  assign n25476 = ~n23504 & ~n25475;
  assign n25477 = ~i_FULL & ~n25476;
  assign n25478 = ~n25474 & ~n25477;
  assign n25479 = ~i_nEMPTY & ~n25478;
  assign n25480 = ~n25466 & ~n25479;
  assign n25481 = ~controllable_BtoS_ACK0 & ~n25480;
  assign n25482 = ~n25440 & ~n25481;
  assign n25483 = n4465 & ~n25482;
  assign n25484 = ~n24894 & ~n25481;
  assign n25485 = ~n4465 & ~n25484;
  assign n25486 = ~n25483 & ~n25485;
  assign n25487 = i_StoB_REQ10 & ~n25486;
  assign n25488 = ~n14495 & ~n15889;
  assign n25489 = ~i_RtoB_ACK0 & ~n25488;
  assign n25490 = ~n24611 & ~n25489;
  assign n25491 = controllable_DEQ & ~n25490;
  assign n25492 = ~n13922 & ~n15908;
  assign n25493 = ~i_RtoB_ACK0 & ~n25492;
  assign n25494 = ~n24617 & ~n25493;
  assign n25495 = ~controllable_DEQ & ~n25494;
  assign n25496 = ~n25491 & ~n25495;
  assign n25497 = i_FULL & ~n25496;
  assign n25498 = ~n14505 & ~n15927;
  assign n25499 = ~i_RtoB_ACK0 & ~n25498;
  assign n25500 = ~n24611 & ~n25499;
  assign n25501 = controllable_DEQ & ~n25500;
  assign n25502 = ~n13936 & ~n15943;
  assign n25503 = ~i_RtoB_ACK0 & ~n25502;
  assign n25504 = ~n24617 & ~n25503;
  assign n25505 = ~controllable_DEQ & ~n25504;
  assign n25506 = ~n25501 & ~n25505;
  assign n25507 = ~i_FULL & ~n25506;
  assign n25508 = ~n25497 & ~n25507;
  assign n25509 = i_nEMPTY & ~n25508;
  assign n25510 = ~n13946 & ~n15980;
  assign n25511 = ~i_RtoB_ACK0 & ~n25510;
  assign n25512 = ~n24637 & ~n25511;
  assign n25513 = ~controllable_DEQ & ~n25512;
  assign n25514 = ~n21593 & ~n25513;
  assign n25515 = i_FULL & ~n25514;
  assign n25516 = ~n14521 & ~n15889;
  assign n25517 = ~i_RtoB_ACK0 & ~n25516;
  assign n25518 = ~n24611 & ~n25517;
  assign n25519 = ~controllable_DEQ & ~n25518;
  assign n25520 = ~n21605 & ~n25519;
  assign n25521 = ~i_FULL & ~n25520;
  assign n25522 = ~n25515 & ~n25521;
  assign n25523 = ~i_nEMPTY & ~n25522;
  assign n25524 = ~n25509 & ~n25523;
  assign n25525 = controllable_BtoS_ACK0 & ~n25524;
  assign n25526 = ~n14533 & ~n16031;
  assign n25527 = ~i_RtoB_ACK0 & ~n25526;
  assign n25528 = ~n24655 & ~n25527;
  assign n25529 = controllable_DEQ & ~n25528;
  assign n25530 = ~n13967 & ~n16050;
  assign n25531 = ~i_RtoB_ACK0 & ~n25530;
  assign n25532 = ~n24661 & ~n25531;
  assign n25533 = ~controllable_DEQ & ~n25532;
  assign n25534 = ~n25529 & ~n25533;
  assign n25535 = i_FULL & ~n25534;
  assign n25536 = ~n14543 & ~n16069;
  assign n25537 = ~i_RtoB_ACK0 & ~n25536;
  assign n25538 = ~n24655 & ~n25537;
  assign n25539 = controllable_DEQ & ~n25538;
  assign n25540 = ~n13981 & ~n16085;
  assign n25541 = ~i_RtoB_ACK0 & ~n25540;
  assign n25542 = ~n24661 & ~n25541;
  assign n25543 = ~controllable_DEQ & ~n25542;
  assign n25544 = ~n25539 & ~n25543;
  assign n25545 = ~i_FULL & ~n25544;
  assign n25546 = ~n25535 & ~n25545;
  assign n25547 = i_nEMPTY & ~n25546;
  assign n25548 = ~n13991 & ~n16122;
  assign n25549 = ~i_RtoB_ACK0 & ~n25548;
  assign n25550 = ~n24681 & ~n25549;
  assign n25551 = ~controllable_DEQ & ~n25550;
  assign n25552 = ~n21649 & ~n25551;
  assign n25553 = i_FULL & ~n25552;
  assign n25554 = ~n14559 & ~n16031;
  assign n25555 = ~i_RtoB_ACK0 & ~n25554;
  assign n25556 = ~n24655 & ~n25555;
  assign n25557 = ~controllable_DEQ & ~n25556;
  assign n25558 = ~n21661 & ~n25557;
  assign n25559 = ~i_FULL & ~n25558;
  assign n25560 = ~n25553 & ~n25559;
  assign n25561 = ~i_nEMPTY & ~n25560;
  assign n25562 = ~n25547 & ~n25561;
  assign n25563 = ~controllable_BtoS_ACK0 & ~n25562;
  assign n25564 = ~n25525 & ~n25563;
  assign n25565 = n4465 & ~n25564;
  assign n25566 = ~n24777 & ~n25565;
  assign n25567 = ~i_StoB_REQ10 & ~n25566;
  assign n25568 = ~n25487 & ~n25567;
  assign n25569 = ~controllable_BtoS_ACK10 & ~n25568;
  assign n25570 = ~n25399 & ~n25569;
  assign n25571 = ~n4464 & ~n25570;
  assign n25572 = ~n25397 & ~n25571;
  assign n25573 = n4463 & ~n25572;
  assign n25574 = ~n12168 & ~n14741;
  assign n25575 = i_RtoB_ACK0 & ~n25574;
  assign n25576 = ~n23527 & ~n25575;
  assign n25577 = controllable_DEQ & ~n25576;
  assign n25578 = ~n12189 & ~n14757;
  assign n25579 = i_RtoB_ACK0 & ~n25578;
  assign n25580 = ~n23533 & ~n25579;
  assign n25581 = ~controllable_DEQ & ~n25580;
  assign n25582 = ~n25577 & ~n25581;
  assign n25583 = i_nEMPTY & ~n25582;
  assign n25584 = ~n23543 & ~n25575;
  assign n25585 = ~controllable_DEQ & ~n25584;
  assign n25586 = ~n23541 & ~n25585;
  assign n25587 = i_FULL & ~n25586;
  assign n25588 = ~n23553 & ~n25575;
  assign n25589 = ~controllable_DEQ & ~n25588;
  assign n25590 = ~n23551 & ~n25589;
  assign n25591 = ~i_FULL & ~n25590;
  assign n25592 = ~n25587 & ~n25591;
  assign n25593 = ~i_nEMPTY & ~n25592;
  assign n25594 = ~n25583 & ~n25593;
  assign n25595 = controllable_BtoS_ACK0 & ~n25594;
  assign n25596 = ~n12261 & ~n16723;
  assign n25597 = i_RtoB_ACK0 & ~n25596;
  assign n25598 = ~n23565 & ~n25597;
  assign n25599 = controllable_DEQ & ~n25598;
  assign n25600 = ~n12279 & ~n16729;
  assign n25601 = i_RtoB_ACK0 & ~n25600;
  assign n25602 = ~n23571 & ~n25601;
  assign n25603 = ~controllable_DEQ & ~n25602;
  assign n25604 = ~n25599 & ~n25603;
  assign n25605 = i_nEMPTY & ~n25604;
  assign n25606 = ~n23581 & ~n25597;
  assign n25607 = ~controllable_DEQ & ~n25606;
  assign n25608 = ~n23579 & ~n25607;
  assign n25609 = i_FULL & ~n25608;
  assign n25610 = ~n23591 & ~n25597;
  assign n25611 = ~controllable_DEQ & ~n25610;
  assign n25612 = ~n23589 & ~n25611;
  assign n25613 = ~i_FULL & ~n25612;
  assign n25614 = ~n25609 & ~n25613;
  assign n25615 = ~i_nEMPTY & ~n25614;
  assign n25616 = ~n25605 & ~n25615;
  assign n25617 = ~controllable_BtoS_ACK0 & ~n25616;
  assign n25618 = ~n25595 & ~n25617;
  assign n25619 = n4465 & ~n25618;
  assign n25620 = ~n23619 & ~n25619;
  assign n25621 = i_StoB_REQ10 & ~n25620;
  assign n25622 = ~n23169 & ~n25621;
  assign n25623 = controllable_BtoS_ACK10 & ~n25622;
  assign n25624 = ~n23873 & ~n25623;
  assign n25625 = n4464 & ~n25624;
  assign n25626 = ~n24127 & ~n25625;
  assign n25627 = ~n4463 & ~n25626;
  assign n25628 = ~n25573 & ~n25627;
  assign n25629 = ~n4462 & ~n25628;
  assign n25630 = ~n25123 & ~n25629;
  assign n25631 = ~n4461 & ~n25630;
  assign n25632 = ~n24133 & ~n25631;
  assign n25633 = ~n4459 & ~n25632;
  assign n25634 = ~n6583 & ~n16780;
  assign n25635 = i_RtoB_ACK0 & ~n25634;
  assign n25636 = ~n6778 & ~n9306;
  assign n25637 = ~controllable_BtoR_REQ0 & ~n25636;
  assign n25638 = ~n14904 & ~n25637;
  assign n25639 = ~i_RtoB_ACK0 & ~n25638;
  assign n25640 = ~n25635 & ~n25639;
  assign n25641 = controllable_DEQ & ~n25640;
  assign n25642 = ~n6791 & ~n16788;
  assign n25643 = i_RtoB_ACK0 & ~n25642;
  assign n25644 = ~n13480 & ~n14923;
  assign n25645 = ~i_RtoB_ACK0 & ~n25644;
  assign n25646 = ~n25643 & ~n25645;
  assign n25647 = ~controllable_DEQ & ~n25646;
  assign n25648 = ~n25641 & ~n25647;
  assign n25649 = i_FULL & ~n25648;
  assign n25650 = ~n6815 & ~n9532;
  assign n25651 = ~controllable_BtoR_REQ0 & ~n25650;
  assign n25652 = ~n14942 & ~n25651;
  assign n25653 = ~i_RtoB_ACK0 & ~n25652;
  assign n25654 = ~n25635 & ~n25653;
  assign n25655 = controllable_DEQ & ~n25654;
  assign n25656 = ~n13494 & ~n14958;
  assign n25657 = ~i_RtoB_ACK0 & ~n25656;
  assign n25658 = ~n25643 & ~n25657;
  assign n25659 = ~controllable_DEQ & ~n25658;
  assign n25660 = ~n25655 & ~n25659;
  assign n25661 = ~i_FULL & ~n25660;
  assign n25662 = ~n25649 & ~n25661;
  assign n25663 = i_nEMPTY & ~n25662;
  assign n25664 = ~n6583 & ~n16806;
  assign n25665 = i_RtoB_ACK0 & ~n25664;
  assign n25666 = ~n13504 & ~n14995;
  assign n25667 = ~i_RtoB_ACK0 & ~n25666;
  assign n25668 = ~n25665 & ~n25667;
  assign n25669 = ~controllable_DEQ & ~n25668;
  assign n25670 = ~n21089 & ~n25669;
  assign n25671 = i_FULL & ~n25670;
  assign n25672 = ~n6873 & ~n9306;
  assign n25673 = ~controllable_BtoR_REQ0 & ~n25672;
  assign n25674 = ~n14904 & ~n25673;
  assign n25675 = ~i_RtoB_ACK0 & ~n25674;
  assign n25676 = ~n25635 & ~n25675;
  assign n25677 = ~controllable_DEQ & ~n25676;
  assign n25678 = ~n21101 & ~n25677;
  assign n25679 = ~i_FULL & ~n25678;
  assign n25680 = ~n25671 & ~n25679;
  assign n25681 = ~i_nEMPTY & ~n25680;
  assign n25682 = ~n25663 & ~n25681;
  assign n25683 = controllable_BtoS_ACK0 & ~n25682;
  assign n25684 = ~n6922 & ~n16825;
  assign n25685 = i_RtoB_ACK0 & ~n25684;
  assign n25686 = ~n6944 & ~n9639;
  assign n25687 = ~controllable_BtoR_REQ0 & ~n25686;
  assign n25688 = ~n15046 & ~n25687;
  assign n25689 = ~i_RtoB_ACK0 & ~n25688;
  assign n25690 = ~n25685 & ~n25689;
  assign n25691 = controllable_DEQ & ~n25690;
  assign n25692 = ~n6957 & ~n16833;
  assign n25693 = i_RtoB_ACK0 & ~n25692;
  assign n25694 = ~n13525 & ~n15065;
  assign n25695 = ~i_RtoB_ACK0 & ~n25694;
  assign n25696 = ~n25693 & ~n25695;
  assign n25697 = ~controllable_DEQ & ~n25696;
  assign n25698 = ~n25691 & ~n25697;
  assign n25699 = i_FULL & ~n25698;
  assign n25700 = ~n6981 & ~n9679;
  assign n25701 = ~controllable_BtoR_REQ0 & ~n25700;
  assign n25702 = ~n15084 & ~n25701;
  assign n25703 = ~i_RtoB_ACK0 & ~n25702;
  assign n25704 = ~n25685 & ~n25703;
  assign n25705 = controllable_DEQ & ~n25704;
  assign n25706 = ~n13539 & ~n15100;
  assign n25707 = ~i_RtoB_ACK0 & ~n25706;
  assign n25708 = ~n25693 & ~n25707;
  assign n25709 = ~controllable_DEQ & ~n25708;
  assign n25710 = ~n25705 & ~n25709;
  assign n25711 = ~i_FULL & ~n25710;
  assign n25712 = ~n25699 & ~n25711;
  assign n25713 = i_nEMPTY & ~n25712;
  assign n25714 = ~n6922 & ~n16851;
  assign n25715 = i_RtoB_ACK0 & ~n25714;
  assign n25716 = ~n13549 & ~n15137;
  assign n25717 = ~i_RtoB_ACK0 & ~n25716;
  assign n25718 = ~n25715 & ~n25717;
  assign n25719 = ~controllable_DEQ & ~n25718;
  assign n25720 = ~n21145 & ~n25719;
  assign n25721 = i_FULL & ~n25720;
  assign n25722 = ~n7039 & ~n9639;
  assign n25723 = ~controllable_BtoR_REQ0 & ~n25722;
  assign n25724 = ~n15046 & ~n25723;
  assign n25725 = ~i_RtoB_ACK0 & ~n25724;
  assign n25726 = ~n25685 & ~n25725;
  assign n25727 = ~controllable_DEQ & ~n25726;
  assign n25728 = ~n21157 & ~n25727;
  assign n25729 = ~i_FULL & ~n25728;
  assign n25730 = ~n25721 & ~n25729;
  assign n25731 = ~i_nEMPTY & ~n25730;
  assign n25732 = ~n25713 & ~n25731;
  assign n25733 = ~controllable_BtoS_ACK0 & ~n25732;
  assign n25734 = ~n25683 & ~n25733;
  assign n25735 = n4465 & ~n25734;
  assign n25736 = ~n7091 & ~n16872;
  assign n25737 = i_RtoB_ACK0 & ~n25736;
  assign n25738 = ~n25365 & ~n25737;
  assign n25739 = controllable_DEQ & ~n25738;
  assign n25740 = ~n7117 & ~n16880;
  assign n25741 = i_RtoB_ACK0 & ~n25740;
  assign n25742 = ~n25369 & ~n25741;
  assign n25743 = ~controllable_DEQ & ~n25742;
  assign n25744 = ~n25739 & ~n25743;
  assign n25745 = i_nEMPTY & ~n25744;
  assign n25746 = ~n7091 & ~n16890;
  assign n25747 = i_RtoB_ACK0 & ~n25746;
  assign n25748 = ~n25375 & ~n25747;
  assign n25749 = ~controllable_DEQ & ~n25748;
  assign n25750 = ~n21187 & ~n25749;
  assign n25751 = i_FULL & ~n25750;
  assign n25752 = ~n25381 & ~n25737;
  assign n25753 = ~controllable_DEQ & ~n25752;
  assign n25754 = ~n21199 & ~n25753;
  assign n25755 = ~i_FULL & ~n25754;
  assign n25756 = ~n25751 & ~n25755;
  assign n25757 = ~i_nEMPTY & ~n25756;
  assign n25758 = ~n25745 & ~n25757;
  assign n25759 = controllable_BtoS_ACK0 & ~n25758;
  assign n25760 = ~n24383 & ~n25759;
  assign n25761 = ~n4465 & ~n25760;
  assign n25762 = ~n25735 & ~n25761;
  assign n25763 = ~i_StoB_REQ10 & ~n25762;
  assign n25764 = ~n24217 & ~n25763;
  assign n25765 = controllable_BtoS_ACK10 & ~n25764;
  assign n25766 = ~n24547 & ~n25763;
  assign n25767 = ~controllable_BtoS_ACK10 & ~n25766;
  assign n25768 = ~n25765 & ~n25767;
  assign n25769 = n4464 & ~n25768;
  assign n25770 = ~n7919 & ~n17188;
  assign n25771 = i_RtoB_ACK0 & ~n25770;
  assign n25772 = ~n25489 & ~n25771;
  assign n25773 = controllable_DEQ & ~n25772;
  assign n25774 = ~n7953 & ~n17196;
  assign n25775 = i_RtoB_ACK0 & ~n25774;
  assign n25776 = ~n25493 & ~n25775;
  assign n25777 = ~controllable_DEQ & ~n25776;
  assign n25778 = ~n25773 & ~n25777;
  assign n25779 = i_FULL & ~n25778;
  assign n25780 = ~n25499 & ~n25771;
  assign n25781 = controllable_DEQ & ~n25780;
  assign n25782 = ~n25503 & ~n25775;
  assign n25783 = ~controllable_DEQ & ~n25782;
  assign n25784 = ~n25781 & ~n25783;
  assign n25785 = ~i_FULL & ~n25784;
  assign n25786 = ~n25779 & ~n25785;
  assign n25787 = i_nEMPTY & ~n25786;
  assign n25788 = ~n7919 & ~n17214;
  assign n25789 = i_RtoB_ACK0 & ~n25788;
  assign n25790 = ~n25511 & ~n25789;
  assign n25791 = ~controllable_DEQ & ~n25790;
  assign n25792 = ~n21593 & ~n25791;
  assign n25793 = i_FULL & ~n25792;
  assign n25794 = ~n25517 & ~n25771;
  assign n25795 = ~controllable_DEQ & ~n25794;
  assign n25796 = ~n21605 & ~n25795;
  assign n25797 = ~i_FULL & ~n25796;
  assign n25798 = ~n25793 & ~n25797;
  assign n25799 = ~i_nEMPTY & ~n25798;
  assign n25800 = ~n25787 & ~n25799;
  assign n25801 = controllable_BtoS_ACK0 & ~n25800;
  assign n25802 = ~n8086 & ~n17233;
  assign n25803 = i_RtoB_ACK0 & ~n25802;
  assign n25804 = ~n25527 & ~n25803;
  assign n25805 = controllable_DEQ & ~n25804;
  assign n25806 = ~n8117 & ~n17241;
  assign n25807 = i_RtoB_ACK0 & ~n25806;
  assign n25808 = ~n25531 & ~n25807;
  assign n25809 = ~controllable_DEQ & ~n25808;
  assign n25810 = ~n25805 & ~n25809;
  assign n25811 = i_FULL & ~n25810;
  assign n25812 = ~n25537 & ~n25803;
  assign n25813 = controllable_DEQ & ~n25812;
  assign n25814 = ~n25541 & ~n25807;
  assign n25815 = ~controllable_DEQ & ~n25814;
  assign n25816 = ~n25813 & ~n25815;
  assign n25817 = ~i_FULL & ~n25816;
  assign n25818 = ~n25811 & ~n25817;
  assign n25819 = i_nEMPTY & ~n25818;
  assign n25820 = ~n8086 & ~n17259;
  assign n25821 = i_RtoB_ACK0 & ~n25820;
  assign n25822 = ~n25549 & ~n25821;
  assign n25823 = ~controllable_DEQ & ~n25822;
  assign n25824 = ~n21649 & ~n25823;
  assign n25825 = i_FULL & ~n25824;
  assign n25826 = ~n25555 & ~n25803;
  assign n25827 = ~controllable_DEQ & ~n25826;
  assign n25828 = ~n21661 & ~n25827;
  assign n25829 = ~i_FULL & ~n25828;
  assign n25830 = ~n25825 & ~n25829;
  assign n25831 = ~i_nEMPTY & ~n25830;
  assign n25832 = ~n25819 & ~n25831;
  assign n25833 = ~controllable_BtoS_ACK0 & ~n25832;
  assign n25834 = ~n25801 & ~n25833;
  assign n25835 = n4465 & ~n25834;
  assign n25836 = ~n24777 & ~n25835;
  assign n25837 = ~i_StoB_REQ10 & ~n25836;
  assign n25838 = ~n24609 & ~n25837;
  assign n25839 = controllable_BtoS_ACK10 & ~n25838;
  assign n25840 = ~n24939 & ~n25837;
  assign n25841 = ~controllable_BtoS_ACK10 & ~n25840;
  assign n25842 = ~n25839 & ~n25841;
  assign n25843 = ~n4464 & ~n25842;
  assign n25844 = ~n25769 & ~n25843;
  assign n25845 = ~n4463 & ~n25844;
  assign n25846 = ~n21983 & ~n25845;
  assign n25847 = n4462 & ~n25846;
  assign n25848 = ~n11147 & ~n18428;
  assign n25849 = i_RtoB_ACK0 & ~n25848;
  assign n25850 = ~n11158 & ~n12172;
  assign n25851 = ~controllable_BtoR_REQ0 & ~n25850;
  assign n25852 = ~n17545 & ~n25851;
  assign n25853 = ~i_RtoB_ACK0 & ~n25852;
  assign n25854 = ~n25849 & ~n25853;
  assign n25855 = controllable_DEQ & ~n25854;
  assign n25856 = ~n11170 & ~n18434;
  assign n25857 = i_RtoB_ACK0 & ~n25856;
  assign n25858 = ~n11168 & ~n12193;
  assign n25859 = ~controllable_BtoR_REQ0 & ~n25858;
  assign n25860 = ~n17562 & ~n25859;
  assign n25861 = ~i_RtoB_ACK0 & ~n25860;
  assign n25862 = ~n25857 & ~n25861;
  assign n25863 = ~controllable_DEQ & ~n25862;
  assign n25864 = ~n25855 & ~n25863;
  assign n25865 = i_nEMPTY & ~n25864;
  assign n25866 = ~n11145 & ~n12216;
  assign n25867 = ~controllable_BtoR_REQ0 & ~n25866;
  assign n25868 = ~n17581 & ~n25867;
  assign n25869 = ~i_RtoB_ACK0 & ~n25868;
  assign n25870 = ~n25849 & ~n25869;
  assign n25871 = ~controllable_DEQ & ~n25870;
  assign n25872 = ~n23063 & ~n25871;
  assign n25873 = i_FULL & ~n25872;
  assign n25874 = ~n12172 & ~n14103;
  assign n25875 = ~controllable_BtoR_REQ0 & ~n25874;
  assign n25876 = ~n17545 & ~n25875;
  assign n25877 = ~i_RtoB_ACK0 & ~n25876;
  assign n25878 = ~n25849 & ~n25877;
  assign n25879 = ~controllable_DEQ & ~n25878;
  assign n25880 = ~n23073 & ~n25879;
  assign n25881 = ~i_FULL & ~n25880;
  assign n25882 = ~n25873 & ~n25881;
  assign n25883 = ~i_nEMPTY & ~n25882;
  assign n25884 = ~n25865 & ~n25883;
  assign n25885 = controllable_BtoS_ACK0 & ~n25884;
  assign n25886 = ~n5340 & ~n18456;
  assign n25887 = i_RtoB_ACK0 & ~n25886;
  assign n25888 = ~n24191 & ~n25887;
  assign n25889 = controllable_DEQ & ~n25888;
  assign n25890 = ~n5363 & ~n18462;
  assign n25891 = i_RtoB_ACK0 & ~n25890;
  assign n25892 = ~n22095 & ~n25891;
  assign n25893 = ~controllable_DEQ & ~n25892;
  assign n25894 = ~n25889 & ~n25893;
  assign n25895 = i_nEMPTY & ~n25894;
  assign n25896 = ~n22117 & ~n25887;
  assign n25897 = ~controllable_DEQ & ~n25896;
  assign n25898 = ~n21031 & ~n25897;
  assign n25899 = i_FULL & ~n25898;
  assign n25900 = ~n24205 & ~n25887;
  assign n25901 = ~controllable_DEQ & ~n25900;
  assign n25902 = ~n21041 & ~n25901;
  assign n25903 = ~i_FULL & ~n25902;
  assign n25904 = ~n25899 & ~n25903;
  assign n25905 = ~i_nEMPTY & ~n25904;
  assign n25906 = ~n25895 & ~n25905;
  assign n25907 = ~controllable_BtoS_ACK0 & ~n25906;
  assign n25908 = ~n25885 & ~n25907;
  assign n25909 = n4465 & ~n25908;
  assign n25910 = ~n24215 & ~n25909;
  assign n25911 = i_StoB_REQ10 & ~n25910;
  assign n25912 = ~n23169 & ~n25911;
  assign n25913 = controllable_BtoS_ACK10 & ~n25912;
  assign n25914 = ~n25395 & ~n25913;
  assign n25915 = n4464 & ~n25914;
  assign n25916 = ~n25571 & ~n25915;
  assign n25917 = ~n4463 & ~n25916;
  assign n25918 = ~n23523 & ~n25917;
  assign n25919 = ~n4462 & ~n25918;
  assign n25920 = ~n25847 & ~n25919;
  assign n25921 = n4461 & ~n25920;
  assign n25922 = ~n8763 & ~n18867;
  assign n25923 = ~controllable_BtoR_REQ0 & ~n25922;
  assign n25924 = ~n14598 & ~n25923;
  assign n25925 = ~i_RtoB_ACK0 & ~n25924;
  assign n25926 = ~n24135 & ~n25925;
  assign n25927 = controllable_DEQ & ~n25926;
  assign n25928 = ~controllable_BtoR_REQ0 & ~n8781;
  assign n25929 = ~n14615 & ~n25928;
  assign n25930 = ~i_RtoB_ACK0 & ~n25929;
  assign n25931 = ~n24141 & ~n25930;
  assign n25932 = ~controllable_DEQ & ~n25931;
  assign n25933 = ~n25927 & ~n25932;
  assign n25934 = i_FULL & ~n25933;
  assign n25935 = ~n5245 & ~n8763;
  assign n25936 = ~controllable_BtoR_REQ0 & ~n25935;
  assign n25937 = ~n14598 & ~n25936;
  assign n25938 = ~i_RtoB_ACK0 & ~n25937;
  assign n25939 = ~n24135 & ~n25938;
  assign n25940 = controllable_DEQ & ~n25939;
  assign n25941 = ~n8782 & ~n18888;
  assign n25942 = ~controllable_BtoR_REQ0 & ~n25941;
  assign n25943 = ~n14615 & ~n25942;
  assign n25944 = ~i_RtoB_ACK0 & ~n25943;
  assign n25945 = ~n24141 & ~n25944;
  assign n25946 = ~controllable_DEQ & ~n25945;
  assign n25947 = ~n25940 & ~n25946;
  assign n25948 = ~i_FULL & ~n25947;
  assign n25949 = ~n25934 & ~n25948;
  assign n25950 = i_nEMPTY & ~n25949;
  assign n25951 = ~controllable_BtoR_REQ0 & ~n8818;
  assign n25952 = ~n14634 & ~n25951;
  assign n25953 = ~i_RtoB_ACK0 & ~n25952;
  assign n25954 = ~n24135 & ~n25953;
  assign n25955 = ~controllable_DEQ & ~n25954;
  assign n25956 = ~n22013 & ~n25955;
  assign n25957 = i_FULL & ~n25956;
  assign n25958 = ~n8763 & ~n18917;
  assign n25959 = ~controllable_BtoR_REQ0 & ~n25958;
  assign n25960 = ~n14598 & ~n25959;
  assign n25961 = ~i_RtoB_ACK0 & ~n25960;
  assign n25962 = ~n24135 & ~n25961;
  assign n25963 = ~controllable_DEQ & ~n25962;
  assign n25964 = ~n22023 & ~n25963;
  assign n25965 = ~i_FULL & ~n25964;
  assign n25966 = ~n25957 & ~n25965;
  assign n25967 = ~i_nEMPTY & ~n25966;
  assign n25968 = ~n25950 & ~n25967;
  assign n25969 = controllable_BtoS_ACK0 & ~n25968;
  assign n25970 = ~n8863 & ~n18931;
  assign n25971 = ~controllable_BtoR_REQ0 & ~n25970;
  assign n25972 = ~n14673 & ~n25971;
  assign n25973 = ~i_RtoB_ACK0 & ~n25972;
  assign n25974 = ~n24161 & ~n25973;
  assign n25975 = controllable_DEQ & ~n25974;
  assign n25976 = ~controllable_BtoR_REQ0 & ~n8884;
  assign n25977 = ~n14690 & ~n25976;
  assign n25978 = ~i_RtoB_ACK0 & ~n25977;
  assign n25979 = ~n24167 & ~n25978;
  assign n25980 = ~controllable_DEQ & ~n25979;
  assign n25981 = ~n25975 & ~n25980;
  assign n25982 = i_FULL & ~n25981;
  assign n25983 = ~n8863 & ~n18948;
  assign n25984 = ~controllable_BtoR_REQ0 & ~n25983;
  assign n25985 = ~n14673 & ~n25984;
  assign n25986 = ~i_RtoB_ACK0 & ~n25985;
  assign n25987 = ~n24161 & ~n25986;
  assign n25988 = controllable_DEQ & ~n25987;
  assign n25989 = ~n8885 & ~n18956;
  assign n25990 = ~controllable_BtoR_REQ0 & ~n25989;
  assign n25991 = ~n14690 & ~n25990;
  assign n25992 = ~i_RtoB_ACK0 & ~n25991;
  assign n25993 = ~n24167 & ~n25992;
  assign n25994 = ~controllable_DEQ & ~n25993;
  assign n25995 = ~n25988 & ~n25994;
  assign n25996 = ~i_FULL & ~n25995;
  assign n25997 = ~n25982 & ~n25996;
  assign n25998 = i_nEMPTY & ~n25997;
  assign n25999 = ~controllable_BtoR_REQ0 & ~n8925;
  assign n26000 = ~n14709 & ~n25999;
  assign n26001 = ~i_RtoB_ACK0 & ~n26000;
  assign n26002 = ~n24161 & ~n26001;
  assign n26003 = ~controllable_DEQ & ~n26002;
  assign n26004 = ~n22063 & ~n26003;
  assign n26005 = i_FULL & ~n26004;
  assign n26006 = ~n8863 & ~n18987;
  assign n26007 = ~controllable_BtoR_REQ0 & ~n26006;
  assign n26008 = ~n14673 & ~n26007;
  assign n26009 = ~i_RtoB_ACK0 & ~n26008;
  assign n26010 = ~n24161 & ~n26009;
  assign n26011 = ~controllable_DEQ & ~n26010;
  assign n26012 = ~n22073 & ~n26011;
  assign n26013 = ~i_FULL & ~n26012;
  assign n26014 = ~n26005 & ~n26013;
  assign n26015 = ~i_nEMPTY & ~n26014;
  assign n26016 = ~n25998 & ~n26015;
  assign n26017 = ~controllable_BtoS_ACK0 & ~n26016;
  assign n26018 = ~n25969 & ~n26017;
  assign n26019 = n4465 & ~n26018;
  assign n26020 = ~n8972 & ~n19003;
  assign n26021 = ~controllable_BtoR_REQ0 & ~n26020;
  assign n26022 = ~n14824 & ~n26021;
  assign n26023 = ~i_RtoB_ACK0 & ~n26022;
  assign n26024 = ~n24189 & ~n26023;
  assign n26025 = controllable_DEQ & ~n26024;
  assign n26026 = ~controllable_BtoR_REQ0 & ~n8990;
  assign n26027 = ~n14841 & ~n26026;
  assign n26028 = ~i_RtoB_ACK0 & ~n26027;
  assign n26029 = ~n24195 & ~n26028;
  assign n26030 = ~controllable_DEQ & ~n26029;
  assign n26031 = ~n26025 & ~n26030;
  assign n26032 = i_FULL & ~n26031;
  assign n26033 = ~n8972 & ~n18948;
  assign n26034 = ~controllable_BtoR_REQ0 & ~n26033;
  assign n26035 = ~n14824 & ~n26034;
  assign n26036 = ~i_RtoB_ACK0 & ~n26035;
  assign n26037 = ~n24189 & ~n26036;
  assign n26038 = controllable_DEQ & ~n26037;
  assign n26039 = ~n8991 & ~n19024;
  assign n26040 = ~controllable_BtoR_REQ0 & ~n26039;
  assign n26041 = ~n14841 & ~n26040;
  assign n26042 = ~i_RtoB_ACK0 & ~n26041;
  assign n26043 = ~n24195 & ~n26042;
  assign n26044 = ~controllable_DEQ & ~n26043;
  assign n26045 = ~n26038 & ~n26044;
  assign n26046 = ~i_FULL & ~n26045;
  assign n26047 = ~n26032 & ~n26046;
  assign n26048 = i_nEMPTY & ~n26047;
  assign n26049 = ~controllable_BtoR_REQ0 & ~n9027;
  assign n26050 = ~n14860 & ~n26049;
  assign n26051 = ~i_RtoB_ACK0 & ~n26050;
  assign n26052 = ~n24189 & ~n26051;
  assign n26053 = ~controllable_DEQ & ~n26052;
  assign n26054 = ~n22115 & ~n26053;
  assign n26055 = i_FULL & ~n26054;
  assign n26056 = ~n8972 & ~n19053;
  assign n26057 = ~controllable_BtoR_REQ0 & ~n26056;
  assign n26058 = ~n14824 & ~n26057;
  assign n26059 = ~i_RtoB_ACK0 & ~n26058;
  assign n26060 = ~n24189 & ~n26059;
  assign n26061 = ~controllable_DEQ & ~n26060;
  assign n26062 = ~n22125 & ~n26061;
  assign n26063 = ~i_FULL & ~n26062;
  assign n26064 = ~n26055 & ~n26063;
  assign n26065 = ~i_nEMPTY & ~n26064;
  assign n26066 = ~n26048 & ~n26065;
  assign n26067 = ~controllable_BtoS_ACK0 & ~n26066;
  assign n26068 = ~n21013 & ~n26067;
  assign n26069 = ~n4465 & ~n26068;
  assign n26070 = ~n26019 & ~n26069;
  assign n26071 = i_StoB_REQ10 & ~n26070;
  assign n26072 = ~n13246 & ~n19078;
  assign n26073 = ~controllable_BtoR_REQ0 & ~n26072;
  assign n26074 = ~n14904 & ~n26073;
  assign n26075 = ~i_RtoB_ACK0 & ~n26074;
  assign n26076 = ~n24219 & ~n26075;
  assign n26077 = controllable_DEQ & ~n26076;
  assign n26078 = ~n13255 & ~n19092;
  assign n26079 = ~controllable_BtoR_REQ0 & ~n26078;
  assign n26080 = ~n14923 & ~n26079;
  assign n26081 = ~i_RtoB_ACK0 & ~n26080;
  assign n26082 = ~n24225 & ~n26081;
  assign n26083 = ~controllable_DEQ & ~n26082;
  assign n26084 = ~n26077 & ~n26083;
  assign n26085 = i_FULL & ~n26084;
  assign n26086 = ~n13265 & ~n19102;
  assign n26087 = ~controllable_BtoR_REQ0 & ~n26086;
  assign n26088 = ~n14942 & ~n26087;
  assign n26089 = ~i_RtoB_ACK0 & ~n26088;
  assign n26090 = ~n24219 & ~n26089;
  assign n26091 = controllable_DEQ & ~n26090;
  assign n26092 = ~n13273 & ~n19110;
  assign n26093 = ~controllable_BtoR_REQ0 & ~n26092;
  assign n26094 = ~n14958 & ~n26093;
  assign n26095 = ~i_RtoB_ACK0 & ~n26094;
  assign n26096 = ~n24225 & ~n26095;
  assign n26097 = ~controllable_DEQ & ~n26096;
  assign n26098 = ~n26091 & ~n26097;
  assign n26099 = ~i_FULL & ~n26098;
  assign n26100 = ~n26085 & ~n26099;
  assign n26101 = i_nEMPTY & ~n26100;
  assign n26102 = ~n13286 & ~n19134;
  assign n26103 = ~controllable_BtoR_REQ0 & ~n26102;
  assign n26104 = ~n14995 & ~n26103;
  assign n26105 = ~i_RtoB_ACK0 & ~n26104;
  assign n26106 = ~n24245 & ~n26105;
  assign n26107 = ~controllable_DEQ & ~n26106;
  assign n26108 = ~n22169 & ~n26107;
  assign n26109 = i_FULL & ~n26108;
  assign n26110 = ~n13246 & ~n19150;
  assign n26111 = ~controllable_BtoR_REQ0 & ~n26110;
  assign n26112 = ~n14904 & ~n26111;
  assign n26113 = ~i_RtoB_ACK0 & ~n26112;
  assign n26114 = ~n24219 & ~n26113;
  assign n26115 = ~controllable_DEQ & ~n26114;
  assign n26116 = ~n22181 & ~n26115;
  assign n26117 = ~i_FULL & ~n26116;
  assign n26118 = ~n26109 & ~n26117;
  assign n26119 = ~i_nEMPTY & ~n26118;
  assign n26120 = ~n26101 & ~n26119;
  assign n26121 = controllable_BtoS_ACK0 & ~n26120;
  assign n26122 = ~n13310 & ~n19171;
  assign n26123 = ~controllable_BtoR_REQ0 & ~n26122;
  assign n26124 = ~n15046 & ~n26123;
  assign n26125 = ~i_RtoB_ACK0 & ~n26124;
  assign n26126 = ~n24263 & ~n26125;
  assign n26127 = controllable_DEQ & ~n26126;
  assign n26128 = ~n13319 & ~n19185;
  assign n26129 = ~controllable_BtoR_REQ0 & ~n26128;
  assign n26130 = ~n15065 & ~n26129;
  assign n26131 = ~i_RtoB_ACK0 & ~n26130;
  assign n26132 = ~n24269 & ~n26131;
  assign n26133 = ~controllable_DEQ & ~n26132;
  assign n26134 = ~n26127 & ~n26133;
  assign n26135 = i_FULL & ~n26134;
  assign n26136 = ~n13329 & ~n19195;
  assign n26137 = ~controllable_BtoR_REQ0 & ~n26136;
  assign n26138 = ~n15084 & ~n26137;
  assign n26139 = ~i_RtoB_ACK0 & ~n26138;
  assign n26140 = ~n24263 & ~n26139;
  assign n26141 = controllable_DEQ & ~n26140;
  assign n26142 = ~n13337 & ~n19203;
  assign n26143 = ~controllable_BtoR_REQ0 & ~n26142;
  assign n26144 = ~n15100 & ~n26143;
  assign n26145 = ~i_RtoB_ACK0 & ~n26144;
  assign n26146 = ~n24269 & ~n26145;
  assign n26147 = ~controllable_DEQ & ~n26146;
  assign n26148 = ~n26141 & ~n26147;
  assign n26149 = ~i_FULL & ~n26148;
  assign n26150 = ~n26135 & ~n26149;
  assign n26151 = i_nEMPTY & ~n26150;
  assign n26152 = ~n13350 & ~n19227;
  assign n26153 = ~controllable_BtoR_REQ0 & ~n26152;
  assign n26154 = ~n15137 & ~n26153;
  assign n26155 = ~i_RtoB_ACK0 & ~n26154;
  assign n26156 = ~n24289 & ~n26155;
  assign n26157 = ~controllable_DEQ & ~n26156;
  assign n26158 = ~n22221 & ~n26157;
  assign n26159 = i_FULL & ~n26158;
  assign n26160 = ~n13310 & ~n19243;
  assign n26161 = ~controllable_BtoR_REQ0 & ~n26160;
  assign n26162 = ~n15046 & ~n26161;
  assign n26163 = ~i_RtoB_ACK0 & ~n26162;
  assign n26164 = ~n24263 & ~n26163;
  assign n26165 = ~controllable_DEQ & ~n26164;
  assign n26166 = ~n22233 & ~n26165;
  assign n26167 = ~i_FULL & ~n26166;
  assign n26168 = ~n26159 & ~n26167;
  assign n26169 = ~i_nEMPTY & ~n26168;
  assign n26170 = ~n26151 & ~n26169;
  assign n26171 = ~controllable_BtoS_ACK0 & ~n26170;
  assign n26172 = ~n26121 & ~n26171;
  assign n26173 = n4465 & ~n26172;
  assign n26174 = ~n13376 & ~n19259;
  assign n26175 = ~controllable_BtoR_REQ0 & ~n26174;
  assign n26176 = ~n15190 & ~n26175;
  assign n26177 = ~i_RtoB_ACK0 & ~n26176;
  assign n26178 = ~n24309 & ~n26177;
  assign n26179 = controllable_DEQ & ~n26178;
  assign n26180 = ~n13385 & ~n19267;
  assign n26181 = ~controllable_BtoR_REQ0 & ~n26180;
  assign n26182 = ~n15209 & ~n26181;
  assign n26183 = ~i_RtoB_ACK0 & ~n26182;
  assign n26184 = ~n24315 & ~n26183;
  assign n26185 = ~controllable_DEQ & ~n26184;
  assign n26186 = ~n26179 & ~n26185;
  assign n26187 = i_nEMPTY & ~n26186;
  assign n26188 = ~n13396 & ~n19283;
  assign n26189 = ~controllable_BtoR_REQ0 & ~n26188;
  assign n26190 = ~n15237 & ~n26189;
  assign n26191 = ~i_RtoB_ACK0 & ~n26190;
  assign n26192 = ~n24323 & ~n26191;
  assign n26193 = ~controllable_DEQ & ~n26192;
  assign n26194 = ~n22263 & ~n26193;
  assign n26195 = i_FULL & ~n26194;
  assign n26196 = ~n13376 & ~n19299;
  assign n26197 = ~controllable_BtoR_REQ0 & ~n26196;
  assign n26198 = ~n15190 & ~n26197;
  assign n26199 = ~i_RtoB_ACK0 & ~n26198;
  assign n26200 = ~n24309 & ~n26199;
  assign n26201 = ~controllable_DEQ & ~n26200;
  assign n26202 = ~n22275 & ~n26201;
  assign n26203 = ~i_FULL & ~n26202;
  assign n26204 = ~n26195 & ~n26203;
  assign n26205 = ~i_nEMPTY & ~n26204;
  assign n26206 = ~n26187 & ~n26205;
  assign n26207 = controllable_BtoS_ACK0 & ~n26206;
  assign n26208 = ~n9881 & ~n19313;
  assign n26209 = ~controllable_BtoR_REQ0 & ~n26208;
  assign n26210 = ~n15281 & ~n26209;
  assign n26211 = ~i_RtoB_ACK0 & ~n26210;
  assign n26212 = ~n24341 & ~n26211;
  assign n26213 = controllable_DEQ & ~n26212;
  assign n26214 = ~n9912 & ~n19321;
  assign n26215 = ~controllable_BtoR_REQ0 & ~n26214;
  assign n26216 = ~n15300 & ~n26215;
  assign n26217 = ~i_RtoB_ACK0 & ~n26216;
  assign n26218 = ~n24347 & ~n26217;
  assign n26219 = ~controllable_DEQ & ~n26218;
  assign n26220 = ~n26213 & ~n26219;
  assign n26221 = i_FULL & ~n26220;
  assign n26222 = ~n9925 & ~n11317;
  assign n26223 = ~controllable_BtoR_REQ0 & ~n26222;
  assign n26224 = ~n15319 & ~n26223;
  assign n26225 = ~i_RtoB_ACK0 & ~n26224;
  assign n26226 = ~n24341 & ~n26225;
  assign n26227 = controllable_DEQ & ~n26226;
  assign n26228 = ~n9935 & ~n19335;
  assign n26229 = ~controllable_BtoR_REQ0 & ~n26228;
  assign n26230 = ~n15335 & ~n26229;
  assign n26231 = ~i_RtoB_ACK0 & ~n26230;
  assign n26232 = ~n24347 & ~n26231;
  assign n26233 = ~controllable_DEQ & ~n26232;
  assign n26234 = ~n26227 & ~n26233;
  assign n26235 = ~i_FULL & ~n26234;
  assign n26236 = ~n26221 & ~n26235;
  assign n26237 = i_nEMPTY & ~n26236;
  assign n26238 = ~n9959 & ~n19351;
  assign n26239 = ~controllable_BtoR_REQ0 & ~n26238;
  assign n26240 = ~n15372 & ~n26239;
  assign n26241 = ~i_RtoB_ACK0 & ~n26240;
  assign n26242 = ~n24367 & ~n26241;
  assign n26243 = ~controllable_DEQ & ~n26242;
  assign n26244 = ~n22315 & ~n26243;
  assign n26245 = i_FULL & ~n26244;
  assign n26246 = ~n9881 & ~n19365;
  assign n26247 = ~controllable_BtoR_REQ0 & ~n26246;
  assign n26248 = ~n15281 & ~n26247;
  assign n26249 = ~i_RtoB_ACK0 & ~n26248;
  assign n26250 = ~n24341 & ~n26249;
  assign n26251 = ~controllable_DEQ & ~n26250;
  assign n26252 = ~n22327 & ~n26251;
  assign n26253 = ~i_FULL & ~n26252;
  assign n26254 = ~n26245 & ~n26253;
  assign n26255 = ~i_nEMPTY & ~n26254;
  assign n26256 = ~n26237 & ~n26255;
  assign n26257 = ~controllable_BtoS_ACK0 & ~n26256;
  assign n26258 = ~n26207 & ~n26257;
  assign n26259 = ~n4465 & ~n26258;
  assign n26260 = ~n26173 & ~n26259;
  assign n26261 = ~i_StoB_REQ10 & ~n26260;
  assign n26262 = ~n26071 & ~n26261;
  assign n26263 = controllable_BtoS_ACK10 & ~n26262;
  assign n26264 = ~n10011 & ~n19386;
  assign n26265 = ~controllable_BtoR_REQ0 & ~n26264;
  assign n26266 = ~n19384 & ~n26265;
  assign n26267 = ~i_RtoB_ACK0 & ~n26266;
  assign n26268 = ~n24391 & ~n26267;
  assign n26269 = controllable_DEQ & ~n26268;
  assign n26270 = ~n9519 & ~n19395;
  assign n26271 = ~controllable_BtoR_REQ0 & ~n26270;
  assign n26272 = ~n19393 & ~n26271;
  assign n26273 = ~i_RtoB_ACK0 & ~n26272;
  assign n26274 = ~n24397 & ~n26273;
  assign n26275 = ~controllable_DEQ & ~n26274;
  assign n26276 = ~n26269 & ~n26275;
  assign n26277 = i_FULL & ~n26276;
  assign n26278 = ~n10031 & ~n11238;
  assign n26279 = ~controllable_BtoR_REQ0 & ~n26278;
  assign n26280 = ~n19404 & ~n26279;
  assign n26281 = ~i_RtoB_ACK0 & ~n26280;
  assign n26282 = ~n24391 & ~n26281;
  assign n26283 = controllable_DEQ & ~n26282;
  assign n26284 = ~n9544 & ~n19411;
  assign n26285 = ~controllable_BtoR_REQ0 & ~n26284;
  assign n26286 = ~n19409 & ~n26285;
  assign n26287 = ~i_RtoB_ACK0 & ~n26286;
  assign n26288 = ~n24397 & ~n26287;
  assign n26289 = ~controllable_DEQ & ~n26288;
  assign n26290 = ~n26283 & ~n26289;
  assign n26291 = ~i_FULL & ~n26290;
  assign n26292 = ~n26277 & ~n26291;
  assign n26293 = i_nEMPTY & ~n26292;
  assign n26294 = ~n9573 & ~n19429;
  assign n26295 = ~controllable_BtoR_REQ0 & ~n26294;
  assign n26296 = ~n19427 & ~n26295;
  assign n26297 = ~i_RtoB_ACK0 & ~n26296;
  assign n26298 = ~n24417 & ~n26297;
  assign n26299 = ~controllable_DEQ & ~n26298;
  assign n26300 = ~n22373 & ~n26299;
  assign n26301 = i_FULL & ~n26300;
  assign n26302 = ~controllable_DEQ & ~n26268;
  assign n26303 = ~n22385 & ~n26302;
  assign n26304 = ~i_FULL & ~n26303;
  assign n26305 = ~n26301 & ~n26304;
  assign n26306 = ~i_nEMPTY & ~n26305;
  assign n26307 = ~n26293 & ~n26306;
  assign n26308 = controllable_BtoS_ACK0 & ~n26307;
  assign n26309 = ~n10084 & ~n19452;
  assign n26310 = ~controllable_BtoR_REQ0 & ~n26309;
  assign n26311 = ~n19450 & ~n26310;
  assign n26312 = ~i_RtoB_ACK0 & ~n26311;
  assign n26313 = ~n24432 & ~n26312;
  assign n26314 = controllable_DEQ & ~n26313;
  assign n26315 = ~n9666 & ~n19461;
  assign n26316 = ~controllable_BtoR_REQ0 & ~n26315;
  assign n26317 = ~n19459 & ~n26316;
  assign n26318 = ~i_RtoB_ACK0 & ~n26317;
  assign n26319 = ~n24438 & ~n26318;
  assign n26320 = ~controllable_DEQ & ~n26319;
  assign n26321 = ~n26314 & ~n26320;
  assign n26322 = i_FULL & ~n26321;
  assign n26323 = ~n10104 & ~n11317;
  assign n26324 = ~controllable_BtoR_REQ0 & ~n26323;
  assign n26325 = ~n19470 & ~n26324;
  assign n26326 = ~i_RtoB_ACK0 & ~n26325;
  assign n26327 = ~n24432 & ~n26326;
  assign n26328 = controllable_DEQ & ~n26327;
  assign n26329 = ~n9691 & ~n19477;
  assign n26330 = ~controllable_BtoR_REQ0 & ~n26329;
  assign n26331 = ~n19475 & ~n26330;
  assign n26332 = ~i_RtoB_ACK0 & ~n26331;
  assign n26333 = ~n24438 & ~n26332;
  assign n26334 = ~controllable_DEQ & ~n26333;
  assign n26335 = ~n26328 & ~n26334;
  assign n26336 = ~i_FULL & ~n26335;
  assign n26337 = ~n26322 & ~n26336;
  assign n26338 = i_nEMPTY & ~n26337;
  assign n26339 = ~n9720 & ~n19495;
  assign n26340 = ~controllable_BtoR_REQ0 & ~n26339;
  assign n26341 = ~n19493 & ~n26340;
  assign n26342 = ~i_RtoB_ACK0 & ~n26341;
  assign n26343 = ~n24458 & ~n26342;
  assign n26344 = ~controllable_DEQ & ~n26343;
  assign n26345 = ~n22422 & ~n26344;
  assign n26346 = i_FULL & ~n26345;
  assign n26347 = ~controllable_DEQ & ~n26313;
  assign n26348 = ~n22434 & ~n26347;
  assign n26349 = ~i_FULL & ~n26348;
  assign n26350 = ~n26346 & ~n26349;
  assign n26351 = ~i_nEMPTY & ~n26350;
  assign n26352 = ~n26338 & ~n26351;
  assign n26353 = ~controllable_BtoS_ACK0 & ~n26352;
  assign n26354 = ~n26308 & ~n26353;
  assign n26355 = n4465 & ~n26354;
  assign n26356 = ~n10151 & ~n11238;
  assign n26357 = ~controllable_BtoR_REQ0 & ~n26356;
  assign n26358 = ~n19518 & ~n26357;
  assign n26359 = ~i_RtoB_ACK0 & ~n26358;
  assign n26360 = ~n24475 & ~n26359;
  assign n26361 = controllable_DEQ & ~n26360;
  assign n26362 = ~n9812 & ~n11248;
  assign n26363 = ~controllable_BtoR_REQ0 & ~n26362;
  assign n26364 = ~n19523 & ~n26363;
  assign n26365 = ~i_RtoB_ACK0 & ~n26364;
  assign n26366 = ~n24481 & ~n26365;
  assign n26367 = ~controllable_DEQ & ~n26366;
  assign n26368 = ~n26361 & ~n26367;
  assign n26369 = i_nEMPTY & ~n26368;
  assign n26370 = ~n9835 & ~n11230;
  assign n26371 = ~controllable_BtoR_REQ0 & ~n26370;
  assign n26372 = ~n19535 & ~n26371;
  assign n26373 = ~i_RtoB_ACK0 & ~n26372;
  assign n26374 = ~n24489 & ~n26373;
  assign n26375 = ~controllable_DEQ & ~n26374;
  assign n26376 = ~n22461 & ~n26375;
  assign n26377 = i_FULL & ~n26376;
  assign n26378 = ~controllable_DEQ & ~n26360;
  assign n26379 = ~n22473 & ~n26378;
  assign n26380 = ~i_FULL & ~n26379;
  assign n26381 = ~n26377 & ~n26380;
  assign n26382 = ~i_nEMPTY & ~n26381;
  assign n26383 = ~n26369 & ~n26382;
  assign n26384 = controllable_BtoS_ACK0 & ~n26383;
  assign n26385 = ~n10198 & ~n19313;
  assign n26386 = ~controllable_BtoR_REQ0 & ~n26385;
  assign n26387 = ~n19554 & ~n26386;
  assign n26388 = ~i_RtoB_ACK0 & ~n26387;
  assign n26389 = ~n24504 & ~n26388;
  assign n26390 = controllable_DEQ & ~n26389;
  assign n26391 = ~n19559 & ~n26215;
  assign n26392 = ~i_RtoB_ACK0 & ~n26391;
  assign n26393 = ~n24510 & ~n26392;
  assign n26394 = ~controllable_DEQ & ~n26393;
  assign n26395 = ~n26390 & ~n26394;
  assign n26396 = i_FULL & ~n26395;
  assign n26397 = ~n10214 & ~n11317;
  assign n26398 = ~controllable_BtoR_REQ0 & ~n26397;
  assign n26399 = ~n19566 & ~n26398;
  assign n26400 = ~i_RtoB_ACK0 & ~n26399;
  assign n26401 = ~n24504 & ~n26400;
  assign n26402 = controllable_DEQ & ~n26401;
  assign n26403 = ~n19571 & ~n26229;
  assign n26404 = ~i_RtoB_ACK0 & ~n26403;
  assign n26405 = ~n24510 & ~n26404;
  assign n26406 = ~controllable_DEQ & ~n26405;
  assign n26407 = ~n26402 & ~n26406;
  assign n26408 = ~i_FULL & ~n26407;
  assign n26409 = ~n26396 & ~n26408;
  assign n26410 = i_nEMPTY & ~n26409;
  assign n26411 = ~n19585 & ~n26239;
  assign n26412 = ~i_RtoB_ACK0 & ~n26411;
  assign n26413 = ~n24530 & ~n26412;
  assign n26414 = ~controllable_DEQ & ~n26413;
  assign n26415 = ~n22510 & ~n26414;
  assign n26416 = i_FULL & ~n26415;
  assign n26417 = ~controllable_DEQ & ~n26389;
  assign n26418 = ~n22522 & ~n26417;
  assign n26419 = ~i_FULL & ~n26418;
  assign n26420 = ~n26416 & ~n26419;
  assign n26421 = ~i_nEMPTY & ~n26420;
  assign n26422 = ~n26410 & ~n26421;
  assign n26423 = ~controllable_BtoS_ACK0 & ~n26422;
  assign n26424 = ~n26384 & ~n26423;
  assign n26425 = ~n4465 & ~n26424;
  assign n26426 = ~n26355 & ~n26425;
  assign n26427 = i_StoB_REQ10 & ~n26426;
  assign n26428 = ~n26261 & ~n26427;
  assign n26429 = ~controllable_BtoS_ACK10 & ~n26428;
  assign n26430 = ~n26263 & ~n26429;
  assign n26431 = n4464 & ~n26430;
  assign n26432 = ~n10265 & ~n19613;
  assign n26433 = ~controllable_BtoR_REQ0 & ~n26432;
  assign n26434 = ~n15732 & ~n26433;
  assign n26435 = ~i_RtoB_ACK0 & ~n26434;
  assign n26436 = ~n24553 & ~n26435;
  assign n26437 = controllable_DEQ & ~n26436;
  assign n26438 = ~controllable_BtoR_REQ0 & ~n10283;
  assign n26439 = ~n15749 & ~n26438;
  assign n26440 = ~i_RtoB_ACK0 & ~n26439;
  assign n26441 = ~n24559 & ~n26440;
  assign n26442 = ~controllable_DEQ & ~n26441;
  assign n26443 = ~n26437 & ~n26442;
  assign n26444 = i_FULL & ~n26443;
  assign n26445 = ~n5245 & ~n10265;
  assign n26446 = ~controllable_BtoR_REQ0 & ~n26445;
  assign n26447 = ~n15732 & ~n26446;
  assign n26448 = ~i_RtoB_ACK0 & ~n26447;
  assign n26449 = ~n24553 & ~n26448;
  assign n26450 = controllable_DEQ & ~n26449;
  assign n26451 = ~n10284 & ~n19634;
  assign n26452 = ~controllable_BtoR_REQ0 & ~n26451;
  assign n26453 = ~n15749 & ~n26452;
  assign n26454 = ~i_RtoB_ACK0 & ~n26453;
  assign n26455 = ~n24559 & ~n26454;
  assign n26456 = ~controllable_DEQ & ~n26455;
  assign n26457 = ~n26450 & ~n26456;
  assign n26458 = ~i_FULL & ~n26457;
  assign n26459 = ~n26444 & ~n26458;
  assign n26460 = i_nEMPTY & ~n26459;
  assign n26461 = ~controllable_BtoR_REQ0 & ~n10320;
  assign n26462 = ~n15768 & ~n26461;
  assign n26463 = ~i_RtoB_ACK0 & ~n26462;
  assign n26464 = ~n24553 & ~n26463;
  assign n26465 = ~controllable_DEQ & ~n26464;
  assign n26466 = ~n22567 & ~n26465;
  assign n26467 = i_FULL & ~n26466;
  assign n26468 = ~n10265 & ~n19663;
  assign n26469 = ~controllable_BtoR_REQ0 & ~n26468;
  assign n26470 = ~n15732 & ~n26469;
  assign n26471 = ~i_RtoB_ACK0 & ~n26470;
  assign n26472 = ~n24553 & ~n26471;
  assign n26473 = ~controllable_DEQ & ~n26472;
  assign n26474 = ~n22577 & ~n26473;
  assign n26475 = ~i_FULL & ~n26474;
  assign n26476 = ~n26467 & ~n26475;
  assign n26477 = ~i_nEMPTY & ~n26476;
  assign n26478 = ~n26460 & ~n26477;
  assign n26479 = controllable_BtoS_ACK0 & ~n26478;
  assign n26480 = ~n10359 & ~n19677;
  assign n26481 = ~controllable_BtoR_REQ0 & ~n26480;
  assign n26482 = ~n15807 & ~n26481;
  assign n26483 = ~i_RtoB_ACK0 & ~n26482;
  assign n26484 = ~n24579 & ~n26483;
  assign n26485 = controllable_DEQ & ~n26484;
  assign n26486 = ~controllable_BtoR_REQ0 & ~n10377;
  assign n26487 = ~n15824 & ~n26486;
  assign n26488 = ~i_RtoB_ACK0 & ~n26487;
  assign n26489 = ~n24585 & ~n26488;
  assign n26490 = ~controllable_DEQ & ~n26489;
  assign n26491 = ~n26485 & ~n26490;
  assign n26492 = i_FULL & ~n26491;
  assign n26493 = ~n10359 & ~n18948;
  assign n26494 = ~controllable_BtoR_REQ0 & ~n26493;
  assign n26495 = ~n15807 & ~n26494;
  assign n26496 = ~i_RtoB_ACK0 & ~n26495;
  assign n26497 = ~n24579 & ~n26496;
  assign n26498 = controllable_DEQ & ~n26497;
  assign n26499 = ~n10378 & ~n19698;
  assign n26500 = ~controllable_BtoR_REQ0 & ~n26499;
  assign n26501 = ~n15824 & ~n26500;
  assign n26502 = ~i_RtoB_ACK0 & ~n26501;
  assign n26503 = ~n24585 & ~n26502;
  assign n26504 = ~controllable_DEQ & ~n26503;
  assign n26505 = ~n26498 & ~n26504;
  assign n26506 = ~i_FULL & ~n26505;
  assign n26507 = ~n26492 & ~n26506;
  assign n26508 = i_nEMPTY & ~n26507;
  assign n26509 = ~controllable_BtoR_REQ0 & ~n10414;
  assign n26510 = ~n15843 & ~n26509;
  assign n26511 = ~i_RtoB_ACK0 & ~n26510;
  assign n26512 = ~n24579 & ~n26511;
  assign n26513 = ~controllable_DEQ & ~n26512;
  assign n26514 = ~n22617 & ~n26513;
  assign n26515 = i_FULL & ~n26514;
  assign n26516 = ~n10359 & ~n19727;
  assign n26517 = ~controllable_BtoR_REQ0 & ~n26516;
  assign n26518 = ~n15807 & ~n26517;
  assign n26519 = ~i_RtoB_ACK0 & ~n26518;
  assign n26520 = ~n24579 & ~n26519;
  assign n26521 = ~controllable_DEQ & ~n26520;
  assign n26522 = ~n22627 & ~n26521;
  assign n26523 = ~i_FULL & ~n26522;
  assign n26524 = ~n26515 & ~n26523;
  assign n26525 = ~i_nEMPTY & ~n26524;
  assign n26526 = ~n26508 & ~n26525;
  assign n26527 = ~controllable_BtoS_ACK0 & ~n26526;
  assign n26528 = ~n26479 & ~n26527;
  assign n26529 = n4465 & ~n26528;
  assign n26530 = ~n21013 & ~n26527;
  assign n26531 = ~n4465 & ~n26530;
  assign n26532 = ~n26529 & ~n26531;
  assign n26533 = i_StoB_REQ10 & ~n26532;
  assign n26534 = ~n13698 & ~n19747;
  assign n26535 = ~controllable_BtoR_REQ0 & ~n26534;
  assign n26536 = ~n15889 & ~n26535;
  assign n26537 = ~i_RtoB_ACK0 & ~n26536;
  assign n26538 = ~n24611 & ~n26537;
  assign n26539 = controllable_DEQ & ~n26538;
  assign n26540 = ~n13707 & ~n19755;
  assign n26541 = ~controllable_BtoR_REQ0 & ~n26540;
  assign n26542 = ~n15908 & ~n26541;
  assign n26543 = ~i_RtoB_ACK0 & ~n26542;
  assign n26544 = ~n24617 & ~n26543;
  assign n26545 = ~controllable_DEQ & ~n26544;
  assign n26546 = ~n26539 & ~n26545;
  assign n26547 = i_FULL & ~n26546;
  assign n26548 = ~n13717 & ~n19765;
  assign n26549 = ~controllable_BtoR_REQ0 & ~n26548;
  assign n26550 = ~n15927 & ~n26549;
  assign n26551 = ~i_RtoB_ACK0 & ~n26550;
  assign n26552 = ~n24611 & ~n26551;
  assign n26553 = controllable_DEQ & ~n26552;
  assign n26554 = ~n13725 & ~n19773;
  assign n26555 = ~controllable_BtoR_REQ0 & ~n26554;
  assign n26556 = ~n15943 & ~n26555;
  assign n26557 = ~i_RtoB_ACK0 & ~n26556;
  assign n26558 = ~n24617 & ~n26557;
  assign n26559 = ~controllable_DEQ & ~n26558;
  assign n26560 = ~n26553 & ~n26559;
  assign n26561 = ~i_FULL & ~n26560;
  assign n26562 = ~n26547 & ~n26561;
  assign n26563 = i_nEMPTY & ~n26562;
  assign n26564 = ~n13738 & ~n19791;
  assign n26565 = ~controllable_BtoR_REQ0 & ~n26564;
  assign n26566 = ~n15980 & ~n26565;
  assign n26567 = ~i_RtoB_ACK0 & ~n26566;
  assign n26568 = ~n24637 & ~n26567;
  assign n26569 = ~controllable_DEQ & ~n26568;
  assign n26570 = ~n22673 & ~n26569;
  assign n26571 = i_FULL & ~n26570;
  assign n26572 = ~n13698 & ~n19807;
  assign n26573 = ~controllable_BtoR_REQ0 & ~n26572;
  assign n26574 = ~n15889 & ~n26573;
  assign n26575 = ~i_RtoB_ACK0 & ~n26574;
  assign n26576 = ~n24611 & ~n26575;
  assign n26577 = ~controllable_DEQ & ~n26576;
  assign n26578 = ~n22685 & ~n26577;
  assign n26579 = ~i_FULL & ~n26578;
  assign n26580 = ~n26571 & ~n26579;
  assign n26581 = ~i_nEMPTY & ~n26580;
  assign n26582 = ~n26563 & ~n26581;
  assign n26583 = controllable_BtoS_ACK0 & ~n26582;
  assign n26584 = ~n13762 & ~n19821;
  assign n26585 = ~controllable_BtoR_REQ0 & ~n26584;
  assign n26586 = ~n16031 & ~n26585;
  assign n26587 = ~i_RtoB_ACK0 & ~n26586;
  assign n26588 = ~n24655 & ~n26587;
  assign n26589 = controllable_DEQ & ~n26588;
  assign n26590 = ~n13771 & ~n19829;
  assign n26591 = ~controllable_BtoR_REQ0 & ~n26590;
  assign n26592 = ~n16050 & ~n26591;
  assign n26593 = ~i_RtoB_ACK0 & ~n26592;
  assign n26594 = ~n24661 & ~n26593;
  assign n26595 = ~controllable_DEQ & ~n26594;
  assign n26596 = ~n26589 & ~n26595;
  assign n26597 = i_FULL & ~n26596;
  assign n26598 = ~n13781 & ~n19839;
  assign n26599 = ~controllable_BtoR_REQ0 & ~n26598;
  assign n26600 = ~n16069 & ~n26599;
  assign n26601 = ~i_RtoB_ACK0 & ~n26600;
  assign n26602 = ~n24655 & ~n26601;
  assign n26603 = controllable_DEQ & ~n26602;
  assign n26604 = ~n13789 & ~n19847;
  assign n26605 = ~controllable_BtoR_REQ0 & ~n26604;
  assign n26606 = ~n16085 & ~n26605;
  assign n26607 = ~i_RtoB_ACK0 & ~n26606;
  assign n26608 = ~n24661 & ~n26607;
  assign n26609 = ~controllable_DEQ & ~n26608;
  assign n26610 = ~n26603 & ~n26609;
  assign n26611 = ~i_FULL & ~n26610;
  assign n26612 = ~n26597 & ~n26611;
  assign n26613 = i_nEMPTY & ~n26612;
  assign n26614 = ~n13802 & ~n19865;
  assign n26615 = ~controllable_BtoR_REQ0 & ~n26614;
  assign n26616 = ~n16122 & ~n26615;
  assign n26617 = ~i_RtoB_ACK0 & ~n26616;
  assign n26618 = ~n24681 & ~n26617;
  assign n26619 = ~controllable_DEQ & ~n26618;
  assign n26620 = ~n22725 & ~n26619;
  assign n26621 = i_FULL & ~n26620;
  assign n26622 = ~n13762 & ~n19881;
  assign n26623 = ~controllable_BtoR_REQ0 & ~n26622;
  assign n26624 = ~n16031 & ~n26623;
  assign n26625 = ~i_RtoB_ACK0 & ~n26624;
  assign n26626 = ~n24655 & ~n26625;
  assign n26627 = ~controllable_DEQ & ~n26626;
  assign n26628 = ~n22737 & ~n26627;
  assign n26629 = ~i_FULL & ~n26628;
  assign n26630 = ~n26621 & ~n26629;
  assign n26631 = ~i_nEMPTY & ~n26630;
  assign n26632 = ~n26613 & ~n26631;
  assign n26633 = ~controllable_BtoS_ACK0 & ~n26632;
  assign n26634 = ~n26583 & ~n26633;
  assign n26635 = n4465 & ~n26634;
  assign n26636 = ~n10719 & ~n11238;
  assign n26637 = ~controllable_BtoR_REQ0 & ~n26636;
  assign n26638 = ~n16175 & ~n26637;
  assign n26639 = ~i_RtoB_ACK0 & ~n26638;
  assign n26640 = ~n24701 & ~n26639;
  assign n26641 = controllable_DEQ & ~n26640;
  assign n26642 = ~n10736 & ~n11248;
  assign n26643 = ~controllable_BtoR_REQ0 & ~n26642;
  assign n26644 = ~n16194 & ~n26643;
  assign n26645 = ~i_RtoB_ACK0 & ~n26644;
  assign n26646 = ~n24707 & ~n26645;
  assign n26647 = ~controllable_DEQ & ~n26646;
  assign n26648 = ~n26641 & ~n26647;
  assign n26649 = i_nEMPTY & ~n26648;
  assign n26650 = ~n10752 & ~n11230;
  assign n26651 = ~controllable_BtoR_REQ0 & ~n26650;
  assign n26652 = ~n16220 & ~n26651;
  assign n26653 = ~i_RtoB_ACK0 & ~n26652;
  assign n26654 = ~n24715 & ~n26653;
  assign n26655 = ~controllable_DEQ & ~n26654;
  assign n26656 = ~n22767 & ~n26655;
  assign n26657 = i_FULL & ~n26656;
  assign n26658 = ~n10719 & ~n11284;
  assign n26659 = ~controllable_BtoR_REQ0 & ~n26658;
  assign n26660 = ~n16175 & ~n26659;
  assign n26661 = ~i_RtoB_ACK0 & ~n26660;
  assign n26662 = ~n24701 & ~n26661;
  assign n26663 = ~controllable_DEQ & ~n26662;
  assign n26664 = ~n22779 & ~n26663;
  assign n26665 = ~i_FULL & ~n26664;
  assign n26666 = ~n26657 & ~n26665;
  assign n26667 = ~i_nEMPTY & ~n26666;
  assign n26668 = ~n26649 & ~n26667;
  assign n26669 = controllable_BtoS_ACK0 & ~n26668;
  assign n26670 = ~n10790 & ~n19931;
  assign n26671 = ~controllable_BtoR_REQ0 & ~n26670;
  assign n26672 = ~n16262 & ~n26671;
  assign n26673 = ~i_RtoB_ACK0 & ~n26672;
  assign n26674 = ~n24733 & ~n26673;
  assign n26675 = controllable_DEQ & ~n26674;
  assign n26676 = ~n10622 & ~n19939;
  assign n26677 = ~controllable_BtoR_REQ0 & ~n26676;
  assign n26678 = ~n16281 & ~n26677;
  assign n26679 = ~i_RtoB_ACK0 & ~n26678;
  assign n26680 = ~n24739 & ~n26679;
  assign n26681 = ~controllable_DEQ & ~n26680;
  assign n26682 = ~n26675 & ~n26681;
  assign n26683 = i_FULL & ~n26682;
  assign n26684 = ~n10816 & ~n11317;
  assign n26685 = ~controllable_BtoR_REQ0 & ~n26684;
  assign n26686 = ~n16300 & ~n26685;
  assign n26687 = ~i_RtoB_ACK0 & ~n26686;
  assign n26688 = ~n24733 & ~n26687;
  assign n26689 = controllable_DEQ & ~n26688;
  assign n26690 = ~n10826 & ~n19953;
  assign n26691 = ~controllable_BtoR_REQ0 & ~n26690;
  assign n26692 = ~n16316 & ~n26691;
  assign n26693 = ~i_RtoB_ACK0 & ~n26692;
  assign n26694 = ~n24739 & ~n26693;
  assign n26695 = ~controllable_DEQ & ~n26694;
  assign n26696 = ~n26689 & ~n26695;
  assign n26697 = ~i_FULL & ~n26696;
  assign n26698 = ~n26683 & ~n26697;
  assign n26699 = i_nEMPTY & ~n26698;
  assign n26700 = ~n10673 & ~n19969;
  assign n26701 = ~controllable_BtoR_REQ0 & ~n26700;
  assign n26702 = ~n16353 & ~n26701;
  assign n26703 = ~i_RtoB_ACK0 & ~n26702;
  assign n26704 = ~n24759 & ~n26703;
  assign n26705 = ~controllable_DEQ & ~n26704;
  assign n26706 = ~n22819 & ~n26705;
  assign n26707 = i_FULL & ~n26706;
  assign n26708 = ~n10790 & ~n19983;
  assign n26709 = ~controllable_BtoR_REQ0 & ~n26708;
  assign n26710 = ~n16262 & ~n26709;
  assign n26711 = ~i_RtoB_ACK0 & ~n26710;
  assign n26712 = ~n24733 & ~n26711;
  assign n26713 = ~controllable_DEQ & ~n26712;
  assign n26714 = ~n22831 & ~n26713;
  assign n26715 = ~i_FULL & ~n26714;
  assign n26716 = ~n26707 & ~n26715;
  assign n26717 = ~i_nEMPTY & ~n26716;
  assign n26718 = ~n26699 & ~n26717;
  assign n26719 = ~controllable_BtoS_ACK0 & ~n26718;
  assign n26720 = ~n26669 & ~n26719;
  assign n26721 = ~n4465 & ~n26720;
  assign n26722 = ~n26635 & ~n26721;
  assign n26723 = ~i_StoB_REQ10 & ~n26722;
  assign n26724 = ~n26533 & ~n26723;
  assign n26725 = controllable_BtoS_ACK10 & ~n26724;
  assign n26726 = ~n10890 & ~n20004;
  assign n26727 = ~controllable_BtoR_REQ0 & ~n26726;
  assign n26728 = ~n20002 & ~n26727;
  assign n26729 = ~i_RtoB_ACK0 & ~n26728;
  assign n26730 = ~n24783 & ~n26729;
  assign n26731 = controllable_DEQ & ~n26730;
  assign n26732 = ~n10495 & ~n20013;
  assign n26733 = ~controllable_BtoR_REQ0 & ~n26732;
  assign n26734 = ~n20011 & ~n26733;
  assign n26735 = ~i_RtoB_ACK0 & ~n26734;
  assign n26736 = ~n24789 & ~n26735;
  assign n26737 = ~controllable_DEQ & ~n26736;
  assign n26738 = ~n26731 & ~n26737;
  assign n26739 = i_FULL & ~n26738;
  assign n26740 = ~n10910 & ~n11238;
  assign n26741 = ~controllable_BtoR_REQ0 & ~n26740;
  assign n26742 = ~n20022 & ~n26741;
  assign n26743 = ~i_RtoB_ACK0 & ~n26742;
  assign n26744 = ~n24783 & ~n26743;
  assign n26745 = controllable_DEQ & ~n26744;
  assign n26746 = ~n10520 & ~n20029;
  assign n26747 = ~controllable_BtoR_REQ0 & ~n26746;
  assign n26748 = ~n20027 & ~n26747;
  assign n26749 = ~i_RtoB_ACK0 & ~n26748;
  assign n26750 = ~n24789 & ~n26749;
  assign n26751 = ~controllable_DEQ & ~n26750;
  assign n26752 = ~n26745 & ~n26751;
  assign n26753 = ~i_FULL & ~n26752;
  assign n26754 = ~n26739 & ~n26753;
  assign n26755 = i_nEMPTY & ~n26754;
  assign n26756 = ~n10546 & ~n20047;
  assign n26757 = ~controllable_BtoR_REQ0 & ~n26756;
  assign n26758 = ~n20045 & ~n26757;
  assign n26759 = ~i_RtoB_ACK0 & ~n26758;
  assign n26760 = ~n24809 & ~n26759;
  assign n26761 = ~controllable_DEQ & ~n26760;
  assign n26762 = ~n22877 & ~n26761;
  assign n26763 = i_FULL & ~n26762;
  assign n26764 = ~controllable_DEQ & ~n26730;
  assign n26765 = ~n22889 & ~n26764;
  assign n26766 = ~i_FULL & ~n26765;
  assign n26767 = ~n26763 & ~n26766;
  assign n26768 = ~i_nEMPTY & ~n26767;
  assign n26769 = ~n26755 & ~n26768;
  assign n26770 = controllable_BtoS_ACK0 & ~n26769;
  assign n26771 = ~n10957 & ~n19931;
  assign n26772 = ~controllable_BtoR_REQ0 & ~n26771;
  assign n26773 = ~n20068 & ~n26772;
  assign n26774 = ~i_RtoB_ACK0 & ~n26773;
  assign n26775 = ~n24824 & ~n26774;
  assign n26776 = controllable_DEQ & ~n26775;
  assign n26777 = ~n20073 & ~n26677;
  assign n26778 = ~i_RtoB_ACK0 & ~n26777;
  assign n26779 = ~n24830 & ~n26778;
  assign n26780 = ~controllable_DEQ & ~n26779;
  assign n26781 = ~n26776 & ~n26780;
  assign n26782 = i_FULL & ~n26781;
  assign n26783 = ~n10977 & ~n11317;
  assign n26784 = ~controllable_BtoR_REQ0 & ~n26783;
  assign n26785 = ~n20080 & ~n26784;
  assign n26786 = ~i_RtoB_ACK0 & ~n26785;
  assign n26787 = ~n24824 & ~n26786;
  assign n26788 = controllable_DEQ & ~n26787;
  assign n26789 = ~n10647 & ~n19953;
  assign n26790 = ~controllable_BtoR_REQ0 & ~n26789;
  assign n26791 = ~n20085 & ~n26790;
  assign n26792 = ~i_RtoB_ACK0 & ~n26791;
  assign n26793 = ~n24830 & ~n26792;
  assign n26794 = ~controllable_DEQ & ~n26793;
  assign n26795 = ~n26788 & ~n26794;
  assign n26796 = ~i_FULL & ~n26795;
  assign n26797 = ~n26782 & ~n26796;
  assign n26798 = i_nEMPTY & ~n26797;
  assign n26799 = ~n20099 & ~n26701;
  assign n26800 = ~i_RtoB_ACK0 & ~n26799;
  assign n26801 = ~n24850 & ~n26800;
  assign n26802 = ~controllable_DEQ & ~n26801;
  assign n26803 = ~n22926 & ~n26802;
  assign n26804 = i_FULL & ~n26803;
  assign n26805 = ~controllable_DEQ & ~n26775;
  assign n26806 = ~n22938 & ~n26805;
  assign n26807 = ~i_FULL & ~n26806;
  assign n26808 = ~n26804 & ~n26807;
  assign n26809 = ~i_nEMPTY & ~n26808;
  assign n26810 = ~n26798 & ~n26809;
  assign n26811 = ~controllable_BtoS_ACK0 & ~n26810;
  assign n26812 = ~n26770 & ~n26811;
  assign n26813 = n4465 & ~n26812;
  assign n26814 = ~n11022 & ~n11238;
  assign n26815 = ~controllable_BtoR_REQ0 & ~n26814;
  assign n26816 = ~n20120 & ~n26815;
  assign n26817 = ~i_RtoB_ACK0 & ~n26816;
  assign n26818 = ~n24867 & ~n26817;
  assign n26819 = controllable_DEQ & ~n26818;
  assign n26820 = ~n20125 & ~n26643;
  assign n26821 = ~i_RtoB_ACK0 & ~n26820;
  assign n26822 = ~n24873 & ~n26821;
  assign n26823 = ~controllable_DEQ & ~n26822;
  assign n26824 = ~n26819 & ~n26823;
  assign n26825 = i_nEMPTY & ~n26824;
  assign n26826 = ~n20137 & ~n26651;
  assign n26827 = ~i_RtoB_ACK0 & ~n26826;
  assign n26828 = ~n24881 & ~n26827;
  assign n26829 = ~controllable_DEQ & ~n26828;
  assign n26830 = ~n22965 & ~n26829;
  assign n26831 = i_FULL & ~n26830;
  assign n26832 = ~controllable_DEQ & ~n26818;
  assign n26833 = ~n22977 & ~n26832;
  assign n26834 = ~i_FULL & ~n26833;
  assign n26835 = ~n26831 & ~n26834;
  assign n26836 = ~i_nEMPTY & ~n26835;
  assign n26837 = ~n26825 & ~n26836;
  assign n26838 = controllable_BtoS_ACK0 & ~n26837;
  assign n26839 = ~n11067 & ~n19931;
  assign n26840 = ~controllable_BtoR_REQ0 & ~n26839;
  assign n26841 = ~n20156 & ~n26840;
  assign n26842 = ~i_RtoB_ACK0 & ~n26841;
  assign n26843 = ~n24896 & ~n26842;
  assign n26844 = controllable_DEQ & ~n26843;
  assign n26845 = ~n20161 & ~n26677;
  assign n26846 = ~i_RtoB_ACK0 & ~n26845;
  assign n26847 = ~n24902 & ~n26846;
  assign n26848 = ~controllable_DEQ & ~n26847;
  assign n26849 = ~n26844 & ~n26848;
  assign n26850 = i_FULL & ~n26849;
  assign n26851 = ~n11083 & ~n11317;
  assign n26852 = ~controllable_BtoR_REQ0 & ~n26851;
  assign n26853 = ~n20168 & ~n26852;
  assign n26854 = ~i_RtoB_ACK0 & ~n26853;
  assign n26855 = ~n24896 & ~n26854;
  assign n26856 = controllable_DEQ & ~n26855;
  assign n26857 = ~n20173 & ~n26691;
  assign n26858 = ~i_RtoB_ACK0 & ~n26857;
  assign n26859 = ~n24902 & ~n26858;
  assign n26860 = ~controllable_DEQ & ~n26859;
  assign n26861 = ~n26856 & ~n26860;
  assign n26862 = ~i_FULL & ~n26861;
  assign n26863 = ~n26850 & ~n26862;
  assign n26864 = i_nEMPTY & ~n26863;
  assign n26865 = ~n20187 & ~n26701;
  assign n26866 = ~i_RtoB_ACK0 & ~n26865;
  assign n26867 = ~n24922 & ~n26866;
  assign n26868 = ~controllable_DEQ & ~n26867;
  assign n26869 = ~n23014 & ~n26868;
  assign n26870 = i_FULL & ~n26869;
  assign n26871 = ~controllable_DEQ & ~n26843;
  assign n26872 = ~n23026 & ~n26871;
  assign n26873 = ~i_FULL & ~n26872;
  assign n26874 = ~n26870 & ~n26873;
  assign n26875 = ~i_nEMPTY & ~n26874;
  assign n26876 = ~n26864 & ~n26875;
  assign n26877 = ~controllable_BtoS_ACK0 & ~n26876;
  assign n26878 = ~n26838 & ~n26877;
  assign n26879 = ~n4465 & ~n26878;
  assign n26880 = ~n26813 & ~n26879;
  assign n26881 = i_StoB_REQ10 & ~n26880;
  assign n26882 = ~n26723 & ~n26881;
  assign n26883 = ~controllable_BtoS_ACK10 & ~n26882;
  assign n26884 = ~n26725 & ~n26883;
  assign n26885 = ~n4464 & ~n26884;
  assign n26886 = ~n26431 & ~n26885;
  assign n26887 = n4463 & ~n26886;
  assign n26888 = ~n9306 & ~n19078;
  assign n26889 = ~controllable_BtoR_REQ0 & ~n26888;
  assign n26890 = ~n14904 & ~n26889;
  assign n26891 = ~i_RtoB_ACK0 & ~n26890;
  assign n26892 = ~n24219 & ~n26891;
  assign n26893 = controllable_DEQ & ~n26892;
  assign n26894 = ~n9519 & ~n19092;
  assign n26895 = ~controllable_BtoR_REQ0 & ~n26894;
  assign n26896 = ~n14923 & ~n26895;
  assign n26897 = ~i_RtoB_ACK0 & ~n26896;
  assign n26898 = ~n24225 & ~n26897;
  assign n26899 = ~controllable_DEQ & ~n26898;
  assign n26900 = ~n26893 & ~n26899;
  assign n26901 = i_FULL & ~n26900;
  assign n26902 = ~n9532 & ~n19102;
  assign n26903 = ~controllable_BtoR_REQ0 & ~n26902;
  assign n26904 = ~n14942 & ~n26903;
  assign n26905 = ~i_RtoB_ACK0 & ~n26904;
  assign n26906 = ~n24219 & ~n26905;
  assign n26907 = controllable_DEQ & ~n26906;
  assign n26908 = ~n9544 & ~n19110;
  assign n26909 = ~controllable_BtoR_REQ0 & ~n26908;
  assign n26910 = ~n14958 & ~n26909;
  assign n26911 = ~i_RtoB_ACK0 & ~n26910;
  assign n26912 = ~n24225 & ~n26911;
  assign n26913 = ~controllable_DEQ & ~n26912;
  assign n26914 = ~n26907 & ~n26913;
  assign n26915 = ~i_FULL & ~n26914;
  assign n26916 = ~n26901 & ~n26915;
  assign n26917 = i_nEMPTY & ~n26916;
  assign n26918 = ~n9573 & ~n19134;
  assign n26919 = ~controllable_BtoR_REQ0 & ~n26918;
  assign n26920 = ~n14995 & ~n26919;
  assign n26921 = ~i_RtoB_ACK0 & ~n26920;
  assign n26922 = ~n24245 & ~n26921;
  assign n26923 = ~controllable_DEQ & ~n26922;
  assign n26924 = ~n22169 & ~n26923;
  assign n26925 = i_FULL & ~n26924;
  assign n26926 = ~n9306 & ~n19150;
  assign n26927 = ~controllable_BtoR_REQ0 & ~n26926;
  assign n26928 = ~n14904 & ~n26927;
  assign n26929 = ~i_RtoB_ACK0 & ~n26928;
  assign n26930 = ~n24219 & ~n26929;
  assign n26931 = ~controllable_DEQ & ~n26930;
  assign n26932 = ~n22181 & ~n26931;
  assign n26933 = ~i_FULL & ~n26932;
  assign n26934 = ~n26925 & ~n26933;
  assign n26935 = ~i_nEMPTY & ~n26934;
  assign n26936 = ~n26917 & ~n26935;
  assign n26937 = controllable_BtoS_ACK0 & ~n26936;
  assign n26938 = ~n9639 & ~n19171;
  assign n26939 = ~controllable_BtoR_REQ0 & ~n26938;
  assign n26940 = ~n15046 & ~n26939;
  assign n26941 = ~i_RtoB_ACK0 & ~n26940;
  assign n26942 = ~n24263 & ~n26941;
  assign n26943 = controllable_DEQ & ~n26942;
  assign n26944 = ~n9666 & ~n19185;
  assign n26945 = ~controllable_BtoR_REQ0 & ~n26944;
  assign n26946 = ~n15065 & ~n26945;
  assign n26947 = ~i_RtoB_ACK0 & ~n26946;
  assign n26948 = ~n24269 & ~n26947;
  assign n26949 = ~controllable_DEQ & ~n26948;
  assign n26950 = ~n26943 & ~n26949;
  assign n26951 = i_FULL & ~n26950;
  assign n26952 = ~n9679 & ~n19195;
  assign n26953 = ~controllable_BtoR_REQ0 & ~n26952;
  assign n26954 = ~n15084 & ~n26953;
  assign n26955 = ~i_RtoB_ACK0 & ~n26954;
  assign n26956 = ~n24263 & ~n26955;
  assign n26957 = controllable_DEQ & ~n26956;
  assign n26958 = ~n9691 & ~n19203;
  assign n26959 = ~controllable_BtoR_REQ0 & ~n26958;
  assign n26960 = ~n15100 & ~n26959;
  assign n26961 = ~i_RtoB_ACK0 & ~n26960;
  assign n26962 = ~n24269 & ~n26961;
  assign n26963 = ~controllable_DEQ & ~n26962;
  assign n26964 = ~n26957 & ~n26963;
  assign n26965 = ~i_FULL & ~n26964;
  assign n26966 = ~n26951 & ~n26965;
  assign n26967 = i_nEMPTY & ~n26966;
  assign n26968 = ~n9720 & ~n19227;
  assign n26969 = ~controllable_BtoR_REQ0 & ~n26968;
  assign n26970 = ~n15137 & ~n26969;
  assign n26971 = ~i_RtoB_ACK0 & ~n26970;
  assign n26972 = ~n24289 & ~n26971;
  assign n26973 = ~controllable_DEQ & ~n26972;
  assign n26974 = ~n22221 & ~n26973;
  assign n26975 = i_FULL & ~n26974;
  assign n26976 = ~n9639 & ~n19243;
  assign n26977 = ~controllable_BtoR_REQ0 & ~n26976;
  assign n26978 = ~n15046 & ~n26977;
  assign n26979 = ~i_RtoB_ACK0 & ~n26978;
  assign n26980 = ~n24263 & ~n26979;
  assign n26981 = ~controllable_DEQ & ~n26980;
  assign n26982 = ~n22233 & ~n26981;
  assign n26983 = ~i_FULL & ~n26982;
  assign n26984 = ~n26975 & ~n26983;
  assign n26985 = ~i_nEMPTY & ~n26984;
  assign n26986 = ~n26967 & ~n26985;
  assign n26987 = ~controllable_BtoS_ACK0 & ~n26986;
  assign n26988 = ~n26937 & ~n26987;
  assign n26989 = n4465 & ~n26988;
  assign n26990 = ~n9791 & ~n19259;
  assign n26991 = ~controllable_BtoR_REQ0 & ~n26990;
  assign n26992 = ~n15190 & ~n26991;
  assign n26993 = ~i_RtoB_ACK0 & ~n26992;
  assign n26994 = ~n24309 & ~n26993;
  assign n26995 = controllable_DEQ & ~n26994;
  assign n26996 = ~n9812 & ~n19267;
  assign n26997 = ~controllable_BtoR_REQ0 & ~n26996;
  assign n26998 = ~n15209 & ~n26997;
  assign n26999 = ~i_RtoB_ACK0 & ~n26998;
  assign n27000 = ~n24315 & ~n26999;
  assign n27001 = ~controllable_DEQ & ~n27000;
  assign n27002 = ~n26995 & ~n27001;
  assign n27003 = i_nEMPTY & ~n27002;
  assign n27004 = ~n9835 & ~n19283;
  assign n27005 = ~controllable_BtoR_REQ0 & ~n27004;
  assign n27006 = ~n15237 & ~n27005;
  assign n27007 = ~i_RtoB_ACK0 & ~n27006;
  assign n27008 = ~n24323 & ~n27007;
  assign n27009 = ~controllable_DEQ & ~n27008;
  assign n27010 = ~n22263 & ~n27009;
  assign n27011 = i_FULL & ~n27010;
  assign n27012 = ~n9791 & ~n19299;
  assign n27013 = ~controllable_BtoR_REQ0 & ~n27012;
  assign n27014 = ~n15190 & ~n27013;
  assign n27015 = ~i_RtoB_ACK0 & ~n27014;
  assign n27016 = ~n24309 & ~n27015;
  assign n27017 = ~controllable_DEQ & ~n27016;
  assign n27018 = ~n22275 & ~n27017;
  assign n27019 = ~i_FULL & ~n27018;
  assign n27020 = ~n27011 & ~n27019;
  assign n27021 = ~i_nEMPTY & ~n27020;
  assign n27022 = ~n27003 & ~n27021;
  assign n27023 = controllable_BtoS_ACK0 & ~n27022;
  assign n27024 = ~n26257 & ~n27023;
  assign n27025 = ~n4465 & ~n27024;
  assign n27026 = ~n26989 & ~n27025;
  assign n27027 = ~i_StoB_REQ10 & ~n27026;
  assign n27028 = ~n26071 & ~n27027;
  assign n27029 = controllable_BtoS_ACK10 & ~n27028;
  assign n27030 = ~n26427 & ~n27027;
  assign n27031 = ~controllable_BtoS_ACK10 & ~n27030;
  assign n27032 = ~n27029 & ~n27031;
  assign n27033 = n4464 & ~n27032;
  assign n27034 = ~n10470 & ~n19747;
  assign n27035 = ~controllable_BtoR_REQ0 & ~n27034;
  assign n27036 = ~n15889 & ~n27035;
  assign n27037 = ~i_RtoB_ACK0 & ~n27036;
  assign n27038 = ~n24611 & ~n27037;
  assign n27039 = controllable_DEQ & ~n27038;
  assign n27040 = ~n10495 & ~n19755;
  assign n27041 = ~controllable_BtoR_REQ0 & ~n27040;
  assign n27042 = ~n15908 & ~n27041;
  assign n27043 = ~i_RtoB_ACK0 & ~n27042;
  assign n27044 = ~n24617 & ~n27043;
  assign n27045 = ~controllable_DEQ & ~n27044;
  assign n27046 = ~n27039 & ~n27045;
  assign n27047 = i_FULL & ~n27046;
  assign n27048 = ~n10508 & ~n19765;
  assign n27049 = ~controllable_BtoR_REQ0 & ~n27048;
  assign n27050 = ~n15927 & ~n27049;
  assign n27051 = ~i_RtoB_ACK0 & ~n27050;
  assign n27052 = ~n24611 & ~n27051;
  assign n27053 = controllable_DEQ & ~n27052;
  assign n27054 = ~n10520 & ~n19773;
  assign n27055 = ~controllable_BtoR_REQ0 & ~n27054;
  assign n27056 = ~n15943 & ~n27055;
  assign n27057 = ~i_RtoB_ACK0 & ~n27056;
  assign n27058 = ~n24617 & ~n27057;
  assign n27059 = ~controllable_DEQ & ~n27058;
  assign n27060 = ~n27053 & ~n27059;
  assign n27061 = ~i_FULL & ~n27060;
  assign n27062 = ~n27047 & ~n27061;
  assign n27063 = i_nEMPTY & ~n27062;
  assign n27064 = ~n10546 & ~n19791;
  assign n27065 = ~controllable_BtoR_REQ0 & ~n27064;
  assign n27066 = ~n15980 & ~n27065;
  assign n27067 = ~i_RtoB_ACK0 & ~n27066;
  assign n27068 = ~n24637 & ~n27067;
  assign n27069 = ~controllable_DEQ & ~n27068;
  assign n27070 = ~n22673 & ~n27069;
  assign n27071 = i_FULL & ~n27070;
  assign n27072 = ~n10470 & ~n19807;
  assign n27073 = ~controllable_BtoR_REQ0 & ~n27072;
  assign n27074 = ~n15889 & ~n27073;
  assign n27075 = ~i_RtoB_ACK0 & ~n27074;
  assign n27076 = ~n24611 & ~n27075;
  assign n27077 = ~controllable_DEQ & ~n27076;
  assign n27078 = ~n22685 & ~n27077;
  assign n27079 = ~i_FULL & ~n27078;
  assign n27080 = ~n27071 & ~n27079;
  assign n27081 = ~i_nEMPTY & ~n27080;
  assign n27082 = ~n27063 & ~n27081;
  assign n27083 = controllable_BtoS_ACK0 & ~n27082;
  assign n27084 = ~n10600 & ~n19821;
  assign n27085 = ~controllable_BtoR_REQ0 & ~n27084;
  assign n27086 = ~n16031 & ~n27085;
  assign n27087 = ~i_RtoB_ACK0 & ~n27086;
  assign n27088 = ~n24655 & ~n27087;
  assign n27089 = controllable_DEQ & ~n27088;
  assign n27090 = ~n10622 & ~n19829;
  assign n27091 = ~controllable_BtoR_REQ0 & ~n27090;
  assign n27092 = ~n16050 & ~n27091;
  assign n27093 = ~i_RtoB_ACK0 & ~n27092;
  assign n27094 = ~n24661 & ~n27093;
  assign n27095 = ~controllable_DEQ & ~n27094;
  assign n27096 = ~n27089 & ~n27095;
  assign n27097 = i_FULL & ~n27096;
  assign n27098 = ~n10635 & ~n19839;
  assign n27099 = ~controllable_BtoR_REQ0 & ~n27098;
  assign n27100 = ~n16069 & ~n27099;
  assign n27101 = ~i_RtoB_ACK0 & ~n27100;
  assign n27102 = ~n24655 & ~n27101;
  assign n27103 = controllable_DEQ & ~n27102;
  assign n27104 = ~n10647 & ~n19847;
  assign n27105 = ~controllable_BtoR_REQ0 & ~n27104;
  assign n27106 = ~n16085 & ~n27105;
  assign n27107 = ~i_RtoB_ACK0 & ~n27106;
  assign n27108 = ~n24661 & ~n27107;
  assign n27109 = ~controllable_DEQ & ~n27108;
  assign n27110 = ~n27103 & ~n27109;
  assign n27111 = ~i_FULL & ~n27110;
  assign n27112 = ~n27097 & ~n27111;
  assign n27113 = i_nEMPTY & ~n27112;
  assign n27114 = ~n10673 & ~n19865;
  assign n27115 = ~controllable_BtoR_REQ0 & ~n27114;
  assign n27116 = ~n16122 & ~n27115;
  assign n27117 = ~i_RtoB_ACK0 & ~n27116;
  assign n27118 = ~n24681 & ~n27117;
  assign n27119 = ~controllable_DEQ & ~n27118;
  assign n27120 = ~n22725 & ~n27119;
  assign n27121 = i_FULL & ~n27120;
  assign n27122 = ~n10600 & ~n19881;
  assign n27123 = ~controllable_BtoR_REQ0 & ~n27122;
  assign n27124 = ~n16031 & ~n27123;
  assign n27125 = ~i_RtoB_ACK0 & ~n27124;
  assign n27126 = ~n24655 & ~n27125;
  assign n27127 = ~controllable_DEQ & ~n27126;
  assign n27128 = ~n22737 & ~n27127;
  assign n27129 = ~i_FULL & ~n27128;
  assign n27130 = ~n27121 & ~n27129;
  assign n27131 = ~i_nEMPTY & ~n27130;
  assign n27132 = ~n27113 & ~n27131;
  assign n27133 = ~controllable_BtoS_ACK0 & ~n27132;
  assign n27134 = ~n27083 & ~n27133;
  assign n27135 = n4465 & ~n27134;
  assign n27136 = ~n26721 & ~n27135;
  assign n27137 = ~i_StoB_REQ10 & ~n27136;
  assign n27138 = ~n26533 & ~n27137;
  assign n27139 = controllable_BtoS_ACK10 & ~n27138;
  assign n27140 = ~n26881 & ~n27137;
  assign n27141 = ~controllable_BtoS_ACK10 & ~n27140;
  assign n27142 = ~n27139 & ~n27141;
  assign n27143 = ~n4464 & ~n27142;
  assign n27144 = ~n27033 & ~n27143;
  assign n27145 = ~n4463 & ~n27144;
  assign n27146 = ~n26887 & ~n27145;
  assign n27147 = n4462 & ~n27146;
  assign n27148 = ~n14075 & ~n20219;
  assign n27149 = ~controllable_BtoR_REQ0 & ~n27148;
  assign n27150 = ~n17545 & ~n27149;
  assign n27151 = ~i_RtoB_ACK0 & ~n27150;
  assign n27152 = ~n25125 & ~n27151;
  assign n27153 = controllable_DEQ & ~n27152;
  assign n27154 = ~n14084 & ~n20229;
  assign n27155 = ~controllable_BtoR_REQ0 & ~n27154;
  assign n27156 = ~n17562 & ~n27155;
  assign n27157 = ~i_RtoB_ACK0 & ~n27156;
  assign n27158 = ~n25131 & ~n27157;
  assign n27159 = ~controllable_DEQ & ~n27158;
  assign n27160 = ~n27153 & ~n27159;
  assign n27161 = i_nEMPTY & ~n27160;
  assign n27162 = ~n14094 & ~n20245;
  assign n27163 = ~controllable_BtoR_REQ0 & ~n27162;
  assign n27164 = ~n17581 & ~n27163;
  assign n27165 = ~i_RtoB_ACK0 & ~n27164;
  assign n27166 = ~n25125 & ~n27165;
  assign n27167 = ~controllable_DEQ & ~n27166;
  assign n27168 = ~n23541 & ~n27167;
  assign n27169 = i_FULL & ~n27168;
  assign n27170 = ~n14075 & ~n20260;
  assign n27171 = ~controllable_BtoR_REQ0 & ~n27170;
  assign n27172 = ~n17545 & ~n27171;
  assign n27173 = ~i_RtoB_ACK0 & ~n27172;
  assign n27174 = ~n25125 & ~n27173;
  assign n27175 = ~controllable_DEQ & ~n27174;
  assign n27176 = ~n23551 & ~n27175;
  assign n27177 = ~i_FULL & ~n27176;
  assign n27178 = ~n27169 & ~n27177;
  assign n27179 = ~i_nEMPTY & ~n27178;
  assign n27180 = ~n27161 & ~n27179;
  assign n27181 = controllable_BtoS_ACK0 & ~n27180;
  assign n27182 = ~n14118 & ~n20274;
  assign n27183 = ~controllable_BtoR_REQ0 & ~n27182;
  assign n27184 = ~n14824 & ~n27183;
  assign n27185 = ~i_RtoB_ACK0 & ~n27184;
  assign n27186 = ~n24189 & ~n27185;
  assign n27187 = controllable_DEQ & ~n27186;
  assign n27188 = ~n14127 & ~n20282;
  assign n27189 = ~controllable_BtoR_REQ0 & ~n27188;
  assign n27190 = ~n14841 & ~n27189;
  assign n27191 = ~i_RtoB_ACK0 & ~n27190;
  assign n27192 = ~n24195 & ~n27191;
  assign n27193 = ~controllable_DEQ & ~n27192;
  assign n27194 = ~n27187 & ~n27193;
  assign n27195 = i_nEMPTY & ~n27194;
  assign n27196 = ~n14137 & ~n20298;
  assign n27197 = ~controllable_BtoR_REQ0 & ~n27196;
  assign n27198 = ~n14860 & ~n27197;
  assign n27199 = ~i_RtoB_ACK0 & ~n27198;
  assign n27200 = ~n24189 & ~n27199;
  assign n27201 = ~controllable_DEQ & ~n27200;
  assign n27202 = ~n23579 & ~n27201;
  assign n27203 = i_FULL & ~n27202;
  assign n27204 = ~n14118 & ~n20313;
  assign n27205 = ~controllable_BtoR_REQ0 & ~n27204;
  assign n27206 = ~n14824 & ~n27205;
  assign n27207 = ~i_RtoB_ACK0 & ~n27206;
  assign n27208 = ~n24189 & ~n27207;
  assign n27209 = ~controllable_DEQ & ~n27208;
  assign n27210 = ~n23589 & ~n27209;
  assign n27211 = ~i_FULL & ~n27210;
  assign n27212 = ~n27203 & ~n27211;
  assign n27213 = ~i_nEMPTY & ~n27212;
  assign n27214 = ~n27195 & ~n27213;
  assign n27215 = ~controllable_BtoS_ACK0 & ~n27214;
  assign n27216 = ~n27181 & ~n27215;
  assign n27217 = n4465 & ~n27216;
  assign n27218 = ~n8991 & ~n20328;
  assign n27219 = ~controllable_BtoR_REQ0 & ~n27218;
  assign n27220 = ~n14841 & ~n27219;
  assign n27221 = ~i_RtoB_ACK0 & ~n27220;
  assign n27222 = ~n24195 & ~n27221;
  assign n27223 = ~controllable_DEQ & ~n27222;
  assign n27224 = ~n26038 & ~n27223;
  assign n27225 = i_nEMPTY & ~n27224;
  assign n27226 = ~n9028 & ~n20337;
  assign n27227 = ~controllable_BtoR_REQ0 & ~n27226;
  assign n27228 = ~n14860 & ~n27227;
  assign n27229 = ~i_RtoB_ACK0 & ~n27228;
  assign n27230 = ~n24189 & ~n27229;
  assign n27231 = ~controllable_DEQ & ~n27230;
  assign n27232 = ~n22115 & ~n27231;
  assign n27233 = i_FULL & ~n27232;
  assign n27234 = ~n8972 & ~n20347;
  assign n27235 = ~controllable_BtoR_REQ0 & ~n27234;
  assign n27236 = ~n14824 & ~n27235;
  assign n27237 = ~i_RtoB_ACK0 & ~n27236;
  assign n27238 = ~n24189 & ~n27237;
  assign n27239 = ~controllable_DEQ & ~n27238;
  assign n27240 = ~n22125 & ~n27239;
  assign n27241 = ~i_FULL & ~n27240;
  assign n27242 = ~n27233 & ~n27241;
  assign n27243 = ~i_nEMPTY & ~n27242;
  assign n27244 = ~n27225 & ~n27243;
  assign n27245 = ~controllable_BtoS_ACK0 & ~n27244;
  assign n27246 = ~n21013 & ~n27245;
  assign n27247 = ~n4465 & ~n27246;
  assign n27248 = ~n27217 & ~n27247;
  assign n27249 = i_StoB_REQ10 & ~n27248;
  assign n27250 = ~n23169 & ~n27249;
  assign n27251 = controllable_BtoS_ACK10 & ~n27250;
  assign n27252 = ~n12363 & ~n20368;
  assign n27253 = ~controllable_BtoR_REQ0 & ~n27252;
  assign n27254 = ~n20366 & ~n27253;
  assign n27255 = ~i_RtoB_ACK0 & ~n27254;
  assign n27256 = ~n25187 & ~n27255;
  assign n27257 = controllable_DEQ & ~n27256;
  assign n27258 = ~n12386 & ~n20377;
  assign n27259 = ~controllable_BtoR_REQ0 & ~n27258;
  assign n27260 = ~n20375 & ~n27259;
  assign n27261 = ~i_RtoB_ACK0 & ~n27260;
  assign n27262 = ~n25193 & ~n27261;
  assign n27263 = ~controllable_DEQ & ~n27262;
  assign n27264 = ~n27257 & ~n27263;
  assign n27265 = i_FULL & ~n27264;
  assign n27266 = ~n11238 & ~n12399;
  assign n27267 = ~controllable_BtoR_REQ0 & ~n27266;
  assign n27268 = ~n20386 & ~n27267;
  assign n27269 = ~i_RtoB_ACK0 & ~n27268;
  assign n27270 = ~n25187 & ~n27269;
  assign n27271 = controllable_DEQ & ~n27270;
  assign n27272 = ~n12409 & ~n20393;
  assign n27273 = ~controllable_BtoR_REQ0 & ~n27272;
  assign n27274 = ~n20391 & ~n27273;
  assign n27275 = ~i_RtoB_ACK0 & ~n27274;
  assign n27276 = ~n25193 & ~n27275;
  assign n27277 = ~controllable_DEQ & ~n27276;
  assign n27278 = ~n27271 & ~n27277;
  assign n27279 = ~i_FULL & ~n27278;
  assign n27280 = ~n27265 & ~n27279;
  assign n27281 = i_nEMPTY & ~n27280;
  assign n27282 = ~n12429 & ~n20411;
  assign n27283 = ~controllable_BtoR_REQ0 & ~n27282;
  assign n27284 = ~n20409 & ~n27283;
  assign n27285 = ~i_RtoB_ACK0 & ~n27284;
  assign n27286 = ~n25213 & ~n27285;
  assign n27287 = ~controllable_DEQ & ~n27286;
  assign n27288 = ~n23653 & ~n27287;
  assign n27289 = i_FULL & ~n27288;
  assign n27290 = ~controllable_DEQ & ~n27256;
  assign n27291 = ~n23665 & ~n27290;
  assign n27292 = ~i_FULL & ~n27291;
  assign n27293 = ~n27289 & ~n27292;
  assign n27294 = ~i_nEMPTY & ~n27293;
  assign n27295 = ~n27281 & ~n27294;
  assign n27296 = controllable_BtoS_ACK0 & ~n27295;
  assign n27297 = ~n12464 & ~n19313;
  assign n27298 = ~controllable_BtoR_REQ0 & ~n27297;
  assign n27299 = ~n20432 & ~n27298;
  assign n27300 = ~i_RtoB_ACK0 & ~n27299;
  assign n27301 = ~n25228 & ~n27300;
  assign n27302 = controllable_DEQ & ~n27301;
  assign n27303 = ~n20437 & ~n26215;
  assign n27304 = ~i_RtoB_ACK0 & ~n27303;
  assign n27305 = ~n25234 & ~n27304;
  assign n27306 = ~controllable_DEQ & ~n27305;
  assign n27307 = ~n27302 & ~n27306;
  assign n27308 = i_FULL & ~n27307;
  assign n27309 = ~n11317 & ~n12490;
  assign n27310 = ~controllable_BtoR_REQ0 & ~n27309;
  assign n27311 = ~n20444 & ~n27310;
  assign n27312 = ~i_RtoB_ACK0 & ~n27311;
  assign n27313 = ~n25228 & ~n27312;
  assign n27314 = controllable_DEQ & ~n27313;
  assign n27315 = ~n12500 & ~n19335;
  assign n27316 = ~controllable_BtoR_REQ0 & ~n27315;
  assign n27317 = ~n20449 & ~n27316;
  assign n27318 = ~i_RtoB_ACK0 & ~n27317;
  assign n27319 = ~n25234 & ~n27318;
  assign n27320 = ~controllable_DEQ & ~n27319;
  assign n27321 = ~n27314 & ~n27320;
  assign n27322 = ~i_FULL & ~n27321;
  assign n27323 = ~n27308 & ~n27322;
  assign n27324 = i_nEMPTY & ~n27323;
  assign n27325 = ~n20463 & ~n26239;
  assign n27326 = ~i_RtoB_ACK0 & ~n27325;
  assign n27327 = ~n25254 & ~n27326;
  assign n27328 = ~controllable_DEQ & ~n27327;
  assign n27329 = ~n23702 & ~n27328;
  assign n27330 = i_FULL & ~n27329;
  assign n27331 = ~controllable_DEQ & ~n27301;
  assign n27332 = ~n23714 & ~n27331;
  assign n27333 = ~i_FULL & ~n27332;
  assign n27334 = ~n27330 & ~n27333;
  assign n27335 = ~i_nEMPTY & ~n27334;
  assign n27336 = ~n27324 & ~n27335;
  assign n27337 = ~controllable_BtoS_ACK0 & ~n27336;
  assign n27338 = ~n27296 & ~n27337;
  assign n27339 = n4465 & ~n27338;
  assign n27340 = ~n26384 & ~n27337;
  assign n27341 = ~n4465 & ~n27340;
  assign n27342 = ~n27339 & ~n27341;
  assign n27343 = i_StoB_REQ10 & ~n27342;
  assign n27344 = ~n12557 & ~n20368;
  assign n27345 = ~controllable_BtoR_REQ0 & ~n27344;
  assign n27346 = ~n17974 & ~n27345;
  assign n27347 = ~i_RtoB_ACK0 & ~n27346;
  assign n27348 = ~n25275 & ~n27347;
  assign n27349 = controllable_DEQ & ~n27348;
  assign n27350 = ~n17993 & ~n27259;
  assign n27351 = ~i_RtoB_ACK0 & ~n27350;
  assign n27352 = ~n25281 & ~n27351;
  assign n27353 = ~controllable_DEQ & ~n27352;
  assign n27354 = ~n27349 & ~n27353;
  assign n27355 = i_FULL & ~n27354;
  assign n27356 = ~n11238 & ~n12583;
  assign n27357 = ~controllable_BtoR_REQ0 & ~n27356;
  assign n27358 = ~n18012 & ~n27357;
  assign n27359 = ~i_RtoB_ACK0 & ~n27358;
  assign n27360 = ~n25275 & ~n27359;
  assign n27361 = controllable_DEQ & ~n27360;
  assign n27362 = ~n12593 & ~n20393;
  assign n27363 = ~controllable_BtoR_REQ0 & ~n27362;
  assign n27364 = ~n18028 & ~n27363;
  assign n27365 = ~i_RtoB_ACK0 & ~n27364;
  assign n27366 = ~n25281 & ~n27365;
  assign n27367 = ~controllable_DEQ & ~n27366;
  assign n27368 = ~n27361 & ~n27367;
  assign n27369 = ~i_FULL & ~n27368;
  assign n27370 = ~n27355 & ~n27369;
  assign n27371 = i_nEMPTY & ~n27370;
  assign n27372 = ~n18065 & ~n27283;
  assign n27373 = ~i_RtoB_ACK0 & ~n27372;
  assign n27374 = ~n25301 & ~n27373;
  assign n27375 = ~controllable_DEQ & ~n27374;
  assign n27376 = ~n23757 & ~n27375;
  assign n27377 = i_FULL & ~n27376;
  assign n27378 = ~n12557 & ~n20525;
  assign n27379 = ~controllable_BtoR_REQ0 & ~n27378;
  assign n27380 = ~n17974 & ~n27379;
  assign n27381 = ~i_RtoB_ACK0 & ~n27380;
  assign n27382 = ~n25275 & ~n27381;
  assign n27383 = ~controllable_DEQ & ~n27382;
  assign n27384 = ~n23769 & ~n27383;
  assign n27385 = ~i_FULL & ~n27384;
  assign n27386 = ~n27377 & ~n27385;
  assign n27387 = ~i_nEMPTY & ~n27386;
  assign n27388 = ~n27371 & ~n27387;
  assign n27389 = controllable_BtoS_ACK0 & ~n27388;
  assign n27390 = ~n12653 & ~n19313;
  assign n27391 = ~controllable_BtoR_REQ0 & ~n27390;
  assign n27392 = ~n18116 & ~n27391;
  assign n27393 = ~i_RtoB_ACK0 & ~n27392;
  assign n27394 = ~n25319 & ~n27393;
  assign n27395 = controllable_DEQ & ~n27394;
  assign n27396 = ~n18135 & ~n26215;
  assign n27397 = ~i_RtoB_ACK0 & ~n27396;
  assign n27398 = ~n25325 & ~n27397;
  assign n27399 = ~controllable_DEQ & ~n27398;
  assign n27400 = ~n27395 & ~n27399;
  assign n27401 = i_FULL & ~n27400;
  assign n27402 = ~n11317 & ~n12679;
  assign n27403 = ~controllable_BtoR_REQ0 & ~n27402;
  assign n27404 = ~n18154 & ~n27403;
  assign n27405 = ~i_RtoB_ACK0 & ~n27404;
  assign n27406 = ~n25319 & ~n27405;
  assign n27407 = controllable_DEQ & ~n27406;
  assign n27408 = ~n12689 & ~n19335;
  assign n27409 = ~controllable_BtoR_REQ0 & ~n27408;
  assign n27410 = ~n18170 & ~n27409;
  assign n27411 = ~i_RtoB_ACK0 & ~n27410;
  assign n27412 = ~n25325 & ~n27411;
  assign n27413 = ~controllable_DEQ & ~n27412;
  assign n27414 = ~n27407 & ~n27413;
  assign n27415 = ~i_FULL & ~n27414;
  assign n27416 = ~n27401 & ~n27415;
  assign n27417 = i_nEMPTY & ~n27416;
  assign n27418 = ~n18207 & ~n26239;
  assign n27419 = ~i_RtoB_ACK0 & ~n27418;
  assign n27420 = ~n25345 & ~n27419;
  assign n27421 = ~controllable_DEQ & ~n27420;
  assign n27422 = ~n23809 & ~n27421;
  assign n27423 = i_FULL & ~n27422;
  assign n27424 = ~n12653 & ~n19365;
  assign n27425 = ~controllable_BtoR_REQ0 & ~n27424;
  assign n27426 = ~n18116 & ~n27425;
  assign n27427 = ~i_RtoB_ACK0 & ~n27426;
  assign n27428 = ~n25319 & ~n27427;
  assign n27429 = ~controllable_DEQ & ~n27428;
  assign n27430 = ~n23821 & ~n27429;
  assign n27431 = ~i_FULL & ~n27430;
  assign n27432 = ~n27423 & ~n27431;
  assign n27433 = ~i_nEMPTY & ~n27432;
  assign n27434 = ~n27417 & ~n27433;
  assign n27435 = ~controllable_BtoS_ACK0 & ~n27434;
  assign n27436 = ~n27389 & ~n27435;
  assign n27437 = n4465 & ~n27436;
  assign n27438 = ~n9791 & ~n11238;
  assign n27439 = ~controllable_BtoR_REQ0 & ~n27438;
  assign n27440 = ~n15190 & ~n27439;
  assign n27441 = ~i_RtoB_ACK0 & ~n27440;
  assign n27442 = ~n24309 & ~n27441;
  assign n27443 = controllable_DEQ & ~n27442;
  assign n27444 = ~n15209 & ~n26363;
  assign n27445 = ~i_RtoB_ACK0 & ~n27444;
  assign n27446 = ~n24315 & ~n27445;
  assign n27447 = ~controllable_DEQ & ~n27446;
  assign n27448 = ~n27443 & ~n27447;
  assign n27449 = i_nEMPTY & ~n27448;
  assign n27450 = ~n15237 & ~n26371;
  assign n27451 = ~i_RtoB_ACK0 & ~n27450;
  assign n27452 = ~n24323 & ~n27451;
  assign n27453 = ~controllable_DEQ & ~n27452;
  assign n27454 = ~n23849 & ~n27453;
  assign n27455 = i_FULL & ~n27454;
  assign n27456 = ~n9791 & ~n11284;
  assign n27457 = ~controllable_BtoR_REQ0 & ~n27456;
  assign n27458 = ~n15190 & ~n27457;
  assign n27459 = ~i_RtoB_ACK0 & ~n27458;
  assign n27460 = ~n24309 & ~n27459;
  assign n27461 = ~controllable_DEQ & ~n27460;
  assign n27462 = ~n23859 & ~n27461;
  assign n27463 = ~i_FULL & ~n27462;
  assign n27464 = ~n27455 & ~n27463;
  assign n27465 = ~i_nEMPTY & ~n27464;
  assign n27466 = ~n27449 & ~n27465;
  assign n27467 = controllable_BtoS_ACK0 & ~n27466;
  assign n27468 = ~n26257 & ~n27467;
  assign n27469 = ~n4465 & ~n27468;
  assign n27470 = ~n27437 & ~n27469;
  assign n27471 = ~i_StoB_REQ10 & ~n27470;
  assign n27472 = ~n27343 & ~n27471;
  assign n27473 = ~controllable_BtoS_ACK10 & ~n27472;
  assign n27474 = ~n27251 & ~n27473;
  assign n27475 = n4464 & ~n27474;
  assign n27476 = ~n5255 & ~n10284;
  assign n27477 = ~controllable_BtoR_REQ0 & ~n27476;
  assign n27478 = ~n15749 & ~n27477;
  assign n27479 = ~i_RtoB_ACK0 & ~n27478;
  assign n27480 = ~n24559 & ~n27479;
  assign n27481 = ~controllable_DEQ & ~n27480;
  assign n27482 = ~n26450 & ~n27481;
  assign n27483 = i_nEMPTY & ~n27482;
  assign n27484 = ~n5232 & ~n10321;
  assign n27485 = ~controllable_BtoR_REQ0 & ~n27484;
  assign n27486 = ~n15768 & ~n27485;
  assign n27487 = ~i_RtoB_ACK0 & ~n27486;
  assign n27488 = ~n24553 & ~n27487;
  assign n27489 = ~controllable_DEQ & ~n27488;
  assign n27490 = ~n22567 & ~n27489;
  assign n27491 = i_FULL & ~n27490;
  assign n27492 = ~n10265 & ~n14799;
  assign n27493 = ~controllable_BtoR_REQ0 & ~n27492;
  assign n27494 = ~n15732 & ~n27493;
  assign n27495 = ~i_RtoB_ACK0 & ~n27494;
  assign n27496 = ~n24553 & ~n27495;
  assign n27497 = ~controllable_DEQ & ~n27496;
  assign n27498 = ~n22577 & ~n27497;
  assign n27499 = ~i_FULL & ~n27498;
  assign n27500 = ~n27491 & ~n27499;
  assign n27501 = ~i_nEMPTY & ~n27500;
  assign n27502 = ~n27483 & ~n27501;
  assign n27503 = controllable_BtoS_ACK0 & ~n27502;
  assign n27504 = ~n10378 & ~n20328;
  assign n27505 = ~controllable_BtoR_REQ0 & ~n27504;
  assign n27506 = ~n15824 & ~n27505;
  assign n27507 = ~i_RtoB_ACK0 & ~n27506;
  assign n27508 = ~n24585 & ~n27507;
  assign n27509 = ~controllable_DEQ & ~n27508;
  assign n27510 = ~n26498 & ~n27509;
  assign n27511 = i_nEMPTY & ~n27510;
  assign n27512 = ~n10415 & ~n20337;
  assign n27513 = ~controllable_BtoR_REQ0 & ~n27512;
  assign n27514 = ~n15843 & ~n27513;
  assign n27515 = ~i_RtoB_ACK0 & ~n27514;
  assign n27516 = ~n24579 & ~n27515;
  assign n27517 = ~controllable_DEQ & ~n27516;
  assign n27518 = ~n22617 & ~n27517;
  assign n27519 = i_FULL & ~n27518;
  assign n27520 = ~n10359 & ~n20347;
  assign n27521 = ~controllable_BtoR_REQ0 & ~n27520;
  assign n27522 = ~n15807 & ~n27521;
  assign n27523 = ~i_RtoB_ACK0 & ~n27522;
  assign n27524 = ~n24579 & ~n27523;
  assign n27525 = ~controllable_DEQ & ~n27524;
  assign n27526 = ~n22627 & ~n27525;
  assign n27527 = ~i_FULL & ~n27526;
  assign n27528 = ~n27519 & ~n27527;
  assign n27529 = ~i_nEMPTY & ~n27528;
  assign n27530 = ~n27511 & ~n27529;
  assign n27531 = ~controllable_BtoS_ACK0 & ~n27530;
  assign n27532 = ~n27503 & ~n27531;
  assign n27533 = n4465 & ~n27532;
  assign n27534 = ~n21013 & ~n27531;
  assign n27535 = ~n4465 & ~n27534;
  assign n27536 = ~n27533 & ~n27535;
  assign n27537 = i_StoB_REQ10 & ~n27536;
  assign n27538 = ~n23169 & ~n27537;
  assign n27539 = controllable_BtoS_ACK10 & ~n27538;
  assign n27540 = ~n12865 & ~n20004;
  assign n27541 = ~controllable_BtoR_REQ0 & ~n27540;
  assign n27542 = ~n20680 & ~n27541;
  assign n27543 = ~i_RtoB_ACK0 & ~n27542;
  assign n27544 = ~n25401 & ~n27543;
  assign n27545 = controllable_DEQ & ~n27544;
  assign n27546 = ~n20685 & ~n26733;
  assign n27547 = ~i_RtoB_ACK0 & ~n27546;
  assign n27548 = ~n25407 & ~n27547;
  assign n27549 = ~controllable_DEQ & ~n27548;
  assign n27550 = ~n27545 & ~n27549;
  assign n27551 = i_FULL & ~n27550;
  assign n27552 = ~n11238 & ~n12891;
  assign n27553 = ~controllable_BtoR_REQ0 & ~n27552;
  assign n27554 = ~n20692 & ~n27553;
  assign n27555 = ~i_RtoB_ACK0 & ~n27554;
  assign n27556 = ~n25401 & ~n27555;
  assign n27557 = controllable_DEQ & ~n27556;
  assign n27558 = ~n12901 & ~n20029;
  assign n27559 = ~controllable_BtoR_REQ0 & ~n27558;
  assign n27560 = ~n20697 & ~n27559;
  assign n27561 = ~i_RtoB_ACK0 & ~n27560;
  assign n27562 = ~n25407 & ~n27561;
  assign n27563 = ~controllable_DEQ & ~n27562;
  assign n27564 = ~n27557 & ~n27563;
  assign n27565 = ~i_FULL & ~n27564;
  assign n27566 = ~n27551 & ~n27565;
  assign n27567 = i_nEMPTY & ~n27566;
  assign n27568 = ~n20711 & ~n26757;
  assign n27569 = ~i_RtoB_ACK0 & ~n27568;
  assign n27570 = ~n25427 & ~n27569;
  assign n27571 = ~controllable_DEQ & ~n27570;
  assign n27572 = ~n23957 & ~n27571;
  assign n27573 = i_FULL & ~n27572;
  assign n27574 = ~controllable_DEQ & ~n27544;
  assign n27575 = ~n23969 & ~n27574;
  assign n27576 = ~i_FULL & ~n27575;
  assign n27577 = ~n27573 & ~n27576;
  assign n27578 = ~i_nEMPTY & ~n27577;
  assign n27579 = ~n27567 & ~n27578;
  assign n27580 = controllable_BtoS_ACK0 & ~n27579;
  assign n27581 = ~n12950 & ~n19931;
  assign n27582 = ~controllable_BtoR_REQ0 & ~n27581;
  assign n27583 = ~n20730 & ~n27582;
  assign n27584 = ~i_RtoB_ACK0 & ~n27583;
  assign n27585 = ~n25442 & ~n27584;
  assign n27586 = controllable_DEQ & ~n27585;
  assign n27587 = ~n20735 & ~n26677;
  assign n27588 = ~i_RtoB_ACK0 & ~n27587;
  assign n27589 = ~n25448 & ~n27588;
  assign n27590 = ~controllable_DEQ & ~n27589;
  assign n27591 = ~n27586 & ~n27590;
  assign n27592 = i_FULL & ~n27591;
  assign n27593 = ~n11317 & ~n12976;
  assign n27594 = ~controllable_BtoR_REQ0 & ~n27593;
  assign n27595 = ~n20742 & ~n27594;
  assign n27596 = ~i_RtoB_ACK0 & ~n27595;
  assign n27597 = ~n25442 & ~n27596;
  assign n27598 = controllable_DEQ & ~n27597;
  assign n27599 = ~n12986 & ~n19953;
  assign n27600 = ~controllable_BtoR_REQ0 & ~n27599;
  assign n27601 = ~n20747 & ~n27600;
  assign n27602 = ~i_RtoB_ACK0 & ~n27601;
  assign n27603 = ~n25448 & ~n27602;
  assign n27604 = ~controllable_DEQ & ~n27603;
  assign n27605 = ~n27598 & ~n27604;
  assign n27606 = ~i_FULL & ~n27605;
  assign n27607 = ~n27592 & ~n27606;
  assign n27608 = i_nEMPTY & ~n27607;
  assign n27609 = ~n20761 & ~n26701;
  assign n27610 = ~i_RtoB_ACK0 & ~n27609;
  assign n27611 = ~n25468 & ~n27610;
  assign n27612 = ~controllable_DEQ & ~n27611;
  assign n27613 = ~n24006 & ~n27612;
  assign n27614 = i_FULL & ~n27613;
  assign n27615 = ~controllable_DEQ & ~n27585;
  assign n27616 = ~n24018 & ~n27615;
  assign n27617 = ~i_FULL & ~n27616;
  assign n27618 = ~n27614 & ~n27617;
  assign n27619 = ~i_nEMPTY & ~n27618;
  assign n27620 = ~n27608 & ~n27619;
  assign n27621 = ~controllable_BtoS_ACK0 & ~n27620;
  assign n27622 = ~n27580 & ~n27621;
  assign n27623 = n4465 & ~n27622;
  assign n27624 = ~n26838 & ~n27621;
  assign n27625 = ~n4465 & ~n27624;
  assign n27626 = ~n27623 & ~n27625;
  assign n27627 = i_StoB_REQ10 & ~n27626;
  assign n27628 = ~n10470 & ~n20004;
  assign n27629 = ~controllable_BtoR_REQ0 & ~n27628;
  assign n27630 = ~n15889 & ~n27629;
  assign n27631 = ~i_RtoB_ACK0 & ~n27630;
  assign n27632 = ~n24611 & ~n27631;
  assign n27633 = controllable_DEQ & ~n27632;
  assign n27634 = ~n15908 & ~n26733;
  assign n27635 = ~i_RtoB_ACK0 & ~n27634;
  assign n27636 = ~n24617 & ~n27635;
  assign n27637 = ~controllable_DEQ & ~n27636;
  assign n27638 = ~n27633 & ~n27637;
  assign n27639 = i_FULL & ~n27638;
  assign n27640 = ~n10508 & ~n11238;
  assign n27641 = ~controllable_BtoR_REQ0 & ~n27640;
  assign n27642 = ~n15927 & ~n27641;
  assign n27643 = ~i_RtoB_ACK0 & ~n27642;
  assign n27644 = ~n24611 & ~n27643;
  assign n27645 = controllable_DEQ & ~n27644;
  assign n27646 = ~n15943 & ~n26747;
  assign n27647 = ~i_RtoB_ACK0 & ~n27646;
  assign n27648 = ~n24617 & ~n27647;
  assign n27649 = ~controllable_DEQ & ~n27648;
  assign n27650 = ~n27645 & ~n27649;
  assign n27651 = ~i_FULL & ~n27650;
  assign n27652 = ~n27639 & ~n27651;
  assign n27653 = i_nEMPTY & ~n27652;
  assign n27654 = ~n15980 & ~n26757;
  assign n27655 = ~i_RtoB_ACK0 & ~n27654;
  assign n27656 = ~n24637 & ~n27655;
  assign n27657 = ~controllable_DEQ & ~n27656;
  assign n27658 = ~n24057 & ~n27657;
  assign n27659 = i_FULL & ~n27658;
  assign n27660 = ~n10470 & ~n20823;
  assign n27661 = ~controllable_BtoR_REQ0 & ~n27660;
  assign n27662 = ~n15889 & ~n27661;
  assign n27663 = ~i_RtoB_ACK0 & ~n27662;
  assign n27664 = ~n24611 & ~n27663;
  assign n27665 = ~controllable_DEQ & ~n27664;
  assign n27666 = ~n24067 & ~n27665;
  assign n27667 = ~i_FULL & ~n27666;
  assign n27668 = ~n27659 & ~n27667;
  assign n27669 = ~i_nEMPTY & ~n27668;
  assign n27670 = ~n27653 & ~n27669;
  assign n27671 = controllable_BtoS_ACK0 & ~n27670;
  assign n27672 = ~n10600 & ~n19931;
  assign n27673 = ~controllable_BtoR_REQ0 & ~n27672;
  assign n27674 = ~n16031 & ~n27673;
  assign n27675 = ~i_RtoB_ACK0 & ~n27674;
  assign n27676 = ~n24655 & ~n27675;
  assign n27677 = controllable_DEQ & ~n27676;
  assign n27678 = ~n16050 & ~n26677;
  assign n27679 = ~i_RtoB_ACK0 & ~n27678;
  assign n27680 = ~n24661 & ~n27679;
  assign n27681 = ~controllable_DEQ & ~n27680;
  assign n27682 = ~n27677 & ~n27681;
  assign n27683 = i_FULL & ~n27682;
  assign n27684 = ~n10635 & ~n11317;
  assign n27685 = ~controllable_BtoR_REQ0 & ~n27684;
  assign n27686 = ~n16069 & ~n27685;
  assign n27687 = ~i_RtoB_ACK0 & ~n27686;
  assign n27688 = ~n24655 & ~n27687;
  assign n27689 = controllable_DEQ & ~n27688;
  assign n27690 = ~n16085 & ~n26790;
  assign n27691 = ~i_RtoB_ACK0 & ~n27690;
  assign n27692 = ~n24661 & ~n27691;
  assign n27693 = ~controllable_DEQ & ~n27692;
  assign n27694 = ~n27689 & ~n27693;
  assign n27695 = ~i_FULL & ~n27694;
  assign n27696 = ~n27683 & ~n27695;
  assign n27697 = i_nEMPTY & ~n27696;
  assign n27698 = ~n16122 & ~n26701;
  assign n27699 = ~i_RtoB_ACK0 & ~n27698;
  assign n27700 = ~n24681 & ~n27699;
  assign n27701 = ~controllable_DEQ & ~n27700;
  assign n27702 = ~n24101 & ~n27701;
  assign n27703 = i_FULL & ~n27702;
  assign n27704 = ~n10600 & ~n19983;
  assign n27705 = ~controllable_BtoR_REQ0 & ~n27704;
  assign n27706 = ~n16031 & ~n27705;
  assign n27707 = ~i_RtoB_ACK0 & ~n27706;
  assign n27708 = ~n24655 & ~n27707;
  assign n27709 = ~controllable_DEQ & ~n27708;
  assign n27710 = ~n24111 & ~n27709;
  assign n27711 = ~i_FULL & ~n27710;
  assign n27712 = ~n27703 & ~n27711;
  assign n27713 = ~i_nEMPTY & ~n27712;
  assign n27714 = ~n27697 & ~n27713;
  assign n27715 = ~controllable_BtoS_ACK0 & ~n27714;
  assign n27716 = ~n27671 & ~n27715;
  assign n27717 = n4465 & ~n27716;
  assign n27718 = ~n26721 & ~n27717;
  assign n27719 = ~i_StoB_REQ10 & ~n27718;
  assign n27720 = ~n27627 & ~n27719;
  assign n27721 = ~controllable_BtoS_ACK10 & ~n27720;
  assign n27722 = ~n27539 & ~n27721;
  assign n27723 = ~n4464 & ~n27722;
  assign n27724 = ~n27475 & ~n27723;
  assign n27725 = n4463 & ~n27724;
  assign n27726 = ~n12172 & ~n20219;
  assign n27727 = ~controllable_BtoR_REQ0 & ~n27726;
  assign n27728 = ~n17545 & ~n27727;
  assign n27729 = ~i_RtoB_ACK0 & ~n27728;
  assign n27730 = ~n25125 & ~n27729;
  assign n27731 = controllable_DEQ & ~n27730;
  assign n27732 = ~n12193 & ~n20229;
  assign n27733 = ~controllable_BtoR_REQ0 & ~n27732;
  assign n27734 = ~n17562 & ~n27733;
  assign n27735 = ~i_RtoB_ACK0 & ~n27734;
  assign n27736 = ~n25131 & ~n27735;
  assign n27737 = ~controllable_DEQ & ~n27736;
  assign n27738 = ~n27731 & ~n27737;
  assign n27739 = i_nEMPTY & ~n27738;
  assign n27740 = ~n12216 & ~n20245;
  assign n27741 = ~controllable_BtoR_REQ0 & ~n27740;
  assign n27742 = ~n17581 & ~n27741;
  assign n27743 = ~i_RtoB_ACK0 & ~n27742;
  assign n27744 = ~n25125 & ~n27743;
  assign n27745 = ~controllable_DEQ & ~n27744;
  assign n27746 = ~n23541 & ~n27745;
  assign n27747 = i_FULL & ~n27746;
  assign n27748 = ~n12172 & ~n20260;
  assign n27749 = ~controllable_BtoR_REQ0 & ~n27748;
  assign n27750 = ~n17545 & ~n27749;
  assign n27751 = ~i_RtoB_ACK0 & ~n27750;
  assign n27752 = ~n25125 & ~n27751;
  assign n27753 = ~controllable_DEQ & ~n27752;
  assign n27754 = ~n23551 & ~n27753;
  assign n27755 = ~i_FULL & ~n27754;
  assign n27756 = ~n27747 & ~n27755;
  assign n27757 = ~i_nEMPTY & ~n27756;
  assign n27758 = ~n27739 & ~n27757;
  assign n27759 = controllable_BtoS_ACK0 & ~n27758;
  assign n27760 = ~n8972 & ~n20274;
  assign n27761 = ~controllable_BtoR_REQ0 & ~n27760;
  assign n27762 = ~n14824 & ~n27761;
  assign n27763 = ~i_RtoB_ACK0 & ~n27762;
  assign n27764 = ~n24189 & ~n27763;
  assign n27765 = controllable_DEQ & ~n27764;
  assign n27766 = ~n8991 & ~n20282;
  assign n27767 = ~controllable_BtoR_REQ0 & ~n27766;
  assign n27768 = ~n14841 & ~n27767;
  assign n27769 = ~i_RtoB_ACK0 & ~n27768;
  assign n27770 = ~n24195 & ~n27769;
  assign n27771 = ~controllable_DEQ & ~n27770;
  assign n27772 = ~n27765 & ~n27771;
  assign n27773 = i_nEMPTY & ~n27772;
  assign n27774 = ~n9028 & ~n20298;
  assign n27775 = ~controllable_BtoR_REQ0 & ~n27774;
  assign n27776 = ~n14860 & ~n27775;
  assign n27777 = ~i_RtoB_ACK0 & ~n27776;
  assign n27778 = ~n24189 & ~n27777;
  assign n27779 = ~controllable_DEQ & ~n27778;
  assign n27780 = ~n23579 & ~n27779;
  assign n27781 = i_FULL & ~n27780;
  assign n27782 = ~n8972 & ~n20313;
  assign n27783 = ~controllable_BtoR_REQ0 & ~n27782;
  assign n27784 = ~n14824 & ~n27783;
  assign n27785 = ~i_RtoB_ACK0 & ~n27784;
  assign n27786 = ~n24189 & ~n27785;
  assign n27787 = ~controllable_DEQ & ~n27786;
  assign n27788 = ~n23589 & ~n27787;
  assign n27789 = ~i_FULL & ~n27788;
  assign n27790 = ~n27781 & ~n27789;
  assign n27791 = ~i_nEMPTY & ~n27790;
  assign n27792 = ~n27773 & ~n27791;
  assign n27793 = ~controllable_BtoS_ACK0 & ~n27792;
  assign n27794 = ~n27759 & ~n27793;
  assign n27795 = n4465 & ~n27794;
  assign n27796 = ~n27247 & ~n27795;
  assign n27797 = i_StoB_REQ10 & ~n27796;
  assign n27798 = ~n23169 & ~n27797;
  assign n27799 = controllable_BtoS_ACK10 & ~n27798;
  assign n27800 = ~n27473 & ~n27799;
  assign n27801 = n4464 & ~n27800;
  assign n27802 = ~n27723 & ~n27801;
  assign n27803 = ~n4463 & ~n27802;
  assign n27804 = ~n27725 & ~n27803;
  assign n27805 = ~n4462 & ~n27804;
  assign n27806 = ~n27147 & ~n27805;
  assign n27807 = ~n4461 & ~n27806;
  assign n27808 = ~n25921 & ~n27807;
  assign n27809 = n4459 & ~n27808;
  assign n27810 = ~n25633 & ~n27809;
  assign n27811 = ~n4455 & ~n27810;
  assign n27812 = ~n20897 & ~n27811;
  assign n27813 = n4445 & ~n27812;
  assign n27814 = controllable_BtoR_REQ1 & ~n18916;
  assign n27815 = ~n18867 & ~n27814;
  assign n27816 = ~controllable_BtoR_REQ0 & ~n27815;
  assign n27817 = ~controllable_BtoR_REQ0 & ~n27816;
  assign n27818 = ~i_RtoB_ACK0 & ~n27817;
  assign n27819 = ~n5236 & ~n27818;
  assign n27820 = controllable_DEQ & ~n27819;
  assign n27821 = ~controllable_BtoR_REQ0 & ~n25928;
  assign n27822 = ~i_RtoB_ACK0 & ~n27821;
  assign n27823 = ~n5259 & ~n27822;
  assign n27824 = ~controllable_DEQ & ~n27823;
  assign n27825 = ~n27820 & ~n27824;
  assign n27826 = i_FULL & ~n27825;
  assign n27827 = ~controllable_BtoR_REQ0 & ~n18887;
  assign n27828 = ~controllable_BtoR_REQ0 & ~n27827;
  assign n27829 = ~i_RtoB_ACK0 & ~n27828;
  assign n27830 = ~n5259 & ~n27829;
  assign n27831 = ~controllable_DEQ & ~n27830;
  assign n27832 = ~n5251 & ~n27831;
  assign n27833 = ~i_FULL & ~n27832;
  assign n27834 = ~n27826 & ~n27833;
  assign n27835 = i_nEMPTY & ~n27834;
  assign n27836 = ~controllable_BtoR_REQ0 & ~n25951;
  assign n27837 = ~i_RtoB_ACK0 & ~n27836;
  assign n27838 = ~n5236 & ~n27837;
  assign n27839 = ~controllable_DEQ & ~n27838;
  assign n27840 = ~n5281 & ~n27839;
  assign n27841 = i_FULL & ~n27840;
  assign n27842 = ~controllable_BtoR_REQ0 & ~n18916;
  assign n27843 = ~controllable_BtoR_REQ0 & ~n27842;
  assign n27844 = ~i_RtoB_ACK0 & ~n27843;
  assign n27845 = ~n5236 & ~n27844;
  assign n27846 = ~controllable_DEQ & ~n27845;
  assign n27847 = ~n5296 & ~n27846;
  assign n27848 = ~i_FULL & ~n27847;
  assign n27849 = ~n27841 & ~n27848;
  assign n27850 = ~i_nEMPTY & ~n27849;
  assign n27851 = ~n27835 & ~n27850;
  assign n27852 = controllable_BtoS_ACK0 & ~n27851;
  assign n27853 = ~i_RtoB_ACK1 & ~n11298;
  assign n27854 = ~i_RtoB_ACK1 & ~n27853;
  assign n27855 = controllable_BtoR_REQ1 & ~n27854;
  assign n27856 = ~n20337 & ~n27855;
  assign n27857 = ~controllable_BtoR_REQ0 & ~n27856;
  assign n27858 = ~controllable_BtoR_REQ0 & ~n27857;
  assign n27859 = i_RtoB_ACK0 & ~n27858;
  assign n27860 = controllable_BtoR_REQ1 & ~n18986;
  assign n27861 = ~n18931 & ~n27860;
  assign n27862 = ~controllable_BtoR_REQ0 & ~n27861;
  assign n27863 = ~controllable_BtoR_REQ0 & ~n27862;
  assign n27864 = ~i_RtoB_ACK0 & ~n27863;
  assign n27865 = ~n27859 & ~n27864;
  assign n27866 = controllable_DEQ & ~n27865;
  assign n27867 = controllable_BtoR_REQ1 & ~n17759;
  assign n27868 = ~n20328 & ~n27867;
  assign n27869 = ~controllable_BtoR_REQ0 & ~n27868;
  assign n27870 = ~controllable_BtoR_REQ0 & ~n27869;
  assign n27871 = i_RtoB_ACK0 & ~n27870;
  assign n27872 = ~controllable_BtoR_REQ0 & ~n25976;
  assign n27873 = ~i_RtoB_ACK0 & ~n27872;
  assign n27874 = ~n27871 & ~n27873;
  assign n27875 = ~controllable_DEQ & ~n27874;
  assign n27876 = ~n27866 & ~n27875;
  assign n27877 = i_FULL & ~n27876;
  assign n27878 = controllable_BtoR_REQ1 & ~n20346;
  assign n27879 = ~n18948 & ~n27878;
  assign n27880 = ~controllable_BtoR_REQ0 & ~n27879;
  assign n27881 = ~controllable_BtoR_REQ0 & ~n27880;
  assign n27882 = ~i_RtoB_ACK0 & ~n27881;
  assign n27883 = ~n27859 & ~n27882;
  assign n27884 = controllable_DEQ & ~n27883;
  assign n27885 = ~controllable_BtoR_REQ0 & ~n18955;
  assign n27886 = ~controllable_BtoR_REQ0 & ~n27885;
  assign n27887 = ~i_RtoB_ACK0 & ~n27886;
  assign n27888 = ~n27871 & ~n27887;
  assign n27889 = ~controllable_DEQ & ~n27888;
  assign n27890 = ~n27884 & ~n27889;
  assign n27891 = ~i_FULL & ~n27890;
  assign n27892 = ~n27877 & ~n27891;
  assign n27893 = i_nEMPTY & ~n27892;
  assign n27894 = controllable_BtoR_REQ1 & ~n17726;
  assign n27895 = ~n8917 & ~n27894;
  assign n27896 = ~controllable_BtoR_REQ0 & ~n27895;
  assign n27897 = ~controllable_BtoR_REQ0 & ~n27896;
  assign n27898 = ~i_RtoB_ACK0 & ~n27897;
  assign n27899 = ~i_RtoB_ACK0 & ~n27898;
  assign n27900 = controllable_DEQ & ~n27899;
  assign n27901 = ~controllable_BtoR_REQ0 & ~n25999;
  assign n27902 = ~i_RtoB_ACK0 & ~n27901;
  assign n27903 = ~n27859 & ~n27902;
  assign n27904 = ~controllable_DEQ & ~n27903;
  assign n27905 = ~n27900 & ~n27904;
  assign n27906 = i_FULL & ~n27905;
  assign n27907 = ~n8936 & ~n27867;
  assign n27908 = ~controllable_BtoR_REQ0 & ~n27907;
  assign n27909 = ~controllable_BtoR_REQ0 & ~n27908;
  assign n27910 = ~i_RtoB_ACK0 & ~n27909;
  assign n27911 = ~i_RtoB_ACK0 & ~n27910;
  assign n27912 = controllable_DEQ & ~n27911;
  assign n27913 = ~controllable_BtoR_REQ0 & ~n18986;
  assign n27914 = ~controllable_BtoR_REQ0 & ~n27913;
  assign n27915 = ~i_RtoB_ACK0 & ~n27914;
  assign n27916 = ~n27859 & ~n27915;
  assign n27917 = ~controllable_DEQ & ~n27916;
  assign n27918 = ~n27912 & ~n27917;
  assign n27919 = ~i_FULL & ~n27918;
  assign n27920 = ~n27906 & ~n27919;
  assign n27921 = ~i_nEMPTY & ~n27920;
  assign n27922 = ~n27893 & ~n27921;
  assign n27923 = ~controllable_BtoS_ACK0 & ~n27922;
  assign n27924 = ~n27852 & ~n27923;
  assign n27925 = n4465 & ~n27924;
  assign n27926 = controllable_BtoR_REQ1 & ~n19052;
  assign n27927 = ~n19003 & ~n27926;
  assign n27928 = ~controllable_BtoR_REQ0 & ~n27927;
  assign n27929 = ~controllable_BtoR_REQ0 & ~n27928;
  assign n27930 = ~i_RtoB_ACK0 & ~n27929;
  assign n27931 = ~n27859 & ~n27930;
  assign n27932 = controllable_DEQ & ~n27931;
  assign n27933 = ~controllable_BtoR_REQ0 & ~n26026;
  assign n27934 = ~i_RtoB_ACK0 & ~n27933;
  assign n27935 = ~n27871 & ~n27934;
  assign n27936 = ~controllable_DEQ & ~n27935;
  assign n27937 = ~n27932 & ~n27936;
  assign n27938 = i_FULL & ~n27937;
  assign n27939 = ~controllable_BtoR_REQ0 & ~n19023;
  assign n27940 = ~controllable_BtoR_REQ0 & ~n27939;
  assign n27941 = ~i_RtoB_ACK0 & ~n27940;
  assign n27942 = ~n27871 & ~n27941;
  assign n27943 = ~controllable_DEQ & ~n27942;
  assign n27944 = ~n27884 & ~n27943;
  assign n27945 = ~i_FULL & ~n27944;
  assign n27946 = ~n27938 & ~n27945;
  assign n27947 = i_nEMPTY & ~n27946;
  assign n27948 = ~controllable_BtoR_REQ0 & ~n26049;
  assign n27949 = ~i_RtoB_ACK0 & ~n27948;
  assign n27950 = ~n27859 & ~n27949;
  assign n27951 = ~controllable_DEQ & ~n27950;
  assign n27952 = ~n27900 & ~n27951;
  assign n27953 = i_FULL & ~n27952;
  assign n27954 = ~controllable_BtoR_REQ0 & ~n19052;
  assign n27955 = ~controllable_BtoR_REQ0 & ~n27954;
  assign n27956 = ~i_RtoB_ACK0 & ~n27955;
  assign n27957 = ~n27859 & ~n27956;
  assign n27958 = ~controllable_DEQ & ~n27957;
  assign n27959 = ~n27912 & ~n27958;
  assign n27960 = ~i_FULL & ~n27959;
  assign n27961 = ~n27953 & ~n27960;
  assign n27962 = ~i_nEMPTY & ~n27961;
  assign n27963 = ~n27947 & ~n27962;
  assign n27964 = ~controllable_BtoS_ACK0 & ~n27963;
  assign n27965 = ~n5307 & ~n27964;
  assign n27966 = ~n4465 & ~n27965;
  assign n27967 = ~n27925 & ~n27966;
  assign n27968 = i_StoB_REQ10 & ~n27967;
  assign n27969 = ~n9599 & ~n9789;
  assign n27970 = controllable_BtoR_REQ1 & ~n27969;
  assign n27971 = ~n19386 & ~n27970;
  assign n27972 = ~controllable_BtoR_REQ0 & ~n27971;
  assign n27973 = ~controllable_BtoR_REQ0 & ~n27972;
  assign n27974 = ~i_RtoB_ACK0 & ~n27973;
  assign n27975 = ~n11234 & ~n27974;
  assign n27976 = controllable_DEQ & ~n27975;
  assign n27977 = ~controllable_BtoR_REQ0 & ~n19394;
  assign n27978 = ~controllable_BtoR_REQ0 & ~n27977;
  assign n27979 = ~i_RtoB_ACK0 & ~n27978;
  assign n27980 = ~n11252 & ~n27979;
  assign n27981 = ~controllable_DEQ & ~n27980;
  assign n27982 = ~n27976 & ~n27981;
  assign n27983 = i_FULL & ~n27982;
  assign n27984 = ~controllable_BtoR_REQ0 & ~n19410;
  assign n27985 = ~controllable_BtoR_REQ0 & ~n27984;
  assign n27986 = ~i_RtoB_ACK0 & ~n27985;
  assign n27987 = ~n11252 & ~n27986;
  assign n27988 = ~controllable_DEQ & ~n27987;
  assign n27989 = ~n11244 & ~n27988;
  assign n27990 = ~i_FULL & ~n27989;
  assign n27991 = ~n27983 & ~n27990;
  assign n27992 = i_nEMPTY & ~n27991;
  assign n27993 = ~controllable_BtoR_REQ0 & ~n19428;
  assign n27994 = ~controllable_BtoR_REQ0 & ~n27993;
  assign n27995 = ~i_RtoB_ACK0 & ~n27994;
  assign n27996 = ~n11234 & ~n27995;
  assign n27997 = ~controllable_DEQ & ~n27996;
  assign n27998 = ~n11269 & ~n27997;
  assign n27999 = i_FULL & ~n27998;
  assign n28000 = ~n9571 & ~n9599;
  assign n28001 = ~controllable_BtoR_REQ1 & ~n28000;
  assign n28002 = ~n27970 & ~n28001;
  assign n28003 = ~controllable_BtoR_REQ0 & ~n28002;
  assign n28004 = ~controllable_BtoR_REQ0 & ~n28003;
  assign n28005 = ~i_RtoB_ACK0 & ~n28004;
  assign n28006 = ~n11234 & ~n28005;
  assign n28007 = ~controllable_DEQ & ~n28006;
  assign n28008 = ~n11282 & ~n28007;
  assign n28009 = ~i_FULL & ~n28008;
  assign n28010 = ~n27999 & ~n28009;
  assign n28011 = ~i_nEMPTY & ~n28010;
  assign n28012 = ~n27992 & ~n28011;
  assign n28013 = controllable_BtoS_ACK0 & ~n28012;
  assign n28014 = ~n9749 & ~n11311;
  assign n28015 = controllable_BtoR_REQ1 & ~n28014;
  assign n28016 = ~n19452 & ~n28015;
  assign n28017 = ~controllable_BtoR_REQ0 & ~n28016;
  assign n28018 = ~controllable_BtoR_REQ0 & ~n28017;
  assign n28019 = ~i_RtoB_ACK0 & ~n28018;
  assign n28020 = ~n11309 & ~n28019;
  assign n28021 = controllable_DEQ & ~n28020;
  assign n28022 = ~controllable_BtoR_REQ0 & ~n19460;
  assign n28023 = ~controllable_BtoR_REQ0 & ~n28022;
  assign n28024 = ~i_RtoB_ACK0 & ~n28023;
  assign n28025 = ~n11332 & ~n28024;
  assign n28026 = ~controllable_DEQ & ~n28025;
  assign n28027 = ~n28021 & ~n28026;
  assign n28028 = i_FULL & ~n28027;
  assign n28029 = ~controllable_BtoR_REQ0 & ~n19476;
  assign n28030 = ~controllable_BtoR_REQ0 & ~n28029;
  assign n28031 = ~i_RtoB_ACK0 & ~n28030;
  assign n28032 = ~n11332 & ~n28031;
  assign n28033 = ~controllable_DEQ & ~n28032;
  assign n28034 = ~n11323 & ~n28033;
  assign n28035 = ~i_FULL & ~n28034;
  assign n28036 = ~n28028 & ~n28035;
  assign n28037 = i_nEMPTY & ~n28036;
  assign n28038 = ~controllable_BtoR_REQ0 & ~n19494;
  assign n28039 = ~controllable_BtoR_REQ0 & ~n28038;
  assign n28040 = ~i_RtoB_ACK0 & ~n28039;
  assign n28041 = ~n11309 & ~n28040;
  assign n28042 = ~controllable_DEQ & ~n28041;
  assign n28043 = ~n11351 & ~n28042;
  assign n28044 = i_FULL & ~n28043;
  assign n28045 = ~n9718 & ~n9749;
  assign n28046 = ~controllable_BtoR_REQ1 & ~n28045;
  assign n28047 = ~n28015 & ~n28046;
  assign n28048 = ~controllable_BtoR_REQ0 & ~n28047;
  assign n28049 = ~controllable_BtoR_REQ0 & ~n28048;
  assign n28050 = ~i_RtoB_ACK0 & ~n28049;
  assign n28051 = ~n11309 & ~n28050;
  assign n28052 = ~controllable_DEQ & ~n28051;
  assign n28053 = ~n11364 & ~n28052;
  assign n28054 = ~i_FULL & ~n28053;
  assign n28055 = ~n28044 & ~n28054;
  assign n28056 = ~i_nEMPTY & ~n28055;
  assign n28057 = ~n28037 & ~n28056;
  assign n28058 = ~controllable_BtoS_ACK0 & ~n28057;
  assign n28059 = ~n28013 & ~n28058;
  assign n28060 = n4465 & ~n28059;
  assign n28061 = ~n9981 & ~n11311;
  assign n28062 = controllable_BtoR_REQ1 & ~n28061;
  assign n28063 = ~n19313 & ~n28062;
  assign n28064 = ~controllable_BtoR_REQ0 & ~n28063;
  assign n28065 = ~controllable_BtoR_REQ0 & ~n28064;
  assign n28066 = ~i_RtoB_ACK0 & ~n28065;
  assign n28067 = ~n11309 & ~n28066;
  assign n28068 = controllable_DEQ & ~n28067;
  assign n28069 = ~controllable_BtoR_REQ0 & ~n19320;
  assign n28070 = ~controllable_BtoR_REQ0 & ~n28069;
  assign n28071 = ~i_RtoB_ACK0 & ~n28070;
  assign n28072 = ~n11332 & ~n28071;
  assign n28073 = ~controllable_DEQ & ~n28072;
  assign n28074 = ~n28068 & ~n28073;
  assign n28075 = i_FULL & ~n28074;
  assign n28076 = ~controllable_BtoR_REQ0 & ~n19334;
  assign n28077 = ~controllable_BtoR_REQ0 & ~n28076;
  assign n28078 = ~i_RtoB_ACK0 & ~n28077;
  assign n28079 = ~n11332 & ~n28078;
  assign n28080 = ~controllable_DEQ & ~n28079;
  assign n28081 = ~n11323 & ~n28080;
  assign n28082 = ~i_FULL & ~n28081;
  assign n28083 = ~n28075 & ~n28082;
  assign n28084 = i_nEMPTY & ~n28083;
  assign n28085 = ~controllable_BtoR_REQ0 & ~n19350;
  assign n28086 = ~controllable_BtoR_REQ0 & ~n28085;
  assign n28087 = ~i_RtoB_ACK0 & ~n28086;
  assign n28088 = ~n11309 & ~n28087;
  assign n28089 = ~controllable_DEQ & ~n28088;
  assign n28090 = ~n11351 & ~n28089;
  assign n28091 = i_FULL & ~n28090;
  assign n28092 = ~n19365 & ~n28062;
  assign n28093 = ~controllable_BtoR_REQ0 & ~n28092;
  assign n28094 = ~controllable_BtoR_REQ0 & ~n28093;
  assign n28095 = ~i_RtoB_ACK0 & ~n28094;
  assign n28096 = ~n11309 & ~n28095;
  assign n28097 = ~controllable_DEQ & ~n28096;
  assign n28098 = ~n11364 & ~n28097;
  assign n28099 = ~i_FULL & ~n28098;
  assign n28100 = ~n28091 & ~n28099;
  assign n28101 = ~i_nEMPTY & ~n28100;
  assign n28102 = ~n28084 & ~n28101;
  assign n28103 = ~controllable_BtoS_ACK0 & ~n28102;
  assign n28104 = ~n11296 & ~n28103;
  assign n28105 = ~n4465 & ~n28104;
  assign n28106 = ~n28060 & ~n28105;
  assign n28107 = ~i_StoB_REQ10 & ~n28106;
  assign n28108 = ~n27968 & ~n28107;
  assign n28109 = controllable_BtoS_ACK10 & ~n28108;
  assign n28110 = controllable_BtoR_REQ1 & ~n17065;
  assign n28111 = ~n11230 & ~n28110;
  assign n28112 = ~controllable_BtoR_REQ0 & ~n28111;
  assign n28113 = ~controllable_BtoR_REQ0 & ~n28112;
  assign n28114 = i_RtoB_ACK0 & ~n28113;
  assign n28115 = ~n9547 & ~n10149;
  assign n28116 = controllable_BtoR_REQ1 & ~n28115;
  assign n28117 = ~n19386 & ~n28116;
  assign n28118 = ~controllable_BtoR_REQ0 & ~n28117;
  assign n28119 = ~controllable_BtoR_REQ0 & ~n28118;
  assign n28120 = ~i_RtoB_ACK0 & ~n28119;
  assign n28121 = ~n28114 & ~n28120;
  assign n28122 = controllable_DEQ & ~n28121;
  assign n28123 = controllable_BtoR_REQ1 & ~n17055;
  assign n28124 = ~n11248 & ~n28123;
  assign n28125 = ~controllable_BtoR_REQ0 & ~n28124;
  assign n28126 = ~controllable_BtoR_REQ0 & ~n28125;
  assign n28127 = i_RtoB_ACK0 & ~n28126;
  assign n28128 = ~n27979 & ~n28127;
  assign n28129 = ~controllable_DEQ & ~n28128;
  assign n28130 = ~n28122 & ~n28129;
  assign n28131 = i_FULL & ~n28130;
  assign n28132 = ~n9813 & ~n10149;
  assign n28133 = controllable_BtoR_REQ1 & ~n28132;
  assign n28134 = ~n11238 & ~n28133;
  assign n28135 = ~controllable_BtoR_REQ0 & ~n28134;
  assign n28136 = ~controllable_BtoR_REQ0 & ~n28135;
  assign n28137 = ~i_RtoB_ACK0 & ~n28136;
  assign n28138 = ~n28114 & ~n28137;
  assign n28139 = controllable_DEQ & ~n28138;
  assign n28140 = ~n27986 & ~n28127;
  assign n28141 = ~controllable_DEQ & ~n28140;
  assign n28142 = ~n28139 & ~n28141;
  assign n28143 = ~i_FULL & ~n28142;
  assign n28144 = ~n28131 & ~n28143;
  assign n28145 = i_nEMPTY & ~n28144;
  assign n28146 = ~n7574 & ~n10047;
  assign n28147 = controllable_BtoR_REQ1 & ~n28146;
  assign n28148 = ~n10049 & ~n28147;
  assign n28149 = ~controllable_BtoR_REQ0 & ~n28148;
  assign n28150 = ~controllable_BtoR_REQ0 & ~n28149;
  assign n28151 = ~i_RtoB_ACK0 & ~n28150;
  assign n28152 = ~i_RtoB_ACK0 & ~n28151;
  assign n28153 = controllable_DEQ & ~n28152;
  assign n28154 = ~n27995 & ~n28114;
  assign n28155 = ~controllable_DEQ & ~n28154;
  assign n28156 = ~n28153 & ~n28155;
  assign n28157 = i_FULL & ~n28156;
  assign n28158 = ~n10061 & ~n28123;
  assign n28159 = ~controllable_BtoR_REQ0 & ~n28158;
  assign n28160 = ~controllable_BtoR_REQ0 & ~n28159;
  assign n28161 = ~i_RtoB_ACK0 & ~n28160;
  assign n28162 = ~i_RtoB_ACK0 & ~n28161;
  assign n28163 = controllable_DEQ & ~n28162;
  assign n28164 = ~controllable_DEQ & ~n28121;
  assign n28165 = ~n28163 & ~n28164;
  assign n28166 = ~i_FULL & ~n28165;
  assign n28167 = ~n28157 & ~n28166;
  assign n28168 = ~i_nEMPTY & ~n28167;
  assign n28169 = ~n28145 & ~n28168;
  assign n28170 = controllable_BtoS_ACK0 & ~n28169;
  assign n28171 = controllable_BtoR_REQ1 & ~n18545;
  assign n28172 = ~n11305 & ~n28171;
  assign n28173 = ~controllable_BtoR_REQ0 & ~n28172;
  assign n28174 = ~controllable_BtoR_REQ0 & ~n28173;
  assign n28175 = i_RtoB_ACK0 & ~n28174;
  assign n28176 = ~n9694 & ~n12462;
  assign n28177 = controllable_BtoR_REQ1 & ~n28176;
  assign n28178 = ~n19452 & ~n28177;
  assign n28179 = ~controllable_BtoR_REQ0 & ~n28178;
  assign n28180 = ~controllable_BtoR_REQ0 & ~n28179;
  assign n28181 = ~i_RtoB_ACK0 & ~n28180;
  assign n28182 = ~n28175 & ~n28181;
  assign n28183 = controllable_DEQ & ~n28182;
  assign n28184 = controllable_BtoR_REQ1 & ~n18527;
  assign n28185 = ~n11328 & ~n28184;
  assign n28186 = ~controllable_BtoR_REQ0 & ~n28185;
  assign n28187 = ~controllable_BtoR_REQ0 & ~n28186;
  assign n28188 = i_RtoB_ACK0 & ~n28187;
  assign n28189 = ~n28024 & ~n28188;
  assign n28190 = ~controllable_DEQ & ~n28189;
  assign n28191 = ~n28183 & ~n28190;
  assign n28192 = i_FULL & ~n28191;
  assign n28193 = ~n9904 & ~n12462;
  assign n28194 = controllable_BtoR_REQ1 & ~n28193;
  assign n28195 = ~n11317 & ~n28194;
  assign n28196 = ~controllable_BtoR_REQ0 & ~n28195;
  assign n28197 = ~controllable_BtoR_REQ0 & ~n28196;
  assign n28198 = ~i_RtoB_ACK0 & ~n28197;
  assign n28199 = ~n28175 & ~n28198;
  assign n28200 = controllable_DEQ & ~n28199;
  assign n28201 = ~n28031 & ~n28188;
  assign n28202 = ~controllable_DEQ & ~n28201;
  assign n28203 = ~n28200 & ~n28202;
  assign n28204 = ~i_FULL & ~n28203;
  assign n28205 = ~n28192 & ~n28204;
  assign n28206 = i_nEMPTY & ~n28205;
  assign n28207 = ~n9949 & ~n11580;
  assign n28208 = controllable_BtoR_REQ1 & ~n28207;
  assign n28209 = ~n9951 & ~n28208;
  assign n28210 = ~controllable_BtoR_REQ0 & ~n28209;
  assign n28211 = ~controllable_BtoR_REQ0 & ~n28210;
  assign n28212 = ~i_RtoB_ACK0 & ~n28211;
  assign n28213 = ~i_RtoB_ACK0 & ~n28212;
  assign n28214 = controllable_DEQ & ~n28213;
  assign n28215 = ~n28040 & ~n28175;
  assign n28216 = ~controllable_DEQ & ~n28215;
  assign n28217 = ~n28214 & ~n28216;
  assign n28218 = i_FULL & ~n28217;
  assign n28219 = ~n9973 & ~n28184;
  assign n28220 = ~controllable_BtoR_REQ0 & ~n28219;
  assign n28221 = ~controllable_BtoR_REQ0 & ~n28220;
  assign n28222 = ~i_RtoB_ACK0 & ~n28221;
  assign n28223 = ~i_RtoB_ACK0 & ~n28222;
  assign n28224 = controllable_DEQ & ~n28223;
  assign n28225 = ~controllable_DEQ & ~n28182;
  assign n28226 = ~n28224 & ~n28225;
  assign n28227 = ~i_FULL & ~n28226;
  assign n28228 = ~n28218 & ~n28227;
  assign n28229 = ~i_nEMPTY & ~n28228;
  assign n28230 = ~n28206 & ~n28229;
  assign n28231 = ~controllable_BtoS_ACK0 & ~n28230;
  assign n28232 = ~n28170 & ~n28231;
  assign n28233 = n4465 & ~n28232;
  assign n28234 = ~n11255 & ~n28127;
  assign n28235 = ~controllable_DEQ & ~n28234;
  assign n28236 = ~n28139 & ~n28235;
  assign n28237 = i_nEMPTY & ~n28236;
  assign n28238 = ~n11272 & ~n28114;
  assign n28239 = ~controllable_DEQ & ~n28238;
  assign n28240 = ~n28153 & ~n28239;
  assign n28241 = i_FULL & ~n28240;
  assign n28242 = ~controllable_DEQ & ~n28138;
  assign n28243 = ~n28163 & ~n28242;
  assign n28244 = ~i_FULL & ~n28243;
  assign n28245 = ~n28241 & ~n28244;
  assign n28246 = ~i_nEMPTY & ~n28245;
  assign n28247 = ~n28237 & ~n28246;
  assign n28248 = controllable_BtoS_ACK0 & ~n28247;
  assign n28249 = ~n9895 & ~n12462;
  assign n28250 = controllable_BtoR_REQ1 & ~n28249;
  assign n28251 = ~n19313 & ~n28250;
  assign n28252 = ~controllable_BtoR_REQ0 & ~n28251;
  assign n28253 = ~controllable_BtoR_REQ0 & ~n28252;
  assign n28254 = ~i_RtoB_ACK0 & ~n28253;
  assign n28255 = ~n28175 & ~n28254;
  assign n28256 = controllable_DEQ & ~n28255;
  assign n28257 = ~n28071 & ~n28188;
  assign n28258 = ~controllable_DEQ & ~n28257;
  assign n28259 = ~n28256 & ~n28258;
  assign n28260 = i_FULL & ~n28259;
  assign n28261 = ~n28078 & ~n28188;
  assign n28262 = ~controllable_DEQ & ~n28261;
  assign n28263 = ~n28200 & ~n28262;
  assign n28264 = ~i_FULL & ~n28263;
  assign n28265 = ~n28260 & ~n28264;
  assign n28266 = i_nEMPTY & ~n28265;
  assign n28267 = ~n28087 & ~n28175;
  assign n28268 = ~controllable_DEQ & ~n28267;
  assign n28269 = ~n28214 & ~n28268;
  assign n28270 = i_FULL & ~n28269;
  assign n28271 = ~controllable_DEQ & ~n28255;
  assign n28272 = ~n28224 & ~n28271;
  assign n28273 = ~i_FULL & ~n28272;
  assign n28274 = ~n28270 & ~n28273;
  assign n28275 = ~i_nEMPTY & ~n28274;
  assign n28276 = ~n28266 & ~n28275;
  assign n28277 = ~controllable_BtoS_ACK0 & ~n28276;
  assign n28278 = ~n28248 & ~n28277;
  assign n28279 = ~n4465 & ~n28278;
  assign n28280 = ~n28233 & ~n28279;
  assign n28281 = i_StoB_REQ10 & ~n28280;
  assign n28282 = ~n28107 & ~n28281;
  assign n28283 = ~controllable_BtoS_ACK10 & ~n28282;
  assign n28284 = ~n28109 & ~n28283;
  assign n28285 = n4464 & ~n28284;
  assign n28286 = controllable_BtoR_REQ1 & ~n19662;
  assign n28287 = ~n19613 & ~n28286;
  assign n28288 = ~controllable_BtoR_REQ0 & ~n28287;
  assign n28289 = ~controllable_BtoR_REQ0 & ~n28288;
  assign n28290 = ~i_RtoB_ACK0 & ~n28289;
  assign n28291 = ~n5236 & ~n28290;
  assign n28292 = controllable_DEQ & ~n28291;
  assign n28293 = ~controllable_BtoR_REQ0 & ~n26438;
  assign n28294 = ~i_RtoB_ACK0 & ~n28293;
  assign n28295 = ~n5259 & ~n28294;
  assign n28296 = ~controllable_DEQ & ~n28295;
  assign n28297 = ~n28292 & ~n28296;
  assign n28298 = i_FULL & ~n28297;
  assign n28299 = ~controllable_BtoR_REQ0 & ~n19633;
  assign n28300 = ~controllable_BtoR_REQ0 & ~n28299;
  assign n28301 = ~i_RtoB_ACK0 & ~n28300;
  assign n28302 = ~n5259 & ~n28301;
  assign n28303 = ~controllable_DEQ & ~n28302;
  assign n28304 = ~n5251 & ~n28303;
  assign n28305 = ~i_FULL & ~n28304;
  assign n28306 = ~n28298 & ~n28305;
  assign n28307 = i_nEMPTY & ~n28306;
  assign n28308 = ~controllable_BtoR_REQ0 & ~n26461;
  assign n28309 = ~i_RtoB_ACK0 & ~n28308;
  assign n28310 = ~n5236 & ~n28309;
  assign n28311 = ~controllable_DEQ & ~n28310;
  assign n28312 = ~n5281 & ~n28311;
  assign n28313 = i_FULL & ~n28312;
  assign n28314 = ~controllable_BtoR_REQ0 & ~n19662;
  assign n28315 = ~controllable_BtoR_REQ0 & ~n28314;
  assign n28316 = ~i_RtoB_ACK0 & ~n28315;
  assign n28317 = ~n5236 & ~n28316;
  assign n28318 = ~controllable_DEQ & ~n28317;
  assign n28319 = ~n5296 & ~n28318;
  assign n28320 = ~i_FULL & ~n28319;
  assign n28321 = ~n28313 & ~n28320;
  assign n28322 = ~i_nEMPTY & ~n28321;
  assign n28323 = ~n28307 & ~n28322;
  assign n28324 = controllable_BtoS_ACK0 & ~n28323;
  assign n28325 = controllable_BtoR_REQ1 & ~n19726;
  assign n28326 = ~n19677 & ~n28325;
  assign n28327 = ~controllable_BtoR_REQ0 & ~n28326;
  assign n28328 = ~controllable_BtoR_REQ0 & ~n28327;
  assign n28329 = ~i_RtoB_ACK0 & ~n28328;
  assign n28330 = ~n27859 & ~n28329;
  assign n28331 = controllable_DEQ & ~n28330;
  assign n28332 = ~controllable_BtoR_REQ0 & ~n26486;
  assign n28333 = ~i_RtoB_ACK0 & ~n28332;
  assign n28334 = ~n27871 & ~n28333;
  assign n28335 = ~controllable_DEQ & ~n28334;
  assign n28336 = ~n28331 & ~n28335;
  assign n28337 = i_FULL & ~n28336;
  assign n28338 = ~controllable_BtoR_REQ0 & ~n19697;
  assign n28339 = ~controllable_BtoR_REQ0 & ~n28338;
  assign n28340 = ~i_RtoB_ACK0 & ~n28339;
  assign n28341 = ~n27871 & ~n28340;
  assign n28342 = ~controllable_DEQ & ~n28341;
  assign n28343 = ~n27884 & ~n28342;
  assign n28344 = ~i_FULL & ~n28343;
  assign n28345 = ~n28337 & ~n28344;
  assign n28346 = i_nEMPTY & ~n28345;
  assign n28347 = ~controllable_BtoR_REQ0 & ~n26509;
  assign n28348 = ~i_RtoB_ACK0 & ~n28347;
  assign n28349 = ~n27859 & ~n28348;
  assign n28350 = ~controllable_DEQ & ~n28349;
  assign n28351 = ~n27900 & ~n28350;
  assign n28352 = i_FULL & ~n28351;
  assign n28353 = ~controllable_BtoR_REQ0 & ~n19726;
  assign n28354 = ~controllable_BtoR_REQ0 & ~n28353;
  assign n28355 = ~i_RtoB_ACK0 & ~n28354;
  assign n28356 = ~n27859 & ~n28355;
  assign n28357 = ~controllable_DEQ & ~n28356;
  assign n28358 = ~n27912 & ~n28357;
  assign n28359 = ~i_FULL & ~n28358;
  assign n28360 = ~n28352 & ~n28359;
  assign n28361 = ~i_nEMPTY & ~n28360;
  assign n28362 = ~n28346 & ~n28361;
  assign n28363 = ~controllable_BtoS_ACK0 & ~n28362;
  assign n28364 = ~n28324 & ~n28363;
  assign n28365 = n4465 & ~n28364;
  assign n28366 = ~n5307 & ~n28363;
  assign n28367 = ~n4465 & ~n28366;
  assign n28368 = ~n28365 & ~n28367;
  assign n28369 = i_StoB_REQ10 & ~n28368;
  assign n28370 = ~n9789 & ~n10568;
  assign n28371 = controllable_BtoR_REQ1 & ~n28370;
  assign n28372 = ~n20004 & ~n28371;
  assign n28373 = ~controllable_BtoR_REQ0 & ~n28372;
  assign n28374 = ~controllable_BtoR_REQ0 & ~n28373;
  assign n28375 = ~i_RtoB_ACK0 & ~n28374;
  assign n28376 = ~n11234 & ~n28375;
  assign n28377 = controllable_DEQ & ~n28376;
  assign n28378 = ~controllable_BtoR_REQ0 & ~n20012;
  assign n28379 = ~controllable_BtoR_REQ0 & ~n28378;
  assign n28380 = ~i_RtoB_ACK0 & ~n28379;
  assign n28381 = ~n11252 & ~n28380;
  assign n28382 = ~controllable_DEQ & ~n28381;
  assign n28383 = ~n28377 & ~n28382;
  assign n28384 = i_FULL & ~n28383;
  assign n28385 = ~controllable_BtoR_REQ0 & ~n20028;
  assign n28386 = ~controllable_BtoR_REQ0 & ~n28385;
  assign n28387 = ~i_RtoB_ACK0 & ~n28386;
  assign n28388 = ~n11252 & ~n28387;
  assign n28389 = ~controllable_DEQ & ~n28388;
  assign n28390 = ~n11244 & ~n28389;
  assign n28391 = ~i_FULL & ~n28390;
  assign n28392 = ~n28384 & ~n28391;
  assign n28393 = i_nEMPTY & ~n28392;
  assign n28394 = ~controllable_BtoR_REQ0 & ~n20046;
  assign n28395 = ~controllable_BtoR_REQ0 & ~n28394;
  assign n28396 = ~i_RtoB_ACK0 & ~n28395;
  assign n28397 = ~n11234 & ~n28396;
  assign n28398 = ~controllable_DEQ & ~n28397;
  assign n28399 = ~n11269 & ~n28398;
  assign n28400 = i_FULL & ~n28399;
  assign n28401 = ~n20823 & ~n28371;
  assign n28402 = ~controllable_BtoR_REQ0 & ~n28401;
  assign n28403 = ~controllable_BtoR_REQ0 & ~n28402;
  assign n28404 = ~i_RtoB_ACK0 & ~n28403;
  assign n28405 = ~n11234 & ~n28404;
  assign n28406 = ~controllable_DEQ & ~n28405;
  assign n28407 = ~n11282 & ~n28406;
  assign n28408 = ~i_FULL & ~n28407;
  assign n28409 = ~n28400 & ~n28408;
  assign n28410 = ~i_nEMPTY & ~n28409;
  assign n28411 = ~n28393 & ~n28410;
  assign n28412 = controllable_BtoS_ACK0 & ~n28411;
  assign n28413 = ~n10695 & ~n11311;
  assign n28414 = controllable_BtoR_REQ1 & ~n28413;
  assign n28415 = ~n19931 & ~n28414;
  assign n28416 = ~controllable_BtoR_REQ0 & ~n28415;
  assign n28417 = ~controllable_BtoR_REQ0 & ~n28416;
  assign n28418 = ~i_RtoB_ACK0 & ~n28417;
  assign n28419 = ~n11309 & ~n28418;
  assign n28420 = controllable_DEQ & ~n28419;
  assign n28421 = ~controllable_BtoR_REQ0 & ~n19938;
  assign n28422 = ~controllable_BtoR_REQ0 & ~n28421;
  assign n28423 = ~i_RtoB_ACK0 & ~n28422;
  assign n28424 = ~n11332 & ~n28423;
  assign n28425 = ~controllable_DEQ & ~n28424;
  assign n28426 = ~n28420 & ~n28425;
  assign n28427 = i_FULL & ~n28426;
  assign n28428 = ~controllable_BtoR_REQ0 & ~n19952;
  assign n28429 = ~controllable_BtoR_REQ0 & ~n28428;
  assign n28430 = ~i_RtoB_ACK0 & ~n28429;
  assign n28431 = ~n11332 & ~n28430;
  assign n28432 = ~controllable_DEQ & ~n28431;
  assign n28433 = ~n11323 & ~n28432;
  assign n28434 = ~i_FULL & ~n28433;
  assign n28435 = ~n28427 & ~n28434;
  assign n28436 = i_nEMPTY & ~n28435;
  assign n28437 = ~controllable_BtoR_REQ0 & ~n19968;
  assign n28438 = ~controllable_BtoR_REQ0 & ~n28437;
  assign n28439 = ~i_RtoB_ACK0 & ~n28438;
  assign n28440 = ~n11309 & ~n28439;
  assign n28441 = ~controllable_DEQ & ~n28440;
  assign n28442 = ~n11351 & ~n28441;
  assign n28443 = i_FULL & ~n28442;
  assign n28444 = ~n19983 & ~n28414;
  assign n28445 = ~controllable_BtoR_REQ0 & ~n28444;
  assign n28446 = ~controllable_BtoR_REQ0 & ~n28445;
  assign n28447 = ~i_RtoB_ACK0 & ~n28446;
  assign n28448 = ~n11309 & ~n28447;
  assign n28449 = ~controllable_DEQ & ~n28448;
  assign n28450 = ~n11364 & ~n28449;
  assign n28451 = ~i_FULL & ~n28450;
  assign n28452 = ~n28443 & ~n28451;
  assign n28453 = ~i_nEMPTY & ~n28452;
  assign n28454 = ~n28436 & ~n28453;
  assign n28455 = ~controllable_BtoS_ACK0 & ~n28454;
  assign n28456 = ~n28412 & ~n28455;
  assign n28457 = n4465 & ~n28456;
  assign n28458 = ~n11296 & ~n28455;
  assign n28459 = ~n4465 & ~n28458;
  assign n28460 = ~n28457 & ~n28459;
  assign n28461 = ~i_StoB_REQ10 & ~n28460;
  assign n28462 = ~n28369 & ~n28461;
  assign n28463 = controllable_BtoS_ACK10 & ~n28462;
  assign n28464 = ~n10149 & ~n10522;
  assign n28465 = controllable_BtoR_REQ1 & ~n28464;
  assign n28466 = ~n20004 & ~n28465;
  assign n28467 = ~controllable_BtoR_REQ0 & ~n28466;
  assign n28468 = ~controllable_BtoR_REQ0 & ~n28467;
  assign n28469 = ~i_RtoB_ACK0 & ~n28468;
  assign n28470 = ~n28114 & ~n28469;
  assign n28471 = controllable_DEQ & ~n28470;
  assign n28472 = ~n28127 & ~n28380;
  assign n28473 = ~controllable_DEQ & ~n28472;
  assign n28474 = ~n28471 & ~n28473;
  assign n28475 = i_FULL & ~n28474;
  assign n28476 = ~n28127 & ~n28387;
  assign n28477 = ~controllable_DEQ & ~n28476;
  assign n28478 = ~n28139 & ~n28477;
  assign n28479 = ~i_FULL & ~n28478;
  assign n28480 = ~n28475 & ~n28479;
  assign n28481 = i_nEMPTY & ~n28480;
  assign n28482 = ~n28114 & ~n28396;
  assign n28483 = ~controllable_DEQ & ~n28482;
  assign n28484 = ~n28153 & ~n28483;
  assign n28485 = i_FULL & ~n28484;
  assign n28486 = ~controllable_DEQ & ~n28470;
  assign n28487 = ~n28163 & ~n28486;
  assign n28488 = ~i_FULL & ~n28487;
  assign n28489 = ~n28485 & ~n28488;
  assign n28490 = ~i_nEMPTY & ~n28489;
  assign n28491 = ~n28481 & ~n28490;
  assign n28492 = controllable_BtoS_ACK0 & ~n28491;
  assign n28493 = ~n10649 & ~n12462;
  assign n28494 = controllable_BtoR_REQ1 & ~n28493;
  assign n28495 = ~n19931 & ~n28494;
  assign n28496 = ~controllable_BtoR_REQ0 & ~n28495;
  assign n28497 = ~controllable_BtoR_REQ0 & ~n28496;
  assign n28498 = ~i_RtoB_ACK0 & ~n28497;
  assign n28499 = ~n28175 & ~n28498;
  assign n28500 = controllable_DEQ & ~n28499;
  assign n28501 = ~n28188 & ~n28423;
  assign n28502 = ~controllable_DEQ & ~n28501;
  assign n28503 = ~n28500 & ~n28502;
  assign n28504 = i_FULL & ~n28503;
  assign n28505 = ~n28188 & ~n28430;
  assign n28506 = ~controllable_DEQ & ~n28505;
  assign n28507 = ~n28200 & ~n28506;
  assign n28508 = ~i_FULL & ~n28507;
  assign n28509 = ~n28504 & ~n28508;
  assign n28510 = i_nEMPTY & ~n28509;
  assign n28511 = ~n28175 & ~n28439;
  assign n28512 = ~controllable_DEQ & ~n28511;
  assign n28513 = ~n28214 & ~n28512;
  assign n28514 = i_FULL & ~n28513;
  assign n28515 = ~controllable_DEQ & ~n28499;
  assign n28516 = ~n28224 & ~n28515;
  assign n28517 = ~i_FULL & ~n28516;
  assign n28518 = ~n28514 & ~n28517;
  assign n28519 = ~i_nEMPTY & ~n28518;
  assign n28520 = ~n28510 & ~n28519;
  assign n28521 = ~controllable_BtoS_ACK0 & ~n28520;
  assign n28522 = ~n28492 & ~n28521;
  assign n28523 = n4465 & ~n28522;
  assign n28524 = ~n28248 & ~n28521;
  assign n28525 = ~n4465 & ~n28524;
  assign n28526 = ~n28523 & ~n28525;
  assign n28527 = i_StoB_REQ10 & ~n28526;
  assign n28528 = ~n28461 & ~n28527;
  assign n28529 = ~controllable_BtoS_ACK10 & ~n28528;
  assign n28530 = ~n28463 & ~n28529;
  assign n28531 = ~n4464 & ~n28530;
  assign n28532 = ~n28285 & ~n28531;
  assign n28533 = n4463 & ~n28532;
  assign n28534 = ~controllable_BtoR_REQ0 & ~n8851;
  assign n28535 = ~controllable_BtoR_REQ0 & ~n28534;
  assign n28536 = ~i_RtoB_ACK0 & ~n28535;
  assign n28537 = ~n27871 & ~n28536;
  assign n28538 = ~controllable_DEQ & ~n28537;
  assign n28539 = ~n27884 & ~n28538;
  assign n28540 = i_nEMPTY & ~n28539;
  assign n28541 = ~controllable_BtoR_REQ0 & ~n8853;
  assign n28542 = ~controllable_BtoR_REQ0 & ~n28541;
  assign n28543 = ~i_RtoB_ACK0 & ~n28542;
  assign n28544 = ~n27859 & ~n28543;
  assign n28545 = ~controllable_DEQ & ~n28544;
  assign n28546 = ~n27900 & ~n28545;
  assign n28547 = i_FULL & ~n28546;
  assign n28548 = ~controllable_BtoR_REQ0 & ~n20346;
  assign n28549 = ~controllable_BtoR_REQ0 & ~n28548;
  assign n28550 = ~i_RtoB_ACK0 & ~n28549;
  assign n28551 = ~n27859 & ~n28550;
  assign n28552 = ~controllable_DEQ & ~n28551;
  assign n28553 = ~n27912 & ~n28552;
  assign n28554 = ~i_FULL & ~n28553;
  assign n28555 = ~n28547 & ~n28554;
  assign n28556 = ~i_nEMPTY & ~n28555;
  assign n28557 = ~n28540 & ~n28556;
  assign n28558 = ~controllable_BtoS_ACK0 & ~n28557;
  assign n28559 = ~n5307 & ~n28558;
  assign n28560 = i_StoB_REQ10 & ~n28559;
  assign n28561 = ~n11380 & ~n28560;
  assign n28562 = controllable_BtoS_ACK10 & ~n28561;
  assign n28563 = ~n11335 & ~n28188;
  assign n28564 = ~controllable_DEQ & ~n28563;
  assign n28565 = ~n28200 & ~n28564;
  assign n28566 = i_nEMPTY & ~n28565;
  assign n28567 = ~n11354 & ~n28175;
  assign n28568 = ~controllable_DEQ & ~n28567;
  assign n28569 = ~n28214 & ~n28568;
  assign n28570 = i_FULL & ~n28569;
  assign n28571 = ~controllable_DEQ & ~n28199;
  assign n28572 = ~n28224 & ~n28571;
  assign n28573 = ~i_FULL & ~n28572;
  assign n28574 = ~n28570 & ~n28573;
  assign n28575 = ~i_nEMPTY & ~n28574;
  assign n28576 = ~n28566 & ~n28575;
  assign n28577 = ~controllable_BtoS_ACK0 & ~n28576;
  assign n28578 = ~n28248 & ~n28577;
  assign n28579 = i_StoB_REQ10 & ~n28578;
  assign n28580 = ~n11380 & ~n28579;
  assign n28581 = ~controllable_BtoS_ACK10 & ~n28580;
  assign n28582 = ~n28562 & ~n28581;
  assign n28583 = ~n4463 & ~n28582;
  assign n28584 = ~n28533 & ~n28583;
  assign n28585 = n4462 & ~n28584;
  assign n28586 = ~n10149 & ~n12370;
  assign n28587 = controllable_BtoR_REQ1 & ~n28586;
  assign n28588 = ~n20368 & ~n28587;
  assign n28589 = ~controllable_BtoR_REQ0 & ~n28588;
  assign n28590 = ~controllable_BtoR_REQ0 & ~n28589;
  assign n28591 = ~i_RtoB_ACK0 & ~n28590;
  assign n28592 = ~n28114 & ~n28591;
  assign n28593 = controllable_DEQ & ~n28592;
  assign n28594 = ~controllable_BtoR_REQ0 & ~n20376;
  assign n28595 = ~controllable_BtoR_REQ0 & ~n28594;
  assign n28596 = ~i_RtoB_ACK0 & ~n28595;
  assign n28597 = ~n28127 & ~n28596;
  assign n28598 = ~controllable_DEQ & ~n28597;
  assign n28599 = ~n28593 & ~n28598;
  assign n28600 = i_FULL & ~n28599;
  assign n28601 = ~controllable_BtoR_REQ0 & ~n20392;
  assign n28602 = ~controllable_BtoR_REQ0 & ~n28601;
  assign n28603 = ~i_RtoB_ACK0 & ~n28602;
  assign n28604 = ~n28127 & ~n28603;
  assign n28605 = ~controllable_DEQ & ~n28604;
  assign n28606 = ~n28139 & ~n28605;
  assign n28607 = ~i_FULL & ~n28606;
  assign n28608 = ~n28600 & ~n28607;
  assign n28609 = i_nEMPTY & ~n28608;
  assign n28610 = ~controllable_BtoR_REQ0 & ~n20410;
  assign n28611 = ~controllable_BtoR_REQ0 & ~n28610;
  assign n28612 = ~i_RtoB_ACK0 & ~n28611;
  assign n28613 = ~n28114 & ~n28612;
  assign n28614 = ~controllable_DEQ & ~n28613;
  assign n28615 = ~n28153 & ~n28614;
  assign n28616 = i_FULL & ~n28615;
  assign n28617 = ~controllable_DEQ & ~n28592;
  assign n28618 = ~n28163 & ~n28617;
  assign n28619 = ~i_FULL & ~n28618;
  assign n28620 = ~n28616 & ~n28619;
  assign n28621 = ~i_nEMPTY & ~n28620;
  assign n28622 = ~n28609 & ~n28621;
  assign n28623 = controllable_BtoS_ACK0 & ~n28622;
  assign n28624 = ~n28277 & ~n28623;
  assign n28625 = n4465 & ~n28624;
  assign n28626 = ~n28279 & ~n28625;
  assign n28627 = i_StoB_REQ10 & ~n28626;
  assign n28628 = ~n9789 & ~n12629;
  assign n28629 = controllable_BtoR_REQ1 & ~n28628;
  assign n28630 = ~n20368 & ~n28629;
  assign n28631 = ~controllable_BtoR_REQ0 & ~n28630;
  assign n28632 = ~controllable_BtoR_REQ0 & ~n28631;
  assign n28633 = ~i_RtoB_ACK0 & ~n28632;
  assign n28634 = ~n11234 & ~n28633;
  assign n28635 = controllable_DEQ & ~n28634;
  assign n28636 = ~n11252 & ~n28596;
  assign n28637 = ~controllable_DEQ & ~n28636;
  assign n28638 = ~n28635 & ~n28637;
  assign n28639 = i_FULL & ~n28638;
  assign n28640 = ~n11252 & ~n28603;
  assign n28641 = ~controllable_DEQ & ~n28640;
  assign n28642 = ~n11244 & ~n28641;
  assign n28643 = ~i_FULL & ~n28642;
  assign n28644 = ~n28639 & ~n28643;
  assign n28645 = i_nEMPTY & ~n28644;
  assign n28646 = ~n11234 & ~n28612;
  assign n28647 = ~controllable_DEQ & ~n28646;
  assign n28648 = ~n11269 & ~n28647;
  assign n28649 = i_FULL & ~n28648;
  assign n28650 = ~n20525 & ~n28629;
  assign n28651 = ~controllable_BtoR_REQ0 & ~n28650;
  assign n28652 = ~controllable_BtoR_REQ0 & ~n28651;
  assign n28653 = ~i_RtoB_ACK0 & ~n28652;
  assign n28654 = ~n11234 & ~n28653;
  assign n28655 = ~controllable_DEQ & ~n28654;
  assign n28656 = ~n11282 & ~n28655;
  assign n28657 = ~i_FULL & ~n28656;
  assign n28658 = ~n28649 & ~n28657;
  assign n28659 = ~i_nEMPTY & ~n28658;
  assign n28660 = ~n28645 & ~n28659;
  assign n28661 = controllable_BtoS_ACK0 & ~n28660;
  assign n28662 = ~n28103 & ~n28661;
  assign n28663 = n4465 & ~n28662;
  assign n28664 = ~n28105 & ~n28663;
  assign n28665 = ~i_StoB_REQ10 & ~n28664;
  assign n28666 = ~n28627 & ~n28665;
  assign n28667 = ~controllable_BtoS_ACK10 & ~n28666;
  assign n28668 = ~n28562 & ~n28667;
  assign n28669 = n4464 & ~n28668;
  assign n28670 = ~n28529 & ~n28562;
  assign n28671 = ~n4464 & ~n28670;
  assign n28672 = ~n28669 & ~n28671;
  assign n28673 = n4463 & ~n28672;
  assign n28674 = ~n28583 & ~n28673;
  assign n28675 = ~n4462 & ~n28674;
  assign n28676 = ~n28585 & ~n28675;
  assign n28677 = ~n4459 & ~n28676;
  assign n28678 = ~n7054 & ~n8835;
  assign n28679 = ~controllable_BtoR_REQ1 & ~n28678;
  assign n28680 = ~controllable_BtoR_REQ1 & ~n28679;
  assign n28681 = controllable_BtoR_REQ0 & ~n28680;
  assign n28682 = ~n18869 & ~n28681;
  assign n28683 = ~i_RtoB_ACK0 & ~n28682;
  assign n28684 = ~n14745 & ~n28683;
  assign n28685 = controllable_DEQ & ~n28684;
  assign n28686 = ~n5038 & ~n7111;
  assign n28687 = ~controllable_BtoR_REQ1 & ~n28686;
  assign n28688 = ~controllable_BtoR_REQ1 & ~n28687;
  assign n28689 = controllable_BtoR_REQ0 & ~n28688;
  assign n28690 = ~n18876 & ~n28689;
  assign n28691 = ~i_RtoB_ACK0 & ~n28690;
  assign n28692 = ~n14761 & ~n28691;
  assign n28693 = ~controllable_DEQ & ~n28692;
  assign n28694 = ~n28685 & ~n28693;
  assign n28695 = i_FULL & ~n28694;
  assign n28696 = ~n7111 & ~n8765;
  assign n28697 = ~controllable_BtoR_REQ1 & ~n28696;
  assign n28698 = ~controllable_BtoR_REQ1 & ~n28697;
  assign n28699 = controllable_BtoR_REQ0 & ~n28698;
  assign n28700 = ~n18890 & ~n28699;
  assign n28701 = ~i_RtoB_ACK0 & ~n28700;
  assign n28702 = ~n14761 & ~n28701;
  assign n28703 = ~controllable_DEQ & ~n28702;
  assign n28704 = ~n14755 & ~n28703;
  assign n28705 = ~i_FULL & ~n28704;
  assign n28706 = ~n28695 & ~n28705;
  assign n28707 = i_nEMPTY & ~n28706;
  assign n28708 = ~n7054 & ~n8817;
  assign n28709 = ~controllable_BtoR_REQ1 & ~n28708;
  assign n28710 = ~controllable_BtoR_REQ1 & ~n28709;
  assign n28711 = controllable_BtoR_REQ0 & ~n28710;
  assign n28712 = ~n18905 & ~n28711;
  assign n28713 = ~i_RtoB_ACK0 & ~n28712;
  assign n28714 = ~n14745 & ~n28713;
  assign n28715 = ~controllable_DEQ & ~n28714;
  assign n28716 = ~n14780 & ~n28715;
  assign n28717 = i_FULL & ~n28716;
  assign n28718 = ~n18919 & ~n28681;
  assign n28719 = ~i_RtoB_ACK0 & ~n28718;
  assign n28720 = ~n14745 & ~n28719;
  assign n28721 = ~controllable_DEQ & ~n28720;
  assign n28722 = ~n14798 & ~n28721;
  assign n28723 = ~i_FULL & ~n28722;
  assign n28724 = ~n28717 & ~n28723;
  assign n28725 = ~i_nEMPTY & ~n28724;
  assign n28726 = ~n28707 & ~n28725;
  assign n28727 = controllable_BtoS_ACK0 & ~n28726;
  assign n28728 = ~n16723 & ~n20339;
  assign n28729 = i_RtoB_ACK0 & ~n28728;
  assign n28730 = ~n8948 & ~n11299;
  assign n28731 = ~controllable_BtoR_REQ1 & ~n28730;
  assign n28732 = ~controllable_BtoR_REQ1 & ~n28731;
  assign n28733 = controllable_BtoR_REQ0 & ~n28732;
  assign n28734 = ~n18933 & ~n28733;
  assign n28735 = ~i_RtoB_ACK0 & ~n28734;
  assign n28736 = ~n28729 & ~n28735;
  assign n28737 = controllable_DEQ & ~n28736;
  assign n28738 = ~n16729 & ~n20330;
  assign n28739 = i_RtoB_ACK0 & ~n28738;
  assign n28740 = ~n5135 & ~n11324;
  assign n28741 = ~controllable_BtoR_REQ1 & ~n28740;
  assign n28742 = ~controllable_BtoR_REQ1 & ~n28741;
  assign n28743 = controllable_BtoR_REQ0 & ~n28742;
  assign n28744 = ~n18940 & ~n28743;
  assign n28745 = ~i_RtoB_ACK0 & ~n28744;
  assign n28746 = ~n28739 & ~n28745;
  assign n28747 = ~controllable_DEQ & ~n28746;
  assign n28748 = ~n28737 & ~n28747;
  assign n28749 = i_FULL & ~n28748;
  assign n28750 = ~n11299 & ~n12317;
  assign n28751 = ~controllable_BtoR_REQ1 & ~n28750;
  assign n28752 = ~controllable_BtoR_REQ1 & ~n28751;
  assign n28753 = controllable_BtoR_REQ0 & ~n28752;
  assign n28754 = ~n18950 & ~n28753;
  assign n28755 = ~i_RtoB_ACK0 & ~n28754;
  assign n28756 = ~n28729 & ~n28755;
  assign n28757 = controllable_DEQ & ~n28756;
  assign n28758 = ~n8866 & ~n11324;
  assign n28759 = ~controllable_BtoR_REQ1 & ~n28758;
  assign n28760 = ~controllable_BtoR_REQ1 & ~n28759;
  assign n28761 = controllable_BtoR_REQ0 & ~n28760;
  assign n28762 = ~n18958 & ~n28761;
  assign n28763 = ~i_RtoB_ACK0 & ~n28762;
  assign n28764 = ~n28739 & ~n28763;
  assign n28765 = ~controllable_DEQ & ~n28764;
  assign n28766 = ~n28757 & ~n28765;
  assign n28767 = ~i_FULL & ~n28766;
  assign n28768 = ~n28749 & ~n28767;
  assign n28769 = i_nEMPTY & ~n28768;
  assign n28770 = ~n17729 & ~n18967;
  assign n28771 = ~i_RtoB_ACK0 & ~n28770;
  assign n28772 = ~i_RtoB_ACK0 & ~n28771;
  assign n28773 = controllable_DEQ & ~n28772;
  assign n28774 = ~n8924 & ~n11299;
  assign n28775 = ~controllable_BtoR_REQ1 & ~n28774;
  assign n28776 = ~controllable_BtoR_REQ1 & ~n28775;
  assign n28777 = controllable_BtoR_REQ0 & ~n28776;
  assign n28778 = ~n18974 & ~n28777;
  assign n28779 = ~i_RtoB_ACK0 & ~n28778;
  assign n28780 = ~n28729 & ~n28779;
  assign n28781 = ~controllable_DEQ & ~n28780;
  assign n28782 = ~n28773 & ~n28781;
  assign n28783 = i_FULL & ~n28782;
  assign n28784 = ~n17762 & ~n18981;
  assign n28785 = ~i_RtoB_ACK0 & ~n28784;
  assign n28786 = ~i_RtoB_ACK0 & ~n28785;
  assign n28787 = controllable_DEQ & ~n28786;
  assign n28788 = ~n18989 & ~n28733;
  assign n28789 = ~i_RtoB_ACK0 & ~n28788;
  assign n28790 = ~n28729 & ~n28789;
  assign n28791 = ~controllable_DEQ & ~n28790;
  assign n28792 = ~n28787 & ~n28791;
  assign n28793 = ~i_FULL & ~n28792;
  assign n28794 = ~n28783 & ~n28793;
  assign n28795 = ~i_nEMPTY & ~n28794;
  assign n28796 = ~n28769 & ~n28795;
  assign n28797 = ~controllable_BtoS_ACK0 & ~n28796;
  assign n28798 = ~n28727 & ~n28797;
  assign n28799 = n4465 & ~n28798;
  assign n28800 = ~n9044 & ~n11299;
  assign n28801 = ~controllable_BtoR_REQ1 & ~n28800;
  assign n28802 = ~controllable_BtoR_REQ1 & ~n28801;
  assign n28803 = controllable_BtoR_REQ0 & ~n28802;
  assign n28804 = ~n19005 & ~n28803;
  assign n28805 = ~i_RtoB_ACK0 & ~n28804;
  assign n28806 = ~n28729 & ~n28805;
  assign n28807 = controllable_DEQ & ~n28806;
  assign n28808 = ~n5349 & ~n11324;
  assign n28809 = ~controllable_BtoR_REQ1 & ~n28808;
  assign n28810 = ~controllable_BtoR_REQ1 & ~n28809;
  assign n28811 = controllable_BtoR_REQ0 & ~n28810;
  assign n28812 = ~n19012 & ~n28811;
  assign n28813 = ~i_RtoB_ACK0 & ~n28812;
  assign n28814 = ~n28739 & ~n28813;
  assign n28815 = ~controllable_DEQ & ~n28814;
  assign n28816 = ~n28807 & ~n28815;
  assign n28817 = i_FULL & ~n28816;
  assign n28818 = ~n8974 & ~n11324;
  assign n28819 = ~controllable_BtoR_REQ1 & ~n28818;
  assign n28820 = ~controllable_BtoR_REQ1 & ~n28819;
  assign n28821 = controllable_BtoR_REQ0 & ~n28820;
  assign n28822 = ~n19026 & ~n28821;
  assign n28823 = ~i_RtoB_ACK0 & ~n28822;
  assign n28824 = ~n28739 & ~n28823;
  assign n28825 = ~controllable_DEQ & ~n28824;
  assign n28826 = ~n28757 & ~n28825;
  assign n28827 = ~i_FULL & ~n28826;
  assign n28828 = ~n28817 & ~n28827;
  assign n28829 = i_nEMPTY & ~n28828;
  assign n28830 = ~n9026 & ~n11299;
  assign n28831 = ~controllable_BtoR_REQ1 & ~n28830;
  assign n28832 = ~controllable_BtoR_REQ1 & ~n28831;
  assign n28833 = controllable_BtoR_REQ0 & ~n28832;
  assign n28834 = ~n19041 & ~n28833;
  assign n28835 = ~i_RtoB_ACK0 & ~n28834;
  assign n28836 = ~n28729 & ~n28835;
  assign n28837 = ~controllable_DEQ & ~n28836;
  assign n28838 = ~n28773 & ~n28837;
  assign n28839 = i_FULL & ~n28838;
  assign n28840 = ~n19055 & ~n28803;
  assign n28841 = ~i_RtoB_ACK0 & ~n28840;
  assign n28842 = ~n28729 & ~n28841;
  assign n28843 = ~controllable_DEQ & ~n28842;
  assign n28844 = ~n28787 & ~n28843;
  assign n28845 = ~i_FULL & ~n28844;
  assign n28846 = ~n28839 & ~n28845;
  assign n28847 = ~i_nEMPTY & ~n28846;
  assign n28848 = ~n28829 & ~n28847;
  assign n28849 = ~controllable_BtoS_ACK0 & ~n28848;
  assign n28850 = ~n14811 & ~n28849;
  assign n28851 = ~n4465 & ~n28850;
  assign n28852 = ~n28799 & ~n28851;
  assign n28853 = i_StoB_REQ10 & ~n28852;
  assign n28854 = ~n9599 & ~n17616;
  assign n28855 = ~controllable_BtoR_REQ1 & ~n28854;
  assign n28856 = ~controllable_BtoR_REQ1 & ~n28855;
  assign n28857 = controllable_BtoR_REQ0 & ~n28856;
  assign n28858 = ~n19388 & ~n28857;
  assign n28859 = ~i_RtoB_ACK0 & ~n28858;
  assign n28860 = ~n17615 & ~n28859;
  assign n28861 = controllable_DEQ & ~n28860;
  assign n28862 = ~n9520 & ~n17631;
  assign n28863 = ~controllable_BtoR_REQ1 & ~n28862;
  assign n28864 = ~controllable_BtoR_REQ1 & ~n28863;
  assign n28865 = controllable_BtoR_REQ0 & ~n28864;
  assign n28866 = ~n19397 & ~n28865;
  assign n28867 = ~i_RtoB_ACK0 & ~n28866;
  assign n28868 = ~n17630 & ~n28867;
  assign n28869 = ~controllable_DEQ & ~n28868;
  assign n28870 = ~n28861 & ~n28869;
  assign n28871 = i_FULL & ~n28870;
  assign n28872 = ~n9547 & ~n17631;
  assign n28873 = ~controllable_BtoR_REQ1 & ~n28872;
  assign n28874 = ~controllable_BtoR_REQ1 & ~n28873;
  assign n28875 = controllable_BtoR_REQ0 & ~n28874;
  assign n28876 = ~n19413 & ~n28875;
  assign n28877 = ~i_RtoB_ACK0 & ~n28876;
  assign n28878 = ~n17630 & ~n28877;
  assign n28879 = ~controllable_DEQ & ~n28878;
  assign n28880 = ~n17626 & ~n28879;
  assign n28881 = ~i_FULL & ~n28880;
  assign n28882 = ~n28871 & ~n28881;
  assign n28883 = i_nEMPTY & ~n28882;
  assign n28884 = ~n9575 & ~n17616;
  assign n28885 = ~controllable_BtoR_REQ1 & ~n28884;
  assign n28886 = ~controllable_BtoR_REQ1 & ~n28885;
  assign n28887 = controllable_BtoR_REQ0 & ~n28886;
  assign n28888 = ~n19431 & ~n28887;
  assign n28889 = ~i_RtoB_ACK0 & ~n28888;
  assign n28890 = ~n17653 & ~n28889;
  assign n28891 = ~controllable_DEQ & ~n28890;
  assign n28892 = ~n17651 & ~n28891;
  assign n28893 = i_FULL & ~n28892;
  assign n28894 = ~controllable_BtoR_REQ1 & ~n28001;
  assign n28895 = ~controllable_BtoR_REQ0 & ~n28894;
  assign n28896 = ~n28857 & ~n28895;
  assign n28897 = ~i_RtoB_ACK0 & ~n28896;
  assign n28898 = ~n17615 & ~n28897;
  assign n28899 = ~controllable_DEQ & ~n28898;
  assign n28900 = ~n17673 & ~n28899;
  assign n28901 = ~i_FULL & ~n28900;
  assign n28902 = ~n28893 & ~n28901;
  assign n28903 = ~i_nEMPTY & ~n28902;
  assign n28904 = ~n28883 & ~n28903;
  assign n28905 = controllable_BtoS_ACK0 & ~n28904;
  assign n28906 = ~n9749 & ~n17695;
  assign n28907 = ~controllable_BtoR_REQ1 & ~n28906;
  assign n28908 = ~controllable_BtoR_REQ1 & ~n28907;
  assign n28909 = controllable_BtoR_REQ0 & ~n28908;
  assign n28910 = ~n19454 & ~n28909;
  assign n28911 = ~i_RtoB_ACK0 & ~n28910;
  assign n28912 = ~n17694 & ~n28911;
  assign n28913 = controllable_DEQ & ~n28912;
  assign n28914 = ~n9667 & ~n17714;
  assign n28915 = ~controllable_BtoR_REQ1 & ~n28914;
  assign n28916 = ~controllable_BtoR_REQ1 & ~n28915;
  assign n28917 = controllable_BtoR_REQ0 & ~n28916;
  assign n28918 = ~n19463 & ~n28917;
  assign n28919 = ~i_RtoB_ACK0 & ~n28918;
  assign n28920 = ~n17713 & ~n28919;
  assign n28921 = ~controllable_DEQ & ~n28920;
  assign n28922 = ~n28913 & ~n28921;
  assign n28923 = i_FULL & ~n28922;
  assign n28924 = ~n9694 & ~n17714;
  assign n28925 = ~controllable_BtoR_REQ1 & ~n28924;
  assign n28926 = ~controllable_BtoR_REQ1 & ~n28925;
  assign n28927 = controllable_BtoR_REQ0 & ~n28926;
  assign n28928 = ~n19479 & ~n28927;
  assign n28929 = ~i_RtoB_ACK0 & ~n28928;
  assign n28930 = ~n17713 & ~n28929;
  assign n28931 = ~controllable_DEQ & ~n28930;
  assign n28932 = ~n17705 & ~n28931;
  assign n28933 = ~i_FULL & ~n28932;
  assign n28934 = ~n28923 & ~n28933;
  assign n28935 = i_nEMPTY & ~n28934;
  assign n28936 = ~n9722 & ~n17695;
  assign n28937 = ~controllable_BtoR_REQ1 & ~n28936;
  assign n28938 = ~controllable_BtoR_REQ1 & ~n28937;
  assign n28939 = controllable_BtoR_REQ0 & ~n28938;
  assign n28940 = ~n19497 & ~n28939;
  assign n28941 = ~i_RtoB_ACK0 & ~n28940;
  assign n28942 = ~n17747 & ~n28941;
  assign n28943 = ~controllable_DEQ & ~n28942;
  assign n28944 = ~n17741 & ~n28943;
  assign n28945 = i_FULL & ~n28944;
  assign n28946 = ~controllable_BtoR_REQ1 & ~n28046;
  assign n28947 = ~controllable_BtoR_REQ0 & ~n28946;
  assign n28948 = ~n28909 & ~n28947;
  assign n28949 = ~i_RtoB_ACK0 & ~n28948;
  assign n28950 = ~n17694 & ~n28949;
  assign n28951 = ~controllable_DEQ & ~n28950;
  assign n28952 = ~n17774 & ~n28951;
  assign n28953 = ~i_FULL & ~n28952;
  assign n28954 = ~n28945 & ~n28953;
  assign n28955 = ~i_nEMPTY & ~n28954;
  assign n28956 = ~n28935 & ~n28955;
  assign n28957 = ~controllable_BtoS_ACK0 & ~n28956;
  assign n28958 = ~n28905 & ~n28957;
  assign n28959 = n4465 & ~n28958;
  assign n28960 = ~n9981 & ~n17695;
  assign n28961 = ~controllable_BtoR_REQ1 & ~n28960;
  assign n28962 = ~controllable_BtoR_REQ1 & ~n28961;
  assign n28963 = controllable_BtoR_REQ0 & ~n28962;
  assign n28964 = ~n19315 & ~n28963;
  assign n28965 = ~i_RtoB_ACK0 & ~n28964;
  assign n28966 = ~n17694 & ~n28965;
  assign n28967 = controllable_DEQ & ~n28966;
  assign n28968 = ~n9913 & ~n17714;
  assign n28969 = ~controllable_BtoR_REQ1 & ~n28968;
  assign n28970 = ~controllable_BtoR_REQ1 & ~n28969;
  assign n28971 = controllable_BtoR_REQ0 & ~n28970;
  assign n28972 = ~n19323 & ~n28971;
  assign n28973 = ~i_RtoB_ACK0 & ~n28972;
  assign n28974 = ~n17713 & ~n28973;
  assign n28975 = ~controllable_DEQ & ~n28974;
  assign n28976 = ~n28967 & ~n28975;
  assign n28977 = i_FULL & ~n28976;
  assign n28978 = ~n9895 & ~n17714;
  assign n28979 = ~controllable_BtoR_REQ1 & ~n28978;
  assign n28980 = ~controllable_BtoR_REQ1 & ~n28979;
  assign n28981 = controllable_BtoR_REQ0 & ~n28980;
  assign n28982 = ~n19337 & ~n28981;
  assign n28983 = ~i_RtoB_ACK0 & ~n28982;
  assign n28984 = ~n17713 & ~n28983;
  assign n28985 = ~controllable_DEQ & ~n28984;
  assign n28986 = ~n17705 & ~n28985;
  assign n28987 = ~i_FULL & ~n28986;
  assign n28988 = ~n28977 & ~n28987;
  assign n28989 = i_nEMPTY & ~n28988;
  assign n28990 = ~n9961 & ~n17695;
  assign n28991 = ~controllable_BtoR_REQ1 & ~n28990;
  assign n28992 = ~controllable_BtoR_REQ1 & ~n28991;
  assign n28993 = controllable_BtoR_REQ0 & ~n28992;
  assign n28994 = ~n19353 & ~n28993;
  assign n28995 = ~i_RtoB_ACK0 & ~n28994;
  assign n28996 = ~n17747 & ~n28995;
  assign n28997 = ~controllable_DEQ & ~n28996;
  assign n28998 = ~n17741 & ~n28997;
  assign n28999 = i_FULL & ~n28998;
  assign n29000 = ~n19367 & ~n28963;
  assign n29001 = ~i_RtoB_ACK0 & ~n29000;
  assign n29002 = ~n17694 & ~n29001;
  assign n29003 = ~controllable_DEQ & ~n29002;
  assign n29004 = ~n17774 & ~n29003;
  assign n29005 = ~i_FULL & ~n29004;
  assign n29006 = ~n28999 & ~n29005;
  assign n29007 = ~i_nEMPTY & ~n29006;
  assign n29008 = ~n28989 & ~n29007;
  assign n29009 = ~controllable_BtoS_ACK0 & ~n29008;
  assign n29010 = ~n17685 & ~n29009;
  assign n29011 = ~n4465 & ~n29010;
  assign n29012 = ~n28959 & ~n29011;
  assign n29013 = ~i_StoB_REQ10 & ~n29012;
  assign n29014 = ~n28853 & ~n29013;
  assign n29015 = controllable_BtoS_ACK10 & ~n29014;
  assign n29016 = ~n17050 & ~n17613;
  assign n29017 = i_RtoB_ACK0 & ~n29016;
  assign n29018 = ~i_RtoB_ACK0 & ~n19387;
  assign n29019 = ~n29017 & ~n29018;
  assign n29020 = controllable_DEQ & ~n29019;
  assign n29021 = ~n17058 & ~n17628;
  assign n29022 = i_RtoB_ACK0 & ~n29021;
  assign n29023 = ~i_RtoB_ACK0 & ~n19396;
  assign n29024 = ~n29022 & ~n29023;
  assign n29025 = ~controllable_DEQ & ~n29024;
  assign n29026 = ~n29020 & ~n29025;
  assign n29027 = i_FULL & ~n29026;
  assign n29028 = ~i_RtoB_ACK0 & ~n17621;
  assign n29029 = ~n29017 & ~n29028;
  assign n29030 = controllable_DEQ & ~n29029;
  assign n29031 = ~i_RtoB_ACK0 & ~n19412;
  assign n29032 = ~n29022 & ~n29031;
  assign n29033 = ~controllable_DEQ & ~n29032;
  assign n29034 = ~n29030 & ~n29033;
  assign n29035 = ~i_FULL & ~n29034;
  assign n29036 = ~n29027 & ~n29035;
  assign n29037 = i_nEMPTY & ~n29036;
  assign n29038 = ~i_RtoB_ACK0 & ~n17646;
  assign n29039 = ~n15604 & ~n29038;
  assign n29040 = controllable_DEQ & ~n29039;
  assign n29041 = ~n17068 & ~n17613;
  assign n29042 = i_RtoB_ACK0 & ~n29041;
  assign n29043 = ~i_RtoB_ACK0 & ~n19430;
  assign n29044 = ~n29042 & ~n29043;
  assign n29045 = ~controllable_DEQ & ~n29044;
  assign n29046 = ~n29040 & ~n29045;
  assign n29047 = i_FULL & ~n29046;
  assign n29048 = ~i_RtoB_ACK0 & ~n17668;
  assign n29049 = ~n15619 & ~n29048;
  assign n29050 = controllable_DEQ & ~n29049;
  assign n29051 = ~controllable_DEQ & ~n29019;
  assign n29052 = ~n29050 & ~n29051;
  assign n29053 = ~i_FULL & ~n29052;
  assign n29054 = ~n29047 & ~n29053;
  assign n29055 = ~i_nEMPTY & ~n29054;
  assign n29056 = ~n29037 & ~n29055;
  assign n29057 = controllable_BtoS_ACK0 & ~n29056;
  assign n29058 = ~n17692 & ~n18522;
  assign n29059 = i_RtoB_ACK0 & ~n29058;
  assign n29060 = ~i_RtoB_ACK0 & ~n19453;
  assign n29061 = ~n29059 & ~n29060;
  assign n29062 = controllable_DEQ & ~n29061;
  assign n29063 = ~n17711 & ~n18530;
  assign n29064 = i_RtoB_ACK0 & ~n29063;
  assign n29065 = ~i_RtoB_ACK0 & ~n19462;
  assign n29066 = ~n29064 & ~n29065;
  assign n29067 = ~controllable_DEQ & ~n29066;
  assign n29068 = ~n29062 & ~n29067;
  assign n29069 = i_FULL & ~n29068;
  assign n29070 = ~i_RtoB_ACK0 & ~n17700;
  assign n29071 = ~n29059 & ~n29070;
  assign n29072 = controllable_DEQ & ~n29071;
  assign n29073 = ~i_RtoB_ACK0 & ~n19478;
  assign n29074 = ~n29064 & ~n29073;
  assign n29075 = ~controllable_DEQ & ~n29074;
  assign n29076 = ~n29072 & ~n29075;
  assign n29077 = ~i_FULL & ~n29076;
  assign n29078 = ~n29069 & ~n29077;
  assign n29079 = i_nEMPTY & ~n29078;
  assign n29080 = ~i_RtoB_ACK0 & ~n17736;
  assign n29081 = ~n17925 & ~n29080;
  assign n29082 = controllable_DEQ & ~n29081;
  assign n29083 = ~n17692 & ~n18548;
  assign n29084 = i_RtoB_ACK0 & ~n29083;
  assign n29085 = ~i_RtoB_ACK0 & ~n19496;
  assign n29086 = ~n29084 & ~n29085;
  assign n29087 = ~controllable_DEQ & ~n29086;
  assign n29088 = ~n29082 & ~n29087;
  assign n29089 = i_FULL & ~n29088;
  assign n29090 = ~i_RtoB_ACK0 & ~n17769;
  assign n29091 = ~n17943 & ~n29090;
  assign n29092 = controllable_DEQ & ~n29091;
  assign n29093 = ~controllable_DEQ & ~n29061;
  assign n29094 = ~n29092 & ~n29093;
  assign n29095 = ~i_FULL & ~n29094;
  assign n29096 = ~n29089 & ~n29095;
  assign n29097 = ~i_nEMPTY & ~n29096;
  assign n29098 = ~n29079 & ~n29097;
  assign n29099 = ~controllable_BtoS_ACK0 & ~n29098;
  assign n29100 = ~n29057 & ~n29099;
  assign n29101 = n4465 & ~n29100;
  assign n29102 = ~i_RtoB_ACK0 & ~n17627;
  assign n29103 = ~n29022 & ~n29102;
  assign n29104 = ~controllable_DEQ & ~n29103;
  assign n29105 = ~n29030 & ~n29104;
  assign n29106 = i_nEMPTY & ~n29105;
  assign n29107 = ~i_RtoB_ACK0 & ~n17612;
  assign n29108 = ~n29042 & ~n29107;
  assign n29109 = ~controllable_DEQ & ~n29108;
  assign n29110 = ~n29040 & ~n29109;
  assign n29111 = i_FULL & ~n29110;
  assign n29112 = ~controllable_DEQ & ~n29029;
  assign n29113 = ~n29050 & ~n29112;
  assign n29114 = ~i_FULL & ~n29113;
  assign n29115 = ~n29111 & ~n29114;
  assign n29116 = ~i_nEMPTY & ~n29115;
  assign n29117 = ~n29106 & ~n29116;
  assign n29118 = controllable_BtoS_ACK0 & ~n29117;
  assign n29119 = ~i_RtoB_ACK0 & ~n19314;
  assign n29120 = ~n29059 & ~n29119;
  assign n29121 = controllable_DEQ & ~n29120;
  assign n29122 = ~i_RtoB_ACK0 & ~n19322;
  assign n29123 = ~n29064 & ~n29122;
  assign n29124 = ~controllable_DEQ & ~n29123;
  assign n29125 = ~n29121 & ~n29124;
  assign n29126 = i_FULL & ~n29125;
  assign n29127 = ~i_RtoB_ACK0 & ~n19336;
  assign n29128 = ~n29064 & ~n29127;
  assign n29129 = ~controllable_DEQ & ~n29128;
  assign n29130 = ~n29072 & ~n29129;
  assign n29131 = ~i_FULL & ~n29130;
  assign n29132 = ~n29126 & ~n29131;
  assign n29133 = i_nEMPTY & ~n29132;
  assign n29134 = ~i_RtoB_ACK0 & ~n19352;
  assign n29135 = ~n29084 & ~n29134;
  assign n29136 = ~controllable_DEQ & ~n29135;
  assign n29137 = ~n29082 & ~n29136;
  assign n29138 = i_FULL & ~n29137;
  assign n29139 = ~controllable_DEQ & ~n29120;
  assign n29140 = ~n29092 & ~n29139;
  assign n29141 = ~i_FULL & ~n29140;
  assign n29142 = ~n29138 & ~n29141;
  assign n29143 = ~i_nEMPTY & ~n29142;
  assign n29144 = ~n29133 & ~n29143;
  assign n29145 = ~controllable_BtoS_ACK0 & ~n29144;
  assign n29146 = ~n29118 & ~n29145;
  assign n29147 = ~n4465 & ~n29146;
  assign n29148 = ~n29101 & ~n29147;
  assign n29149 = i_StoB_REQ10 & ~n29148;
  assign n29150 = ~n29013 & ~n29149;
  assign n29151 = ~controllable_BtoS_ACK10 & ~n29150;
  assign n29152 = ~n29015 & ~n29151;
  assign n29153 = n4464 & ~n29152;
  assign n29154 = ~n7054 & ~n10337;
  assign n29155 = ~controllable_BtoR_REQ1 & ~n29154;
  assign n29156 = ~controllable_BtoR_REQ1 & ~n29155;
  assign n29157 = controllable_BtoR_REQ0 & ~n29156;
  assign n29158 = ~n19615 & ~n29157;
  assign n29159 = ~i_RtoB_ACK0 & ~n29158;
  assign n29160 = ~n14745 & ~n29159;
  assign n29161 = controllable_DEQ & ~n29160;
  assign n29162 = ~n7111 & ~n7716;
  assign n29163 = ~controllable_BtoR_REQ1 & ~n29162;
  assign n29164 = ~controllable_BtoR_REQ1 & ~n29163;
  assign n29165 = controllable_BtoR_REQ0 & ~n29164;
  assign n29166 = ~n19622 & ~n29165;
  assign n29167 = ~i_RtoB_ACK0 & ~n29166;
  assign n29168 = ~n14761 & ~n29167;
  assign n29169 = ~controllable_DEQ & ~n29168;
  assign n29170 = ~n29161 & ~n29169;
  assign n29171 = i_FULL & ~n29170;
  assign n29172 = ~n7111 & ~n10267;
  assign n29173 = ~controllable_BtoR_REQ1 & ~n29172;
  assign n29174 = ~controllable_BtoR_REQ1 & ~n29173;
  assign n29175 = controllable_BtoR_REQ0 & ~n29174;
  assign n29176 = ~n19636 & ~n29175;
  assign n29177 = ~i_RtoB_ACK0 & ~n29176;
  assign n29178 = ~n14761 & ~n29177;
  assign n29179 = ~controllable_DEQ & ~n29178;
  assign n29180 = ~n14755 & ~n29179;
  assign n29181 = ~i_FULL & ~n29180;
  assign n29182 = ~n29171 & ~n29181;
  assign n29183 = i_nEMPTY & ~n29182;
  assign n29184 = ~n7054 & ~n10319;
  assign n29185 = ~controllable_BtoR_REQ1 & ~n29184;
  assign n29186 = ~controllable_BtoR_REQ1 & ~n29185;
  assign n29187 = controllable_BtoR_REQ0 & ~n29186;
  assign n29188 = ~n19651 & ~n29187;
  assign n29189 = ~i_RtoB_ACK0 & ~n29188;
  assign n29190 = ~n14745 & ~n29189;
  assign n29191 = ~controllable_DEQ & ~n29190;
  assign n29192 = ~n14780 & ~n29191;
  assign n29193 = i_FULL & ~n29192;
  assign n29194 = ~n19665 & ~n29157;
  assign n29195 = ~i_RtoB_ACK0 & ~n29194;
  assign n29196 = ~n14745 & ~n29195;
  assign n29197 = ~controllable_DEQ & ~n29196;
  assign n29198 = ~n14798 & ~n29197;
  assign n29199 = ~i_FULL & ~n29198;
  assign n29200 = ~n29193 & ~n29199;
  assign n29201 = ~i_nEMPTY & ~n29200;
  assign n29202 = ~n29183 & ~n29201;
  assign n29203 = controllable_BtoS_ACK0 & ~n29202;
  assign n29204 = ~n10431 & ~n11299;
  assign n29205 = ~controllable_BtoR_REQ1 & ~n29204;
  assign n29206 = ~controllable_BtoR_REQ1 & ~n29205;
  assign n29207 = controllable_BtoR_REQ0 & ~n29206;
  assign n29208 = ~n19679 & ~n29207;
  assign n29209 = ~i_RtoB_ACK0 & ~n29208;
  assign n29210 = ~n28729 & ~n29209;
  assign n29211 = controllable_DEQ & ~n29210;
  assign n29212 = ~n7808 & ~n11324;
  assign n29213 = ~controllable_BtoR_REQ1 & ~n29212;
  assign n29214 = ~controllable_BtoR_REQ1 & ~n29213;
  assign n29215 = controllable_BtoR_REQ0 & ~n29214;
  assign n29216 = ~n19686 & ~n29215;
  assign n29217 = ~i_RtoB_ACK0 & ~n29216;
  assign n29218 = ~n28739 & ~n29217;
  assign n29219 = ~controllable_DEQ & ~n29218;
  assign n29220 = ~n29211 & ~n29219;
  assign n29221 = i_FULL & ~n29220;
  assign n29222 = ~n10361 & ~n11324;
  assign n29223 = ~controllable_BtoR_REQ1 & ~n29222;
  assign n29224 = ~controllable_BtoR_REQ1 & ~n29223;
  assign n29225 = controllable_BtoR_REQ0 & ~n29224;
  assign n29226 = ~n19700 & ~n29225;
  assign n29227 = ~i_RtoB_ACK0 & ~n29226;
  assign n29228 = ~n28739 & ~n29227;
  assign n29229 = ~controllable_DEQ & ~n29228;
  assign n29230 = ~n28757 & ~n29229;
  assign n29231 = ~i_FULL & ~n29230;
  assign n29232 = ~n29221 & ~n29231;
  assign n29233 = i_nEMPTY & ~n29232;
  assign n29234 = ~n10413 & ~n11299;
  assign n29235 = ~controllable_BtoR_REQ1 & ~n29234;
  assign n29236 = ~controllable_BtoR_REQ1 & ~n29235;
  assign n29237 = controllable_BtoR_REQ0 & ~n29236;
  assign n29238 = ~n19715 & ~n29237;
  assign n29239 = ~i_RtoB_ACK0 & ~n29238;
  assign n29240 = ~n28729 & ~n29239;
  assign n29241 = ~controllable_DEQ & ~n29240;
  assign n29242 = ~n28773 & ~n29241;
  assign n29243 = i_FULL & ~n29242;
  assign n29244 = ~n19729 & ~n29207;
  assign n29245 = ~i_RtoB_ACK0 & ~n29244;
  assign n29246 = ~n28729 & ~n29245;
  assign n29247 = ~controllable_DEQ & ~n29246;
  assign n29248 = ~n28787 & ~n29247;
  assign n29249 = ~i_FULL & ~n29248;
  assign n29250 = ~n29243 & ~n29249;
  assign n29251 = ~i_nEMPTY & ~n29250;
  assign n29252 = ~n29233 & ~n29251;
  assign n29253 = ~controllable_BtoS_ACK0 & ~n29252;
  assign n29254 = ~n29203 & ~n29253;
  assign n29255 = n4465 & ~n29254;
  assign n29256 = ~n14811 & ~n29253;
  assign n29257 = ~n4465 & ~n29256;
  assign n29258 = ~n29255 & ~n29257;
  assign n29259 = i_StoB_REQ10 & ~n29258;
  assign n29260 = ~n10568 & ~n17616;
  assign n29261 = ~controllable_BtoR_REQ1 & ~n29260;
  assign n29262 = ~controllable_BtoR_REQ1 & ~n29261;
  assign n29263 = controllable_BtoR_REQ0 & ~n29262;
  assign n29264 = ~n20006 & ~n29263;
  assign n29265 = ~i_RtoB_ACK0 & ~n29264;
  assign n29266 = ~n17615 & ~n29265;
  assign n29267 = controllable_DEQ & ~n29266;
  assign n29268 = ~n10496 & ~n17631;
  assign n29269 = ~controllable_BtoR_REQ1 & ~n29268;
  assign n29270 = ~controllable_BtoR_REQ1 & ~n29269;
  assign n29271 = controllable_BtoR_REQ0 & ~n29270;
  assign n29272 = ~n20015 & ~n29271;
  assign n29273 = ~i_RtoB_ACK0 & ~n29272;
  assign n29274 = ~n17630 & ~n29273;
  assign n29275 = ~controllable_DEQ & ~n29274;
  assign n29276 = ~n29267 & ~n29275;
  assign n29277 = i_FULL & ~n29276;
  assign n29278 = ~n10522 & ~n17631;
  assign n29279 = ~controllable_BtoR_REQ1 & ~n29278;
  assign n29280 = ~controllable_BtoR_REQ1 & ~n29279;
  assign n29281 = controllable_BtoR_REQ0 & ~n29280;
  assign n29282 = ~n20031 & ~n29281;
  assign n29283 = ~i_RtoB_ACK0 & ~n29282;
  assign n29284 = ~n17630 & ~n29283;
  assign n29285 = ~controllable_DEQ & ~n29284;
  assign n29286 = ~n17626 & ~n29285;
  assign n29287 = ~i_FULL & ~n29286;
  assign n29288 = ~n29277 & ~n29287;
  assign n29289 = i_nEMPTY & ~n29288;
  assign n29290 = ~n10548 & ~n17616;
  assign n29291 = ~controllable_BtoR_REQ1 & ~n29290;
  assign n29292 = ~controllable_BtoR_REQ1 & ~n29291;
  assign n29293 = controllable_BtoR_REQ0 & ~n29292;
  assign n29294 = ~n20049 & ~n29293;
  assign n29295 = ~i_RtoB_ACK0 & ~n29294;
  assign n29296 = ~n17653 & ~n29295;
  assign n29297 = ~controllable_DEQ & ~n29296;
  assign n29298 = ~n17651 & ~n29297;
  assign n29299 = i_FULL & ~n29298;
  assign n29300 = ~n20825 & ~n29263;
  assign n29301 = ~i_RtoB_ACK0 & ~n29300;
  assign n29302 = ~n17615 & ~n29301;
  assign n29303 = ~controllable_DEQ & ~n29302;
  assign n29304 = ~n17673 & ~n29303;
  assign n29305 = ~i_FULL & ~n29304;
  assign n29306 = ~n29299 & ~n29305;
  assign n29307 = ~i_nEMPTY & ~n29306;
  assign n29308 = ~n29289 & ~n29307;
  assign n29309 = controllable_BtoS_ACK0 & ~n29308;
  assign n29310 = ~n10695 & ~n17695;
  assign n29311 = ~controllable_BtoR_REQ1 & ~n29310;
  assign n29312 = ~controllable_BtoR_REQ1 & ~n29311;
  assign n29313 = controllable_BtoR_REQ0 & ~n29312;
  assign n29314 = ~n19933 & ~n29313;
  assign n29315 = ~i_RtoB_ACK0 & ~n29314;
  assign n29316 = ~n17694 & ~n29315;
  assign n29317 = controllable_DEQ & ~n29316;
  assign n29318 = ~n10623 & ~n17714;
  assign n29319 = ~controllable_BtoR_REQ1 & ~n29318;
  assign n29320 = ~controllable_BtoR_REQ1 & ~n29319;
  assign n29321 = controllable_BtoR_REQ0 & ~n29320;
  assign n29322 = ~n19941 & ~n29321;
  assign n29323 = ~i_RtoB_ACK0 & ~n29322;
  assign n29324 = ~n17713 & ~n29323;
  assign n29325 = ~controllable_DEQ & ~n29324;
  assign n29326 = ~n29317 & ~n29325;
  assign n29327 = i_FULL & ~n29326;
  assign n29328 = ~n10649 & ~n17714;
  assign n29329 = ~controllable_BtoR_REQ1 & ~n29328;
  assign n29330 = ~controllable_BtoR_REQ1 & ~n29329;
  assign n29331 = controllable_BtoR_REQ0 & ~n29330;
  assign n29332 = ~n19955 & ~n29331;
  assign n29333 = ~i_RtoB_ACK0 & ~n29332;
  assign n29334 = ~n17713 & ~n29333;
  assign n29335 = ~controllable_DEQ & ~n29334;
  assign n29336 = ~n17705 & ~n29335;
  assign n29337 = ~i_FULL & ~n29336;
  assign n29338 = ~n29327 & ~n29337;
  assign n29339 = i_nEMPTY & ~n29338;
  assign n29340 = ~n10675 & ~n17695;
  assign n29341 = ~controllable_BtoR_REQ1 & ~n29340;
  assign n29342 = ~controllable_BtoR_REQ1 & ~n29341;
  assign n29343 = controllable_BtoR_REQ0 & ~n29342;
  assign n29344 = ~n19971 & ~n29343;
  assign n29345 = ~i_RtoB_ACK0 & ~n29344;
  assign n29346 = ~n17747 & ~n29345;
  assign n29347 = ~controllable_DEQ & ~n29346;
  assign n29348 = ~n17741 & ~n29347;
  assign n29349 = i_FULL & ~n29348;
  assign n29350 = ~n19985 & ~n29313;
  assign n29351 = ~i_RtoB_ACK0 & ~n29350;
  assign n29352 = ~n17694 & ~n29351;
  assign n29353 = ~controllable_DEQ & ~n29352;
  assign n29354 = ~n17774 & ~n29353;
  assign n29355 = ~i_FULL & ~n29354;
  assign n29356 = ~n29349 & ~n29355;
  assign n29357 = ~i_nEMPTY & ~n29356;
  assign n29358 = ~n29339 & ~n29357;
  assign n29359 = ~controllable_BtoS_ACK0 & ~n29358;
  assign n29360 = ~n29309 & ~n29359;
  assign n29361 = n4465 & ~n29360;
  assign n29362 = ~n17685 & ~n29359;
  assign n29363 = ~n4465 & ~n29362;
  assign n29364 = ~n29361 & ~n29363;
  assign n29365 = ~i_StoB_REQ10 & ~n29364;
  assign n29366 = ~n29259 & ~n29365;
  assign n29367 = controllable_BtoS_ACK10 & ~n29366;
  assign n29368 = ~i_RtoB_ACK0 & ~n20005;
  assign n29369 = ~n29017 & ~n29368;
  assign n29370 = controllable_DEQ & ~n29369;
  assign n29371 = ~i_RtoB_ACK0 & ~n20014;
  assign n29372 = ~n29022 & ~n29371;
  assign n29373 = ~controllable_DEQ & ~n29372;
  assign n29374 = ~n29370 & ~n29373;
  assign n29375 = i_FULL & ~n29374;
  assign n29376 = ~i_RtoB_ACK0 & ~n20030;
  assign n29377 = ~n29022 & ~n29376;
  assign n29378 = ~controllable_DEQ & ~n29377;
  assign n29379 = ~n29030 & ~n29378;
  assign n29380 = ~i_FULL & ~n29379;
  assign n29381 = ~n29375 & ~n29380;
  assign n29382 = i_nEMPTY & ~n29381;
  assign n29383 = ~i_RtoB_ACK0 & ~n20048;
  assign n29384 = ~n29042 & ~n29383;
  assign n29385 = ~controllable_DEQ & ~n29384;
  assign n29386 = ~n29040 & ~n29385;
  assign n29387 = i_FULL & ~n29386;
  assign n29388 = ~controllable_DEQ & ~n29369;
  assign n29389 = ~n29050 & ~n29388;
  assign n29390 = ~i_FULL & ~n29389;
  assign n29391 = ~n29387 & ~n29390;
  assign n29392 = ~i_nEMPTY & ~n29391;
  assign n29393 = ~n29382 & ~n29392;
  assign n29394 = controllable_BtoS_ACK0 & ~n29393;
  assign n29395 = ~i_RtoB_ACK0 & ~n19932;
  assign n29396 = ~n29059 & ~n29395;
  assign n29397 = controllable_DEQ & ~n29396;
  assign n29398 = ~i_RtoB_ACK0 & ~n19940;
  assign n29399 = ~n29064 & ~n29398;
  assign n29400 = ~controllable_DEQ & ~n29399;
  assign n29401 = ~n29397 & ~n29400;
  assign n29402 = i_FULL & ~n29401;
  assign n29403 = ~i_RtoB_ACK0 & ~n19954;
  assign n29404 = ~n29064 & ~n29403;
  assign n29405 = ~controllable_DEQ & ~n29404;
  assign n29406 = ~n29072 & ~n29405;
  assign n29407 = ~i_FULL & ~n29406;
  assign n29408 = ~n29402 & ~n29407;
  assign n29409 = i_nEMPTY & ~n29408;
  assign n29410 = ~i_RtoB_ACK0 & ~n19970;
  assign n29411 = ~n29084 & ~n29410;
  assign n29412 = ~controllable_DEQ & ~n29411;
  assign n29413 = ~n29082 & ~n29412;
  assign n29414 = i_FULL & ~n29413;
  assign n29415 = ~controllable_DEQ & ~n29396;
  assign n29416 = ~n29092 & ~n29415;
  assign n29417 = ~i_FULL & ~n29416;
  assign n29418 = ~n29414 & ~n29417;
  assign n29419 = ~i_nEMPTY & ~n29418;
  assign n29420 = ~n29409 & ~n29419;
  assign n29421 = ~controllable_BtoS_ACK0 & ~n29420;
  assign n29422 = ~n29394 & ~n29421;
  assign n29423 = n4465 & ~n29422;
  assign n29424 = ~n29118 & ~n29421;
  assign n29425 = ~n4465 & ~n29424;
  assign n29426 = ~n29423 & ~n29425;
  assign n29427 = i_StoB_REQ10 & ~n29426;
  assign n29428 = ~n29365 & ~n29427;
  assign n29429 = ~controllable_BtoS_ACK10 & ~n29428;
  assign n29430 = ~n29367 & ~n29429;
  assign n29431 = ~n4464 & ~n29430;
  assign n29432 = ~n29153 & ~n29431;
  assign n29433 = n4462 & ~n29432;
  assign n29434 = ~n8876 & ~n11324;
  assign n29435 = ~controllable_BtoR_REQ1 & ~n29434;
  assign n29436 = ~controllable_BtoR_REQ1 & ~n29435;
  assign n29437 = controllable_BtoR_REQ0 & ~n29436;
  assign n29438 = ~n20330 & ~n29437;
  assign n29439 = ~i_RtoB_ACK0 & ~n29438;
  assign n29440 = ~n28739 & ~n29439;
  assign n29441 = ~controllable_DEQ & ~n29440;
  assign n29442 = ~n28757 & ~n29441;
  assign n29443 = i_nEMPTY & ~n29442;
  assign n29444 = ~n8854 & ~n11299;
  assign n29445 = ~controllable_BtoR_REQ1 & ~n29444;
  assign n29446 = ~controllable_BtoR_REQ1 & ~n29445;
  assign n29447 = controllable_BtoR_REQ0 & ~n29446;
  assign n29448 = ~n20339 & ~n29447;
  assign n29449 = ~i_RtoB_ACK0 & ~n29448;
  assign n29450 = ~n28729 & ~n29449;
  assign n29451 = ~controllable_DEQ & ~n29450;
  assign n29452 = ~n28773 & ~n29451;
  assign n29453 = i_FULL & ~n29452;
  assign n29454 = ~n20349 & ~n28753;
  assign n29455 = ~i_RtoB_ACK0 & ~n29454;
  assign n29456 = ~n28729 & ~n29455;
  assign n29457 = ~controllable_DEQ & ~n29456;
  assign n29458 = ~n28787 & ~n29457;
  assign n29459 = ~i_FULL & ~n29458;
  assign n29460 = ~n29453 & ~n29459;
  assign n29461 = ~i_nEMPTY & ~n29460;
  assign n29462 = ~n29443 & ~n29461;
  assign n29463 = ~controllable_BtoS_ACK0 & ~n29462;
  assign n29464 = ~n14811 & ~n29463;
  assign n29465 = i_StoB_REQ10 & ~n29464;
  assign n29466 = ~n17788 & ~n29465;
  assign n29467 = controllable_BtoS_ACK10 & ~n29466;
  assign n29468 = ~i_RtoB_ACK0 & ~n20369;
  assign n29469 = ~n29017 & ~n29468;
  assign n29470 = controllable_DEQ & ~n29469;
  assign n29471 = ~i_RtoB_ACK0 & ~n20378;
  assign n29472 = ~n29022 & ~n29471;
  assign n29473 = ~controllable_DEQ & ~n29472;
  assign n29474 = ~n29470 & ~n29473;
  assign n29475 = i_FULL & ~n29474;
  assign n29476 = ~i_RtoB_ACK0 & ~n20394;
  assign n29477 = ~n29022 & ~n29476;
  assign n29478 = ~controllable_DEQ & ~n29477;
  assign n29479 = ~n29030 & ~n29478;
  assign n29480 = ~i_FULL & ~n29479;
  assign n29481 = ~n29475 & ~n29480;
  assign n29482 = i_nEMPTY & ~n29481;
  assign n29483 = ~i_RtoB_ACK0 & ~n20412;
  assign n29484 = ~n29042 & ~n29483;
  assign n29485 = ~controllable_DEQ & ~n29484;
  assign n29486 = ~n29040 & ~n29485;
  assign n29487 = i_FULL & ~n29486;
  assign n29488 = ~controllable_DEQ & ~n29469;
  assign n29489 = ~n29050 & ~n29488;
  assign n29490 = ~i_FULL & ~n29489;
  assign n29491 = ~n29487 & ~n29490;
  assign n29492 = ~i_nEMPTY & ~n29491;
  assign n29493 = ~n29482 & ~n29492;
  assign n29494 = controllable_BtoS_ACK0 & ~n29493;
  assign n29495 = ~n29145 & ~n29494;
  assign n29496 = n4465 & ~n29495;
  assign n29497 = ~n29147 & ~n29496;
  assign n29498 = i_StoB_REQ10 & ~n29497;
  assign n29499 = ~n12629 & ~n17616;
  assign n29500 = ~controllable_BtoR_REQ1 & ~n29499;
  assign n29501 = ~controllable_BtoR_REQ1 & ~n29500;
  assign n29502 = controllable_BtoR_REQ0 & ~n29501;
  assign n29503 = ~n20370 & ~n29502;
  assign n29504 = ~i_RtoB_ACK0 & ~n29503;
  assign n29505 = ~n17615 & ~n29504;
  assign n29506 = controllable_DEQ & ~n29505;
  assign n29507 = ~n12387 & ~n17631;
  assign n29508 = ~controllable_BtoR_REQ1 & ~n29507;
  assign n29509 = ~controllable_BtoR_REQ1 & ~n29508;
  assign n29510 = controllable_BtoR_REQ0 & ~n29509;
  assign n29511 = ~n20379 & ~n29510;
  assign n29512 = ~i_RtoB_ACK0 & ~n29511;
  assign n29513 = ~n17630 & ~n29512;
  assign n29514 = ~controllable_DEQ & ~n29513;
  assign n29515 = ~n29506 & ~n29514;
  assign n29516 = i_FULL & ~n29515;
  assign n29517 = ~n12370 & ~n17631;
  assign n29518 = ~controllable_BtoR_REQ1 & ~n29517;
  assign n29519 = ~controllable_BtoR_REQ1 & ~n29518;
  assign n29520 = controllable_BtoR_REQ0 & ~n29519;
  assign n29521 = ~n20395 & ~n29520;
  assign n29522 = ~i_RtoB_ACK0 & ~n29521;
  assign n29523 = ~n17630 & ~n29522;
  assign n29524 = ~controllable_DEQ & ~n29523;
  assign n29525 = ~n17626 & ~n29524;
  assign n29526 = ~i_FULL & ~n29525;
  assign n29527 = ~n29516 & ~n29526;
  assign n29528 = i_nEMPTY & ~n29527;
  assign n29529 = ~n12431 & ~n17616;
  assign n29530 = ~controllable_BtoR_REQ1 & ~n29529;
  assign n29531 = ~controllable_BtoR_REQ1 & ~n29530;
  assign n29532 = controllable_BtoR_REQ0 & ~n29531;
  assign n29533 = ~n20413 & ~n29532;
  assign n29534 = ~i_RtoB_ACK0 & ~n29533;
  assign n29535 = ~n17653 & ~n29534;
  assign n29536 = ~controllable_DEQ & ~n29535;
  assign n29537 = ~n17651 & ~n29536;
  assign n29538 = i_FULL & ~n29537;
  assign n29539 = ~n20527 & ~n29502;
  assign n29540 = ~i_RtoB_ACK0 & ~n29539;
  assign n29541 = ~n17615 & ~n29540;
  assign n29542 = ~controllable_DEQ & ~n29541;
  assign n29543 = ~n17673 & ~n29542;
  assign n29544 = ~i_FULL & ~n29543;
  assign n29545 = ~n29538 & ~n29544;
  assign n29546 = ~i_nEMPTY & ~n29545;
  assign n29547 = ~n29528 & ~n29546;
  assign n29548 = controllable_BtoS_ACK0 & ~n29547;
  assign n29549 = ~n29009 & ~n29548;
  assign n29550 = n4465 & ~n29549;
  assign n29551 = ~n29011 & ~n29550;
  assign n29552 = ~i_StoB_REQ10 & ~n29551;
  assign n29553 = ~n29498 & ~n29552;
  assign n29554 = ~controllable_BtoS_ACK10 & ~n29553;
  assign n29555 = ~n29467 & ~n29554;
  assign n29556 = n4464 & ~n29555;
  assign n29557 = ~n29429 & ~n29467;
  assign n29558 = ~n4464 & ~n29557;
  assign n29559 = ~n29556 & ~n29558;
  assign n29560 = ~n4462 & ~n29559;
  assign n29561 = ~n29433 & ~n29560;
  assign n29562 = n4461 & ~n29561;
  assign n29563 = ~i_RtoB_ACK0 & ~n17710;
  assign n29564 = ~n29064 & ~n29563;
  assign n29565 = ~controllable_DEQ & ~n29564;
  assign n29566 = ~n29072 & ~n29565;
  assign n29567 = i_nEMPTY & ~n29566;
  assign n29568 = ~i_RtoB_ACK0 & ~n17691;
  assign n29569 = ~n29084 & ~n29568;
  assign n29570 = ~controllable_DEQ & ~n29569;
  assign n29571 = ~n29082 & ~n29570;
  assign n29572 = i_FULL & ~n29571;
  assign n29573 = ~controllable_DEQ & ~n29071;
  assign n29574 = ~n29092 & ~n29573;
  assign n29575 = ~i_FULL & ~n29574;
  assign n29576 = ~n29572 & ~n29575;
  assign n29577 = ~i_nEMPTY & ~n29576;
  assign n29578 = ~n29567 & ~n29577;
  assign n29579 = ~controllable_BtoS_ACK0 & ~n29578;
  assign n29580 = ~n29118 & ~n29579;
  assign n29581 = i_StoB_REQ10 & ~n29580;
  assign n29582 = ~n17788 & ~n29581;
  assign n29583 = ~controllable_BtoS_ACK10 & ~n29582;
  assign n29584 = ~n29467 & ~n29583;
  assign n29585 = ~n4461 & ~n29584;
  assign n29586 = ~n29562 & ~n29585;
  assign n29587 = n4459 & ~n29586;
  assign n29588 = ~n28677 & ~n29587;
  assign n29589 = n4455 & ~n29588;
  assign n29590 = ~n27816 & ~n28681;
  assign n29591 = ~i_RtoB_ACK0 & ~n29590;
  assign n29592 = ~n20977 & ~n29591;
  assign n29593 = controllable_DEQ & ~n29592;
  assign n29594 = ~n25928 & ~n28689;
  assign n29595 = ~i_RtoB_ACK0 & ~n29594;
  assign n29596 = ~n20983 & ~n29595;
  assign n29597 = ~controllable_DEQ & ~n29596;
  assign n29598 = ~n29593 & ~n29597;
  assign n29599 = i_FULL & ~n29598;
  assign n29600 = ~n27827 & ~n28699;
  assign n29601 = ~i_RtoB_ACK0 & ~n29600;
  assign n29602 = ~n20983 & ~n29601;
  assign n29603 = ~controllable_DEQ & ~n29602;
  assign n29604 = ~n20981 & ~n29603;
  assign n29605 = ~i_FULL & ~n29604;
  assign n29606 = ~n29599 & ~n29605;
  assign n29607 = i_nEMPTY & ~n29606;
  assign n29608 = ~n25951 & ~n28711;
  assign n29609 = ~i_RtoB_ACK0 & ~n29608;
  assign n29610 = ~n20977 & ~n29609;
  assign n29611 = ~controllable_DEQ & ~n29610;
  assign n29612 = ~n20993 & ~n29611;
  assign n29613 = i_FULL & ~n29612;
  assign n29614 = ~n27842 & ~n28681;
  assign n29615 = ~i_RtoB_ACK0 & ~n29614;
  assign n29616 = ~n20977 & ~n29615;
  assign n29617 = ~controllable_DEQ & ~n29616;
  assign n29618 = ~n21003 & ~n29617;
  assign n29619 = ~i_FULL & ~n29618;
  assign n29620 = ~n29613 & ~n29619;
  assign n29621 = ~i_nEMPTY & ~n29620;
  assign n29622 = ~n29607 & ~n29621;
  assign n29623 = controllable_BtoS_ACK0 & ~n29622;
  assign n29624 = ~n16723 & ~n27857;
  assign n29625 = i_RtoB_ACK0 & ~n29624;
  assign n29626 = ~n27862 & ~n28733;
  assign n29627 = ~i_RtoB_ACK0 & ~n29626;
  assign n29628 = ~n29625 & ~n29627;
  assign n29629 = controllable_DEQ & ~n29628;
  assign n29630 = ~n16729 & ~n27869;
  assign n29631 = i_RtoB_ACK0 & ~n29630;
  assign n29632 = ~n25976 & ~n28743;
  assign n29633 = ~i_RtoB_ACK0 & ~n29632;
  assign n29634 = ~n29631 & ~n29633;
  assign n29635 = ~controllable_DEQ & ~n29634;
  assign n29636 = ~n29629 & ~n29635;
  assign n29637 = i_FULL & ~n29636;
  assign n29638 = ~n27880 & ~n28753;
  assign n29639 = ~i_RtoB_ACK0 & ~n29638;
  assign n29640 = ~n29625 & ~n29639;
  assign n29641 = controllable_DEQ & ~n29640;
  assign n29642 = ~n27885 & ~n28761;
  assign n29643 = ~i_RtoB_ACK0 & ~n29642;
  assign n29644 = ~n29631 & ~n29643;
  assign n29645 = ~controllable_DEQ & ~n29644;
  assign n29646 = ~n29641 & ~n29645;
  assign n29647 = ~i_FULL & ~n29646;
  assign n29648 = ~n29637 & ~n29647;
  assign n29649 = i_nEMPTY & ~n29648;
  assign n29650 = ~n17729 & ~n27896;
  assign n29651 = ~i_RtoB_ACK0 & ~n29650;
  assign n29652 = ~i_RtoB_ACK0 & ~n29651;
  assign n29653 = controllable_DEQ & ~n29652;
  assign n29654 = ~n25999 & ~n28777;
  assign n29655 = ~i_RtoB_ACK0 & ~n29654;
  assign n29656 = ~n29625 & ~n29655;
  assign n29657 = ~controllable_DEQ & ~n29656;
  assign n29658 = ~n29653 & ~n29657;
  assign n29659 = i_FULL & ~n29658;
  assign n29660 = ~n17762 & ~n27908;
  assign n29661 = ~i_RtoB_ACK0 & ~n29660;
  assign n29662 = ~i_RtoB_ACK0 & ~n29661;
  assign n29663 = controllable_DEQ & ~n29662;
  assign n29664 = ~n27913 & ~n28733;
  assign n29665 = ~i_RtoB_ACK0 & ~n29664;
  assign n29666 = ~n29625 & ~n29665;
  assign n29667 = ~controllable_DEQ & ~n29666;
  assign n29668 = ~n29663 & ~n29667;
  assign n29669 = ~i_FULL & ~n29668;
  assign n29670 = ~n29659 & ~n29669;
  assign n29671 = ~i_nEMPTY & ~n29670;
  assign n29672 = ~n29649 & ~n29671;
  assign n29673 = ~controllable_BtoS_ACK0 & ~n29672;
  assign n29674 = ~n29623 & ~n29673;
  assign n29675 = n4465 & ~n29674;
  assign n29676 = ~n27928 & ~n28803;
  assign n29677 = ~i_RtoB_ACK0 & ~n29676;
  assign n29678 = ~n29625 & ~n29677;
  assign n29679 = controllable_DEQ & ~n29678;
  assign n29680 = ~n26026 & ~n28811;
  assign n29681 = ~i_RtoB_ACK0 & ~n29680;
  assign n29682 = ~n29631 & ~n29681;
  assign n29683 = ~controllable_DEQ & ~n29682;
  assign n29684 = ~n29679 & ~n29683;
  assign n29685 = i_FULL & ~n29684;
  assign n29686 = ~n27939 & ~n28821;
  assign n29687 = ~i_RtoB_ACK0 & ~n29686;
  assign n29688 = ~n29631 & ~n29687;
  assign n29689 = ~controllable_DEQ & ~n29688;
  assign n29690 = ~n29641 & ~n29689;
  assign n29691 = ~i_FULL & ~n29690;
  assign n29692 = ~n29685 & ~n29691;
  assign n29693 = i_nEMPTY & ~n29692;
  assign n29694 = ~n26049 & ~n28833;
  assign n29695 = ~i_RtoB_ACK0 & ~n29694;
  assign n29696 = ~n29625 & ~n29695;
  assign n29697 = ~controllable_DEQ & ~n29696;
  assign n29698 = ~n29653 & ~n29697;
  assign n29699 = i_FULL & ~n29698;
  assign n29700 = ~n27954 & ~n28803;
  assign n29701 = ~i_RtoB_ACK0 & ~n29700;
  assign n29702 = ~n29625 & ~n29701;
  assign n29703 = ~controllable_DEQ & ~n29702;
  assign n29704 = ~n29663 & ~n29703;
  assign n29705 = ~i_FULL & ~n29704;
  assign n29706 = ~n29699 & ~n29705;
  assign n29707 = ~i_nEMPTY & ~n29706;
  assign n29708 = ~n29693 & ~n29707;
  assign n29709 = ~controllable_BtoS_ACK0 & ~n29708;
  assign n29710 = ~n21013 & ~n29709;
  assign n29711 = ~n4465 & ~n29710;
  assign n29712 = ~n29675 & ~n29711;
  assign n29713 = i_StoB_REQ10 & ~n29712;
  assign n29714 = ~n27972 & ~n28857;
  assign n29715 = ~i_RtoB_ACK0 & ~n29714;
  assign n29716 = ~n23089 & ~n29715;
  assign n29717 = controllable_DEQ & ~n29716;
  assign n29718 = ~n27977 & ~n28865;
  assign n29719 = ~i_RtoB_ACK0 & ~n29718;
  assign n29720 = ~n23095 & ~n29719;
  assign n29721 = ~controllable_DEQ & ~n29720;
  assign n29722 = ~n29717 & ~n29721;
  assign n29723 = i_FULL & ~n29722;
  assign n29724 = ~n27984 & ~n28875;
  assign n29725 = ~i_RtoB_ACK0 & ~n29724;
  assign n29726 = ~n23095 & ~n29725;
  assign n29727 = ~controllable_DEQ & ~n29726;
  assign n29728 = ~n23093 & ~n29727;
  assign n29729 = ~i_FULL & ~n29728;
  assign n29730 = ~n29723 & ~n29729;
  assign n29731 = i_nEMPTY & ~n29730;
  assign n29732 = ~n27993 & ~n28887;
  assign n29733 = ~i_RtoB_ACK0 & ~n29732;
  assign n29734 = ~n23107 & ~n29733;
  assign n29735 = ~controllable_DEQ & ~n29734;
  assign n29736 = ~n23105 & ~n29735;
  assign n29737 = i_FULL & ~n29736;
  assign n29738 = ~n28003 & ~n28857;
  assign n29739 = ~i_RtoB_ACK0 & ~n29738;
  assign n29740 = ~n23089 & ~n29739;
  assign n29741 = ~controllable_DEQ & ~n29740;
  assign n29742 = ~n23117 & ~n29741;
  assign n29743 = ~i_FULL & ~n29742;
  assign n29744 = ~n29737 & ~n29743;
  assign n29745 = ~i_nEMPTY & ~n29744;
  assign n29746 = ~n29731 & ~n29745;
  assign n29747 = controllable_BtoS_ACK0 & ~n29746;
  assign n29748 = ~n28017 & ~n28909;
  assign n29749 = ~i_RtoB_ACK0 & ~n29748;
  assign n29750 = ~n23129 & ~n29749;
  assign n29751 = controllable_DEQ & ~n29750;
  assign n29752 = ~n28022 & ~n28917;
  assign n29753 = ~i_RtoB_ACK0 & ~n29752;
  assign n29754 = ~n23135 & ~n29753;
  assign n29755 = ~controllable_DEQ & ~n29754;
  assign n29756 = ~n29751 & ~n29755;
  assign n29757 = i_FULL & ~n29756;
  assign n29758 = ~n28029 & ~n28927;
  assign n29759 = ~i_RtoB_ACK0 & ~n29758;
  assign n29760 = ~n23135 & ~n29759;
  assign n29761 = ~controllable_DEQ & ~n29760;
  assign n29762 = ~n23133 & ~n29761;
  assign n29763 = ~i_FULL & ~n29762;
  assign n29764 = ~n29757 & ~n29763;
  assign n29765 = i_nEMPTY & ~n29764;
  assign n29766 = ~n28038 & ~n28939;
  assign n29767 = ~i_RtoB_ACK0 & ~n29766;
  assign n29768 = ~n23147 & ~n29767;
  assign n29769 = ~controllable_DEQ & ~n29768;
  assign n29770 = ~n23145 & ~n29769;
  assign n29771 = i_FULL & ~n29770;
  assign n29772 = ~n28048 & ~n28909;
  assign n29773 = ~i_RtoB_ACK0 & ~n29772;
  assign n29774 = ~n23129 & ~n29773;
  assign n29775 = ~controllable_DEQ & ~n29774;
  assign n29776 = ~n23157 & ~n29775;
  assign n29777 = ~i_FULL & ~n29776;
  assign n29778 = ~n29771 & ~n29777;
  assign n29779 = ~i_nEMPTY & ~n29778;
  assign n29780 = ~n29765 & ~n29779;
  assign n29781 = ~controllable_BtoS_ACK0 & ~n29780;
  assign n29782 = ~n29747 & ~n29781;
  assign n29783 = n4465 & ~n29782;
  assign n29784 = ~n28064 & ~n28963;
  assign n29785 = ~i_RtoB_ACK0 & ~n29784;
  assign n29786 = ~n23129 & ~n29785;
  assign n29787 = controllable_DEQ & ~n29786;
  assign n29788 = ~n28069 & ~n28971;
  assign n29789 = ~i_RtoB_ACK0 & ~n29788;
  assign n29790 = ~n23135 & ~n29789;
  assign n29791 = ~controllable_DEQ & ~n29790;
  assign n29792 = ~n29787 & ~n29791;
  assign n29793 = i_FULL & ~n29792;
  assign n29794 = ~n28076 & ~n28981;
  assign n29795 = ~i_RtoB_ACK0 & ~n29794;
  assign n29796 = ~n23135 & ~n29795;
  assign n29797 = ~controllable_DEQ & ~n29796;
  assign n29798 = ~n23133 & ~n29797;
  assign n29799 = ~i_FULL & ~n29798;
  assign n29800 = ~n29793 & ~n29799;
  assign n29801 = i_nEMPTY & ~n29800;
  assign n29802 = ~n28085 & ~n28993;
  assign n29803 = ~i_RtoB_ACK0 & ~n29802;
  assign n29804 = ~n23147 & ~n29803;
  assign n29805 = ~controllable_DEQ & ~n29804;
  assign n29806 = ~n23145 & ~n29805;
  assign n29807 = i_FULL & ~n29806;
  assign n29808 = ~n28093 & ~n28963;
  assign n29809 = ~i_RtoB_ACK0 & ~n29808;
  assign n29810 = ~n23129 & ~n29809;
  assign n29811 = ~controllable_DEQ & ~n29810;
  assign n29812 = ~n23157 & ~n29811;
  assign n29813 = ~i_FULL & ~n29812;
  assign n29814 = ~n29807 & ~n29813;
  assign n29815 = ~i_nEMPTY & ~n29814;
  assign n29816 = ~n29801 & ~n29815;
  assign n29817 = ~controllable_BtoS_ACK0 & ~n29816;
  assign n29818 = ~n23127 & ~n29817;
  assign n29819 = ~n4465 & ~n29818;
  assign n29820 = ~n29783 & ~n29819;
  assign n29821 = ~i_StoB_REQ10 & ~n29820;
  assign n29822 = ~n29713 & ~n29821;
  assign n29823 = controllable_BtoS_ACK10 & ~n29822;
  assign n29824 = ~n17050 & ~n28112;
  assign n29825 = i_RtoB_ACK0 & ~n29824;
  assign n29826 = controllable_BtoR_REQ0 & ~n19387;
  assign n29827 = ~n28118 & ~n29826;
  assign n29828 = ~i_RtoB_ACK0 & ~n29827;
  assign n29829 = ~n29825 & ~n29828;
  assign n29830 = controllable_DEQ & ~n29829;
  assign n29831 = ~n17058 & ~n28125;
  assign n29832 = i_RtoB_ACK0 & ~n29831;
  assign n29833 = controllable_BtoR_REQ0 & ~n19396;
  assign n29834 = ~n27977 & ~n29833;
  assign n29835 = ~i_RtoB_ACK0 & ~n29834;
  assign n29836 = ~n29832 & ~n29835;
  assign n29837 = ~controllable_DEQ & ~n29836;
  assign n29838 = ~n29830 & ~n29837;
  assign n29839 = i_FULL & ~n29838;
  assign n29840 = controllable_BtoR_REQ0 & ~n17621;
  assign n29841 = ~n28135 & ~n29840;
  assign n29842 = ~i_RtoB_ACK0 & ~n29841;
  assign n29843 = ~n29825 & ~n29842;
  assign n29844 = controllable_DEQ & ~n29843;
  assign n29845 = controllable_BtoR_REQ0 & ~n19412;
  assign n29846 = ~n27984 & ~n29845;
  assign n29847 = ~i_RtoB_ACK0 & ~n29846;
  assign n29848 = ~n29832 & ~n29847;
  assign n29849 = ~controllable_DEQ & ~n29848;
  assign n29850 = ~n29844 & ~n29849;
  assign n29851 = ~i_FULL & ~n29850;
  assign n29852 = ~n29839 & ~n29851;
  assign n29853 = i_nEMPTY & ~n29852;
  assign n29854 = controllable_BtoR_REQ0 & ~n17646;
  assign n29855 = ~n28149 & ~n29854;
  assign n29856 = ~i_RtoB_ACK0 & ~n29855;
  assign n29857 = ~n15604 & ~n29856;
  assign n29858 = controllable_DEQ & ~n29857;
  assign n29859 = ~n17068 & ~n28112;
  assign n29860 = i_RtoB_ACK0 & ~n29859;
  assign n29861 = controllable_BtoR_REQ0 & ~n19430;
  assign n29862 = ~n27993 & ~n29861;
  assign n29863 = ~i_RtoB_ACK0 & ~n29862;
  assign n29864 = ~n29860 & ~n29863;
  assign n29865 = ~controllable_DEQ & ~n29864;
  assign n29866 = ~n29858 & ~n29865;
  assign n29867 = i_FULL & ~n29866;
  assign n29868 = controllable_BtoR_REQ0 & ~n17668;
  assign n29869 = ~n28159 & ~n29868;
  assign n29870 = ~i_RtoB_ACK0 & ~n29869;
  assign n29871 = ~n15619 & ~n29870;
  assign n29872 = controllable_DEQ & ~n29871;
  assign n29873 = ~controllable_DEQ & ~n29829;
  assign n29874 = ~n29872 & ~n29873;
  assign n29875 = ~i_FULL & ~n29874;
  assign n29876 = ~n29867 & ~n29875;
  assign n29877 = ~i_nEMPTY & ~n29876;
  assign n29878 = ~n29853 & ~n29877;
  assign n29879 = controllable_BtoS_ACK0 & ~n29878;
  assign n29880 = ~n18522 & ~n28173;
  assign n29881 = i_RtoB_ACK0 & ~n29880;
  assign n29882 = controllable_BtoR_REQ0 & ~n19453;
  assign n29883 = ~n28179 & ~n29882;
  assign n29884 = ~i_RtoB_ACK0 & ~n29883;
  assign n29885 = ~n29881 & ~n29884;
  assign n29886 = controllable_DEQ & ~n29885;
  assign n29887 = ~n18530 & ~n28186;
  assign n29888 = i_RtoB_ACK0 & ~n29887;
  assign n29889 = controllable_BtoR_REQ0 & ~n19462;
  assign n29890 = ~n28022 & ~n29889;
  assign n29891 = ~i_RtoB_ACK0 & ~n29890;
  assign n29892 = ~n29888 & ~n29891;
  assign n29893 = ~controllable_DEQ & ~n29892;
  assign n29894 = ~n29886 & ~n29893;
  assign n29895 = i_FULL & ~n29894;
  assign n29896 = controllable_BtoR_REQ0 & ~n17700;
  assign n29897 = ~n28196 & ~n29896;
  assign n29898 = ~i_RtoB_ACK0 & ~n29897;
  assign n29899 = ~n29881 & ~n29898;
  assign n29900 = controllable_DEQ & ~n29899;
  assign n29901 = controllable_BtoR_REQ0 & ~n19478;
  assign n29902 = ~n28029 & ~n29901;
  assign n29903 = ~i_RtoB_ACK0 & ~n29902;
  assign n29904 = ~n29888 & ~n29903;
  assign n29905 = ~controllable_DEQ & ~n29904;
  assign n29906 = ~n29900 & ~n29905;
  assign n29907 = ~i_FULL & ~n29906;
  assign n29908 = ~n29895 & ~n29907;
  assign n29909 = i_nEMPTY & ~n29908;
  assign n29910 = controllable_BtoR_REQ0 & ~n17736;
  assign n29911 = ~n28210 & ~n29910;
  assign n29912 = ~i_RtoB_ACK0 & ~n29911;
  assign n29913 = ~n17925 & ~n29912;
  assign n29914 = controllable_DEQ & ~n29913;
  assign n29915 = ~n18548 & ~n28173;
  assign n29916 = i_RtoB_ACK0 & ~n29915;
  assign n29917 = controllable_BtoR_REQ0 & ~n19496;
  assign n29918 = ~n28038 & ~n29917;
  assign n29919 = ~i_RtoB_ACK0 & ~n29918;
  assign n29920 = ~n29916 & ~n29919;
  assign n29921 = ~controllable_DEQ & ~n29920;
  assign n29922 = ~n29914 & ~n29921;
  assign n29923 = i_FULL & ~n29922;
  assign n29924 = controllable_BtoR_REQ0 & ~n17769;
  assign n29925 = ~n28220 & ~n29924;
  assign n29926 = ~i_RtoB_ACK0 & ~n29925;
  assign n29927 = ~n17943 & ~n29926;
  assign n29928 = controllable_DEQ & ~n29927;
  assign n29929 = ~controllable_DEQ & ~n29885;
  assign n29930 = ~n29928 & ~n29929;
  assign n29931 = ~i_FULL & ~n29930;
  assign n29932 = ~n29923 & ~n29931;
  assign n29933 = ~i_nEMPTY & ~n29932;
  assign n29934 = ~n29909 & ~n29933;
  assign n29935 = ~controllable_BtoS_ACK0 & ~n29934;
  assign n29936 = ~n29879 & ~n29935;
  assign n29937 = n4465 & ~n29936;
  assign n29938 = controllable_BtoR_REQ0 & ~n17627;
  assign n29939 = ~n11253 & ~n29938;
  assign n29940 = ~i_RtoB_ACK0 & ~n29939;
  assign n29941 = ~n29832 & ~n29940;
  assign n29942 = ~controllable_DEQ & ~n29941;
  assign n29943 = ~n29844 & ~n29942;
  assign n29944 = i_nEMPTY & ~n29943;
  assign n29945 = controllable_BtoR_REQ0 & ~n17612;
  assign n29946 = ~n11270 & ~n29945;
  assign n29947 = ~i_RtoB_ACK0 & ~n29946;
  assign n29948 = ~n29860 & ~n29947;
  assign n29949 = ~controllable_DEQ & ~n29948;
  assign n29950 = ~n29858 & ~n29949;
  assign n29951 = i_FULL & ~n29950;
  assign n29952 = ~controllable_DEQ & ~n29843;
  assign n29953 = ~n29872 & ~n29952;
  assign n29954 = ~i_FULL & ~n29953;
  assign n29955 = ~n29951 & ~n29954;
  assign n29956 = ~i_nEMPTY & ~n29955;
  assign n29957 = ~n29944 & ~n29956;
  assign n29958 = controllable_BtoS_ACK0 & ~n29957;
  assign n29959 = controllable_BtoR_REQ0 & ~n19314;
  assign n29960 = ~n28252 & ~n29959;
  assign n29961 = ~i_RtoB_ACK0 & ~n29960;
  assign n29962 = ~n29881 & ~n29961;
  assign n29963 = controllable_DEQ & ~n29962;
  assign n29964 = controllable_BtoR_REQ0 & ~n19322;
  assign n29965 = ~n28069 & ~n29964;
  assign n29966 = ~i_RtoB_ACK0 & ~n29965;
  assign n29967 = ~n29888 & ~n29966;
  assign n29968 = ~controllable_DEQ & ~n29967;
  assign n29969 = ~n29963 & ~n29968;
  assign n29970 = i_FULL & ~n29969;
  assign n29971 = controllable_BtoR_REQ0 & ~n19336;
  assign n29972 = ~n28076 & ~n29971;
  assign n29973 = ~i_RtoB_ACK0 & ~n29972;
  assign n29974 = ~n29888 & ~n29973;
  assign n29975 = ~controllable_DEQ & ~n29974;
  assign n29976 = ~n29900 & ~n29975;
  assign n29977 = ~i_FULL & ~n29976;
  assign n29978 = ~n29970 & ~n29977;
  assign n29979 = i_nEMPTY & ~n29978;
  assign n29980 = controllable_BtoR_REQ0 & ~n19352;
  assign n29981 = ~n28085 & ~n29980;
  assign n29982 = ~i_RtoB_ACK0 & ~n29981;
  assign n29983 = ~n29916 & ~n29982;
  assign n29984 = ~controllable_DEQ & ~n29983;
  assign n29985 = ~n29914 & ~n29984;
  assign n29986 = i_FULL & ~n29985;
  assign n29987 = ~controllable_DEQ & ~n29962;
  assign n29988 = ~n29928 & ~n29987;
  assign n29989 = ~i_FULL & ~n29988;
  assign n29990 = ~n29986 & ~n29989;
  assign n29991 = ~i_nEMPTY & ~n29990;
  assign n29992 = ~n29979 & ~n29991;
  assign n29993 = ~controllable_BtoS_ACK0 & ~n29992;
  assign n29994 = ~n29958 & ~n29993;
  assign n29995 = ~n4465 & ~n29994;
  assign n29996 = ~n29937 & ~n29995;
  assign n29997 = i_StoB_REQ10 & ~n29996;
  assign n29998 = ~n29821 & ~n29997;
  assign n29999 = ~controllable_BtoS_ACK10 & ~n29998;
  assign n30000 = ~n29823 & ~n29999;
  assign n30001 = n4464 & ~n30000;
  assign n30002 = ~n28288 & ~n29157;
  assign n30003 = ~i_RtoB_ACK0 & ~n30002;
  assign n30004 = ~n20977 & ~n30003;
  assign n30005 = controllable_DEQ & ~n30004;
  assign n30006 = ~n26438 & ~n29165;
  assign n30007 = ~i_RtoB_ACK0 & ~n30006;
  assign n30008 = ~n20983 & ~n30007;
  assign n30009 = ~controllable_DEQ & ~n30008;
  assign n30010 = ~n30005 & ~n30009;
  assign n30011 = i_FULL & ~n30010;
  assign n30012 = ~n28299 & ~n29175;
  assign n30013 = ~i_RtoB_ACK0 & ~n30012;
  assign n30014 = ~n20983 & ~n30013;
  assign n30015 = ~controllable_DEQ & ~n30014;
  assign n30016 = ~n20981 & ~n30015;
  assign n30017 = ~i_FULL & ~n30016;
  assign n30018 = ~n30011 & ~n30017;
  assign n30019 = i_nEMPTY & ~n30018;
  assign n30020 = ~n26461 & ~n29187;
  assign n30021 = ~i_RtoB_ACK0 & ~n30020;
  assign n30022 = ~n20977 & ~n30021;
  assign n30023 = ~controllable_DEQ & ~n30022;
  assign n30024 = ~n20993 & ~n30023;
  assign n30025 = i_FULL & ~n30024;
  assign n30026 = ~n28314 & ~n29157;
  assign n30027 = ~i_RtoB_ACK0 & ~n30026;
  assign n30028 = ~n20977 & ~n30027;
  assign n30029 = ~controllable_DEQ & ~n30028;
  assign n30030 = ~n21003 & ~n30029;
  assign n30031 = ~i_FULL & ~n30030;
  assign n30032 = ~n30025 & ~n30031;
  assign n30033 = ~i_nEMPTY & ~n30032;
  assign n30034 = ~n30019 & ~n30033;
  assign n30035 = controllable_BtoS_ACK0 & ~n30034;
  assign n30036 = ~n28327 & ~n29207;
  assign n30037 = ~i_RtoB_ACK0 & ~n30036;
  assign n30038 = ~n29625 & ~n30037;
  assign n30039 = controllable_DEQ & ~n30038;
  assign n30040 = ~n26486 & ~n29215;
  assign n30041 = ~i_RtoB_ACK0 & ~n30040;
  assign n30042 = ~n29631 & ~n30041;
  assign n30043 = ~controllable_DEQ & ~n30042;
  assign n30044 = ~n30039 & ~n30043;
  assign n30045 = i_FULL & ~n30044;
  assign n30046 = ~n28338 & ~n29225;
  assign n30047 = ~i_RtoB_ACK0 & ~n30046;
  assign n30048 = ~n29631 & ~n30047;
  assign n30049 = ~controllable_DEQ & ~n30048;
  assign n30050 = ~n29641 & ~n30049;
  assign n30051 = ~i_FULL & ~n30050;
  assign n30052 = ~n30045 & ~n30051;
  assign n30053 = i_nEMPTY & ~n30052;
  assign n30054 = ~n26509 & ~n29237;
  assign n30055 = ~i_RtoB_ACK0 & ~n30054;
  assign n30056 = ~n29625 & ~n30055;
  assign n30057 = ~controllable_DEQ & ~n30056;
  assign n30058 = ~n29653 & ~n30057;
  assign n30059 = i_FULL & ~n30058;
  assign n30060 = ~n28353 & ~n29207;
  assign n30061 = ~i_RtoB_ACK0 & ~n30060;
  assign n30062 = ~n29625 & ~n30061;
  assign n30063 = ~controllable_DEQ & ~n30062;
  assign n30064 = ~n29663 & ~n30063;
  assign n30065 = ~i_FULL & ~n30064;
  assign n30066 = ~n30059 & ~n30065;
  assign n30067 = ~i_nEMPTY & ~n30066;
  assign n30068 = ~n30053 & ~n30067;
  assign n30069 = ~controllable_BtoS_ACK0 & ~n30068;
  assign n30070 = ~n30035 & ~n30069;
  assign n30071 = n4465 & ~n30070;
  assign n30072 = ~n21013 & ~n30069;
  assign n30073 = ~n4465 & ~n30072;
  assign n30074 = ~n30071 & ~n30073;
  assign n30075 = i_StoB_REQ10 & ~n30074;
  assign n30076 = ~n28373 & ~n29263;
  assign n30077 = ~i_RtoB_ACK0 & ~n30076;
  assign n30078 = ~n23089 & ~n30077;
  assign n30079 = controllable_DEQ & ~n30078;
  assign n30080 = ~n28378 & ~n29271;
  assign n30081 = ~i_RtoB_ACK0 & ~n30080;
  assign n30082 = ~n23095 & ~n30081;
  assign n30083 = ~controllable_DEQ & ~n30082;
  assign n30084 = ~n30079 & ~n30083;
  assign n30085 = i_FULL & ~n30084;
  assign n30086 = ~n28385 & ~n29281;
  assign n30087 = ~i_RtoB_ACK0 & ~n30086;
  assign n30088 = ~n23095 & ~n30087;
  assign n30089 = ~controllable_DEQ & ~n30088;
  assign n30090 = ~n23093 & ~n30089;
  assign n30091 = ~i_FULL & ~n30090;
  assign n30092 = ~n30085 & ~n30091;
  assign n30093 = i_nEMPTY & ~n30092;
  assign n30094 = ~n28394 & ~n29293;
  assign n30095 = ~i_RtoB_ACK0 & ~n30094;
  assign n30096 = ~n23107 & ~n30095;
  assign n30097 = ~controllable_DEQ & ~n30096;
  assign n30098 = ~n23105 & ~n30097;
  assign n30099 = i_FULL & ~n30098;
  assign n30100 = ~n28402 & ~n29263;
  assign n30101 = ~i_RtoB_ACK0 & ~n30100;
  assign n30102 = ~n23089 & ~n30101;
  assign n30103 = ~controllable_DEQ & ~n30102;
  assign n30104 = ~n23117 & ~n30103;
  assign n30105 = ~i_FULL & ~n30104;
  assign n30106 = ~n30099 & ~n30105;
  assign n30107 = ~i_nEMPTY & ~n30106;
  assign n30108 = ~n30093 & ~n30107;
  assign n30109 = controllable_BtoS_ACK0 & ~n30108;
  assign n30110 = ~n28416 & ~n29313;
  assign n30111 = ~i_RtoB_ACK0 & ~n30110;
  assign n30112 = ~n23129 & ~n30111;
  assign n30113 = controllable_DEQ & ~n30112;
  assign n30114 = ~n28421 & ~n29321;
  assign n30115 = ~i_RtoB_ACK0 & ~n30114;
  assign n30116 = ~n23135 & ~n30115;
  assign n30117 = ~controllable_DEQ & ~n30116;
  assign n30118 = ~n30113 & ~n30117;
  assign n30119 = i_FULL & ~n30118;
  assign n30120 = ~n28428 & ~n29331;
  assign n30121 = ~i_RtoB_ACK0 & ~n30120;
  assign n30122 = ~n23135 & ~n30121;
  assign n30123 = ~controllable_DEQ & ~n30122;
  assign n30124 = ~n23133 & ~n30123;
  assign n30125 = ~i_FULL & ~n30124;
  assign n30126 = ~n30119 & ~n30125;
  assign n30127 = i_nEMPTY & ~n30126;
  assign n30128 = ~n28437 & ~n29343;
  assign n30129 = ~i_RtoB_ACK0 & ~n30128;
  assign n30130 = ~n23147 & ~n30129;
  assign n30131 = ~controllable_DEQ & ~n30130;
  assign n30132 = ~n23145 & ~n30131;
  assign n30133 = i_FULL & ~n30132;
  assign n30134 = ~n28445 & ~n29313;
  assign n30135 = ~i_RtoB_ACK0 & ~n30134;
  assign n30136 = ~n23129 & ~n30135;
  assign n30137 = ~controllable_DEQ & ~n30136;
  assign n30138 = ~n23157 & ~n30137;
  assign n30139 = ~i_FULL & ~n30138;
  assign n30140 = ~n30133 & ~n30139;
  assign n30141 = ~i_nEMPTY & ~n30140;
  assign n30142 = ~n30127 & ~n30141;
  assign n30143 = ~controllable_BtoS_ACK0 & ~n30142;
  assign n30144 = ~n30109 & ~n30143;
  assign n30145 = n4465 & ~n30144;
  assign n30146 = ~n23127 & ~n30143;
  assign n30147 = ~n4465 & ~n30146;
  assign n30148 = ~n30145 & ~n30147;
  assign n30149 = ~i_StoB_REQ10 & ~n30148;
  assign n30150 = ~n30075 & ~n30149;
  assign n30151 = controllable_BtoS_ACK10 & ~n30150;
  assign n30152 = controllable_BtoR_REQ0 & ~n20005;
  assign n30153 = ~n28467 & ~n30152;
  assign n30154 = ~i_RtoB_ACK0 & ~n30153;
  assign n30155 = ~n29825 & ~n30154;
  assign n30156 = controllable_DEQ & ~n30155;
  assign n30157 = controllable_BtoR_REQ0 & ~n20014;
  assign n30158 = ~n28378 & ~n30157;
  assign n30159 = ~i_RtoB_ACK0 & ~n30158;
  assign n30160 = ~n29832 & ~n30159;
  assign n30161 = ~controllable_DEQ & ~n30160;
  assign n30162 = ~n30156 & ~n30161;
  assign n30163 = i_FULL & ~n30162;
  assign n30164 = controllable_BtoR_REQ0 & ~n20030;
  assign n30165 = ~n28385 & ~n30164;
  assign n30166 = ~i_RtoB_ACK0 & ~n30165;
  assign n30167 = ~n29832 & ~n30166;
  assign n30168 = ~controllable_DEQ & ~n30167;
  assign n30169 = ~n29844 & ~n30168;
  assign n30170 = ~i_FULL & ~n30169;
  assign n30171 = ~n30163 & ~n30170;
  assign n30172 = i_nEMPTY & ~n30171;
  assign n30173 = controllable_BtoR_REQ0 & ~n20048;
  assign n30174 = ~n28394 & ~n30173;
  assign n30175 = ~i_RtoB_ACK0 & ~n30174;
  assign n30176 = ~n29860 & ~n30175;
  assign n30177 = ~controllable_DEQ & ~n30176;
  assign n30178 = ~n29858 & ~n30177;
  assign n30179 = i_FULL & ~n30178;
  assign n30180 = ~controllable_DEQ & ~n30155;
  assign n30181 = ~n29872 & ~n30180;
  assign n30182 = ~i_FULL & ~n30181;
  assign n30183 = ~n30179 & ~n30182;
  assign n30184 = ~i_nEMPTY & ~n30183;
  assign n30185 = ~n30172 & ~n30184;
  assign n30186 = controllable_BtoS_ACK0 & ~n30185;
  assign n30187 = controllable_BtoR_REQ0 & ~n19932;
  assign n30188 = ~n28496 & ~n30187;
  assign n30189 = ~i_RtoB_ACK0 & ~n30188;
  assign n30190 = ~n29881 & ~n30189;
  assign n30191 = controllable_DEQ & ~n30190;
  assign n30192 = controllable_BtoR_REQ0 & ~n19940;
  assign n30193 = ~n28421 & ~n30192;
  assign n30194 = ~i_RtoB_ACK0 & ~n30193;
  assign n30195 = ~n29888 & ~n30194;
  assign n30196 = ~controllable_DEQ & ~n30195;
  assign n30197 = ~n30191 & ~n30196;
  assign n30198 = i_FULL & ~n30197;
  assign n30199 = controllable_BtoR_REQ0 & ~n19954;
  assign n30200 = ~n28428 & ~n30199;
  assign n30201 = ~i_RtoB_ACK0 & ~n30200;
  assign n30202 = ~n29888 & ~n30201;
  assign n30203 = ~controllable_DEQ & ~n30202;
  assign n30204 = ~n29900 & ~n30203;
  assign n30205 = ~i_FULL & ~n30204;
  assign n30206 = ~n30198 & ~n30205;
  assign n30207 = i_nEMPTY & ~n30206;
  assign n30208 = controllable_BtoR_REQ0 & ~n19970;
  assign n30209 = ~n28437 & ~n30208;
  assign n30210 = ~i_RtoB_ACK0 & ~n30209;
  assign n30211 = ~n29916 & ~n30210;
  assign n30212 = ~controllable_DEQ & ~n30211;
  assign n30213 = ~n29914 & ~n30212;
  assign n30214 = i_FULL & ~n30213;
  assign n30215 = ~controllable_DEQ & ~n30190;
  assign n30216 = ~n29928 & ~n30215;
  assign n30217 = ~i_FULL & ~n30216;
  assign n30218 = ~n30214 & ~n30217;
  assign n30219 = ~i_nEMPTY & ~n30218;
  assign n30220 = ~n30207 & ~n30219;
  assign n30221 = ~controllable_BtoS_ACK0 & ~n30220;
  assign n30222 = ~n30186 & ~n30221;
  assign n30223 = n4465 & ~n30222;
  assign n30224 = ~n29958 & ~n30221;
  assign n30225 = ~n4465 & ~n30224;
  assign n30226 = ~n30223 & ~n30225;
  assign n30227 = i_StoB_REQ10 & ~n30226;
  assign n30228 = ~n30149 & ~n30227;
  assign n30229 = ~controllable_BtoS_ACK10 & ~n30228;
  assign n30230 = ~n30151 & ~n30229;
  assign n30231 = ~n4464 & ~n30230;
  assign n30232 = ~n30001 & ~n30231;
  assign n30233 = n4463 & ~n30232;
  assign n30234 = ~n5247 & ~n28681;
  assign n30235 = ~i_RtoB_ACK0 & ~n30234;
  assign n30236 = ~n20977 & ~n30235;
  assign n30237 = controllable_DEQ & ~n30236;
  assign n30238 = ~n5260 & ~n28689;
  assign n30239 = ~i_RtoB_ACK0 & ~n30238;
  assign n30240 = ~n20983 & ~n30239;
  assign n30241 = ~controllable_DEQ & ~n30240;
  assign n30242 = ~n30237 & ~n30241;
  assign n30243 = i_FULL & ~n30242;
  assign n30244 = ~n5260 & ~n28699;
  assign n30245 = ~i_RtoB_ACK0 & ~n30244;
  assign n30246 = ~n20983 & ~n30245;
  assign n30247 = ~controllable_DEQ & ~n30246;
  assign n30248 = ~n20981 & ~n30247;
  assign n30249 = ~i_FULL & ~n30248;
  assign n30250 = ~n30243 & ~n30249;
  assign n30251 = i_nEMPTY & ~n30250;
  assign n30252 = ~n5282 & ~n28711;
  assign n30253 = ~i_RtoB_ACK0 & ~n30252;
  assign n30254 = ~n20977 & ~n30253;
  assign n30255 = ~controllable_DEQ & ~n30254;
  assign n30256 = ~n20993 & ~n30255;
  assign n30257 = i_FULL & ~n30256;
  assign n30258 = ~n5297 & ~n28681;
  assign n30259 = ~i_RtoB_ACK0 & ~n30258;
  assign n30260 = ~n20977 & ~n30259;
  assign n30261 = ~controllable_DEQ & ~n30260;
  assign n30262 = ~n21003 & ~n30261;
  assign n30263 = ~i_FULL & ~n30262;
  assign n30264 = ~n30257 & ~n30263;
  assign n30265 = ~i_nEMPTY & ~n30264;
  assign n30266 = ~n30251 & ~n30265;
  assign n30267 = controllable_BtoS_ACK0 & ~n30266;
  assign n30268 = ~n27880 & ~n28733;
  assign n30269 = ~i_RtoB_ACK0 & ~n30268;
  assign n30270 = ~n29625 & ~n30269;
  assign n30271 = controllable_DEQ & ~n30270;
  assign n30272 = ~n28534 & ~n28743;
  assign n30273 = ~i_RtoB_ACK0 & ~n30272;
  assign n30274 = ~n29631 & ~n30273;
  assign n30275 = ~controllable_DEQ & ~n30274;
  assign n30276 = ~n30271 & ~n30275;
  assign n30277 = i_FULL & ~n30276;
  assign n30278 = ~n28534 & ~n28761;
  assign n30279 = ~i_RtoB_ACK0 & ~n30278;
  assign n30280 = ~n29631 & ~n30279;
  assign n30281 = ~controllable_DEQ & ~n30280;
  assign n30282 = ~n29641 & ~n30281;
  assign n30283 = ~i_FULL & ~n30282;
  assign n30284 = ~n30277 & ~n30283;
  assign n30285 = i_nEMPTY & ~n30284;
  assign n30286 = ~n28541 & ~n28777;
  assign n30287 = ~i_RtoB_ACK0 & ~n30286;
  assign n30288 = ~n29625 & ~n30287;
  assign n30289 = ~controllable_DEQ & ~n30288;
  assign n30290 = ~n29653 & ~n30289;
  assign n30291 = i_FULL & ~n30290;
  assign n30292 = ~n28548 & ~n28733;
  assign n30293 = ~i_RtoB_ACK0 & ~n30292;
  assign n30294 = ~n29625 & ~n30293;
  assign n30295 = ~controllable_DEQ & ~n30294;
  assign n30296 = ~n29663 & ~n30295;
  assign n30297 = ~i_FULL & ~n30296;
  assign n30298 = ~n30291 & ~n30297;
  assign n30299 = ~i_nEMPTY & ~n30298;
  assign n30300 = ~n30285 & ~n30299;
  assign n30301 = ~controllable_BtoS_ACK0 & ~n30300;
  assign n30302 = ~n30267 & ~n30301;
  assign n30303 = n4465 & ~n30302;
  assign n30304 = ~n27880 & ~n28803;
  assign n30305 = ~i_RtoB_ACK0 & ~n30304;
  assign n30306 = ~n29625 & ~n30305;
  assign n30307 = controllable_DEQ & ~n30306;
  assign n30308 = ~n28534 & ~n28811;
  assign n30309 = ~i_RtoB_ACK0 & ~n30308;
  assign n30310 = ~n29631 & ~n30309;
  assign n30311 = ~controllable_DEQ & ~n30310;
  assign n30312 = ~n30307 & ~n30311;
  assign n30313 = i_FULL & ~n30312;
  assign n30314 = ~n28534 & ~n28821;
  assign n30315 = ~i_RtoB_ACK0 & ~n30314;
  assign n30316 = ~n29631 & ~n30315;
  assign n30317 = ~controllable_DEQ & ~n30316;
  assign n30318 = ~n29641 & ~n30317;
  assign n30319 = ~i_FULL & ~n30318;
  assign n30320 = ~n30313 & ~n30319;
  assign n30321 = i_nEMPTY & ~n30320;
  assign n30322 = ~n28541 & ~n28833;
  assign n30323 = ~i_RtoB_ACK0 & ~n30322;
  assign n30324 = ~n29625 & ~n30323;
  assign n30325 = ~controllable_DEQ & ~n30324;
  assign n30326 = ~n29653 & ~n30325;
  assign n30327 = i_FULL & ~n30326;
  assign n30328 = ~n28548 & ~n28803;
  assign n30329 = ~i_RtoB_ACK0 & ~n30328;
  assign n30330 = ~n29625 & ~n30329;
  assign n30331 = ~controllable_DEQ & ~n30330;
  assign n30332 = ~n29663 & ~n30331;
  assign n30333 = ~i_FULL & ~n30332;
  assign n30334 = ~n30327 & ~n30333;
  assign n30335 = ~i_nEMPTY & ~n30334;
  assign n30336 = ~n30321 & ~n30335;
  assign n30337 = ~controllable_BtoS_ACK0 & ~n30336;
  assign n30338 = ~n21013 & ~n30337;
  assign n30339 = ~n4465 & ~n30338;
  assign n30340 = ~n30303 & ~n30339;
  assign n30341 = i_StoB_REQ10 & ~n30340;
  assign n30342 = ~n11240 & ~n28857;
  assign n30343 = ~i_RtoB_ACK0 & ~n30342;
  assign n30344 = ~n23089 & ~n30343;
  assign n30345 = controllable_DEQ & ~n30344;
  assign n30346 = ~n11253 & ~n28865;
  assign n30347 = ~i_RtoB_ACK0 & ~n30346;
  assign n30348 = ~n23095 & ~n30347;
  assign n30349 = ~controllable_DEQ & ~n30348;
  assign n30350 = ~n30345 & ~n30349;
  assign n30351 = i_FULL & ~n30350;
  assign n30352 = ~n11253 & ~n28875;
  assign n30353 = ~i_RtoB_ACK0 & ~n30352;
  assign n30354 = ~n23095 & ~n30353;
  assign n30355 = ~controllable_DEQ & ~n30354;
  assign n30356 = ~n23093 & ~n30355;
  assign n30357 = ~i_FULL & ~n30356;
  assign n30358 = ~n30351 & ~n30357;
  assign n30359 = i_nEMPTY & ~n30358;
  assign n30360 = ~n11270 & ~n28887;
  assign n30361 = ~i_RtoB_ACK0 & ~n30360;
  assign n30362 = ~n23107 & ~n30361;
  assign n30363 = ~controllable_DEQ & ~n30362;
  assign n30364 = ~n23105 & ~n30363;
  assign n30365 = i_FULL & ~n30364;
  assign n30366 = ~n11286 & ~n28857;
  assign n30367 = ~i_RtoB_ACK0 & ~n30366;
  assign n30368 = ~n23089 & ~n30367;
  assign n30369 = ~controllable_DEQ & ~n30368;
  assign n30370 = ~n23117 & ~n30369;
  assign n30371 = ~i_FULL & ~n30370;
  assign n30372 = ~n30365 & ~n30371;
  assign n30373 = ~i_nEMPTY & ~n30372;
  assign n30374 = ~n30359 & ~n30373;
  assign n30375 = controllable_BtoS_ACK0 & ~n30374;
  assign n30376 = ~n11319 & ~n28909;
  assign n30377 = ~i_RtoB_ACK0 & ~n30376;
  assign n30378 = ~n23129 & ~n30377;
  assign n30379 = controllable_DEQ & ~n30378;
  assign n30380 = ~n11333 & ~n28917;
  assign n30381 = ~i_RtoB_ACK0 & ~n30380;
  assign n30382 = ~n23135 & ~n30381;
  assign n30383 = ~controllable_DEQ & ~n30382;
  assign n30384 = ~n30379 & ~n30383;
  assign n30385 = i_FULL & ~n30384;
  assign n30386 = ~n11333 & ~n28927;
  assign n30387 = ~i_RtoB_ACK0 & ~n30386;
  assign n30388 = ~n23135 & ~n30387;
  assign n30389 = ~controllable_DEQ & ~n30388;
  assign n30390 = ~n23133 & ~n30389;
  assign n30391 = ~i_FULL & ~n30390;
  assign n30392 = ~n30385 & ~n30391;
  assign n30393 = i_nEMPTY & ~n30392;
  assign n30394 = ~n11352 & ~n28939;
  assign n30395 = ~i_RtoB_ACK0 & ~n30394;
  assign n30396 = ~n23147 & ~n30395;
  assign n30397 = ~controllable_DEQ & ~n30396;
  assign n30398 = ~n23145 & ~n30397;
  assign n30399 = i_FULL & ~n30398;
  assign n30400 = ~n11368 & ~n28909;
  assign n30401 = ~i_RtoB_ACK0 & ~n30400;
  assign n30402 = ~n23129 & ~n30401;
  assign n30403 = ~controllable_DEQ & ~n30402;
  assign n30404 = ~n23157 & ~n30403;
  assign n30405 = ~i_FULL & ~n30404;
  assign n30406 = ~n30399 & ~n30405;
  assign n30407 = ~i_nEMPTY & ~n30406;
  assign n30408 = ~n30393 & ~n30407;
  assign n30409 = ~controllable_BtoS_ACK0 & ~n30408;
  assign n30410 = ~n30375 & ~n30409;
  assign n30411 = n4465 & ~n30410;
  assign n30412 = ~n11319 & ~n28963;
  assign n30413 = ~i_RtoB_ACK0 & ~n30412;
  assign n30414 = ~n23129 & ~n30413;
  assign n30415 = controllable_DEQ & ~n30414;
  assign n30416 = ~n11333 & ~n28971;
  assign n30417 = ~i_RtoB_ACK0 & ~n30416;
  assign n30418 = ~n23135 & ~n30417;
  assign n30419 = ~controllable_DEQ & ~n30418;
  assign n30420 = ~n30415 & ~n30419;
  assign n30421 = i_FULL & ~n30420;
  assign n30422 = ~n11333 & ~n28981;
  assign n30423 = ~i_RtoB_ACK0 & ~n30422;
  assign n30424 = ~n23135 & ~n30423;
  assign n30425 = ~controllable_DEQ & ~n30424;
  assign n30426 = ~n23133 & ~n30425;
  assign n30427 = ~i_FULL & ~n30426;
  assign n30428 = ~n30421 & ~n30427;
  assign n30429 = i_nEMPTY & ~n30428;
  assign n30430 = ~n11352 & ~n28993;
  assign n30431 = ~i_RtoB_ACK0 & ~n30430;
  assign n30432 = ~n23147 & ~n30431;
  assign n30433 = ~controllable_DEQ & ~n30432;
  assign n30434 = ~n23145 & ~n30433;
  assign n30435 = i_FULL & ~n30434;
  assign n30436 = ~n11368 & ~n28963;
  assign n30437 = ~i_RtoB_ACK0 & ~n30436;
  assign n30438 = ~n23129 & ~n30437;
  assign n30439 = ~controllable_DEQ & ~n30438;
  assign n30440 = ~n23157 & ~n30439;
  assign n30441 = ~i_FULL & ~n30440;
  assign n30442 = ~n30435 & ~n30441;
  assign n30443 = ~i_nEMPTY & ~n30442;
  assign n30444 = ~n30429 & ~n30443;
  assign n30445 = ~controllable_BtoS_ACK0 & ~n30444;
  assign n30446 = ~n23127 & ~n30445;
  assign n30447 = ~n4465 & ~n30446;
  assign n30448 = ~n30411 & ~n30447;
  assign n30449 = ~i_StoB_REQ10 & ~n30448;
  assign n30450 = ~n30341 & ~n30449;
  assign n30451 = controllable_BtoS_ACK10 & ~n30450;
  assign n30452 = ~n28135 & ~n29826;
  assign n30453 = ~i_RtoB_ACK0 & ~n30452;
  assign n30454 = ~n29825 & ~n30453;
  assign n30455 = controllable_DEQ & ~n30454;
  assign n30456 = ~n11253 & ~n29833;
  assign n30457 = ~i_RtoB_ACK0 & ~n30456;
  assign n30458 = ~n29832 & ~n30457;
  assign n30459 = ~controllable_DEQ & ~n30458;
  assign n30460 = ~n30455 & ~n30459;
  assign n30461 = i_FULL & ~n30460;
  assign n30462 = ~n11253 & ~n29845;
  assign n30463 = ~i_RtoB_ACK0 & ~n30462;
  assign n30464 = ~n29832 & ~n30463;
  assign n30465 = ~controllable_DEQ & ~n30464;
  assign n30466 = ~n29844 & ~n30465;
  assign n30467 = ~i_FULL & ~n30466;
  assign n30468 = ~n30461 & ~n30467;
  assign n30469 = i_nEMPTY & ~n30468;
  assign n30470 = ~n11270 & ~n29861;
  assign n30471 = ~i_RtoB_ACK0 & ~n30470;
  assign n30472 = ~n29860 & ~n30471;
  assign n30473 = ~controllable_DEQ & ~n30472;
  assign n30474 = ~n29858 & ~n30473;
  assign n30475 = i_FULL & ~n30474;
  assign n30476 = ~controllable_DEQ & ~n30454;
  assign n30477 = ~n29872 & ~n30476;
  assign n30478 = ~i_FULL & ~n30477;
  assign n30479 = ~n30475 & ~n30478;
  assign n30480 = ~i_nEMPTY & ~n30479;
  assign n30481 = ~n30469 & ~n30480;
  assign n30482 = controllable_BtoS_ACK0 & ~n30481;
  assign n30483 = ~n28196 & ~n29882;
  assign n30484 = ~i_RtoB_ACK0 & ~n30483;
  assign n30485 = ~n29881 & ~n30484;
  assign n30486 = controllable_DEQ & ~n30485;
  assign n30487 = ~n11333 & ~n29889;
  assign n30488 = ~i_RtoB_ACK0 & ~n30487;
  assign n30489 = ~n29888 & ~n30488;
  assign n30490 = ~controllable_DEQ & ~n30489;
  assign n30491 = ~n30486 & ~n30490;
  assign n30492 = i_FULL & ~n30491;
  assign n30493 = ~n11333 & ~n29901;
  assign n30494 = ~i_RtoB_ACK0 & ~n30493;
  assign n30495 = ~n29888 & ~n30494;
  assign n30496 = ~controllable_DEQ & ~n30495;
  assign n30497 = ~n29900 & ~n30496;
  assign n30498 = ~i_FULL & ~n30497;
  assign n30499 = ~n30492 & ~n30498;
  assign n30500 = i_nEMPTY & ~n30499;
  assign n30501 = ~n11352 & ~n29917;
  assign n30502 = ~i_RtoB_ACK0 & ~n30501;
  assign n30503 = ~n29916 & ~n30502;
  assign n30504 = ~controllable_DEQ & ~n30503;
  assign n30505 = ~n29914 & ~n30504;
  assign n30506 = i_FULL & ~n30505;
  assign n30507 = ~controllable_DEQ & ~n30485;
  assign n30508 = ~n29928 & ~n30507;
  assign n30509 = ~i_FULL & ~n30508;
  assign n30510 = ~n30506 & ~n30509;
  assign n30511 = ~i_nEMPTY & ~n30510;
  assign n30512 = ~n30500 & ~n30511;
  assign n30513 = ~controllable_BtoS_ACK0 & ~n30512;
  assign n30514 = ~n30482 & ~n30513;
  assign n30515 = n4465 & ~n30514;
  assign n30516 = ~n28196 & ~n29959;
  assign n30517 = ~i_RtoB_ACK0 & ~n30516;
  assign n30518 = ~n29881 & ~n30517;
  assign n30519 = controllable_DEQ & ~n30518;
  assign n30520 = ~n11333 & ~n29964;
  assign n30521 = ~i_RtoB_ACK0 & ~n30520;
  assign n30522 = ~n29888 & ~n30521;
  assign n30523 = ~controllable_DEQ & ~n30522;
  assign n30524 = ~n30519 & ~n30523;
  assign n30525 = i_FULL & ~n30524;
  assign n30526 = ~n11333 & ~n29971;
  assign n30527 = ~i_RtoB_ACK0 & ~n30526;
  assign n30528 = ~n29888 & ~n30527;
  assign n30529 = ~controllable_DEQ & ~n30528;
  assign n30530 = ~n29900 & ~n30529;
  assign n30531 = ~i_FULL & ~n30530;
  assign n30532 = ~n30525 & ~n30531;
  assign n30533 = i_nEMPTY & ~n30532;
  assign n30534 = ~n11352 & ~n29980;
  assign n30535 = ~i_RtoB_ACK0 & ~n30534;
  assign n30536 = ~n29916 & ~n30535;
  assign n30537 = ~controllable_DEQ & ~n30536;
  assign n30538 = ~n29914 & ~n30537;
  assign n30539 = i_FULL & ~n30538;
  assign n30540 = ~controllable_DEQ & ~n30518;
  assign n30541 = ~n29928 & ~n30540;
  assign n30542 = ~i_FULL & ~n30541;
  assign n30543 = ~n30539 & ~n30542;
  assign n30544 = ~i_nEMPTY & ~n30543;
  assign n30545 = ~n30533 & ~n30544;
  assign n30546 = ~controllable_BtoS_ACK0 & ~n30545;
  assign n30547 = ~n29958 & ~n30546;
  assign n30548 = ~n4465 & ~n30547;
  assign n30549 = ~n30515 & ~n30548;
  assign n30550 = i_StoB_REQ10 & ~n30549;
  assign n30551 = ~n30449 & ~n30550;
  assign n30552 = ~controllable_BtoS_ACK10 & ~n30551;
  assign n30553 = ~n30451 & ~n30552;
  assign n30554 = n4464 & ~n30553;
  assign n30555 = ~n5247 & ~n29157;
  assign n30556 = ~i_RtoB_ACK0 & ~n30555;
  assign n30557 = ~n20977 & ~n30556;
  assign n30558 = controllable_DEQ & ~n30557;
  assign n30559 = ~n5260 & ~n29165;
  assign n30560 = ~i_RtoB_ACK0 & ~n30559;
  assign n30561 = ~n20983 & ~n30560;
  assign n30562 = ~controllable_DEQ & ~n30561;
  assign n30563 = ~n30558 & ~n30562;
  assign n30564 = i_FULL & ~n30563;
  assign n30565 = ~n5260 & ~n29175;
  assign n30566 = ~i_RtoB_ACK0 & ~n30565;
  assign n30567 = ~n20983 & ~n30566;
  assign n30568 = ~controllable_DEQ & ~n30567;
  assign n30569 = ~n20981 & ~n30568;
  assign n30570 = ~i_FULL & ~n30569;
  assign n30571 = ~n30564 & ~n30570;
  assign n30572 = i_nEMPTY & ~n30571;
  assign n30573 = ~n5282 & ~n29187;
  assign n30574 = ~i_RtoB_ACK0 & ~n30573;
  assign n30575 = ~n20977 & ~n30574;
  assign n30576 = ~controllable_DEQ & ~n30575;
  assign n30577 = ~n20993 & ~n30576;
  assign n30578 = i_FULL & ~n30577;
  assign n30579 = ~n5297 & ~n29157;
  assign n30580 = ~i_RtoB_ACK0 & ~n30579;
  assign n30581 = ~n20977 & ~n30580;
  assign n30582 = ~controllable_DEQ & ~n30581;
  assign n30583 = ~n21003 & ~n30582;
  assign n30584 = ~i_FULL & ~n30583;
  assign n30585 = ~n30578 & ~n30584;
  assign n30586 = ~i_nEMPTY & ~n30585;
  assign n30587 = ~n30572 & ~n30586;
  assign n30588 = controllable_BtoS_ACK0 & ~n30587;
  assign n30589 = ~n27880 & ~n29207;
  assign n30590 = ~i_RtoB_ACK0 & ~n30589;
  assign n30591 = ~n29625 & ~n30590;
  assign n30592 = controllable_DEQ & ~n30591;
  assign n30593 = ~n28534 & ~n29215;
  assign n30594 = ~i_RtoB_ACK0 & ~n30593;
  assign n30595 = ~n29631 & ~n30594;
  assign n30596 = ~controllable_DEQ & ~n30595;
  assign n30597 = ~n30592 & ~n30596;
  assign n30598 = i_FULL & ~n30597;
  assign n30599 = ~n28534 & ~n29225;
  assign n30600 = ~i_RtoB_ACK0 & ~n30599;
  assign n30601 = ~n29631 & ~n30600;
  assign n30602 = ~controllable_DEQ & ~n30601;
  assign n30603 = ~n29641 & ~n30602;
  assign n30604 = ~i_FULL & ~n30603;
  assign n30605 = ~n30598 & ~n30604;
  assign n30606 = i_nEMPTY & ~n30605;
  assign n30607 = ~n28541 & ~n29237;
  assign n30608 = ~i_RtoB_ACK0 & ~n30607;
  assign n30609 = ~n29625 & ~n30608;
  assign n30610 = ~controllable_DEQ & ~n30609;
  assign n30611 = ~n29653 & ~n30610;
  assign n30612 = i_FULL & ~n30611;
  assign n30613 = ~n28548 & ~n29207;
  assign n30614 = ~i_RtoB_ACK0 & ~n30613;
  assign n30615 = ~n29625 & ~n30614;
  assign n30616 = ~controllable_DEQ & ~n30615;
  assign n30617 = ~n29663 & ~n30616;
  assign n30618 = ~i_FULL & ~n30617;
  assign n30619 = ~n30612 & ~n30618;
  assign n30620 = ~i_nEMPTY & ~n30619;
  assign n30621 = ~n30606 & ~n30620;
  assign n30622 = ~controllable_BtoS_ACK0 & ~n30621;
  assign n30623 = ~n30588 & ~n30622;
  assign n30624 = n4465 & ~n30623;
  assign n30625 = ~n21013 & ~n30622;
  assign n30626 = ~n4465 & ~n30625;
  assign n30627 = ~n30624 & ~n30626;
  assign n30628 = i_StoB_REQ10 & ~n30627;
  assign n30629 = ~n11240 & ~n29263;
  assign n30630 = ~i_RtoB_ACK0 & ~n30629;
  assign n30631 = ~n23089 & ~n30630;
  assign n30632 = controllable_DEQ & ~n30631;
  assign n30633 = ~n11253 & ~n29271;
  assign n30634 = ~i_RtoB_ACK0 & ~n30633;
  assign n30635 = ~n23095 & ~n30634;
  assign n30636 = ~controllable_DEQ & ~n30635;
  assign n30637 = ~n30632 & ~n30636;
  assign n30638 = i_FULL & ~n30637;
  assign n30639 = ~n11253 & ~n29281;
  assign n30640 = ~i_RtoB_ACK0 & ~n30639;
  assign n30641 = ~n23095 & ~n30640;
  assign n30642 = ~controllable_DEQ & ~n30641;
  assign n30643 = ~n23093 & ~n30642;
  assign n30644 = ~i_FULL & ~n30643;
  assign n30645 = ~n30638 & ~n30644;
  assign n30646 = i_nEMPTY & ~n30645;
  assign n30647 = ~n11270 & ~n29293;
  assign n30648 = ~i_RtoB_ACK0 & ~n30647;
  assign n30649 = ~n23107 & ~n30648;
  assign n30650 = ~controllable_DEQ & ~n30649;
  assign n30651 = ~n23105 & ~n30650;
  assign n30652 = i_FULL & ~n30651;
  assign n30653 = ~n11286 & ~n29263;
  assign n30654 = ~i_RtoB_ACK0 & ~n30653;
  assign n30655 = ~n23089 & ~n30654;
  assign n30656 = ~controllable_DEQ & ~n30655;
  assign n30657 = ~n23117 & ~n30656;
  assign n30658 = ~i_FULL & ~n30657;
  assign n30659 = ~n30652 & ~n30658;
  assign n30660 = ~i_nEMPTY & ~n30659;
  assign n30661 = ~n30646 & ~n30660;
  assign n30662 = controllable_BtoS_ACK0 & ~n30661;
  assign n30663 = ~n11319 & ~n29313;
  assign n30664 = ~i_RtoB_ACK0 & ~n30663;
  assign n30665 = ~n23129 & ~n30664;
  assign n30666 = controllable_DEQ & ~n30665;
  assign n30667 = ~n11333 & ~n29321;
  assign n30668 = ~i_RtoB_ACK0 & ~n30667;
  assign n30669 = ~n23135 & ~n30668;
  assign n30670 = ~controllable_DEQ & ~n30669;
  assign n30671 = ~n30666 & ~n30670;
  assign n30672 = i_FULL & ~n30671;
  assign n30673 = ~n11333 & ~n29331;
  assign n30674 = ~i_RtoB_ACK0 & ~n30673;
  assign n30675 = ~n23135 & ~n30674;
  assign n30676 = ~controllable_DEQ & ~n30675;
  assign n30677 = ~n23133 & ~n30676;
  assign n30678 = ~i_FULL & ~n30677;
  assign n30679 = ~n30672 & ~n30678;
  assign n30680 = i_nEMPTY & ~n30679;
  assign n30681 = ~n11352 & ~n29343;
  assign n30682 = ~i_RtoB_ACK0 & ~n30681;
  assign n30683 = ~n23147 & ~n30682;
  assign n30684 = ~controllable_DEQ & ~n30683;
  assign n30685 = ~n23145 & ~n30684;
  assign n30686 = i_FULL & ~n30685;
  assign n30687 = ~n11368 & ~n29313;
  assign n30688 = ~i_RtoB_ACK0 & ~n30687;
  assign n30689 = ~n23129 & ~n30688;
  assign n30690 = ~controllable_DEQ & ~n30689;
  assign n30691 = ~n23157 & ~n30690;
  assign n30692 = ~i_FULL & ~n30691;
  assign n30693 = ~n30686 & ~n30692;
  assign n30694 = ~i_nEMPTY & ~n30693;
  assign n30695 = ~n30680 & ~n30694;
  assign n30696 = ~controllable_BtoS_ACK0 & ~n30695;
  assign n30697 = ~n30662 & ~n30696;
  assign n30698 = n4465 & ~n30697;
  assign n30699 = ~n23127 & ~n30696;
  assign n30700 = ~n4465 & ~n30699;
  assign n30701 = ~n30698 & ~n30700;
  assign n30702 = ~i_StoB_REQ10 & ~n30701;
  assign n30703 = ~n30628 & ~n30702;
  assign n30704 = controllable_BtoS_ACK10 & ~n30703;
  assign n30705 = ~n28135 & ~n30152;
  assign n30706 = ~i_RtoB_ACK0 & ~n30705;
  assign n30707 = ~n29825 & ~n30706;
  assign n30708 = controllable_DEQ & ~n30707;
  assign n30709 = ~n11253 & ~n30157;
  assign n30710 = ~i_RtoB_ACK0 & ~n30709;
  assign n30711 = ~n29832 & ~n30710;
  assign n30712 = ~controllable_DEQ & ~n30711;
  assign n30713 = ~n30708 & ~n30712;
  assign n30714 = i_FULL & ~n30713;
  assign n30715 = ~n11253 & ~n30164;
  assign n30716 = ~i_RtoB_ACK0 & ~n30715;
  assign n30717 = ~n29832 & ~n30716;
  assign n30718 = ~controllable_DEQ & ~n30717;
  assign n30719 = ~n29844 & ~n30718;
  assign n30720 = ~i_FULL & ~n30719;
  assign n30721 = ~n30714 & ~n30720;
  assign n30722 = i_nEMPTY & ~n30721;
  assign n30723 = ~n11270 & ~n30173;
  assign n30724 = ~i_RtoB_ACK0 & ~n30723;
  assign n30725 = ~n29860 & ~n30724;
  assign n30726 = ~controllable_DEQ & ~n30725;
  assign n30727 = ~n29858 & ~n30726;
  assign n30728 = i_FULL & ~n30727;
  assign n30729 = ~controllable_DEQ & ~n30707;
  assign n30730 = ~n29872 & ~n30729;
  assign n30731 = ~i_FULL & ~n30730;
  assign n30732 = ~n30728 & ~n30731;
  assign n30733 = ~i_nEMPTY & ~n30732;
  assign n30734 = ~n30722 & ~n30733;
  assign n30735 = controllable_BtoS_ACK0 & ~n30734;
  assign n30736 = ~n28196 & ~n30187;
  assign n30737 = ~i_RtoB_ACK0 & ~n30736;
  assign n30738 = ~n29881 & ~n30737;
  assign n30739 = controllable_DEQ & ~n30738;
  assign n30740 = ~n11333 & ~n30192;
  assign n30741 = ~i_RtoB_ACK0 & ~n30740;
  assign n30742 = ~n29888 & ~n30741;
  assign n30743 = ~controllable_DEQ & ~n30742;
  assign n30744 = ~n30739 & ~n30743;
  assign n30745 = i_FULL & ~n30744;
  assign n30746 = ~n11333 & ~n30199;
  assign n30747 = ~i_RtoB_ACK0 & ~n30746;
  assign n30748 = ~n29888 & ~n30747;
  assign n30749 = ~controllable_DEQ & ~n30748;
  assign n30750 = ~n29900 & ~n30749;
  assign n30751 = ~i_FULL & ~n30750;
  assign n30752 = ~n30745 & ~n30751;
  assign n30753 = i_nEMPTY & ~n30752;
  assign n30754 = ~n11352 & ~n30208;
  assign n30755 = ~i_RtoB_ACK0 & ~n30754;
  assign n30756 = ~n29916 & ~n30755;
  assign n30757 = ~controllable_DEQ & ~n30756;
  assign n30758 = ~n29914 & ~n30757;
  assign n30759 = i_FULL & ~n30758;
  assign n30760 = ~controllable_DEQ & ~n30738;
  assign n30761 = ~n29928 & ~n30760;
  assign n30762 = ~i_FULL & ~n30761;
  assign n30763 = ~n30759 & ~n30762;
  assign n30764 = ~i_nEMPTY & ~n30763;
  assign n30765 = ~n30753 & ~n30764;
  assign n30766 = ~controllable_BtoS_ACK0 & ~n30765;
  assign n30767 = ~n30735 & ~n30766;
  assign n30768 = n4465 & ~n30767;
  assign n30769 = ~n29958 & ~n30766;
  assign n30770 = ~n4465 & ~n30769;
  assign n30771 = ~n30768 & ~n30770;
  assign n30772 = i_StoB_REQ10 & ~n30771;
  assign n30773 = ~n30702 & ~n30772;
  assign n30774 = ~controllable_BtoS_ACK10 & ~n30773;
  assign n30775 = ~n30704 & ~n30774;
  assign n30776 = ~n4464 & ~n30775;
  assign n30777 = ~n30554 & ~n30776;
  assign n30778 = ~n4463 & ~n30777;
  assign n30779 = ~n30233 & ~n30778;
  assign n30780 = n4462 & ~n30779;
  assign n30781 = ~n28534 & ~n29437;
  assign n30782 = ~i_RtoB_ACK0 & ~n30781;
  assign n30783 = ~n29631 & ~n30782;
  assign n30784 = ~controllable_DEQ & ~n30783;
  assign n30785 = ~n29641 & ~n30784;
  assign n30786 = i_nEMPTY & ~n30785;
  assign n30787 = ~n28541 & ~n29447;
  assign n30788 = ~i_RtoB_ACK0 & ~n30787;
  assign n30789 = ~n29625 & ~n30788;
  assign n30790 = ~controllable_DEQ & ~n30789;
  assign n30791 = ~n29653 & ~n30790;
  assign n30792 = i_FULL & ~n30791;
  assign n30793 = ~n28548 & ~n28753;
  assign n30794 = ~i_RtoB_ACK0 & ~n30793;
  assign n30795 = ~n29625 & ~n30794;
  assign n30796 = ~controllable_DEQ & ~n30795;
  assign n30797 = ~n29663 & ~n30796;
  assign n30798 = ~i_FULL & ~n30797;
  assign n30799 = ~n30792 & ~n30798;
  assign n30800 = ~i_nEMPTY & ~n30799;
  assign n30801 = ~n30786 & ~n30800;
  assign n30802 = ~controllable_BtoS_ACK0 & ~n30801;
  assign n30803 = ~n21013 & ~n30802;
  assign n30804 = i_StoB_REQ10 & ~n30803;
  assign n30805 = ~n23169 & ~n30804;
  assign n30806 = controllable_BtoS_ACK10 & ~n30805;
  assign n30807 = controllable_BtoR_REQ0 & ~n20369;
  assign n30808 = ~n28589 & ~n30807;
  assign n30809 = ~i_RtoB_ACK0 & ~n30808;
  assign n30810 = ~n29825 & ~n30809;
  assign n30811 = controllable_DEQ & ~n30810;
  assign n30812 = controllable_BtoR_REQ0 & ~n20378;
  assign n30813 = ~n28594 & ~n30812;
  assign n30814 = ~i_RtoB_ACK0 & ~n30813;
  assign n30815 = ~n29832 & ~n30814;
  assign n30816 = ~controllable_DEQ & ~n30815;
  assign n30817 = ~n30811 & ~n30816;
  assign n30818 = i_FULL & ~n30817;
  assign n30819 = controllable_BtoR_REQ0 & ~n20394;
  assign n30820 = ~n28601 & ~n30819;
  assign n30821 = ~i_RtoB_ACK0 & ~n30820;
  assign n30822 = ~n29832 & ~n30821;
  assign n30823 = ~controllable_DEQ & ~n30822;
  assign n30824 = ~n29844 & ~n30823;
  assign n30825 = ~i_FULL & ~n30824;
  assign n30826 = ~n30818 & ~n30825;
  assign n30827 = i_nEMPTY & ~n30826;
  assign n30828 = controllable_BtoR_REQ0 & ~n20412;
  assign n30829 = ~n28610 & ~n30828;
  assign n30830 = ~i_RtoB_ACK0 & ~n30829;
  assign n30831 = ~n29860 & ~n30830;
  assign n30832 = ~controllable_DEQ & ~n30831;
  assign n30833 = ~n29858 & ~n30832;
  assign n30834 = i_FULL & ~n30833;
  assign n30835 = ~controllable_DEQ & ~n30810;
  assign n30836 = ~n29872 & ~n30835;
  assign n30837 = ~i_FULL & ~n30836;
  assign n30838 = ~n30834 & ~n30837;
  assign n30839 = ~i_nEMPTY & ~n30838;
  assign n30840 = ~n30827 & ~n30839;
  assign n30841 = controllable_BtoS_ACK0 & ~n30840;
  assign n30842 = ~n29993 & ~n30841;
  assign n30843 = n4465 & ~n30842;
  assign n30844 = ~n29995 & ~n30843;
  assign n30845 = i_StoB_REQ10 & ~n30844;
  assign n30846 = ~n28631 & ~n29502;
  assign n30847 = ~i_RtoB_ACK0 & ~n30846;
  assign n30848 = ~n23089 & ~n30847;
  assign n30849 = controllable_DEQ & ~n30848;
  assign n30850 = ~n28594 & ~n29510;
  assign n30851 = ~i_RtoB_ACK0 & ~n30850;
  assign n30852 = ~n23095 & ~n30851;
  assign n30853 = ~controllable_DEQ & ~n30852;
  assign n30854 = ~n30849 & ~n30853;
  assign n30855 = i_FULL & ~n30854;
  assign n30856 = ~n28601 & ~n29520;
  assign n30857 = ~i_RtoB_ACK0 & ~n30856;
  assign n30858 = ~n23095 & ~n30857;
  assign n30859 = ~controllable_DEQ & ~n30858;
  assign n30860 = ~n23093 & ~n30859;
  assign n30861 = ~i_FULL & ~n30860;
  assign n30862 = ~n30855 & ~n30861;
  assign n30863 = i_nEMPTY & ~n30862;
  assign n30864 = ~n28610 & ~n29532;
  assign n30865 = ~i_RtoB_ACK0 & ~n30864;
  assign n30866 = ~n23107 & ~n30865;
  assign n30867 = ~controllable_DEQ & ~n30866;
  assign n30868 = ~n23105 & ~n30867;
  assign n30869 = i_FULL & ~n30868;
  assign n30870 = ~n28651 & ~n29502;
  assign n30871 = ~i_RtoB_ACK0 & ~n30870;
  assign n30872 = ~n23089 & ~n30871;
  assign n30873 = ~controllable_DEQ & ~n30872;
  assign n30874 = ~n23117 & ~n30873;
  assign n30875 = ~i_FULL & ~n30874;
  assign n30876 = ~n30869 & ~n30875;
  assign n30877 = ~i_nEMPTY & ~n30876;
  assign n30878 = ~n30863 & ~n30877;
  assign n30879 = controllable_BtoS_ACK0 & ~n30878;
  assign n30880 = ~n29817 & ~n30879;
  assign n30881 = n4465 & ~n30880;
  assign n30882 = ~n29819 & ~n30881;
  assign n30883 = ~i_StoB_REQ10 & ~n30882;
  assign n30884 = ~n30845 & ~n30883;
  assign n30885 = ~controllable_BtoS_ACK10 & ~n30884;
  assign n30886 = ~n30806 & ~n30885;
  assign n30887 = n4464 & ~n30886;
  assign n30888 = ~n30229 & ~n30806;
  assign n30889 = ~n4464 & ~n30888;
  assign n30890 = ~n30887 & ~n30889;
  assign n30891 = n4463 & ~n30890;
  assign n30892 = ~n28135 & ~n30807;
  assign n30893 = ~i_RtoB_ACK0 & ~n30892;
  assign n30894 = ~n29825 & ~n30893;
  assign n30895 = controllable_DEQ & ~n30894;
  assign n30896 = ~n11253 & ~n30812;
  assign n30897 = ~i_RtoB_ACK0 & ~n30896;
  assign n30898 = ~n29832 & ~n30897;
  assign n30899 = ~controllable_DEQ & ~n30898;
  assign n30900 = ~n30895 & ~n30899;
  assign n30901 = i_FULL & ~n30900;
  assign n30902 = ~n11253 & ~n30819;
  assign n30903 = ~i_RtoB_ACK0 & ~n30902;
  assign n30904 = ~n29832 & ~n30903;
  assign n30905 = ~controllable_DEQ & ~n30904;
  assign n30906 = ~n29844 & ~n30905;
  assign n30907 = ~i_FULL & ~n30906;
  assign n30908 = ~n30901 & ~n30907;
  assign n30909 = i_nEMPTY & ~n30908;
  assign n30910 = ~n11270 & ~n30828;
  assign n30911 = ~i_RtoB_ACK0 & ~n30910;
  assign n30912 = ~n29860 & ~n30911;
  assign n30913 = ~controllable_DEQ & ~n30912;
  assign n30914 = ~n29858 & ~n30913;
  assign n30915 = i_FULL & ~n30914;
  assign n30916 = ~controllable_DEQ & ~n30894;
  assign n30917 = ~n29872 & ~n30916;
  assign n30918 = ~i_FULL & ~n30917;
  assign n30919 = ~n30915 & ~n30918;
  assign n30920 = ~i_nEMPTY & ~n30919;
  assign n30921 = ~n30909 & ~n30920;
  assign n30922 = controllable_BtoS_ACK0 & ~n30921;
  assign n30923 = ~n30546 & ~n30922;
  assign n30924 = n4465 & ~n30923;
  assign n30925 = ~n30548 & ~n30924;
  assign n30926 = i_StoB_REQ10 & ~n30925;
  assign n30927 = ~n11240 & ~n29502;
  assign n30928 = ~i_RtoB_ACK0 & ~n30927;
  assign n30929 = ~n23089 & ~n30928;
  assign n30930 = controllable_DEQ & ~n30929;
  assign n30931 = ~n11253 & ~n29510;
  assign n30932 = ~i_RtoB_ACK0 & ~n30931;
  assign n30933 = ~n23095 & ~n30932;
  assign n30934 = ~controllable_DEQ & ~n30933;
  assign n30935 = ~n30930 & ~n30934;
  assign n30936 = i_FULL & ~n30935;
  assign n30937 = ~n11253 & ~n29520;
  assign n30938 = ~i_RtoB_ACK0 & ~n30937;
  assign n30939 = ~n23095 & ~n30938;
  assign n30940 = ~controllable_DEQ & ~n30939;
  assign n30941 = ~n23093 & ~n30940;
  assign n30942 = ~i_FULL & ~n30941;
  assign n30943 = ~n30936 & ~n30942;
  assign n30944 = i_nEMPTY & ~n30943;
  assign n30945 = ~n11270 & ~n29532;
  assign n30946 = ~i_RtoB_ACK0 & ~n30945;
  assign n30947 = ~n23107 & ~n30946;
  assign n30948 = ~controllable_DEQ & ~n30947;
  assign n30949 = ~n23105 & ~n30948;
  assign n30950 = i_FULL & ~n30949;
  assign n30951 = ~n11286 & ~n29502;
  assign n30952 = ~i_RtoB_ACK0 & ~n30951;
  assign n30953 = ~n23089 & ~n30952;
  assign n30954 = ~controllable_DEQ & ~n30953;
  assign n30955 = ~n23117 & ~n30954;
  assign n30956 = ~i_FULL & ~n30955;
  assign n30957 = ~n30950 & ~n30956;
  assign n30958 = ~i_nEMPTY & ~n30957;
  assign n30959 = ~n30944 & ~n30958;
  assign n30960 = controllable_BtoS_ACK0 & ~n30959;
  assign n30961 = ~n30445 & ~n30960;
  assign n30962 = n4465 & ~n30961;
  assign n30963 = ~n30447 & ~n30962;
  assign n30964 = ~i_StoB_REQ10 & ~n30963;
  assign n30965 = ~n30926 & ~n30964;
  assign n30966 = ~controllable_BtoS_ACK10 & ~n30965;
  assign n30967 = ~n30806 & ~n30966;
  assign n30968 = n4464 & ~n30967;
  assign n30969 = ~n30774 & ~n30806;
  assign n30970 = ~n4464 & ~n30969;
  assign n30971 = ~n30968 & ~n30970;
  assign n30972 = ~n4463 & ~n30971;
  assign n30973 = ~n30891 & ~n30972;
  assign n30974 = ~n4462 & ~n30973;
  assign n30975 = ~n30780 & ~n30974;
  assign n30976 = n4461 & ~n30975;
  assign n30977 = ~n14749 & ~n27816;
  assign n30978 = ~i_RtoB_ACK0 & ~n30977;
  assign n30979 = ~n20977 & ~n30978;
  assign n30980 = controllable_DEQ & ~n30979;
  assign n30981 = ~n14765 & ~n25928;
  assign n30982 = ~i_RtoB_ACK0 & ~n30981;
  assign n30983 = ~n20983 & ~n30982;
  assign n30984 = ~controllable_DEQ & ~n30983;
  assign n30985 = ~n30980 & ~n30984;
  assign n30986 = i_FULL & ~n30985;
  assign n30987 = ~n14765 & ~n27827;
  assign n30988 = ~i_RtoB_ACK0 & ~n30987;
  assign n30989 = ~n20983 & ~n30988;
  assign n30990 = ~controllable_DEQ & ~n30989;
  assign n30991 = ~n20981 & ~n30990;
  assign n30992 = ~i_FULL & ~n30991;
  assign n30993 = ~n30986 & ~n30992;
  assign n30994 = i_nEMPTY & ~n30993;
  assign n30995 = ~n14784 & ~n25951;
  assign n30996 = ~i_RtoB_ACK0 & ~n30995;
  assign n30997 = ~n20977 & ~n30996;
  assign n30998 = ~controllable_DEQ & ~n30997;
  assign n30999 = ~n20993 & ~n30998;
  assign n31000 = i_FULL & ~n30999;
  assign n31001 = ~n14749 & ~n27842;
  assign n31002 = ~i_RtoB_ACK0 & ~n31001;
  assign n31003 = ~n20977 & ~n31002;
  assign n31004 = ~controllable_DEQ & ~n31003;
  assign n31005 = ~n21003 & ~n31004;
  assign n31006 = ~i_FULL & ~n31005;
  assign n31007 = ~n31000 & ~n31006;
  assign n31008 = ~i_nEMPTY & ~n31007;
  assign n31009 = ~n30994 & ~n31008;
  assign n31010 = controllable_BtoS_ACK0 & ~n31009;
  assign n31011 = ~n27862 & ~n28753;
  assign n31012 = ~i_RtoB_ACK0 & ~n31011;
  assign n31013 = ~n29625 & ~n31012;
  assign n31014 = controllable_DEQ & ~n31013;
  assign n31015 = ~n25976 & ~n29437;
  assign n31016 = ~i_RtoB_ACK0 & ~n31015;
  assign n31017 = ~n29631 & ~n31016;
  assign n31018 = ~controllable_DEQ & ~n31017;
  assign n31019 = ~n31014 & ~n31018;
  assign n31020 = i_FULL & ~n31019;
  assign n31021 = ~n27885 & ~n29437;
  assign n31022 = ~i_RtoB_ACK0 & ~n31021;
  assign n31023 = ~n29631 & ~n31022;
  assign n31024 = ~controllable_DEQ & ~n31023;
  assign n31025 = ~n29641 & ~n31024;
  assign n31026 = ~i_FULL & ~n31025;
  assign n31027 = ~n31020 & ~n31026;
  assign n31028 = i_nEMPTY & ~n31027;
  assign n31029 = ~n25999 & ~n29447;
  assign n31030 = ~i_RtoB_ACK0 & ~n31029;
  assign n31031 = ~n29625 & ~n31030;
  assign n31032 = ~controllable_DEQ & ~n31031;
  assign n31033 = ~n29653 & ~n31032;
  assign n31034 = i_FULL & ~n31033;
  assign n31035 = ~n27913 & ~n28753;
  assign n31036 = ~i_RtoB_ACK0 & ~n31035;
  assign n31037 = ~n29625 & ~n31036;
  assign n31038 = ~controllable_DEQ & ~n31037;
  assign n31039 = ~n29663 & ~n31038;
  assign n31040 = ~i_FULL & ~n31039;
  assign n31041 = ~n31034 & ~n31040;
  assign n31042 = ~i_nEMPTY & ~n31041;
  assign n31043 = ~n31028 & ~n31042;
  assign n31044 = ~controllable_BtoS_ACK0 & ~n31043;
  assign n31045 = ~n31010 & ~n31044;
  assign n31046 = n4465 & ~n31045;
  assign n31047 = ~n27928 & ~n28753;
  assign n31048 = ~i_RtoB_ACK0 & ~n31047;
  assign n31049 = ~n29625 & ~n31048;
  assign n31050 = controllable_DEQ & ~n31049;
  assign n31051 = ~n26026 & ~n29437;
  assign n31052 = ~i_RtoB_ACK0 & ~n31051;
  assign n31053 = ~n29631 & ~n31052;
  assign n31054 = ~controllable_DEQ & ~n31053;
  assign n31055 = ~n31050 & ~n31054;
  assign n31056 = i_FULL & ~n31055;
  assign n31057 = ~n27939 & ~n29437;
  assign n31058 = ~i_RtoB_ACK0 & ~n31057;
  assign n31059 = ~n29631 & ~n31058;
  assign n31060 = ~controllable_DEQ & ~n31059;
  assign n31061 = ~n29641 & ~n31060;
  assign n31062 = ~i_FULL & ~n31061;
  assign n31063 = ~n31056 & ~n31062;
  assign n31064 = i_nEMPTY & ~n31063;
  assign n31065 = ~n26049 & ~n29447;
  assign n31066 = ~i_RtoB_ACK0 & ~n31065;
  assign n31067 = ~n29625 & ~n31066;
  assign n31068 = ~controllable_DEQ & ~n31067;
  assign n31069 = ~n29653 & ~n31068;
  assign n31070 = i_FULL & ~n31069;
  assign n31071 = ~n27954 & ~n28753;
  assign n31072 = ~i_RtoB_ACK0 & ~n31071;
  assign n31073 = ~n29625 & ~n31072;
  assign n31074 = ~controllable_DEQ & ~n31073;
  assign n31075 = ~n29663 & ~n31074;
  assign n31076 = ~i_FULL & ~n31075;
  assign n31077 = ~n31070 & ~n31076;
  assign n31078 = ~i_nEMPTY & ~n31077;
  assign n31079 = ~n31064 & ~n31078;
  assign n31080 = ~controllable_BtoS_ACK0 & ~n31079;
  assign n31081 = ~n21013 & ~n31080;
  assign n31082 = ~n4465 & ~n31081;
  assign n31083 = ~n31046 & ~n31082;
  assign n31084 = i_StoB_REQ10 & ~n31083;
  assign n31085 = ~n17620 & ~n27972;
  assign n31086 = ~i_RtoB_ACK0 & ~n31085;
  assign n31087 = ~n23089 & ~n31086;
  assign n31088 = controllable_DEQ & ~n31087;
  assign n31089 = ~n17635 & ~n27977;
  assign n31090 = ~i_RtoB_ACK0 & ~n31089;
  assign n31091 = ~n23095 & ~n31090;
  assign n31092 = ~controllable_DEQ & ~n31091;
  assign n31093 = ~n31088 & ~n31092;
  assign n31094 = i_FULL & ~n31093;
  assign n31095 = ~n17635 & ~n27984;
  assign n31096 = ~i_RtoB_ACK0 & ~n31095;
  assign n31097 = ~n23095 & ~n31096;
  assign n31098 = ~controllable_DEQ & ~n31097;
  assign n31099 = ~n23093 & ~n31098;
  assign n31100 = ~i_FULL & ~n31099;
  assign n31101 = ~n31094 & ~n31100;
  assign n31102 = i_nEMPTY & ~n31101;
  assign n31103 = ~n17657 & ~n27993;
  assign n31104 = ~i_RtoB_ACK0 & ~n31103;
  assign n31105 = ~n23107 & ~n31104;
  assign n31106 = ~controllable_DEQ & ~n31105;
  assign n31107 = ~n23105 & ~n31106;
  assign n31108 = i_FULL & ~n31107;
  assign n31109 = ~n17620 & ~n28003;
  assign n31110 = ~i_RtoB_ACK0 & ~n31109;
  assign n31111 = ~n23089 & ~n31110;
  assign n31112 = ~controllable_DEQ & ~n31111;
  assign n31113 = ~n23117 & ~n31112;
  assign n31114 = ~i_FULL & ~n31113;
  assign n31115 = ~n31108 & ~n31114;
  assign n31116 = ~i_nEMPTY & ~n31115;
  assign n31117 = ~n31102 & ~n31116;
  assign n31118 = controllable_BtoS_ACK0 & ~n31117;
  assign n31119 = ~n17699 & ~n28017;
  assign n31120 = ~i_RtoB_ACK0 & ~n31119;
  assign n31121 = ~n23129 & ~n31120;
  assign n31122 = controllable_DEQ & ~n31121;
  assign n31123 = ~n17718 & ~n28022;
  assign n31124 = ~i_RtoB_ACK0 & ~n31123;
  assign n31125 = ~n23135 & ~n31124;
  assign n31126 = ~controllable_DEQ & ~n31125;
  assign n31127 = ~n31122 & ~n31126;
  assign n31128 = i_FULL & ~n31127;
  assign n31129 = ~n17718 & ~n28029;
  assign n31130 = ~i_RtoB_ACK0 & ~n31129;
  assign n31131 = ~n23135 & ~n31130;
  assign n31132 = ~controllable_DEQ & ~n31131;
  assign n31133 = ~n23133 & ~n31132;
  assign n31134 = ~i_FULL & ~n31133;
  assign n31135 = ~n31128 & ~n31134;
  assign n31136 = i_nEMPTY & ~n31135;
  assign n31137 = ~n17751 & ~n28038;
  assign n31138 = ~i_RtoB_ACK0 & ~n31137;
  assign n31139 = ~n23147 & ~n31138;
  assign n31140 = ~controllable_DEQ & ~n31139;
  assign n31141 = ~n23145 & ~n31140;
  assign n31142 = i_FULL & ~n31141;
  assign n31143 = ~n17699 & ~n28048;
  assign n31144 = ~i_RtoB_ACK0 & ~n31143;
  assign n31145 = ~n23129 & ~n31144;
  assign n31146 = ~controllable_DEQ & ~n31145;
  assign n31147 = ~n23157 & ~n31146;
  assign n31148 = ~i_FULL & ~n31147;
  assign n31149 = ~n31142 & ~n31148;
  assign n31150 = ~i_nEMPTY & ~n31149;
  assign n31151 = ~n31136 & ~n31150;
  assign n31152 = ~controllable_BtoS_ACK0 & ~n31151;
  assign n31153 = ~n31118 & ~n31152;
  assign n31154 = n4465 & ~n31153;
  assign n31155 = ~n17699 & ~n28064;
  assign n31156 = ~i_RtoB_ACK0 & ~n31155;
  assign n31157 = ~n23129 & ~n31156;
  assign n31158 = controllable_DEQ & ~n31157;
  assign n31159 = ~n17718 & ~n28069;
  assign n31160 = ~i_RtoB_ACK0 & ~n31159;
  assign n31161 = ~n23135 & ~n31160;
  assign n31162 = ~controllable_DEQ & ~n31161;
  assign n31163 = ~n31158 & ~n31162;
  assign n31164 = i_FULL & ~n31163;
  assign n31165 = ~n17718 & ~n28076;
  assign n31166 = ~i_RtoB_ACK0 & ~n31165;
  assign n31167 = ~n23135 & ~n31166;
  assign n31168 = ~controllable_DEQ & ~n31167;
  assign n31169 = ~n23133 & ~n31168;
  assign n31170 = ~i_FULL & ~n31169;
  assign n31171 = ~n31164 & ~n31170;
  assign n31172 = i_nEMPTY & ~n31171;
  assign n31173 = ~n17751 & ~n28085;
  assign n31174 = ~i_RtoB_ACK0 & ~n31173;
  assign n31175 = ~n23147 & ~n31174;
  assign n31176 = ~controllable_DEQ & ~n31175;
  assign n31177 = ~n23145 & ~n31176;
  assign n31178 = i_FULL & ~n31177;
  assign n31179 = ~n17699 & ~n28093;
  assign n31180 = ~i_RtoB_ACK0 & ~n31179;
  assign n31181 = ~n23129 & ~n31180;
  assign n31182 = ~controllable_DEQ & ~n31181;
  assign n31183 = ~n23157 & ~n31182;
  assign n31184 = ~i_FULL & ~n31183;
  assign n31185 = ~n31178 & ~n31184;
  assign n31186 = ~i_nEMPTY & ~n31185;
  assign n31187 = ~n31172 & ~n31186;
  assign n31188 = ~controllable_BtoS_ACK0 & ~n31187;
  assign n31189 = ~n23127 & ~n31188;
  assign n31190 = ~n4465 & ~n31189;
  assign n31191 = ~n31154 & ~n31190;
  assign n31192 = ~i_StoB_REQ10 & ~n31191;
  assign n31193 = ~n31084 & ~n31192;
  assign n31194 = controllable_BtoS_ACK10 & ~n31193;
  assign n31195 = ~n28118 & ~n29840;
  assign n31196 = ~i_RtoB_ACK0 & ~n31195;
  assign n31197 = ~n29825 & ~n31196;
  assign n31198 = controllable_DEQ & ~n31197;
  assign n31199 = ~n27977 & ~n29938;
  assign n31200 = ~i_RtoB_ACK0 & ~n31199;
  assign n31201 = ~n29832 & ~n31200;
  assign n31202 = ~controllable_DEQ & ~n31201;
  assign n31203 = ~n31198 & ~n31202;
  assign n31204 = i_FULL & ~n31203;
  assign n31205 = ~n27984 & ~n29938;
  assign n31206 = ~i_RtoB_ACK0 & ~n31205;
  assign n31207 = ~n29832 & ~n31206;
  assign n31208 = ~controllable_DEQ & ~n31207;
  assign n31209 = ~n29844 & ~n31208;
  assign n31210 = ~i_FULL & ~n31209;
  assign n31211 = ~n31204 & ~n31210;
  assign n31212 = i_nEMPTY & ~n31211;
  assign n31213 = ~n27993 & ~n29945;
  assign n31214 = ~i_RtoB_ACK0 & ~n31213;
  assign n31215 = ~n29860 & ~n31214;
  assign n31216 = ~controllable_DEQ & ~n31215;
  assign n31217 = ~n29858 & ~n31216;
  assign n31218 = i_FULL & ~n31217;
  assign n31219 = ~controllable_DEQ & ~n31197;
  assign n31220 = ~n29872 & ~n31219;
  assign n31221 = ~i_FULL & ~n31220;
  assign n31222 = ~n31218 & ~n31221;
  assign n31223 = ~i_nEMPTY & ~n31222;
  assign n31224 = ~n31212 & ~n31223;
  assign n31225 = controllable_BtoS_ACK0 & ~n31224;
  assign n31226 = ~n28179 & ~n29896;
  assign n31227 = ~i_RtoB_ACK0 & ~n31226;
  assign n31228 = ~n29881 & ~n31227;
  assign n31229 = controllable_DEQ & ~n31228;
  assign n31230 = controllable_BtoR_REQ0 & ~n17710;
  assign n31231 = ~n28022 & ~n31230;
  assign n31232 = ~i_RtoB_ACK0 & ~n31231;
  assign n31233 = ~n29888 & ~n31232;
  assign n31234 = ~controllable_DEQ & ~n31233;
  assign n31235 = ~n31229 & ~n31234;
  assign n31236 = i_FULL & ~n31235;
  assign n31237 = ~n28029 & ~n31230;
  assign n31238 = ~i_RtoB_ACK0 & ~n31237;
  assign n31239 = ~n29888 & ~n31238;
  assign n31240 = ~controllable_DEQ & ~n31239;
  assign n31241 = ~n29900 & ~n31240;
  assign n31242 = ~i_FULL & ~n31241;
  assign n31243 = ~n31236 & ~n31242;
  assign n31244 = i_nEMPTY & ~n31243;
  assign n31245 = controllable_BtoR_REQ0 & ~n17691;
  assign n31246 = ~n28038 & ~n31245;
  assign n31247 = ~i_RtoB_ACK0 & ~n31246;
  assign n31248 = ~n29916 & ~n31247;
  assign n31249 = ~controllable_DEQ & ~n31248;
  assign n31250 = ~n29914 & ~n31249;
  assign n31251 = i_FULL & ~n31250;
  assign n31252 = ~controllable_DEQ & ~n31228;
  assign n31253 = ~n29928 & ~n31252;
  assign n31254 = ~i_FULL & ~n31253;
  assign n31255 = ~n31251 & ~n31254;
  assign n31256 = ~i_nEMPTY & ~n31255;
  assign n31257 = ~n31244 & ~n31256;
  assign n31258 = ~controllable_BtoS_ACK0 & ~n31257;
  assign n31259 = ~n31225 & ~n31258;
  assign n31260 = n4465 & ~n31259;
  assign n31261 = ~n28252 & ~n29896;
  assign n31262 = ~i_RtoB_ACK0 & ~n31261;
  assign n31263 = ~n29881 & ~n31262;
  assign n31264 = controllable_DEQ & ~n31263;
  assign n31265 = ~n28069 & ~n31230;
  assign n31266 = ~i_RtoB_ACK0 & ~n31265;
  assign n31267 = ~n29888 & ~n31266;
  assign n31268 = ~controllable_DEQ & ~n31267;
  assign n31269 = ~n31264 & ~n31268;
  assign n31270 = i_FULL & ~n31269;
  assign n31271 = ~n28076 & ~n31230;
  assign n31272 = ~i_RtoB_ACK0 & ~n31271;
  assign n31273 = ~n29888 & ~n31272;
  assign n31274 = ~controllable_DEQ & ~n31273;
  assign n31275 = ~n29900 & ~n31274;
  assign n31276 = ~i_FULL & ~n31275;
  assign n31277 = ~n31270 & ~n31276;
  assign n31278 = i_nEMPTY & ~n31277;
  assign n31279 = ~n28085 & ~n31245;
  assign n31280 = ~i_RtoB_ACK0 & ~n31279;
  assign n31281 = ~n29916 & ~n31280;
  assign n31282 = ~controllable_DEQ & ~n31281;
  assign n31283 = ~n29914 & ~n31282;
  assign n31284 = i_FULL & ~n31283;
  assign n31285 = ~controllable_DEQ & ~n31263;
  assign n31286 = ~n29928 & ~n31285;
  assign n31287 = ~i_FULL & ~n31286;
  assign n31288 = ~n31284 & ~n31287;
  assign n31289 = ~i_nEMPTY & ~n31288;
  assign n31290 = ~n31278 & ~n31289;
  assign n31291 = ~controllable_BtoS_ACK0 & ~n31290;
  assign n31292 = ~n29958 & ~n31291;
  assign n31293 = ~n4465 & ~n31292;
  assign n31294 = ~n31260 & ~n31293;
  assign n31295 = i_StoB_REQ10 & ~n31294;
  assign n31296 = ~n31192 & ~n31295;
  assign n31297 = ~controllable_BtoS_ACK10 & ~n31296;
  assign n31298 = ~n31194 & ~n31297;
  assign n31299 = n4464 & ~n31298;
  assign n31300 = ~n14749 & ~n28288;
  assign n31301 = ~i_RtoB_ACK0 & ~n31300;
  assign n31302 = ~n20977 & ~n31301;
  assign n31303 = controllable_DEQ & ~n31302;
  assign n31304 = ~n14765 & ~n26438;
  assign n31305 = ~i_RtoB_ACK0 & ~n31304;
  assign n31306 = ~n20983 & ~n31305;
  assign n31307 = ~controllable_DEQ & ~n31306;
  assign n31308 = ~n31303 & ~n31307;
  assign n31309 = i_FULL & ~n31308;
  assign n31310 = ~n14765 & ~n28299;
  assign n31311 = ~i_RtoB_ACK0 & ~n31310;
  assign n31312 = ~n20983 & ~n31311;
  assign n31313 = ~controllable_DEQ & ~n31312;
  assign n31314 = ~n20981 & ~n31313;
  assign n31315 = ~i_FULL & ~n31314;
  assign n31316 = ~n31309 & ~n31315;
  assign n31317 = i_nEMPTY & ~n31316;
  assign n31318 = ~n14784 & ~n26461;
  assign n31319 = ~i_RtoB_ACK0 & ~n31318;
  assign n31320 = ~n20977 & ~n31319;
  assign n31321 = ~controllable_DEQ & ~n31320;
  assign n31322 = ~n20993 & ~n31321;
  assign n31323 = i_FULL & ~n31322;
  assign n31324 = ~n14749 & ~n28314;
  assign n31325 = ~i_RtoB_ACK0 & ~n31324;
  assign n31326 = ~n20977 & ~n31325;
  assign n31327 = ~controllable_DEQ & ~n31326;
  assign n31328 = ~n21003 & ~n31327;
  assign n31329 = ~i_FULL & ~n31328;
  assign n31330 = ~n31323 & ~n31329;
  assign n31331 = ~i_nEMPTY & ~n31330;
  assign n31332 = ~n31317 & ~n31331;
  assign n31333 = controllable_BtoS_ACK0 & ~n31332;
  assign n31334 = ~n28327 & ~n28753;
  assign n31335 = ~i_RtoB_ACK0 & ~n31334;
  assign n31336 = ~n29625 & ~n31335;
  assign n31337 = controllable_DEQ & ~n31336;
  assign n31338 = ~n26486 & ~n29437;
  assign n31339 = ~i_RtoB_ACK0 & ~n31338;
  assign n31340 = ~n29631 & ~n31339;
  assign n31341 = ~controllable_DEQ & ~n31340;
  assign n31342 = ~n31337 & ~n31341;
  assign n31343 = i_FULL & ~n31342;
  assign n31344 = ~n28338 & ~n29437;
  assign n31345 = ~i_RtoB_ACK0 & ~n31344;
  assign n31346 = ~n29631 & ~n31345;
  assign n31347 = ~controllable_DEQ & ~n31346;
  assign n31348 = ~n29641 & ~n31347;
  assign n31349 = ~i_FULL & ~n31348;
  assign n31350 = ~n31343 & ~n31349;
  assign n31351 = i_nEMPTY & ~n31350;
  assign n31352 = ~n26509 & ~n29447;
  assign n31353 = ~i_RtoB_ACK0 & ~n31352;
  assign n31354 = ~n29625 & ~n31353;
  assign n31355 = ~controllable_DEQ & ~n31354;
  assign n31356 = ~n29653 & ~n31355;
  assign n31357 = i_FULL & ~n31356;
  assign n31358 = ~n28353 & ~n28753;
  assign n31359 = ~i_RtoB_ACK0 & ~n31358;
  assign n31360 = ~n29625 & ~n31359;
  assign n31361 = ~controllable_DEQ & ~n31360;
  assign n31362 = ~n29663 & ~n31361;
  assign n31363 = ~i_FULL & ~n31362;
  assign n31364 = ~n31357 & ~n31363;
  assign n31365 = ~i_nEMPTY & ~n31364;
  assign n31366 = ~n31351 & ~n31365;
  assign n31367 = ~controllable_BtoS_ACK0 & ~n31366;
  assign n31368 = ~n31333 & ~n31367;
  assign n31369 = n4465 & ~n31368;
  assign n31370 = ~n21013 & ~n31367;
  assign n31371 = ~n4465 & ~n31370;
  assign n31372 = ~n31369 & ~n31371;
  assign n31373 = i_StoB_REQ10 & ~n31372;
  assign n31374 = ~n17620 & ~n28373;
  assign n31375 = ~i_RtoB_ACK0 & ~n31374;
  assign n31376 = ~n23089 & ~n31375;
  assign n31377 = controllable_DEQ & ~n31376;
  assign n31378 = ~n17635 & ~n28378;
  assign n31379 = ~i_RtoB_ACK0 & ~n31378;
  assign n31380 = ~n23095 & ~n31379;
  assign n31381 = ~controllable_DEQ & ~n31380;
  assign n31382 = ~n31377 & ~n31381;
  assign n31383 = i_FULL & ~n31382;
  assign n31384 = ~n17635 & ~n28385;
  assign n31385 = ~i_RtoB_ACK0 & ~n31384;
  assign n31386 = ~n23095 & ~n31385;
  assign n31387 = ~controllable_DEQ & ~n31386;
  assign n31388 = ~n23093 & ~n31387;
  assign n31389 = ~i_FULL & ~n31388;
  assign n31390 = ~n31383 & ~n31389;
  assign n31391 = i_nEMPTY & ~n31390;
  assign n31392 = ~n17657 & ~n28394;
  assign n31393 = ~i_RtoB_ACK0 & ~n31392;
  assign n31394 = ~n23107 & ~n31393;
  assign n31395 = ~controllable_DEQ & ~n31394;
  assign n31396 = ~n23105 & ~n31395;
  assign n31397 = i_FULL & ~n31396;
  assign n31398 = ~n17620 & ~n28402;
  assign n31399 = ~i_RtoB_ACK0 & ~n31398;
  assign n31400 = ~n23089 & ~n31399;
  assign n31401 = ~controllable_DEQ & ~n31400;
  assign n31402 = ~n23117 & ~n31401;
  assign n31403 = ~i_FULL & ~n31402;
  assign n31404 = ~n31397 & ~n31403;
  assign n31405 = ~i_nEMPTY & ~n31404;
  assign n31406 = ~n31391 & ~n31405;
  assign n31407 = controllable_BtoS_ACK0 & ~n31406;
  assign n31408 = ~n17699 & ~n28416;
  assign n31409 = ~i_RtoB_ACK0 & ~n31408;
  assign n31410 = ~n23129 & ~n31409;
  assign n31411 = controllable_DEQ & ~n31410;
  assign n31412 = ~n17718 & ~n28421;
  assign n31413 = ~i_RtoB_ACK0 & ~n31412;
  assign n31414 = ~n23135 & ~n31413;
  assign n31415 = ~controllable_DEQ & ~n31414;
  assign n31416 = ~n31411 & ~n31415;
  assign n31417 = i_FULL & ~n31416;
  assign n31418 = ~n17718 & ~n28428;
  assign n31419 = ~i_RtoB_ACK0 & ~n31418;
  assign n31420 = ~n23135 & ~n31419;
  assign n31421 = ~controllable_DEQ & ~n31420;
  assign n31422 = ~n23133 & ~n31421;
  assign n31423 = ~i_FULL & ~n31422;
  assign n31424 = ~n31417 & ~n31423;
  assign n31425 = i_nEMPTY & ~n31424;
  assign n31426 = ~n17751 & ~n28437;
  assign n31427 = ~i_RtoB_ACK0 & ~n31426;
  assign n31428 = ~n23147 & ~n31427;
  assign n31429 = ~controllable_DEQ & ~n31428;
  assign n31430 = ~n23145 & ~n31429;
  assign n31431 = i_FULL & ~n31430;
  assign n31432 = ~n17699 & ~n28445;
  assign n31433 = ~i_RtoB_ACK0 & ~n31432;
  assign n31434 = ~n23129 & ~n31433;
  assign n31435 = ~controllable_DEQ & ~n31434;
  assign n31436 = ~n23157 & ~n31435;
  assign n31437 = ~i_FULL & ~n31436;
  assign n31438 = ~n31431 & ~n31437;
  assign n31439 = ~i_nEMPTY & ~n31438;
  assign n31440 = ~n31425 & ~n31439;
  assign n31441 = ~controllable_BtoS_ACK0 & ~n31440;
  assign n31442 = ~n31407 & ~n31441;
  assign n31443 = n4465 & ~n31442;
  assign n31444 = ~n23127 & ~n31441;
  assign n31445 = ~n4465 & ~n31444;
  assign n31446 = ~n31443 & ~n31445;
  assign n31447 = ~i_StoB_REQ10 & ~n31446;
  assign n31448 = ~n31373 & ~n31447;
  assign n31449 = controllable_BtoS_ACK10 & ~n31448;
  assign n31450 = ~n28467 & ~n29840;
  assign n31451 = ~i_RtoB_ACK0 & ~n31450;
  assign n31452 = ~n29825 & ~n31451;
  assign n31453 = controllable_DEQ & ~n31452;
  assign n31454 = ~n28378 & ~n29938;
  assign n31455 = ~i_RtoB_ACK0 & ~n31454;
  assign n31456 = ~n29832 & ~n31455;
  assign n31457 = ~controllable_DEQ & ~n31456;
  assign n31458 = ~n31453 & ~n31457;
  assign n31459 = i_FULL & ~n31458;
  assign n31460 = ~n28385 & ~n29938;
  assign n31461 = ~i_RtoB_ACK0 & ~n31460;
  assign n31462 = ~n29832 & ~n31461;
  assign n31463 = ~controllable_DEQ & ~n31462;
  assign n31464 = ~n29844 & ~n31463;
  assign n31465 = ~i_FULL & ~n31464;
  assign n31466 = ~n31459 & ~n31465;
  assign n31467 = i_nEMPTY & ~n31466;
  assign n31468 = ~n28394 & ~n29945;
  assign n31469 = ~i_RtoB_ACK0 & ~n31468;
  assign n31470 = ~n29860 & ~n31469;
  assign n31471 = ~controllable_DEQ & ~n31470;
  assign n31472 = ~n29858 & ~n31471;
  assign n31473 = i_FULL & ~n31472;
  assign n31474 = ~controllable_DEQ & ~n31452;
  assign n31475 = ~n29872 & ~n31474;
  assign n31476 = ~i_FULL & ~n31475;
  assign n31477 = ~n31473 & ~n31476;
  assign n31478 = ~i_nEMPTY & ~n31477;
  assign n31479 = ~n31467 & ~n31478;
  assign n31480 = controllable_BtoS_ACK0 & ~n31479;
  assign n31481 = ~n28496 & ~n29896;
  assign n31482 = ~i_RtoB_ACK0 & ~n31481;
  assign n31483 = ~n29881 & ~n31482;
  assign n31484 = controllable_DEQ & ~n31483;
  assign n31485 = ~n28421 & ~n31230;
  assign n31486 = ~i_RtoB_ACK0 & ~n31485;
  assign n31487 = ~n29888 & ~n31486;
  assign n31488 = ~controllable_DEQ & ~n31487;
  assign n31489 = ~n31484 & ~n31488;
  assign n31490 = i_FULL & ~n31489;
  assign n31491 = ~n28428 & ~n31230;
  assign n31492 = ~i_RtoB_ACK0 & ~n31491;
  assign n31493 = ~n29888 & ~n31492;
  assign n31494 = ~controllable_DEQ & ~n31493;
  assign n31495 = ~n29900 & ~n31494;
  assign n31496 = ~i_FULL & ~n31495;
  assign n31497 = ~n31490 & ~n31496;
  assign n31498 = i_nEMPTY & ~n31497;
  assign n31499 = ~n28437 & ~n31245;
  assign n31500 = ~i_RtoB_ACK0 & ~n31499;
  assign n31501 = ~n29916 & ~n31500;
  assign n31502 = ~controllable_DEQ & ~n31501;
  assign n31503 = ~n29914 & ~n31502;
  assign n31504 = i_FULL & ~n31503;
  assign n31505 = ~controllable_DEQ & ~n31483;
  assign n31506 = ~n29928 & ~n31505;
  assign n31507 = ~i_FULL & ~n31506;
  assign n31508 = ~n31504 & ~n31507;
  assign n31509 = ~i_nEMPTY & ~n31508;
  assign n31510 = ~n31498 & ~n31509;
  assign n31511 = ~controllable_BtoS_ACK0 & ~n31510;
  assign n31512 = ~n31480 & ~n31511;
  assign n31513 = n4465 & ~n31512;
  assign n31514 = ~n29958 & ~n31511;
  assign n31515 = ~n4465 & ~n31514;
  assign n31516 = ~n31513 & ~n31515;
  assign n31517 = i_StoB_REQ10 & ~n31516;
  assign n31518 = ~n31447 & ~n31517;
  assign n31519 = ~controllable_BtoS_ACK10 & ~n31518;
  assign n31520 = ~n31449 & ~n31519;
  assign n31521 = ~n4464 & ~n31520;
  assign n31522 = ~n31299 & ~n31521;
  assign n31523 = n4463 & ~n31522;
  assign n31524 = ~n11333 & ~n31230;
  assign n31525 = ~i_RtoB_ACK0 & ~n31524;
  assign n31526 = ~n29888 & ~n31525;
  assign n31527 = ~controllable_DEQ & ~n31526;
  assign n31528 = ~n29900 & ~n31527;
  assign n31529 = i_nEMPTY & ~n31528;
  assign n31530 = ~n11352 & ~n31245;
  assign n31531 = ~i_RtoB_ACK0 & ~n31530;
  assign n31532 = ~n29916 & ~n31531;
  assign n31533 = ~controllable_DEQ & ~n31532;
  assign n31534 = ~n29914 & ~n31533;
  assign n31535 = i_FULL & ~n31534;
  assign n31536 = ~controllable_DEQ & ~n29899;
  assign n31537 = ~n29928 & ~n31536;
  assign n31538 = ~i_FULL & ~n31537;
  assign n31539 = ~n31535 & ~n31538;
  assign n31540 = ~i_nEMPTY & ~n31539;
  assign n31541 = ~n31529 & ~n31540;
  assign n31542 = ~controllable_BtoS_ACK0 & ~n31541;
  assign n31543 = ~n29958 & ~n31542;
  assign n31544 = i_StoB_REQ10 & ~n31543;
  assign n31545 = ~n23169 & ~n31544;
  assign n31546 = ~controllable_BtoS_ACK10 & ~n31545;
  assign n31547 = ~n30806 & ~n31546;
  assign n31548 = ~n4463 & ~n31547;
  assign n31549 = ~n31523 & ~n31548;
  assign n31550 = n4462 & ~n31549;
  assign n31551 = ~n28589 & ~n29840;
  assign n31552 = ~i_RtoB_ACK0 & ~n31551;
  assign n31553 = ~n29825 & ~n31552;
  assign n31554 = controllable_DEQ & ~n31553;
  assign n31555 = ~n28594 & ~n29938;
  assign n31556 = ~i_RtoB_ACK0 & ~n31555;
  assign n31557 = ~n29832 & ~n31556;
  assign n31558 = ~controllable_DEQ & ~n31557;
  assign n31559 = ~n31554 & ~n31558;
  assign n31560 = i_FULL & ~n31559;
  assign n31561 = ~n28601 & ~n29938;
  assign n31562 = ~i_RtoB_ACK0 & ~n31561;
  assign n31563 = ~n29832 & ~n31562;
  assign n31564 = ~controllable_DEQ & ~n31563;
  assign n31565 = ~n29844 & ~n31564;
  assign n31566 = ~i_FULL & ~n31565;
  assign n31567 = ~n31560 & ~n31566;
  assign n31568 = i_nEMPTY & ~n31567;
  assign n31569 = ~n28610 & ~n29945;
  assign n31570 = ~i_RtoB_ACK0 & ~n31569;
  assign n31571 = ~n29860 & ~n31570;
  assign n31572 = ~controllable_DEQ & ~n31571;
  assign n31573 = ~n29858 & ~n31572;
  assign n31574 = i_FULL & ~n31573;
  assign n31575 = ~controllable_DEQ & ~n31553;
  assign n31576 = ~n29872 & ~n31575;
  assign n31577 = ~i_FULL & ~n31576;
  assign n31578 = ~n31574 & ~n31577;
  assign n31579 = ~i_nEMPTY & ~n31578;
  assign n31580 = ~n31568 & ~n31579;
  assign n31581 = controllable_BtoS_ACK0 & ~n31580;
  assign n31582 = ~n31291 & ~n31581;
  assign n31583 = n4465 & ~n31582;
  assign n31584 = ~n31293 & ~n31583;
  assign n31585 = i_StoB_REQ10 & ~n31584;
  assign n31586 = ~n17620 & ~n28631;
  assign n31587 = ~i_RtoB_ACK0 & ~n31586;
  assign n31588 = ~n23089 & ~n31587;
  assign n31589 = controllable_DEQ & ~n31588;
  assign n31590 = ~n17635 & ~n28594;
  assign n31591 = ~i_RtoB_ACK0 & ~n31590;
  assign n31592 = ~n23095 & ~n31591;
  assign n31593 = ~controllable_DEQ & ~n31592;
  assign n31594 = ~n31589 & ~n31593;
  assign n31595 = i_FULL & ~n31594;
  assign n31596 = ~n17635 & ~n28601;
  assign n31597 = ~i_RtoB_ACK0 & ~n31596;
  assign n31598 = ~n23095 & ~n31597;
  assign n31599 = ~controllable_DEQ & ~n31598;
  assign n31600 = ~n23093 & ~n31599;
  assign n31601 = ~i_FULL & ~n31600;
  assign n31602 = ~n31595 & ~n31601;
  assign n31603 = i_nEMPTY & ~n31602;
  assign n31604 = ~n17657 & ~n28610;
  assign n31605 = ~i_RtoB_ACK0 & ~n31604;
  assign n31606 = ~n23107 & ~n31605;
  assign n31607 = ~controllable_DEQ & ~n31606;
  assign n31608 = ~n23105 & ~n31607;
  assign n31609 = i_FULL & ~n31608;
  assign n31610 = ~n17620 & ~n28651;
  assign n31611 = ~i_RtoB_ACK0 & ~n31610;
  assign n31612 = ~n23089 & ~n31611;
  assign n31613 = ~controllable_DEQ & ~n31612;
  assign n31614 = ~n23117 & ~n31613;
  assign n31615 = ~i_FULL & ~n31614;
  assign n31616 = ~n31609 & ~n31615;
  assign n31617 = ~i_nEMPTY & ~n31616;
  assign n31618 = ~n31603 & ~n31617;
  assign n31619 = controllable_BtoS_ACK0 & ~n31618;
  assign n31620 = ~n31188 & ~n31619;
  assign n31621 = n4465 & ~n31620;
  assign n31622 = ~n31190 & ~n31621;
  assign n31623 = ~i_StoB_REQ10 & ~n31622;
  assign n31624 = ~n31585 & ~n31623;
  assign n31625 = ~controllable_BtoS_ACK10 & ~n31624;
  assign n31626 = ~n30806 & ~n31625;
  assign n31627 = n4464 & ~n31626;
  assign n31628 = ~n30806 & ~n31519;
  assign n31629 = ~n4464 & ~n31628;
  assign n31630 = ~n31627 & ~n31629;
  assign n31631 = n4463 & ~n31630;
  assign n31632 = ~n31548 & ~n31631;
  assign n31633 = ~n4462 & ~n31632;
  assign n31634 = ~n31550 & ~n31633;
  assign n31635 = ~n4461 & ~n31634;
  assign n31636 = ~n30976 & ~n31635;
  assign n31637 = ~n4459 & ~n31636;
  assign n31638 = ~n5242 & ~n18867;
  assign n31639 = ~controllable_BtoR_REQ0 & ~n31638;
  assign n31640 = ~n28681 & ~n31639;
  assign n31641 = ~i_RtoB_ACK0 & ~n31640;
  assign n31642 = ~n20977 & ~n31641;
  assign n31643 = controllable_DEQ & ~n31642;
  assign n31644 = controllable_BtoR_REQ1 & ~n5229;
  assign n31645 = ~n18874 & ~n31644;
  assign n31646 = ~controllable_BtoR_REQ0 & ~n31645;
  assign n31647 = ~n28689 & ~n31646;
  assign n31648 = ~i_RtoB_ACK0 & ~n31647;
  assign n31649 = ~n20983 & ~n31648;
  assign n31650 = ~controllable_DEQ & ~n31649;
  assign n31651 = ~n31643 & ~n31650;
  assign n31652 = i_FULL & ~n31651;
  assign n31653 = ~n18888 & ~n31644;
  assign n31654 = ~controllable_BtoR_REQ0 & ~n31653;
  assign n31655 = ~n28699 & ~n31654;
  assign n31656 = ~i_RtoB_ACK0 & ~n31655;
  assign n31657 = ~n20983 & ~n31656;
  assign n31658 = ~controllable_DEQ & ~n31657;
  assign n31659 = ~n20981 & ~n31658;
  assign n31660 = ~i_FULL & ~n31659;
  assign n31661 = ~n31652 & ~n31660;
  assign n31662 = i_nEMPTY & ~n31661;
  assign n31663 = controllable_BtoR_REQ1 & ~n5231;
  assign n31664 = ~n18903 & ~n31663;
  assign n31665 = ~controllable_BtoR_REQ0 & ~n31664;
  assign n31666 = ~n28711 & ~n31665;
  assign n31667 = ~i_RtoB_ACK0 & ~n31666;
  assign n31668 = ~n20977 & ~n31667;
  assign n31669 = ~controllable_DEQ & ~n31668;
  assign n31670 = ~n20993 & ~n31669;
  assign n31671 = i_FULL & ~n31670;
  assign n31672 = ~n5242 & ~n18917;
  assign n31673 = ~controllable_BtoR_REQ0 & ~n31672;
  assign n31674 = ~n28681 & ~n31673;
  assign n31675 = ~i_RtoB_ACK0 & ~n31674;
  assign n31676 = ~n20977 & ~n31675;
  assign n31677 = ~controllable_DEQ & ~n31676;
  assign n31678 = ~n21003 & ~n31677;
  assign n31679 = ~i_FULL & ~n31678;
  assign n31680 = ~n31671 & ~n31679;
  assign n31681 = ~i_nEMPTY & ~n31680;
  assign n31682 = ~n31662 & ~n31681;
  assign n31683 = controllable_BtoS_ACK0 & ~n31682;
  assign n31684 = ~n18931 & ~n27878;
  assign n31685 = ~controllable_BtoR_REQ0 & ~n31684;
  assign n31686 = ~n28733 & ~n31685;
  assign n31687 = ~i_RtoB_ACK0 & ~n31686;
  assign n31688 = ~n29625 & ~n31687;
  assign n31689 = controllable_DEQ & ~n31688;
  assign n31690 = controllable_BtoR_REQ1 & ~n8851;
  assign n31691 = ~n18938 & ~n31690;
  assign n31692 = ~controllable_BtoR_REQ0 & ~n31691;
  assign n31693 = ~n28743 & ~n31692;
  assign n31694 = ~i_RtoB_ACK0 & ~n31693;
  assign n31695 = ~n29631 & ~n31694;
  assign n31696 = ~controllable_DEQ & ~n31695;
  assign n31697 = ~n31689 & ~n31696;
  assign n31698 = i_FULL & ~n31697;
  assign n31699 = ~n18956 & ~n31690;
  assign n31700 = ~controllable_BtoR_REQ0 & ~n31699;
  assign n31701 = ~n28761 & ~n31700;
  assign n31702 = ~i_RtoB_ACK0 & ~n31701;
  assign n31703 = ~n29631 & ~n31702;
  assign n31704 = ~controllable_DEQ & ~n31703;
  assign n31705 = ~n29641 & ~n31704;
  assign n31706 = ~i_FULL & ~n31705;
  assign n31707 = ~n31698 & ~n31706;
  assign n31708 = i_nEMPTY & ~n31707;
  assign n31709 = controllable_BtoR_REQ1 & ~n8853;
  assign n31710 = ~n18972 & ~n31709;
  assign n31711 = ~controllable_BtoR_REQ0 & ~n31710;
  assign n31712 = ~n28777 & ~n31711;
  assign n31713 = ~i_RtoB_ACK0 & ~n31712;
  assign n31714 = ~n29625 & ~n31713;
  assign n31715 = ~controllable_DEQ & ~n31714;
  assign n31716 = ~n29653 & ~n31715;
  assign n31717 = i_FULL & ~n31716;
  assign n31718 = ~n18987 & ~n27878;
  assign n31719 = ~controllable_BtoR_REQ0 & ~n31718;
  assign n31720 = ~n28733 & ~n31719;
  assign n31721 = ~i_RtoB_ACK0 & ~n31720;
  assign n31722 = ~n29625 & ~n31721;
  assign n31723 = ~controllable_DEQ & ~n31722;
  assign n31724 = ~n29663 & ~n31723;
  assign n31725 = ~i_FULL & ~n31724;
  assign n31726 = ~n31717 & ~n31725;
  assign n31727 = ~i_nEMPTY & ~n31726;
  assign n31728 = ~n31708 & ~n31727;
  assign n31729 = ~controllable_BtoS_ACK0 & ~n31728;
  assign n31730 = ~n31683 & ~n31729;
  assign n31731 = n4465 & ~n31730;
  assign n31732 = ~n19003 & ~n27878;
  assign n31733 = ~controllable_BtoR_REQ0 & ~n31732;
  assign n31734 = ~n28803 & ~n31733;
  assign n31735 = ~i_RtoB_ACK0 & ~n31734;
  assign n31736 = ~n29625 & ~n31735;
  assign n31737 = controllable_DEQ & ~n31736;
  assign n31738 = ~n19010 & ~n31690;
  assign n31739 = ~controllable_BtoR_REQ0 & ~n31738;
  assign n31740 = ~n28811 & ~n31739;
  assign n31741 = ~i_RtoB_ACK0 & ~n31740;
  assign n31742 = ~n29631 & ~n31741;
  assign n31743 = ~controllable_DEQ & ~n31742;
  assign n31744 = ~n31737 & ~n31743;
  assign n31745 = i_FULL & ~n31744;
  assign n31746 = ~n19024 & ~n31690;
  assign n31747 = ~controllable_BtoR_REQ0 & ~n31746;
  assign n31748 = ~n28821 & ~n31747;
  assign n31749 = ~i_RtoB_ACK0 & ~n31748;
  assign n31750 = ~n29631 & ~n31749;
  assign n31751 = ~controllable_DEQ & ~n31750;
  assign n31752 = ~n29641 & ~n31751;
  assign n31753 = ~i_FULL & ~n31752;
  assign n31754 = ~n31745 & ~n31753;
  assign n31755 = i_nEMPTY & ~n31754;
  assign n31756 = ~n19039 & ~n31709;
  assign n31757 = ~controllable_BtoR_REQ0 & ~n31756;
  assign n31758 = ~n28833 & ~n31757;
  assign n31759 = ~i_RtoB_ACK0 & ~n31758;
  assign n31760 = ~n29625 & ~n31759;
  assign n31761 = ~controllable_DEQ & ~n31760;
  assign n31762 = ~n29653 & ~n31761;
  assign n31763 = i_FULL & ~n31762;
  assign n31764 = ~n19053 & ~n27878;
  assign n31765 = ~controllable_BtoR_REQ0 & ~n31764;
  assign n31766 = ~n28803 & ~n31765;
  assign n31767 = ~i_RtoB_ACK0 & ~n31766;
  assign n31768 = ~n29625 & ~n31767;
  assign n31769 = ~controllable_DEQ & ~n31768;
  assign n31770 = ~n29663 & ~n31769;
  assign n31771 = ~i_FULL & ~n31770;
  assign n31772 = ~n31763 & ~n31771;
  assign n31773 = ~i_nEMPTY & ~n31772;
  assign n31774 = ~n31755 & ~n31773;
  assign n31775 = ~controllable_BtoS_ACK0 & ~n31774;
  assign n31776 = ~n21013 & ~n31775;
  assign n31777 = ~n4465 & ~n31776;
  assign n31778 = ~n31731 & ~n31777;
  assign n31779 = i_StoB_REQ10 & ~n31778;
  assign n31780 = ~n11236 & ~n19386;
  assign n31781 = ~controllable_BtoR_REQ0 & ~n31780;
  assign n31782 = ~n28857 & ~n31781;
  assign n31783 = ~i_RtoB_ACK0 & ~n31782;
  assign n31784 = ~n23089 & ~n31783;
  assign n31785 = controllable_DEQ & ~n31784;
  assign n31786 = controllable_BtoR_REQ1 & ~n9301;
  assign n31787 = ~n19395 & ~n31786;
  assign n31788 = ~controllable_BtoR_REQ0 & ~n31787;
  assign n31789 = ~n28865 & ~n31788;
  assign n31790 = ~i_RtoB_ACK0 & ~n31789;
  assign n31791 = ~n23095 & ~n31790;
  assign n31792 = ~controllable_DEQ & ~n31791;
  assign n31793 = ~n31785 & ~n31792;
  assign n31794 = i_FULL & ~n31793;
  assign n31795 = ~n19411 & ~n31786;
  assign n31796 = ~controllable_BtoR_REQ0 & ~n31795;
  assign n31797 = ~n28875 & ~n31796;
  assign n31798 = ~i_RtoB_ACK0 & ~n31797;
  assign n31799 = ~n23095 & ~n31798;
  assign n31800 = ~controllable_DEQ & ~n31799;
  assign n31801 = ~n23093 & ~n31800;
  assign n31802 = ~i_FULL & ~n31801;
  assign n31803 = ~n31794 & ~n31802;
  assign n31804 = i_nEMPTY & ~n31803;
  assign n31805 = controllable_BtoR_REQ1 & ~n9570;
  assign n31806 = ~n19429 & ~n31805;
  assign n31807 = ~controllable_BtoR_REQ0 & ~n31806;
  assign n31808 = ~n28887 & ~n31807;
  assign n31809 = ~i_RtoB_ACK0 & ~n31808;
  assign n31810 = ~n23107 & ~n31809;
  assign n31811 = ~controllable_DEQ & ~n31810;
  assign n31812 = ~n23105 & ~n31811;
  assign n31813 = i_FULL & ~n31812;
  assign n31814 = ~n11236 & ~n28001;
  assign n31815 = ~controllable_BtoR_REQ0 & ~n31814;
  assign n31816 = ~n28857 & ~n31815;
  assign n31817 = ~i_RtoB_ACK0 & ~n31816;
  assign n31818 = ~n23089 & ~n31817;
  assign n31819 = ~controllable_DEQ & ~n31818;
  assign n31820 = ~n23117 & ~n31819;
  assign n31821 = ~i_FULL & ~n31820;
  assign n31822 = ~n31813 & ~n31821;
  assign n31823 = ~i_nEMPTY & ~n31822;
  assign n31824 = ~n31804 & ~n31823;
  assign n31825 = controllable_BtoS_ACK0 & ~n31824;
  assign n31826 = ~n11315 & ~n19452;
  assign n31827 = ~controllable_BtoR_REQ0 & ~n31826;
  assign n31828 = ~n28909 & ~n31827;
  assign n31829 = ~i_RtoB_ACK0 & ~n31828;
  assign n31830 = ~n23129 & ~n31829;
  assign n31831 = controllable_DEQ & ~n31830;
  assign n31832 = controllable_BtoR_REQ1 & ~n9634;
  assign n31833 = ~n19461 & ~n31832;
  assign n31834 = ~controllable_BtoR_REQ0 & ~n31833;
  assign n31835 = ~n28917 & ~n31834;
  assign n31836 = ~i_RtoB_ACK0 & ~n31835;
  assign n31837 = ~n23135 & ~n31836;
  assign n31838 = ~controllable_DEQ & ~n31837;
  assign n31839 = ~n31831 & ~n31838;
  assign n31840 = i_FULL & ~n31839;
  assign n31841 = ~n19477 & ~n31832;
  assign n31842 = ~controllable_BtoR_REQ0 & ~n31841;
  assign n31843 = ~n28927 & ~n31842;
  assign n31844 = ~i_RtoB_ACK0 & ~n31843;
  assign n31845 = ~n23135 & ~n31844;
  assign n31846 = ~controllable_DEQ & ~n31845;
  assign n31847 = ~n23133 & ~n31846;
  assign n31848 = ~i_FULL & ~n31847;
  assign n31849 = ~n31840 & ~n31848;
  assign n31850 = i_nEMPTY & ~n31849;
  assign n31851 = controllable_BtoR_REQ1 & ~n9717;
  assign n31852 = ~n19495 & ~n31851;
  assign n31853 = ~controllable_BtoR_REQ0 & ~n31852;
  assign n31854 = ~n28939 & ~n31853;
  assign n31855 = ~i_RtoB_ACK0 & ~n31854;
  assign n31856 = ~n23147 & ~n31855;
  assign n31857 = ~controllable_DEQ & ~n31856;
  assign n31858 = ~n23145 & ~n31857;
  assign n31859 = i_FULL & ~n31858;
  assign n31860 = ~n11315 & ~n28046;
  assign n31861 = ~controllable_BtoR_REQ0 & ~n31860;
  assign n31862 = ~n28909 & ~n31861;
  assign n31863 = ~i_RtoB_ACK0 & ~n31862;
  assign n31864 = ~n23129 & ~n31863;
  assign n31865 = ~controllable_DEQ & ~n31864;
  assign n31866 = ~n23157 & ~n31865;
  assign n31867 = ~i_FULL & ~n31866;
  assign n31868 = ~n31859 & ~n31867;
  assign n31869 = ~i_nEMPTY & ~n31868;
  assign n31870 = ~n31850 & ~n31869;
  assign n31871 = ~controllable_BtoS_ACK0 & ~n31870;
  assign n31872 = ~n31825 & ~n31871;
  assign n31873 = n4465 & ~n31872;
  assign n31874 = ~n11315 & ~n19313;
  assign n31875 = ~controllable_BtoR_REQ0 & ~n31874;
  assign n31876 = ~n28963 & ~n31875;
  assign n31877 = ~i_RtoB_ACK0 & ~n31876;
  assign n31878 = ~n23129 & ~n31877;
  assign n31879 = controllable_DEQ & ~n31878;
  assign n31880 = ~n19321 & ~n31832;
  assign n31881 = ~controllable_BtoR_REQ0 & ~n31880;
  assign n31882 = ~n28971 & ~n31881;
  assign n31883 = ~i_RtoB_ACK0 & ~n31882;
  assign n31884 = ~n23135 & ~n31883;
  assign n31885 = ~controllable_DEQ & ~n31884;
  assign n31886 = ~n31879 & ~n31885;
  assign n31887 = i_FULL & ~n31886;
  assign n31888 = ~n19335 & ~n31832;
  assign n31889 = ~controllable_BtoR_REQ0 & ~n31888;
  assign n31890 = ~n28981 & ~n31889;
  assign n31891 = ~i_RtoB_ACK0 & ~n31890;
  assign n31892 = ~n23135 & ~n31891;
  assign n31893 = ~controllable_DEQ & ~n31892;
  assign n31894 = ~n23133 & ~n31893;
  assign n31895 = ~i_FULL & ~n31894;
  assign n31896 = ~n31887 & ~n31895;
  assign n31897 = i_nEMPTY & ~n31896;
  assign n31898 = ~n19351 & ~n31851;
  assign n31899 = ~controllable_BtoR_REQ0 & ~n31898;
  assign n31900 = ~n28993 & ~n31899;
  assign n31901 = ~i_RtoB_ACK0 & ~n31900;
  assign n31902 = ~n23147 & ~n31901;
  assign n31903 = ~controllable_DEQ & ~n31902;
  assign n31904 = ~n23145 & ~n31903;
  assign n31905 = i_FULL & ~n31904;
  assign n31906 = ~n11315 & ~n19365;
  assign n31907 = ~controllable_BtoR_REQ0 & ~n31906;
  assign n31908 = ~n28963 & ~n31907;
  assign n31909 = ~i_RtoB_ACK0 & ~n31908;
  assign n31910 = ~n23129 & ~n31909;
  assign n31911 = ~controllable_DEQ & ~n31910;
  assign n31912 = ~n23157 & ~n31911;
  assign n31913 = ~i_FULL & ~n31912;
  assign n31914 = ~n31905 & ~n31913;
  assign n31915 = ~i_nEMPTY & ~n31914;
  assign n31916 = ~n31897 & ~n31915;
  assign n31917 = ~controllable_BtoS_ACK0 & ~n31916;
  assign n31918 = ~n23127 & ~n31917;
  assign n31919 = ~n4465 & ~n31918;
  assign n31920 = ~n31873 & ~n31919;
  assign n31921 = ~i_StoB_REQ10 & ~n31920;
  assign n31922 = ~n31779 & ~n31921;
  assign n31923 = controllable_BtoS_ACK10 & ~n31922;
  assign n31924 = ~n19386 & ~n28133;
  assign n31925 = ~controllable_BtoR_REQ0 & ~n31924;
  assign n31926 = ~n29826 & ~n31925;
  assign n31927 = ~i_RtoB_ACK0 & ~n31926;
  assign n31928 = ~n29825 & ~n31927;
  assign n31929 = controllable_DEQ & ~n31928;
  assign n31930 = ~n29833 & ~n31788;
  assign n31931 = ~i_RtoB_ACK0 & ~n31930;
  assign n31932 = ~n29832 & ~n31931;
  assign n31933 = ~controllable_DEQ & ~n31932;
  assign n31934 = ~n31929 & ~n31933;
  assign n31935 = i_FULL & ~n31934;
  assign n31936 = ~n29845 & ~n31796;
  assign n31937 = ~i_RtoB_ACK0 & ~n31936;
  assign n31938 = ~n29832 & ~n31937;
  assign n31939 = ~controllable_DEQ & ~n31938;
  assign n31940 = ~n29844 & ~n31939;
  assign n31941 = ~i_FULL & ~n31940;
  assign n31942 = ~n31935 & ~n31941;
  assign n31943 = i_nEMPTY & ~n31942;
  assign n31944 = ~n29861 & ~n31807;
  assign n31945 = ~i_RtoB_ACK0 & ~n31944;
  assign n31946 = ~n29860 & ~n31945;
  assign n31947 = ~controllable_DEQ & ~n31946;
  assign n31948 = ~n29858 & ~n31947;
  assign n31949 = i_FULL & ~n31948;
  assign n31950 = ~controllable_DEQ & ~n31928;
  assign n31951 = ~n29872 & ~n31950;
  assign n31952 = ~i_FULL & ~n31951;
  assign n31953 = ~n31949 & ~n31952;
  assign n31954 = ~i_nEMPTY & ~n31953;
  assign n31955 = ~n31943 & ~n31954;
  assign n31956 = controllable_BtoS_ACK0 & ~n31955;
  assign n31957 = ~n19452 & ~n28194;
  assign n31958 = ~controllable_BtoR_REQ0 & ~n31957;
  assign n31959 = ~n29882 & ~n31958;
  assign n31960 = ~i_RtoB_ACK0 & ~n31959;
  assign n31961 = ~n29881 & ~n31960;
  assign n31962 = controllable_DEQ & ~n31961;
  assign n31963 = ~n29889 & ~n31834;
  assign n31964 = ~i_RtoB_ACK0 & ~n31963;
  assign n31965 = ~n29888 & ~n31964;
  assign n31966 = ~controllable_DEQ & ~n31965;
  assign n31967 = ~n31962 & ~n31966;
  assign n31968 = i_FULL & ~n31967;
  assign n31969 = ~n29901 & ~n31842;
  assign n31970 = ~i_RtoB_ACK0 & ~n31969;
  assign n31971 = ~n29888 & ~n31970;
  assign n31972 = ~controllable_DEQ & ~n31971;
  assign n31973 = ~n29900 & ~n31972;
  assign n31974 = ~i_FULL & ~n31973;
  assign n31975 = ~n31968 & ~n31974;
  assign n31976 = i_nEMPTY & ~n31975;
  assign n31977 = ~n29917 & ~n31853;
  assign n31978 = ~i_RtoB_ACK0 & ~n31977;
  assign n31979 = ~n29916 & ~n31978;
  assign n31980 = ~controllable_DEQ & ~n31979;
  assign n31981 = ~n29914 & ~n31980;
  assign n31982 = i_FULL & ~n31981;
  assign n31983 = ~controllable_DEQ & ~n31961;
  assign n31984 = ~n29928 & ~n31983;
  assign n31985 = ~i_FULL & ~n31984;
  assign n31986 = ~n31982 & ~n31985;
  assign n31987 = ~i_nEMPTY & ~n31986;
  assign n31988 = ~n31976 & ~n31987;
  assign n31989 = ~controllable_BtoS_ACK0 & ~n31988;
  assign n31990 = ~n31956 & ~n31989;
  assign n31991 = n4465 & ~n31990;
  assign n31992 = ~n19313 & ~n28194;
  assign n31993 = ~controllable_BtoR_REQ0 & ~n31992;
  assign n31994 = ~n29959 & ~n31993;
  assign n31995 = ~i_RtoB_ACK0 & ~n31994;
  assign n31996 = ~n29881 & ~n31995;
  assign n31997 = controllable_DEQ & ~n31996;
  assign n31998 = ~n29964 & ~n31881;
  assign n31999 = ~i_RtoB_ACK0 & ~n31998;
  assign n32000 = ~n29888 & ~n31999;
  assign n32001 = ~controllable_DEQ & ~n32000;
  assign n32002 = ~n31997 & ~n32001;
  assign n32003 = i_FULL & ~n32002;
  assign n32004 = ~n29971 & ~n31889;
  assign n32005 = ~i_RtoB_ACK0 & ~n32004;
  assign n32006 = ~n29888 & ~n32005;
  assign n32007 = ~controllable_DEQ & ~n32006;
  assign n32008 = ~n29900 & ~n32007;
  assign n32009 = ~i_FULL & ~n32008;
  assign n32010 = ~n32003 & ~n32009;
  assign n32011 = i_nEMPTY & ~n32010;
  assign n32012 = ~n29980 & ~n31899;
  assign n32013 = ~i_RtoB_ACK0 & ~n32012;
  assign n32014 = ~n29916 & ~n32013;
  assign n32015 = ~controllable_DEQ & ~n32014;
  assign n32016 = ~n29914 & ~n32015;
  assign n32017 = i_FULL & ~n32016;
  assign n32018 = ~controllable_DEQ & ~n31996;
  assign n32019 = ~n29928 & ~n32018;
  assign n32020 = ~i_FULL & ~n32019;
  assign n32021 = ~n32017 & ~n32020;
  assign n32022 = ~i_nEMPTY & ~n32021;
  assign n32023 = ~n32011 & ~n32022;
  assign n32024 = ~controllable_BtoS_ACK0 & ~n32023;
  assign n32025 = ~n29958 & ~n32024;
  assign n32026 = ~n4465 & ~n32025;
  assign n32027 = ~n31991 & ~n32026;
  assign n32028 = i_StoB_REQ10 & ~n32027;
  assign n32029 = ~n31921 & ~n32028;
  assign n32030 = ~controllable_BtoS_ACK10 & ~n32029;
  assign n32031 = ~n31923 & ~n32030;
  assign n32032 = n4464 & ~n32031;
  assign n32033 = ~n5242 & ~n19613;
  assign n32034 = ~controllable_BtoR_REQ0 & ~n32033;
  assign n32035 = ~n29157 & ~n32034;
  assign n32036 = ~i_RtoB_ACK0 & ~n32035;
  assign n32037 = ~n20977 & ~n32036;
  assign n32038 = controllable_DEQ & ~n32037;
  assign n32039 = ~n19620 & ~n31644;
  assign n32040 = ~controllable_BtoR_REQ0 & ~n32039;
  assign n32041 = ~n29165 & ~n32040;
  assign n32042 = ~i_RtoB_ACK0 & ~n32041;
  assign n32043 = ~n20983 & ~n32042;
  assign n32044 = ~controllable_DEQ & ~n32043;
  assign n32045 = ~n32038 & ~n32044;
  assign n32046 = i_FULL & ~n32045;
  assign n32047 = ~n19634 & ~n31644;
  assign n32048 = ~controllable_BtoR_REQ0 & ~n32047;
  assign n32049 = ~n29175 & ~n32048;
  assign n32050 = ~i_RtoB_ACK0 & ~n32049;
  assign n32051 = ~n20983 & ~n32050;
  assign n32052 = ~controllable_DEQ & ~n32051;
  assign n32053 = ~n20981 & ~n32052;
  assign n32054 = ~i_FULL & ~n32053;
  assign n32055 = ~n32046 & ~n32054;
  assign n32056 = i_nEMPTY & ~n32055;
  assign n32057 = ~n19649 & ~n31663;
  assign n32058 = ~controllable_BtoR_REQ0 & ~n32057;
  assign n32059 = ~n29187 & ~n32058;
  assign n32060 = ~i_RtoB_ACK0 & ~n32059;
  assign n32061 = ~n20977 & ~n32060;
  assign n32062 = ~controllable_DEQ & ~n32061;
  assign n32063 = ~n20993 & ~n32062;
  assign n32064 = i_FULL & ~n32063;
  assign n32065 = ~n5242 & ~n19663;
  assign n32066 = ~controllable_BtoR_REQ0 & ~n32065;
  assign n32067 = ~n29157 & ~n32066;
  assign n32068 = ~i_RtoB_ACK0 & ~n32067;
  assign n32069 = ~n20977 & ~n32068;
  assign n32070 = ~controllable_DEQ & ~n32069;
  assign n32071 = ~n21003 & ~n32070;
  assign n32072 = ~i_FULL & ~n32071;
  assign n32073 = ~n32064 & ~n32072;
  assign n32074 = ~i_nEMPTY & ~n32073;
  assign n32075 = ~n32056 & ~n32074;
  assign n32076 = controllable_BtoS_ACK0 & ~n32075;
  assign n32077 = ~n19677 & ~n27878;
  assign n32078 = ~controllable_BtoR_REQ0 & ~n32077;
  assign n32079 = ~n29207 & ~n32078;
  assign n32080 = ~i_RtoB_ACK0 & ~n32079;
  assign n32081 = ~n29625 & ~n32080;
  assign n32082 = controllable_DEQ & ~n32081;
  assign n32083 = ~n19684 & ~n31690;
  assign n32084 = ~controllable_BtoR_REQ0 & ~n32083;
  assign n32085 = ~n29215 & ~n32084;
  assign n32086 = ~i_RtoB_ACK0 & ~n32085;
  assign n32087 = ~n29631 & ~n32086;
  assign n32088 = ~controllable_DEQ & ~n32087;
  assign n32089 = ~n32082 & ~n32088;
  assign n32090 = i_FULL & ~n32089;
  assign n32091 = ~n19698 & ~n31690;
  assign n32092 = ~controllable_BtoR_REQ0 & ~n32091;
  assign n32093 = ~n29225 & ~n32092;
  assign n32094 = ~i_RtoB_ACK0 & ~n32093;
  assign n32095 = ~n29631 & ~n32094;
  assign n32096 = ~controllable_DEQ & ~n32095;
  assign n32097 = ~n29641 & ~n32096;
  assign n32098 = ~i_FULL & ~n32097;
  assign n32099 = ~n32090 & ~n32098;
  assign n32100 = i_nEMPTY & ~n32099;
  assign n32101 = ~n19713 & ~n31709;
  assign n32102 = ~controllable_BtoR_REQ0 & ~n32101;
  assign n32103 = ~n29237 & ~n32102;
  assign n32104 = ~i_RtoB_ACK0 & ~n32103;
  assign n32105 = ~n29625 & ~n32104;
  assign n32106 = ~controllable_DEQ & ~n32105;
  assign n32107 = ~n29653 & ~n32106;
  assign n32108 = i_FULL & ~n32107;
  assign n32109 = ~n19727 & ~n27878;
  assign n32110 = ~controllable_BtoR_REQ0 & ~n32109;
  assign n32111 = ~n29207 & ~n32110;
  assign n32112 = ~i_RtoB_ACK0 & ~n32111;
  assign n32113 = ~n29625 & ~n32112;
  assign n32114 = ~controllable_DEQ & ~n32113;
  assign n32115 = ~n29663 & ~n32114;
  assign n32116 = ~i_FULL & ~n32115;
  assign n32117 = ~n32108 & ~n32116;
  assign n32118 = ~i_nEMPTY & ~n32117;
  assign n32119 = ~n32100 & ~n32118;
  assign n32120 = ~controllable_BtoS_ACK0 & ~n32119;
  assign n32121 = ~n32076 & ~n32120;
  assign n32122 = n4465 & ~n32121;
  assign n32123 = ~n21013 & ~n32120;
  assign n32124 = ~n4465 & ~n32123;
  assign n32125 = ~n32122 & ~n32124;
  assign n32126 = i_StoB_REQ10 & ~n32125;
  assign n32127 = ~n11236 & ~n20004;
  assign n32128 = ~controllable_BtoR_REQ0 & ~n32127;
  assign n32129 = ~n29263 & ~n32128;
  assign n32130 = ~i_RtoB_ACK0 & ~n32129;
  assign n32131 = ~n23089 & ~n32130;
  assign n32132 = controllable_DEQ & ~n32131;
  assign n32133 = ~n20013 & ~n31786;
  assign n32134 = ~controllable_BtoR_REQ0 & ~n32133;
  assign n32135 = ~n29271 & ~n32134;
  assign n32136 = ~i_RtoB_ACK0 & ~n32135;
  assign n32137 = ~n23095 & ~n32136;
  assign n32138 = ~controllable_DEQ & ~n32137;
  assign n32139 = ~n32132 & ~n32138;
  assign n32140 = i_FULL & ~n32139;
  assign n32141 = ~n20029 & ~n31786;
  assign n32142 = ~controllable_BtoR_REQ0 & ~n32141;
  assign n32143 = ~n29281 & ~n32142;
  assign n32144 = ~i_RtoB_ACK0 & ~n32143;
  assign n32145 = ~n23095 & ~n32144;
  assign n32146 = ~controllable_DEQ & ~n32145;
  assign n32147 = ~n23093 & ~n32146;
  assign n32148 = ~i_FULL & ~n32147;
  assign n32149 = ~n32140 & ~n32148;
  assign n32150 = i_nEMPTY & ~n32149;
  assign n32151 = ~n20047 & ~n31805;
  assign n32152 = ~controllable_BtoR_REQ0 & ~n32151;
  assign n32153 = ~n29293 & ~n32152;
  assign n32154 = ~i_RtoB_ACK0 & ~n32153;
  assign n32155 = ~n23107 & ~n32154;
  assign n32156 = ~controllable_DEQ & ~n32155;
  assign n32157 = ~n23105 & ~n32156;
  assign n32158 = i_FULL & ~n32157;
  assign n32159 = ~n11236 & ~n20823;
  assign n32160 = ~controllable_BtoR_REQ0 & ~n32159;
  assign n32161 = ~n29263 & ~n32160;
  assign n32162 = ~i_RtoB_ACK0 & ~n32161;
  assign n32163 = ~n23089 & ~n32162;
  assign n32164 = ~controllable_DEQ & ~n32163;
  assign n32165 = ~n23117 & ~n32164;
  assign n32166 = ~i_FULL & ~n32165;
  assign n32167 = ~n32158 & ~n32166;
  assign n32168 = ~i_nEMPTY & ~n32167;
  assign n32169 = ~n32150 & ~n32168;
  assign n32170 = controllable_BtoS_ACK0 & ~n32169;
  assign n32171 = ~n11315 & ~n19931;
  assign n32172 = ~controllable_BtoR_REQ0 & ~n32171;
  assign n32173 = ~n29313 & ~n32172;
  assign n32174 = ~i_RtoB_ACK0 & ~n32173;
  assign n32175 = ~n23129 & ~n32174;
  assign n32176 = controllable_DEQ & ~n32175;
  assign n32177 = ~n19939 & ~n31832;
  assign n32178 = ~controllable_BtoR_REQ0 & ~n32177;
  assign n32179 = ~n29321 & ~n32178;
  assign n32180 = ~i_RtoB_ACK0 & ~n32179;
  assign n32181 = ~n23135 & ~n32180;
  assign n32182 = ~controllable_DEQ & ~n32181;
  assign n32183 = ~n32176 & ~n32182;
  assign n32184 = i_FULL & ~n32183;
  assign n32185 = ~n19953 & ~n31832;
  assign n32186 = ~controllable_BtoR_REQ0 & ~n32185;
  assign n32187 = ~n29331 & ~n32186;
  assign n32188 = ~i_RtoB_ACK0 & ~n32187;
  assign n32189 = ~n23135 & ~n32188;
  assign n32190 = ~controllable_DEQ & ~n32189;
  assign n32191 = ~n23133 & ~n32190;
  assign n32192 = ~i_FULL & ~n32191;
  assign n32193 = ~n32184 & ~n32192;
  assign n32194 = i_nEMPTY & ~n32193;
  assign n32195 = ~n19969 & ~n31851;
  assign n32196 = ~controllable_BtoR_REQ0 & ~n32195;
  assign n32197 = ~n29343 & ~n32196;
  assign n32198 = ~i_RtoB_ACK0 & ~n32197;
  assign n32199 = ~n23147 & ~n32198;
  assign n32200 = ~controllable_DEQ & ~n32199;
  assign n32201 = ~n23145 & ~n32200;
  assign n32202 = i_FULL & ~n32201;
  assign n32203 = ~n11315 & ~n19983;
  assign n32204 = ~controllable_BtoR_REQ0 & ~n32203;
  assign n32205 = ~n29313 & ~n32204;
  assign n32206 = ~i_RtoB_ACK0 & ~n32205;
  assign n32207 = ~n23129 & ~n32206;
  assign n32208 = ~controllable_DEQ & ~n32207;
  assign n32209 = ~n23157 & ~n32208;
  assign n32210 = ~i_FULL & ~n32209;
  assign n32211 = ~n32202 & ~n32210;
  assign n32212 = ~i_nEMPTY & ~n32211;
  assign n32213 = ~n32194 & ~n32212;
  assign n32214 = ~controllable_BtoS_ACK0 & ~n32213;
  assign n32215 = ~n32170 & ~n32214;
  assign n32216 = n4465 & ~n32215;
  assign n32217 = ~n23127 & ~n32214;
  assign n32218 = ~n4465 & ~n32217;
  assign n32219 = ~n32216 & ~n32218;
  assign n32220 = ~i_StoB_REQ10 & ~n32219;
  assign n32221 = ~n32126 & ~n32220;
  assign n32222 = controllable_BtoS_ACK10 & ~n32221;
  assign n32223 = ~n20004 & ~n28133;
  assign n32224 = ~controllable_BtoR_REQ0 & ~n32223;
  assign n32225 = ~n30152 & ~n32224;
  assign n32226 = ~i_RtoB_ACK0 & ~n32225;
  assign n32227 = ~n29825 & ~n32226;
  assign n32228 = controllable_DEQ & ~n32227;
  assign n32229 = ~n30157 & ~n32134;
  assign n32230 = ~i_RtoB_ACK0 & ~n32229;
  assign n32231 = ~n29832 & ~n32230;
  assign n32232 = ~controllable_DEQ & ~n32231;
  assign n32233 = ~n32228 & ~n32232;
  assign n32234 = i_FULL & ~n32233;
  assign n32235 = ~n30164 & ~n32142;
  assign n32236 = ~i_RtoB_ACK0 & ~n32235;
  assign n32237 = ~n29832 & ~n32236;
  assign n32238 = ~controllable_DEQ & ~n32237;
  assign n32239 = ~n29844 & ~n32238;
  assign n32240 = ~i_FULL & ~n32239;
  assign n32241 = ~n32234 & ~n32240;
  assign n32242 = i_nEMPTY & ~n32241;
  assign n32243 = ~n30173 & ~n32152;
  assign n32244 = ~i_RtoB_ACK0 & ~n32243;
  assign n32245 = ~n29860 & ~n32244;
  assign n32246 = ~controllable_DEQ & ~n32245;
  assign n32247 = ~n29858 & ~n32246;
  assign n32248 = i_FULL & ~n32247;
  assign n32249 = ~controllable_DEQ & ~n32227;
  assign n32250 = ~n29872 & ~n32249;
  assign n32251 = ~i_FULL & ~n32250;
  assign n32252 = ~n32248 & ~n32251;
  assign n32253 = ~i_nEMPTY & ~n32252;
  assign n32254 = ~n32242 & ~n32253;
  assign n32255 = controllable_BtoS_ACK0 & ~n32254;
  assign n32256 = ~n19931 & ~n28194;
  assign n32257 = ~controllable_BtoR_REQ0 & ~n32256;
  assign n32258 = ~n30187 & ~n32257;
  assign n32259 = ~i_RtoB_ACK0 & ~n32258;
  assign n32260 = ~n29881 & ~n32259;
  assign n32261 = controllable_DEQ & ~n32260;
  assign n32262 = ~n30192 & ~n32178;
  assign n32263 = ~i_RtoB_ACK0 & ~n32262;
  assign n32264 = ~n29888 & ~n32263;
  assign n32265 = ~controllable_DEQ & ~n32264;
  assign n32266 = ~n32261 & ~n32265;
  assign n32267 = i_FULL & ~n32266;
  assign n32268 = ~n30199 & ~n32186;
  assign n32269 = ~i_RtoB_ACK0 & ~n32268;
  assign n32270 = ~n29888 & ~n32269;
  assign n32271 = ~controllable_DEQ & ~n32270;
  assign n32272 = ~n29900 & ~n32271;
  assign n32273 = ~i_FULL & ~n32272;
  assign n32274 = ~n32267 & ~n32273;
  assign n32275 = i_nEMPTY & ~n32274;
  assign n32276 = ~n30208 & ~n32196;
  assign n32277 = ~i_RtoB_ACK0 & ~n32276;
  assign n32278 = ~n29916 & ~n32277;
  assign n32279 = ~controllable_DEQ & ~n32278;
  assign n32280 = ~n29914 & ~n32279;
  assign n32281 = i_FULL & ~n32280;
  assign n32282 = ~controllable_DEQ & ~n32260;
  assign n32283 = ~n29928 & ~n32282;
  assign n32284 = ~i_FULL & ~n32283;
  assign n32285 = ~n32281 & ~n32284;
  assign n32286 = ~i_nEMPTY & ~n32285;
  assign n32287 = ~n32275 & ~n32286;
  assign n32288 = ~controllable_BtoS_ACK0 & ~n32287;
  assign n32289 = ~n32255 & ~n32288;
  assign n32290 = n4465 & ~n32289;
  assign n32291 = ~n29958 & ~n32288;
  assign n32292 = ~n4465 & ~n32291;
  assign n32293 = ~n32290 & ~n32292;
  assign n32294 = i_StoB_REQ10 & ~n32293;
  assign n32295 = ~n32220 & ~n32294;
  assign n32296 = ~controllable_BtoS_ACK10 & ~n32295;
  assign n32297 = ~n32222 & ~n32296;
  assign n32298 = ~n4464 & ~n32297;
  assign n32299 = ~n32032 & ~n32298;
  assign n32300 = ~n4463 & ~n32299;
  assign n32301 = ~n30233 & ~n32300;
  assign n32302 = n4462 & ~n32301;
  assign n32303 = ~n20368 & ~n28133;
  assign n32304 = ~controllable_BtoR_REQ0 & ~n32303;
  assign n32305 = ~n30807 & ~n32304;
  assign n32306 = ~i_RtoB_ACK0 & ~n32305;
  assign n32307 = ~n29825 & ~n32306;
  assign n32308 = controllable_DEQ & ~n32307;
  assign n32309 = ~n20377 & ~n31786;
  assign n32310 = ~controllable_BtoR_REQ0 & ~n32309;
  assign n32311 = ~n30812 & ~n32310;
  assign n32312 = ~i_RtoB_ACK0 & ~n32311;
  assign n32313 = ~n29832 & ~n32312;
  assign n32314 = ~controllable_DEQ & ~n32313;
  assign n32315 = ~n32308 & ~n32314;
  assign n32316 = i_FULL & ~n32315;
  assign n32317 = ~n20393 & ~n31786;
  assign n32318 = ~controllable_BtoR_REQ0 & ~n32317;
  assign n32319 = ~n30819 & ~n32318;
  assign n32320 = ~i_RtoB_ACK0 & ~n32319;
  assign n32321 = ~n29832 & ~n32320;
  assign n32322 = ~controllable_DEQ & ~n32321;
  assign n32323 = ~n29844 & ~n32322;
  assign n32324 = ~i_FULL & ~n32323;
  assign n32325 = ~n32316 & ~n32324;
  assign n32326 = i_nEMPTY & ~n32325;
  assign n32327 = ~n20411 & ~n31805;
  assign n32328 = ~controllable_BtoR_REQ0 & ~n32327;
  assign n32329 = ~n30828 & ~n32328;
  assign n32330 = ~i_RtoB_ACK0 & ~n32329;
  assign n32331 = ~n29860 & ~n32330;
  assign n32332 = ~controllable_DEQ & ~n32331;
  assign n32333 = ~n29858 & ~n32332;
  assign n32334 = i_FULL & ~n32333;
  assign n32335 = ~controllable_DEQ & ~n32307;
  assign n32336 = ~n29872 & ~n32335;
  assign n32337 = ~i_FULL & ~n32336;
  assign n32338 = ~n32334 & ~n32337;
  assign n32339 = ~i_nEMPTY & ~n32338;
  assign n32340 = ~n32326 & ~n32339;
  assign n32341 = controllable_BtoS_ACK0 & ~n32340;
  assign n32342 = ~n32024 & ~n32341;
  assign n32343 = n4465 & ~n32342;
  assign n32344 = ~n32026 & ~n32343;
  assign n32345 = i_StoB_REQ10 & ~n32344;
  assign n32346 = ~n11236 & ~n20368;
  assign n32347 = ~controllable_BtoR_REQ0 & ~n32346;
  assign n32348 = ~n29502 & ~n32347;
  assign n32349 = ~i_RtoB_ACK0 & ~n32348;
  assign n32350 = ~n23089 & ~n32349;
  assign n32351 = controllable_DEQ & ~n32350;
  assign n32352 = ~n29510 & ~n32310;
  assign n32353 = ~i_RtoB_ACK0 & ~n32352;
  assign n32354 = ~n23095 & ~n32353;
  assign n32355 = ~controllable_DEQ & ~n32354;
  assign n32356 = ~n32351 & ~n32355;
  assign n32357 = i_FULL & ~n32356;
  assign n32358 = ~n29520 & ~n32318;
  assign n32359 = ~i_RtoB_ACK0 & ~n32358;
  assign n32360 = ~n23095 & ~n32359;
  assign n32361 = ~controllable_DEQ & ~n32360;
  assign n32362 = ~n23093 & ~n32361;
  assign n32363 = ~i_FULL & ~n32362;
  assign n32364 = ~n32357 & ~n32363;
  assign n32365 = i_nEMPTY & ~n32364;
  assign n32366 = ~n29532 & ~n32328;
  assign n32367 = ~i_RtoB_ACK0 & ~n32366;
  assign n32368 = ~n23107 & ~n32367;
  assign n32369 = ~controllable_DEQ & ~n32368;
  assign n32370 = ~n23105 & ~n32369;
  assign n32371 = i_FULL & ~n32370;
  assign n32372 = ~n11236 & ~n20525;
  assign n32373 = ~controllable_BtoR_REQ0 & ~n32372;
  assign n32374 = ~n29502 & ~n32373;
  assign n32375 = ~i_RtoB_ACK0 & ~n32374;
  assign n32376 = ~n23089 & ~n32375;
  assign n32377 = ~controllable_DEQ & ~n32376;
  assign n32378 = ~n23117 & ~n32377;
  assign n32379 = ~i_FULL & ~n32378;
  assign n32380 = ~n32371 & ~n32379;
  assign n32381 = ~i_nEMPTY & ~n32380;
  assign n32382 = ~n32365 & ~n32381;
  assign n32383 = controllable_BtoS_ACK0 & ~n32382;
  assign n32384 = ~n31917 & ~n32383;
  assign n32385 = n4465 & ~n32384;
  assign n32386 = ~n31919 & ~n32385;
  assign n32387 = ~i_StoB_REQ10 & ~n32386;
  assign n32388 = ~n32345 & ~n32387;
  assign n32389 = ~controllable_BtoS_ACK10 & ~n32388;
  assign n32390 = ~n30806 & ~n32389;
  assign n32391 = n4464 & ~n32390;
  assign n32392 = ~n30806 & ~n32296;
  assign n32393 = ~n4464 & ~n32392;
  assign n32394 = ~n32391 & ~n32393;
  assign n32395 = ~n4463 & ~n32394;
  assign n32396 = ~n30891 & ~n32395;
  assign n32397 = ~n4462 & ~n32396;
  assign n32398 = ~n32302 & ~n32397;
  assign n32399 = n4461 & ~n32398;
  assign n32400 = ~n5245 & ~n27814;
  assign n32401 = ~controllable_BtoR_REQ0 & ~n32400;
  assign n32402 = ~n14749 & ~n32401;
  assign n32403 = ~i_RtoB_ACK0 & ~n32402;
  assign n32404 = ~n20977 & ~n32403;
  assign n32405 = controllable_DEQ & ~n32404;
  assign n32406 = ~n5255 & ~n8782;
  assign n32407 = ~controllable_BtoR_REQ0 & ~n32406;
  assign n32408 = ~n14765 & ~n32407;
  assign n32409 = ~i_RtoB_ACK0 & ~n32408;
  assign n32410 = ~n20983 & ~n32409;
  assign n32411 = ~controllable_DEQ & ~n32410;
  assign n32412 = ~n32405 & ~n32411;
  assign n32413 = i_FULL & ~n32412;
  assign n32414 = controllable_BtoR_REQ1 & ~n18887;
  assign n32415 = ~n5255 & ~n32414;
  assign n32416 = ~controllable_BtoR_REQ0 & ~n32415;
  assign n32417 = ~n14765 & ~n32416;
  assign n32418 = ~i_RtoB_ACK0 & ~n32417;
  assign n32419 = ~n20983 & ~n32418;
  assign n32420 = ~controllable_DEQ & ~n32419;
  assign n32421 = ~n20981 & ~n32420;
  assign n32422 = ~i_FULL & ~n32421;
  assign n32423 = ~n32413 & ~n32422;
  assign n32424 = i_nEMPTY & ~n32423;
  assign n32425 = ~n5232 & ~n8819;
  assign n32426 = ~controllable_BtoR_REQ0 & ~n32425;
  assign n32427 = ~n14784 & ~n32426;
  assign n32428 = ~i_RtoB_ACK0 & ~n32427;
  assign n32429 = ~n20977 & ~n32428;
  assign n32430 = ~controllable_DEQ & ~n32429;
  assign n32431 = ~n20993 & ~n32430;
  assign n32432 = i_FULL & ~n32431;
  assign n32433 = ~n14799 & ~n27814;
  assign n32434 = ~controllable_BtoR_REQ0 & ~n32433;
  assign n32435 = ~n14749 & ~n32434;
  assign n32436 = ~i_RtoB_ACK0 & ~n32435;
  assign n32437 = ~n20977 & ~n32436;
  assign n32438 = ~controllable_DEQ & ~n32437;
  assign n32439 = ~n21003 & ~n32438;
  assign n32440 = ~i_FULL & ~n32439;
  assign n32441 = ~n32432 & ~n32440;
  assign n32442 = ~i_nEMPTY & ~n32441;
  assign n32443 = ~n32424 & ~n32442;
  assign n32444 = controllable_BtoS_ACK0 & ~n32443;
  assign n32445 = ~n18948 & ~n27860;
  assign n32446 = ~controllable_BtoR_REQ0 & ~n32445;
  assign n32447 = ~n28753 & ~n32446;
  assign n32448 = ~i_RtoB_ACK0 & ~n32447;
  assign n32449 = ~n29625 & ~n32448;
  assign n32450 = controllable_DEQ & ~n32449;
  assign n32451 = ~n8885 & ~n20328;
  assign n32452 = ~controllable_BtoR_REQ0 & ~n32451;
  assign n32453 = ~n29437 & ~n32452;
  assign n32454 = ~i_RtoB_ACK0 & ~n32453;
  assign n32455 = ~n29631 & ~n32454;
  assign n32456 = ~controllable_DEQ & ~n32455;
  assign n32457 = ~n32450 & ~n32456;
  assign n32458 = i_FULL & ~n32457;
  assign n32459 = controllable_BtoR_REQ1 & ~n18955;
  assign n32460 = ~n20328 & ~n32459;
  assign n32461 = ~controllable_BtoR_REQ0 & ~n32460;
  assign n32462 = ~n29437 & ~n32461;
  assign n32463 = ~i_RtoB_ACK0 & ~n32462;
  assign n32464 = ~n29631 & ~n32463;
  assign n32465 = ~controllable_DEQ & ~n32464;
  assign n32466 = ~n29641 & ~n32465;
  assign n32467 = ~i_FULL & ~n32466;
  assign n32468 = ~n32458 & ~n32467;
  assign n32469 = i_nEMPTY & ~n32468;
  assign n32470 = ~n8926 & ~n20337;
  assign n32471 = ~controllable_BtoR_REQ0 & ~n32470;
  assign n32472 = ~n29447 & ~n32471;
  assign n32473 = ~i_RtoB_ACK0 & ~n32472;
  assign n32474 = ~n29625 & ~n32473;
  assign n32475 = ~controllable_DEQ & ~n32474;
  assign n32476 = ~n29653 & ~n32475;
  assign n32477 = i_FULL & ~n32476;
  assign n32478 = ~n20347 & ~n27860;
  assign n32479 = ~controllable_BtoR_REQ0 & ~n32478;
  assign n32480 = ~n28753 & ~n32479;
  assign n32481 = ~i_RtoB_ACK0 & ~n32480;
  assign n32482 = ~n29625 & ~n32481;
  assign n32483 = ~controllable_DEQ & ~n32482;
  assign n32484 = ~n29663 & ~n32483;
  assign n32485 = ~i_FULL & ~n32484;
  assign n32486 = ~n32477 & ~n32485;
  assign n32487 = ~i_nEMPTY & ~n32486;
  assign n32488 = ~n32469 & ~n32487;
  assign n32489 = ~controllable_BtoS_ACK0 & ~n32488;
  assign n32490 = ~n32444 & ~n32489;
  assign n32491 = n4465 & ~n32490;
  assign n32492 = ~n18948 & ~n27926;
  assign n32493 = ~controllable_BtoR_REQ0 & ~n32492;
  assign n32494 = ~n28753 & ~n32493;
  assign n32495 = ~i_RtoB_ACK0 & ~n32494;
  assign n32496 = ~n29625 & ~n32495;
  assign n32497 = controllable_DEQ & ~n32496;
  assign n32498 = ~n27219 & ~n29437;
  assign n32499 = ~i_RtoB_ACK0 & ~n32498;
  assign n32500 = ~n29631 & ~n32499;
  assign n32501 = ~controllable_DEQ & ~n32500;
  assign n32502 = ~n32497 & ~n32501;
  assign n32503 = i_FULL & ~n32502;
  assign n32504 = controllable_BtoR_REQ1 & ~n19023;
  assign n32505 = ~n20328 & ~n32504;
  assign n32506 = ~controllable_BtoR_REQ0 & ~n32505;
  assign n32507 = ~n29437 & ~n32506;
  assign n32508 = ~i_RtoB_ACK0 & ~n32507;
  assign n32509 = ~n29631 & ~n32508;
  assign n32510 = ~controllable_DEQ & ~n32509;
  assign n32511 = ~n29641 & ~n32510;
  assign n32512 = ~i_FULL & ~n32511;
  assign n32513 = ~n32503 & ~n32512;
  assign n32514 = i_nEMPTY & ~n32513;
  assign n32515 = ~n27227 & ~n29447;
  assign n32516 = ~i_RtoB_ACK0 & ~n32515;
  assign n32517 = ~n29625 & ~n32516;
  assign n32518 = ~controllable_DEQ & ~n32517;
  assign n32519 = ~n29653 & ~n32518;
  assign n32520 = i_FULL & ~n32519;
  assign n32521 = ~n20347 & ~n27926;
  assign n32522 = ~controllable_BtoR_REQ0 & ~n32521;
  assign n32523 = ~n28753 & ~n32522;
  assign n32524 = ~i_RtoB_ACK0 & ~n32523;
  assign n32525 = ~n29625 & ~n32524;
  assign n32526 = ~controllable_DEQ & ~n32525;
  assign n32527 = ~n29663 & ~n32526;
  assign n32528 = ~i_FULL & ~n32527;
  assign n32529 = ~n32520 & ~n32528;
  assign n32530 = ~i_nEMPTY & ~n32529;
  assign n32531 = ~n32514 & ~n32530;
  assign n32532 = ~controllable_BtoS_ACK0 & ~n32531;
  assign n32533 = ~n21013 & ~n32532;
  assign n32534 = ~n4465 & ~n32533;
  assign n32535 = ~n32491 & ~n32534;
  assign n32536 = i_StoB_REQ10 & ~n32535;
  assign n32537 = ~n11238 & ~n27970;
  assign n32538 = ~controllable_BtoR_REQ0 & ~n32537;
  assign n32539 = ~n17620 & ~n32538;
  assign n32540 = ~i_RtoB_ACK0 & ~n32539;
  assign n32541 = ~n23089 & ~n32540;
  assign n32542 = controllable_DEQ & ~n32541;
  assign n32543 = controllable_BtoR_REQ1 & ~n19394;
  assign n32544 = ~n11248 & ~n32543;
  assign n32545 = ~controllable_BtoR_REQ0 & ~n32544;
  assign n32546 = ~n17635 & ~n32545;
  assign n32547 = ~i_RtoB_ACK0 & ~n32546;
  assign n32548 = ~n23095 & ~n32547;
  assign n32549 = ~controllable_DEQ & ~n32548;
  assign n32550 = ~n32542 & ~n32549;
  assign n32551 = i_FULL & ~n32550;
  assign n32552 = controllable_BtoR_REQ1 & ~n19410;
  assign n32553 = ~n11248 & ~n32552;
  assign n32554 = ~controllable_BtoR_REQ0 & ~n32553;
  assign n32555 = ~n17635 & ~n32554;
  assign n32556 = ~i_RtoB_ACK0 & ~n32555;
  assign n32557 = ~n23095 & ~n32556;
  assign n32558 = ~controllable_DEQ & ~n32557;
  assign n32559 = ~n23093 & ~n32558;
  assign n32560 = ~i_FULL & ~n32559;
  assign n32561 = ~n32551 & ~n32560;
  assign n32562 = i_nEMPTY & ~n32561;
  assign n32563 = controllable_BtoR_REQ1 & ~n19428;
  assign n32564 = ~n11230 & ~n32563;
  assign n32565 = ~controllable_BtoR_REQ0 & ~n32564;
  assign n32566 = ~n17657 & ~n32565;
  assign n32567 = ~i_RtoB_ACK0 & ~n32566;
  assign n32568 = ~n23107 & ~n32567;
  assign n32569 = ~controllable_DEQ & ~n32568;
  assign n32570 = ~n23105 & ~n32569;
  assign n32571 = i_FULL & ~n32570;
  assign n32572 = ~n11284 & ~n27970;
  assign n32573 = ~controllable_BtoR_REQ0 & ~n32572;
  assign n32574 = ~n17620 & ~n32573;
  assign n32575 = ~i_RtoB_ACK0 & ~n32574;
  assign n32576 = ~n23089 & ~n32575;
  assign n32577 = ~controllable_DEQ & ~n32576;
  assign n32578 = ~n23117 & ~n32577;
  assign n32579 = ~i_FULL & ~n32578;
  assign n32580 = ~n32571 & ~n32579;
  assign n32581 = ~i_nEMPTY & ~n32580;
  assign n32582 = ~n32562 & ~n32581;
  assign n32583 = controllable_BtoS_ACK0 & ~n32582;
  assign n32584 = ~n11317 & ~n28015;
  assign n32585 = ~controllable_BtoR_REQ0 & ~n32584;
  assign n32586 = ~n17699 & ~n32585;
  assign n32587 = ~i_RtoB_ACK0 & ~n32586;
  assign n32588 = ~n23129 & ~n32587;
  assign n32589 = controllable_DEQ & ~n32588;
  assign n32590 = controllable_BtoR_REQ1 & ~n19460;
  assign n32591 = ~n11328 & ~n32590;
  assign n32592 = ~controllable_BtoR_REQ0 & ~n32591;
  assign n32593 = ~n17718 & ~n32592;
  assign n32594 = ~i_RtoB_ACK0 & ~n32593;
  assign n32595 = ~n23135 & ~n32594;
  assign n32596 = ~controllable_DEQ & ~n32595;
  assign n32597 = ~n32589 & ~n32596;
  assign n32598 = i_FULL & ~n32597;
  assign n32599 = controllable_BtoR_REQ1 & ~n19476;
  assign n32600 = ~n11328 & ~n32599;
  assign n32601 = ~controllable_BtoR_REQ0 & ~n32600;
  assign n32602 = ~n17718 & ~n32601;
  assign n32603 = ~i_RtoB_ACK0 & ~n32602;
  assign n32604 = ~n23135 & ~n32603;
  assign n32605 = ~controllable_DEQ & ~n32604;
  assign n32606 = ~n23133 & ~n32605;
  assign n32607 = ~i_FULL & ~n32606;
  assign n32608 = ~n32598 & ~n32607;
  assign n32609 = i_nEMPTY & ~n32608;
  assign n32610 = controllable_BtoR_REQ1 & ~n19494;
  assign n32611 = ~n11305 & ~n32610;
  assign n32612 = ~controllable_BtoR_REQ0 & ~n32611;
  assign n32613 = ~n17751 & ~n32612;
  assign n32614 = ~i_RtoB_ACK0 & ~n32613;
  assign n32615 = ~n23147 & ~n32614;
  assign n32616 = ~controllable_DEQ & ~n32615;
  assign n32617 = ~n23145 & ~n32616;
  assign n32618 = i_FULL & ~n32617;
  assign n32619 = ~n11366 & ~n28015;
  assign n32620 = ~controllable_BtoR_REQ0 & ~n32619;
  assign n32621 = ~n17699 & ~n32620;
  assign n32622 = ~i_RtoB_ACK0 & ~n32621;
  assign n32623 = ~n23129 & ~n32622;
  assign n32624 = ~controllable_DEQ & ~n32623;
  assign n32625 = ~n23157 & ~n32624;
  assign n32626 = ~i_FULL & ~n32625;
  assign n32627 = ~n32618 & ~n32626;
  assign n32628 = ~i_nEMPTY & ~n32627;
  assign n32629 = ~n32609 & ~n32628;
  assign n32630 = ~controllable_BtoS_ACK0 & ~n32629;
  assign n32631 = ~n32583 & ~n32630;
  assign n32632 = n4465 & ~n32631;
  assign n32633 = ~n11317 & ~n28062;
  assign n32634 = ~controllable_BtoR_REQ0 & ~n32633;
  assign n32635 = ~n17699 & ~n32634;
  assign n32636 = ~i_RtoB_ACK0 & ~n32635;
  assign n32637 = ~n23129 & ~n32636;
  assign n32638 = controllable_DEQ & ~n32637;
  assign n32639 = controllable_BtoR_REQ1 & ~n19320;
  assign n32640 = ~n11328 & ~n32639;
  assign n32641 = ~controllable_BtoR_REQ0 & ~n32640;
  assign n32642 = ~n17718 & ~n32641;
  assign n32643 = ~i_RtoB_ACK0 & ~n32642;
  assign n32644 = ~n23135 & ~n32643;
  assign n32645 = ~controllable_DEQ & ~n32644;
  assign n32646 = ~n32638 & ~n32645;
  assign n32647 = i_FULL & ~n32646;
  assign n32648 = controllable_BtoR_REQ1 & ~n19334;
  assign n32649 = ~n11328 & ~n32648;
  assign n32650 = ~controllable_BtoR_REQ0 & ~n32649;
  assign n32651 = ~n17718 & ~n32650;
  assign n32652 = ~i_RtoB_ACK0 & ~n32651;
  assign n32653 = ~n23135 & ~n32652;
  assign n32654 = ~controllable_DEQ & ~n32653;
  assign n32655 = ~n23133 & ~n32654;
  assign n32656 = ~i_FULL & ~n32655;
  assign n32657 = ~n32647 & ~n32656;
  assign n32658 = i_nEMPTY & ~n32657;
  assign n32659 = controllable_BtoR_REQ1 & ~n19350;
  assign n32660 = ~n11305 & ~n32659;
  assign n32661 = ~controllable_BtoR_REQ0 & ~n32660;
  assign n32662 = ~n17751 & ~n32661;
  assign n32663 = ~i_RtoB_ACK0 & ~n32662;
  assign n32664 = ~n23147 & ~n32663;
  assign n32665 = ~controllable_DEQ & ~n32664;
  assign n32666 = ~n23145 & ~n32665;
  assign n32667 = i_FULL & ~n32666;
  assign n32668 = ~n11366 & ~n28062;
  assign n32669 = ~controllable_BtoR_REQ0 & ~n32668;
  assign n32670 = ~n17699 & ~n32669;
  assign n32671 = ~i_RtoB_ACK0 & ~n32670;
  assign n32672 = ~n23129 & ~n32671;
  assign n32673 = ~controllable_DEQ & ~n32672;
  assign n32674 = ~n23157 & ~n32673;
  assign n32675 = ~i_FULL & ~n32674;
  assign n32676 = ~n32667 & ~n32675;
  assign n32677 = ~i_nEMPTY & ~n32676;
  assign n32678 = ~n32658 & ~n32677;
  assign n32679 = ~controllable_BtoS_ACK0 & ~n32678;
  assign n32680 = ~n23127 & ~n32679;
  assign n32681 = ~n4465 & ~n32680;
  assign n32682 = ~n32632 & ~n32681;
  assign n32683 = ~i_StoB_REQ10 & ~n32682;
  assign n32684 = ~n32536 & ~n32683;
  assign n32685 = controllable_BtoS_ACK10 & ~n32684;
  assign n32686 = ~n11238 & ~n28116;
  assign n32687 = ~controllable_BtoR_REQ0 & ~n32686;
  assign n32688 = ~n29840 & ~n32687;
  assign n32689 = ~i_RtoB_ACK0 & ~n32688;
  assign n32690 = ~n29825 & ~n32689;
  assign n32691 = controllable_DEQ & ~n32690;
  assign n32692 = ~n29938 & ~n32545;
  assign n32693 = ~i_RtoB_ACK0 & ~n32692;
  assign n32694 = ~n29832 & ~n32693;
  assign n32695 = ~controllable_DEQ & ~n32694;
  assign n32696 = ~n32691 & ~n32695;
  assign n32697 = i_FULL & ~n32696;
  assign n32698 = ~n29938 & ~n32554;
  assign n32699 = ~i_RtoB_ACK0 & ~n32698;
  assign n32700 = ~n29832 & ~n32699;
  assign n32701 = ~controllable_DEQ & ~n32700;
  assign n32702 = ~n29844 & ~n32701;
  assign n32703 = ~i_FULL & ~n32702;
  assign n32704 = ~n32697 & ~n32703;
  assign n32705 = i_nEMPTY & ~n32704;
  assign n32706 = ~n29945 & ~n32565;
  assign n32707 = ~i_RtoB_ACK0 & ~n32706;
  assign n32708 = ~n29860 & ~n32707;
  assign n32709 = ~controllable_DEQ & ~n32708;
  assign n32710 = ~n29858 & ~n32709;
  assign n32711 = i_FULL & ~n32710;
  assign n32712 = ~controllable_DEQ & ~n32690;
  assign n32713 = ~n29872 & ~n32712;
  assign n32714 = ~i_FULL & ~n32713;
  assign n32715 = ~n32711 & ~n32714;
  assign n32716 = ~i_nEMPTY & ~n32715;
  assign n32717 = ~n32705 & ~n32716;
  assign n32718 = controllable_BtoS_ACK0 & ~n32717;
  assign n32719 = ~n11317 & ~n28177;
  assign n32720 = ~controllable_BtoR_REQ0 & ~n32719;
  assign n32721 = ~n29896 & ~n32720;
  assign n32722 = ~i_RtoB_ACK0 & ~n32721;
  assign n32723 = ~n29881 & ~n32722;
  assign n32724 = controllable_DEQ & ~n32723;
  assign n32725 = ~n31230 & ~n32592;
  assign n32726 = ~i_RtoB_ACK0 & ~n32725;
  assign n32727 = ~n29888 & ~n32726;
  assign n32728 = ~controllable_DEQ & ~n32727;
  assign n32729 = ~n32724 & ~n32728;
  assign n32730 = i_FULL & ~n32729;
  assign n32731 = ~n31230 & ~n32601;
  assign n32732 = ~i_RtoB_ACK0 & ~n32731;
  assign n32733 = ~n29888 & ~n32732;
  assign n32734 = ~controllable_DEQ & ~n32733;
  assign n32735 = ~n29900 & ~n32734;
  assign n32736 = ~i_FULL & ~n32735;
  assign n32737 = ~n32730 & ~n32736;
  assign n32738 = i_nEMPTY & ~n32737;
  assign n32739 = ~n31245 & ~n32612;
  assign n32740 = ~i_RtoB_ACK0 & ~n32739;
  assign n32741 = ~n29916 & ~n32740;
  assign n32742 = ~controllable_DEQ & ~n32741;
  assign n32743 = ~n29914 & ~n32742;
  assign n32744 = i_FULL & ~n32743;
  assign n32745 = ~controllable_DEQ & ~n32723;
  assign n32746 = ~n29928 & ~n32745;
  assign n32747 = ~i_FULL & ~n32746;
  assign n32748 = ~n32744 & ~n32747;
  assign n32749 = ~i_nEMPTY & ~n32748;
  assign n32750 = ~n32738 & ~n32749;
  assign n32751 = ~controllable_BtoS_ACK0 & ~n32750;
  assign n32752 = ~n32718 & ~n32751;
  assign n32753 = n4465 & ~n32752;
  assign n32754 = ~n11317 & ~n28250;
  assign n32755 = ~controllable_BtoR_REQ0 & ~n32754;
  assign n32756 = ~n29896 & ~n32755;
  assign n32757 = ~i_RtoB_ACK0 & ~n32756;
  assign n32758 = ~n29881 & ~n32757;
  assign n32759 = controllable_DEQ & ~n32758;
  assign n32760 = ~n31230 & ~n32641;
  assign n32761 = ~i_RtoB_ACK0 & ~n32760;
  assign n32762 = ~n29888 & ~n32761;
  assign n32763 = ~controllable_DEQ & ~n32762;
  assign n32764 = ~n32759 & ~n32763;
  assign n32765 = i_FULL & ~n32764;
  assign n32766 = ~n31230 & ~n32650;
  assign n32767 = ~i_RtoB_ACK0 & ~n32766;
  assign n32768 = ~n29888 & ~n32767;
  assign n32769 = ~controllable_DEQ & ~n32768;
  assign n32770 = ~n29900 & ~n32769;
  assign n32771 = ~i_FULL & ~n32770;
  assign n32772 = ~n32765 & ~n32771;
  assign n32773 = i_nEMPTY & ~n32772;
  assign n32774 = ~n31245 & ~n32661;
  assign n32775 = ~i_RtoB_ACK0 & ~n32774;
  assign n32776 = ~n29916 & ~n32775;
  assign n32777 = ~controllable_DEQ & ~n32776;
  assign n32778 = ~n29914 & ~n32777;
  assign n32779 = i_FULL & ~n32778;
  assign n32780 = ~controllable_DEQ & ~n32758;
  assign n32781 = ~n29928 & ~n32780;
  assign n32782 = ~i_FULL & ~n32781;
  assign n32783 = ~n32779 & ~n32782;
  assign n32784 = ~i_nEMPTY & ~n32783;
  assign n32785 = ~n32773 & ~n32784;
  assign n32786 = ~controllable_BtoS_ACK0 & ~n32785;
  assign n32787 = ~n29958 & ~n32786;
  assign n32788 = ~n4465 & ~n32787;
  assign n32789 = ~n32753 & ~n32788;
  assign n32790 = i_StoB_REQ10 & ~n32789;
  assign n32791 = ~n32683 & ~n32790;
  assign n32792 = ~controllable_BtoS_ACK10 & ~n32791;
  assign n32793 = ~n32685 & ~n32792;
  assign n32794 = n4464 & ~n32793;
  assign n32795 = ~n5245 & ~n28286;
  assign n32796 = ~controllable_BtoR_REQ0 & ~n32795;
  assign n32797 = ~n14749 & ~n32796;
  assign n32798 = ~i_RtoB_ACK0 & ~n32797;
  assign n32799 = ~n20977 & ~n32798;
  assign n32800 = controllable_DEQ & ~n32799;
  assign n32801 = ~n14765 & ~n27477;
  assign n32802 = ~i_RtoB_ACK0 & ~n32801;
  assign n32803 = ~n20983 & ~n32802;
  assign n32804 = ~controllable_DEQ & ~n32803;
  assign n32805 = ~n32800 & ~n32804;
  assign n32806 = i_FULL & ~n32805;
  assign n32807 = controllable_BtoR_REQ1 & ~n19633;
  assign n32808 = ~n5255 & ~n32807;
  assign n32809 = ~controllable_BtoR_REQ0 & ~n32808;
  assign n32810 = ~n14765 & ~n32809;
  assign n32811 = ~i_RtoB_ACK0 & ~n32810;
  assign n32812 = ~n20983 & ~n32811;
  assign n32813 = ~controllable_DEQ & ~n32812;
  assign n32814 = ~n20981 & ~n32813;
  assign n32815 = ~i_FULL & ~n32814;
  assign n32816 = ~n32806 & ~n32815;
  assign n32817 = i_nEMPTY & ~n32816;
  assign n32818 = ~n14784 & ~n27485;
  assign n32819 = ~i_RtoB_ACK0 & ~n32818;
  assign n32820 = ~n20977 & ~n32819;
  assign n32821 = ~controllable_DEQ & ~n32820;
  assign n32822 = ~n20993 & ~n32821;
  assign n32823 = i_FULL & ~n32822;
  assign n32824 = ~n14799 & ~n28286;
  assign n32825 = ~controllable_BtoR_REQ0 & ~n32824;
  assign n32826 = ~n14749 & ~n32825;
  assign n32827 = ~i_RtoB_ACK0 & ~n32826;
  assign n32828 = ~n20977 & ~n32827;
  assign n32829 = ~controllable_DEQ & ~n32828;
  assign n32830 = ~n21003 & ~n32829;
  assign n32831 = ~i_FULL & ~n32830;
  assign n32832 = ~n32823 & ~n32831;
  assign n32833 = ~i_nEMPTY & ~n32832;
  assign n32834 = ~n32817 & ~n32833;
  assign n32835 = controllable_BtoS_ACK0 & ~n32834;
  assign n32836 = ~n18948 & ~n28325;
  assign n32837 = ~controllable_BtoR_REQ0 & ~n32836;
  assign n32838 = ~n28753 & ~n32837;
  assign n32839 = ~i_RtoB_ACK0 & ~n32838;
  assign n32840 = ~n29625 & ~n32839;
  assign n32841 = controllable_DEQ & ~n32840;
  assign n32842 = ~n27505 & ~n29437;
  assign n32843 = ~i_RtoB_ACK0 & ~n32842;
  assign n32844 = ~n29631 & ~n32843;
  assign n32845 = ~controllable_DEQ & ~n32844;
  assign n32846 = ~n32841 & ~n32845;
  assign n32847 = i_FULL & ~n32846;
  assign n32848 = controllable_BtoR_REQ1 & ~n19697;
  assign n32849 = ~n20328 & ~n32848;
  assign n32850 = ~controllable_BtoR_REQ0 & ~n32849;
  assign n32851 = ~n29437 & ~n32850;
  assign n32852 = ~i_RtoB_ACK0 & ~n32851;
  assign n32853 = ~n29631 & ~n32852;
  assign n32854 = ~controllable_DEQ & ~n32853;
  assign n32855 = ~n29641 & ~n32854;
  assign n32856 = ~i_FULL & ~n32855;
  assign n32857 = ~n32847 & ~n32856;
  assign n32858 = i_nEMPTY & ~n32857;
  assign n32859 = ~n27513 & ~n29447;
  assign n32860 = ~i_RtoB_ACK0 & ~n32859;
  assign n32861 = ~n29625 & ~n32860;
  assign n32862 = ~controllable_DEQ & ~n32861;
  assign n32863 = ~n29653 & ~n32862;
  assign n32864 = i_FULL & ~n32863;
  assign n32865 = ~n20347 & ~n28325;
  assign n32866 = ~controllable_BtoR_REQ0 & ~n32865;
  assign n32867 = ~n28753 & ~n32866;
  assign n32868 = ~i_RtoB_ACK0 & ~n32867;
  assign n32869 = ~n29625 & ~n32868;
  assign n32870 = ~controllable_DEQ & ~n32869;
  assign n32871 = ~n29663 & ~n32870;
  assign n32872 = ~i_FULL & ~n32871;
  assign n32873 = ~n32864 & ~n32872;
  assign n32874 = ~i_nEMPTY & ~n32873;
  assign n32875 = ~n32858 & ~n32874;
  assign n32876 = ~controllable_BtoS_ACK0 & ~n32875;
  assign n32877 = ~n32835 & ~n32876;
  assign n32878 = n4465 & ~n32877;
  assign n32879 = ~n21013 & ~n32876;
  assign n32880 = ~n4465 & ~n32879;
  assign n32881 = ~n32878 & ~n32880;
  assign n32882 = i_StoB_REQ10 & ~n32881;
  assign n32883 = ~n11238 & ~n28371;
  assign n32884 = ~controllable_BtoR_REQ0 & ~n32883;
  assign n32885 = ~n17620 & ~n32884;
  assign n32886 = ~i_RtoB_ACK0 & ~n32885;
  assign n32887 = ~n23089 & ~n32886;
  assign n32888 = controllable_DEQ & ~n32887;
  assign n32889 = controllable_BtoR_REQ1 & ~n20012;
  assign n32890 = ~n11248 & ~n32889;
  assign n32891 = ~controllable_BtoR_REQ0 & ~n32890;
  assign n32892 = ~n17635 & ~n32891;
  assign n32893 = ~i_RtoB_ACK0 & ~n32892;
  assign n32894 = ~n23095 & ~n32893;
  assign n32895 = ~controllable_DEQ & ~n32894;
  assign n32896 = ~n32888 & ~n32895;
  assign n32897 = i_FULL & ~n32896;
  assign n32898 = controllable_BtoR_REQ1 & ~n20028;
  assign n32899 = ~n11248 & ~n32898;
  assign n32900 = ~controllable_BtoR_REQ0 & ~n32899;
  assign n32901 = ~n17635 & ~n32900;
  assign n32902 = ~i_RtoB_ACK0 & ~n32901;
  assign n32903 = ~n23095 & ~n32902;
  assign n32904 = ~controllable_DEQ & ~n32903;
  assign n32905 = ~n23093 & ~n32904;
  assign n32906 = ~i_FULL & ~n32905;
  assign n32907 = ~n32897 & ~n32906;
  assign n32908 = i_nEMPTY & ~n32907;
  assign n32909 = controllable_BtoR_REQ1 & ~n20046;
  assign n32910 = ~n11230 & ~n32909;
  assign n32911 = ~controllable_BtoR_REQ0 & ~n32910;
  assign n32912 = ~n17657 & ~n32911;
  assign n32913 = ~i_RtoB_ACK0 & ~n32912;
  assign n32914 = ~n23107 & ~n32913;
  assign n32915 = ~controllable_DEQ & ~n32914;
  assign n32916 = ~n23105 & ~n32915;
  assign n32917 = i_FULL & ~n32916;
  assign n32918 = ~n11284 & ~n28371;
  assign n32919 = ~controllable_BtoR_REQ0 & ~n32918;
  assign n32920 = ~n17620 & ~n32919;
  assign n32921 = ~i_RtoB_ACK0 & ~n32920;
  assign n32922 = ~n23089 & ~n32921;
  assign n32923 = ~controllable_DEQ & ~n32922;
  assign n32924 = ~n23117 & ~n32923;
  assign n32925 = ~i_FULL & ~n32924;
  assign n32926 = ~n32917 & ~n32925;
  assign n32927 = ~i_nEMPTY & ~n32926;
  assign n32928 = ~n32908 & ~n32927;
  assign n32929 = controllable_BtoS_ACK0 & ~n32928;
  assign n32930 = ~n11317 & ~n28414;
  assign n32931 = ~controllable_BtoR_REQ0 & ~n32930;
  assign n32932 = ~n17699 & ~n32931;
  assign n32933 = ~i_RtoB_ACK0 & ~n32932;
  assign n32934 = ~n23129 & ~n32933;
  assign n32935 = controllable_DEQ & ~n32934;
  assign n32936 = controllable_BtoR_REQ1 & ~n19938;
  assign n32937 = ~n11328 & ~n32936;
  assign n32938 = ~controllable_BtoR_REQ0 & ~n32937;
  assign n32939 = ~n17718 & ~n32938;
  assign n32940 = ~i_RtoB_ACK0 & ~n32939;
  assign n32941 = ~n23135 & ~n32940;
  assign n32942 = ~controllable_DEQ & ~n32941;
  assign n32943 = ~n32935 & ~n32942;
  assign n32944 = i_FULL & ~n32943;
  assign n32945 = controllable_BtoR_REQ1 & ~n19952;
  assign n32946 = ~n11328 & ~n32945;
  assign n32947 = ~controllable_BtoR_REQ0 & ~n32946;
  assign n32948 = ~n17718 & ~n32947;
  assign n32949 = ~i_RtoB_ACK0 & ~n32948;
  assign n32950 = ~n23135 & ~n32949;
  assign n32951 = ~controllable_DEQ & ~n32950;
  assign n32952 = ~n23133 & ~n32951;
  assign n32953 = ~i_FULL & ~n32952;
  assign n32954 = ~n32944 & ~n32953;
  assign n32955 = i_nEMPTY & ~n32954;
  assign n32956 = controllable_BtoR_REQ1 & ~n19968;
  assign n32957 = ~n11305 & ~n32956;
  assign n32958 = ~controllable_BtoR_REQ0 & ~n32957;
  assign n32959 = ~n17751 & ~n32958;
  assign n32960 = ~i_RtoB_ACK0 & ~n32959;
  assign n32961 = ~n23147 & ~n32960;
  assign n32962 = ~controllable_DEQ & ~n32961;
  assign n32963 = ~n23145 & ~n32962;
  assign n32964 = i_FULL & ~n32963;
  assign n32965 = ~n11366 & ~n28414;
  assign n32966 = ~controllable_BtoR_REQ0 & ~n32965;
  assign n32967 = ~n17699 & ~n32966;
  assign n32968 = ~i_RtoB_ACK0 & ~n32967;
  assign n32969 = ~n23129 & ~n32968;
  assign n32970 = ~controllable_DEQ & ~n32969;
  assign n32971 = ~n23157 & ~n32970;
  assign n32972 = ~i_FULL & ~n32971;
  assign n32973 = ~n32964 & ~n32972;
  assign n32974 = ~i_nEMPTY & ~n32973;
  assign n32975 = ~n32955 & ~n32974;
  assign n32976 = ~controllable_BtoS_ACK0 & ~n32975;
  assign n32977 = ~n32929 & ~n32976;
  assign n32978 = n4465 & ~n32977;
  assign n32979 = ~n23127 & ~n32976;
  assign n32980 = ~n4465 & ~n32979;
  assign n32981 = ~n32978 & ~n32980;
  assign n32982 = ~i_StoB_REQ10 & ~n32981;
  assign n32983 = ~n32882 & ~n32982;
  assign n32984 = controllable_BtoS_ACK10 & ~n32983;
  assign n32985 = ~n11238 & ~n28465;
  assign n32986 = ~controllable_BtoR_REQ0 & ~n32985;
  assign n32987 = ~n29840 & ~n32986;
  assign n32988 = ~i_RtoB_ACK0 & ~n32987;
  assign n32989 = ~n29825 & ~n32988;
  assign n32990 = controllable_DEQ & ~n32989;
  assign n32991 = ~n29938 & ~n32891;
  assign n32992 = ~i_RtoB_ACK0 & ~n32991;
  assign n32993 = ~n29832 & ~n32992;
  assign n32994 = ~controllable_DEQ & ~n32993;
  assign n32995 = ~n32990 & ~n32994;
  assign n32996 = i_FULL & ~n32995;
  assign n32997 = ~n29938 & ~n32900;
  assign n32998 = ~i_RtoB_ACK0 & ~n32997;
  assign n32999 = ~n29832 & ~n32998;
  assign n33000 = ~controllable_DEQ & ~n32999;
  assign n33001 = ~n29844 & ~n33000;
  assign n33002 = ~i_FULL & ~n33001;
  assign n33003 = ~n32996 & ~n33002;
  assign n33004 = i_nEMPTY & ~n33003;
  assign n33005 = ~n29945 & ~n32911;
  assign n33006 = ~i_RtoB_ACK0 & ~n33005;
  assign n33007 = ~n29860 & ~n33006;
  assign n33008 = ~controllable_DEQ & ~n33007;
  assign n33009 = ~n29858 & ~n33008;
  assign n33010 = i_FULL & ~n33009;
  assign n33011 = ~controllable_DEQ & ~n32989;
  assign n33012 = ~n29872 & ~n33011;
  assign n33013 = ~i_FULL & ~n33012;
  assign n33014 = ~n33010 & ~n33013;
  assign n33015 = ~i_nEMPTY & ~n33014;
  assign n33016 = ~n33004 & ~n33015;
  assign n33017 = controllable_BtoS_ACK0 & ~n33016;
  assign n33018 = ~n11317 & ~n28494;
  assign n33019 = ~controllable_BtoR_REQ0 & ~n33018;
  assign n33020 = ~n29896 & ~n33019;
  assign n33021 = ~i_RtoB_ACK0 & ~n33020;
  assign n33022 = ~n29881 & ~n33021;
  assign n33023 = controllable_DEQ & ~n33022;
  assign n33024 = ~n31230 & ~n32938;
  assign n33025 = ~i_RtoB_ACK0 & ~n33024;
  assign n33026 = ~n29888 & ~n33025;
  assign n33027 = ~controllable_DEQ & ~n33026;
  assign n33028 = ~n33023 & ~n33027;
  assign n33029 = i_FULL & ~n33028;
  assign n33030 = ~n31230 & ~n32947;
  assign n33031 = ~i_RtoB_ACK0 & ~n33030;
  assign n33032 = ~n29888 & ~n33031;
  assign n33033 = ~controllable_DEQ & ~n33032;
  assign n33034 = ~n29900 & ~n33033;
  assign n33035 = ~i_FULL & ~n33034;
  assign n33036 = ~n33029 & ~n33035;
  assign n33037 = i_nEMPTY & ~n33036;
  assign n33038 = ~n31245 & ~n32958;
  assign n33039 = ~i_RtoB_ACK0 & ~n33038;
  assign n33040 = ~n29916 & ~n33039;
  assign n33041 = ~controllable_DEQ & ~n33040;
  assign n33042 = ~n29914 & ~n33041;
  assign n33043 = i_FULL & ~n33042;
  assign n33044 = ~controllable_DEQ & ~n33022;
  assign n33045 = ~n29928 & ~n33044;
  assign n33046 = ~i_FULL & ~n33045;
  assign n33047 = ~n33043 & ~n33046;
  assign n33048 = ~i_nEMPTY & ~n33047;
  assign n33049 = ~n33037 & ~n33048;
  assign n33050 = ~controllable_BtoS_ACK0 & ~n33049;
  assign n33051 = ~n33017 & ~n33050;
  assign n33052 = n4465 & ~n33051;
  assign n33053 = ~n29958 & ~n33050;
  assign n33054 = ~n4465 & ~n33053;
  assign n33055 = ~n33052 & ~n33054;
  assign n33056 = i_StoB_REQ10 & ~n33055;
  assign n33057 = ~n32982 & ~n33056;
  assign n33058 = ~controllable_BtoS_ACK10 & ~n33057;
  assign n33059 = ~n32984 & ~n33058;
  assign n33060 = ~n4464 & ~n33059;
  assign n33061 = ~n32794 & ~n33060;
  assign n33062 = n4463 & ~n33061;
  assign n33063 = ~n31548 & ~n33062;
  assign n33064 = n4462 & ~n33063;
  assign n33065 = ~n11238 & ~n28587;
  assign n33066 = ~controllable_BtoR_REQ0 & ~n33065;
  assign n33067 = ~n29840 & ~n33066;
  assign n33068 = ~i_RtoB_ACK0 & ~n33067;
  assign n33069 = ~n29825 & ~n33068;
  assign n33070 = controllable_DEQ & ~n33069;
  assign n33071 = controllable_BtoR_REQ1 & ~n20376;
  assign n33072 = ~n11248 & ~n33071;
  assign n33073 = ~controllable_BtoR_REQ0 & ~n33072;
  assign n33074 = ~n29938 & ~n33073;
  assign n33075 = ~i_RtoB_ACK0 & ~n33074;
  assign n33076 = ~n29832 & ~n33075;
  assign n33077 = ~controllable_DEQ & ~n33076;
  assign n33078 = ~n33070 & ~n33077;
  assign n33079 = i_FULL & ~n33078;
  assign n33080 = controllable_BtoR_REQ1 & ~n20392;
  assign n33081 = ~n11248 & ~n33080;
  assign n33082 = ~controllable_BtoR_REQ0 & ~n33081;
  assign n33083 = ~n29938 & ~n33082;
  assign n33084 = ~i_RtoB_ACK0 & ~n33083;
  assign n33085 = ~n29832 & ~n33084;
  assign n33086 = ~controllable_DEQ & ~n33085;
  assign n33087 = ~n29844 & ~n33086;
  assign n33088 = ~i_FULL & ~n33087;
  assign n33089 = ~n33079 & ~n33088;
  assign n33090 = i_nEMPTY & ~n33089;
  assign n33091 = controllable_BtoR_REQ1 & ~n20410;
  assign n33092 = ~n11230 & ~n33091;
  assign n33093 = ~controllable_BtoR_REQ0 & ~n33092;
  assign n33094 = ~n29945 & ~n33093;
  assign n33095 = ~i_RtoB_ACK0 & ~n33094;
  assign n33096 = ~n29860 & ~n33095;
  assign n33097 = ~controllable_DEQ & ~n33096;
  assign n33098 = ~n29858 & ~n33097;
  assign n33099 = i_FULL & ~n33098;
  assign n33100 = ~controllable_DEQ & ~n33069;
  assign n33101 = ~n29872 & ~n33100;
  assign n33102 = ~i_FULL & ~n33101;
  assign n33103 = ~n33099 & ~n33102;
  assign n33104 = ~i_nEMPTY & ~n33103;
  assign n33105 = ~n33090 & ~n33104;
  assign n33106 = controllable_BtoS_ACK0 & ~n33105;
  assign n33107 = ~n32786 & ~n33106;
  assign n33108 = n4465 & ~n33107;
  assign n33109 = ~n32788 & ~n33108;
  assign n33110 = i_StoB_REQ10 & ~n33109;
  assign n33111 = ~n11238 & ~n28629;
  assign n33112 = ~controllable_BtoR_REQ0 & ~n33111;
  assign n33113 = ~n17620 & ~n33112;
  assign n33114 = ~i_RtoB_ACK0 & ~n33113;
  assign n33115 = ~n23089 & ~n33114;
  assign n33116 = controllable_DEQ & ~n33115;
  assign n33117 = ~n17635 & ~n33073;
  assign n33118 = ~i_RtoB_ACK0 & ~n33117;
  assign n33119 = ~n23095 & ~n33118;
  assign n33120 = ~controllable_DEQ & ~n33119;
  assign n33121 = ~n33116 & ~n33120;
  assign n33122 = i_FULL & ~n33121;
  assign n33123 = ~n17635 & ~n33082;
  assign n33124 = ~i_RtoB_ACK0 & ~n33123;
  assign n33125 = ~n23095 & ~n33124;
  assign n33126 = ~controllable_DEQ & ~n33125;
  assign n33127 = ~n23093 & ~n33126;
  assign n33128 = ~i_FULL & ~n33127;
  assign n33129 = ~n33122 & ~n33128;
  assign n33130 = i_nEMPTY & ~n33129;
  assign n33131 = ~n17657 & ~n33093;
  assign n33132 = ~i_RtoB_ACK0 & ~n33131;
  assign n33133 = ~n23107 & ~n33132;
  assign n33134 = ~controllable_DEQ & ~n33133;
  assign n33135 = ~n23105 & ~n33134;
  assign n33136 = i_FULL & ~n33135;
  assign n33137 = ~n11284 & ~n28629;
  assign n33138 = ~controllable_BtoR_REQ0 & ~n33137;
  assign n33139 = ~n17620 & ~n33138;
  assign n33140 = ~i_RtoB_ACK0 & ~n33139;
  assign n33141 = ~n23089 & ~n33140;
  assign n33142 = ~controllable_DEQ & ~n33141;
  assign n33143 = ~n23117 & ~n33142;
  assign n33144 = ~i_FULL & ~n33143;
  assign n33145 = ~n33136 & ~n33144;
  assign n33146 = ~i_nEMPTY & ~n33145;
  assign n33147 = ~n33130 & ~n33146;
  assign n33148 = controllable_BtoS_ACK0 & ~n33147;
  assign n33149 = ~n32679 & ~n33148;
  assign n33150 = n4465 & ~n33149;
  assign n33151 = ~n32681 & ~n33150;
  assign n33152 = ~i_StoB_REQ10 & ~n33151;
  assign n33153 = ~n33110 & ~n33152;
  assign n33154 = ~controllable_BtoS_ACK10 & ~n33153;
  assign n33155 = ~n30806 & ~n33154;
  assign n33156 = n4464 & ~n33155;
  assign n33157 = ~n30806 & ~n33058;
  assign n33158 = ~n4464 & ~n33157;
  assign n33159 = ~n33156 & ~n33158;
  assign n33160 = n4463 & ~n33159;
  assign n33161 = ~n31548 & ~n33160;
  assign n33162 = ~n4462 & ~n33161;
  assign n33163 = ~n33064 & ~n33162;
  assign n33164 = ~n4461 & ~n33163;
  assign n33165 = ~n32399 & ~n33164;
  assign n33166 = n4459 & ~n33165;
  assign n33167 = ~n31637 & ~n33166;
  assign n33168 = ~n4455 & ~n33167;
  assign n33169 = ~n29589 & ~n33168;
  assign n33170 = ~n4445 & ~n33169;
  assign n33171 = ~n27813 & ~n33170;
  assign n33172 = n4442 & ~n33171;
  assign n33173 = ~n4459 & ~n28582;
  assign n33174 = n4459 & ~n29584;
  assign n33175 = ~n33173 & ~n33174;
  assign n33176 = n4455 & ~n33175;
  assign n33177 = ~n4455 & ~n31547;
  assign n33178 = ~n33176 & ~n33177;
  assign n33179 = ~n4442 & ~n33178;
  assign n33180 = ~n33172 & ~n33179;
  assign n33181 = ~n4438 & ~n33180;
  assign n33182 = ~n4438 & ~n33181;
  assign n33183 = n4386 & ~n33182;
  assign n33184 = ~controllable_DEQ & ~n5045;
  assign n33185 = ~n5091 & ~n33184;
  assign n33186 = ~i_FULL & ~n33185;
  assign n33187 = ~n5083 & ~n33186;
  assign n33188 = ~i_nEMPTY & ~n33187;
  assign n33189 = ~n5061 & ~n33188;
  assign n33190 = controllable_BtoS_ACK0 & ~n33189;
  assign n33191 = ~controllable_DEQ & ~n5142;
  assign n33192 = ~n5188 & ~n33191;
  assign n33193 = ~i_FULL & ~n33192;
  assign n33194 = ~n5180 & ~n33193;
  assign n33195 = ~i_nEMPTY & ~n33194;
  assign n33196 = ~n5158 & ~n33195;
  assign n33197 = ~controllable_BtoS_ACK0 & ~n33196;
  assign n33198 = ~n33190 & ~n33197;
  assign n33199 = n4465 & ~n33198;
  assign n33200 = ~controllable_DEQ & ~n5250;
  assign n33201 = ~n5296 & ~n33200;
  assign n33202 = ~i_FULL & ~n33201;
  assign n33203 = ~n5288 & ~n33202;
  assign n33204 = ~i_nEMPTY & ~n33203;
  assign n33205 = ~n5266 & ~n33204;
  assign n33206 = controllable_BtoS_ACK0 & ~n33205;
  assign n33207 = ~controllable_DEQ & ~n5356;
  assign n33208 = ~n5402 & ~n33207;
  assign n33209 = ~i_FULL & ~n33208;
  assign n33210 = ~n5394 & ~n33209;
  assign n33211 = ~i_nEMPTY & ~n33210;
  assign n33212 = ~n5372 & ~n33211;
  assign n33213 = ~controllable_BtoS_ACK0 & ~n33212;
  assign n33214 = ~n33206 & ~n33213;
  assign n33215 = ~n4465 & ~n33214;
  assign n33216 = ~n33199 & ~n33215;
  assign n33217 = i_StoB_REQ10 & ~n33216;
  assign n33218 = ~controllable_DEQ & ~n6783;
  assign n33219 = ~n6871 & ~n33218;
  assign n33220 = ~i_FULL & ~n33219;
  assign n33221 = ~n6863 & ~n33220;
  assign n33222 = ~i_nEMPTY & ~n33221;
  assign n33223 = ~n6834 & ~n33222;
  assign n33224 = controllable_BtoS_ACK0 & ~n33223;
  assign n33225 = ~controllable_DEQ & ~n6949;
  assign n33226 = ~n7037 & ~n33225;
  assign n33227 = ~i_FULL & ~n33226;
  assign n33228 = ~n7029 & ~n33227;
  assign n33229 = ~i_nEMPTY & ~n33228;
  assign n33230 = ~n7000 & ~n33229;
  assign n33231 = ~controllable_BtoS_ACK0 & ~n33230;
  assign n33232 = ~n33224 & ~n33231;
  assign n33233 = n4465 & ~n33232;
  assign n33234 = ~controllable_DEQ & ~n7109;
  assign n33235 = ~n7157 & ~n33234;
  assign n33236 = ~i_FULL & ~n33235;
  assign n33237 = ~n7149 & ~n33236;
  assign n33238 = ~i_nEMPTY & ~n33237;
  assign n33239 = ~n7126 & ~n33238;
  assign n33240 = controllable_BtoS_ACK0 & ~n33239;
  assign n33241 = ~controllable_DEQ & ~n7275;
  assign n33242 = ~n7363 & ~n33241;
  assign n33243 = ~i_FULL & ~n33242;
  assign n33244 = ~n7355 & ~n33243;
  assign n33245 = ~i_nEMPTY & ~n33244;
  assign n33246 = ~n7326 & ~n33245;
  assign n33247 = ~controllable_BtoS_ACK0 & ~n33246;
  assign n33248 = ~n33240 & ~n33247;
  assign n33249 = ~n4465 & ~n33248;
  assign n33250 = ~n33233 & ~n33249;
  assign n33251 = ~i_StoB_REQ10 & ~n33250;
  assign n33252 = ~n33217 & ~n33251;
  assign n33253 = controllable_BtoS_ACK10 & ~n33252;
  assign n33254 = ~n7683 & ~n33251;
  assign n33255 = ~controllable_BtoS_ACK10 & ~n33254;
  assign n33256 = ~n33253 & ~n33255;
  assign n33257 = n4464 & ~n33256;
  assign n33258 = ~controllable_DEQ & ~n7723;
  assign n33259 = ~n7769 & ~n33258;
  assign n33260 = ~i_FULL & ~n33259;
  assign n33261 = ~n7761 & ~n33260;
  assign n33262 = ~i_nEMPTY & ~n33261;
  assign n33263 = ~n7739 & ~n33262;
  assign n33264 = controllable_BtoS_ACK0 & ~n33263;
  assign n33265 = ~controllable_DEQ & ~n7815;
  assign n33266 = ~n7861 & ~n33265;
  assign n33267 = ~i_FULL & ~n33266;
  assign n33268 = ~n7853 & ~n33267;
  assign n33269 = ~i_nEMPTY & ~n33268;
  assign n33270 = ~n7831 & ~n33269;
  assign n33271 = ~controllable_BtoS_ACK0 & ~n33270;
  assign n33272 = ~n33264 & ~n33271;
  assign n33273 = n4465 & ~n33272;
  assign n33274 = ~n33206 & ~n33271;
  assign n33275 = ~n4465 & ~n33274;
  assign n33276 = ~n33273 & ~n33275;
  assign n33277 = i_StoB_REQ10 & ~n33276;
  assign n33278 = ~controllable_DEQ & ~n7945;
  assign n33279 = ~n8033 & ~n33278;
  assign n33280 = ~i_FULL & ~n33279;
  assign n33281 = ~n8025 & ~n33280;
  assign n33282 = ~i_nEMPTY & ~n33281;
  assign n33283 = ~n7996 & ~n33282;
  assign n33284 = controllable_BtoS_ACK0 & ~n33283;
  assign n33285 = ~controllable_DEQ & ~n8109;
  assign n33286 = ~n8197 & ~n33285;
  assign n33287 = ~i_FULL & ~n33286;
  assign n33288 = ~n8189 & ~n33287;
  assign n33289 = ~i_nEMPTY & ~n33288;
  assign n33290 = ~n8160 & ~n33289;
  assign n33291 = ~controllable_BtoS_ACK0 & ~n33290;
  assign n33292 = ~n33284 & ~n33291;
  assign n33293 = n4465 & ~n33292;
  assign n33294 = ~controllable_DEQ & ~n8247;
  assign n33295 = ~n8293 & ~n33294;
  assign n33296 = ~i_FULL & ~n33295;
  assign n33297 = ~n8285 & ~n33296;
  assign n33298 = ~i_nEMPTY & ~n33297;
  assign n33299 = ~n8263 & ~n33298;
  assign n33300 = controllable_BtoS_ACK0 & ~n33299;
  assign n33301 = ~controllable_DEQ & ~n8350;
  assign n33302 = ~n8433 & ~n33301;
  assign n33303 = ~i_FULL & ~n33302;
  assign n33304 = ~n8425 & ~n33303;
  assign n33305 = ~i_nEMPTY & ~n33304;
  assign n33306 = ~n8399 & ~n33305;
  assign n33307 = ~controllable_BtoS_ACK0 & ~n33306;
  assign n33308 = ~n33300 & ~n33307;
  assign n33309 = ~n4465 & ~n33308;
  assign n33310 = ~n33293 & ~n33309;
  assign n33311 = ~i_StoB_REQ10 & ~n33310;
  assign n33312 = ~n33277 & ~n33311;
  assign n33313 = controllable_BtoS_ACK10 & ~n33312;
  assign n33314 = ~n8748 & ~n33311;
  assign n33315 = ~controllable_BtoS_ACK10 & ~n33314;
  assign n33316 = ~n33313 & ~n33315;
  assign n33317 = ~n4464 & ~n33316;
  assign n33318 = ~n33257 & ~n33317;
  assign n33319 = n4463 & ~n33318;
  assign n33320 = ~controllable_DEQ & ~n8772;
  assign n33321 = ~n8833 & ~n33320;
  assign n33322 = ~i_FULL & ~n33321;
  assign n33323 = ~n8827 & ~n33322;
  assign n33324 = ~i_nEMPTY & ~n33323;
  assign n33325 = ~n8810 & ~n33324;
  assign n33326 = controllable_BtoS_ACK0 & ~n33325;
  assign n33327 = ~controllable_DEQ & ~n8873;
  assign n33328 = ~n8942 & ~n33327;
  assign n33329 = ~i_FULL & ~n33328;
  assign n33330 = ~n8934 & ~n33329;
  assign n33331 = ~i_nEMPTY & ~n33330;
  assign n33332 = ~n8913 & ~n33331;
  assign n33333 = ~controllable_BtoS_ACK0 & ~n33332;
  assign n33334 = ~n33326 & ~n33333;
  assign n33335 = n4465 & ~n33334;
  assign n33336 = ~controllable_DEQ & ~n8981;
  assign n33337 = ~n9042 & ~n33336;
  assign n33338 = ~i_FULL & ~n33337;
  assign n33339 = ~n9036 & ~n33338;
  assign n33340 = ~i_nEMPTY & ~n33339;
  assign n33341 = ~n9019 & ~n33340;
  assign n33342 = ~controllable_BtoS_ACK0 & ~n33341;
  assign n33343 = ~n33206 & ~n33342;
  assign n33344 = ~n4465 & ~n33343;
  assign n33345 = ~n33335 & ~n33344;
  assign n33346 = i_StoB_REQ10 & ~n33345;
  assign n33347 = ~controllable_DEQ & ~n9508;
  assign n33348 = ~n9593 & ~n33347;
  assign n33349 = ~i_FULL & ~n33348;
  assign n33350 = ~n9585 & ~n33349;
  assign n33351 = ~i_nEMPTY & ~n33350;
  assign n33352 = ~n9559 & ~n33351;
  assign n33353 = controllable_BtoS_ACK0 & ~n33352;
  assign n33354 = ~controllable_DEQ & ~n9655;
  assign n33355 = ~n9740 & ~n33354;
  assign n33356 = ~i_FULL & ~n33355;
  assign n33357 = ~n9732 & ~n33356;
  assign n33358 = ~i_nEMPTY & ~n33357;
  assign n33359 = ~n9706 & ~n33358;
  assign n33360 = ~controllable_BtoS_ACK0 & ~n33359;
  assign n33361 = ~n33353 & ~n33360;
  assign n33362 = n4465 & ~n33361;
  assign n33363 = ~controllable_DEQ & ~n9801;
  assign n33364 = ~n9854 & ~n33363;
  assign n33365 = ~i_FULL & ~n33364;
  assign n33366 = ~n9846 & ~n33365;
  assign n33367 = ~i_nEMPTY & ~n33366;
  assign n33368 = ~n9823 & ~n33367;
  assign n33369 = controllable_BtoS_ACK0 & ~n33368;
  assign n33370 = ~controllable_DEQ & ~n9902;
  assign n33371 = ~n9979 & ~n33370;
  assign n33372 = ~i_FULL & ~n33371;
  assign n33373 = ~n9971 & ~n33372;
  assign n33374 = ~i_nEMPTY & ~n33373;
  assign n33375 = ~n9947 & ~n33374;
  assign n33376 = ~controllable_BtoS_ACK0 & ~n33375;
  assign n33377 = ~n33369 & ~n33376;
  assign n33378 = ~n4465 & ~n33377;
  assign n33379 = ~n33362 & ~n33378;
  assign n33380 = ~i_StoB_REQ10 & ~n33379;
  assign n33381 = ~n33346 & ~n33380;
  assign n33382 = controllable_BtoS_ACK10 & ~n33381;
  assign n33383 = ~n10253 & ~n33380;
  assign n33384 = ~controllable_BtoS_ACK10 & ~n33383;
  assign n33385 = ~n33382 & ~n33384;
  assign n33386 = n4464 & ~n33385;
  assign n33387 = ~controllable_DEQ & ~n10274;
  assign n33388 = ~n10335 & ~n33387;
  assign n33389 = ~i_FULL & ~n33388;
  assign n33390 = ~n10329 & ~n33389;
  assign n33391 = ~i_nEMPTY & ~n33390;
  assign n33392 = ~n10312 & ~n33391;
  assign n33393 = controllable_BtoS_ACK0 & ~n33392;
  assign n33394 = ~controllable_DEQ & ~n10368;
  assign n33395 = ~n10429 & ~n33394;
  assign n33396 = ~i_FULL & ~n33395;
  assign n33397 = ~n10423 & ~n33396;
  assign n33398 = ~i_nEMPTY & ~n33397;
  assign n33399 = ~n10406 & ~n33398;
  assign n33400 = ~controllable_BtoS_ACK0 & ~n33399;
  assign n33401 = ~n33393 & ~n33400;
  assign n33402 = n4465 & ~n33401;
  assign n33403 = ~n33206 & ~n33400;
  assign n33404 = ~n4465 & ~n33403;
  assign n33405 = ~n33402 & ~n33404;
  assign n33406 = i_StoB_REQ10 & ~n33405;
  assign n33407 = ~controllable_DEQ & ~n10485;
  assign n33408 = ~n10566 & ~n33407;
  assign n33409 = ~i_FULL & ~n33408;
  assign n33410 = ~n10558 & ~n33409;
  assign n33411 = ~i_nEMPTY & ~n33410;
  assign n33412 = ~n10534 & ~n33411;
  assign n33413 = controllable_BtoS_ACK0 & ~n33412;
  assign n33414 = ~controllable_DEQ & ~n10612;
  assign n33415 = ~n10693 & ~n33414;
  assign n33416 = ~i_FULL & ~n33415;
  assign n33417 = ~n10685 & ~n33416;
  assign n33418 = ~i_nEMPTY & ~n33417;
  assign n33419 = ~n10661 & ~n33418;
  assign n33420 = ~controllable_BtoS_ACK0 & ~n33419;
  assign n33421 = ~n33413 & ~n33420;
  assign n33422 = n4465 & ~n33421;
  assign n33423 = ~controllable_DEQ & ~n10726;
  assign n33424 = ~n10766 & ~n33423;
  assign n33425 = ~i_FULL & ~n33424;
  assign n33426 = ~n10760 & ~n33425;
  assign n33427 = ~i_nEMPTY & ~n33426;
  assign n33428 = ~n10744 & ~n33427;
  assign n33429 = controllable_BtoS_ACK0 & ~n33428;
  assign n33430 = ~controllable_DEQ & ~n10797;
  assign n33431 = ~n10860 & ~n33430;
  assign n33432 = ~i_FULL & ~n33431;
  assign n33433 = ~n10854 & ~n33432;
  assign n33434 = ~i_nEMPTY & ~n33433;
  assign n33435 = ~n10838 & ~n33434;
  assign n33436 = ~controllable_BtoS_ACK0 & ~n33435;
  assign n33437 = ~n33429 & ~n33436;
  assign n33438 = ~n4465 & ~n33437;
  assign n33439 = ~n33422 & ~n33438;
  assign n33440 = ~i_StoB_REQ10 & ~n33439;
  assign n33441 = ~n33406 & ~n33440;
  assign n33442 = controllable_BtoS_ACK10 & ~n33441;
  assign n33443 = ~n11122 & ~n33440;
  assign n33444 = ~controllable_BtoS_ACK10 & ~n33443;
  assign n33445 = ~n33442 & ~n33444;
  assign n33446 = ~n4464 & ~n33445;
  assign n33447 = ~n33386 & ~n33446;
  assign n33448 = ~n4463 & ~n33447;
  assign n33449 = ~n33319 & ~n33448;
  assign n33450 = n4462 & ~n33449;
  assign n33451 = ~controllable_DEQ & ~n11163;
  assign n33452 = ~n11209 & ~n33451;
  assign n33453 = ~i_FULL & ~n33452;
  assign n33454 = ~n11201 & ~n33453;
  assign n33455 = ~i_nEMPTY & ~n33454;
  assign n33456 = ~n11179 & ~n33455;
  assign n33457 = controllable_BtoS_ACK0 & ~n33456;
  assign n33458 = ~n33213 & ~n33457;
  assign n33459 = n4465 & ~n33458;
  assign n33460 = ~n33215 & ~n33459;
  assign n33461 = i_StoB_REQ10 & ~n33460;
  assign n33462 = ~controllable_DEQ & ~n11243;
  assign n33463 = ~n11282 & ~n33462;
  assign n33464 = ~i_FULL & ~n33463;
  assign n33465 = ~n11276 & ~n33464;
  assign n33466 = ~i_nEMPTY & ~n33465;
  assign n33467 = ~n11259 & ~n33466;
  assign n33468 = controllable_BtoS_ACK0 & ~n33467;
  assign n33469 = ~controllable_DEQ & ~n11322;
  assign n33470 = ~n11364 & ~n33469;
  assign n33471 = ~i_FULL & ~n33470;
  assign n33472 = ~n11358 & ~n33471;
  assign n33473 = ~i_nEMPTY & ~n33472;
  assign n33474 = ~n11339 & ~n33473;
  assign n33475 = ~controllable_BtoS_ACK0 & ~n33474;
  assign n33476 = ~n33468 & ~n33475;
  assign n33477 = ~i_StoB_REQ10 & ~n33476;
  assign n33478 = ~n33461 & ~n33477;
  assign n33479 = controllable_BtoS_ACK10 & ~n33478;
  assign n33480 = ~controllable_DEQ & ~n11673;
  assign n33481 = ~n11756 & ~n33480;
  assign n33482 = ~i_FULL & ~n33481;
  assign n33483 = ~n11748 & ~n33482;
  assign n33484 = ~i_nEMPTY & ~n33483;
  assign n33485 = ~n11722 & ~n33484;
  assign n33486 = controllable_BtoS_ACK0 & ~n33485;
  assign n33487 = ~controllable_DEQ & ~n11820;
  assign n33488 = ~n11903 & ~n33487;
  assign n33489 = ~i_FULL & ~n33488;
  assign n33490 = ~n11895 & ~n33489;
  assign n33491 = ~i_nEMPTY & ~n33490;
  assign n33492 = ~n11869 & ~n33491;
  assign n33493 = ~controllable_BtoS_ACK0 & ~n33492;
  assign n33494 = ~n33486 & ~n33493;
  assign n33495 = n4465 & ~n33494;
  assign n33496 = ~n33249 & ~n33495;
  assign n33497 = ~i_StoB_REQ10 & ~n33496;
  assign n33498 = ~n11623 & ~n33497;
  assign n33499 = ~controllable_BtoS_ACK10 & ~n33498;
  assign n33500 = ~n33479 & ~n33499;
  assign n33501 = n4464 & ~n33500;
  assign n33502 = ~n33277 & ~n33477;
  assign n33503 = controllable_BtoS_ACK10 & ~n33502;
  assign n33504 = ~n12149 & ~n33311;
  assign n33505 = ~controllable_BtoS_ACK10 & ~n33504;
  assign n33506 = ~n33503 & ~n33505;
  assign n33507 = ~n4464 & ~n33506;
  assign n33508 = ~n33501 & ~n33507;
  assign n33509 = n4463 & ~n33508;
  assign n33510 = ~controllable_DEQ & ~n12182;
  assign n33511 = ~n12234 & ~n33510;
  assign n33512 = ~i_FULL & ~n33511;
  assign n33513 = ~n12226 & ~n33512;
  assign n33514 = ~i_nEMPTY & ~n33513;
  assign n33515 = ~n12203 & ~n33514;
  assign n33516 = controllable_BtoS_ACK0 & ~n33515;
  assign n33517 = ~controllable_DEQ & ~n12273;
  assign n33518 = ~n12315 & ~n33517;
  assign n33519 = ~i_FULL & ~n33518;
  assign n33520 = ~n12307 & ~n33519;
  assign n33521 = ~i_nEMPTY & ~n33520;
  assign n33522 = ~n12289 & ~n33521;
  assign n33523 = ~controllable_BtoS_ACK0 & ~n33522;
  assign n33524 = ~n33516 & ~n33523;
  assign n33525 = n4465 & ~n33524;
  assign n33526 = ~controllable_DEQ & ~n9006;
  assign n33527 = ~n9042 & ~n33526;
  assign n33528 = ~i_FULL & ~n33527;
  assign n33529 = ~n12341 & ~n33528;
  assign n33530 = ~i_nEMPTY & ~n33529;
  assign n33531 = ~n12337 & ~n33530;
  assign n33532 = ~controllable_BtoS_ACK0 & ~n33531;
  assign n33533 = ~n33206 & ~n33532;
  assign n33534 = ~n4465 & ~n33533;
  assign n33535 = ~n33525 & ~n33534;
  assign n33536 = i_StoB_REQ10 & ~n33535;
  assign n33537 = ~n33477 & ~n33536;
  assign n33538 = controllable_BtoS_ACK10 & ~n33537;
  assign n33539 = ~controllable_DEQ & ~n12564;
  assign n33540 = ~n12627 & ~n33539;
  assign n33541 = ~i_FULL & ~n33540;
  assign n33542 = ~n12621 & ~n33541;
  assign n33543 = ~i_nEMPTY & ~n33542;
  assign n33544 = ~n12605 & ~n33543;
  assign n33545 = controllable_BtoS_ACK0 & ~n33544;
  assign n33546 = ~controllable_DEQ & ~n12660;
  assign n33547 = ~n12723 & ~n33546;
  assign n33548 = ~i_FULL & ~n33547;
  assign n33549 = ~n12717 & ~n33548;
  assign n33550 = ~i_nEMPTY & ~n33549;
  assign n33551 = ~n12701 & ~n33550;
  assign n33552 = ~controllable_BtoS_ACK0 & ~n33551;
  assign n33553 = ~n33545 & ~n33552;
  assign n33554 = n4465 & ~n33553;
  assign n33555 = ~controllable_DEQ & ~n12748;
  assign n33556 = ~n12773 & ~n33555;
  assign n33557 = ~i_FULL & ~n33556;
  assign n33558 = ~n12767 & ~n33557;
  assign n33559 = ~i_nEMPTY & ~n33558;
  assign n33560 = ~n12757 & ~n33559;
  assign n33561 = controllable_BtoS_ACK0 & ~n33560;
  assign n33562 = ~n33376 & ~n33561;
  assign n33563 = ~n4465 & ~n33562;
  assign n33564 = ~n33554 & ~n33563;
  assign n33565 = ~i_StoB_REQ10 & ~n33564;
  assign n33566 = ~n12547 & ~n33565;
  assign n33567 = ~controllable_BtoS_ACK10 & ~n33566;
  assign n33568 = ~n33538 & ~n33567;
  assign n33569 = n4464 & ~n33568;
  assign n33570 = ~controllable_DEQ & ~n10299;
  assign n33571 = ~n10335 & ~n33570;
  assign n33572 = ~i_FULL & ~n33571;
  assign n33573 = ~n12805 & ~n33572;
  assign n33574 = ~i_nEMPTY & ~n33573;
  assign n33575 = ~n12797 & ~n33574;
  assign n33576 = controllable_BtoS_ACK0 & ~n33575;
  assign n33577 = ~controllable_DEQ & ~n10393;
  assign n33578 = ~n10429 & ~n33577;
  assign n33579 = ~i_FULL & ~n33578;
  assign n33580 = ~n12835 & ~n33579;
  assign n33581 = ~i_nEMPTY & ~n33580;
  assign n33582 = ~n12827 & ~n33581;
  assign n33583 = ~controllable_BtoS_ACK0 & ~n33582;
  assign n33584 = ~n33576 & ~n33583;
  assign n33585 = n4465 & ~n33584;
  assign n33586 = ~n33206 & ~n33583;
  assign n33587 = ~n4465 & ~n33586;
  assign n33588 = ~n33585 & ~n33587;
  assign n33589 = i_StoB_REQ10 & ~n33588;
  assign n33590 = ~n33477 & ~n33589;
  assign n33591 = controllable_BtoS_ACK10 & ~n33590;
  assign n33592 = ~controllable_DEQ & ~n13042;
  assign n33593 = ~n13079 & ~n33592;
  assign n33594 = ~i_FULL & ~n33593;
  assign n33595 = ~n13073 & ~n33594;
  assign n33596 = ~i_nEMPTY & ~n33595;
  assign n33597 = ~n13063 & ~n33596;
  assign n33598 = controllable_BtoS_ACK0 & ~n33597;
  assign n33599 = ~controllable_DEQ & ~n13096;
  assign n33600 = ~n13133 & ~n33599;
  assign n33601 = ~i_FULL & ~n33600;
  assign n33602 = ~n13127 & ~n33601;
  assign n33603 = ~i_nEMPTY & ~n33602;
  assign n33604 = ~n13117 & ~n33603;
  assign n33605 = ~controllable_BtoS_ACK0 & ~n33604;
  assign n33606 = ~n33598 & ~n33605;
  assign n33607 = n4465 & ~n33606;
  assign n33608 = ~n33438 & ~n33607;
  assign n33609 = ~i_StoB_REQ10 & ~n33608;
  assign n33610 = ~n13033 & ~n33609;
  assign n33611 = ~controllable_BtoS_ACK10 & ~n33610;
  assign n33612 = ~n33591 & ~n33611;
  assign n33613 = ~n4464 & ~n33612;
  assign n33614 = ~n33569 & ~n33613;
  assign n33615 = ~n4463 & ~n33614;
  assign n33616 = ~n33509 & ~n33615;
  assign n33617 = ~n4462 & ~n33616;
  assign n33618 = ~n33450 & ~n33617;
  assign n33619 = n4461 & ~n33618;
  assign n33620 = ~controllable_DEQ & ~n13160;
  assign n33621 = ~n5091 & ~n33620;
  assign n33622 = ~i_FULL & ~n33621;
  assign n33623 = ~n13169 & ~n33622;
  assign n33624 = ~i_nEMPTY & ~n33623;
  assign n33625 = ~n13165 & ~n33624;
  assign n33626 = controllable_BtoS_ACK0 & ~n33625;
  assign n33627 = ~controllable_DEQ & ~n13187;
  assign n33628 = ~n5188 & ~n33627;
  assign n33629 = ~i_FULL & ~n33628;
  assign n33630 = ~n13196 & ~n33629;
  assign n33631 = ~i_nEMPTY & ~n33630;
  assign n33632 = ~n13192 & ~n33631;
  assign n33633 = ~controllable_BtoS_ACK0 & ~n33632;
  assign n33634 = ~n33626 & ~n33633;
  assign n33635 = n4465 & ~n33634;
  assign n33636 = ~controllable_DEQ & ~n13216;
  assign n33637 = ~n5402 & ~n33636;
  assign n33638 = ~i_FULL & ~n33637;
  assign n33639 = ~n13225 & ~n33638;
  assign n33640 = ~i_nEMPTY & ~n33639;
  assign n33641 = ~n13221 & ~n33640;
  assign n33642 = ~controllable_BtoS_ACK0 & ~n33641;
  assign n33643 = ~n33206 & ~n33642;
  assign n33644 = ~n4465 & ~n33643;
  assign n33645 = ~n33635 & ~n33644;
  assign n33646 = i_StoB_REQ10 & ~n33645;
  assign n33647 = ~controllable_DEQ & ~n13251;
  assign n33648 = ~n6871 & ~n33647;
  assign n33649 = ~i_FULL & ~n33648;
  assign n33650 = ~n13294 & ~n33649;
  assign n33651 = ~i_nEMPTY & ~n33650;
  assign n33652 = ~n13283 & ~n33651;
  assign n33653 = controllable_BtoS_ACK0 & ~n33652;
  assign n33654 = ~controllable_DEQ & ~n13315;
  assign n33655 = ~n7037 & ~n33654;
  assign n33656 = ~i_FULL & ~n33655;
  assign n33657 = ~n13358 & ~n33656;
  assign n33658 = ~i_nEMPTY & ~n33657;
  assign n33659 = ~n13347 & ~n33658;
  assign n33660 = ~controllable_BtoS_ACK0 & ~n33659;
  assign n33661 = ~n33653 & ~n33660;
  assign n33662 = n4465 & ~n33661;
  assign n33663 = ~controllable_DEQ & ~n13381;
  assign n33664 = ~n7157 & ~n33663;
  assign n33665 = ~i_FULL & ~n33664;
  assign n33666 = ~n13404 & ~n33665;
  assign n33667 = ~i_nEMPTY & ~n33666;
  assign n33668 = ~n13393 & ~n33667;
  assign n33669 = controllable_BtoS_ACK0 & ~n33668;
  assign n33670 = ~controllable_DEQ & ~n13421;
  assign n33671 = ~n7363 & ~n33670;
  assign n33672 = ~i_FULL & ~n33671;
  assign n33673 = ~n13454 & ~n33672;
  assign n33674 = ~i_nEMPTY & ~n33673;
  assign n33675 = ~n13446 & ~n33674;
  assign n33676 = ~controllable_BtoS_ACK0 & ~n33675;
  assign n33677 = ~n33669 & ~n33676;
  assign n33678 = ~n4465 & ~n33677;
  assign n33679 = ~n33662 & ~n33678;
  assign n33680 = ~i_StoB_REQ10 & ~n33679;
  assign n33681 = ~n33646 & ~n33680;
  assign n33682 = controllable_BtoS_ACK10 & ~n33681;
  assign n33683 = ~n13630 & ~n33680;
  assign n33684 = ~controllable_BtoS_ACK10 & ~n33683;
  assign n33685 = ~n33682 & ~n33684;
  assign n33686 = n4464 & ~n33685;
  assign n33687 = ~controllable_DEQ & ~n13639;
  assign n33688 = ~n7769 & ~n33687;
  assign n33689 = ~i_FULL & ~n33688;
  assign n33690 = ~n13648 & ~n33689;
  assign n33691 = ~i_nEMPTY & ~n33690;
  assign n33692 = ~n13644 & ~n33691;
  assign n33693 = controllable_BtoS_ACK0 & ~n33692;
  assign n33694 = ~controllable_DEQ & ~n13666;
  assign n33695 = ~n7861 & ~n33694;
  assign n33696 = ~i_FULL & ~n33695;
  assign n33697 = ~n13675 & ~n33696;
  assign n33698 = ~i_nEMPTY & ~n33697;
  assign n33699 = ~n13671 & ~n33698;
  assign n33700 = ~controllable_BtoS_ACK0 & ~n33699;
  assign n33701 = ~n33693 & ~n33700;
  assign n33702 = n4465 & ~n33701;
  assign n33703 = ~n33206 & ~n33700;
  assign n33704 = ~n4465 & ~n33703;
  assign n33705 = ~n33702 & ~n33704;
  assign n33706 = i_StoB_REQ10 & ~n33705;
  assign n33707 = ~controllable_DEQ & ~n13703;
  assign n33708 = ~n8033 & ~n33707;
  assign n33709 = ~i_FULL & ~n33708;
  assign n33710 = ~n13746 & ~n33709;
  assign n33711 = ~i_nEMPTY & ~n33710;
  assign n33712 = ~n13735 & ~n33711;
  assign n33713 = controllable_BtoS_ACK0 & ~n33712;
  assign n33714 = ~controllable_DEQ & ~n13767;
  assign n33715 = ~n8197 & ~n33714;
  assign n33716 = ~i_FULL & ~n33715;
  assign n33717 = ~n13810 & ~n33716;
  assign n33718 = ~i_nEMPTY & ~n33717;
  assign n33719 = ~n13799 & ~n33718;
  assign n33720 = ~controllable_BtoS_ACK0 & ~n33719;
  assign n33721 = ~n33713 & ~n33720;
  assign n33722 = n4465 & ~n33721;
  assign n33723 = ~controllable_DEQ & ~n13829;
  assign n33724 = ~n8293 & ~n33723;
  assign n33725 = ~i_FULL & ~n33724;
  assign n33726 = ~n13846 & ~n33725;
  assign n33727 = ~i_nEMPTY & ~n33726;
  assign n33728 = ~n13838 & ~n33727;
  assign n33729 = controllable_BtoS_ACK0 & ~n33728;
  assign n33730 = ~controllable_DEQ & ~n13863;
  assign n33731 = ~n8433 & ~n33730;
  assign n33732 = ~i_FULL & ~n33731;
  assign n33733 = ~n13896 & ~n33732;
  assign n33734 = ~i_nEMPTY & ~n33733;
  assign n33735 = ~n13888 & ~n33734;
  assign n33736 = ~controllable_BtoS_ACK0 & ~n33735;
  assign n33737 = ~n33729 & ~n33736;
  assign n33738 = ~n4465 & ~n33737;
  assign n33739 = ~n33722 & ~n33738;
  assign n33740 = ~i_StoB_REQ10 & ~n33739;
  assign n33741 = ~n33706 & ~n33740;
  assign n33742 = controllable_BtoS_ACK10 & ~n33741;
  assign n33743 = ~n14064 & ~n33740;
  assign n33744 = ~controllable_BtoS_ACK10 & ~n33743;
  assign n33745 = ~n33742 & ~n33744;
  assign n33746 = ~n4464 & ~n33745;
  assign n33747 = ~n33686 & ~n33746;
  assign n33748 = n4463 & ~n33747;
  assign n33749 = ~n33448 & ~n33748;
  assign n33750 = n4462 & ~n33749;
  assign n33751 = ~controllable_DEQ & ~n14080;
  assign n33752 = ~n11209 & ~n33751;
  assign n33753 = ~i_FULL & ~n33752;
  assign n33754 = ~n14102 & ~n33753;
  assign n33755 = ~i_nEMPTY & ~n33754;
  assign n33756 = ~n14092 & ~n33755;
  assign n33757 = controllable_BtoS_ACK0 & ~n33756;
  assign n33758 = ~controllable_DEQ & ~n14123;
  assign n33759 = ~n5402 & ~n33758;
  assign n33760 = ~i_FULL & ~n33759;
  assign n33761 = ~n14145 & ~n33760;
  assign n33762 = ~i_nEMPTY & ~n33761;
  assign n33763 = ~n14135 & ~n33762;
  assign n33764 = ~controllable_BtoS_ACK0 & ~n33763;
  assign n33765 = ~n33757 & ~n33764;
  assign n33766 = n4465 & ~n33765;
  assign n33767 = ~n33644 & ~n33766;
  assign n33768 = i_StoB_REQ10 & ~n33767;
  assign n33769 = ~n33477 & ~n33768;
  assign n33770 = controllable_BtoS_ACK10 & ~n33769;
  assign n33771 = ~controllable_DEQ & ~n14264;
  assign n33772 = ~n11756 & ~n33771;
  assign n33773 = ~i_FULL & ~n33772;
  assign n33774 = ~n14297 & ~n33773;
  assign n33775 = ~i_nEMPTY & ~n33774;
  assign n33776 = ~n14289 & ~n33775;
  assign n33777 = controllable_BtoS_ACK0 & ~n33776;
  assign n33778 = ~controllable_DEQ & ~n14314;
  assign n33779 = ~n11903 & ~n33778;
  assign n33780 = ~i_FULL & ~n33779;
  assign n33781 = ~n14347 & ~n33780;
  assign n33782 = ~i_nEMPTY & ~n33781;
  assign n33783 = ~n14339 & ~n33782;
  assign n33784 = ~controllable_BtoS_ACK0 & ~n33783;
  assign n33785 = ~n33777 & ~n33784;
  assign n33786 = n4465 & ~n33785;
  assign n33787 = ~controllable_DEQ & ~n14366;
  assign n33788 = ~n7157 & ~n33787;
  assign n33789 = ~i_FULL & ~n33788;
  assign n33790 = ~n14375 & ~n33789;
  assign n33791 = ~i_nEMPTY & ~n33790;
  assign n33792 = ~n14371 & ~n33791;
  assign n33793 = controllable_BtoS_ACK0 & ~n33792;
  assign n33794 = ~n33676 & ~n33793;
  assign n33795 = ~n4465 & ~n33794;
  assign n33796 = ~n33786 & ~n33795;
  assign n33797 = ~i_StoB_REQ10 & ~n33796;
  assign n33798 = ~n14259 & ~n33797;
  assign n33799 = ~controllable_BtoS_ACK10 & ~n33798;
  assign n33800 = ~n33770 & ~n33799;
  assign n33801 = n4464 & ~n33800;
  assign n33802 = ~n33477 & ~n33706;
  assign n33803 = controllable_BtoS_ACK10 & ~n33802;
  assign n33804 = ~controllable_DEQ & ~n14498;
  assign n33805 = ~n8033 & ~n33804;
  assign n33806 = ~i_FULL & ~n33805;
  assign n33807 = ~n14519 & ~n33806;
  assign n33808 = ~i_nEMPTY & ~n33807;
  assign n33809 = ~n14515 & ~n33808;
  assign n33810 = controllable_BtoS_ACK0 & ~n33809;
  assign n33811 = ~controllable_DEQ & ~n14536;
  assign n33812 = ~n8197 & ~n33811;
  assign n33813 = ~i_FULL & ~n33812;
  assign n33814 = ~n14557 & ~n33813;
  assign n33815 = ~i_nEMPTY & ~n33814;
  assign n33816 = ~n14553 & ~n33815;
  assign n33817 = ~controllable_BtoS_ACK0 & ~n33816;
  assign n33818 = ~n33810 & ~n33817;
  assign n33819 = n4465 & ~n33818;
  assign n33820 = ~n33738 & ~n33819;
  assign n33821 = ~i_StoB_REQ10 & ~n33820;
  assign n33822 = ~n14493 & ~n33821;
  assign n33823 = ~controllable_BtoS_ACK10 & ~n33822;
  assign n33824 = ~n33803 & ~n33823;
  assign n33825 = ~n4464 & ~n33824;
  assign n33826 = ~n33801 & ~n33825;
  assign n33827 = n4463 & ~n33826;
  assign n33828 = ~n33615 & ~n33827;
  assign n33829 = ~n4462 & ~n33828;
  assign n33830 = ~n33750 & ~n33829;
  assign n33831 = ~n4461 & ~n33830;
  assign n33832 = ~n33619 & ~n33831;
  assign n33833 = ~n4459 & ~n33832;
  assign n33834 = ~controllable_DEQ & ~n14603;
  assign n33835 = ~n14648 & ~n33834;
  assign n33836 = ~i_FULL & ~n33835;
  assign n33837 = ~n14640 & ~n33836;
  assign n33838 = ~i_nEMPTY & ~n33837;
  assign n33839 = ~n14621 & ~n33838;
  assign n33840 = controllable_BtoS_ACK0 & ~n33839;
  assign n33841 = ~controllable_DEQ & ~n14678;
  assign n33842 = ~n14723 & ~n33841;
  assign n33843 = ~i_FULL & ~n33842;
  assign n33844 = ~n14715 & ~n33843;
  assign n33845 = ~i_nEMPTY & ~n33844;
  assign n33846 = ~n14696 & ~n33845;
  assign n33847 = ~controllable_BtoS_ACK0 & ~n33846;
  assign n33848 = ~n33840 & ~n33847;
  assign n33849 = n4465 & ~n33848;
  assign n33850 = ~controllable_DEQ & ~n14754;
  assign n33851 = ~n14798 & ~n33850;
  assign n33852 = ~i_FULL & ~n33851;
  assign n33853 = ~n14790 & ~n33852;
  assign n33854 = ~i_nEMPTY & ~n33853;
  assign n33855 = ~n14771 & ~n33854;
  assign n33856 = controllable_BtoS_ACK0 & ~n33855;
  assign n33857 = ~controllable_DEQ & ~n14829;
  assign n33858 = ~n14874 & ~n33857;
  assign n33859 = ~i_FULL & ~n33858;
  assign n33860 = ~n14866 & ~n33859;
  assign n33861 = ~i_nEMPTY & ~n33860;
  assign n33862 = ~n14847 & ~n33861;
  assign n33863 = ~controllable_BtoS_ACK0 & ~n33862;
  assign n33864 = ~n33856 & ~n33863;
  assign n33865 = ~n4465 & ~n33864;
  assign n33866 = ~n33849 & ~n33865;
  assign n33867 = i_StoB_REQ10 & ~n33866;
  assign n33868 = ~controllable_DEQ & ~n14909;
  assign n33869 = ~n15020 & ~n33868;
  assign n33870 = ~i_FULL & ~n33869;
  assign n33871 = ~n15003 & ~n33870;
  assign n33872 = ~i_nEMPTY & ~n33871;
  assign n33873 = ~n14968 & ~n33872;
  assign n33874 = controllable_BtoS_ACK0 & ~n33873;
  assign n33875 = ~controllable_DEQ & ~n15051;
  assign n33876 = ~n15162 & ~n33875;
  assign n33877 = ~i_FULL & ~n33876;
  assign n33878 = ~n15145 & ~n33877;
  assign n33879 = ~i_nEMPTY & ~n33878;
  assign n33880 = ~n15110 & ~n33879;
  assign n33881 = ~controllable_BtoS_ACK0 & ~n33880;
  assign n33882 = ~n33874 & ~n33881;
  assign n33883 = n4465 & ~n33882;
  assign n33884 = ~controllable_DEQ & ~n15195;
  assign n33885 = ~n15255 & ~n33884;
  assign n33886 = ~i_FULL & ~n33885;
  assign n33887 = ~n15243 & ~n33886;
  assign n33888 = ~i_nEMPTY & ~n33887;
  assign n33889 = ~n15215 & ~n33888;
  assign n33890 = controllable_BtoS_ACK0 & ~n33889;
  assign n33891 = ~controllable_DEQ & ~n15286;
  assign n33892 = ~n15397 & ~n33891;
  assign n33893 = ~i_FULL & ~n33892;
  assign n33894 = ~n15380 & ~n33893;
  assign n33895 = ~i_nEMPTY & ~n33894;
  assign n33896 = ~n15345 & ~n33895;
  assign n33897 = ~controllable_BtoS_ACK0 & ~n33896;
  assign n33898 = ~n33890 & ~n33897;
  assign n33899 = ~n4465 & ~n33898;
  assign n33900 = ~n33883 & ~n33899;
  assign n33901 = ~i_StoB_REQ10 & ~n33900;
  assign n33902 = ~n33867 & ~n33901;
  assign n33903 = controllable_BtoS_ACK10 & ~n33902;
  assign n33904 = ~n15715 & ~n33901;
  assign n33905 = ~controllable_BtoS_ACK10 & ~n33904;
  assign n33906 = ~n33903 & ~n33905;
  assign n33907 = n4464 & ~n33906;
  assign n33908 = ~controllable_DEQ & ~n15737;
  assign n33909 = ~n15782 & ~n33908;
  assign n33910 = ~i_FULL & ~n33909;
  assign n33911 = ~n15774 & ~n33910;
  assign n33912 = ~i_nEMPTY & ~n33911;
  assign n33913 = ~n15755 & ~n33912;
  assign n33914 = controllable_BtoS_ACK0 & ~n33913;
  assign n33915 = ~controllable_DEQ & ~n15812;
  assign n33916 = ~n15857 & ~n33915;
  assign n33917 = ~i_FULL & ~n33916;
  assign n33918 = ~n15849 & ~n33917;
  assign n33919 = ~i_nEMPTY & ~n33918;
  assign n33920 = ~n15830 & ~n33919;
  assign n33921 = ~controllable_BtoS_ACK0 & ~n33920;
  assign n33922 = ~n33914 & ~n33921;
  assign n33923 = n4465 & ~n33922;
  assign n33924 = ~n33856 & ~n33921;
  assign n33925 = ~n4465 & ~n33924;
  assign n33926 = ~n33923 & ~n33925;
  assign n33927 = i_StoB_REQ10 & ~n33926;
  assign n33928 = ~controllable_DEQ & ~n15894;
  assign n33929 = ~n16005 & ~n33928;
  assign n33930 = ~i_FULL & ~n33929;
  assign n33931 = ~n15988 & ~n33930;
  assign n33932 = ~i_nEMPTY & ~n33931;
  assign n33933 = ~n15953 & ~n33932;
  assign n33934 = controllable_BtoS_ACK0 & ~n33933;
  assign n33935 = ~controllable_DEQ & ~n16036;
  assign n33936 = ~n16147 & ~n33935;
  assign n33937 = ~i_FULL & ~n33936;
  assign n33938 = ~n16130 & ~n33937;
  assign n33939 = ~i_nEMPTY & ~n33938;
  assign n33940 = ~n16095 & ~n33939;
  assign n33941 = ~controllable_BtoS_ACK0 & ~n33940;
  assign n33942 = ~n33934 & ~n33941;
  assign n33943 = n4465 & ~n33942;
  assign n33944 = ~controllable_DEQ & ~n16180;
  assign n33945 = ~n16236 & ~n33944;
  assign n33946 = ~i_FULL & ~n33945;
  assign n33947 = ~n16226 & ~n33946;
  assign n33948 = ~i_nEMPTY & ~n33947;
  assign n33949 = ~n16200 & ~n33948;
  assign n33950 = controllable_BtoS_ACK0 & ~n33949;
  assign n33951 = ~controllable_DEQ & ~n16267;
  assign n33952 = ~n16378 & ~n33951;
  assign n33953 = ~i_FULL & ~n33952;
  assign n33954 = ~n16361 & ~n33953;
  assign n33955 = ~i_nEMPTY & ~n33954;
  assign n33956 = ~n16326 & ~n33955;
  assign n33957 = ~controllable_BtoS_ACK0 & ~n33956;
  assign n33958 = ~n33950 & ~n33957;
  assign n33959 = ~n4465 & ~n33958;
  assign n33960 = ~n33943 & ~n33959;
  assign n33961 = ~i_StoB_REQ10 & ~n33960;
  assign n33962 = ~n33927 & ~n33961;
  assign n33963 = controllable_BtoS_ACK10 & ~n33962;
  assign n33964 = ~n16691 & ~n33961;
  assign n33965 = ~controllable_BtoS_ACK10 & ~n33964;
  assign n33966 = ~n33963 & ~n33965;
  assign n33967 = ~n4464 & ~n33966;
  assign n33968 = ~n33907 & ~n33967;
  assign n33969 = n4463 & ~n33968;
  assign n33970 = ~controllable_DEQ & ~n16700;
  assign n33971 = ~n14648 & ~n33970;
  assign n33972 = ~i_FULL & ~n33971;
  assign n33973 = ~n16711 & ~n33972;
  assign n33974 = ~i_nEMPTY & ~n33973;
  assign n33975 = ~n16707 & ~n33974;
  assign n33976 = controllable_BtoS_ACK0 & ~n33975;
  assign n33977 = ~controllable_DEQ & ~n16726;
  assign n33978 = ~n14723 & ~n33977;
  assign n33979 = ~i_FULL & ~n33978;
  assign n33980 = ~n16739 & ~n33979;
  assign n33981 = ~i_nEMPTY & ~n33980;
  assign n33982 = ~n16735 & ~n33981;
  assign n33983 = ~controllable_BtoS_ACK0 & ~n33982;
  assign n33984 = ~n33976 & ~n33983;
  assign n33985 = n4465 & ~n33984;
  assign n33986 = ~controllable_DEQ & ~n16752;
  assign n33987 = ~n14874 & ~n33986;
  assign n33988 = ~i_FULL & ~n33987;
  assign n33989 = ~n16763 & ~n33988;
  assign n33990 = ~i_nEMPTY & ~n33989;
  assign n33991 = ~n16759 & ~n33990;
  assign n33992 = ~controllable_BtoS_ACK0 & ~n33991;
  assign n33993 = ~n33856 & ~n33992;
  assign n33994 = ~n4465 & ~n33993;
  assign n33995 = ~n33985 & ~n33994;
  assign n33996 = i_StoB_REQ10 & ~n33995;
  assign n33997 = ~controllable_DEQ & ~n16783;
  assign n33998 = ~n15020 & ~n33997;
  assign n33999 = ~i_FULL & ~n33998;
  assign n34000 = ~n16812 & ~n33999;
  assign n34001 = ~i_nEMPTY & ~n34000;
  assign n34002 = ~n16802 & ~n34001;
  assign n34003 = controllable_BtoS_ACK0 & ~n34002;
  assign n34004 = ~controllable_DEQ & ~n16828;
  assign n34005 = ~n15162 & ~n34004;
  assign n34006 = ~i_FULL & ~n34005;
  assign n34007 = ~n16857 & ~n34006;
  assign n34008 = ~i_nEMPTY & ~n34007;
  assign n34009 = ~n16847 & ~n34008;
  assign n34010 = ~controllable_BtoS_ACK0 & ~n34009;
  assign n34011 = ~n34003 & ~n34010;
  assign n34012 = n4465 & ~n34011;
  assign n34013 = ~controllable_DEQ & ~n16875;
  assign n34014 = ~n15255 & ~n34013;
  assign n34015 = ~i_FULL & ~n34014;
  assign n34016 = ~n16896 & ~n34015;
  assign n34017 = ~i_nEMPTY & ~n34016;
  assign n34018 = ~n16886 & ~n34017;
  assign n34019 = controllable_BtoS_ACK0 & ~n34018;
  assign n34020 = ~controllable_DEQ & ~n16912;
  assign n34021 = ~n15397 & ~n34020;
  assign n34022 = ~i_FULL & ~n34021;
  assign n34023 = ~n16941 & ~n34022;
  assign n34024 = ~i_nEMPTY & ~n34023;
  assign n34025 = ~n16931 & ~n34024;
  assign n34026 = ~controllable_BtoS_ACK0 & ~n34025;
  assign n34027 = ~n34019 & ~n34026;
  assign n34028 = ~n4465 & ~n34027;
  assign n34029 = ~n34012 & ~n34028;
  assign n34030 = ~i_StoB_REQ10 & ~n34029;
  assign n34031 = ~n33996 & ~n34030;
  assign n34032 = controllable_BtoS_ACK10 & ~n34031;
  assign n34033 = ~n17129 & ~n34030;
  assign n34034 = ~controllable_BtoS_ACK10 & ~n34033;
  assign n34035 = ~n34032 & ~n34034;
  assign n34036 = n4464 & ~n34035;
  assign n34037 = ~controllable_DEQ & ~n17136;
  assign n34038 = ~n15782 & ~n34037;
  assign n34039 = ~i_FULL & ~n34038;
  assign n34040 = ~n17147 & ~n34039;
  assign n34041 = ~i_nEMPTY & ~n34040;
  assign n34042 = ~n17143 & ~n34041;
  assign n34043 = controllable_BtoS_ACK0 & ~n34042;
  assign n34044 = ~controllable_DEQ & ~n17158;
  assign n34045 = ~n15857 & ~n34044;
  assign n34046 = ~i_FULL & ~n34045;
  assign n34047 = ~n17169 & ~n34046;
  assign n34048 = ~i_nEMPTY & ~n34047;
  assign n34049 = ~n17165 & ~n34048;
  assign n34050 = ~controllable_BtoS_ACK0 & ~n34049;
  assign n34051 = ~n34043 & ~n34050;
  assign n34052 = n4465 & ~n34051;
  assign n34053 = ~n33856 & ~n34050;
  assign n34054 = ~n4465 & ~n34053;
  assign n34055 = ~n34052 & ~n34054;
  assign n34056 = i_StoB_REQ10 & ~n34055;
  assign n34057 = ~controllable_DEQ & ~n17191;
  assign n34058 = ~n16005 & ~n34057;
  assign n34059 = ~i_FULL & ~n34058;
  assign n34060 = ~n17220 & ~n34059;
  assign n34061 = ~i_nEMPTY & ~n34060;
  assign n34062 = ~n17210 & ~n34061;
  assign n34063 = controllable_BtoS_ACK0 & ~n34062;
  assign n34064 = ~controllable_DEQ & ~n17236;
  assign n34065 = ~n16147 & ~n34064;
  assign n34066 = ~i_FULL & ~n34065;
  assign n34067 = ~n17265 & ~n34066;
  assign n34068 = ~i_nEMPTY & ~n34067;
  assign n34069 = ~n17255 & ~n34068;
  assign n34070 = ~controllable_BtoS_ACK0 & ~n34069;
  assign n34071 = ~n34063 & ~n34070;
  assign n34072 = n4465 & ~n34071;
  assign n34073 = ~controllable_DEQ & ~n17283;
  assign n34074 = ~n16236 & ~n34073;
  assign n34075 = ~i_FULL & ~n34074;
  assign n34076 = ~n17304 & ~n34075;
  assign n34077 = ~i_nEMPTY & ~n34076;
  assign n34078 = ~n17294 & ~n34077;
  assign n34079 = controllable_BtoS_ACK0 & ~n34078;
  assign n34080 = ~controllable_DEQ & ~n17320;
  assign n34081 = ~n16378 & ~n34080;
  assign n34082 = ~i_FULL & ~n34081;
  assign n34083 = ~n17349 & ~n34082;
  assign n34084 = ~i_nEMPTY & ~n34083;
  assign n34085 = ~n17339 & ~n34084;
  assign n34086 = ~controllable_BtoS_ACK0 & ~n34085;
  assign n34087 = ~n34079 & ~n34086;
  assign n34088 = ~n4465 & ~n34087;
  assign n34089 = ~n34072 & ~n34088;
  assign n34090 = ~i_StoB_REQ10 & ~n34089;
  assign n34091 = ~n34056 & ~n34090;
  assign n34092 = controllable_BtoS_ACK10 & ~n34091;
  assign n34093 = ~n17524 & ~n34090;
  assign n34094 = ~controllable_BtoS_ACK10 & ~n34093;
  assign n34095 = ~n34092 & ~n34094;
  assign n34096 = ~n4464 & ~n34095;
  assign n34097 = ~n34036 & ~n34096;
  assign n34098 = ~n4463 & ~n34097;
  assign n34099 = ~n33969 & ~n34098;
  assign n34100 = n4462 & ~n34099;
  assign n34101 = ~controllable_DEQ & ~n17550;
  assign n34102 = ~n17595 & ~n34101;
  assign n34103 = ~i_FULL & ~n34102;
  assign n34104 = ~n17587 & ~n34103;
  assign n34105 = ~i_nEMPTY & ~n34104;
  assign n34106 = ~n17568 & ~n34105;
  assign n34107 = controllable_BtoS_ACK0 & ~n34106;
  assign n34108 = ~n33863 & ~n34107;
  assign n34109 = n4465 & ~n34108;
  assign n34110 = ~n33865 & ~n34109;
  assign n34111 = i_StoB_REQ10 & ~n34110;
  assign n34112 = ~controllable_DEQ & ~n17625;
  assign n34113 = ~n17673 & ~n34112;
  assign n34114 = ~i_FULL & ~n34113;
  assign n34115 = ~n17663 & ~n34114;
  assign n34116 = ~i_nEMPTY & ~n34115;
  assign n34117 = ~n17641 & ~n34116;
  assign n34118 = controllable_BtoS_ACK0 & ~n34117;
  assign n34119 = ~controllable_DEQ & ~n17704;
  assign n34120 = ~n17774 & ~n34119;
  assign n34121 = ~i_FULL & ~n34120;
  assign n34122 = ~n17757 & ~n34121;
  assign n34123 = ~i_nEMPTY & ~n34122;
  assign n34124 = ~n17724 & ~n34123;
  assign n34125 = ~controllable_BtoS_ACK0 & ~n34124;
  assign n34126 = ~n34118 & ~n34125;
  assign n34127 = ~i_StoB_REQ10 & ~n34126;
  assign n34128 = ~n34111 & ~n34127;
  assign n34129 = controllable_BtoS_ACK10 & ~n34128;
  assign n34130 = ~controllable_DEQ & ~n17979;
  assign n34131 = ~n18090 & ~n34130;
  assign n34132 = ~i_FULL & ~n34131;
  assign n34133 = ~n18073 & ~n34132;
  assign n34134 = ~i_nEMPTY & ~n34133;
  assign n34135 = ~n18038 & ~n34134;
  assign n34136 = controllable_BtoS_ACK0 & ~n34135;
  assign n34137 = ~controllable_DEQ & ~n18121;
  assign n34138 = ~n18232 & ~n34137;
  assign n34139 = ~i_FULL & ~n34138;
  assign n34140 = ~n18215 & ~n34139;
  assign n34141 = ~i_nEMPTY & ~n34140;
  assign n34142 = ~n18180 & ~n34141;
  assign n34143 = ~controllable_BtoS_ACK0 & ~n34142;
  assign n34144 = ~n34136 & ~n34143;
  assign n34145 = n4465 & ~n34144;
  assign n34146 = ~n33899 & ~n34145;
  assign n34147 = ~i_StoB_REQ10 & ~n34146;
  assign n34148 = ~n17960 & ~n34147;
  assign n34149 = ~controllable_BtoS_ACK10 & ~n34148;
  assign n34150 = ~n34129 & ~n34149;
  assign n34151 = n4464 & ~n34150;
  assign n34152 = ~n33927 & ~n34127;
  assign n34153 = controllable_BtoS_ACK10 & ~n34152;
  assign n34154 = ~n18418 & ~n33961;
  assign n34155 = ~controllable_BtoS_ACK10 & ~n34154;
  assign n34156 = ~n34153 & ~n34155;
  assign n34157 = ~n4464 & ~n34156;
  assign n34158 = ~n34151 & ~n34157;
  assign n34159 = n4463 & ~n34158;
  assign n34160 = ~controllable_DEQ & ~n18431;
  assign n34161 = ~n17595 & ~n34160;
  assign n34162 = ~i_FULL & ~n34161;
  assign n34163 = ~n18444 & ~n34162;
  assign n34164 = ~i_nEMPTY & ~n34163;
  assign n34165 = ~n18440 & ~n34164;
  assign n34166 = controllable_BtoS_ACK0 & ~n34165;
  assign n34167 = ~controllable_DEQ & ~n18459;
  assign n34168 = ~n14874 & ~n34167;
  assign n34169 = ~i_FULL & ~n34168;
  assign n34170 = ~n18472 & ~n34169;
  assign n34171 = ~i_nEMPTY & ~n34170;
  assign n34172 = ~n18468 & ~n34171;
  assign n34173 = ~controllable_BtoS_ACK0 & ~n34172;
  assign n34174 = ~n34166 & ~n34173;
  assign n34175 = n4465 & ~n34174;
  assign n34176 = ~n33994 & ~n34175;
  assign n34177 = i_StoB_REQ10 & ~n34176;
  assign n34178 = ~n34127 & ~n34177;
  assign n34179 = controllable_BtoS_ACK10 & ~n34178;
  assign n34180 = ~controllable_DEQ & ~n18575;
  assign n34181 = ~n18090 & ~n34180;
  assign n34182 = ~i_FULL & ~n34181;
  assign n34183 = ~n18604 & ~n34182;
  assign n34184 = ~i_nEMPTY & ~n34183;
  assign n34185 = ~n18594 & ~n34184;
  assign n34186 = controllable_BtoS_ACK0 & ~n34185;
  assign n34187 = ~controllable_DEQ & ~n18620;
  assign n34188 = ~n18232 & ~n34187;
  assign n34189 = ~i_FULL & ~n34188;
  assign n34190 = ~n18649 & ~n34189;
  assign n34191 = ~i_nEMPTY & ~n34190;
  assign n34192 = ~n18639 & ~n34191;
  assign n34193 = ~controllable_BtoS_ACK0 & ~n34192;
  assign n34194 = ~n34186 & ~n34193;
  assign n34195 = n4465 & ~n34194;
  assign n34196 = ~controllable_DEQ & ~n18662;
  assign n34197 = ~n15255 & ~n34196;
  assign n34198 = ~i_FULL & ~n34197;
  assign n34199 = ~n18675 & ~n34198;
  assign n34200 = ~i_nEMPTY & ~n34199;
  assign n34201 = ~n18669 & ~n34200;
  assign n34202 = controllable_BtoS_ACK0 & ~n34201;
  assign n34203 = ~n34026 & ~n34202;
  assign n34204 = ~n4465 & ~n34203;
  assign n34205 = ~n34195 & ~n34204;
  assign n34206 = ~i_StoB_REQ10 & ~n34205;
  assign n34207 = ~n18567 & ~n34206;
  assign n34208 = ~controllable_BtoS_ACK10 & ~n34207;
  assign n34209 = ~n34179 & ~n34208;
  assign n34210 = n4464 & ~n34209;
  assign n34211 = ~n34056 & ~n34127;
  assign n34212 = controllable_BtoS_ACK10 & ~n34211;
  assign n34213 = ~controllable_DEQ & ~n18769;
  assign n34214 = ~n16005 & ~n34213;
  assign n34215 = ~i_FULL & ~n34214;
  assign n34216 = ~n18798 & ~n34215;
  assign n34217 = ~i_nEMPTY & ~n34216;
  assign n34218 = ~n18788 & ~n34217;
  assign n34219 = controllable_BtoS_ACK0 & ~n34218;
  assign n34220 = ~controllable_DEQ & ~n18814;
  assign n34221 = ~n16147 & ~n34220;
  assign n34222 = ~i_FULL & ~n34221;
  assign n34223 = ~n18843 & ~n34222;
  assign n34224 = ~i_nEMPTY & ~n34223;
  assign n34225 = ~n18833 & ~n34224;
  assign n34226 = ~controllable_BtoS_ACK0 & ~n34225;
  assign n34227 = ~n34219 & ~n34226;
  assign n34228 = n4465 & ~n34227;
  assign n34229 = ~n34088 & ~n34228;
  assign n34230 = ~i_StoB_REQ10 & ~n34229;
  assign n34231 = ~n18761 & ~n34230;
  assign n34232 = ~controllable_BtoS_ACK10 & ~n34231;
  assign n34233 = ~n34212 & ~n34232;
  assign n34234 = ~n4464 & ~n34233;
  assign n34235 = ~n34210 & ~n34234;
  assign n34236 = ~n4463 & ~n34235;
  assign n34237 = ~n34159 & ~n34236;
  assign n34238 = ~n4462 & ~n34237;
  assign n34239 = ~n34100 & ~n34238;
  assign n34240 = n4461 & ~n34239;
  assign n34241 = ~controllable_DEQ & ~n18872;
  assign n34242 = ~n18915 & ~n34241;
  assign n34243 = ~i_FULL & ~n34242;
  assign n34244 = ~n18911 & ~n34243;
  assign n34245 = ~i_nEMPTY & ~n34244;
  assign n34246 = ~n18898 & ~n34245;
  assign n34247 = controllable_BtoS_ACK0 & ~n34246;
  assign n34248 = ~controllable_DEQ & ~n18936;
  assign n34249 = ~n18985 & ~n34248;
  assign n34250 = ~i_FULL & ~n34249;
  assign n34251 = ~n18980 & ~n34250;
  assign n34252 = ~i_nEMPTY & ~n34251;
  assign n34253 = ~n18966 & ~n34252;
  assign n34254 = ~controllable_BtoS_ACK0 & ~n34253;
  assign n34255 = ~n34247 & ~n34254;
  assign n34256 = n4465 & ~n34255;
  assign n34257 = ~controllable_DEQ & ~n19008;
  assign n34258 = ~n19051 & ~n34257;
  assign n34259 = ~i_FULL & ~n34258;
  assign n34260 = ~n19047 & ~n34259;
  assign n34261 = ~i_nEMPTY & ~n34260;
  assign n34262 = ~n19034 & ~n34261;
  assign n34263 = ~controllable_BtoS_ACK0 & ~n34262;
  assign n34264 = ~n33856 & ~n34263;
  assign n34265 = ~n4465 & ~n34264;
  assign n34266 = ~n34256 & ~n34265;
  assign n34267 = i_StoB_REQ10 & ~n34266;
  assign n34268 = ~controllable_DEQ & ~n19083;
  assign n34269 = ~n19148 & ~n34268;
  assign n34270 = ~i_FULL & ~n34269;
  assign n34271 = ~n19142 & ~n34270;
  assign n34272 = ~i_nEMPTY & ~n34271;
  assign n34273 = ~n19120 & ~n34272;
  assign n34274 = controllable_BtoS_ACK0 & ~n34273;
  assign n34275 = ~controllable_DEQ & ~n19176;
  assign n34276 = ~n19241 & ~n34275;
  assign n34277 = ~i_FULL & ~n34276;
  assign n34278 = ~n19235 & ~n34277;
  assign n34279 = ~i_nEMPTY & ~n34278;
  assign n34280 = ~n19213 & ~n34279;
  assign n34281 = ~controllable_BtoS_ACK0 & ~n34280;
  assign n34282 = ~n34274 & ~n34281;
  assign n34283 = n4465 & ~n34282;
  assign n34284 = ~controllable_DEQ & ~n19264;
  assign n34285 = ~n19297 & ~n34284;
  assign n34286 = ~i_FULL & ~n34285;
  assign n34287 = ~n19291 & ~n34286;
  assign n34288 = ~i_nEMPTY & ~n34287;
  assign n34289 = ~n19275 & ~n34288;
  assign n34290 = controllable_BtoS_ACK0 & ~n34289;
  assign n34291 = ~controllable_DEQ & ~n19318;
  assign n34292 = ~n19363 & ~n34291;
  assign n34293 = ~i_FULL & ~n34292;
  assign n34294 = ~n19359 & ~n34293;
  assign n34295 = ~i_nEMPTY & ~n34294;
  assign n34296 = ~n19345 & ~n34295;
  assign n34297 = ~controllable_BtoS_ACK0 & ~n34296;
  assign n34298 = ~n34290 & ~n34297;
  assign n34299 = ~n4465 & ~n34298;
  assign n34300 = ~n34283 & ~n34299;
  assign n34301 = ~i_StoB_REQ10 & ~n34300;
  assign n34302 = ~n34267 & ~n34301;
  assign n34303 = controllable_BtoS_ACK10 & ~n34302;
  assign n34304 = ~n19607 & ~n34301;
  assign n34305 = ~controllable_BtoS_ACK10 & ~n34304;
  assign n34306 = ~n34303 & ~n34305;
  assign n34307 = n4464 & ~n34306;
  assign n34308 = ~controllable_DEQ & ~n19618;
  assign n34309 = ~n19661 & ~n34308;
  assign n34310 = ~i_FULL & ~n34309;
  assign n34311 = ~n19657 & ~n34310;
  assign n34312 = ~i_nEMPTY & ~n34311;
  assign n34313 = ~n19644 & ~n34312;
  assign n34314 = controllable_BtoS_ACK0 & ~n34313;
  assign n34315 = ~controllable_DEQ & ~n19682;
  assign n34316 = ~n19725 & ~n34315;
  assign n34317 = ~i_FULL & ~n34316;
  assign n34318 = ~n19721 & ~n34317;
  assign n34319 = ~i_nEMPTY & ~n34318;
  assign n34320 = ~n19708 & ~n34319;
  assign n34321 = ~controllable_BtoS_ACK0 & ~n34320;
  assign n34322 = ~n34314 & ~n34321;
  assign n34323 = n4465 & ~n34322;
  assign n34324 = ~n33856 & ~n34321;
  assign n34325 = ~n4465 & ~n34324;
  assign n34326 = ~n34323 & ~n34325;
  assign n34327 = i_StoB_REQ10 & ~n34326;
  assign n34328 = ~controllable_DEQ & ~n19752;
  assign n34329 = ~n19805 & ~n34328;
  assign n34330 = ~i_FULL & ~n34329;
  assign n34331 = ~n19799 & ~n34330;
  assign n34332 = ~i_nEMPTY & ~n34331;
  assign n34333 = ~n19783 & ~n34332;
  assign n34334 = controllable_BtoS_ACK0 & ~n34333;
  assign n34335 = ~controllable_DEQ & ~n19826;
  assign n34336 = ~n19879 & ~n34335;
  assign n34337 = ~i_FULL & ~n34336;
  assign n34338 = ~n19873 & ~n34337;
  assign n34339 = ~i_nEMPTY & ~n34338;
  assign n34340 = ~n19857 & ~n34339;
  assign n34341 = ~controllable_BtoS_ACK0 & ~n34340;
  assign n34342 = ~n34334 & ~n34341;
  assign n34343 = n4465 & ~n34342;
  assign n34344 = ~controllable_DEQ & ~n19898;
  assign n34345 = ~n19919 & ~n34344;
  assign n34346 = ~i_FULL & ~n34345;
  assign n34347 = ~n19915 & ~n34346;
  assign n34348 = ~i_nEMPTY & ~n34347;
  assign n34349 = ~n19905 & ~n34348;
  assign n34350 = controllable_BtoS_ACK0 & ~n34349;
  assign n34351 = ~controllable_DEQ & ~n19936;
  assign n34352 = ~n19981 & ~n34351;
  assign n34353 = ~i_FULL & ~n34352;
  assign n34354 = ~n19977 & ~n34353;
  assign n34355 = ~i_nEMPTY & ~n34354;
  assign n34356 = ~n19963 & ~n34355;
  assign n34357 = ~controllable_BtoS_ACK0 & ~n34356;
  assign n34358 = ~n34350 & ~n34357;
  assign n34359 = ~n4465 & ~n34358;
  assign n34360 = ~n34343 & ~n34359;
  assign n34361 = ~i_StoB_REQ10 & ~n34360;
  assign n34362 = ~n34327 & ~n34361;
  assign n34363 = controllable_BtoS_ACK10 & ~n34362;
  assign n34364 = ~n20209 & ~n34361;
  assign n34365 = ~controllable_BtoS_ACK10 & ~n34364;
  assign n34366 = ~n34363 & ~n34365;
  assign n34367 = ~n4464 & ~n34366;
  assign n34368 = ~n34307 & ~n34367;
  assign n34369 = n4462 & ~n34368;
  assign n34370 = ~controllable_DEQ & ~n20224;
  assign n34371 = ~n20258 & ~n34370;
  assign n34372 = ~i_FULL & ~n34371;
  assign n34373 = ~n20253 & ~n34372;
  assign n34374 = ~i_nEMPTY & ~n34373;
  assign n34375 = ~n20237 & ~n34374;
  assign n34376 = controllable_BtoS_ACK0 & ~n34375;
  assign n34377 = ~controllable_DEQ & ~n20279;
  assign n34378 = ~n20311 & ~n34377;
  assign n34379 = ~i_FULL & ~n34378;
  assign n34380 = ~n20306 & ~n34379;
  assign n34381 = ~i_nEMPTY & ~n34380;
  assign n34382 = ~n20290 & ~n34381;
  assign n34383 = ~controllable_BtoS_ACK0 & ~n34382;
  assign n34384 = ~n34376 & ~n34383;
  assign n34385 = n4465 & ~n34384;
  assign n34386 = ~controllable_DEQ & ~n19021;
  assign n34387 = ~n19051 & ~n34386;
  assign n34388 = ~i_FULL & ~n34387;
  assign n34389 = ~n20345 & ~n34388;
  assign n34390 = ~i_nEMPTY & ~n34389;
  assign n34391 = ~n20336 & ~n34390;
  assign n34392 = ~controllable_BtoS_ACK0 & ~n34391;
  assign n34393 = ~n33856 & ~n34392;
  assign n34394 = ~n4465 & ~n34393;
  assign n34395 = ~n34385 & ~n34394;
  assign n34396 = i_StoB_REQ10 & ~n34395;
  assign n34397 = ~n34127 & ~n34396;
  assign n34398 = controllable_BtoS_ACK10 & ~n34397;
  assign n34399 = ~controllable_DEQ & ~n20490;
  assign n34400 = ~n20523 & ~n34399;
  assign n34401 = ~i_FULL & ~n34400;
  assign n34402 = ~n20519 & ~n34401;
  assign n34403 = ~i_nEMPTY & ~n34402;
  assign n34404 = ~n20509 & ~n34403;
  assign n34405 = controllable_BtoS_ACK0 & ~n34404;
  assign n34406 = ~controllable_DEQ & ~n20540;
  assign n34407 = ~n20573 & ~n34406;
  assign n34408 = ~i_FULL & ~n34407;
  assign n34409 = ~n20569 & ~n34408;
  assign n34410 = ~i_nEMPTY & ~n34409;
  assign n34411 = ~n20559 & ~n34410;
  assign n34412 = ~controllable_BtoS_ACK0 & ~n34411;
  assign n34413 = ~n34405 & ~n34412;
  assign n34414 = n4465 & ~n34413;
  assign n34415 = ~controllable_DEQ & ~n20588;
  assign n34416 = ~n20609 & ~n34415;
  assign n34417 = ~i_FULL & ~n34416;
  assign n34418 = ~n20605 & ~n34417;
  assign n34419 = ~i_nEMPTY & ~n34418;
  assign n34420 = ~n20595 & ~n34419;
  assign n34421 = controllable_BtoS_ACK0 & ~n34420;
  assign n34422 = ~n34297 & ~n34421;
  assign n34423 = ~n4465 & ~n34422;
  assign n34424 = ~n34414 & ~n34423;
  assign n34425 = ~i_StoB_REQ10 & ~n34424;
  assign n34426 = ~n20487 & ~n34425;
  assign n34427 = ~controllable_BtoS_ACK10 & ~n34426;
  assign n34428 = ~n34398 & ~n34427;
  assign n34429 = n4464 & ~n34428;
  assign n34430 = ~controllable_DEQ & ~n19631;
  assign n34431 = ~n19661 & ~n34430;
  assign n34432 = ~i_FULL & ~n34431;
  assign n34433 = ~n20639 & ~n34432;
  assign n34434 = ~i_nEMPTY & ~n34433;
  assign n34435 = ~n20633 & ~n34434;
  assign n34436 = controllable_BtoS_ACK0 & ~n34435;
  assign n34437 = ~controllable_DEQ & ~n19695;
  assign n34438 = ~n19725 & ~n34437;
  assign n34439 = ~i_FULL & ~n34438;
  assign n34440 = ~n20661 & ~n34439;
  assign n34441 = ~i_nEMPTY & ~n34440;
  assign n34442 = ~n20655 & ~n34441;
  assign n34443 = ~controllable_BtoS_ACK0 & ~n34442;
  assign n34444 = ~n34436 & ~n34443;
  assign n34445 = n4465 & ~n34444;
  assign n34446 = ~n33856 & ~n34443;
  assign n34447 = ~n4465 & ~n34446;
  assign n34448 = ~n34445 & ~n34447;
  assign n34449 = i_StoB_REQ10 & ~n34448;
  assign n34450 = ~n34127 & ~n34449;
  assign n34451 = controllable_BtoS_ACK10 & ~n34450;
  assign n34452 = ~controllable_DEQ & ~n20788;
  assign n34453 = ~n20821 & ~n34452;
  assign n34454 = ~i_FULL & ~n34453;
  assign n34455 = ~n20817 & ~n34454;
  assign n34456 = ~i_nEMPTY & ~n34455;
  assign n34457 = ~n20807 & ~n34456;
  assign n34458 = controllable_BtoS_ACK0 & ~n34457;
  assign n34459 = ~controllable_DEQ & ~n20838;
  assign n34460 = ~n20871 & ~n34459;
  assign n34461 = ~i_FULL & ~n34460;
  assign n34462 = ~n20867 & ~n34461;
  assign n34463 = ~i_nEMPTY & ~n34462;
  assign n34464 = ~n20857 & ~n34463;
  assign n34465 = ~controllable_BtoS_ACK0 & ~n34464;
  assign n34466 = ~n34458 & ~n34465;
  assign n34467 = n4465 & ~n34466;
  assign n34468 = ~n34359 & ~n34467;
  assign n34469 = ~i_StoB_REQ10 & ~n34468;
  assign n34470 = ~n20785 & ~n34469;
  assign n34471 = ~controllable_BtoS_ACK10 & ~n34470;
  assign n34472 = ~n34451 & ~n34471;
  assign n34473 = ~n4464 & ~n34472;
  assign n34474 = ~n34429 & ~n34473;
  assign n34475 = ~n4462 & ~n34474;
  assign n34476 = ~n34369 & ~n34475;
  assign n34477 = ~n4461 & ~n34476;
  assign n34478 = ~n34240 & ~n34477;
  assign n34479 = n4459 & ~n34478;
  assign n34480 = ~n33833 & ~n34479;
  assign n34481 = n4455 & ~n34480;
  assign n34482 = ~controllable_DEQ & ~n20902;
  assign n34483 = ~n20925 & ~n34482;
  assign n34484 = ~i_FULL & ~n34483;
  assign n34485 = ~n20921 & ~n34484;
  assign n34486 = ~i_nEMPTY & ~n34485;
  assign n34487 = ~n20911 & ~n34486;
  assign n34488 = controllable_BtoS_ACK0 & ~n34487;
  assign n34489 = ~controllable_DEQ & ~n20940;
  assign n34490 = ~n20963 & ~n34489;
  assign n34491 = ~i_FULL & ~n34490;
  assign n34492 = ~n20959 & ~n34491;
  assign n34493 = ~i_nEMPTY & ~n34492;
  assign n34494 = ~n20949 & ~n34493;
  assign n34495 = ~controllable_BtoS_ACK0 & ~n34494;
  assign n34496 = ~n34488 & ~n34495;
  assign n34497 = n4465 & ~n34496;
  assign n34498 = ~controllable_DEQ & ~n20980;
  assign n34499 = ~n21003 & ~n34498;
  assign n34500 = ~i_FULL & ~n34499;
  assign n34501 = ~n20999 & ~n34500;
  assign n34502 = ~i_nEMPTY & ~n34501;
  assign n34503 = ~n20989 & ~n34502;
  assign n34504 = controllable_BtoS_ACK0 & ~n34503;
  assign n34505 = ~controllable_DEQ & ~n21018;
  assign n34506 = ~n21041 & ~n34505;
  assign n34507 = ~i_FULL & ~n34506;
  assign n34508 = ~n21037 & ~n34507;
  assign n34509 = ~i_nEMPTY & ~n34508;
  assign n34510 = ~n21027 & ~n34509;
  assign n34511 = ~controllable_BtoS_ACK0 & ~n34510;
  assign n34512 = ~n34504 & ~n34511;
  assign n34513 = ~n4465 & ~n34512;
  assign n34514 = ~n34497 & ~n34513;
  assign n34515 = i_StoB_REQ10 & ~n34514;
  assign n34516 = ~controllable_DEQ & ~n21060;
  assign n34517 = ~n21101 & ~n34516;
  assign n34518 = ~i_FULL & ~n34517;
  assign n34519 = ~n21097 & ~n34518;
  assign n34520 = ~i_nEMPTY & ~n34519;
  assign n34521 = ~n21085 & ~n34520;
  assign n34522 = controllable_BtoS_ACK0 & ~n34521;
  assign n34523 = ~controllable_DEQ & ~n21116;
  assign n34524 = ~n21157 & ~n34523;
  assign n34525 = ~i_FULL & ~n34524;
  assign n34526 = ~n21153 & ~n34525;
  assign n34527 = ~i_nEMPTY & ~n34526;
  assign n34528 = ~n21141 & ~n34527;
  assign n34529 = ~controllable_BtoS_ACK0 & ~n34528;
  assign n34530 = ~n34522 & ~n34529;
  assign n34531 = n4465 & ~n34530;
  assign n34532 = ~controllable_DEQ & ~n21174;
  assign n34533 = ~n21199 & ~n34532;
  assign n34534 = ~i_FULL & ~n34533;
  assign n34535 = ~n21195 & ~n34534;
  assign n34536 = ~i_nEMPTY & ~n34535;
  assign n34537 = ~n21183 & ~n34536;
  assign n34538 = controllable_BtoS_ACK0 & ~n34537;
  assign n34539 = ~controllable_DEQ & ~n21214;
  assign n34540 = ~n21255 & ~n34539;
  assign n34541 = ~i_FULL & ~n34540;
  assign n34542 = ~n21251 & ~n34541;
  assign n34543 = ~i_nEMPTY & ~n34542;
  assign n34544 = ~n21239 & ~n34543;
  assign n34545 = ~controllable_BtoS_ACK0 & ~n34544;
  assign n34546 = ~n34538 & ~n34545;
  assign n34547 = ~n4465 & ~n34546;
  assign n34548 = ~n34531 & ~n34547;
  assign n34549 = ~i_StoB_REQ10 & ~n34548;
  assign n34550 = ~n34515 & ~n34549;
  assign n34551 = controllable_BtoS_ACK10 & ~n34550;
  assign n34552 = ~n21473 & ~n34549;
  assign n34553 = ~controllable_BtoS_ACK10 & ~n34552;
  assign n34554 = ~n34551 & ~n34553;
  assign n34555 = n4464 & ~n34554;
  assign n34556 = ~controllable_DEQ & ~n21482;
  assign n34557 = ~n21505 & ~n34556;
  assign n34558 = ~i_FULL & ~n34557;
  assign n34559 = ~n21501 & ~n34558;
  assign n34560 = ~i_nEMPTY & ~n34559;
  assign n34561 = ~n21491 & ~n34560;
  assign n34562 = controllable_BtoS_ACK0 & ~n34561;
  assign n34563 = ~controllable_DEQ & ~n21520;
  assign n34564 = ~n21543 & ~n34563;
  assign n34565 = ~i_FULL & ~n34564;
  assign n34566 = ~n21539 & ~n34565;
  assign n34567 = ~i_nEMPTY & ~n34566;
  assign n34568 = ~n21529 & ~n34567;
  assign n34569 = ~controllable_BtoS_ACK0 & ~n34568;
  assign n34570 = ~n34562 & ~n34569;
  assign n34571 = n4465 & ~n34570;
  assign n34572 = ~n34504 & ~n34569;
  assign n34573 = ~n4465 & ~n34572;
  assign n34574 = ~n34571 & ~n34573;
  assign n34575 = i_StoB_REQ10 & ~n34574;
  assign n34576 = ~controllable_DEQ & ~n21564;
  assign n34577 = ~n21605 & ~n34576;
  assign n34578 = ~i_FULL & ~n34577;
  assign n34579 = ~n21601 & ~n34578;
  assign n34580 = ~i_nEMPTY & ~n34579;
  assign n34581 = ~n21589 & ~n34580;
  assign n34582 = controllable_BtoS_ACK0 & ~n34581;
  assign n34583 = ~controllable_DEQ & ~n21620;
  assign n34584 = ~n21661 & ~n34583;
  assign n34585 = ~i_FULL & ~n34584;
  assign n34586 = ~n21657 & ~n34585;
  assign n34587 = ~i_nEMPTY & ~n34586;
  assign n34588 = ~n21645 & ~n34587;
  assign n34589 = ~controllable_BtoS_ACK0 & ~n34588;
  assign n34590 = ~n34582 & ~n34589;
  assign n34591 = n4465 & ~n34590;
  assign n34592 = ~controllable_DEQ & ~n21678;
  assign n34593 = ~n21703 & ~n34592;
  assign n34594 = ~i_FULL & ~n34593;
  assign n34595 = ~n21699 & ~n34594;
  assign n34596 = ~i_nEMPTY & ~n34595;
  assign n34597 = ~n21687 & ~n34596;
  assign n34598 = controllable_BtoS_ACK0 & ~n34597;
  assign n34599 = ~controllable_DEQ & ~n21718;
  assign n34600 = ~n21759 & ~n34599;
  assign n34601 = ~i_FULL & ~n34600;
  assign n34602 = ~n21755 & ~n34601;
  assign n34603 = ~i_nEMPTY & ~n34602;
  assign n34604 = ~n21743 & ~n34603;
  assign n34605 = ~controllable_BtoS_ACK0 & ~n34604;
  assign n34606 = ~n34598 & ~n34605;
  assign n34607 = ~n4465 & ~n34606;
  assign n34608 = ~n34591 & ~n34607;
  assign n34609 = ~i_StoB_REQ10 & ~n34608;
  assign n34610 = ~n34575 & ~n34609;
  assign n34611 = controllable_BtoS_ACK10 & ~n34610;
  assign n34612 = ~n21977 & ~n34609;
  assign n34613 = ~controllable_BtoS_ACK10 & ~n34612;
  assign n34614 = ~n34611 & ~n34613;
  assign n34615 = ~n4464 & ~n34614;
  assign n34616 = ~n34555 & ~n34615;
  assign n34617 = n4463 & ~n34616;
  assign n34618 = ~controllable_DEQ & ~n21988;
  assign n34619 = ~n22023 & ~n34618;
  assign n34620 = ~i_FULL & ~n34619;
  assign n34621 = ~n22019 & ~n34620;
  assign n34622 = ~i_nEMPTY & ~n34621;
  assign n34623 = ~n22009 & ~n34622;
  assign n34624 = controllable_BtoS_ACK0 & ~n34623;
  assign n34625 = ~controllable_DEQ & ~n22038;
  assign n34626 = ~n22073 & ~n34625;
  assign n34627 = ~i_FULL & ~n34626;
  assign n34628 = ~n22069 & ~n34627;
  assign n34629 = ~i_nEMPTY & ~n34628;
  assign n34630 = ~n22059 & ~n34629;
  assign n34631 = ~controllable_BtoS_ACK0 & ~n34630;
  assign n34632 = ~n34624 & ~n34631;
  assign n34633 = n4465 & ~n34632;
  assign n34634 = ~controllable_DEQ & ~n22090;
  assign n34635 = ~n22125 & ~n34634;
  assign n34636 = ~i_FULL & ~n34635;
  assign n34637 = ~n22121 & ~n34636;
  assign n34638 = ~i_nEMPTY & ~n34637;
  assign n34639 = ~n22111 & ~n34638;
  assign n34640 = ~controllable_BtoS_ACK0 & ~n34639;
  assign n34641 = ~n34504 & ~n34640;
  assign n34642 = ~n4465 & ~n34641;
  assign n34643 = ~n34633 & ~n34642;
  assign n34644 = i_StoB_REQ10 & ~n34643;
  assign n34645 = ~controllable_DEQ & ~n22144;
  assign n34646 = ~n22181 & ~n34645;
  assign n34647 = ~i_FULL & ~n34646;
  assign n34648 = ~n22177 & ~n34647;
  assign n34649 = ~i_nEMPTY & ~n34648;
  assign n34650 = ~n22165 & ~n34649;
  assign n34651 = controllable_BtoS_ACK0 & ~n34650;
  assign n34652 = ~controllable_DEQ & ~n22196;
  assign n34653 = ~n22233 & ~n34652;
  assign n34654 = ~i_FULL & ~n34653;
  assign n34655 = ~n22229 & ~n34654;
  assign n34656 = ~i_nEMPTY & ~n34655;
  assign n34657 = ~n22217 & ~n34656;
  assign n34658 = ~controllable_BtoS_ACK0 & ~n34657;
  assign n34659 = ~n34651 & ~n34658;
  assign n34660 = n4465 & ~n34659;
  assign n34661 = ~controllable_DEQ & ~n22250;
  assign n34662 = ~n22275 & ~n34661;
  assign n34663 = ~i_FULL & ~n34662;
  assign n34664 = ~n22271 & ~n34663;
  assign n34665 = ~i_nEMPTY & ~n34664;
  assign n34666 = ~n22259 & ~n34665;
  assign n34667 = controllable_BtoS_ACK0 & ~n34666;
  assign n34668 = ~controllable_DEQ & ~n22290;
  assign n34669 = ~n22327 & ~n34668;
  assign n34670 = ~i_FULL & ~n34669;
  assign n34671 = ~n22323 & ~n34670;
  assign n34672 = ~i_nEMPTY & ~n34671;
  assign n34673 = ~n22311 & ~n34672;
  assign n34674 = ~controllable_BtoS_ACK0 & ~n34673;
  assign n34675 = ~n34667 & ~n34674;
  assign n34676 = ~n4465 & ~n34675;
  assign n34677 = ~n34660 & ~n34676;
  assign n34678 = ~i_StoB_REQ10 & ~n34677;
  assign n34679 = ~n34644 & ~n34678;
  assign n34680 = controllable_BtoS_ACK10 & ~n34679;
  assign n34681 = ~n22533 & ~n34678;
  assign n34682 = ~controllable_BtoS_ACK10 & ~n34681;
  assign n34683 = ~n34680 & ~n34682;
  assign n34684 = n4464 & ~n34683;
  assign n34685 = ~controllable_DEQ & ~n22542;
  assign n34686 = ~n22577 & ~n34685;
  assign n34687 = ~i_FULL & ~n34686;
  assign n34688 = ~n22573 & ~n34687;
  assign n34689 = ~i_nEMPTY & ~n34688;
  assign n34690 = ~n22563 & ~n34689;
  assign n34691 = controllable_BtoS_ACK0 & ~n34690;
  assign n34692 = ~controllable_DEQ & ~n22592;
  assign n34693 = ~n22627 & ~n34692;
  assign n34694 = ~i_FULL & ~n34693;
  assign n34695 = ~n22623 & ~n34694;
  assign n34696 = ~i_nEMPTY & ~n34695;
  assign n34697 = ~n22613 & ~n34696;
  assign n34698 = ~controllable_BtoS_ACK0 & ~n34697;
  assign n34699 = ~n34691 & ~n34698;
  assign n34700 = n4465 & ~n34699;
  assign n34701 = ~n34504 & ~n34698;
  assign n34702 = ~n4465 & ~n34701;
  assign n34703 = ~n34700 & ~n34702;
  assign n34704 = i_StoB_REQ10 & ~n34703;
  assign n34705 = ~controllable_DEQ & ~n22648;
  assign n34706 = ~n22685 & ~n34705;
  assign n34707 = ~i_FULL & ~n34706;
  assign n34708 = ~n22681 & ~n34707;
  assign n34709 = ~i_nEMPTY & ~n34708;
  assign n34710 = ~n22669 & ~n34709;
  assign n34711 = controllable_BtoS_ACK0 & ~n34710;
  assign n34712 = ~controllable_DEQ & ~n22700;
  assign n34713 = ~n22737 & ~n34712;
  assign n34714 = ~i_FULL & ~n34713;
  assign n34715 = ~n22733 & ~n34714;
  assign n34716 = ~i_nEMPTY & ~n34715;
  assign n34717 = ~n22721 & ~n34716;
  assign n34718 = ~controllable_BtoS_ACK0 & ~n34717;
  assign n34719 = ~n34711 & ~n34718;
  assign n34720 = n4465 & ~n34719;
  assign n34721 = ~controllable_DEQ & ~n22754;
  assign n34722 = ~n22779 & ~n34721;
  assign n34723 = ~i_FULL & ~n34722;
  assign n34724 = ~n22775 & ~n34723;
  assign n34725 = ~i_nEMPTY & ~n34724;
  assign n34726 = ~n22763 & ~n34725;
  assign n34727 = controllable_BtoS_ACK0 & ~n34726;
  assign n34728 = ~controllable_DEQ & ~n22794;
  assign n34729 = ~n22831 & ~n34728;
  assign n34730 = ~i_FULL & ~n34729;
  assign n34731 = ~n22827 & ~n34730;
  assign n34732 = ~i_nEMPTY & ~n34731;
  assign n34733 = ~n22815 & ~n34732;
  assign n34734 = ~controllable_BtoS_ACK0 & ~n34733;
  assign n34735 = ~n34727 & ~n34734;
  assign n34736 = ~n4465 & ~n34735;
  assign n34737 = ~n34720 & ~n34736;
  assign n34738 = ~i_StoB_REQ10 & ~n34737;
  assign n34739 = ~n34704 & ~n34738;
  assign n34740 = controllable_BtoS_ACK10 & ~n34739;
  assign n34741 = ~n23037 & ~n34738;
  assign n34742 = ~controllable_BtoS_ACK10 & ~n34741;
  assign n34743 = ~n34740 & ~n34742;
  assign n34744 = ~n4464 & ~n34743;
  assign n34745 = ~n34684 & ~n34744;
  assign n34746 = ~n4463 & ~n34745;
  assign n34747 = ~n34617 & ~n34746;
  assign n34748 = n4462 & ~n34747;
  assign n34749 = ~controllable_DEQ & ~n23050;
  assign n34750 = ~n23073 & ~n34749;
  assign n34751 = ~i_FULL & ~n34750;
  assign n34752 = ~n23069 & ~n34751;
  assign n34753 = ~i_nEMPTY & ~n34752;
  assign n34754 = ~n23059 & ~n34753;
  assign n34755 = controllable_BtoS_ACK0 & ~n34754;
  assign n34756 = ~n34511 & ~n34755;
  assign n34757 = n4465 & ~n34756;
  assign n34758 = ~n34513 & ~n34757;
  assign n34759 = i_StoB_REQ10 & ~n34758;
  assign n34760 = ~controllable_DEQ & ~n23092;
  assign n34761 = ~n23117 & ~n34760;
  assign n34762 = ~i_FULL & ~n34761;
  assign n34763 = ~n23113 & ~n34762;
  assign n34764 = ~i_nEMPTY & ~n34763;
  assign n34765 = ~n23101 & ~n34764;
  assign n34766 = controllable_BtoS_ACK0 & ~n34765;
  assign n34767 = ~controllable_DEQ & ~n23132;
  assign n34768 = ~n23157 & ~n34767;
  assign n34769 = ~i_FULL & ~n34768;
  assign n34770 = ~n23153 & ~n34769;
  assign n34771 = ~i_nEMPTY & ~n34770;
  assign n34772 = ~n23141 & ~n34771;
  assign n34773 = ~controllable_BtoS_ACK0 & ~n34772;
  assign n34774 = ~n34766 & ~n34773;
  assign n34775 = ~i_StoB_REQ10 & ~n34774;
  assign n34776 = ~n34759 & ~n34775;
  assign n34777 = controllable_BtoS_ACK10 & ~n34776;
  assign n34778 = ~controllable_DEQ & ~n23288;
  assign n34779 = ~n23329 & ~n34778;
  assign n34780 = ~i_FULL & ~n34779;
  assign n34781 = ~n23325 & ~n34780;
  assign n34782 = ~i_nEMPTY & ~n34781;
  assign n34783 = ~n23313 & ~n34782;
  assign n34784 = controllable_BtoS_ACK0 & ~n34783;
  assign n34785 = ~controllable_DEQ & ~n23344;
  assign n34786 = ~n23385 & ~n34785;
  assign n34787 = ~i_FULL & ~n34786;
  assign n34788 = ~n23381 & ~n34787;
  assign n34789 = ~i_nEMPTY & ~n34788;
  assign n34790 = ~n23369 & ~n34789;
  assign n34791 = ~controllable_BtoS_ACK0 & ~n34790;
  assign n34792 = ~n34784 & ~n34791;
  assign n34793 = n4465 & ~n34792;
  assign n34794 = ~n34547 & ~n34793;
  assign n34795 = ~i_StoB_REQ10 & ~n34794;
  assign n34796 = ~n23283 & ~n34795;
  assign n34797 = ~controllable_BtoS_ACK10 & ~n34796;
  assign n34798 = ~n34777 & ~n34797;
  assign n34799 = n4464 & ~n34798;
  assign n34800 = ~n34575 & ~n34775;
  assign n34801 = controllable_BtoS_ACK10 & ~n34800;
  assign n34802 = ~n23517 & ~n34609;
  assign n34803 = ~controllable_BtoS_ACK10 & ~n34802;
  assign n34804 = ~n34801 & ~n34803;
  assign n34805 = ~n4464 & ~n34804;
  assign n34806 = ~n34799 & ~n34805;
  assign n34807 = n4463 & ~n34806;
  assign n34808 = ~controllable_DEQ & ~n23528;
  assign n34809 = ~n23551 & ~n34808;
  assign n34810 = ~i_FULL & ~n34809;
  assign n34811 = ~n23547 & ~n34810;
  assign n34812 = ~i_nEMPTY & ~n34811;
  assign n34813 = ~n23537 & ~n34812;
  assign n34814 = controllable_BtoS_ACK0 & ~n34813;
  assign n34815 = ~controllable_DEQ & ~n23566;
  assign n34816 = ~n23589 & ~n34815;
  assign n34817 = ~i_FULL & ~n34816;
  assign n34818 = ~n23585 & ~n34817;
  assign n34819 = ~i_nEMPTY & ~n34818;
  assign n34820 = ~n23575 & ~n34819;
  assign n34821 = ~controllable_BtoS_ACK0 & ~n34820;
  assign n34822 = ~n34814 & ~n34821;
  assign n34823 = n4465 & ~n34822;
  assign n34824 = ~controllable_DEQ & ~n22102;
  assign n34825 = ~n22125 & ~n34824;
  assign n34826 = ~i_FULL & ~n34825;
  assign n34827 = ~n23609 & ~n34826;
  assign n34828 = ~i_nEMPTY & ~n34827;
  assign n34829 = ~n23605 & ~n34828;
  assign n34830 = ~controllable_BtoS_ACK0 & ~n34829;
  assign n34831 = ~n34504 & ~n34830;
  assign n34832 = ~n4465 & ~n34831;
  assign n34833 = ~n34823 & ~n34832;
  assign n34834 = i_StoB_REQ10 & ~n34833;
  assign n34835 = ~n34775 & ~n34834;
  assign n34836 = controllable_BtoS_ACK10 & ~n34835;
  assign n34837 = ~controllable_DEQ & ~n23732;
  assign n34838 = ~n23769 & ~n34837;
  assign n34839 = ~i_FULL & ~n34838;
  assign n34840 = ~n23765 & ~n34839;
  assign n34841 = ~i_nEMPTY & ~n34840;
  assign n34842 = ~n23753 & ~n34841;
  assign n34843 = controllable_BtoS_ACK0 & ~n34842;
  assign n34844 = ~controllable_DEQ & ~n23784;
  assign n34845 = ~n23821 & ~n34844;
  assign n34846 = ~i_FULL & ~n34845;
  assign n34847 = ~n23817 & ~n34846;
  assign n34848 = ~i_nEMPTY & ~n34847;
  assign n34849 = ~n23805 & ~n34848;
  assign n34850 = ~controllable_BtoS_ACK0 & ~n34849;
  assign n34851 = ~n34843 & ~n34850;
  assign n34852 = n4465 & ~n34851;
  assign n34853 = ~controllable_DEQ & ~n23838;
  assign n34854 = ~n23859 & ~n34853;
  assign n34855 = ~i_FULL & ~n34854;
  assign n34856 = ~n23855 & ~n34855;
  assign n34857 = ~i_nEMPTY & ~n34856;
  assign n34858 = ~n23845 & ~n34857;
  assign n34859 = controllable_BtoS_ACK0 & ~n34858;
  assign n34860 = ~n34674 & ~n34859;
  assign n34861 = ~n4465 & ~n34860;
  assign n34862 = ~n34852 & ~n34861;
  assign n34863 = ~i_StoB_REQ10 & ~n34862;
  assign n34864 = ~n23727 & ~n34863;
  assign n34865 = ~controllable_BtoS_ACK10 & ~n34864;
  assign n34866 = ~n34836 & ~n34865;
  assign n34867 = n4464 & ~n34866;
  assign n34868 = ~controllable_DEQ & ~n22554;
  assign n34869 = ~n22577 & ~n34868;
  assign n34870 = ~i_FULL & ~n34869;
  assign n34871 = ~n23887 & ~n34870;
  assign n34872 = ~i_nEMPTY & ~n34871;
  assign n34873 = ~n23881 & ~n34872;
  assign n34874 = controllable_BtoS_ACK0 & ~n34873;
  assign n34875 = ~controllable_DEQ & ~n22604;
  assign n34876 = ~n22627 & ~n34875;
  assign n34877 = ~i_FULL & ~n34876;
  assign n34878 = ~n23909 & ~n34877;
  assign n34879 = ~i_nEMPTY & ~n34878;
  assign n34880 = ~n23903 & ~n34879;
  assign n34881 = ~controllable_BtoS_ACK0 & ~n34880;
  assign n34882 = ~n34874 & ~n34881;
  assign n34883 = n4465 & ~n34882;
  assign n34884 = ~n34504 & ~n34881;
  assign n34885 = ~n4465 & ~n34884;
  assign n34886 = ~n34883 & ~n34885;
  assign n34887 = i_StoB_REQ10 & ~n34886;
  assign n34888 = ~n34775 & ~n34887;
  assign n34889 = controllable_BtoS_ACK10 & ~n34888;
  assign n34890 = ~controllable_DEQ & ~n24036;
  assign n34891 = ~n24067 & ~n34890;
  assign n34892 = ~i_FULL & ~n34891;
  assign n34893 = ~n24063 & ~n34892;
  assign n34894 = ~i_nEMPTY & ~n34893;
  assign n34895 = ~n24053 & ~n34894;
  assign n34896 = controllable_BtoS_ACK0 & ~n34895;
  assign n34897 = ~controllable_DEQ & ~n24080;
  assign n34898 = ~n24111 & ~n34897;
  assign n34899 = ~i_FULL & ~n34898;
  assign n34900 = ~n24107 & ~n34899;
  assign n34901 = ~i_nEMPTY & ~n34900;
  assign n34902 = ~n24097 & ~n34901;
  assign n34903 = ~controllable_BtoS_ACK0 & ~n34902;
  assign n34904 = ~n34896 & ~n34903;
  assign n34905 = n4465 & ~n34904;
  assign n34906 = ~n34736 & ~n34905;
  assign n34907 = ~i_StoB_REQ10 & ~n34906;
  assign n34908 = ~n24031 & ~n34907;
  assign n34909 = ~controllable_BtoS_ACK10 & ~n34908;
  assign n34910 = ~n34889 & ~n34909;
  assign n34911 = ~n4464 & ~n34910;
  assign n34912 = ~n34867 & ~n34911;
  assign n34913 = ~n4463 & ~n34912;
  assign n34914 = ~n34807 & ~n34913;
  assign n34915 = ~n4462 & ~n34914;
  assign n34916 = ~n34748 & ~n34915;
  assign n34917 = n4461 & ~n34916;
  assign n34918 = ~controllable_DEQ & ~n24138;
  assign n34919 = ~n20925 & ~n34918;
  assign n34920 = ~i_FULL & ~n34919;
  assign n34921 = ~n24149 & ~n34920;
  assign n34922 = ~i_nEMPTY & ~n34921;
  assign n34923 = ~n24145 & ~n34922;
  assign n34924 = controllable_BtoS_ACK0 & ~n34923;
  assign n34925 = ~controllable_DEQ & ~n24164;
  assign n34926 = ~n20963 & ~n34925;
  assign n34927 = ~i_FULL & ~n34926;
  assign n34928 = ~n24175 & ~n34927;
  assign n34929 = ~i_nEMPTY & ~n34928;
  assign n34930 = ~n24171 & ~n34929;
  assign n34931 = ~controllable_BtoS_ACK0 & ~n34930;
  assign n34932 = ~n34924 & ~n34931;
  assign n34933 = n4465 & ~n34932;
  assign n34934 = ~controllable_DEQ & ~n24192;
  assign n34935 = ~n21041 & ~n34934;
  assign n34936 = ~i_FULL & ~n34935;
  assign n34937 = ~n24203 & ~n34936;
  assign n34938 = ~i_nEMPTY & ~n34937;
  assign n34939 = ~n24199 & ~n34938;
  assign n34940 = ~controllable_BtoS_ACK0 & ~n34939;
  assign n34941 = ~n34504 & ~n34940;
  assign n34942 = ~n4465 & ~n34941;
  assign n34943 = ~n34933 & ~n34942;
  assign n34944 = i_StoB_REQ10 & ~n34943;
  assign n34945 = ~controllable_DEQ & ~n24222;
  assign n34946 = ~n21101 & ~n34945;
  assign n34947 = ~i_FULL & ~n34946;
  assign n34948 = ~n24251 & ~n34947;
  assign n34949 = ~i_nEMPTY & ~n34948;
  assign n34950 = ~n24243 & ~n34949;
  assign n34951 = controllable_BtoS_ACK0 & ~n34950;
  assign n34952 = ~controllable_DEQ & ~n24266;
  assign n34953 = ~n21157 & ~n34952;
  assign n34954 = ~i_FULL & ~n34953;
  assign n34955 = ~n24295 & ~n34954;
  assign n34956 = ~i_nEMPTY & ~n34955;
  assign n34957 = ~n24287 & ~n34956;
  assign n34958 = ~controllable_BtoS_ACK0 & ~n34957;
  assign n34959 = ~n34951 & ~n34958;
  assign n34960 = n4465 & ~n34959;
  assign n34961 = ~controllable_DEQ & ~n24312;
  assign n34962 = ~n21199 & ~n34961;
  assign n34963 = ~i_FULL & ~n34962;
  assign n34964 = ~n24329 & ~n34963;
  assign n34965 = ~i_nEMPTY & ~n34964;
  assign n34966 = ~n24321 & ~n34965;
  assign n34967 = controllable_BtoS_ACK0 & ~n34966;
  assign n34968 = ~controllable_DEQ & ~n24344;
  assign n34969 = ~n21255 & ~n34968;
  assign n34970 = ~i_FULL & ~n34969;
  assign n34971 = ~n24373 & ~n34970;
  assign n34972 = ~i_nEMPTY & ~n34971;
  assign n34973 = ~n24365 & ~n34972;
  assign n34974 = ~controllable_BtoS_ACK0 & ~n34973;
  assign n34975 = ~n34967 & ~n34974;
  assign n34976 = ~n4465 & ~n34975;
  assign n34977 = ~n34960 & ~n34976;
  assign n34978 = ~i_StoB_REQ10 & ~n34977;
  assign n34979 = ~n34944 & ~n34978;
  assign n34980 = controllable_BtoS_ACK10 & ~n34979;
  assign n34981 = ~n24547 & ~n34978;
  assign n34982 = ~controllable_BtoS_ACK10 & ~n34981;
  assign n34983 = ~n34980 & ~n34982;
  assign n34984 = n4464 & ~n34983;
  assign n34985 = ~controllable_DEQ & ~n24556;
  assign n34986 = ~n21505 & ~n34985;
  assign n34987 = ~i_FULL & ~n34986;
  assign n34988 = ~n24567 & ~n34987;
  assign n34989 = ~i_nEMPTY & ~n34988;
  assign n34990 = ~n24563 & ~n34989;
  assign n34991 = controllable_BtoS_ACK0 & ~n34990;
  assign n34992 = ~controllable_DEQ & ~n24582;
  assign n34993 = ~n21543 & ~n34992;
  assign n34994 = ~i_FULL & ~n34993;
  assign n34995 = ~n24593 & ~n34994;
  assign n34996 = ~i_nEMPTY & ~n34995;
  assign n34997 = ~n24589 & ~n34996;
  assign n34998 = ~controllable_BtoS_ACK0 & ~n34997;
  assign n34999 = ~n34991 & ~n34998;
  assign n35000 = n4465 & ~n34999;
  assign n35001 = ~n34504 & ~n34998;
  assign n35002 = ~n4465 & ~n35001;
  assign n35003 = ~n35000 & ~n35002;
  assign n35004 = i_StoB_REQ10 & ~n35003;
  assign n35005 = ~controllable_DEQ & ~n24614;
  assign n35006 = ~n21605 & ~n35005;
  assign n35007 = ~i_FULL & ~n35006;
  assign n35008 = ~n24643 & ~n35007;
  assign n35009 = ~i_nEMPTY & ~n35008;
  assign n35010 = ~n24635 & ~n35009;
  assign n35011 = controllable_BtoS_ACK0 & ~n35010;
  assign n35012 = ~controllable_DEQ & ~n24658;
  assign n35013 = ~n21661 & ~n35012;
  assign n35014 = ~i_FULL & ~n35013;
  assign n35015 = ~n24687 & ~n35014;
  assign n35016 = ~i_nEMPTY & ~n35015;
  assign n35017 = ~n24679 & ~n35016;
  assign n35018 = ~controllable_BtoS_ACK0 & ~n35017;
  assign n35019 = ~n35011 & ~n35018;
  assign n35020 = n4465 & ~n35019;
  assign n35021 = ~controllable_DEQ & ~n24704;
  assign n35022 = ~n21703 & ~n35021;
  assign n35023 = ~i_FULL & ~n35022;
  assign n35024 = ~n24721 & ~n35023;
  assign n35025 = ~i_nEMPTY & ~n35024;
  assign n35026 = ~n24713 & ~n35025;
  assign n35027 = controllable_BtoS_ACK0 & ~n35026;
  assign n35028 = ~controllable_DEQ & ~n24736;
  assign n35029 = ~n21759 & ~n35028;
  assign n35030 = ~i_FULL & ~n35029;
  assign n35031 = ~n24765 & ~n35030;
  assign n35032 = ~i_nEMPTY & ~n35031;
  assign n35033 = ~n24757 & ~n35032;
  assign n35034 = ~controllable_BtoS_ACK0 & ~n35033;
  assign n35035 = ~n35027 & ~n35034;
  assign n35036 = ~n4465 & ~n35035;
  assign n35037 = ~n35020 & ~n35036;
  assign n35038 = ~i_StoB_REQ10 & ~n35037;
  assign n35039 = ~n35004 & ~n35038;
  assign n35040 = controllable_BtoS_ACK10 & ~n35039;
  assign n35041 = ~n24939 & ~n35038;
  assign n35042 = ~controllable_BtoS_ACK10 & ~n35041;
  assign n35043 = ~n35040 & ~n35042;
  assign n35044 = ~n4464 & ~n35043;
  assign n35045 = ~n34984 & ~n35044;
  assign n35046 = n4463 & ~n35045;
  assign n35047 = ~controllable_DEQ & ~n24948;
  assign n35048 = ~n22181 & ~n35047;
  assign n35049 = ~i_FULL & ~n35048;
  assign n35050 = ~n24969 & ~n35049;
  assign n35051 = ~i_nEMPTY & ~n35050;
  assign n35052 = ~n24963 & ~n35051;
  assign n35053 = controllable_BtoS_ACK0 & ~n35052;
  assign n35054 = ~controllable_DEQ & ~n24980;
  assign n35055 = ~n22233 & ~n35054;
  assign n35056 = ~i_FULL & ~n35055;
  assign n35057 = ~n25001 & ~n35056;
  assign n35058 = ~i_nEMPTY & ~n35057;
  assign n35059 = ~n24995 & ~n35058;
  assign n35060 = ~controllable_BtoS_ACK0 & ~n35059;
  assign n35061 = ~n35053 & ~n35060;
  assign n35062 = n4465 & ~n35061;
  assign n35063 = ~controllable_DEQ & ~n25014;
  assign n35064 = ~n22275 & ~n35063;
  assign n35065 = ~i_FULL & ~n35064;
  assign n35066 = ~n25027 & ~n35065;
  assign n35067 = ~i_nEMPTY & ~n35066;
  assign n35068 = ~n25021 & ~n35067;
  assign n35069 = controllable_BtoS_ACK0 & ~n35068;
  assign n35070 = ~n34674 & ~n35069;
  assign n35071 = ~n4465 & ~n35070;
  assign n35072 = ~n35062 & ~n35071;
  assign n35073 = ~i_StoB_REQ10 & ~n35072;
  assign n35074 = ~n34644 & ~n35073;
  assign n35075 = controllable_BtoS_ACK10 & ~n35074;
  assign n35076 = ~n22533 & ~n35073;
  assign n35077 = ~controllable_BtoS_ACK10 & ~n35076;
  assign n35078 = ~n35075 & ~n35077;
  assign n35079 = n4464 & ~n35078;
  assign n35080 = ~controllable_DEQ & ~n25048;
  assign n35081 = ~n22685 & ~n35080;
  assign n35082 = ~i_FULL & ~n35081;
  assign n35083 = ~n25069 & ~n35082;
  assign n35084 = ~i_nEMPTY & ~n35083;
  assign n35085 = ~n25063 & ~n35084;
  assign n35086 = controllable_BtoS_ACK0 & ~n35085;
  assign n35087 = ~controllable_DEQ & ~n25080;
  assign n35088 = ~n22737 & ~n35087;
  assign n35089 = ~i_FULL & ~n35088;
  assign n35090 = ~n25101 & ~n35089;
  assign n35091 = ~i_nEMPTY & ~n35090;
  assign n35092 = ~n25095 & ~n35091;
  assign n35093 = ~controllable_BtoS_ACK0 & ~n35092;
  assign n35094 = ~n35086 & ~n35093;
  assign n35095 = n4465 & ~n35094;
  assign n35096 = ~n34736 & ~n35095;
  assign n35097 = ~i_StoB_REQ10 & ~n35096;
  assign n35098 = ~n34704 & ~n35097;
  assign n35099 = controllable_BtoS_ACK10 & ~n35098;
  assign n35100 = ~n23037 & ~n35097;
  assign n35101 = ~controllable_BtoS_ACK10 & ~n35100;
  assign n35102 = ~n35099 & ~n35101;
  assign n35103 = ~n4464 & ~n35102;
  assign n35104 = ~n35079 & ~n35103;
  assign n35105 = ~n4463 & ~n35104;
  assign n35106 = ~n35046 & ~n35105;
  assign n35107 = n4462 & ~n35106;
  assign n35108 = ~controllable_DEQ & ~n25128;
  assign n35109 = ~n23073 & ~n35108;
  assign n35110 = ~i_FULL & ~n35109;
  assign n35111 = ~n25143 & ~n35110;
  assign n35112 = ~i_nEMPTY & ~n35111;
  assign n35113 = ~n25137 & ~n35112;
  assign n35114 = controllable_BtoS_ACK0 & ~n35113;
  assign n35115 = ~controllable_DEQ & ~n25156;
  assign n35116 = ~n21041 & ~n35115;
  assign n35117 = ~i_FULL & ~n35116;
  assign n35118 = ~n25169 & ~n35117;
  assign n35119 = ~i_nEMPTY & ~n35118;
  assign n35120 = ~n25163 & ~n35119;
  assign n35121 = ~controllable_BtoS_ACK0 & ~n35120;
  assign n35122 = ~n35114 & ~n35121;
  assign n35123 = n4465 & ~n35122;
  assign n35124 = ~n34942 & ~n35123;
  assign n35125 = i_StoB_REQ10 & ~n35124;
  assign n35126 = ~n34775 & ~n35125;
  assign n35127 = controllable_BtoS_ACK10 & ~n35126;
  assign n35128 = ~controllable_DEQ & ~n25278;
  assign n35129 = ~n23329 & ~n35128;
  assign n35130 = ~i_FULL & ~n35129;
  assign n35131 = ~n25307 & ~n35130;
  assign n35132 = ~i_nEMPTY & ~n35131;
  assign n35133 = ~n25299 & ~n35132;
  assign n35134 = controllable_BtoS_ACK0 & ~n35133;
  assign n35135 = ~controllable_DEQ & ~n25322;
  assign n35136 = ~n23385 & ~n35135;
  assign n35137 = ~i_FULL & ~n35136;
  assign n35138 = ~n25351 & ~n35137;
  assign n35139 = ~i_nEMPTY & ~n35138;
  assign n35140 = ~n25343 & ~n35139;
  assign n35141 = ~controllable_BtoS_ACK0 & ~n35140;
  assign n35142 = ~n35134 & ~n35141;
  assign n35143 = n4465 & ~n35142;
  assign n35144 = ~controllable_DEQ & ~n25366;
  assign n35145 = ~n21199 & ~n35144;
  assign n35146 = ~i_FULL & ~n35145;
  assign n35147 = ~n25379 & ~n35146;
  assign n35148 = ~i_nEMPTY & ~n35147;
  assign n35149 = ~n25373 & ~n35148;
  assign n35150 = controllable_BtoS_ACK0 & ~n35149;
  assign n35151 = ~n34974 & ~n35150;
  assign n35152 = ~n4465 & ~n35151;
  assign n35153 = ~n35143 & ~n35152;
  assign n35154 = ~i_StoB_REQ10 & ~n35153;
  assign n35155 = ~n25273 & ~n35154;
  assign n35156 = ~controllable_BtoS_ACK10 & ~n35155;
  assign n35157 = ~n35127 & ~n35156;
  assign n35158 = n4464 & ~n35157;
  assign n35159 = ~n34775 & ~n35004;
  assign n35160 = controllable_BtoS_ACK10 & ~n35159;
  assign n35161 = ~controllable_DEQ & ~n25490;
  assign n35162 = ~n21605 & ~n35161;
  assign n35163 = ~i_FULL & ~n35162;
  assign n35164 = ~n25515 & ~n35163;
  assign n35165 = ~i_nEMPTY & ~n35164;
  assign n35166 = ~n25509 & ~n35165;
  assign n35167 = controllable_BtoS_ACK0 & ~n35166;
  assign n35168 = ~controllable_DEQ & ~n25528;
  assign n35169 = ~n21661 & ~n35168;
  assign n35170 = ~i_FULL & ~n35169;
  assign n35171 = ~n25553 & ~n35170;
  assign n35172 = ~i_nEMPTY & ~n35171;
  assign n35173 = ~n25547 & ~n35172;
  assign n35174 = ~controllable_BtoS_ACK0 & ~n35173;
  assign n35175 = ~n35167 & ~n35174;
  assign n35176 = n4465 & ~n35175;
  assign n35177 = ~n35036 & ~n35176;
  assign n35178 = ~i_StoB_REQ10 & ~n35177;
  assign n35179 = ~n25487 & ~n35178;
  assign n35180 = ~controllable_BtoS_ACK10 & ~n35179;
  assign n35181 = ~n35160 & ~n35180;
  assign n35182 = ~n4464 & ~n35181;
  assign n35183 = ~n35158 & ~n35182;
  assign n35184 = n4463 & ~n35183;
  assign n35185 = ~controllable_DEQ & ~n25576;
  assign n35186 = ~n23551 & ~n35185;
  assign n35187 = ~i_FULL & ~n35186;
  assign n35188 = ~n25587 & ~n35187;
  assign n35189 = ~i_nEMPTY & ~n35188;
  assign n35190 = ~n25583 & ~n35189;
  assign n35191 = controllable_BtoS_ACK0 & ~n35190;
  assign n35192 = ~controllable_DEQ & ~n25598;
  assign n35193 = ~n23589 & ~n35192;
  assign n35194 = ~i_FULL & ~n35193;
  assign n35195 = ~n25609 & ~n35194;
  assign n35196 = ~i_nEMPTY & ~n35195;
  assign n35197 = ~n25605 & ~n35196;
  assign n35198 = ~controllable_BtoS_ACK0 & ~n35197;
  assign n35199 = ~n35191 & ~n35198;
  assign n35200 = n4465 & ~n35199;
  assign n35201 = ~n34832 & ~n35200;
  assign n35202 = i_StoB_REQ10 & ~n35201;
  assign n35203 = ~n34775 & ~n35202;
  assign n35204 = controllable_BtoS_ACK10 & ~n35203;
  assign n35205 = ~n34865 & ~n35204;
  assign n35206 = n4464 & ~n35205;
  assign n35207 = ~n34911 & ~n35206;
  assign n35208 = ~n4463 & ~n35207;
  assign n35209 = ~n35184 & ~n35208;
  assign n35210 = ~n4462 & ~n35209;
  assign n35211 = ~n35107 & ~n35210;
  assign n35212 = ~n4461 & ~n35211;
  assign n35213 = ~n34917 & ~n35212;
  assign n35214 = ~n4459 & ~n35213;
  assign n35215 = ~controllable_DEQ & ~n25640;
  assign n35216 = ~n21101 & ~n35215;
  assign n35217 = ~i_FULL & ~n35216;
  assign n35218 = ~n25671 & ~n35217;
  assign n35219 = ~i_nEMPTY & ~n35218;
  assign n35220 = ~n25663 & ~n35219;
  assign n35221 = controllable_BtoS_ACK0 & ~n35220;
  assign n35222 = ~controllable_DEQ & ~n25690;
  assign n35223 = ~n21157 & ~n35222;
  assign n35224 = ~i_FULL & ~n35223;
  assign n35225 = ~n25721 & ~n35224;
  assign n35226 = ~i_nEMPTY & ~n35225;
  assign n35227 = ~n25713 & ~n35226;
  assign n35228 = ~controllable_BtoS_ACK0 & ~n35227;
  assign n35229 = ~n35221 & ~n35228;
  assign n35230 = n4465 & ~n35229;
  assign n35231 = ~controllable_DEQ & ~n25738;
  assign n35232 = ~n21199 & ~n35231;
  assign n35233 = ~i_FULL & ~n35232;
  assign n35234 = ~n25751 & ~n35233;
  assign n35235 = ~i_nEMPTY & ~n35234;
  assign n35236 = ~n25745 & ~n35235;
  assign n35237 = controllable_BtoS_ACK0 & ~n35236;
  assign n35238 = ~n34974 & ~n35237;
  assign n35239 = ~n4465 & ~n35238;
  assign n35240 = ~n35230 & ~n35239;
  assign n35241 = ~i_StoB_REQ10 & ~n35240;
  assign n35242 = ~n34944 & ~n35241;
  assign n35243 = controllable_BtoS_ACK10 & ~n35242;
  assign n35244 = ~n24547 & ~n35241;
  assign n35245 = ~controllable_BtoS_ACK10 & ~n35244;
  assign n35246 = ~n35243 & ~n35245;
  assign n35247 = n4464 & ~n35246;
  assign n35248 = ~controllable_DEQ & ~n25772;
  assign n35249 = ~n21605 & ~n35248;
  assign n35250 = ~i_FULL & ~n35249;
  assign n35251 = ~n25793 & ~n35250;
  assign n35252 = ~i_nEMPTY & ~n35251;
  assign n35253 = ~n25787 & ~n35252;
  assign n35254 = controllable_BtoS_ACK0 & ~n35253;
  assign n35255 = ~controllable_DEQ & ~n25804;
  assign n35256 = ~n21661 & ~n35255;
  assign n35257 = ~i_FULL & ~n35256;
  assign n35258 = ~n25825 & ~n35257;
  assign n35259 = ~i_nEMPTY & ~n35258;
  assign n35260 = ~n25819 & ~n35259;
  assign n35261 = ~controllable_BtoS_ACK0 & ~n35260;
  assign n35262 = ~n35254 & ~n35261;
  assign n35263 = n4465 & ~n35262;
  assign n35264 = ~n35036 & ~n35263;
  assign n35265 = ~i_StoB_REQ10 & ~n35264;
  assign n35266 = ~n35004 & ~n35265;
  assign n35267 = controllable_BtoS_ACK10 & ~n35266;
  assign n35268 = ~n24939 & ~n35265;
  assign n35269 = ~controllable_BtoS_ACK10 & ~n35268;
  assign n35270 = ~n35267 & ~n35269;
  assign n35271 = ~n4464 & ~n35270;
  assign n35272 = ~n35247 & ~n35271;
  assign n35273 = ~n4463 & ~n35272;
  assign n35274 = ~n34617 & ~n35273;
  assign n35275 = n4462 & ~n35274;
  assign n35276 = ~controllable_DEQ & ~n25854;
  assign n35277 = ~n23073 & ~n35276;
  assign n35278 = ~i_FULL & ~n35277;
  assign n35279 = ~n25873 & ~n35278;
  assign n35280 = ~i_nEMPTY & ~n35279;
  assign n35281 = ~n25865 & ~n35280;
  assign n35282 = controllable_BtoS_ACK0 & ~n35281;
  assign n35283 = ~controllable_DEQ & ~n25888;
  assign n35284 = ~n21041 & ~n35283;
  assign n35285 = ~i_FULL & ~n35284;
  assign n35286 = ~n25899 & ~n35285;
  assign n35287 = ~i_nEMPTY & ~n35286;
  assign n35288 = ~n25895 & ~n35287;
  assign n35289 = ~controllable_BtoS_ACK0 & ~n35288;
  assign n35290 = ~n35282 & ~n35289;
  assign n35291 = n4465 & ~n35290;
  assign n35292 = ~n34942 & ~n35291;
  assign n35293 = i_StoB_REQ10 & ~n35292;
  assign n35294 = ~n34775 & ~n35293;
  assign n35295 = controllable_BtoS_ACK10 & ~n35294;
  assign n35296 = ~n35156 & ~n35295;
  assign n35297 = n4464 & ~n35296;
  assign n35298 = ~n35182 & ~n35297;
  assign n35299 = ~n4463 & ~n35298;
  assign n35300 = ~n34807 & ~n35299;
  assign n35301 = ~n4462 & ~n35300;
  assign n35302 = ~n35275 & ~n35301;
  assign n35303 = n4461 & ~n35302;
  assign n35304 = ~controllable_DEQ & ~n25926;
  assign n35305 = ~n22023 & ~n35304;
  assign n35306 = ~i_FULL & ~n35305;
  assign n35307 = ~n25957 & ~n35306;
  assign n35308 = ~i_nEMPTY & ~n35307;
  assign n35309 = ~n25950 & ~n35308;
  assign n35310 = controllable_BtoS_ACK0 & ~n35309;
  assign n35311 = ~controllable_DEQ & ~n25974;
  assign n35312 = ~n22073 & ~n35311;
  assign n35313 = ~i_FULL & ~n35312;
  assign n35314 = ~n26005 & ~n35313;
  assign n35315 = ~i_nEMPTY & ~n35314;
  assign n35316 = ~n25998 & ~n35315;
  assign n35317 = ~controllable_BtoS_ACK0 & ~n35316;
  assign n35318 = ~n35310 & ~n35317;
  assign n35319 = n4465 & ~n35318;
  assign n35320 = ~controllable_DEQ & ~n26024;
  assign n35321 = ~n22125 & ~n35320;
  assign n35322 = ~i_FULL & ~n35321;
  assign n35323 = ~n26055 & ~n35322;
  assign n35324 = ~i_nEMPTY & ~n35323;
  assign n35325 = ~n26048 & ~n35324;
  assign n35326 = ~controllable_BtoS_ACK0 & ~n35325;
  assign n35327 = ~n34504 & ~n35326;
  assign n35328 = ~n4465 & ~n35327;
  assign n35329 = ~n35319 & ~n35328;
  assign n35330 = i_StoB_REQ10 & ~n35329;
  assign n35331 = ~controllable_DEQ & ~n26076;
  assign n35332 = ~n22181 & ~n35331;
  assign n35333 = ~i_FULL & ~n35332;
  assign n35334 = ~n26109 & ~n35333;
  assign n35335 = ~i_nEMPTY & ~n35334;
  assign n35336 = ~n26101 & ~n35335;
  assign n35337 = controllable_BtoS_ACK0 & ~n35336;
  assign n35338 = ~controllable_DEQ & ~n26126;
  assign n35339 = ~n22233 & ~n35338;
  assign n35340 = ~i_FULL & ~n35339;
  assign n35341 = ~n26159 & ~n35340;
  assign n35342 = ~i_nEMPTY & ~n35341;
  assign n35343 = ~n26151 & ~n35342;
  assign n35344 = ~controllable_BtoS_ACK0 & ~n35343;
  assign n35345 = ~n35337 & ~n35344;
  assign n35346 = n4465 & ~n35345;
  assign n35347 = ~controllable_DEQ & ~n26178;
  assign n35348 = ~n22275 & ~n35347;
  assign n35349 = ~i_FULL & ~n35348;
  assign n35350 = ~n26195 & ~n35349;
  assign n35351 = ~i_nEMPTY & ~n35350;
  assign n35352 = ~n26187 & ~n35351;
  assign n35353 = controllable_BtoS_ACK0 & ~n35352;
  assign n35354 = ~controllable_DEQ & ~n26212;
  assign n35355 = ~n22327 & ~n35354;
  assign n35356 = ~i_FULL & ~n35355;
  assign n35357 = ~n26245 & ~n35356;
  assign n35358 = ~i_nEMPTY & ~n35357;
  assign n35359 = ~n26237 & ~n35358;
  assign n35360 = ~controllable_BtoS_ACK0 & ~n35359;
  assign n35361 = ~n35353 & ~n35360;
  assign n35362 = ~n4465 & ~n35361;
  assign n35363 = ~n35346 & ~n35362;
  assign n35364 = ~i_StoB_REQ10 & ~n35363;
  assign n35365 = ~n35330 & ~n35364;
  assign n35366 = controllable_BtoS_ACK10 & ~n35365;
  assign n35367 = ~n26427 & ~n35364;
  assign n35368 = ~controllable_BtoS_ACK10 & ~n35367;
  assign n35369 = ~n35366 & ~n35368;
  assign n35370 = n4464 & ~n35369;
  assign n35371 = ~controllable_DEQ & ~n26436;
  assign n35372 = ~n22577 & ~n35371;
  assign n35373 = ~i_FULL & ~n35372;
  assign n35374 = ~n26467 & ~n35373;
  assign n35375 = ~i_nEMPTY & ~n35374;
  assign n35376 = ~n26460 & ~n35375;
  assign n35377 = controllable_BtoS_ACK0 & ~n35376;
  assign n35378 = ~controllable_DEQ & ~n26484;
  assign n35379 = ~n22627 & ~n35378;
  assign n35380 = ~i_FULL & ~n35379;
  assign n35381 = ~n26515 & ~n35380;
  assign n35382 = ~i_nEMPTY & ~n35381;
  assign n35383 = ~n26508 & ~n35382;
  assign n35384 = ~controllable_BtoS_ACK0 & ~n35383;
  assign n35385 = ~n35377 & ~n35384;
  assign n35386 = n4465 & ~n35385;
  assign n35387 = ~n34504 & ~n35384;
  assign n35388 = ~n4465 & ~n35387;
  assign n35389 = ~n35386 & ~n35388;
  assign n35390 = i_StoB_REQ10 & ~n35389;
  assign n35391 = ~controllable_DEQ & ~n26538;
  assign n35392 = ~n22685 & ~n35391;
  assign n35393 = ~i_FULL & ~n35392;
  assign n35394 = ~n26571 & ~n35393;
  assign n35395 = ~i_nEMPTY & ~n35394;
  assign n35396 = ~n26563 & ~n35395;
  assign n35397 = controllable_BtoS_ACK0 & ~n35396;
  assign n35398 = ~controllable_DEQ & ~n26588;
  assign n35399 = ~n22737 & ~n35398;
  assign n35400 = ~i_FULL & ~n35399;
  assign n35401 = ~n26621 & ~n35400;
  assign n35402 = ~i_nEMPTY & ~n35401;
  assign n35403 = ~n26613 & ~n35402;
  assign n35404 = ~controllable_BtoS_ACK0 & ~n35403;
  assign n35405 = ~n35397 & ~n35404;
  assign n35406 = n4465 & ~n35405;
  assign n35407 = ~controllable_DEQ & ~n26640;
  assign n35408 = ~n22779 & ~n35407;
  assign n35409 = ~i_FULL & ~n35408;
  assign n35410 = ~n26657 & ~n35409;
  assign n35411 = ~i_nEMPTY & ~n35410;
  assign n35412 = ~n26649 & ~n35411;
  assign n35413 = controllable_BtoS_ACK0 & ~n35412;
  assign n35414 = ~controllable_DEQ & ~n26674;
  assign n35415 = ~n22831 & ~n35414;
  assign n35416 = ~i_FULL & ~n35415;
  assign n35417 = ~n26707 & ~n35416;
  assign n35418 = ~i_nEMPTY & ~n35417;
  assign n35419 = ~n26699 & ~n35418;
  assign n35420 = ~controllable_BtoS_ACK0 & ~n35419;
  assign n35421 = ~n35413 & ~n35420;
  assign n35422 = ~n4465 & ~n35421;
  assign n35423 = ~n35406 & ~n35422;
  assign n35424 = ~i_StoB_REQ10 & ~n35423;
  assign n35425 = ~n35390 & ~n35424;
  assign n35426 = controllable_BtoS_ACK10 & ~n35425;
  assign n35427 = ~n26881 & ~n35424;
  assign n35428 = ~controllable_BtoS_ACK10 & ~n35427;
  assign n35429 = ~n35426 & ~n35428;
  assign n35430 = ~n4464 & ~n35429;
  assign n35431 = ~n35370 & ~n35430;
  assign n35432 = n4463 & ~n35431;
  assign n35433 = ~controllable_DEQ & ~n26892;
  assign n35434 = ~n22181 & ~n35433;
  assign n35435 = ~i_FULL & ~n35434;
  assign n35436 = ~n26925 & ~n35435;
  assign n35437 = ~i_nEMPTY & ~n35436;
  assign n35438 = ~n26917 & ~n35437;
  assign n35439 = controllable_BtoS_ACK0 & ~n35438;
  assign n35440 = ~controllable_DEQ & ~n26942;
  assign n35441 = ~n22233 & ~n35440;
  assign n35442 = ~i_FULL & ~n35441;
  assign n35443 = ~n26975 & ~n35442;
  assign n35444 = ~i_nEMPTY & ~n35443;
  assign n35445 = ~n26967 & ~n35444;
  assign n35446 = ~controllable_BtoS_ACK0 & ~n35445;
  assign n35447 = ~n35439 & ~n35446;
  assign n35448 = n4465 & ~n35447;
  assign n35449 = ~controllable_DEQ & ~n26994;
  assign n35450 = ~n22275 & ~n35449;
  assign n35451 = ~i_FULL & ~n35450;
  assign n35452 = ~n27011 & ~n35451;
  assign n35453 = ~i_nEMPTY & ~n35452;
  assign n35454 = ~n27003 & ~n35453;
  assign n35455 = controllable_BtoS_ACK0 & ~n35454;
  assign n35456 = ~n35360 & ~n35455;
  assign n35457 = ~n4465 & ~n35456;
  assign n35458 = ~n35448 & ~n35457;
  assign n35459 = ~i_StoB_REQ10 & ~n35458;
  assign n35460 = ~n35330 & ~n35459;
  assign n35461 = controllable_BtoS_ACK10 & ~n35460;
  assign n35462 = ~n26427 & ~n35459;
  assign n35463 = ~controllable_BtoS_ACK10 & ~n35462;
  assign n35464 = ~n35461 & ~n35463;
  assign n35465 = n4464 & ~n35464;
  assign n35466 = ~controllable_DEQ & ~n27038;
  assign n35467 = ~n22685 & ~n35466;
  assign n35468 = ~i_FULL & ~n35467;
  assign n35469 = ~n27071 & ~n35468;
  assign n35470 = ~i_nEMPTY & ~n35469;
  assign n35471 = ~n27063 & ~n35470;
  assign n35472 = controllable_BtoS_ACK0 & ~n35471;
  assign n35473 = ~controllable_DEQ & ~n27088;
  assign n35474 = ~n22737 & ~n35473;
  assign n35475 = ~i_FULL & ~n35474;
  assign n35476 = ~n27121 & ~n35475;
  assign n35477 = ~i_nEMPTY & ~n35476;
  assign n35478 = ~n27113 & ~n35477;
  assign n35479 = ~controllable_BtoS_ACK0 & ~n35478;
  assign n35480 = ~n35472 & ~n35479;
  assign n35481 = n4465 & ~n35480;
  assign n35482 = ~n35422 & ~n35481;
  assign n35483 = ~i_StoB_REQ10 & ~n35482;
  assign n35484 = ~n35390 & ~n35483;
  assign n35485 = controllable_BtoS_ACK10 & ~n35484;
  assign n35486 = ~n26881 & ~n35483;
  assign n35487 = ~controllable_BtoS_ACK10 & ~n35486;
  assign n35488 = ~n35485 & ~n35487;
  assign n35489 = ~n4464 & ~n35488;
  assign n35490 = ~n35465 & ~n35489;
  assign n35491 = ~n4463 & ~n35490;
  assign n35492 = ~n35432 & ~n35491;
  assign n35493 = n4462 & ~n35492;
  assign n35494 = ~controllable_DEQ & ~n27152;
  assign n35495 = ~n23551 & ~n35494;
  assign n35496 = ~i_FULL & ~n35495;
  assign n35497 = ~n27169 & ~n35496;
  assign n35498 = ~i_nEMPTY & ~n35497;
  assign n35499 = ~n27161 & ~n35498;
  assign n35500 = controllable_BtoS_ACK0 & ~n35499;
  assign n35501 = ~controllable_DEQ & ~n27186;
  assign n35502 = ~n23589 & ~n35501;
  assign n35503 = ~i_FULL & ~n35502;
  assign n35504 = ~n27203 & ~n35503;
  assign n35505 = ~i_nEMPTY & ~n35504;
  assign n35506 = ~n27195 & ~n35505;
  assign n35507 = ~controllable_BtoS_ACK0 & ~n35506;
  assign n35508 = ~n35500 & ~n35507;
  assign n35509 = n4465 & ~n35508;
  assign n35510 = ~controllable_DEQ & ~n26037;
  assign n35511 = ~n22125 & ~n35510;
  assign n35512 = ~i_FULL & ~n35511;
  assign n35513 = ~n27233 & ~n35512;
  assign n35514 = ~i_nEMPTY & ~n35513;
  assign n35515 = ~n27225 & ~n35514;
  assign n35516 = ~controllable_BtoS_ACK0 & ~n35515;
  assign n35517 = ~n34504 & ~n35516;
  assign n35518 = ~n4465 & ~n35517;
  assign n35519 = ~n35509 & ~n35518;
  assign n35520 = i_StoB_REQ10 & ~n35519;
  assign n35521 = ~n34775 & ~n35520;
  assign n35522 = controllable_BtoS_ACK10 & ~n35521;
  assign n35523 = ~controllable_DEQ & ~n27348;
  assign n35524 = ~n23769 & ~n35523;
  assign n35525 = ~i_FULL & ~n35524;
  assign n35526 = ~n27377 & ~n35525;
  assign n35527 = ~i_nEMPTY & ~n35526;
  assign n35528 = ~n27371 & ~n35527;
  assign n35529 = controllable_BtoS_ACK0 & ~n35528;
  assign n35530 = ~controllable_DEQ & ~n27394;
  assign n35531 = ~n23821 & ~n35530;
  assign n35532 = ~i_FULL & ~n35531;
  assign n35533 = ~n27423 & ~n35532;
  assign n35534 = ~i_nEMPTY & ~n35533;
  assign n35535 = ~n27417 & ~n35534;
  assign n35536 = ~controllable_BtoS_ACK0 & ~n35535;
  assign n35537 = ~n35529 & ~n35536;
  assign n35538 = n4465 & ~n35537;
  assign n35539 = ~controllable_DEQ & ~n27442;
  assign n35540 = ~n23859 & ~n35539;
  assign n35541 = ~i_FULL & ~n35540;
  assign n35542 = ~n27455 & ~n35541;
  assign n35543 = ~i_nEMPTY & ~n35542;
  assign n35544 = ~n27449 & ~n35543;
  assign n35545 = controllable_BtoS_ACK0 & ~n35544;
  assign n35546 = ~n35360 & ~n35545;
  assign n35547 = ~n4465 & ~n35546;
  assign n35548 = ~n35538 & ~n35547;
  assign n35549 = ~i_StoB_REQ10 & ~n35548;
  assign n35550 = ~n27343 & ~n35549;
  assign n35551 = ~controllable_BtoS_ACK10 & ~n35550;
  assign n35552 = ~n35522 & ~n35551;
  assign n35553 = n4464 & ~n35552;
  assign n35554 = ~controllable_DEQ & ~n26449;
  assign n35555 = ~n22577 & ~n35554;
  assign n35556 = ~i_FULL & ~n35555;
  assign n35557 = ~n27491 & ~n35556;
  assign n35558 = ~i_nEMPTY & ~n35557;
  assign n35559 = ~n27483 & ~n35558;
  assign n35560 = controllable_BtoS_ACK0 & ~n35559;
  assign n35561 = ~controllable_DEQ & ~n26497;
  assign n35562 = ~n22627 & ~n35561;
  assign n35563 = ~i_FULL & ~n35562;
  assign n35564 = ~n27519 & ~n35563;
  assign n35565 = ~i_nEMPTY & ~n35564;
  assign n35566 = ~n27511 & ~n35565;
  assign n35567 = ~controllable_BtoS_ACK0 & ~n35566;
  assign n35568 = ~n35560 & ~n35567;
  assign n35569 = n4465 & ~n35568;
  assign n35570 = ~n34504 & ~n35567;
  assign n35571 = ~n4465 & ~n35570;
  assign n35572 = ~n35569 & ~n35571;
  assign n35573 = i_StoB_REQ10 & ~n35572;
  assign n35574 = ~n34775 & ~n35573;
  assign n35575 = controllable_BtoS_ACK10 & ~n35574;
  assign n35576 = ~controllable_DEQ & ~n27632;
  assign n35577 = ~n24067 & ~n35576;
  assign n35578 = ~i_FULL & ~n35577;
  assign n35579 = ~n27659 & ~n35578;
  assign n35580 = ~i_nEMPTY & ~n35579;
  assign n35581 = ~n27653 & ~n35580;
  assign n35582 = controllable_BtoS_ACK0 & ~n35581;
  assign n35583 = ~controllable_DEQ & ~n27676;
  assign n35584 = ~n24111 & ~n35583;
  assign n35585 = ~i_FULL & ~n35584;
  assign n35586 = ~n27703 & ~n35585;
  assign n35587 = ~i_nEMPTY & ~n35586;
  assign n35588 = ~n27697 & ~n35587;
  assign n35589 = ~controllable_BtoS_ACK0 & ~n35588;
  assign n35590 = ~n35582 & ~n35589;
  assign n35591 = n4465 & ~n35590;
  assign n35592 = ~n35422 & ~n35591;
  assign n35593 = ~i_StoB_REQ10 & ~n35592;
  assign n35594 = ~n27627 & ~n35593;
  assign n35595 = ~controllable_BtoS_ACK10 & ~n35594;
  assign n35596 = ~n35575 & ~n35595;
  assign n35597 = ~n4464 & ~n35596;
  assign n35598 = ~n35553 & ~n35597;
  assign n35599 = n4463 & ~n35598;
  assign n35600 = ~controllable_DEQ & ~n27730;
  assign n35601 = ~n23551 & ~n35600;
  assign n35602 = ~i_FULL & ~n35601;
  assign n35603 = ~n27747 & ~n35602;
  assign n35604 = ~i_nEMPTY & ~n35603;
  assign n35605 = ~n27739 & ~n35604;
  assign n35606 = controllable_BtoS_ACK0 & ~n35605;
  assign n35607 = ~controllable_DEQ & ~n27764;
  assign n35608 = ~n23589 & ~n35607;
  assign n35609 = ~i_FULL & ~n35608;
  assign n35610 = ~n27781 & ~n35609;
  assign n35611 = ~i_nEMPTY & ~n35610;
  assign n35612 = ~n27773 & ~n35611;
  assign n35613 = ~controllable_BtoS_ACK0 & ~n35612;
  assign n35614 = ~n35606 & ~n35613;
  assign n35615 = n4465 & ~n35614;
  assign n35616 = ~n35518 & ~n35615;
  assign n35617 = i_StoB_REQ10 & ~n35616;
  assign n35618 = ~n34775 & ~n35617;
  assign n35619 = controllable_BtoS_ACK10 & ~n35618;
  assign n35620 = ~n35551 & ~n35619;
  assign n35621 = n4464 & ~n35620;
  assign n35622 = ~n35597 & ~n35621;
  assign n35623 = ~n4463 & ~n35622;
  assign n35624 = ~n35599 & ~n35623;
  assign n35625 = ~n4462 & ~n35624;
  assign n35626 = ~n35493 & ~n35625;
  assign n35627 = ~n4461 & ~n35626;
  assign n35628 = ~n35303 & ~n35627;
  assign n35629 = n4459 & ~n35628;
  assign n35630 = ~n35214 & ~n35629;
  assign n35631 = ~n4455 & ~n35630;
  assign n35632 = ~n34481 & ~n35631;
  assign n35633 = n4445 & ~n35632;
  assign n35634 = ~controllable_DEQ & ~n27819;
  assign n35635 = ~n5296 & ~n35634;
  assign n35636 = ~i_FULL & ~n35635;
  assign n35637 = ~n27841 & ~n35636;
  assign n35638 = ~i_nEMPTY & ~n35637;
  assign n35639 = ~n27835 & ~n35638;
  assign n35640 = controllable_BtoS_ACK0 & ~n35639;
  assign n35641 = ~controllable_DEQ & ~n27865;
  assign n35642 = ~n27912 & ~n35641;
  assign n35643 = ~i_FULL & ~n35642;
  assign n35644 = ~n27906 & ~n35643;
  assign n35645 = ~i_nEMPTY & ~n35644;
  assign n35646 = ~n27893 & ~n35645;
  assign n35647 = ~controllable_BtoS_ACK0 & ~n35646;
  assign n35648 = ~n35640 & ~n35647;
  assign n35649 = n4465 & ~n35648;
  assign n35650 = ~controllable_DEQ & ~n27931;
  assign n35651 = ~n27912 & ~n35650;
  assign n35652 = ~i_FULL & ~n35651;
  assign n35653 = ~n27953 & ~n35652;
  assign n35654 = ~i_nEMPTY & ~n35653;
  assign n35655 = ~n27947 & ~n35654;
  assign n35656 = ~controllable_BtoS_ACK0 & ~n35655;
  assign n35657 = ~n33206 & ~n35656;
  assign n35658 = ~n4465 & ~n35657;
  assign n35659 = ~n35649 & ~n35658;
  assign n35660 = i_StoB_REQ10 & ~n35659;
  assign n35661 = ~controllable_DEQ & ~n27975;
  assign n35662 = ~n11282 & ~n35661;
  assign n35663 = ~i_FULL & ~n35662;
  assign n35664 = ~n27999 & ~n35663;
  assign n35665 = ~i_nEMPTY & ~n35664;
  assign n35666 = ~n27992 & ~n35665;
  assign n35667 = controllable_BtoS_ACK0 & ~n35666;
  assign n35668 = ~controllable_DEQ & ~n28020;
  assign n35669 = ~n11364 & ~n35668;
  assign n35670 = ~i_FULL & ~n35669;
  assign n35671 = ~n28044 & ~n35670;
  assign n35672 = ~i_nEMPTY & ~n35671;
  assign n35673 = ~n28037 & ~n35672;
  assign n35674 = ~controllable_BtoS_ACK0 & ~n35673;
  assign n35675 = ~n35667 & ~n35674;
  assign n35676 = n4465 & ~n35675;
  assign n35677 = ~controllable_DEQ & ~n28067;
  assign n35678 = ~n11364 & ~n35677;
  assign n35679 = ~i_FULL & ~n35678;
  assign n35680 = ~n28091 & ~n35679;
  assign n35681 = ~i_nEMPTY & ~n35680;
  assign n35682 = ~n28084 & ~n35681;
  assign n35683 = ~controllable_BtoS_ACK0 & ~n35682;
  assign n35684 = ~n33468 & ~n35683;
  assign n35685 = ~n4465 & ~n35684;
  assign n35686 = ~n35676 & ~n35685;
  assign n35687 = ~i_StoB_REQ10 & ~n35686;
  assign n35688 = ~n35660 & ~n35687;
  assign n35689 = controllable_BtoS_ACK10 & ~n35688;
  assign n35690 = ~n28281 & ~n35687;
  assign n35691 = ~controllable_BtoS_ACK10 & ~n35690;
  assign n35692 = ~n35689 & ~n35691;
  assign n35693 = n4464 & ~n35692;
  assign n35694 = ~controllable_DEQ & ~n28291;
  assign n35695 = ~n5296 & ~n35694;
  assign n35696 = ~i_FULL & ~n35695;
  assign n35697 = ~n28313 & ~n35696;
  assign n35698 = ~i_nEMPTY & ~n35697;
  assign n35699 = ~n28307 & ~n35698;
  assign n35700 = controllable_BtoS_ACK0 & ~n35699;
  assign n35701 = ~controllable_DEQ & ~n28330;
  assign n35702 = ~n27912 & ~n35701;
  assign n35703 = ~i_FULL & ~n35702;
  assign n35704 = ~n28352 & ~n35703;
  assign n35705 = ~i_nEMPTY & ~n35704;
  assign n35706 = ~n28346 & ~n35705;
  assign n35707 = ~controllable_BtoS_ACK0 & ~n35706;
  assign n35708 = ~n35700 & ~n35707;
  assign n35709 = n4465 & ~n35708;
  assign n35710 = ~n33206 & ~n35707;
  assign n35711 = ~n4465 & ~n35710;
  assign n35712 = ~n35709 & ~n35711;
  assign n35713 = i_StoB_REQ10 & ~n35712;
  assign n35714 = ~controllable_DEQ & ~n28376;
  assign n35715 = ~n11282 & ~n35714;
  assign n35716 = ~i_FULL & ~n35715;
  assign n35717 = ~n28400 & ~n35716;
  assign n35718 = ~i_nEMPTY & ~n35717;
  assign n35719 = ~n28393 & ~n35718;
  assign n35720 = controllable_BtoS_ACK0 & ~n35719;
  assign n35721 = ~controllable_DEQ & ~n28419;
  assign n35722 = ~n11364 & ~n35721;
  assign n35723 = ~i_FULL & ~n35722;
  assign n35724 = ~n28443 & ~n35723;
  assign n35725 = ~i_nEMPTY & ~n35724;
  assign n35726 = ~n28436 & ~n35725;
  assign n35727 = ~controllable_BtoS_ACK0 & ~n35726;
  assign n35728 = ~n35720 & ~n35727;
  assign n35729 = n4465 & ~n35728;
  assign n35730 = ~n33468 & ~n35727;
  assign n35731 = ~n4465 & ~n35730;
  assign n35732 = ~n35729 & ~n35731;
  assign n35733 = ~i_StoB_REQ10 & ~n35732;
  assign n35734 = ~n35713 & ~n35733;
  assign n35735 = controllable_BtoS_ACK10 & ~n35734;
  assign n35736 = ~n28527 & ~n35733;
  assign n35737 = ~controllable_BtoS_ACK10 & ~n35736;
  assign n35738 = ~n35735 & ~n35737;
  assign n35739 = ~n4464 & ~n35738;
  assign n35740 = ~n35693 & ~n35739;
  assign n35741 = n4463 & ~n35740;
  assign n35742 = ~controllable_DEQ & ~n27883;
  assign n35743 = ~n27912 & ~n35742;
  assign n35744 = ~i_FULL & ~n35743;
  assign n35745 = ~n28547 & ~n35744;
  assign n35746 = ~i_nEMPTY & ~n35745;
  assign n35747 = ~n28540 & ~n35746;
  assign n35748 = ~controllable_BtoS_ACK0 & ~n35747;
  assign n35749 = ~n33206 & ~n35748;
  assign n35750 = i_StoB_REQ10 & ~n35749;
  assign n35751 = ~n33477 & ~n35750;
  assign n35752 = controllable_BtoS_ACK10 & ~n35751;
  assign n35753 = ~n28579 & ~n33477;
  assign n35754 = ~controllable_BtoS_ACK10 & ~n35753;
  assign n35755 = ~n35752 & ~n35754;
  assign n35756 = ~n4463 & ~n35755;
  assign n35757 = ~n35741 & ~n35756;
  assign n35758 = n4462 & ~n35757;
  assign n35759 = ~controllable_DEQ & ~n28634;
  assign n35760 = ~n11282 & ~n35759;
  assign n35761 = ~i_FULL & ~n35760;
  assign n35762 = ~n28649 & ~n35761;
  assign n35763 = ~i_nEMPTY & ~n35762;
  assign n35764 = ~n28645 & ~n35763;
  assign n35765 = controllable_BtoS_ACK0 & ~n35764;
  assign n35766 = ~n35683 & ~n35765;
  assign n35767 = n4465 & ~n35766;
  assign n35768 = ~n35685 & ~n35767;
  assign n35769 = ~i_StoB_REQ10 & ~n35768;
  assign n35770 = ~n28627 & ~n35769;
  assign n35771 = ~controllable_BtoS_ACK10 & ~n35770;
  assign n35772 = ~n35752 & ~n35771;
  assign n35773 = n4464 & ~n35772;
  assign n35774 = ~n35737 & ~n35752;
  assign n35775 = ~n4464 & ~n35774;
  assign n35776 = ~n35773 & ~n35775;
  assign n35777 = n4463 & ~n35776;
  assign n35778 = ~n35756 & ~n35777;
  assign n35779 = ~n4462 & ~n35778;
  assign n35780 = ~n35758 & ~n35779;
  assign n35781 = ~n4459 & ~n35780;
  assign n35782 = ~controllable_DEQ & ~n28684;
  assign n35783 = ~n14798 & ~n35782;
  assign n35784 = ~i_FULL & ~n35783;
  assign n35785 = ~n28717 & ~n35784;
  assign n35786 = ~i_nEMPTY & ~n35785;
  assign n35787 = ~n28707 & ~n35786;
  assign n35788 = controllable_BtoS_ACK0 & ~n35787;
  assign n35789 = ~controllable_DEQ & ~n28736;
  assign n35790 = ~n28787 & ~n35789;
  assign n35791 = ~i_FULL & ~n35790;
  assign n35792 = ~n28783 & ~n35791;
  assign n35793 = ~i_nEMPTY & ~n35792;
  assign n35794 = ~n28769 & ~n35793;
  assign n35795 = ~controllable_BtoS_ACK0 & ~n35794;
  assign n35796 = ~n35788 & ~n35795;
  assign n35797 = n4465 & ~n35796;
  assign n35798 = ~controllable_DEQ & ~n28806;
  assign n35799 = ~n28787 & ~n35798;
  assign n35800 = ~i_FULL & ~n35799;
  assign n35801 = ~n28839 & ~n35800;
  assign n35802 = ~i_nEMPTY & ~n35801;
  assign n35803 = ~n28829 & ~n35802;
  assign n35804 = ~controllable_BtoS_ACK0 & ~n35803;
  assign n35805 = ~n33856 & ~n35804;
  assign n35806 = ~n4465 & ~n35805;
  assign n35807 = ~n35797 & ~n35806;
  assign n35808 = i_StoB_REQ10 & ~n35807;
  assign n35809 = ~controllable_DEQ & ~n28860;
  assign n35810 = ~n17673 & ~n35809;
  assign n35811 = ~i_FULL & ~n35810;
  assign n35812 = ~n28893 & ~n35811;
  assign n35813 = ~i_nEMPTY & ~n35812;
  assign n35814 = ~n28883 & ~n35813;
  assign n35815 = controllable_BtoS_ACK0 & ~n35814;
  assign n35816 = ~controllable_DEQ & ~n28912;
  assign n35817 = ~n17774 & ~n35816;
  assign n35818 = ~i_FULL & ~n35817;
  assign n35819 = ~n28945 & ~n35818;
  assign n35820 = ~i_nEMPTY & ~n35819;
  assign n35821 = ~n28935 & ~n35820;
  assign n35822 = ~controllable_BtoS_ACK0 & ~n35821;
  assign n35823 = ~n35815 & ~n35822;
  assign n35824 = n4465 & ~n35823;
  assign n35825 = ~controllable_DEQ & ~n28966;
  assign n35826 = ~n17774 & ~n35825;
  assign n35827 = ~i_FULL & ~n35826;
  assign n35828 = ~n28999 & ~n35827;
  assign n35829 = ~i_nEMPTY & ~n35828;
  assign n35830 = ~n28989 & ~n35829;
  assign n35831 = ~controllable_BtoS_ACK0 & ~n35830;
  assign n35832 = ~n34118 & ~n35831;
  assign n35833 = ~n4465 & ~n35832;
  assign n35834 = ~n35824 & ~n35833;
  assign n35835 = ~i_StoB_REQ10 & ~n35834;
  assign n35836 = ~n35808 & ~n35835;
  assign n35837 = controllable_BtoS_ACK10 & ~n35836;
  assign n35838 = ~n29149 & ~n35835;
  assign n35839 = ~controllable_BtoS_ACK10 & ~n35838;
  assign n35840 = ~n35837 & ~n35839;
  assign n35841 = n4464 & ~n35840;
  assign n35842 = ~controllable_DEQ & ~n29160;
  assign n35843 = ~n14798 & ~n35842;
  assign n35844 = ~i_FULL & ~n35843;
  assign n35845 = ~n29193 & ~n35844;
  assign n35846 = ~i_nEMPTY & ~n35845;
  assign n35847 = ~n29183 & ~n35846;
  assign n35848 = controllable_BtoS_ACK0 & ~n35847;
  assign n35849 = ~controllable_DEQ & ~n29210;
  assign n35850 = ~n28787 & ~n35849;
  assign n35851 = ~i_FULL & ~n35850;
  assign n35852 = ~n29243 & ~n35851;
  assign n35853 = ~i_nEMPTY & ~n35852;
  assign n35854 = ~n29233 & ~n35853;
  assign n35855 = ~controllable_BtoS_ACK0 & ~n35854;
  assign n35856 = ~n35848 & ~n35855;
  assign n35857 = n4465 & ~n35856;
  assign n35858 = ~n33856 & ~n35855;
  assign n35859 = ~n4465 & ~n35858;
  assign n35860 = ~n35857 & ~n35859;
  assign n35861 = i_StoB_REQ10 & ~n35860;
  assign n35862 = ~controllable_DEQ & ~n29266;
  assign n35863 = ~n17673 & ~n35862;
  assign n35864 = ~i_FULL & ~n35863;
  assign n35865 = ~n29299 & ~n35864;
  assign n35866 = ~i_nEMPTY & ~n35865;
  assign n35867 = ~n29289 & ~n35866;
  assign n35868 = controllable_BtoS_ACK0 & ~n35867;
  assign n35869 = ~controllable_DEQ & ~n29316;
  assign n35870 = ~n17774 & ~n35869;
  assign n35871 = ~i_FULL & ~n35870;
  assign n35872 = ~n29349 & ~n35871;
  assign n35873 = ~i_nEMPTY & ~n35872;
  assign n35874 = ~n29339 & ~n35873;
  assign n35875 = ~controllable_BtoS_ACK0 & ~n35874;
  assign n35876 = ~n35868 & ~n35875;
  assign n35877 = n4465 & ~n35876;
  assign n35878 = ~n34118 & ~n35875;
  assign n35879 = ~n4465 & ~n35878;
  assign n35880 = ~n35877 & ~n35879;
  assign n35881 = ~i_StoB_REQ10 & ~n35880;
  assign n35882 = ~n35861 & ~n35881;
  assign n35883 = controllable_BtoS_ACK10 & ~n35882;
  assign n35884 = ~n29427 & ~n35881;
  assign n35885 = ~controllable_BtoS_ACK10 & ~n35884;
  assign n35886 = ~n35883 & ~n35885;
  assign n35887 = ~n4464 & ~n35886;
  assign n35888 = ~n35841 & ~n35887;
  assign n35889 = n4462 & ~n35888;
  assign n35890 = ~controllable_DEQ & ~n28756;
  assign n35891 = ~n28787 & ~n35890;
  assign n35892 = ~i_FULL & ~n35891;
  assign n35893 = ~n29453 & ~n35892;
  assign n35894 = ~i_nEMPTY & ~n35893;
  assign n35895 = ~n29443 & ~n35894;
  assign n35896 = ~controllable_BtoS_ACK0 & ~n35895;
  assign n35897 = ~n33856 & ~n35896;
  assign n35898 = i_StoB_REQ10 & ~n35897;
  assign n35899 = ~n34127 & ~n35898;
  assign n35900 = controllable_BtoS_ACK10 & ~n35899;
  assign n35901 = ~controllable_DEQ & ~n29505;
  assign n35902 = ~n17673 & ~n35901;
  assign n35903 = ~i_FULL & ~n35902;
  assign n35904 = ~n29538 & ~n35903;
  assign n35905 = ~i_nEMPTY & ~n35904;
  assign n35906 = ~n29528 & ~n35905;
  assign n35907 = controllable_BtoS_ACK0 & ~n35906;
  assign n35908 = ~n35831 & ~n35907;
  assign n35909 = n4465 & ~n35908;
  assign n35910 = ~n35833 & ~n35909;
  assign n35911 = ~i_StoB_REQ10 & ~n35910;
  assign n35912 = ~n29498 & ~n35911;
  assign n35913 = ~controllable_BtoS_ACK10 & ~n35912;
  assign n35914 = ~n35900 & ~n35913;
  assign n35915 = n4464 & ~n35914;
  assign n35916 = ~n35885 & ~n35900;
  assign n35917 = ~n4464 & ~n35916;
  assign n35918 = ~n35915 & ~n35917;
  assign n35919 = ~n4462 & ~n35918;
  assign n35920 = ~n35889 & ~n35919;
  assign n35921 = n4461 & ~n35920;
  assign n35922 = ~n29581 & ~n34127;
  assign n35923 = ~controllable_BtoS_ACK10 & ~n35922;
  assign n35924 = ~n35900 & ~n35923;
  assign n35925 = ~n4461 & ~n35924;
  assign n35926 = ~n35921 & ~n35925;
  assign n35927 = n4459 & ~n35926;
  assign n35928 = ~n35781 & ~n35927;
  assign n35929 = n4455 & ~n35928;
  assign n35930 = ~controllable_DEQ & ~n29592;
  assign n35931 = ~n21003 & ~n35930;
  assign n35932 = ~i_FULL & ~n35931;
  assign n35933 = ~n29613 & ~n35932;
  assign n35934 = ~i_nEMPTY & ~n35933;
  assign n35935 = ~n29607 & ~n35934;
  assign n35936 = controllable_BtoS_ACK0 & ~n35935;
  assign n35937 = ~controllable_DEQ & ~n29628;
  assign n35938 = ~n29663 & ~n35937;
  assign n35939 = ~i_FULL & ~n35938;
  assign n35940 = ~n29659 & ~n35939;
  assign n35941 = ~i_nEMPTY & ~n35940;
  assign n35942 = ~n29649 & ~n35941;
  assign n35943 = ~controllable_BtoS_ACK0 & ~n35942;
  assign n35944 = ~n35936 & ~n35943;
  assign n35945 = n4465 & ~n35944;
  assign n35946 = ~controllable_DEQ & ~n29678;
  assign n35947 = ~n29663 & ~n35946;
  assign n35948 = ~i_FULL & ~n35947;
  assign n35949 = ~n29699 & ~n35948;
  assign n35950 = ~i_nEMPTY & ~n35949;
  assign n35951 = ~n29693 & ~n35950;
  assign n35952 = ~controllable_BtoS_ACK0 & ~n35951;
  assign n35953 = ~n34504 & ~n35952;
  assign n35954 = ~n4465 & ~n35953;
  assign n35955 = ~n35945 & ~n35954;
  assign n35956 = i_StoB_REQ10 & ~n35955;
  assign n35957 = ~controllable_DEQ & ~n29716;
  assign n35958 = ~n23117 & ~n35957;
  assign n35959 = ~i_FULL & ~n35958;
  assign n35960 = ~n29737 & ~n35959;
  assign n35961 = ~i_nEMPTY & ~n35960;
  assign n35962 = ~n29731 & ~n35961;
  assign n35963 = controllable_BtoS_ACK0 & ~n35962;
  assign n35964 = ~controllable_DEQ & ~n29750;
  assign n35965 = ~n23157 & ~n35964;
  assign n35966 = ~i_FULL & ~n35965;
  assign n35967 = ~n29771 & ~n35966;
  assign n35968 = ~i_nEMPTY & ~n35967;
  assign n35969 = ~n29765 & ~n35968;
  assign n35970 = ~controllable_BtoS_ACK0 & ~n35969;
  assign n35971 = ~n35963 & ~n35970;
  assign n35972 = n4465 & ~n35971;
  assign n35973 = ~controllable_DEQ & ~n29786;
  assign n35974 = ~n23157 & ~n35973;
  assign n35975 = ~i_FULL & ~n35974;
  assign n35976 = ~n29807 & ~n35975;
  assign n35977 = ~i_nEMPTY & ~n35976;
  assign n35978 = ~n29801 & ~n35977;
  assign n35979 = ~controllable_BtoS_ACK0 & ~n35978;
  assign n35980 = ~n34766 & ~n35979;
  assign n35981 = ~n4465 & ~n35980;
  assign n35982 = ~n35972 & ~n35981;
  assign n35983 = ~i_StoB_REQ10 & ~n35982;
  assign n35984 = ~n35956 & ~n35983;
  assign n35985 = controllable_BtoS_ACK10 & ~n35984;
  assign n35986 = ~n29997 & ~n35983;
  assign n35987 = ~controllable_BtoS_ACK10 & ~n35986;
  assign n35988 = ~n35985 & ~n35987;
  assign n35989 = n4464 & ~n35988;
  assign n35990 = ~controllable_DEQ & ~n30004;
  assign n35991 = ~n21003 & ~n35990;
  assign n35992 = ~i_FULL & ~n35991;
  assign n35993 = ~n30025 & ~n35992;
  assign n35994 = ~i_nEMPTY & ~n35993;
  assign n35995 = ~n30019 & ~n35994;
  assign n35996 = controllable_BtoS_ACK0 & ~n35995;
  assign n35997 = ~controllable_DEQ & ~n30038;
  assign n35998 = ~n29663 & ~n35997;
  assign n35999 = ~i_FULL & ~n35998;
  assign n36000 = ~n30059 & ~n35999;
  assign n36001 = ~i_nEMPTY & ~n36000;
  assign n36002 = ~n30053 & ~n36001;
  assign n36003 = ~controllable_BtoS_ACK0 & ~n36002;
  assign n36004 = ~n35996 & ~n36003;
  assign n36005 = n4465 & ~n36004;
  assign n36006 = ~n34504 & ~n36003;
  assign n36007 = ~n4465 & ~n36006;
  assign n36008 = ~n36005 & ~n36007;
  assign n36009 = i_StoB_REQ10 & ~n36008;
  assign n36010 = ~controllable_DEQ & ~n30078;
  assign n36011 = ~n23117 & ~n36010;
  assign n36012 = ~i_FULL & ~n36011;
  assign n36013 = ~n30099 & ~n36012;
  assign n36014 = ~i_nEMPTY & ~n36013;
  assign n36015 = ~n30093 & ~n36014;
  assign n36016 = controllable_BtoS_ACK0 & ~n36015;
  assign n36017 = ~controllable_DEQ & ~n30112;
  assign n36018 = ~n23157 & ~n36017;
  assign n36019 = ~i_FULL & ~n36018;
  assign n36020 = ~n30133 & ~n36019;
  assign n36021 = ~i_nEMPTY & ~n36020;
  assign n36022 = ~n30127 & ~n36021;
  assign n36023 = ~controllable_BtoS_ACK0 & ~n36022;
  assign n36024 = ~n36016 & ~n36023;
  assign n36025 = n4465 & ~n36024;
  assign n36026 = ~n34766 & ~n36023;
  assign n36027 = ~n4465 & ~n36026;
  assign n36028 = ~n36025 & ~n36027;
  assign n36029 = ~i_StoB_REQ10 & ~n36028;
  assign n36030 = ~n36009 & ~n36029;
  assign n36031 = controllable_BtoS_ACK10 & ~n36030;
  assign n36032 = ~n30227 & ~n36029;
  assign n36033 = ~controllable_BtoS_ACK10 & ~n36032;
  assign n36034 = ~n36031 & ~n36033;
  assign n36035 = ~n4464 & ~n36034;
  assign n36036 = ~n35989 & ~n36035;
  assign n36037 = n4463 & ~n36036;
  assign n36038 = ~controllable_DEQ & ~n30236;
  assign n36039 = ~n21003 & ~n36038;
  assign n36040 = ~i_FULL & ~n36039;
  assign n36041 = ~n30257 & ~n36040;
  assign n36042 = ~i_nEMPTY & ~n36041;
  assign n36043 = ~n30251 & ~n36042;
  assign n36044 = controllable_BtoS_ACK0 & ~n36043;
  assign n36045 = ~controllable_DEQ & ~n30270;
  assign n36046 = ~n29663 & ~n36045;
  assign n36047 = ~i_FULL & ~n36046;
  assign n36048 = ~n30291 & ~n36047;
  assign n36049 = ~i_nEMPTY & ~n36048;
  assign n36050 = ~n30285 & ~n36049;
  assign n36051 = ~controllable_BtoS_ACK0 & ~n36050;
  assign n36052 = ~n36044 & ~n36051;
  assign n36053 = n4465 & ~n36052;
  assign n36054 = ~controllable_DEQ & ~n30306;
  assign n36055 = ~n29663 & ~n36054;
  assign n36056 = ~i_FULL & ~n36055;
  assign n36057 = ~n30327 & ~n36056;
  assign n36058 = ~i_nEMPTY & ~n36057;
  assign n36059 = ~n30321 & ~n36058;
  assign n36060 = ~controllable_BtoS_ACK0 & ~n36059;
  assign n36061 = ~n34504 & ~n36060;
  assign n36062 = ~n4465 & ~n36061;
  assign n36063 = ~n36053 & ~n36062;
  assign n36064 = i_StoB_REQ10 & ~n36063;
  assign n36065 = ~controllable_DEQ & ~n30344;
  assign n36066 = ~n23117 & ~n36065;
  assign n36067 = ~i_FULL & ~n36066;
  assign n36068 = ~n30365 & ~n36067;
  assign n36069 = ~i_nEMPTY & ~n36068;
  assign n36070 = ~n30359 & ~n36069;
  assign n36071 = controllable_BtoS_ACK0 & ~n36070;
  assign n36072 = ~controllable_DEQ & ~n30378;
  assign n36073 = ~n23157 & ~n36072;
  assign n36074 = ~i_FULL & ~n36073;
  assign n36075 = ~n30399 & ~n36074;
  assign n36076 = ~i_nEMPTY & ~n36075;
  assign n36077 = ~n30393 & ~n36076;
  assign n36078 = ~controllable_BtoS_ACK0 & ~n36077;
  assign n36079 = ~n36071 & ~n36078;
  assign n36080 = n4465 & ~n36079;
  assign n36081 = ~controllable_DEQ & ~n30414;
  assign n36082 = ~n23157 & ~n36081;
  assign n36083 = ~i_FULL & ~n36082;
  assign n36084 = ~n30435 & ~n36083;
  assign n36085 = ~i_nEMPTY & ~n36084;
  assign n36086 = ~n30429 & ~n36085;
  assign n36087 = ~controllable_BtoS_ACK0 & ~n36086;
  assign n36088 = ~n34766 & ~n36087;
  assign n36089 = ~n4465 & ~n36088;
  assign n36090 = ~n36080 & ~n36089;
  assign n36091 = ~i_StoB_REQ10 & ~n36090;
  assign n36092 = ~n36064 & ~n36091;
  assign n36093 = controllable_BtoS_ACK10 & ~n36092;
  assign n36094 = ~n30550 & ~n36091;
  assign n36095 = ~controllable_BtoS_ACK10 & ~n36094;
  assign n36096 = ~n36093 & ~n36095;
  assign n36097 = n4464 & ~n36096;
  assign n36098 = ~controllable_DEQ & ~n30557;
  assign n36099 = ~n21003 & ~n36098;
  assign n36100 = ~i_FULL & ~n36099;
  assign n36101 = ~n30578 & ~n36100;
  assign n36102 = ~i_nEMPTY & ~n36101;
  assign n36103 = ~n30572 & ~n36102;
  assign n36104 = controllable_BtoS_ACK0 & ~n36103;
  assign n36105 = ~controllable_DEQ & ~n30591;
  assign n36106 = ~n29663 & ~n36105;
  assign n36107 = ~i_FULL & ~n36106;
  assign n36108 = ~n30612 & ~n36107;
  assign n36109 = ~i_nEMPTY & ~n36108;
  assign n36110 = ~n30606 & ~n36109;
  assign n36111 = ~controllable_BtoS_ACK0 & ~n36110;
  assign n36112 = ~n36104 & ~n36111;
  assign n36113 = n4465 & ~n36112;
  assign n36114 = ~n34504 & ~n36111;
  assign n36115 = ~n4465 & ~n36114;
  assign n36116 = ~n36113 & ~n36115;
  assign n36117 = i_StoB_REQ10 & ~n36116;
  assign n36118 = ~controllable_DEQ & ~n30631;
  assign n36119 = ~n23117 & ~n36118;
  assign n36120 = ~i_FULL & ~n36119;
  assign n36121 = ~n30652 & ~n36120;
  assign n36122 = ~i_nEMPTY & ~n36121;
  assign n36123 = ~n30646 & ~n36122;
  assign n36124 = controllable_BtoS_ACK0 & ~n36123;
  assign n36125 = ~controllable_DEQ & ~n30665;
  assign n36126 = ~n23157 & ~n36125;
  assign n36127 = ~i_FULL & ~n36126;
  assign n36128 = ~n30686 & ~n36127;
  assign n36129 = ~i_nEMPTY & ~n36128;
  assign n36130 = ~n30680 & ~n36129;
  assign n36131 = ~controllable_BtoS_ACK0 & ~n36130;
  assign n36132 = ~n36124 & ~n36131;
  assign n36133 = n4465 & ~n36132;
  assign n36134 = ~n34766 & ~n36131;
  assign n36135 = ~n4465 & ~n36134;
  assign n36136 = ~n36133 & ~n36135;
  assign n36137 = ~i_StoB_REQ10 & ~n36136;
  assign n36138 = ~n36117 & ~n36137;
  assign n36139 = controllable_BtoS_ACK10 & ~n36138;
  assign n36140 = ~n30772 & ~n36137;
  assign n36141 = ~controllable_BtoS_ACK10 & ~n36140;
  assign n36142 = ~n36139 & ~n36141;
  assign n36143 = ~n4464 & ~n36142;
  assign n36144 = ~n36097 & ~n36143;
  assign n36145 = ~n4463 & ~n36144;
  assign n36146 = ~n36037 & ~n36145;
  assign n36147 = n4462 & ~n36146;
  assign n36148 = ~controllable_DEQ & ~n29640;
  assign n36149 = ~n29663 & ~n36148;
  assign n36150 = ~i_FULL & ~n36149;
  assign n36151 = ~n30792 & ~n36150;
  assign n36152 = ~i_nEMPTY & ~n36151;
  assign n36153 = ~n30786 & ~n36152;
  assign n36154 = ~controllable_BtoS_ACK0 & ~n36153;
  assign n36155 = ~n34504 & ~n36154;
  assign n36156 = i_StoB_REQ10 & ~n36155;
  assign n36157 = ~n34775 & ~n36156;
  assign n36158 = controllable_BtoS_ACK10 & ~n36157;
  assign n36159 = ~controllable_DEQ & ~n30848;
  assign n36160 = ~n23117 & ~n36159;
  assign n36161 = ~i_FULL & ~n36160;
  assign n36162 = ~n30869 & ~n36161;
  assign n36163 = ~i_nEMPTY & ~n36162;
  assign n36164 = ~n30863 & ~n36163;
  assign n36165 = controllable_BtoS_ACK0 & ~n36164;
  assign n36166 = ~n35979 & ~n36165;
  assign n36167 = n4465 & ~n36166;
  assign n36168 = ~n35981 & ~n36167;
  assign n36169 = ~i_StoB_REQ10 & ~n36168;
  assign n36170 = ~n30845 & ~n36169;
  assign n36171 = ~controllable_BtoS_ACK10 & ~n36170;
  assign n36172 = ~n36158 & ~n36171;
  assign n36173 = n4464 & ~n36172;
  assign n36174 = ~n36033 & ~n36158;
  assign n36175 = ~n4464 & ~n36174;
  assign n36176 = ~n36173 & ~n36175;
  assign n36177 = n4463 & ~n36176;
  assign n36178 = ~controllable_DEQ & ~n30929;
  assign n36179 = ~n23117 & ~n36178;
  assign n36180 = ~i_FULL & ~n36179;
  assign n36181 = ~n30950 & ~n36180;
  assign n36182 = ~i_nEMPTY & ~n36181;
  assign n36183 = ~n30944 & ~n36182;
  assign n36184 = controllable_BtoS_ACK0 & ~n36183;
  assign n36185 = ~n36087 & ~n36184;
  assign n36186 = n4465 & ~n36185;
  assign n36187 = ~n36089 & ~n36186;
  assign n36188 = ~i_StoB_REQ10 & ~n36187;
  assign n36189 = ~n30926 & ~n36188;
  assign n36190 = ~controllable_BtoS_ACK10 & ~n36189;
  assign n36191 = ~n36158 & ~n36190;
  assign n36192 = n4464 & ~n36191;
  assign n36193 = ~n36141 & ~n36158;
  assign n36194 = ~n4464 & ~n36193;
  assign n36195 = ~n36192 & ~n36194;
  assign n36196 = ~n4463 & ~n36195;
  assign n36197 = ~n36177 & ~n36196;
  assign n36198 = ~n4462 & ~n36197;
  assign n36199 = ~n36147 & ~n36198;
  assign n36200 = n4461 & ~n36199;
  assign n36201 = ~controllable_DEQ & ~n30979;
  assign n36202 = ~n21003 & ~n36201;
  assign n36203 = ~i_FULL & ~n36202;
  assign n36204 = ~n31000 & ~n36203;
  assign n36205 = ~i_nEMPTY & ~n36204;
  assign n36206 = ~n30994 & ~n36205;
  assign n36207 = controllable_BtoS_ACK0 & ~n36206;
  assign n36208 = ~controllable_DEQ & ~n31013;
  assign n36209 = ~n29663 & ~n36208;
  assign n36210 = ~i_FULL & ~n36209;
  assign n36211 = ~n31034 & ~n36210;
  assign n36212 = ~i_nEMPTY & ~n36211;
  assign n36213 = ~n31028 & ~n36212;
  assign n36214 = ~controllable_BtoS_ACK0 & ~n36213;
  assign n36215 = ~n36207 & ~n36214;
  assign n36216 = n4465 & ~n36215;
  assign n36217 = ~controllable_DEQ & ~n31049;
  assign n36218 = ~n29663 & ~n36217;
  assign n36219 = ~i_FULL & ~n36218;
  assign n36220 = ~n31070 & ~n36219;
  assign n36221 = ~i_nEMPTY & ~n36220;
  assign n36222 = ~n31064 & ~n36221;
  assign n36223 = ~controllable_BtoS_ACK0 & ~n36222;
  assign n36224 = ~n34504 & ~n36223;
  assign n36225 = ~n4465 & ~n36224;
  assign n36226 = ~n36216 & ~n36225;
  assign n36227 = i_StoB_REQ10 & ~n36226;
  assign n36228 = ~controllable_DEQ & ~n31087;
  assign n36229 = ~n23117 & ~n36228;
  assign n36230 = ~i_FULL & ~n36229;
  assign n36231 = ~n31108 & ~n36230;
  assign n36232 = ~i_nEMPTY & ~n36231;
  assign n36233 = ~n31102 & ~n36232;
  assign n36234 = controllable_BtoS_ACK0 & ~n36233;
  assign n36235 = ~controllable_DEQ & ~n31121;
  assign n36236 = ~n23157 & ~n36235;
  assign n36237 = ~i_FULL & ~n36236;
  assign n36238 = ~n31142 & ~n36237;
  assign n36239 = ~i_nEMPTY & ~n36238;
  assign n36240 = ~n31136 & ~n36239;
  assign n36241 = ~controllable_BtoS_ACK0 & ~n36240;
  assign n36242 = ~n36234 & ~n36241;
  assign n36243 = n4465 & ~n36242;
  assign n36244 = ~controllable_DEQ & ~n31157;
  assign n36245 = ~n23157 & ~n36244;
  assign n36246 = ~i_FULL & ~n36245;
  assign n36247 = ~n31178 & ~n36246;
  assign n36248 = ~i_nEMPTY & ~n36247;
  assign n36249 = ~n31172 & ~n36248;
  assign n36250 = ~controllable_BtoS_ACK0 & ~n36249;
  assign n36251 = ~n34766 & ~n36250;
  assign n36252 = ~n4465 & ~n36251;
  assign n36253 = ~n36243 & ~n36252;
  assign n36254 = ~i_StoB_REQ10 & ~n36253;
  assign n36255 = ~n36227 & ~n36254;
  assign n36256 = controllable_BtoS_ACK10 & ~n36255;
  assign n36257 = ~n31295 & ~n36254;
  assign n36258 = ~controllable_BtoS_ACK10 & ~n36257;
  assign n36259 = ~n36256 & ~n36258;
  assign n36260 = n4464 & ~n36259;
  assign n36261 = ~controllable_DEQ & ~n31302;
  assign n36262 = ~n21003 & ~n36261;
  assign n36263 = ~i_FULL & ~n36262;
  assign n36264 = ~n31323 & ~n36263;
  assign n36265 = ~i_nEMPTY & ~n36264;
  assign n36266 = ~n31317 & ~n36265;
  assign n36267 = controllable_BtoS_ACK0 & ~n36266;
  assign n36268 = ~controllable_DEQ & ~n31336;
  assign n36269 = ~n29663 & ~n36268;
  assign n36270 = ~i_FULL & ~n36269;
  assign n36271 = ~n31357 & ~n36270;
  assign n36272 = ~i_nEMPTY & ~n36271;
  assign n36273 = ~n31351 & ~n36272;
  assign n36274 = ~controllable_BtoS_ACK0 & ~n36273;
  assign n36275 = ~n36267 & ~n36274;
  assign n36276 = n4465 & ~n36275;
  assign n36277 = ~n34504 & ~n36274;
  assign n36278 = ~n4465 & ~n36277;
  assign n36279 = ~n36276 & ~n36278;
  assign n36280 = i_StoB_REQ10 & ~n36279;
  assign n36281 = ~controllable_DEQ & ~n31376;
  assign n36282 = ~n23117 & ~n36281;
  assign n36283 = ~i_FULL & ~n36282;
  assign n36284 = ~n31397 & ~n36283;
  assign n36285 = ~i_nEMPTY & ~n36284;
  assign n36286 = ~n31391 & ~n36285;
  assign n36287 = controllable_BtoS_ACK0 & ~n36286;
  assign n36288 = ~controllable_DEQ & ~n31410;
  assign n36289 = ~n23157 & ~n36288;
  assign n36290 = ~i_FULL & ~n36289;
  assign n36291 = ~n31431 & ~n36290;
  assign n36292 = ~i_nEMPTY & ~n36291;
  assign n36293 = ~n31425 & ~n36292;
  assign n36294 = ~controllable_BtoS_ACK0 & ~n36293;
  assign n36295 = ~n36287 & ~n36294;
  assign n36296 = n4465 & ~n36295;
  assign n36297 = ~n34766 & ~n36294;
  assign n36298 = ~n4465 & ~n36297;
  assign n36299 = ~n36296 & ~n36298;
  assign n36300 = ~i_StoB_REQ10 & ~n36299;
  assign n36301 = ~n36280 & ~n36300;
  assign n36302 = controllable_BtoS_ACK10 & ~n36301;
  assign n36303 = ~n31517 & ~n36300;
  assign n36304 = ~controllable_BtoS_ACK10 & ~n36303;
  assign n36305 = ~n36302 & ~n36304;
  assign n36306 = ~n4464 & ~n36305;
  assign n36307 = ~n36260 & ~n36306;
  assign n36308 = n4463 & ~n36307;
  assign n36309 = ~n31544 & ~n34775;
  assign n36310 = ~controllable_BtoS_ACK10 & ~n36309;
  assign n36311 = ~n36158 & ~n36310;
  assign n36312 = ~n4463 & ~n36311;
  assign n36313 = ~n36308 & ~n36312;
  assign n36314 = n4462 & ~n36313;
  assign n36315 = ~controllable_DEQ & ~n31588;
  assign n36316 = ~n23117 & ~n36315;
  assign n36317 = ~i_FULL & ~n36316;
  assign n36318 = ~n31609 & ~n36317;
  assign n36319 = ~i_nEMPTY & ~n36318;
  assign n36320 = ~n31603 & ~n36319;
  assign n36321 = controllable_BtoS_ACK0 & ~n36320;
  assign n36322 = ~n36250 & ~n36321;
  assign n36323 = n4465 & ~n36322;
  assign n36324 = ~n36252 & ~n36323;
  assign n36325 = ~i_StoB_REQ10 & ~n36324;
  assign n36326 = ~n31585 & ~n36325;
  assign n36327 = ~controllable_BtoS_ACK10 & ~n36326;
  assign n36328 = ~n36158 & ~n36327;
  assign n36329 = n4464 & ~n36328;
  assign n36330 = ~n36158 & ~n36304;
  assign n36331 = ~n4464 & ~n36330;
  assign n36332 = ~n36329 & ~n36331;
  assign n36333 = n4463 & ~n36332;
  assign n36334 = ~n36312 & ~n36333;
  assign n36335 = ~n4462 & ~n36334;
  assign n36336 = ~n36314 & ~n36335;
  assign n36337 = ~n4461 & ~n36336;
  assign n36338 = ~n36200 & ~n36337;
  assign n36339 = ~n4459 & ~n36338;
  assign n36340 = ~controllable_DEQ & ~n31642;
  assign n36341 = ~n21003 & ~n36340;
  assign n36342 = ~i_FULL & ~n36341;
  assign n36343 = ~n31671 & ~n36342;
  assign n36344 = ~i_nEMPTY & ~n36343;
  assign n36345 = ~n31662 & ~n36344;
  assign n36346 = controllable_BtoS_ACK0 & ~n36345;
  assign n36347 = ~controllable_DEQ & ~n31688;
  assign n36348 = ~n29663 & ~n36347;
  assign n36349 = ~i_FULL & ~n36348;
  assign n36350 = ~n31717 & ~n36349;
  assign n36351 = ~i_nEMPTY & ~n36350;
  assign n36352 = ~n31708 & ~n36351;
  assign n36353 = ~controllable_BtoS_ACK0 & ~n36352;
  assign n36354 = ~n36346 & ~n36353;
  assign n36355 = n4465 & ~n36354;
  assign n36356 = ~controllable_DEQ & ~n31736;
  assign n36357 = ~n29663 & ~n36356;
  assign n36358 = ~i_FULL & ~n36357;
  assign n36359 = ~n31763 & ~n36358;
  assign n36360 = ~i_nEMPTY & ~n36359;
  assign n36361 = ~n31755 & ~n36360;
  assign n36362 = ~controllable_BtoS_ACK0 & ~n36361;
  assign n36363 = ~n34504 & ~n36362;
  assign n36364 = ~n4465 & ~n36363;
  assign n36365 = ~n36355 & ~n36364;
  assign n36366 = i_StoB_REQ10 & ~n36365;
  assign n36367 = ~controllable_DEQ & ~n31784;
  assign n36368 = ~n23117 & ~n36367;
  assign n36369 = ~i_FULL & ~n36368;
  assign n36370 = ~n31813 & ~n36369;
  assign n36371 = ~i_nEMPTY & ~n36370;
  assign n36372 = ~n31804 & ~n36371;
  assign n36373 = controllable_BtoS_ACK0 & ~n36372;
  assign n36374 = ~controllable_DEQ & ~n31830;
  assign n36375 = ~n23157 & ~n36374;
  assign n36376 = ~i_FULL & ~n36375;
  assign n36377 = ~n31859 & ~n36376;
  assign n36378 = ~i_nEMPTY & ~n36377;
  assign n36379 = ~n31850 & ~n36378;
  assign n36380 = ~controllable_BtoS_ACK0 & ~n36379;
  assign n36381 = ~n36373 & ~n36380;
  assign n36382 = n4465 & ~n36381;
  assign n36383 = ~controllable_DEQ & ~n31878;
  assign n36384 = ~n23157 & ~n36383;
  assign n36385 = ~i_FULL & ~n36384;
  assign n36386 = ~n31905 & ~n36385;
  assign n36387 = ~i_nEMPTY & ~n36386;
  assign n36388 = ~n31897 & ~n36387;
  assign n36389 = ~controllable_BtoS_ACK0 & ~n36388;
  assign n36390 = ~n34766 & ~n36389;
  assign n36391 = ~n4465 & ~n36390;
  assign n36392 = ~n36382 & ~n36391;
  assign n36393 = ~i_StoB_REQ10 & ~n36392;
  assign n36394 = ~n36366 & ~n36393;
  assign n36395 = controllable_BtoS_ACK10 & ~n36394;
  assign n36396 = ~n32028 & ~n36393;
  assign n36397 = ~controllable_BtoS_ACK10 & ~n36396;
  assign n36398 = ~n36395 & ~n36397;
  assign n36399 = n4464 & ~n36398;
  assign n36400 = ~controllable_DEQ & ~n32037;
  assign n36401 = ~n21003 & ~n36400;
  assign n36402 = ~i_FULL & ~n36401;
  assign n36403 = ~n32064 & ~n36402;
  assign n36404 = ~i_nEMPTY & ~n36403;
  assign n36405 = ~n32056 & ~n36404;
  assign n36406 = controllable_BtoS_ACK0 & ~n36405;
  assign n36407 = ~controllable_DEQ & ~n32081;
  assign n36408 = ~n29663 & ~n36407;
  assign n36409 = ~i_FULL & ~n36408;
  assign n36410 = ~n32108 & ~n36409;
  assign n36411 = ~i_nEMPTY & ~n36410;
  assign n36412 = ~n32100 & ~n36411;
  assign n36413 = ~controllable_BtoS_ACK0 & ~n36412;
  assign n36414 = ~n36406 & ~n36413;
  assign n36415 = n4465 & ~n36414;
  assign n36416 = ~n34504 & ~n36413;
  assign n36417 = ~n4465 & ~n36416;
  assign n36418 = ~n36415 & ~n36417;
  assign n36419 = i_StoB_REQ10 & ~n36418;
  assign n36420 = ~controllable_DEQ & ~n32131;
  assign n36421 = ~n23117 & ~n36420;
  assign n36422 = ~i_FULL & ~n36421;
  assign n36423 = ~n32158 & ~n36422;
  assign n36424 = ~i_nEMPTY & ~n36423;
  assign n36425 = ~n32150 & ~n36424;
  assign n36426 = controllable_BtoS_ACK0 & ~n36425;
  assign n36427 = ~controllable_DEQ & ~n32175;
  assign n36428 = ~n23157 & ~n36427;
  assign n36429 = ~i_FULL & ~n36428;
  assign n36430 = ~n32202 & ~n36429;
  assign n36431 = ~i_nEMPTY & ~n36430;
  assign n36432 = ~n32194 & ~n36431;
  assign n36433 = ~controllable_BtoS_ACK0 & ~n36432;
  assign n36434 = ~n36426 & ~n36433;
  assign n36435 = n4465 & ~n36434;
  assign n36436 = ~n34766 & ~n36433;
  assign n36437 = ~n4465 & ~n36436;
  assign n36438 = ~n36435 & ~n36437;
  assign n36439 = ~i_StoB_REQ10 & ~n36438;
  assign n36440 = ~n36419 & ~n36439;
  assign n36441 = controllable_BtoS_ACK10 & ~n36440;
  assign n36442 = ~n32294 & ~n36439;
  assign n36443 = ~controllable_BtoS_ACK10 & ~n36442;
  assign n36444 = ~n36441 & ~n36443;
  assign n36445 = ~n4464 & ~n36444;
  assign n36446 = ~n36399 & ~n36445;
  assign n36447 = ~n4463 & ~n36446;
  assign n36448 = ~n36037 & ~n36447;
  assign n36449 = n4462 & ~n36448;
  assign n36450 = ~controllable_DEQ & ~n32350;
  assign n36451 = ~n23117 & ~n36450;
  assign n36452 = ~i_FULL & ~n36451;
  assign n36453 = ~n32371 & ~n36452;
  assign n36454 = ~i_nEMPTY & ~n36453;
  assign n36455 = ~n32365 & ~n36454;
  assign n36456 = controllable_BtoS_ACK0 & ~n36455;
  assign n36457 = ~n36389 & ~n36456;
  assign n36458 = n4465 & ~n36457;
  assign n36459 = ~n36391 & ~n36458;
  assign n36460 = ~i_StoB_REQ10 & ~n36459;
  assign n36461 = ~n32345 & ~n36460;
  assign n36462 = ~controllable_BtoS_ACK10 & ~n36461;
  assign n36463 = ~n36158 & ~n36462;
  assign n36464 = n4464 & ~n36463;
  assign n36465 = ~n36158 & ~n36443;
  assign n36466 = ~n4464 & ~n36465;
  assign n36467 = ~n36464 & ~n36466;
  assign n36468 = ~n4463 & ~n36467;
  assign n36469 = ~n36177 & ~n36468;
  assign n36470 = ~n4462 & ~n36469;
  assign n36471 = ~n36449 & ~n36470;
  assign n36472 = n4461 & ~n36471;
  assign n36473 = ~controllable_DEQ & ~n32404;
  assign n36474 = ~n21003 & ~n36473;
  assign n36475 = ~i_FULL & ~n36474;
  assign n36476 = ~n32432 & ~n36475;
  assign n36477 = ~i_nEMPTY & ~n36476;
  assign n36478 = ~n32424 & ~n36477;
  assign n36479 = controllable_BtoS_ACK0 & ~n36478;
  assign n36480 = ~controllable_DEQ & ~n32449;
  assign n36481 = ~n29663 & ~n36480;
  assign n36482 = ~i_FULL & ~n36481;
  assign n36483 = ~n32477 & ~n36482;
  assign n36484 = ~i_nEMPTY & ~n36483;
  assign n36485 = ~n32469 & ~n36484;
  assign n36486 = ~controllable_BtoS_ACK0 & ~n36485;
  assign n36487 = ~n36479 & ~n36486;
  assign n36488 = n4465 & ~n36487;
  assign n36489 = ~controllable_DEQ & ~n32496;
  assign n36490 = ~n29663 & ~n36489;
  assign n36491 = ~i_FULL & ~n36490;
  assign n36492 = ~n32520 & ~n36491;
  assign n36493 = ~i_nEMPTY & ~n36492;
  assign n36494 = ~n32514 & ~n36493;
  assign n36495 = ~controllable_BtoS_ACK0 & ~n36494;
  assign n36496 = ~n34504 & ~n36495;
  assign n36497 = ~n4465 & ~n36496;
  assign n36498 = ~n36488 & ~n36497;
  assign n36499 = i_StoB_REQ10 & ~n36498;
  assign n36500 = ~controllable_DEQ & ~n32541;
  assign n36501 = ~n23117 & ~n36500;
  assign n36502 = ~i_FULL & ~n36501;
  assign n36503 = ~n32571 & ~n36502;
  assign n36504 = ~i_nEMPTY & ~n36503;
  assign n36505 = ~n32562 & ~n36504;
  assign n36506 = controllable_BtoS_ACK0 & ~n36505;
  assign n36507 = ~controllable_DEQ & ~n32588;
  assign n36508 = ~n23157 & ~n36507;
  assign n36509 = ~i_FULL & ~n36508;
  assign n36510 = ~n32618 & ~n36509;
  assign n36511 = ~i_nEMPTY & ~n36510;
  assign n36512 = ~n32609 & ~n36511;
  assign n36513 = ~controllable_BtoS_ACK0 & ~n36512;
  assign n36514 = ~n36506 & ~n36513;
  assign n36515 = n4465 & ~n36514;
  assign n36516 = ~controllable_DEQ & ~n32637;
  assign n36517 = ~n23157 & ~n36516;
  assign n36518 = ~i_FULL & ~n36517;
  assign n36519 = ~n32667 & ~n36518;
  assign n36520 = ~i_nEMPTY & ~n36519;
  assign n36521 = ~n32658 & ~n36520;
  assign n36522 = ~controllable_BtoS_ACK0 & ~n36521;
  assign n36523 = ~n34766 & ~n36522;
  assign n36524 = ~n4465 & ~n36523;
  assign n36525 = ~n36515 & ~n36524;
  assign n36526 = ~i_StoB_REQ10 & ~n36525;
  assign n36527 = ~n36499 & ~n36526;
  assign n36528 = controllable_BtoS_ACK10 & ~n36527;
  assign n36529 = ~n32790 & ~n36526;
  assign n36530 = ~controllable_BtoS_ACK10 & ~n36529;
  assign n36531 = ~n36528 & ~n36530;
  assign n36532 = n4464 & ~n36531;
  assign n36533 = ~controllable_DEQ & ~n32799;
  assign n36534 = ~n21003 & ~n36533;
  assign n36535 = ~i_FULL & ~n36534;
  assign n36536 = ~n32823 & ~n36535;
  assign n36537 = ~i_nEMPTY & ~n36536;
  assign n36538 = ~n32817 & ~n36537;
  assign n36539 = controllable_BtoS_ACK0 & ~n36538;
  assign n36540 = ~controllable_DEQ & ~n32840;
  assign n36541 = ~n29663 & ~n36540;
  assign n36542 = ~i_FULL & ~n36541;
  assign n36543 = ~n32864 & ~n36542;
  assign n36544 = ~i_nEMPTY & ~n36543;
  assign n36545 = ~n32858 & ~n36544;
  assign n36546 = ~controllable_BtoS_ACK0 & ~n36545;
  assign n36547 = ~n36539 & ~n36546;
  assign n36548 = n4465 & ~n36547;
  assign n36549 = ~n34504 & ~n36546;
  assign n36550 = ~n4465 & ~n36549;
  assign n36551 = ~n36548 & ~n36550;
  assign n36552 = i_StoB_REQ10 & ~n36551;
  assign n36553 = ~controllable_DEQ & ~n32887;
  assign n36554 = ~n23117 & ~n36553;
  assign n36555 = ~i_FULL & ~n36554;
  assign n36556 = ~n32917 & ~n36555;
  assign n36557 = ~i_nEMPTY & ~n36556;
  assign n36558 = ~n32908 & ~n36557;
  assign n36559 = controllable_BtoS_ACK0 & ~n36558;
  assign n36560 = ~controllable_DEQ & ~n32934;
  assign n36561 = ~n23157 & ~n36560;
  assign n36562 = ~i_FULL & ~n36561;
  assign n36563 = ~n32964 & ~n36562;
  assign n36564 = ~i_nEMPTY & ~n36563;
  assign n36565 = ~n32955 & ~n36564;
  assign n36566 = ~controllable_BtoS_ACK0 & ~n36565;
  assign n36567 = ~n36559 & ~n36566;
  assign n36568 = n4465 & ~n36567;
  assign n36569 = ~n34766 & ~n36566;
  assign n36570 = ~n4465 & ~n36569;
  assign n36571 = ~n36568 & ~n36570;
  assign n36572 = ~i_StoB_REQ10 & ~n36571;
  assign n36573 = ~n36552 & ~n36572;
  assign n36574 = controllable_BtoS_ACK10 & ~n36573;
  assign n36575 = ~n33056 & ~n36572;
  assign n36576 = ~controllable_BtoS_ACK10 & ~n36575;
  assign n36577 = ~n36574 & ~n36576;
  assign n36578 = ~n4464 & ~n36577;
  assign n36579 = ~n36532 & ~n36578;
  assign n36580 = n4463 & ~n36579;
  assign n36581 = ~n36312 & ~n36580;
  assign n36582 = n4462 & ~n36581;
  assign n36583 = ~controllable_DEQ & ~n33115;
  assign n36584 = ~n23117 & ~n36583;
  assign n36585 = ~i_FULL & ~n36584;
  assign n36586 = ~n33136 & ~n36585;
  assign n36587 = ~i_nEMPTY & ~n36586;
  assign n36588 = ~n33130 & ~n36587;
  assign n36589 = controllable_BtoS_ACK0 & ~n36588;
  assign n36590 = ~n36522 & ~n36589;
  assign n36591 = n4465 & ~n36590;
  assign n36592 = ~n36524 & ~n36591;
  assign n36593 = ~i_StoB_REQ10 & ~n36592;
  assign n36594 = ~n33110 & ~n36593;
  assign n36595 = ~controllable_BtoS_ACK10 & ~n36594;
  assign n36596 = ~n36158 & ~n36595;
  assign n36597 = n4464 & ~n36596;
  assign n36598 = ~n36158 & ~n36576;
  assign n36599 = ~n4464 & ~n36598;
  assign n36600 = ~n36597 & ~n36599;
  assign n36601 = n4463 & ~n36600;
  assign n36602 = ~n36312 & ~n36601;
  assign n36603 = ~n4462 & ~n36602;
  assign n36604 = ~n36582 & ~n36603;
  assign n36605 = ~n4461 & ~n36604;
  assign n36606 = ~n36472 & ~n36605;
  assign n36607 = n4459 & ~n36606;
  assign n36608 = ~n36339 & ~n36607;
  assign n36609 = ~n4455 & ~n36608;
  assign n36610 = ~n35929 & ~n36609;
  assign n36611 = ~n4445 & ~n36610;
  assign n36612 = ~n35633 & ~n36611;
  assign n36613 = n4442 & ~n36612;
  assign n36614 = ~n4459 & ~n35755;
  assign n36615 = n4459 & ~n35924;
  assign n36616 = ~n36614 & ~n36615;
  assign n36617 = n4455 & ~n36616;
  assign n36618 = ~n4455 & ~n36311;
  assign n36619 = ~n36617 & ~n36618;
  assign n36620 = ~n4442 & ~n36619;
  assign n36621 = ~n36613 & ~n36620;
  assign n36622 = ~n4438 & ~n36621;
  assign n36623 = ~n4438 & ~n36622;
  assign n36624 = ~n4386 & ~n36623;
  assign n36625 = ~n33183 & ~n36624;
  assign n36626 = n4384 & n36625;
  assign n36627 = n4384 & ~n36626;
  assign n36628 = n4244 & ~n36627;
  assign n36629 = ~n11224 & ~n11921;
  assign n36630 = controllable_BtoS_ACK10 & ~n36629;
  assign n36631 = ~i_StoB_REQ14 & ~n8455;
  assign n36632 = controllable_BtoS_ACK14 & ~n36631;
  assign n36633 = ~controllable_BtoS_ACK14 & ~n8454;
  assign n36634 = ~n36632 & ~n36633;
  assign n36635 = controllable_ENQ & ~n36634;
  assign n36636 = controllable_ENQ & ~n36635;
  assign n36637 = i_RtoB_ACK1 & ~n36636;
  assign n36638 = ~i_RtoB_ACK1 & ~n11649;
  assign n36639 = ~n36637 & ~n36638;
  assign n36640 = controllable_BtoR_REQ1 & ~n36639;
  assign n36641 = ~n11650 & ~n36640;
  assign n36642 = ~controllable_BtoR_REQ0 & ~n36641;
  assign n36643 = ~controllable_BtoR_REQ0 & ~n36642;
  assign n36644 = i_RtoB_ACK0 & ~n36643;
  assign n36645 = ~controllable_ENQ & ~n36634;
  assign n36646 = ~n11402 & ~n36645;
  assign n36647 = i_RtoB_ACK1 & ~n36646;
  assign n36648 = ~n11666 & ~n36647;
  assign n36649 = controllable_BtoR_REQ1 & ~n36648;
  assign n36650 = ~n11668 & ~n36649;
  assign n36651 = ~controllable_BtoR_REQ0 & ~n36650;
  assign n36652 = ~controllable_BtoR_REQ0 & ~n36651;
  assign n36653 = ~i_RtoB_ACK0 & ~n36652;
  assign n36654 = ~n36644 & ~n36653;
  assign n36655 = controllable_DEQ & ~n36654;
  assign n36656 = i_RtoB_ACK1 & ~n36634;
  assign n36657 = ~n11701 & ~n36656;
  assign n36658 = controllable_BtoR_REQ1 & ~n36657;
  assign n36659 = ~n11679 & ~n36658;
  assign n36660 = ~controllable_BtoR_REQ0 & ~n36659;
  assign n36661 = ~controllable_BtoR_REQ0 & ~n36660;
  assign n36662 = i_RtoB_ACK0 & ~n36661;
  assign n36663 = ~n11690 & ~n36662;
  assign n36664 = ~controllable_DEQ & ~n36663;
  assign n36665 = ~n36655 & ~n36664;
  assign n36666 = i_FULL & ~n36665;
  assign n36667 = ~n11648 & ~n36645;
  assign n36668 = i_RtoB_ACK1 & ~n36667;
  assign n36669 = ~n11701 & ~n36668;
  assign n36670 = controllable_BtoR_REQ1 & ~n36669;
  assign n36671 = ~n11703 & ~n36670;
  assign n36672 = ~controllable_BtoR_REQ0 & ~n36671;
  assign n36673 = ~controllable_BtoR_REQ0 & ~n36672;
  assign n36674 = ~i_RtoB_ACK0 & ~n36673;
  assign n36675 = ~n36644 & ~n36674;
  assign n36676 = controllable_DEQ & ~n36675;
  assign n36677 = ~n11716 & ~n36662;
  assign n36678 = ~controllable_DEQ & ~n36677;
  assign n36679 = ~n36676 & ~n36678;
  assign n36680 = ~i_FULL & ~n36679;
  assign n36681 = ~n36666 & ~n36680;
  assign n36682 = i_nEMPTY & ~n36681;
  assign n36683 = ~controllable_ENQ & ~n36645;
  assign n36684 = i_RtoB_ACK1 & ~n36683;
  assign n36685 = ~n11730 & ~n36684;
  assign n36686 = controllable_BtoR_REQ1 & ~n36685;
  assign n36687 = ~n11732 & ~n36686;
  assign n36688 = ~controllable_BtoR_REQ0 & ~n36687;
  assign n36689 = ~controllable_BtoR_REQ0 & ~n36688;
  assign n36690 = ~i_RtoB_ACK0 & ~n36689;
  assign n36691 = ~i_RtoB_ACK0 & ~n36690;
  assign n36692 = controllable_DEQ & ~n36691;
  assign n36693 = ~n11744 & ~n36644;
  assign n36694 = ~controllable_DEQ & ~n36693;
  assign n36695 = ~n36692 & ~n36694;
  assign n36696 = i_FULL & ~n36695;
  assign n36697 = ~n11750 & ~n36658;
  assign n36698 = ~controllable_BtoR_REQ0 & ~n36697;
  assign n36699 = ~controllable_BtoR_REQ0 & ~n36698;
  assign n36700 = ~i_RtoB_ACK0 & ~n36699;
  assign n36701 = ~i_RtoB_ACK0 & ~n36700;
  assign n36702 = controllable_DEQ & ~n36701;
  assign n36703 = ~controllable_DEQ & ~n36654;
  assign n36704 = ~n36702 & ~n36703;
  assign n36705 = ~i_FULL & ~n36704;
  assign n36706 = ~n36696 & ~n36705;
  assign n36707 = ~i_nEMPTY & ~n36706;
  assign n36708 = ~n36682 & ~n36707;
  assign n36709 = controllable_BtoS_ACK0 & ~n36708;
  assign n36710 = ~i_StoB_REQ14 & ~n8534;
  assign n36711 = controllable_BtoS_ACK14 & ~n36710;
  assign n36712 = ~controllable_BtoS_ACK14 & ~n7187;
  assign n36713 = ~n36711 & ~n36712;
  assign n36714 = controllable_ENQ & ~n36713;
  assign n36715 = controllable_ENQ & ~n36714;
  assign n36716 = i_RtoB_ACK1 & ~n36715;
  assign n36717 = ~i_RtoB_ACK1 & ~n11796;
  assign n36718 = ~n36716 & ~n36717;
  assign n36719 = controllable_BtoR_REQ1 & ~n36718;
  assign n36720 = ~n11797 & ~n36719;
  assign n36721 = ~controllable_BtoR_REQ0 & ~n36720;
  assign n36722 = ~controllable_BtoR_REQ0 & ~n36721;
  assign n36723 = i_RtoB_ACK0 & ~n36722;
  assign n36724 = ~controllable_ENQ & ~n36713;
  assign n36725 = ~n7256 & ~n36724;
  assign n36726 = i_RtoB_ACK1 & ~n36725;
  assign n36727 = ~n11813 & ~n36726;
  assign n36728 = controllable_BtoR_REQ1 & ~n36727;
  assign n36729 = ~n11815 & ~n36728;
  assign n36730 = ~controllable_BtoR_REQ0 & ~n36729;
  assign n36731 = ~controllable_BtoR_REQ0 & ~n36730;
  assign n36732 = ~i_RtoB_ACK0 & ~n36731;
  assign n36733 = ~n36723 & ~n36732;
  assign n36734 = controllable_DEQ & ~n36733;
  assign n36735 = i_RtoB_ACK1 & ~n36713;
  assign n36736 = ~n11848 & ~n36735;
  assign n36737 = controllable_BtoR_REQ1 & ~n36736;
  assign n36738 = ~n11826 & ~n36737;
  assign n36739 = ~controllable_BtoR_REQ0 & ~n36738;
  assign n36740 = ~controllable_BtoR_REQ0 & ~n36739;
  assign n36741 = i_RtoB_ACK0 & ~n36740;
  assign n36742 = ~n11837 & ~n36741;
  assign n36743 = ~controllable_DEQ & ~n36742;
  assign n36744 = ~n36734 & ~n36743;
  assign n36745 = i_FULL & ~n36744;
  assign n36746 = ~n11795 & ~n36724;
  assign n36747 = i_RtoB_ACK1 & ~n36746;
  assign n36748 = ~n11848 & ~n36747;
  assign n36749 = controllable_BtoR_REQ1 & ~n36748;
  assign n36750 = ~n11850 & ~n36749;
  assign n36751 = ~controllable_BtoR_REQ0 & ~n36750;
  assign n36752 = ~controllable_BtoR_REQ0 & ~n36751;
  assign n36753 = ~i_RtoB_ACK0 & ~n36752;
  assign n36754 = ~n36723 & ~n36753;
  assign n36755 = controllable_DEQ & ~n36754;
  assign n36756 = ~n11863 & ~n36741;
  assign n36757 = ~controllable_DEQ & ~n36756;
  assign n36758 = ~n36755 & ~n36757;
  assign n36759 = ~i_FULL & ~n36758;
  assign n36760 = ~n36745 & ~n36759;
  assign n36761 = i_nEMPTY & ~n36760;
  assign n36762 = ~controllable_ENQ & ~n36724;
  assign n36763 = i_RtoB_ACK1 & ~n36762;
  assign n36764 = ~n11877 & ~n36763;
  assign n36765 = controllable_BtoR_REQ1 & ~n36764;
  assign n36766 = ~n11879 & ~n36765;
  assign n36767 = ~controllable_BtoR_REQ0 & ~n36766;
  assign n36768 = ~controllable_BtoR_REQ0 & ~n36767;
  assign n36769 = ~i_RtoB_ACK0 & ~n36768;
  assign n36770 = ~i_RtoB_ACK0 & ~n36769;
  assign n36771 = controllable_DEQ & ~n36770;
  assign n36772 = ~n11891 & ~n36723;
  assign n36773 = ~controllable_DEQ & ~n36772;
  assign n36774 = ~n36771 & ~n36773;
  assign n36775 = i_FULL & ~n36774;
  assign n36776 = ~n11897 & ~n36737;
  assign n36777 = ~controllable_BtoR_REQ0 & ~n36776;
  assign n36778 = ~controllable_BtoR_REQ0 & ~n36777;
  assign n36779 = ~i_RtoB_ACK0 & ~n36778;
  assign n36780 = ~i_RtoB_ACK0 & ~n36779;
  assign n36781 = controllable_DEQ & ~n36780;
  assign n36782 = ~controllable_DEQ & ~n36733;
  assign n36783 = ~n36781 & ~n36782;
  assign n36784 = ~i_FULL & ~n36783;
  assign n36785 = ~n36775 & ~n36784;
  assign n36786 = ~i_nEMPTY & ~n36785;
  assign n36787 = ~n36761 & ~n36786;
  assign n36788 = ~controllable_BtoS_ACK0 & ~n36787;
  assign n36789 = ~n36709 & ~n36788;
  assign n36790 = n4465 & ~n36789;
  assign n36791 = ~n7681 & ~n36790;
  assign n36792 = i_StoB_REQ10 & ~n36791;
  assign n36793 = ~n11921 & ~n36792;
  assign n36794 = ~controllable_BtoS_ACK10 & ~n36793;
  assign n36795 = ~n36630 & ~n36794;
  assign n36796 = n4464 & ~n36795;
  assign n36797 = ~n8752 & ~n36796;
  assign n36798 = n4463 & ~n36797;
  assign n36799 = ~n4477 & ~n9064;
  assign n36800 = n4476 & ~n36799;
  assign n36801 = ~n9067 & ~n36800;
  assign n36802 = ~i_StoB_REQ3 & ~n36801;
  assign n36803 = ~i_StoB_REQ3 & ~n36802;
  assign n36804 = controllable_BtoS_ACK3 & ~n36803;
  assign n36805 = ~controllable_BtoS_ACK3 & ~n36801;
  assign n36806 = ~n36804 & ~n36805;
  assign n36807 = n4475 & ~n36806;
  assign n36808 = ~n9076 & ~n36807;
  assign n36809 = ~i_StoB_REQ4 & ~n36808;
  assign n36810 = ~i_StoB_REQ4 & ~n36809;
  assign n36811 = controllable_BtoS_ACK4 & ~n36810;
  assign n36812 = ~controllable_BtoS_ACK4 & ~n36808;
  assign n36813 = ~n36811 & ~n36812;
  assign n36814 = n4474 & ~n36813;
  assign n36815 = ~n9085 & ~n36814;
  assign n36816 = ~i_StoB_REQ5 & ~n36815;
  assign n36817 = ~i_StoB_REQ5 & ~n36816;
  assign n36818 = controllable_BtoS_ACK5 & ~n36817;
  assign n36819 = ~controllable_BtoS_ACK5 & ~n36815;
  assign n36820 = ~n36818 & ~n36819;
  assign n36821 = n4473 & ~n36820;
  assign n36822 = ~n9094 & ~n36821;
  assign n36823 = ~i_StoB_REQ8 & ~n36822;
  assign n36824 = ~i_StoB_REQ8 & ~n36823;
  assign n36825 = controllable_BtoS_ACK8 & ~n36824;
  assign n36826 = ~controllable_BtoS_ACK8 & ~n36822;
  assign n36827 = ~n36825 & ~n36826;
  assign n36828 = n4472 & ~n36827;
  assign n36829 = ~n9103 & ~n36828;
  assign n36830 = n4471 & ~n36829;
  assign n36831 = ~n4584 & ~n36830;
  assign n36832 = ~i_StoB_REQ6 & ~n36831;
  assign n36833 = ~i_StoB_REQ6 & ~n36832;
  assign n36834 = controllable_BtoS_ACK6 & ~n36833;
  assign n36835 = ~controllable_BtoS_ACK6 & ~n36831;
  assign n36836 = ~n36834 & ~n36835;
  assign n36837 = ~i_StoB_REQ7 & ~n36836;
  assign n36838 = ~i_StoB_REQ7 & ~n36837;
  assign n36839 = controllable_BtoS_ACK7 & ~n36838;
  assign n36840 = ~controllable_BtoS_ACK7 & ~n36836;
  assign n36841 = ~n36839 & ~n36840;
  assign n36842 = n4470 & ~n36841;
  assign n36843 = ~n9120 & ~n36842;
  assign n36844 = n4469 & ~n36843;
  assign n36845 = ~n4627 & ~n36844;
  assign n36846 = ~i_StoB_REQ9 & ~n36845;
  assign n36847 = ~i_StoB_REQ9 & ~n36846;
  assign n36848 = controllable_BtoS_ACK9 & ~n36847;
  assign n36849 = ~controllable_BtoS_ACK9 & ~n36845;
  assign n36850 = ~n36848 & ~n36849;
  assign n36851 = n4468 & ~n36850;
  assign n36852 = ~n4648 & ~n36851;
  assign n36853 = ~i_StoB_REQ11 & ~n36852;
  assign n36854 = ~i_StoB_REQ11 & ~n36853;
  assign n36855 = controllable_BtoS_ACK11 & ~n36854;
  assign n36856 = ~controllable_BtoS_ACK11 & ~n36852;
  assign n36857 = ~n36855 & ~n36856;
  assign n36858 = n4467 & ~n36857;
  assign n36859 = ~n4670 & ~n36858;
  assign n36860 = ~i_StoB_REQ12 & ~n36859;
  assign n36861 = ~i_StoB_REQ12 & ~n36860;
  assign n36862 = controllable_BtoS_ACK12 & ~n36861;
  assign n36863 = ~controllable_BtoS_ACK12 & ~n36859;
  assign n36864 = ~n36862 & ~n36863;
  assign n36865 = ~controllable_BtoS_ACK13 & ~n36864;
  assign n36866 = ~controllable_BtoS_ACK13 & ~n36865;
  assign n36867 = i_StoB_REQ13 & ~n36866;
  assign n36868 = ~i_StoB_REQ13 & ~n36864;
  assign n36869 = ~n36867 & ~n36868;
  assign n36870 = n4466 & ~n36869;
  assign n36871 = ~n9769 & ~n36870;
  assign n36872 = ~i_StoB_REQ0 & ~n36871;
  assign n36873 = ~i_StoB_REQ0 & ~n36872;
  assign n36874 = ~i_StoB_REQ14 & ~n36873;
  assign n36875 = ~i_StoB_REQ14 & ~n36874;
  assign n36876 = controllable_BtoS_ACK14 & ~n36875;
  assign n36877 = ~controllable_BtoS_ACK14 & ~n36873;
  assign n36878 = ~n36876 & ~n36877;
  assign n36879 = ~i_RtoB_ACK1 & ~n36878;
  assign n36880 = ~n12184 & ~n36879;
  assign n36881 = ~controllable_BtoR_REQ1 & ~n36880;
  assign n36882 = ~n11167 & ~n36881;
  assign n36883 = ~controllable_BtoR_REQ0 & ~n36882;
  assign n36884 = ~controllable_BtoR_REQ0 & ~n36883;
  assign n36885 = i_RtoB_ACK0 & ~n36884;
  assign n36886 = i_RtoB_ACK1 & ~n36878;
  assign n36887 = ~n11156 & ~n36886;
  assign n36888 = controllable_BtoR_REQ1 & ~n36887;
  assign n36889 = ~n11168 & ~n36888;
  assign n36890 = ~controllable_BtoR_REQ0 & ~n36889;
  assign n36891 = ~controllable_BtoR_REQ0 & ~n36890;
  assign n36892 = ~i_RtoB_ACK0 & ~n36891;
  assign n36893 = ~n36885 & ~n36892;
  assign n36894 = ~controllable_DEQ & ~n36893;
  assign n36895 = ~n12183 & ~n36894;
  assign n36896 = i_FULL & ~n36895;
  assign n36897 = ~controllable_ENQ & ~n36878;
  assign n36898 = ~n11143 & ~n36897;
  assign n36899 = ~i_RtoB_ACK1 & ~n36898;
  assign n36900 = ~n12184 & ~n36899;
  assign n36901 = ~controllable_BtoR_REQ1 & ~n36900;
  assign n36902 = ~n36888 & ~n36901;
  assign n36903 = ~controllable_BtoR_REQ0 & ~n36902;
  assign n36904 = ~controllable_BtoR_REQ0 & ~n36903;
  assign n36905 = ~i_RtoB_ACK0 & ~n36904;
  assign n36906 = ~n36885 & ~n36905;
  assign n36907 = ~controllable_DEQ & ~n36906;
  assign n36908 = ~n12183 & ~n36907;
  assign n36909 = ~i_FULL & ~n36908;
  assign n36910 = ~n36896 & ~n36909;
  assign n36911 = i_nEMPTY & ~n36910;
  assign n36912 = controllable_ENQ & ~n36878;
  assign n36913 = controllable_ENQ & ~n36912;
  assign n36914 = ~i_RtoB_ACK1 & ~n36913;
  assign n36915 = ~n11150 & ~n36914;
  assign n36916 = ~controllable_BtoR_REQ1 & ~n36915;
  assign n36917 = ~n11138 & ~n36916;
  assign n36918 = ~controllable_BtoR_REQ0 & ~n36917;
  assign n36919 = ~controllable_BtoR_REQ0 & ~n36918;
  assign n36920 = i_RtoB_ACK0 & ~n36919;
  assign n36921 = i_RtoB_ACK1 & ~n36913;
  assign n36922 = ~n12214 & ~n36921;
  assign n36923 = controllable_BtoR_REQ1 & ~n36922;
  assign n36924 = ~n11145 & ~n36923;
  assign n36925 = ~controllable_BtoR_REQ0 & ~n36924;
  assign n36926 = ~controllable_BtoR_REQ0 & ~n36925;
  assign n36927 = ~i_RtoB_ACK0 & ~n36926;
  assign n36928 = ~n36920 & ~n36927;
  assign n36929 = ~controllable_DEQ & ~n36928;
  assign n36930 = ~n12213 & ~n36929;
  assign n36931 = i_FULL & ~n36930;
  assign n36932 = ~n11153 & ~n36921;
  assign n36933 = controllable_BtoR_REQ1 & ~n36932;
  assign n36934 = ~n4477 & ~n5621;
  assign n36935 = n4476 & ~n36934;
  assign n36936 = ~n4476 & ~n4696;
  assign n36937 = ~n36935 & ~n36936;
  assign n36938 = ~i_StoB_REQ3 & ~n36937;
  assign n36939 = ~i_StoB_REQ3 & ~n36938;
  assign n36940 = controllable_BtoS_ACK3 & ~n36939;
  assign n36941 = i_StoB_REQ3 & ~n36801;
  assign n36942 = ~n36938 & ~n36941;
  assign n36943 = ~controllable_BtoS_ACK3 & ~n36942;
  assign n36944 = ~n36940 & ~n36943;
  assign n36945 = n4475 & ~n36944;
  assign n36946 = ~n4475 & ~n4744;
  assign n36947 = ~n36945 & ~n36946;
  assign n36948 = ~i_StoB_REQ4 & ~n36947;
  assign n36949 = ~i_StoB_REQ4 & ~n36948;
  assign n36950 = controllable_BtoS_ACK4 & ~n36949;
  assign n36951 = i_StoB_REQ4 & ~n36808;
  assign n36952 = ~n36948 & ~n36951;
  assign n36953 = ~controllable_BtoS_ACK4 & ~n36952;
  assign n36954 = ~n36950 & ~n36953;
  assign n36955 = n4474 & ~n36954;
  assign n36956 = ~n4474 & ~n4771;
  assign n36957 = ~n36955 & ~n36956;
  assign n36958 = ~i_StoB_REQ5 & ~n36957;
  assign n36959 = ~i_StoB_REQ5 & ~n36958;
  assign n36960 = controllable_BtoS_ACK5 & ~n36959;
  assign n36961 = i_StoB_REQ5 & ~n36815;
  assign n36962 = ~n36958 & ~n36961;
  assign n36963 = ~controllable_BtoS_ACK5 & ~n36962;
  assign n36964 = ~n36960 & ~n36963;
  assign n36965 = n4473 & ~n36964;
  assign n36966 = ~n4473 & ~n4798;
  assign n36967 = ~n36965 & ~n36966;
  assign n36968 = ~i_StoB_REQ8 & ~n36967;
  assign n36969 = ~i_StoB_REQ8 & ~n36968;
  assign n36970 = controllable_BtoS_ACK8 & ~n36969;
  assign n36971 = i_StoB_REQ8 & ~n36822;
  assign n36972 = ~n36968 & ~n36971;
  assign n36973 = ~controllable_BtoS_ACK8 & ~n36972;
  assign n36974 = ~n36970 & ~n36973;
  assign n36975 = n4472 & ~n36974;
  assign n36976 = ~n4472 & ~n4818;
  assign n36977 = ~n36975 & ~n36976;
  assign n36978 = n4471 & ~n36977;
  assign n36979 = ~n4819 & ~n36978;
  assign n36980 = ~i_StoB_REQ6 & ~n36979;
  assign n36981 = ~i_StoB_REQ6 & ~n36980;
  assign n36982 = controllable_BtoS_ACK6 & ~n36981;
  assign n36983 = i_StoB_REQ6 & ~n36831;
  assign n36984 = ~n36980 & ~n36983;
  assign n36985 = ~controllable_BtoS_ACK6 & ~n36984;
  assign n36986 = ~n36982 & ~n36985;
  assign n36987 = ~i_StoB_REQ7 & ~n36986;
  assign n36988 = ~i_StoB_REQ7 & ~n36987;
  assign n36989 = controllable_BtoS_ACK7 & ~n36988;
  assign n36990 = i_StoB_REQ7 & ~n36836;
  assign n36991 = ~n36987 & ~n36990;
  assign n36992 = ~controllable_BtoS_ACK7 & ~n36991;
  assign n36993 = ~n36989 & ~n36992;
  assign n36994 = n4470 & ~n36993;
  assign n36995 = ~n4470 & ~n4875;
  assign n36996 = ~n36994 & ~n36995;
  assign n36997 = n4469 & ~n36996;
  assign n36998 = ~n4876 & ~n36997;
  assign n36999 = ~i_StoB_REQ9 & ~n36998;
  assign n37000 = ~i_StoB_REQ9 & ~n36999;
  assign n37001 = controllable_BtoS_ACK9 & ~n37000;
  assign n37002 = i_StoB_REQ9 & ~n36845;
  assign n37003 = ~n36999 & ~n37002;
  assign n37004 = ~controllable_BtoS_ACK9 & ~n37003;
  assign n37005 = ~n37001 & ~n37004;
  assign n37006 = n4468 & ~n37005;
  assign n37007 = ~n4901 & ~n37006;
  assign n37008 = ~i_StoB_REQ11 & ~n37007;
  assign n37009 = ~i_StoB_REQ11 & ~n37008;
  assign n37010 = controllable_BtoS_ACK11 & ~n37009;
  assign n37011 = i_StoB_REQ11 & ~n36852;
  assign n37012 = ~n37008 & ~n37011;
  assign n37013 = ~controllable_BtoS_ACK11 & ~n37012;
  assign n37014 = ~n37010 & ~n37013;
  assign n37015 = n4467 & ~n37014;
  assign n37016 = ~n4931 & ~n37015;
  assign n37017 = ~i_StoB_REQ12 & ~n37016;
  assign n37018 = ~i_StoB_REQ12 & ~n37017;
  assign n37019 = controllable_BtoS_ACK12 & ~n37018;
  assign n37020 = i_StoB_REQ12 & ~n36859;
  assign n37021 = ~n37017 & ~n37020;
  assign n37022 = ~controllable_BtoS_ACK12 & ~n37021;
  assign n37023 = ~n37019 & ~n37022;
  assign n37024 = ~i_StoB_REQ13 & ~n37023;
  assign n37025 = ~n36867 & ~n37024;
  assign n37026 = n4466 & ~n37025;
  assign n37027 = ~n4466 & ~n5206;
  assign n37028 = ~n37026 & ~n37027;
  assign n37029 = ~i_StoB_REQ0 & ~n37028;
  assign n37030 = ~i_StoB_REQ0 & ~n37029;
  assign n37031 = ~i_StoB_REQ14 & ~n37030;
  assign n37032 = ~i_StoB_REQ14 & ~n37031;
  assign n37033 = controllable_BtoS_ACK14 & ~n37032;
  assign n37034 = i_StoB_REQ14 & ~n36873;
  assign n37035 = ~n37031 & ~n37034;
  assign n37036 = ~controllable_BtoS_ACK14 & ~n37035;
  assign n37037 = ~n37033 & ~n37036;
  assign n37038 = ~controllable_ENQ & ~n37037;
  assign n37039 = ~n11143 & ~n37038;
  assign n37040 = ~i_RtoB_ACK1 & ~n37039;
  assign n37041 = ~n11150 & ~n37040;
  assign n37042 = ~controllable_BtoR_REQ1 & ~n37041;
  assign n37043 = ~n36933 & ~n37042;
  assign n37044 = ~controllable_BtoR_REQ0 & ~n37043;
  assign n37045 = ~controllable_BtoR_REQ0 & ~n37044;
  assign n37046 = ~i_RtoB_ACK0 & ~n37045;
  assign n37047 = ~n36920 & ~n37046;
  assign n37048 = ~controllable_DEQ & ~n37047;
  assign n37049 = ~n12234 & ~n37048;
  assign n37050 = ~i_FULL & ~n37049;
  assign n37051 = ~n36931 & ~n37050;
  assign n37052 = ~i_nEMPTY & ~n37051;
  assign n37053 = ~n36911 & ~n37052;
  assign n37054 = controllable_BtoS_ACK0 & ~n37053;
  assign n37055 = ~i_StoB_REQ14 & ~n36871;
  assign n37056 = ~i_StoB_REQ14 & ~n37055;
  assign n37057 = controllable_BtoS_ACK14 & ~n37056;
  assign n37058 = ~controllable_BtoS_ACK14 & ~n36871;
  assign n37059 = ~n37057 & ~n37058;
  assign n37060 = ~i_RtoB_ACK1 & ~n37059;
  assign n37061 = ~n8983 & ~n37060;
  assign n37062 = ~controllable_BtoR_REQ1 & ~n37061;
  assign n37063 = ~n5360 & ~n37062;
  assign n37064 = ~controllable_BtoR_REQ0 & ~n37063;
  assign n37065 = ~controllable_BtoR_REQ0 & ~n37064;
  assign n37066 = i_RtoB_ACK0 & ~n37065;
  assign n37067 = i_RtoB_ACK1 & ~n37059;
  assign n37068 = ~n5349 & ~n37067;
  assign n37069 = controllable_BtoR_REQ1 & ~n37068;
  assign n37070 = ~n5361 & ~n37069;
  assign n37071 = ~controllable_BtoR_REQ0 & ~n37070;
  assign n37072 = ~controllable_BtoR_REQ0 & ~n37071;
  assign n37073 = ~i_RtoB_ACK0 & ~n37072;
  assign n37074 = ~n37066 & ~n37073;
  assign n37075 = ~controllable_DEQ & ~n37074;
  assign n37076 = ~n12274 & ~n37075;
  assign n37077 = i_FULL & ~n37076;
  assign n37078 = ~controllable_ENQ & ~n37059;
  assign n37079 = ~n5336 & ~n37078;
  assign n37080 = ~i_RtoB_ACK1 & ~n37079;
  assign n37081 = ~n8983 & ~n37080;
  assign n37082 = ~controllable_BtoR_REQ1 & ~n37081;
  assign n37083 = ~n37069 & ~n37082;
  assign n37084 = ~controllable_BtoR_REQ0 & ~n37083;
  assign n37085 = ~controllable_BtoR_REQ0 & ~n37084;
  assign n37086 = ~i_RtoB_ACK0 & ~n37085;
  assign n37087 = ~n37066 & ~n37086;
  assign n37088 = ~controllable_DEQ & ~n37087;
  assign n37089 = ~n12274 & ~n37088;
  assign n37090 = ~i_FULL & ~n37089;
  assign n37091 = ~n37077 & ~n37090;
  assign n37092 = i_nEMPTY & ~n37091;
  assign n37093 = controllable_ENQ & ~n37059;
  assign n37094 = controllable_ENQ & ~n37093;
  assign n37095 = ~i_RtoB_ACK1 & ~n37094;
  assign n37096 = ~n5343 & ~n37095;
  assign n37097 = ~controllable_BtoR_REQ1 & ~n37096;
  assign n37098 = ~n5330 & ~n37097;
  assign n37099 = ~controllable_BtoR_REQ0 & ~n37098;
  assign n37100 = ~controllable_BtoR_REQ0 & ~n37099;
  assign n37101 = i_RtoB_ACK0 & ~n37100;
  assign n37102 = i_RtoB_ACK1 & ~n37094;
  assign n37103 = ~n9026 & ~n37102;
  assign n37104 = controllable_BtoR_REQ1 & ~n37103;
  assign n37105 = ~n5338 & ~n37104;
  assign n37106 = ~controllable_BtoR_REQ0 & ~n37105;
  assign n37107 = ~controllable_BtoR_REQ0 & ~n37106;
  assign n37108 = ~i_RtoB_ACK0 & ~n37107;
  assign n37109 = ~n37101 & ~n37108;
  assign n37110 = ~controllable_DEQ & ~n37109;
  assign n37111 = ~n12299 & ~n37110;
  assign n37112 = i_FULL & ~n37111;
  assign n37113 = ~n5346 & ~n37102;
  assign n37114 = controllable_BtoR_REQ1 & ~n37113;
  assign n37115 = i_StoB_REQ0 & ~n36871;
  assign n37116 = ~n37029 & ~n37115;
  assign n37117 = ~i_StoB_REQ14 & ~n37116;
  assign n37118 = ~i_StoB_REQ14 & ~n37117;
  assign n37119 = controllable_BtoS_ACK14 & ~n37118;
  assign n37120 = i_StoB_REQ14 & ~n36871;
  assign n37121 = ~n37117 & ~n37120;
  assign n37122 = ~controllable_BtoS_ACK14 & ~n37121;
  assign n37123 = ~n37119 & ~n37122;
  assign n37124 = ~controllable_ENQ & ~n37123;
  assign n37125 = ~n5336 & ~n37124;
  assign n37126 = ~i_RtoB_ACK1 & ~n37125;
  assign n37127 = ~n5343 & ~n37126;
  assign n37128 = ~controllable_BtoR_REQ1 & ~n37127;
  assign n37129 = ~n37114 & ~n37128;
  assign n37130 = ~controllable_BtoR_REQ0 & ~n37129;
  assign n37131 = ~controllable_BtoR_REQ0 & ~n37130;
  assign n37132 = ~i_RtoB_ACK0 & ~n37131;
  assign n37133 = ~n37101 & ~n37132;
  assign n37134 = ~controllable_DEQ & ~n37133;
  assign n37135 = ~n12315 & ~n37134;
  assign n37136 = ~i_FULL & ~n37135;
  assign n37137 = ~n37112 & ~n37136;
  assign n37138 = ~i_nEMPTY & ~n37137;
  assign n37139 = ~n37092 & ~n37138;
  assign n37140 = ~controllable_BtoS_ACK0 & ~n37139;
  assign n37141 = ~n37054 & ~n37140;
  assign n37142 = n4465 & ~n37141;
  assign n37143 = ~n8997 & ~n9007;
  assign n37144 = i_FULL & ~n37143;
  assign n37145 = ~n9017 & ~n37144;
  assign n37146 = i_nEMPTY & ~n37145;
  assign n37147 = ~n9056 & ~n37146;
  assign n37148 = ~controllable_BtoS_ACK0 & ~n37147;
  assign n37149 = ~n5307 & ~n37148;
  assign n37150 = ~n4465 & ~n37149;
  assign n37151 = ~n37142 & ~n37150;
  assign n37152 = i_StoB_REQ10 & ~n37151;
  assign n37153 = ~n7054 & ~n11641;
  assign n37154 = controllable_BtoR_REQ1 & ~n37153;
  assign n37155 = i_StoB_REQ12 & ~n9137;
  assign n37156 = i_StoB_REQ11 & ~n9129;
  assign n37157 = i_StoB_REQ9 & ~n9121;
  assign n37158 = i_StoB_REQ6 & ~n9104;
  assign n37159 = ~n6217 & ~n9155;
  assign n37160 = n4476 & ~n37159;
  assign n37161 = ~n9166 & ~n37160;
  assign n37162 = ~i_StoB_REQ3 & ~n37161;
  assign n37163 = ~n9175 & ~n37162;
  assign n37164 = controllable_BtoS_ACK3 & ~n37163;
  assign n37165 = ~n6250 & ~n37162;
  assign n37166 = ~controllable_BtoS_ACK3 & ~n37165;
  assign n37167 = ~n37164 & ~n37166;
  assign n37168 = n4475 & ~n37167;
  assign n37169 = ~n9179 & ~n37168;
  assign n37170 = ~i_StoB_REQ4 & ~n37169;
  assign n37171 = ~n9188 & ~n37170;
  assign n37172 = controllable_BtoS_ACK4 & ~n37171;
  assign n37173 = ~n6283 & ~n37170;
  assign n37174 = ~controllable_BtoS_ACK4 & ~n37173;
  assign n37175 = ~n37172 & ~n37174;
  assign n37176 = n4474 & ~n37175;
  assign n37177 = ~n9192 & ~n37176;
  assign n37178 = ~i_StoB_REQ5 & ~n37177;
  assign n37179 = ~n9201 & ~n37178;
  assign n37180 = controllable_BtoS_ACK5 & ~n37179;
  assign n37181 = ~n6316 & ~n37178;
  assign n37182 = ~controllable_BtoS_ACK5 & ~n37181;
  assign n37183 = ~n37180 & ~n37182;
  assign n37184 = n4473 & ~n37183;
  assign n37185 = ~n9205 & ~n37184;
  assign n37186 = ~i_StoB_REQ8 & ~n37185;
  assign n37187 = ~n9214 & ~n37186;
  assign n37188 = controllable_BtoS_ACK8 & ~n37187;
  assign n37189 = ~n6341 & ~n37186;
  assign n37190 = ~controllable_BtoS_ACK8 & ~n37189;
  assign n37191 = ~n37188 & ~n37190;
  assign n37192 = n4472 & ~n37191;
  assign n37193 = ~n9218 & ~n37192;
  assign n37194 = n4471 & ~n37193;
  assign n37195 = ~n6022 & ~n37194;
  assign n37196 = ~i_StoB_REQ6 & ~n37195;
  assign n37197 = ~n37158 & ~n37196;
  assign n37198 = controllable_BtoS_ACK6 & ~n37197;
  assign n37199 = ~n6377 & ~n37196;
  assign n37200 = ~controllable_BtoS_ACK6 & ~n37199;
  assign n37201 = ~n37198 & ~n37200;
  assign n37202 = ~i_StoB_REQ7 & ~n37201;
  assign n37203 = ~n9235 & ~n37202;
  assign n37204 = controllable_BtoS_ACK7 & ~n37203;
  assign n37205 = ~n6404 & ~n37202;
  assign n37206 = ~controllable_BtoS_ACK7 & ~n37205;
  assign n37207 = ~n37204 & ~n37206;
  assign n37208 = n4470 & ~n37207;
  assign n37209 = ~n9239 & ~n37208;
  assign n37210 = n4469 & ~n37209;
  assign n37211 = ~n6095 & ~n37210;
  assign n37212 = ~i_StoB_REQ9 & ~n37211;
  assign n37213 = ~n37157 & ~n37212;
  assign n37214 = controllable_BtoS_ACK9 & ~n37213;
  assign n37215 = ~n6432 & ~n37212;
  assign n37216 = ~controllable_BtoS_ACK9 & ~n37215;
  assign n37217 = ~n37214 & ~n37216;
  assign n37218 = n4468 & ~n37217;
  assign n37219 = ~n6130 & ~n37218;
  assign n37220 = ~i_StoB_REQ11 & ~n37219;
  assign n37221 = ~n37156 & ~n37220;
  assign n37222 = controllable_BtoS_ACK11 & ~n37221;
  assign n37223 = ~n6462 & ~n37220;
  assign n37224 = ~controllable_BtoS_ACK11 & ~n37223;
  assign n37225 = ~n37222 & ~n37224;
  assign n37226 = n4467 & ~n37225;
  assign n37227 = ~n6168 & ~n37226;
  assign n37228 = ~i_StoB_REQ12 & ~n37227;
  assign n37229 = ~n37155 & ~n37228;
  assign n37230 = controllable_BtoS_ACK12 & ~n37229;
  assign n37231 = ~n6505 & ~n37228;
  assign n37232 = ~controllable_BtoS_ACK12 & ~n37231;
  assign n37233 = ~n37230 & ~n37232;
  assign n37234 = ~i_StoB_REQ13 & ~n37233;
  assign n37235 = ~n9278 & ~n37234;
  assign n37236 = n4466 & ~n37235;
  assign n37237 = ~n9280 & ~n37236;
  assign n37238 = ~i_StoB_REQ0 & ~n37237;
  assign n37239 = ~n9771 & ~n37238;
  assign n37240 = ~i_StoB_REQ14 & ~n37239;
  assign n37241 = ~n10454 & ~n37240;
  assign n37242 = controllable_BtoS_ACK14 & ~n37241;
  assign n37243 = ~n9287 & ~n37240;
  assign n37244 = ~controllable_BtoS_ACK14 & ~n37243;
  assign n37245 = ~n37242 & ~n37244;
  assign n37246 = controllable_ENQ & ~n37245;
  assign n37247 = controllable_ENQ & ~n37246;
  assign n37248 = ~i_RtoB_ACK1 & ~n37247;
  assign n37249 = ~n11663 & ~n37248;
  assign n37250 = ~controllable_BtoR_REQ1 & ~n37249;
  assign n37251 = ~n37154 & ~n37250;
  assign n37252 = ~controllable_BtoR_REQ0 & ~n37251;
  assign n37253 = ~controllable_BtoR_REQ0 & ~n37252;
  assign n37254 = i_RtoB_ACK0 & ~n37253;
  assign n37255 = ~n9789 & ~n11660;
  assign n37256 = controllable_BtoR_REQ1 & ~n37255;
  assign n37257 = ~controllable_ENQ & ~n37245;
  assign n37258 = ~n9302 & ~n37257;
  assign n37259 = ~i_RtoB_ACK1 & ~n37258;
  assign n37260 = ~n11663 & ~n37259;
  assign n37261 = ~controllable_BtoR_REQ1 & ~n37260;
  assign n37262 = ~n37256 & ~n37261;
  assign n37263 = ~controllable_BtoR_REQ0 & ~n37262;
  assign n37264 = ~controllable_BtoR_REQ0 & ~n37263;
  assign n37265 = ~i_RtoB_ACK0 & ~n37264;
  assign n37266 = ~n37254 & ~n37265;
  assign n37267 = controllable_DEQ & ~n37266;
  assign n37268 = controllable_BtoS_ACK13 & ~n36864;
  assign n37269 = ~n4477 & ~n9164;
  assign n37270 = n4476 & ~n37269;
  assign n37271 = ~n4476 & n5863;
  assign n37272 = ~n37270 & ~n37271;
  assign n37273 = ~i_StoB_REQ3 & ~n37272;
  assign n37274 = ~n36941 & ~n37273;
  assign n37275 = controllable_BtoS_ACK3 & ~n37274;
  assign n37276 = ~controllable_BtoS_ACK3 & ~n37272;
  assign n37277 = ~n37275 & ~n37276;
  assign n37278 = n4475 & ~n37277;
  assign n37279 = ~n4475 & ~n5921;
  assign n37280 = ~n37278 & ~n37279;
  assign n37281 = ~i_StoB_REQ4 & ~n37280;
  assign n37282 = ~n36951 & ~n37281;
  assign n37283 = controllable_BtoS_ACK4 & ~n37282;
  assign n37284 = ~controllable_BtoS_ACK4 & ~n37280;
  assign n37285 = ~n37283 & ~n37284;
  assign n37286 = n4474 & ~n37285;
  assign n37287 = ~n4474 & ~n5956;
  assign n37288 = ~n37286 & ~n37287;
  assign n37289 = ~i_StoB_REQ5 & ~n37288;
  assign n37290 = ~n36961 & ~n37289;
  assign n37291 = controllable_BtoS_ACK5 & ~n37290;
  assign n37292 = ~controllable_BtoS_ACK5 & ~n37288;
  assign n37293 = ~n37291 & ~n37292;
  assign n37294 = n4473 & ~n37293;
  assign n37295 = ~n4473 & ~n5991;
  assign n37296 = ~n37294 & ~n37295;
  assign n37297 = ~i_StoB_REQ8 & ~n37296;
  assign n37298 = ~n36971 & ~n37297;
  assign n37299 = controllable_BtoS_ACK8 & ~n37298;
  assign n37300 = ~controllable_BtoS_ACK8 & ~n37296;
  assign n37301 = ~n37299 & ~n37300;
  assign n37302 = n4472 & ~n37301;
  assign n37303 = ~n4472 & ~n6021;
  assign n37304 = ~n37302 & ~n37303;
  assign n37305 = n4471 & ~n37304;
  assign n37306 = ~n6022 & ~n37305;
  assign n37307 = ~i_StoB_REQ6 & ~n37306;
  assign n37308 = ~n36983 & ~n37307;
  assign n37309 = controllable_BtoS_ACK6 & ~n37308;
  assign n37310 = ~controllable_BtoS_ACK6 & ~n37306;
  assign n37311 = ~n37309 & ~n37310;
  assign n37312 = ~i_StoB_REQ7 & ~n37311;
  assign n37313 = ~n36990 & ~n37312;
  assign n37314 = controllable_BtoS_ACK7 & ~n37313;
  assign n37315 = ~controllable_BtoS_ACK7 & ~n37311;
  assign n37316 = ~n37314 & ~n37315;
  assign n37317 = n4470 & ~n37316;
  assign n37318 = ~n4470 & ~n6094;
  assign n37319 = ~n37317 & ~n37318;
  assign n37320 = n4469 & ~n37319;
  assign n37321 = ~n6095 & ~n37320;
  assign n37322 = ~i_StoB_REQ9 & ~n37321;
  assign n37323 = ~n37002 & ~n37322;
  assign n37324 = controllable_BtoS_ACK9 & ~n37323;
  assign n37325 = ~controllable_BtoS_ACK9 & ~n37321;
  assign n37326 = ~n37324 & ~n37325;
  assign n37327 = n4468 & ~n37326;
  assign n37328 = ~n6130 & ~n37327;
  assign n37329 = ~i_StoB_REQ11 & ~n37328;
  assign n37330 = ~n37011 & ~n37329;
  assign n37331 = controllable_BtoS_ACK11 & ~n37330;
  assign n37332 = ~controllable_BtoS_ACK11 & ~n37328;
  assign n37333 = ~n37331 & ~n37332;
  assign n37334 = n4467 & ~n37333;
  assign n37335 = ~n6168 & ~n37334;
  assign n37336 = ~i_StoB_REQ12 & ~n37335;
  assign n37337 = ~n37020 & ~n37336;
  assign n37338 = controllable_BtoS_ACK12 & ~n37337;
  assign n37339 = ~controllable_BtoS_ACK12 & ~n37335;
  assign n37340 = ~n37338 & ~n37339;
  assign n37341 = ~controllable_BtoS_ACK13 & ~n37340;
  assign n37342 = ~n37268 & ~n37341;
  assign n37343 = i_StoB_REQ13 & ~n37342;
  assign n37344 = ~n9138 & ~n36858;
  assign n37345 = i_StoB_REQ12 & ~n37344;
  assign n37346 = ~n9142 & ~n36851;
  assign n37347 = i_StoB_REQ11 & ~n37346;
  assign n37348 = ~n9146 & ~n36844;
  assign n37349 = i_StoB_REQ9 & ~n37348;
  assign n37350 = ~n9150 & ~n36830;
  assign n37351 = i_StoB_REQ6 & ~n37350;
  assign n37352 = ~n4477 & ~n9155;
  assign n37353 = n4476 & ~n37352;
  assign n37354 = ~n9166 & ~n37353;
  assign n37355 = ~i_StoB_REQ3 & ~n37354;
  assign n37356 = ~n36941 & ~n37355;
  assign n37357 = controllable_BtoS_ACK3 & ~n37356;
  assign n37358 = i_StoB_REQ3 & ~n37272;
  assign n37359 = ~n37355 & ~n37358;
  assign n37360 = ~controllable_BtoS_ACK3 & ~n37359;
  assign n37361 = ~n37357 & ~n37360;
  assign n37362 = n4475 & ~n37361;
  assign n37363 = ~n9179 & ~n37362;
  assign n37364 = ~i_StoB_REQ4 & ~n37363;
  assign n37365 = ~n36951 & ~n37364;
  assign n37366 = controllable_BtoS_ACK4 & ~n37365;
  assign n37367 = i_StoB_REQ4 & ~n37280;
  assign n37368 = ~n37364 & ~n37367;
  assign n37369 = ~controllable_BtoS_ACK4 & ~n37368;
  assign n37370 = ~n37366 & ~n37369;
  assign n37371 = n4474 & ~n37370;
  assign n37372 = ~n9192 & ~n37371;
  assign n37373 = ~i_StoB_REQ5 & ~n37372;
  assign n37374 = ~n36961 & ~n37373;
  assign n37375 = controllable_BtoS_ACK5 & ~n37374;
  assign n37376 = i_StoB_REQ5 & ~n37288;
  assign n37377 = ~n37373 & ~n37376;
  assign n37378 = ~controllable_BtoS_ACK5 & ~n37377;
  assign n37379 = ~n37375 & ~n37378;
  assign n37380 = n4473 & ~n37379;
  assign n37381 = ~n9205 & ~n37380;
  assign n37382 = ~i_StoB_REQ8 & ~n37381;
  assign n37383 = ~n36971 & ~n37382;
  assign n37384 = controllable_BtoS_ACK8 & ~n37383;
  assign n37385 = i_StoB_REQ8 & ~n37296;
  assign n37386 = ~n37382 & ~n37385;
  assign n37387 = ~controllable_BtoS_ACK8 & ~n37386;
  assign n37388 = ~n37384 & ~n37387;
  assign n37389 = n4472 & ~n37388;
  assign n37390 = ~n9218 & ~n37389;
  assign n37391 = n4471 & ~n37390;
  assign n37392 = ~n6022 & ~n37391;
  assign n37393 = ~i_StoB_REQ6 & ~n37392;
  assign n37394 = ~n37351 & ~n37393;
  assign n37395 = controllable_BtoS_ACK6 & ~n37394;
  assign n37396 = i_StoB_REQ6 & ~n37306;
  assign n37397 = ~n37393 & ~n37396;
  assign n37398 = ~controllable_BtoS_ACK6 & ~n37397;
  assign n37399 = ~n37395 & ~n37398;
  assign n37400 = ~i_StoB_REQ7 & ~n37399;
  assign n37401 = ~n36990 & ~n37400;
  assign n37402 = controllable_BtoS_ACK7 & ~n37401;
  assign n37403 = i_StoB_REQ7 & ~n37311;
  assign n37404 = ~n37400 & ~n37403;
  assign n37405 = ~controllable_BtoS_ACK7 & ~n37404;
  assign n37406 = ~n37402 & ~n37405;
  assign n37407 = n4470 & ~n37406;
  assign n37408 = ~n9239 & ~n37407;
  assign n37409 = n4469 & ~n37408;
  assign n37410 = ~n6095 & ~n37409;
  assign n37411 = ~i_StoB_REQ9 & ~n37410;
  assign n37412 = ~n37349 & ~n37411;
  assign n37413 = controllable_BtoS_ACK9 & ~n37412;
  assign n37414 = i_StoB_REQ9 & ~n37321;
  assign n37415 = ~n37411 & ~n37414;
  assign n37416 = ~controllable_BtoS_ACK9 & ~n37415;
  assign n37417 = ~n37413 & ~n37416;
  assign n37418 = n4468 & ~n37417;
  assign n37419 = ~n6130 & ~n37418;
  assign n37420 = ~i_StoB_REQ11 & ~n37419;
  assign n37421 = ~n37347 & ~n37420;
  assign n37422 = controllable_BtoS_ACK11 & ~n37421;
  assign n37423 = i_StoB_REQ11 & ~n37328;
  assign n37424 = ~n37420 & ~n37423;
  assign n37425 = ~controllable_BtoS_ACK11 & ~n37424;
  assign n37426 = ~n37422 & ~n37425;
  assign n37427 = n4467 & ~n37426;
  assign n37428 = ~n6168 & ~n37427;
  assign n37429 = ~i_StoB_REQ12 & ~n37428;
  assign n37430 = ~n37345 & ~n37429;
  assign n37431 = controllable_BtoS_ACK12 & ~n37430;
  assign n37432 = i_StoB_REQ12 & ~n37335;
  assign n37433 = ~n37429 & ~n37432;
  assign n37434 = ~controllable_BtoS_ACK12 & ~n37433;
  assign n37435 = ~n37431 & ~n37434;
  assign n37436 = ~i_StoB_REQ13 & ~n37435;
  assign n37437 = ~n37343 & ~n37436;
  assign n37438 = n4466 & ~n37437;
  assign n37439 = ~n9280 & ~n37438;
  assign n37440 = ~i_StoB_REQ0 & ~n37439;
  assign n37441 = ~n37115 & ~n37440;
  assign n37442 = ~i_StoB_REQ14 & ~n37441;
  assign n37443 = ~n37034 & ~n37442;
  assign n37444 = controllable_BtoS_ACK14 & ~n37443;
  assign n37445 = ~i_StoB_REQ13 & ~n37340;
  assign n37446 = ~n37343 & ~n37445;
  assign n37447 = n4466 & ~n37446;
  assign n37448 = ~n4466 & ~n7070;
  assign n37449 = ~n37447 & ~n37448;
  assign n37450 = ~i_StoB_REQ0 & ~n37449;
  assign n37451 = ~n37115 & ~n37450;
  assign n37452 = i_StoB_REQ14 & ~n37451;
  assign n37453 = ~n37442 & ~n37452;
  assign n37454 = ~controllable_BtoS_ACK14 & ~n37453;
  assign n37455 = ~n37444 & ~n37454;
  assign n37456 = ~i_RtoB_ACK1 & ~n37455;
  assign n37457 = ~n11684 & ~n37456;
  assign n37458 = ~controllable_BtoR_REQ1 & ~n37457;
  assign n37459 = ~n11678 & ~n37458;
  assign n37460 = ~controllable_BtoR_REQ0 & ~n37459;
  assign n37461 = ~controllable_BtoR_REQ0 & ~n37460;
  assign n37462 = i_RtoB_ACK0 & ~n37461;
  assign n37463 = ~i_StoB_REQ14 & ~n37451;
  assign n37464 = ~n37034 & ~n37463;
  assign n37465 = controllable_BtoS_ACK14 & ~n37464;
  assign n37466 = ~controllable_BtoS_ACK14 & ~n37451;
  assign n37467 = ~n37465 & ~n37466;
  assign n37468 = i_RtoB_ACK1 & ~n37467;
  assign n37469 = ~n11429 & ~n37468;
  assign n37470 = controllable_BtoR_REQ1 & ~n37469;
  assign n37471 = ~n12573 & ~n37470;
  assign n37472 = ~controllable_BtoR_REQ0 & ~n37471;
  assign n37473 = ~controllable_BtoR_REQ0 & ~n37472;
  assign n37474 = ~i_RtoB_ACK0 & ~n37473;
  assign n37475 = ~n37462 & ~n37474;
  assign n37476 = ~controllable_DEQ & ~n37475;
  assign n37477 = ~n37267 & ~n37476;
  assign n37478 = i_FULL & ~n37477;
  assign n37479 = ~n9789 & ~n11698;
  assign n37480 = controllable_BtoR_REQ1 & ~n37479;
  assign n37481 = ~n37261 & ~n37480;
  assign n37482 = ~controllable_BtoR_REQ0 & ~n37481;
  assign n37483 = ~controllable_BtoR_REQ0 & ~n37482;
  assign n37484 = ~i_RtoB_ACK0 & ~n37483;
  assign n37485 = ~n37254 & ~n37484;
  assign n37486 = controllable_DEQ & ~n37485;
  assign n37487 = ~n11666 & ~n37468;
  assign n37488 = controllable_BtoR_REQ1 & ~n37487;
  assign n37489 = ~controllable_ENQ & ~n37467;
  assign n37490 = ~n12368 & ~n37489;
  assign n37491 = ~i_RtoB_ACK1 & ~n37490;
  assign n37492 = ~n11684 & ~n37491;
  assign n37493 = ~controllable_BtoR_REQ1 & ~n37492;
  assign n37494 = ~n37488 & ~n37493;
  assign n37495 = ~controllable_BtoR_REQ0 & ~n37494;
  assign n37496 = ~controllable_BtoR_REQ0 & ~n37495;
  assign n37497 = ~i_RtoB_ACK0 & ~n37496;
  assign n37498 = ~n37462 & ~n37497;
  assign n37499 = ~controllable_DEQ & ~n37498;
  assign n37500 = ~n37486 & ~n37499;
  assign n37501 = ~i_FULL & ~n37500;
  assign n37502 = ~n37478 & ~n37501;
  assign n37503 = i_nEMPTY & ~n37502;
  assign n37504 = ~n7127 & ~n11726;
  assign n37505 = controllable_BtoR_REQ1 & ~n37504;
  assign n37506 = ~controllable_ENQ & ~n37257;
  assign n37507 = ~i_RtoB_ACK1 & ~n37506;
  assign n37508 = ~i_RtoB_ACK1 & ~n37507;
  assign n37509 = ~controllable_BtoR_REQ1 & ~n37508;
  assign n37510 = ~n37505 & ~n37509;
  assign n37511 = ~controllable_BtoR_REQ0 & ~n37510;
  assign n37512 = ~controllable_BtoR_REQ0 & ~n37511;
  assign n37513 = ~i_RtoB_ACK0 & ~n37512;
  assign n37514 = ~i_RtoB_ACK0 & ~n37513;
  assign n37515 = controllable_DEQ & ~n37514;
  assign n37516 = controllable_ENQ & ~n37455;
  assign n37517 = controllable_ENQ & ~n37516;
  assign n37518 = ~i_RtoB_ACK1 & ~n37517;
  assign n37519 = ~n11663 & ~n37518;
  assign n37520 = ~controllable_BtoR_REQ1 & ~n37519;
  assign n37521 = ~n11643 & ~n37520;
  assign n37522 = ~controllable_BtoR_REQ0 & ~n37521;
  assign n37523 = ~controllable_BtoR_REQ0 & ~n37522;
  assign n37524 = i_RtoB_ACK0 & ~n37523;
  assign n37525 = controllable_ENQ & ~n37467;
  assign n37526 = controllable_ENQ & ~n37525;
  assign n37527 = i_RtoB_ACK1 & ~n37526;
  assign n37528 = ~n11479 & ~n37527;
  assign n37529 = controllable_BtoR_REQ1 & ~n37528;
  assign n37530 = ~n12613 & ~n37529;
  assign n37531 = ~controllable_BtoR_REQ0 & ~n37530;
  assign n37532 = ~controllable_BtoR_REQ0 & ~n37531;
  assign n37533 = ~i_RtoB_ACK0 & ~n37532;
  assign n37534 = ~n37524 & ~n37533;
  assign n37535 = ~controllable_DEQ & ~n37534;
  assign n37536 = ~n37515 & ~n37535;
  assign n37537 = i_FULL & ~n37536;
  assign n37538 = ~n7111 & ~n11676;
  assign n37539 = controllable_BtoR_REQ1 & ~n37538;
  assign n37540 = ~i_RtoB_ACK1 & ~n37245;
  assign n37541 = ~i_RtoB_ACK1 & ~n37540;
  assign n37542 = ~controllable_BtoR_REQ1 & ~n37541;
  assign n37543 = ~n37539 & ~n37542;
  assign n37544 = ~controllable_BtoR_REQ0 & ~n37543;
  assign n37545 = ~controllable_BtoR_REQ0 & ~n37544;
  assign n37546 = ~i_RtoB_ACK0 & ~n37545;
  assign n37547 = ~i_RtoB_ACK0 & ~n37546;
  assign n37548 = controllable_DEQ & ~n37547;
  assign n37549 = ~n11655 & ~n37525;
  assign n37550 = i_RtoB_ACK1 & ~n37549;
  assign n37551 = ~n11660 & ~n37550;
  assign n37552 = controllable_BtoR_REQ1 & ~n37551;
  assign n37553 = i_StoB_REQ14 & ~n37030;
  assign n37554 = i_StoB_REQ0 & ~n37028;
  assign n37555 = controllable_BtoS_ACK13 & ~n37023;
  assign n37556 = ~n37341 & ~n37555;
  assign n37557 = i_StoB_REQ13 & ~n37556;
  assign n37558 = i_StoB_REQ12 & ~n37016;
  assign n37559 = i_StoB_REQ11 & ~n37007;
  assign n37560 = i_StoB_REQ9 & ~n36998;
  assign n37561 = i_StoB_REQ7 & ~n36986;
  assign n37562 = i_StoB_REQ6 & ~n36979;
  assign n37563 = i_StoB_REQ8 & ~n36967;
  assign n37564 = i_StoB_REQ5 & ~n36957;
  assign n37565 = i_StoB_REQ4 & ~n36947;
  assign n37566 = i_StoB_REQ3 & ~n36937;
  assign n37567 = ~n4477 & ~n6216;
  assign n37568 = ~n4477 & ~n37567;
  assign n37569 = n4476 & ~n37568;
  assign n37570 = ~n4476 & ~n6216;
  assign n37571 = ~n37569 & ~n37570;
  assign n37572 = ~i_StoB_REQ3 & ~n37571;
  assign n37573 = ~n37566 & ~n37572;
  assign n37574 = controllable_BtoS_ACK3 & ~n37573;
  assign n37575 = ~n37358 & ~n37572;
  assign n37576 = ~controllable_BtoS_ACK3 & ~n37575;
  assign n37577 = ~n37574 & ~n37576;
  assign n37578 = n4475 & ~n37577;
  assign n37579 = ~n4475 & ~n6253;
  assign n37580 = ~n37578 & ~n37579;
  assign n37581 = ~i_StoB_REQ4 & ~n37580;
  assign n37582 = ~n37565 & ~n37581;
  assign n37583 = controllable_BtoS_ACK4 & ~n37582;
  assign n37584 = ~n37367 & ~n37581;
  assign n37585 = ~controllable_BtoS_ACK4 & ~n37584;
  assign n37586 = ~n37583 & ~n37585;
  assign n37587 = n4474 & ~n37586;
  assign n37588 = ~n4474 & ~n6286;
  assign n37589 = ~n37587 & ~n37588;
  assign n37590 = ~i_StoB_REQ5 & ~n37589;
  assign n37591 = ~n37564 & ~n37590;
  assign n37592 = controllable_BtoS_ACK5 & ~n37591;
  assign n37593 = ~n37376 & ~n37590;
  assign n37594 = ~controllable_BtoS_ACK5 & ~n37593;
  assign n37595 = ~n37592 & ~n37594;
  assign n37596 = n4473 & ~n37595;
  assign n37597 = ~n4473 & ~n6319;
  assign n37598 = ~n37596 & ~n37597;
  assign n37599 = ~i_StoB_REQ8 & ~n37598;
  assign n37600 = ~n37563 & ~n37599;
  assign n37601 = controllable_BtoS_ACK8 & ~n37600;
  assign n37602 = ~n37385 & ~n37599;
  assign n37603 = ~controllable_BtoS_ACK8 & ~n37602;
  assign n37604 = ~n37601 & ~n37603;
  assign n37605 = n4472 & ~n37604;
  assign n37606 = ~n4472 & ~n6344;
  assign n37607 = ~n37605 & ~n37606;
  assign n37608 = n4471 & ~n37607;
  assign n37609 = ~n6345 & ~n37608;
  assign n37610 = ~i_StoB_REQ6 & ~n37609;
  assign n37611 = ~n37562 & ~n37610;
  assign n37612 = controllable_BtoS_ACK6 & ~n37611;
  assign n37613 = ~n37396 & ~n37610;
  assign n37614 = ~controllable_BtoS_ACK6 & ~n37613;
  assign n37615 = ~n37612 & ~n37614;
  assign n37616 = ~i_StoB_REQ7 & ~n37615;
  assign n37617 = ~n37561 & ~n37616;
  assign n37618 = controllable_BtoS_ACK7 & ~n37617;
  assign n37619 = ~n37403 & ~n37616;
  assign n37620 = ~controllable_BtoS_ACK7 & ~n37619;
  assign n37621 = ~n37618 & ~n37620;
  assign n37622 = n4470 & ~n37621;
  assign n37623 = ~n4470 & ~n6407;
  assign n37624 = ~n37622 & ~n37623;
  assign n37625 = n4469 & ~n37624;
  assign n37626 = ~n6408 & ~n37625;
  assign n37627 = ~i_StoB_REQ9 & ~n37626;
  assign n37628 = ~n37560 & ~n37627;
  assign n37629 = controllable_BtoS_ACK9 & ~n37628;
  assign n37630 = ~n37414 & ~n37627;
  assign n37631 = ~controllable_BtoS_ACK9 & ~n37630;
  assign n37632 = ~n37629 & ~n37631;
  assign n37633 = n4468 & ~n37632;
  assign n37634 = ~n6436 & ~n37633;
  assign n37635 = ~i_StoB_REQ11 & ~n37634;
  assign n37636 = ~n37559 & ~n37635;
  assign n37637 = controllable_BtoS_ACK11 & ~n37636;
  assign n37638 = ~n37423 & ~n37635;
  assign n37639 = ~controllable_BtoS_ACK11 & ~n37638;
  assign n37640 = ~n37637 & ~n37639;
  assign n37641 = n4467 & ~n37640;
  assign n37642 = ~n6466 & ~n37641;
  assign n37643 = ~i_StoB_REQ12 & ~n37642;
  assign n37644 = ~n37558 & ~n37643;
  assign n37645 = controllable_BtoS_ACK12 & ~n37644;
  assign n37646 = ~n37432 & ~n37643;
  assign n37647 = ~controllable_BtoS_ACK12 & ~n37646;
  assign n37648 = ~n37645 & ~n37647;
  assign n37649 = ~i_StoB_REQ13 & ~n37648;
  assign n37650 = ~n37557 & ~n37649;
  assign n37651 = n4466 & ~n37650;
  assign n37652 = ~n4466 & ~n7061;
  assign n37653 = ~n37651 & ~n37652;
  assign n37654 = ~i_StoB_REQ0 & ~n37653;
  assign n37655 = ~n37554 & ~n37654;
  assign n37656 = ~i_StoB_REQ14 & ~n37655;
  assign n37657 = ~n37553 & ~n37656;
  assign n37658 = controllable_BtoS_ACK14 & ~n37657;
  assign n37659 = ~n37452 & ~n37656;
  assign n37660 = ~controllable_BtoS_ACK14 & ~n37659;
  assign n37661 = ~n37658 & ~n37660;
  assign n37662 = ~controllable_ENQ & ~n37661;
  assign n37663 = ~n12368 & ~n37662;
  assign n37664 = ~i_RtoB_ACK1 & ~n37663;
  assign n37665 = ~n11663 & ~n37664;
  assign n37666 = ~controllable_BtoR_REQ1 & ~n37665;
  assign n37667 = ~n37552 & ~n37666;
  assign n37668 = ~controllable_BtoR_REQ0 & ~n37667;
  assign n37669 = ~controllable_BtoR_REQ0 & ~n37668;
  assign n37670 = ~i_RtoB_ACK0 & ~n37669;
  assign n37671 = ~n37524 & ~n37670;
  assign n37672 = ~controllable_DEQ & ~n37671;
  assign n37673 = ~n37548 & ~n37672;
  assign n37674 = ~i_FULL & ~n37673;
  assign n37675 = ~n37537 & ~n37674;
  assign n37676 = ~i_nEMPTY & ~n37675;
  assign n37677 = ~n37503 & ~n37676;
  assign n37678 = controllable_BtoS_ACK0 & ~n37677;
  assign n37679 = ~n11299 & ~n11788;
  assign n37680 = controllable_BtoR_REQ1 & ~n37679;
  assign n37681 = ~n8058 & ~n37238;
  assign n37682 = ~i_StoB_REQ14 & ~n37681;
  assign n37683 = ~n10584 & ~n37682;
  assign n37684 = controllable_BtoS_ACK14 & ~n37683;
  assign n37685 = ~n9618 & ~n37682;
  assign n37686 = ~controllable_BtoS_ACK14 & ~n37685;
  assign n37687 = ~n37684 & ~n37686;
  assign n37688 = controllable_ENQ & ~n37687;
  assign n37689 = controllable_ENQ & ~n37688;
  assign n37690 = ~i_RtoB_ACK1 & ~n37689;
  assign n37691 = ~n11810 & ~n37690;
  assign n37692 = ~controllable_BtoR_REQ1 & ~n37691;
  assign n37693 = ~n37680 & ~n37692;
  assign n37694 = ~controllable_BtoR_REQ0 & ~n37693;
  assign n37695 = ~controllable_BtoR_REQ0 & ~n37694;
  assign n37696 = i_RtoB_ACK0 & ~n37695;
  assign n37697 = ~n11311 & ~n11807;
  assign n37698 = controllable_BtoR_REQ1 & ~n37697;
  assign n37699 = ~controllable_ENQ & ~n37687;
  assign n37700 = ~n9635 & ~n37699;
  assign n37701 = ~i_RtoB_ACK1 & ~n37700;
  assign n37702 = ~n11810 & ~n37701;
  assign n37703 = ~controllable_BtoR_REQ1 & ~n37702;
  assign n37704 = ~n37698 & ~n37703;
  assign n37705 = ~controllable_BtoR_REQ0 & ~n37704;
  assign n37706 = ~controllable_BtoR_REQ0 & ~n37705;
  assign n37707 = ~i_RtoB_ACK0 & ~n37706;
  assign n37708 = ~n37696 & ~n37707;
  assign n37709 = controllable_DEQ & ~n37708;
  assign n37710 = i_StoB_REQ0 & ~n37449;
  assign n37711 = ~n37440 & ~n37710;
  assign n37712 = ~i_StoB_REQ14 & ~n37711;
  assign n37713 = ~n37120 & ~n37712;
  assign n37714 = controllable_BtoS_ACK14 & ~n37713;
  assign n37715 = i_StoB_REQ14 & ~n37449;
  assign n37716 = ~n37712 & ~n37715;
  assign n37717 = ~controllable_BtoS_ACK14 & ~n37716;
  assign n37718 = ~n37714 & ~n37717;
  assign n37719 = ~i_RtoB_ACK1 & ~n37718;
  assign n37720 = ~n11831 & ~n37719;
  assign n37721 = ~controllable_BtoR_REQ1 & ~n37720;
  assign n37722 = ~n11825 & ~n37721;
  assign n37723 = ~controllable_BtoR_REQ0 & ~n37722;
  assign n37724 = ~controllable_BtoR_REQ0 & ~n37723;
  assign n37725 = i_RtoB_ACK0 & ~n37724;
  assign n37726 = ~i_StoB_REQ14 & ~n37449;
  assign n37727 = ~n37120 & ~n37726;
  assign n37728 = controllable_BtoS_ACK14 & ~n37727;
  assign n37729 = ~controllable_BtoS_ACK14 & ~n37449;
  assign n37730 = ~n37728 & ~n37729;
  assign n37731 = i_RtoB_ACK1 & ~n37730;
  assign n37732 = ~n7288 & ~n37731;
  assign n37733 = controllable_BtoR_REQ1 & ~n37732;
  assign n37734 = ~n12669 & ~n37733;
  assign n37735 = ~controllable_BtoR_REQ0 & ~n37734;
  assign n37736 = ~controllable_BtoR_REQ0 & ~n37735;
  assign n37737 = ~i_RtoB_ACK0 & ~n37736;
  assign n37738 = ~n37725 & ~n37737;
  assign n37739 = ~controllable_DEQ & ~n37738;
  assign n37740 = ~n37709 & ~n37739;
  assign n37741 = i_FULL & ~n37740;
  assign n37742 = ~n11311 & ~n11845;
  assign n37743 = controllable_BtoR_REQ1 & ~n37742;
  assign n37744 = ~n37703 & ~n37743;
  assign n37745 = ~controllable_BtoR_REQ0 & ~n37744;
  assign n37746 = ~controllable_BtoR_REQ0 & ~n37745;
  assign n37747 = ~i_RtoB_ACK0 & ~n37746;
  assign n37748 = ~n37696 & ~n37747;
  assign n37749 = controllable_DEQ & ~n37748;
  assign n37750 = ~n11813 & ~n37731;
  assign n37751 = controllable_BtoR_REQ1 & ~n37750;
  assign n37752 = ~controllable_ENQ & ~n37730;
  assign n37753 = ~n9893 & ~n37752;
  assign n37754 = ~i_RtoB_ACK1 & ~n37753;
  assign n37755 = ~n11831 & ~n37754;
  assign n37756 = ~controllable_BtoR_REQ1 & ~n37755;
  assign n37757 = ~n37751 & ~n37756;
  assign n37758 = ~controllable_BtoR_REQ0 & ~n37757;
  assign n37759 = ~controllable_BtoR_REQ0 & ~n37758;
  assign n37760 = ~i_RtoB_ACK0 & ~n37759;
  assign n37761 = ~n37725 & ~n37760;
  assign n37762 = ~controllable_DEQ & ~n37761;
  assign n37763 = ~n37749 & ~n37762;
  assign n37764 = ~i_FULL & ~n37763;
  assign n37765 = ~n37741 & ~n37764;
  assign n37766 = i_nEMPTY & ~n37765;
  assign n37767 = ~n11341 & ~n11873;
  assign n37768 = controllable_BtoR_REQ1 & ~n37767;
  assign n37769 = ~controllable_ENQ & ~n37699;
  assign n37770 = ~i_RtoB_ACK1 & ~n37769;
  assign n37771 = ~i_RtoB_ACK1 & ~n37770;
  assign n37772 = ~controllable_BtoR_REQ1 & ~n37771;
  assign n37773 = ~n37768 & ~n37772;
  assign n37774 = ~controllable_BtoR_REQ0 & ~n37773;
  assign n37775 = ~controllable_BtoR_REQ0 & ~n37774;
  assign n37776 = ~i_RtoB_ACK0 & ~n37775;
  assign n37777 = ~i_RtoB_ACK0 & ~n37776;
  assign n37778 = controllable_DEQ & ~n37777;
  assign n37779 = controllable_ENQ & ~n37718;
  assign n37780 = controllable_ENQ & ~n37779;
  assign n37781 = ~i_RtoB_ACK1 & ~n37780;
  assign n37782 = ~n11810 & ~n37781;
  assign n37783 = ~controllable_BtoR_REQ1 & ~n37782;
  assign n37784 = ~n11790 & ~n37783;
  assign n37785 = ~controllable_BtoR_REQ0 & ~n37784;
  assign n37786 = ~controllable_BtoR_REQ0 & ~n37785;
  assign n37787 = i_RtoB_ACK0 & ~n37786;
  assign n37788 = controllable_ENQ & ~n37730;
  assign n37789 = controllable_ENQ & ~n37788;
  assign n37790 = i_RtoB_ACK1 & ~n37789;
  assign n37791 = ~n7345 & ~n37790;
  assign n37792 = controllable_BtoR_REQ1 & ~n37791;
  assign n37793 = ~n12709 & ~n37792;
  assign n37794 = ~controllable_BtoR_REQ0 & ~n37793;
  assign n37795 = ~controllable_BtoR_REQ0 & ~n37794;
  assign n37796 = ~i_RtoB_ACK0 & ~n37795;
  assign n37797 = ~n37787 & ~n37796;
  assign n37798 = ~controllable_DEQ & ~n37797;
  assign n37799 = ~n37778 & ~n37798;
  assign n37800 = i_FULL & ~n37799;
  assign n37801 = ~n11324 & ~n11823;
  assign n37802 = controllable_BtoR_REQ1 & ~n37801;
  assign n37803 = ~i_RtoB_ACK1 & ~n37687;
  assign n37804 = ~i_RtoB_ACK1 & ~n37803;
  assign n37805 = ~controllable_BtoR_REQ1 & ~n37804;
  assign n37806 = ~n37802 & ~n37805;
  assign n37807 = ~controllable_BtoR_REQ0 & ~n37806;
  assign n37808 = ~controllable_BtoR_REQ0 & ~n37807;
  assign n37809 = ~i_RtoB_ACK0 & ~n37808;
  assign n37810 = ~i_RtoB_ACK0 & ~n37809;
  assign n37811 = controllable_DEQ & ~n37810;
  assign n37812 = ~n11802 & ~n37788;
  assign n37813 = i_RtoB_ACK1 & ~n37812;
  assign n37814 = ~n11807 & ~n37813;
  assign n37815 = controllable_BtoR_REQ1 & ~n37814;
  assign n37816 = i_StoB_REQ14 & ~n37116;
  assign n37817 = ~n37654 & ~n37710;
  assign n37818 = ~i_StoB_REQ14 & ~n37817;
  assign n37819 = ~n37816 & ~n37818;
  assign n37820 = controllable_BtoS_ACK14 & ~n37819;
  assign n37821 = ~n37715 & ~n37818;
  assign n37822 = ~controllable_BtoS_ACK14 & ~n37821;
  assign n37823 = ~n37820 & ~n37822;
  assign n37824 = ~controllable_ENQ & ~n37823;
  assign n37825 = ~n9893 & ~n37824;
  assign n37826 = ~i_RtoB_ACK1 & ~n37825;
  assign n37827 = ~n11810 & ~n37826;
  assign n37828 = ~controllable_BtoR_REQ1 & ~n37827;
  assign n37829 = ~n37815 & ~n37828;
  assign n37830 = ~controllable_BtoR_REQ0 & ~n37829;
  assign n37831 = ~controllable_BtoR_REQ0 & ~n37830;
  assign n37832 = ~i_RtoB_ACK0 & ~n37831;
  assign n37833 = ~n37787 & ~n37832;
  assign n37834 = ~controllable_DEQ & ~n37833;
  assign n37835 = ~n37811 & ~n37834;
  assign n37836 = ~i_FULL & ~n37835;
  assign n37837 = ~n37800 & ~n37836;
  assign n37838 = ~i_nEMPTY & ~n37837;
  assign n37839 = ~n37766 & ~n37838;
  assign n37840 = ~controllable_BtoS_ACK0 & ~n37839;
  assign n37841 = ~n37678 & ~n37840;
  assign n37842 = n4465 & ~n37841;
  assign n37843 = ~n7232 & ~n11299;
  assign n37844 = controllable_BtoR_REQ1 & ~n37843;
  assign n37845 = ~n9873 & ~n37844;
  assign n37846 = ~controllable_BtoR_REQ0 & ~n37845;
  assign n37847 = ~controllable_BtoR_REQ0 & ~n37846;
  assign n37848 = i_RtoB_ACK0 & ~n37847;
  assign n37849 = ~n7262 & ~n11311;
  assign n37850 = controllable_BtoR_REQ1 & ~n37849;
  assign n37851 = ~n9927 & ~n37850;
  assign n37852 = ~controllable_BtoR_REQ0 & ~n37851;
  assign n37853 = ~controllable_BtoR_REQ0 & ~n37852;
  assign n37854 = ~i_RtoB_ACK0 & ~n37853;
  assign n37855 = ~n37848 & ~n37854;
  assign n37856 = controllable_DEQ & ~n37855;
  assign n37857 = ~n9921 & ~n37856;
  assign n37858 = i_FULL & ~n37857;
  assign n37859 = ~n7302 & ~n11311;
  assign n37860 = controllable_BtoR_REQ1 & ~n37859;
  assign n37861 = ~n9927 & ~n37860;
  assign n37862 = ~controllable_BtoR_REQ0 & ~n37861;
  assign n37863 = ~controllable_BtoR_REQ0 & ~n37862;
  assign n37864 = ~i_RtoB_ACK0 & ~n37863;
  assign n37865 = ~n37848 & ~n37864;
  assign n37866 = controllable_DEQ & ~n37865;
  assign n37867 = ~n9943 & ~n37866;
  assign n37868 = ~i_FULL & ~n37867;
  assign n37869 = ~n37858 & ~n37868;
  assign n37870 = i_nEMPTY & ~n37869;
  assign n37871 = ~n7330 & ~n11341;
  assign n37872 = controllable_BtoR_REQ1 & ~n37871;
  assign n37873 = ~n9951 & ~n37872;
  assign n37874 = ~controllable_BtoR_REQ0 & ~n37873;
  assign n37875 = ~controllable_BtoR_REQ0 & ~n37874;
  assign n37876 = ~i_RtoB_ACK0 & ~n37875;
  assign n37877 = ~i_RtoB_ACK0 & ~n37876;
  assign n37878 = controllable_DEQ & ~n37877;
  assign n37879 = ~n9969 & ~n37878;
  assign n37880 = i_FULL & ~n37879;
  assign n37881 = ~n7278 & ~n11324;
  assign n37882 = controllable_BtoR_REQ1 & ~n37881;
  assign n37883 = ~n9973 & ~n37882;
  assign n37884 = ~controllable_BtoR_REQ0 & ~n37883;
  assign n37885 = ~controllable_BtoR_REQ0 & ~n37884;
  assign n37886 = ~i_RtoB_ACK0 & ~n37885;
  assign n37887 = ~i_RtoB_ACK0 & ~n37886;
  assign n37888 = controllable_DEQ & ~n37887;
  assign n37889 = ~n9989 & ~n37888;
  assign n37890 = ~i_FULL & ~n37889;
  assign n37891 = ~n37880 & ~n37890;
  assign n37892 = ~i_nEMPTY & ~n37891;
  assign n37893 = ~n37870 & ~n37892;
  assign n37894 = ~controllable_BtoS_ACK0 & ~n37893;
  assign n37895 = ~n9870 & ~n37894;
  assign n37896 = ~n4465 & ~n37895;
  assign n37897 = ~n37842 & ~n37896;
  assign n37898 = ~i_StoB_REQ10 & ~n37897;
  assign n37899 = ~n37152 & ~n37898;
  assign n37900 = controllable_BtoS_ACK10 & ~n37899;
  assign n37901 = ~n5237 & ~n36638;
  assign n37902 = controllable_BtoR_REQ1 & ~n37901;
  assign n37903 = ~n12549 & ~n37902;
  assign n37904 = ~controllable_BtoR_REQ0 & ~n37903;
  assign n37905 = ~controllable_BtoR_REQ0 & ~n37904;
  assign n37906 = i_RtoB_ACK0 & ~n37905;
  assign n37907 = ~n10149 & ~n11666;
  assign n37908 = controllable_BtoR_REQ1 & ~n37907;
  assign n37909 = ~n12585 & ~n37908;
  assign n37910 = ~controllable_BtoR_REQ0 & ~n37909;
  assign n37911 = ~controllable_BtoR_REQ0 & ~n37910;
  assign n37912 = ~i_RtoB_ACK0 & ~n37911;
  assign n37913 = ~n37906 & ~n37912;
  assign n37914 = controllable_DEQ & ~n37913;
  assign n37915 = ~i_RtoB_ACK1 & ~n37467;
  assign n37916 = ~n11684 & ~n37915;
  assign n37917 = ~controllable_BtoR_REQ1 & ~n37916;
  assign n37918 = ~n36658 & ~n37917;
  assign n37919 = ~controllable_BtoR_REQ0 & ~n37918;
  assign n37920 = ~controllable_BtoR_REQ0 & ~n37919;
  assign n37921 = i_RtoB_ACK0 & ~n37920;
  assign n37922 = ~n37474 & ~n37921;
  assign n37923 = ~controllable_DEQ & ~n37922;
  assign n37924 = ~n37914 & ~n37923;
  assign n37925 = i_FULL & ~n37924;
  assign n37926 = ~n10149 & ~n11701;
  assign n37927 = controllable_BtoR_REQ1 & ~n37926;
  assign n37928 = ~n12585 & ~n37927;
  assign n37929 = ~controllable_BtoR_REQ0 & ~n37928;
  assign n37930 = ~controllable_BtoR_REQ0 & ~n37929;
  assign n37931 = ~i_RtoB_ACK0 & ~n37930;
  assign n37932 = ~n37906 & ~n37931;
  assign n37933 = controllable_DEQ & ~n37932;
  assign n37934 = ~n37497 & ~n37921;
  assign n37935 = ~controllable_DEQ & ~n37934;
  assign n37936 = ~n37933 & ~n37935;
  assign n37937 = ~i_FULL & ~n37936;
  assign n37938 = ~n37925 & ~n37937;
  assign n37939 = i_nEMPTY & ~n37938;
  assign n37940 = ~n7574 & ~n11730;
  assign n37941 = controllable_BtoR_REQ1 & ~n37940;
  assign n37942 = ~n10049 & ~n37941;
  assign n37943 = ~controllable_BtoR_REQ0 & ~n37942;
  assign n37944 = ~controllable_BtoR_REQ0 & ~n37943;
  assign n37945 = ~i_RtoB_ACK0 & ~n37944;
  assign n37946 = ~i_RtoB_ACK0 & ~n37945;
  assign n37947 = controllable_DEQ & ~n37946;
  assign n37948 = ~i_RtoB_ACK1 & ~n37526;
  assign n37949 = ~n11663 & ~n37948;
  assign n37950 = ~controllable_BtoR_REQ1 & ~n37949;
  assign n37951 = ~n36640 & ~n37950;
  assign n37952 = ~controllable_BtoR_REQ0 & ~n37951;
  assign n37953 = ~controllable_BtoR_REQ0 & ~n37952;
  assign n37954 = i_RtoB_ACK0 & ~n37953;
  assign n37955 = ~n37533 & ~n37954;
  assign n37956 = ~controllable_DEQ & ~n37955;
  assign n37957 = ~n37947 & ~n37956;
  assign n37958 = i_FULL & ~n37957;
  assign n37959 = ~n7563 & ~n11701;
  assign n37960 = controllable_BtoR_REQ1 & ~n37959;
  assign n37961 = ~n10061 & ~n37960;
  assign n37962 = ~controllable_BtoR_REQ0 & ~n37961;
  assign n37963 = ~controllable_BtoR_REQ0 & ~n37962;
  assign n37964 = ~i_RtoB_ACK0 & ~n37963;
  assign n37965 = ~i_RtoB_ACK0 & ~n37964;
  assign n37966 = controllable_DEQ & ~n37965;
  assign n37967 = ~n36645 & ~n37525;
  assign n37968 = i_RtoB_ACK1 & ~n37967;
  assign n37969 = ~n11666 & ~n37968;
  assign n37970 = controllable_BtoR_REQ1 & ~n37969;
  assign n37971 = ~n11663 & ~n37491;
  assign n37972 = ~controllable_BtoR_REQ1 & ~n37971;
  assign n37973 = ~n37970 & ~n37972;
  assign n37974 = ~controllable_BtoR_REQ0 & ~n37973;
  assign n37975 = ~controllable_BtoR_REQ0 & ~n37974;
  assign n37976 = ~i_RtoB_ACK0 & ~n37975;
  assign n37977 = ~n37954 & ~n37976;
  assign n37978 = ~controllable_DEQ & ~n37977;
  assign n37979 = ~n37966 & ~n37978;
  assign n37980 = ~i_FULL & ~n37979;
  assign n37981 = ~n37958 & ~n37980;
  assign n37982 = ~i_nEMPTY & ~n37981;
  assign n37983 = ~n37939 & ~n37982;
  assign n37984 = controllable_BtoS_ACK0 & ~n37983;
  assign n37985 = ~n8861 & ~n36717;
  assign n37986 = controllable_BtoR_REQ1 & ~n37985;
  assign n37987 = ~n12645 & ~n37986;
  assign n37988 = ~controllable_BtoR_REQ0 & ~n37987;
  assign n37989 = ~controllable_BtoR_REQ0 & ~n37988;
  assign n37990 = i_RtoB_ACK0 & ~n37989;
  assign n37991 = ~n11813 & ~n12462;
  assign n37992 = controllable_BtoR_REQ1 & ~n37991;
  assign n37993 = ~n12681 & ~n37992;
  assign n37994 = ~controllable_BtoR_REQ0 & ~n37993;
  assign n37995 = ~controllable_BtoR_REQ0 & ~n37994;
  assign n37996 = ~i_RtoB_ACK0 & ~n37995;
  assign n37997 = ~n37990 & ~n37996;
  assign n37998 = controllable_DEQ & ~n37997;
  assign n37999 = ~i_RtoB_ACK1 & ~n37730;
  assign n38000 = ~n11831 & ~n37999;
  assign n38001 = ~controllable_BtoR_REQ1 & ~n38000;
  assign n38002 = ~n36737 & ~n38001;
  assign n38003 = ~controllable_BtoR_REQ0 & ~n38002;
  assign n38004 = ~controllable_BtoR_REQ0 & ~n38003;
  assign n38005 = i_RtoB_ACK0 & ~n38004;
  assign n38006 = ~n37737 & ~n38005;
  assign n38007 = ~controllable_DEQ & ~n38006;
  assign n38008 = ~n37998 & ~n38007;
  assign n38009 = i_FULL & ~n38008;
  assign n38010 = ~n11848 & ~n12462;
  assign n38011 = controllable_BtoR_REQ1 & ~n38010;
  assign n38012 = ~n12681 & ~n38011;
  assign n38013 = ~controllable_BtoR_REQ0 & ~n38012;
  assign n38014 = ~controllable_BtoR_REQ0 & ~n38013;
  assign n38015 = ~i_RtoB_ACK0 & ~n38014;
  assign n38016 = ~n37990 & ~n38015;
  assign n38017 = controllable_DEQ & ~n38016;
  assign n38018 = ~n37760 & ~n38005;
  assign n38019 = ~controllable_DEQ & ~n38018;
  assign n38020 = ~n38017 & ~n38019;
  assign n38021 = ~i_FULL & ~n38020;
  assign n38022 = ~n38009 & ~n38021;
  assign n38023 = i_nEMPTY & ~n38022;
  assign n38024 = ~n11580 & ~n11877;
  assign n38025 = controllable_BtoR_REQ1 & ~n38024;
  assign n38026 = ~n9951 & ~n38025;
  assign n38027 = ~controllable_BtoR_REQ0 & ~n38026;
  assign n38028 = ~controllable_BtoR_REQ0 & ~n38027;
  assign n38029 = ~i_RtoB_ACK0 & ~n38028;
  assign n38030 = ~i_RtoB_ACK0 & ~n38029;
  assign n38031 = controllable_DEQ & ~n38030;
  assign n38032 = ~i_RtoB_ACK1 & ~n37789;
  assign n38033 = ~n11810 & ~n38032;
  assign n38034 = ~controllable_BtoR_REQ1 & ~n38033;
  assign n38035 = ~n36719 & ~n38034;
  assign n38036 = ~controllable_BtoR_REQ0 & ~n38035;
  assign n38037 = ~controllable_BtoR_REQ0 & ~n38036;
  assign n38038 = i_RtoB_ACK0 & ~n38037;
  assign n38039 = ~n37796 & ~n38038;
  assign n38040 = ~controllable_DEQ & ~n38039;
  assign n38041 = ~n38031 & ~n38040;
  assign n38042 = i_FULL & ~n38041;
  assign n38043 = ~n8883 & ~n11848;
  assign n38044 = controllable_BtoR_REQ1 & ~n38043;
  assign n38045 = ~n9973 & ~n38044;
  assign n38046 = ~controllable_BtoR_REQ0 & ~n38045;
  assign n38047 = ~controllable_BtoR_REQ0 & ~n38046;
  assign n38048 = ~i_RtoB_ACK0 & ~n38047;
  assign n38049 = ~i_RtoB_ACK0 & ~n38048;
  assign n38050 = controllable_DEQ & ~n38049;
  assign n38051 = ~n36724 & ~n37788;
  assign n38052 = i_RtoB_ACK1 & ~n38051;
  assign n38053 = ~n11813 & ~n38052;
  assign n38054 = controllable_BtoR_REQ1 & ~n38053;
  assign n38055 = ~n11810 & ~n37754;
  assign n38056 = ~controllable_BtoR_REQ1 & ~n38055;
  assign n38057 = ~n38054 & ~n38056;
  assign n38058 = ~controllable_BtoR_REQ0 & ~n38057;
  assign n38059 = ~controllable_BtoR_REQ0 & ~n38058;
  assign n38060 = ~i_RtoB_ACK0 & ~n38059;
  assign n38061 = ~n38038 & ~n38060;
  assign n38062 = ~controllable_DEQ & ~n38061;
  assign n38063 = ~n38050 & ~n38062;
  assign n38064 = ~i_FULL & ~n38063;
  assign n38065 = ~n38042 & ~n38064;
  assign n38066 = ~i_nEMPTY & ~n38065;
  assign n38067 = ~n38023 & ~n38066;
  assign n38068 = ~controllable_BtoS_ACK0 & ~n38067;
  assign n38069 = ~n37984 & ~n38068;
  assign n38070 = n4465 & ~n38069;
  assign n38071 = ~n7608 & ~n8861;
  assign n38072 = controllable_BtoR_REQ1 & ~n38071;
  assign n38073 = ~n9873 & ~n38072;
  assign n38074 = ~controllable_BtoR_REQ0 & ~n38073;
  assign n38075 = ~controllable_BtoR_REQ0 & ~n38074;
  assign n38076 = i_RtoB_ACK0 & ~n38075;
  assign n38077 = ~n7268 & ~n12462;
  assign n38078 = controllable_BtoR_REQ1 & ~n38077;
  assign n38079 = ~n9927 & ~n38078;
  assign n38080 = ~controllable_BtoR_REQ0 & ~n38079;
  assign n38081 = ~controllable_BtoR_REQ0 & ~n38080;
  assign n38082 = ~i_RtoB_ACK0 & ~n38081;
  assign n38083 = ~n38076 & ~n38082;
  assign n38084 = controllable_DEQ & ~n38083;
  assign n38085 = ~n10210 & ~n38084;
  assign n38086 = i_FULL & ~n38085;
  assign n38087 = ~n7305 & ~n12462;
  assign n38088 = controllable_BtoR_REQ1 & ~n38087;
  assign n38089 = ~n9927 & ~n38088;
  assign n38090 = ~controllable_BtoR_REQ0 & ~n38089;
  assign n38091 = ~controllable_BtoR_REQ0 & ~n38090;
  assign n38092 = ~i_RtoB_ACK0 & ~n38091;
  assign n38093 = ~n38076 & ~n38092;
  assign n38094 = controllable_DEQ & ~n38093;
  assign n38095 = ~n10222 & ~n38094;
  assign n38096 = ~i_FULL & ~n38095;
  assign n38097 = ~n38086 & ~n38096;
  assign n38098 = i_nEMPTY & ~n38097;
  assign n38099 = ~n7334 & ~n11580;
  assign n38100 = controllable_BtoR_REQ1 & ~n38099;
  assign n38101 = ~n9951 & ~n38100;
  assign n38102 = ~controllable_BtoR_REQ0 & ~n38101;
  assign n38103 = ~controllable_BtoR_REQ0 & ~n38102;
  assign n38104 = ~i_RtoB_ACK0 & ~n38103;
  assign n38105 = ~i_RtoB_ACK0 & ~n38104;
  assign n38106 = controllable_DEQ & ~n38105;
  assign n38107 = ~n10234 & ~n38106;
  assign n38108 = i_FULL & ~n38107;
  assign n38109 = ~n7305 & ~n8883;
  assign n38110 = controllable_BtoR_REQ1 & ~n38109;
  assign n38111 = ~n9973 & ~n38110;
  assign n38112 = ~controllable_BtoR_REQ0 & ~n38111;
  assign n38113 = ~controllable_BtoR_REQ0 & ~n38112;
  assign n38114 = ~i_RtoB_ACK0 & ~n38113;
  assign n38115 = ~i_RtoB_ACK0 & ~n38114;
  assign n38116 = controllable_DEQ & ~n38115;
  assign n38117 = ~n10243 & ~n38116;
  assign n38118 = ~i_FULL & ~n38117;
  assign n38119 = ~n38108 & ~n38118;
  assign n38120 = ~i_nEMPTY & ~n38119;
  assign n38121 = ~n38098 & ~n38120;
  assign n38122 = ~controllable_BtoS_ACK0 & ~n38121;
  assign n38123 = ~n10190 & ~n38122;
  assign n38124 = ~n4465 & ~n38123;
  assign n38125 = ~n38070 & ~n38124;
  assign n38126 = i_StoB_REQ10 & ~n38125;
  assign n38127 = ~n37898 & ~n38126;
  assign n38128 = ~controllable_BtoS_ACK10 & ~n38127;
  assign n38129 = ~n37900 & ~n38128;
  assign n38130 = n4464 & ~n38129;
  assign n38131 = ~n10290 & ~n10300;
  assign n38132 = i_FULL & ~n38131;
  assign n38133 = ~n10310 & ~n38132;
  assign n38134 = i_nEMPTY & ~n38133;
  assign n38135 = ~n10349 & ~n38134;
  assign n38136 = controllable_BtoS_ACK0 & ~n38135;
  assign n38137 = ~n10384 & ~n10394;
  assign n38138 = i_FULL & ~n38137;
  assign n38139 = ~n10404 & ~n38138;
  assign n38140 = i_nEMPTY & ~n38139;
  assign n38141 = ~n10443 & ~n38140;
  assign n38142 = ~controllable_BtoS_ACK0 & ~n38141;
  assign n38143 = ~n38136 & ~n38142;
  assign n38144 = n4465 & ~n38143;
  assign n38145 = ~n5307 & ~n38142;
  assign n38146 = ~n4465 & ~n38145;
  assign n38147 = ~n38144 & ~n38146;
  assign n38148 = i_StoB_REQ10 & ~n38147;
  assign n38149 = ~n7054 & ~n7903;
  assign n38150 = controllable_BtoR_REQ1 & ~n38149;
  assign n38151 = ~n10462 & ~n38150;
  assign n38152 = ~controllable_BtoR_REQ0 & ~n38151;
  assign n38153 = ~controllable_BtoR_REQ0 & ~n38152;
  assign n38154 = i_RtoB_ACK0 & ~n38153;
  assign n38155 = ~n7932 & ~n9789;
  assign n38156 = controllable_BtoR_REQ1 & ~n38155;
  assign n38157 = ~n10512 & ~n38156;
  assign n38158 = ~controllable_BtoR_REQ0 & ~n38157;
  assign n38159 = ~controllable_BtoR_REQ0 & ~n38158;
  assign n38160 = ~i_RtoB_ACK0 & ~n38159;
  assign n38161 = ~n38154 & ~n38160;
  assign n38162 = controllable_DEQ & ~n38161;
  assign n38163 = ~n10504 & ~n38162;
  assign n38164 = i_FULL & ~n38163;
  assign n38165 = ~n7972 & ~n9789;
  assign n38166 = controllable_BtoR_REQ1 & ~n38165;
  assign n38167 = ~n10512 & ~n38166;
  assign n38168 = ~controllable_BtoR_REQ0 & ~n38167;
  assign n38169 = ~controllable_BtoR_REQ0 & ~n38168;
  assign n38170 = ~i_RtoB_ACK0 & ~n38169;
  assign n38171 = ~n38154 & ~n38170;
  assign n38172 = controllable_DEQ & ~n38171;
  assign n38173 = ~n10530 & ~n38172;
  assign n38174 = ~i_FULL & ~n38173;
  assign n38175 = ~n38164 & ~n38174;
  assign n38176 = i_nEMPTY & ~n38175;
  assign n38177 = ~n7127 & ~n8000;
  assign n38178 = controllable_BtoR_REQ1 & ~n38177;
  assign n38179 = ~n10538 & ~n38178;
  assign n38180 = ~controllable_BtoR_REQ0 & ~n38179;
  assign n38181 = ~controllable_BtoR_REQ0 & ~n38180;
  assign n38182 = ~i_RtoB_ACK0 & ~n38181;
  assign n38183 = ~i_RtoB_ACK0 & ~n38182;
  assign n38184 = controllable_DEQ & ~n38183;
  assign n38185 = ~n10556 & ~n38184;
  assign n38186 = i_FULL & ~n38185;
  assign n38187 = ~n7111 & ~n7948;
  assign n38188 = controllable_BtoR_REQ1 & ~n38187;
  assign n38189 = ~n10560 & ~n38188;
  assign n38190 = ~controllable_BtoR_REQ0 & ~n38189;
  assign n38191 = ~controllable_BtoR_REQ0 & ~n38190;
  assign n38192 = ~i_RtoB_ACK0 & ~n38191;
  assign n38193 = ~i_RtoB_ACK0 & ~n38192;
  assign n38194 = controllable_DEQ & ~n38193;
  assign n38195 = ~n10576 & ~n38194;
  assign n38196 = ~i_FULL & ~n38195;
  assign n38197 = ~n38186 & ~n38196;
  assign n38198 = ~i_nEMPTY & ~n38197;
  assign n38199 = ~n38176 & ~n38198;
  assign n38200 = controllable_BtoS_ACK0 & ~n38199;
  assign n38201 = ~n8072 & ~n11299;
  assign n38202 = controllable_BtoR_REQ1 & ~n38201;
  assign n38203 = ~n10592 & ~n38202;
  assign n38204 = ~controllable_BtoR_REQ0 & ~n38203;
  assign n38205 = ~controllable_BtoR_REQ0 & ~n38204;
  assign n38206 = i_RtoB_ACK0 & ~n38205;
  assign n38207 = ~n8096 & ~n11311;
  assign n38208 = controllable_BtoR_REQ1 & ~n38207;
  assign n38209 = ~n10639 & ~n38208;
  assign n38210 = ~controllable_BtoR_REQ0 & ~n38209;
  assign n38211 = ~controllable_BtoR_REQ0 & ~n38210;
  assign n38212 = ~i_RtoB_ACK0 & ~n38211;
  assign n38213 = ~n38206 & ~n38212;
  assign n38214 = controllable_DEQ & ~n38213;
  assign n38215 = ~n10631 & ~n38214;
  assign n38216 = i_FULL & ~n38215;
  assign n38217 = ~n8136 & ~n11311;
  assign n38218 = controllable_BtoR_REQ1 & ~n38217;
  assign n38219 = ~n10639 & ~n38218;
  assign n38220 = ~controllable_BtoR_REQ0 & ~n38219;
  assign n38221 = ~controllable_BtoR_REQ0 & ~n38220;
  assign n38222 = ~i_RtoB_ACK0 & ~n38221;
  assign n38223 = ~n38206 & ~n38222;
  assign n38224 = controllable_DEQ & ~n38223;
  assign n38225 = ~n10657 & ~n38224;
  assign n38226 = ~i_FULL & ~n38225;
  assign n38227 = ~n38216 & ~n38226;
  assign n38228 = i_nEMPTY & ~n38227;
  assign n38229 = ~n8164 & ~n11341;
  assign n38230 = controllable_BtoR_REQ1 & ~n38229;
  assign n38231 = ~n10665 & ~n38230;
  assign n38232 = ~controllable_BtoR_REQ0 & ~n38231;
  assign n38233 = ~controllable_BtoR_REQ0 & ~n38232;
  assign n38234 = ~i_RtoB_ACK0 & ~n38233;
  assign n38235 = ~i_RtoB_ACK0 & ~n38234;
  assign n38236 = controllable_DEQ & ~n38235;
  assign n38237 = ~n10683 & ~n38236;
  assign n38238 = i_FULL & ~n38237;
  assign n38239 = ~n8112 & ~n11324;
  assign n38240 = controllable_BtoR_REQ1 & ~n38239;
  assign n38241 = ~n10687 & ~n38240;
  assign n38242 = ~controllable_BtoR_REQ0 & ~n38241;
  assign n38243 = ~controllable_BtoR_REQ0 & ~n38242;
  assign n38244 = ~i_RtoB_ACK0 & ~n38243;
  assign n38245 = ~i_RtoB_ACK0 & ~n38244;
  assign n38246 = controllable_DEQ & ~n38245;
  assign n38247 = ~n10703 & ~n38246;
  assign n38248 = ~i_FULL & ~n38247;
  assign n38249 = ~n38238 & ~n38248;
  assign n38250 = ~i_nEMPTY & ~n38249;
  assign n38251 = ~n38228 & ~n38250;
  assign n38252 = ~controllable_BtoS_ACK0 & ~n38251;
  assign n38253 = ~n38200 & ~n38252;
  assign n38254 = n4465 & ~n38253;
  assign n38255 = ~n8319 & ~n11299;
  assign n38256 = controllable_BtoR_REQ1 & ~n38255;
  assign n38257 = ~n10782 & ~n38256;
  assign n38258 = ~controllable_BtoR_REQ0 & ~n38257;
  assign n38259 = ~controllable_BtoR_REQ0 & ~n38258;
  assign n38260 = i_RtoB_ACK0 & ~n38259;
  assign n38261 = ~n8337 & ~n11311;
  assign n38262 = controllable_BtoR_REQ1 & ~n38261;
  assign n38263 = ~n10818 & ~n38262;
  assign n38264 = ~controllable_BtoR_REQ0 & ~n38263;
  assign n38265 = ~controllable_BtoR_REQ0 & ~n38264;
  assign n38266 = ~i_RtoB_ACK0 & ~n38265;
  assign n38267 = ~n38260 & ~n38266;
  assign n38268 = controllable_DEQ & ~n38267;
  assign n38269 = ~n10812 & ~n38268;
  assign n38270 = i_FULL & ~n38269;
  assign n38271 = ~n8375 & ~n11311;
  assign n38272 = controllable_BtoR_REQ1 & ~n38271;
  assign n38273 = ~n10818 & ~n38272;
  assign n38274 = ~controllable_BtoR_REQ0 & ~n38273;
  assign n38275 = ~controllable_BtoR_REQ0 & ~n38274;
  assign n38276 = ~i_RtoB_ACK0 & ~n38275;
  assign n38277 = ~n38260 & ~n38276;
  assign n38278 = controllable_DEQ & ~n38277;
  assign n38279 = ~n10834 & ~n38278;
  assign n38280 = ~i_FULL & ~n38279;
  assign n38281 = ~n38270 & ~n38280;
  assign n38282 = i_nEMPTY & ~n38281;
  assign n38283 = ~n8403 & ~n11341;
  assign n38284 = controllable_BtoR_REQ1 & ~n38283;
  assign n38285 = ~n9951 & ~n38284;
  assign n38286 = ~controllable_BtoR_REQ0 & ~n38285;
  assign n38287 = ~controllable_BtoR_REQ0 & ~n38286;
  assign n38288 = ~i_RtoB_ACK0 & ~n38287;
  assign n38289 = ~i_RtoB_ACK0 & ~n38288;
  assign n38290 = controllable_DEQ & ~n38289;
  assign n38291 = ~n10852 & ~n38290;
  assign n38292 = i_FULL & ~n38291;
  assign n38293 = ~n8353 & ~n11324;
  assign n38294 = controllable_BtoR_REQ1 & ~n38293;
  assign n38295 = ~n9973 & ~n38294;
  assign n38296 = ~controllable_BtoR_REQ0 & ~n38295;
  assign n38297 = ~controllable_BtoR_REQ0 & ~n38296;
  assign n38298 = ~i_RtoB_ACK0 & ~n38297;
  assign n38299 = ~i_RtoB_ACK0 & ~n38298;
  assign n38300 = controllable_DEQ & ~n38299;
  assign n38301 = ~n10868 & ~n38300;
  assign n38302 = ~i_FULL & ~n38301;
  assign n38303 = ~n38292 & ~n38302;
  assign n38304 = ~i_nEMPTY & ~n38303;
  assign n38305 = ~n38282 & ~n38304;
  assign n38306 = ~controllable_BtoS_ACK0 & ~n38305;
  assign n38307 = ~n10780 & ~n38306;
  assign n38308 = ~n4465 & ~n38307;
  assign n38309 = ~n38254 & ~n38308;
  assign n38310 = ~i_StoB_REQ10 & ~n38309;
  assign n38311 = ~n38148 & ~n38310;
  assign n38312 = controllable_BtoS_ACK10 & ~n38311;
  assign n38313 = ~n5237 & ~n8462;
  assign n38314 = controllable_BtoR_REQ1 & ~n38313;
  assign n38315 = ~n10882 & ~n38314;
  assign n38316 = ~controllable_BtoR_REQ0 & ~n38315;
  assign n38317 = ~controllable_BtoR_REQ0 & ~n38316;
  assign n38318 = i_RtoB_ACK0 & ~n38317;
  assign n38319 = ~n7938 & ~n10149;
  assign n38320 = controllable_BtoR_REQ1 & ~n38319;
  assign n38321 = ~n10912 & ~n38320;
  assign n38322 = ~controllable_BtoR_REQ0 & ~n38321;
  assign n38323 = ~controllable_BtoR_REQ0 & ~n38322;
  assign n38324 = ~i_RtoB_ACK0 & ~n38323;
  assign n38325 = ~n38318 & ~n38324;
  assign n38326 = controllable_DEQ & ~n38325;
  assign n38327 = ~n10906 & ~n38326;
  assign n38328 = i_FULL & ~n38327;
  assign n38329 = ~n7975 & ~n10149;
  assign n38330 = controllable_BtoR_REQ1 & ~n38329;
  assign n38331 = ~n10912 & ~n38330;
  assign n38332 = ~controllable_BtoR_REQ0 & ~n38331;
  assign n38333 = ~controllable_BtoR_REQ0 & ~n38332;
  assign n38334 = ~i_RtoB_ACK0 & ~n38333;
  assign n38335 = ~n38318 & ~n38334;
  assign n38336 = controllable_DEQ & ~n38335;
  assign n38337 = ~n10920 & ~n38336;
  assign n38338 = ~i_FULL & ~n38337;
  assign n38339 = ~n38328 & ~n38338;
  assign n38340 = i_nEMPTY & ~n38339;
  assign n38341 = ~n7574 & ~n8004;
  assign n38342 = controllable_BtoR_REQ1 & ~n38341;
  assign n38343 = ~n10049 & ~n38342;
  assign n38344 = ~controllable_BtoR_REQ0 & ~n38343;
  assign n38345 = ~controllable_BtoR_REQ0 & ~n38344;
  assign n38346 = ~i_RtoB_ACK0 & ~n38345;
  assign n38347 = ~i_RtoB_ACK0 & ~n38346;
  assign n38348 = controllable_DEQ & ~n38347;
  assign n38349 = ~n10932 & ~n38348;
  assign n38350 = i_FULL & ~n38349;
  assign n38351 = ~n7563 & ~n7975;
  assign n38352 = controllable_BtoR_REQ1 & ~n38351;
  assign n38353 = ~n10061 & ~n38352;
  assign n38354 = ~controllable_BtoR_REQ0 & ~n38353;
  assign n38355 = ~controllable_BtoR_REQ0 & ~n38354;
  assign n38356 = ~i_RtoB_ACK0 & ~n38355;
  assign n38357 = ~i_RtoB_ACK0 & ~n38356;
  assign n38358 = controllable_DEQ & ~n38357;
  assign n38359 = ~n10941 & ~n38358;
  assign n38360 = ~i_FULL & ~n38359;
  assign n38361 = ~n38350 & ~n38360;
  assign n38362 = ~i_nEMPTY & ~n38361;
  assign n38363 = ~n38340 & ~n38362;
  assign n38364 = controllable_BtoS_ACK0 & ~n38363;
  assign n38365 = ~n8541 & ~n8861;
  assign n38366 = controllable_BtoR_REQ1 & ~n38365;
  assign n38367 = ~n10949 & ~n38366;
  assign n38368 = ~controllable_BtoR_REQ0 & ~n38367;
  assign n38369 = ~controllable_BtoR_REQ0 & ~n38368;
  assign n38370 = i_RtoB_ACK0 & ~n38369;
  assign n38371 = ~n8102 & ~n12462;
  assign n38372 = controllable_BtoR_REQ1 & ~n38371;
  assign n38373 = ~n10979 & ~n38372;
  assign n38374 = ~controllable_BtoR_REQ0 & ~n38373;
  assign n38375 = ~controllable_BtoR_REQ0 & ~n38374;
  assign n38376 = ~i_RtoB_ACK0 & ~n38375;
  assign n38377 = ~n38370 & ~n38376;
  assign n38378 = controllable_DEQ & ~n38377;
  assign n38379 = ~n10973 & ~n38378;
  assign n38380 = i_FULL & ~n38379;
  assign n38381 = ~n8139 & ~n12462;
  assign n38382 = controllable_BtoR_REQ1 & ~n38381;
  assign n38383 = ~n10979 & ~n38382;
  assign n38384 = ~controllable_BtoR_REQ0 & ~n38383;
  assign n38385 = ~controllable_BtoR_REQ0 & ~n38384;
  assign n38386 = ~i_RtoB_ACK0 & ~n38385;
  assign n38387 = ~n38370 & ~n38386;
  assign n38388 = controllable_DEQ & ~n38387;
  assign n38389 = ~n10987 & ~n38388;
  assign n38390 = ~i_FULL & ~n38389;
  assign n38391 = ~n38380 & ~n38390;
  assign n38392 = i_nEMPTY & ~n38391;
  assign n38393 = ~n8168 & ~n11580;
  assign n38394 = controllable_BtoR_REQ1 & ~n38393;
  assign n38395 = ~n9951 & ~n38394;
  assign n38396 = ~controllable_BtoR_REQ0 & ~n38395;
  assign n38397 = ~controllable_BtoR_REQ0 & ~n38396;
  assign n38398 = ~i_RtoB_ACK0 & ~n38397;
  assign n38399 = ~i_RtoB_ACK0 & ~n38398;
  assign n38400 = controllable_DEQ & ~n38399;
  assign n38401 = ~n10999 & ~n38400;
  assign n38402 = i_FULL & ~n38401;
  assign n38403 = ~n8139 & ~n8883;
  assign n38404 = controllable_BtoR_REQ1 & ~n38403;
  assign n38405 = ~n9973 & ~n38404;
  assign n38406 = ~controllable_BtoR_REQ0 & ~n38405;
  assign n38407 = ~controllable_BtoR_REQ0 & ~n38406;
  assign n38408 = ~i_RtoB_ACK0 & ~n38407;
  assign n38409 = ~i_RtoB_ACK0 & ~n38408;
  assign n38410 = controllable_DEQ & ~n38409;
  assign n38411 = ~n11008 & ~n38410;
  assign n38412 = ~i_FULL & ~n38411;
  assign n38413 = ~n38402 & ~n38412;
  assign n38414 = ~i_nEMPTY & ~n38413;
  assign n38415 = ~n38392 & ~n38414;
  assign n38416 = ~controllable_BtoS_ACK0 & ~n38415;
  assign n38417 = ~n38364 & ~n38416;
  assign n38418 = n4465 & ~n38417;
  assign n38419 = ~n8673 & ~n8861;
  assign n38420 = controllable_BtoR_REQ1 & ~n38419;
  assign n38421 = ~n10782 & ~n38420;
  assign n38422 = ~controllable_BtoR_REQ0 & ~n38421;
  assign n38423 = ~controllable_BtoR_REQ0 & ~n38422;
  assign n38424 = i_RtoB_ACK0 & ~n38423;
  assign n38425 = ~n8343 & ~n12462;
  assign n38426 = controllable_BtoR_REQ1 & ~n38425;
  assign n38427 = ~n10818 & ~n38426;
  assign n38428 = ~controllable_BtoR_REQ0 & ~n38427;
  assign n38429 = ~controllable_BtoR_REQ0 & ~n38428;
  assign n38430 = ~i_RtoB_ACK0 & ~n38429;
  assign n38431 = ~n38424 & ~n38430;
  assign n38432 = controllable_DEQ & ~n38431;
  assign n38433 = ~n11079 & ~n38432;
  assign n38434 = i_FULL & ~n38433;
  assign n38435 = ~n8378 & ~n12462;
  assign n38436 = controllable_BtoR_REQ1 & ~n38435;
  assign n38437 = ~n10818 & ~n38436;
  assign n38438 = ~controllable_BtoR_REQ0 & ~n38437;
  assign n38439 = ~controllable_BtoR_REQ0 & ~n38438;
  assign n38440 = ~i_RtoB_ACK0 & ~n38439;
  assign n38441 = ~n38424 & ~n38440;
  assign n38442 = controllable_DEQ & ~n38441;
  assign n38443 = ~n11091 & ~n38442;
  assign n38444 = ~i_FULL & ~n38443;
  assign n38445 = ~n38434 & ~n38444;
  assign n38446 = i_nEMPTY & ~n38445;
  assign n38447 = ~n8407 & ~n11580;
  assign n38448 = controllable_BtoR_REQ1 & ~n38447;
  assign n38449 = ~n9951 & ~n38448;
  assign n38450 = ~controllable_BtoR_REQ0 & ~n38449;
  assign n38451 = ~controllable_BtoR_REQ0 & ~n38450;
  assign n38452 = ~i_RtoB_ACK0 & ~n38451;
  assign n38453 = ~i_RtoB_ACK0 & ~n38452;
  assign n38454 = controllable_DEQ & ~n38453;
  assign n38455 = ~n11103 & ~n38454;
  assign n38456 = i_FULL & ~n38455;
  assign n38457 = ~n8378 & ~n8883;
  assign n38458 = controllable_BtoR_REQ1 & ~n38457;
  assign n38459 = ~n9973 & ~n38458;
  assign n38460 = ~controllable_BtoR_REQ0 & ~n38459;
  assign n38461 = ~controllable_BtoR_REQ0 & ~n38460;
  assign n38462 = ~i_RtoB_ACK0 & ~n38461;
  assign n38463 = ~i_RtoB_ACK0 & ~n38462;
  assign n38464 = controllable_DEQ & ~n38463;
  assign n38465 = ~n11112 & ~n38464;
  assign n38466 = ~i_FULL & ~n38465;
  assign n38467 = ~n38456 & ~n38466;
  assign n38468 = ~i_nEMPTY & ~n38467;
  assign n38469 = ~n38446 & ~n38468;
  assign n38470 = ~controllable_BtoS_ACK0 & ~n38469;
  assign n38471 = ~n11059 & ~n38470;
  assign n38472 = ~n4465 & ~n38471;
  assign n38473 = ~n38418 & ~n38472;
  assign n38474 = i_StoB_REQ10 & ~n38473;
  assign n38475 = ~n38310 & ~n38474;
  assign n38476 = ~controllable_BtoS_ACK10 & ~n38475;
  assign n38477 = ~n38312 & ~n38476;
  assign n38478 = ~n4464 & ~n38477;
  assign n38479 = ~n38130 & ~n38478;
  assign n38480 = ~n4463 & ~n38479;
  assign n38481 = ~n36798 & ~n38480;
  assign n38482 = n4462 & ~n38481;
  assign n38483 = ~n12363 & ~n12401;
  assign n38484 = ~controllable_BtoR_REQ0 & ~n38483;
  assign n38485 = ~controllable_BtoR_REQ0 & ~n38484;
  assign n38486 = ~i_RtoB_ACK0 & ~n38485;
  assign n38487 = ~n12361 & ~n38486;
  assign n38488 = controllable_DEQ & ~n38487;
  assign n38489 = ~n12395 & ~n38488;
  assign n38490 = i_FULL & ~n38489;
  assign n38491 = ~n12419 & ~n38490;
  assign n38492 = i_nEMPTY & ~n38491;
  assign n38493 = ~n12452 & ~n38492;
  assign n38494 = controllable_BtoS_ACK0 & ~n38493;
  assign n38495 = ~n12464 & ~n12492;
  assign n38496 = ~controllable_BtoR_REQ0 & ~n38495;
  assign n38497 = ~controllable_BtoR_REQ0 & ~n38496;
  assign n38498 = ~i_RtoB_ACK0 & ~n38497;
  assign n38499 = ~n12460 & ~n38498;
  assign n38500 = controllable_DEQ & ~n38499;
  assign n38501 = ~n12486 & ~n38500;
  assign n38502 = i_FULL & ~n38501;
  assign n38503 = ~n12510 & ~n38502;
  assign n38504 = i_nEMPTY & ~n38503;
  assign n38505 = ~n12539 & ~n38504;
  assign n38506 = ~controllable_BtoS_ACK0 & ~n38505;
  assign n38507 = ~n38494 & ~n38506;
  assign n38508 = n4465 & ~n38507;
  assign n38509 = ~n10190 & ~n38506;
  assign n38510 = ~n4465 & ~n38509;
  assign n38511 = ~n38508 & ~n38510;
  assign n38512 = i_StoB_REQ10 & ~n38511;
  assign n38513 = ~n12549 & ~n37154;
  assign n38514 = ~controllable_BtoR_REQ0 & ~n38513;
  assign n38515 = ~controllable_BtoR_REQ0 & ~n38514;
  assign n38516 = i_RtoB_ACK0 & ~n38515;
  assign n38517 = ~n12585 & ~n37256;
  assign n38518 = ~controllable_BtoR_REQ0 & ~n38517;
  assign n38519 = ~controllable_BtoR_REQ0 & ~n38518;
  assign n38520 = ~i_RtoB_ACK0 & ~n38519;
  assign n38521 = ~n38516 & ~n38520;
  assign n38522 = controllable_DEQ & ~n38521;
  assign n38523 = ~n12579 & ~n38522;
  assign n38524 = i_FULL & ~n38523;
  assign n38525 = ~n12585 & ~n37480;
  assign n38526 = ~controllable_BtoR_REQ0 & ~n38525;
  assign n38527 = ~controllable_BtoR_REQ0 & ~n38526;
  assign n38528 = ~i_RtoB_ACK0 & ~n38527;
  assign n38529 = ~n38516 & ~n38528;
  assign n38530 = controllable_DEQ & ~n38529;
  assign n38531 = ~n12601 & ~n38530;
  assign n38532 = ~i_FULL & ~n38531;
  assign n38533 = ~n38524 & ~n38532;
  assign n38534 = i_nEMPTY & ~n38533;
  assign n38535 = ~n10049 & ~n37505;
  assign n38536 = ~controllable_BtoR_REQ0 & ~n38535;
  assign n38537 = ~controllable_BtoR_REQ0 & ~n38536;
  assign n38538 = ~i_RtoB_ACK0 & ~n38537;
  assign n38539 = ~i_RtoB_ACK0 & ~n38538;
  assign n38540 = controllable_DEQ & ~n38539;
  assign n38541 = ~n12619 & ~n38540;
  assign n38542 = i_FULL & ~n38541;
  assign n38543 = ~n10061 & ~n37539;
  assign n38544 = ~controllable_BtoR_REQ0 & ~n38543;
  assign n38545 = ~controllable_BtoR_REQ0 & ~n38544;
  assign n38546 = ~i_RtoB_ACK0 & ~n38545;
  assign n38547 = ~i_RtoB_ACK0 & ~n38546;
  assign n38548 = controllable_DEQ & ~n38547;
  assign n38549 = ~n12637 & ~n38548;
  assign n38550 = ~i_FULL & ~n38549;
  assign n38551 = ~n38542 & ~n38550;
  assign n38552 = ~i_nEMPTY & ~n38551;
  assign n38553 = ~n38534 & ~n38552;
  assign n38554 = controllable_BtoS_ACK0 & ~n38553;
  assign n38555 = ~n12645 & ~n37680;
  assign n38556 = ~controllable_BtoR_REQ0 & ~n38555;
  assign n38557 = ~controllable_BtoR_REQ0 & ~n38556;
  assign n38558 = i_RtoB_ACK0 & ~n38557;
  assign n38559 = ~n12681 & ~n37698;
  assign n38560 = ~controllable_BtoR_REQ0 & ~n38559;
  assign n38561 = ~controllable_BtoR_REQ0 & ~n38560;
  assign n38562 = ~i_RtoB_ACK0 & ~n38561;
  assign n38563 = ~n38558 & ~n38562;
  assign n38564 = controllable_DEQ & ~n38563;
  assign n38565 = ~n12675 & ~n38564;
  assign n38566 = i_FULL & ~n38565;
  assign n38567 = ~n12681 & ~n37743;
  assign n38568 = ~controllable_BtoR_REQ0 & ~n38567;
  assign n38569 = ~controllable_BtoR_REQ0 & ~n38568;
  assign n38570 = ~i_RtoB_ACK0 & ~n38569;
  assign n38571 = ~n38558 & ~n38570;
  assign n38572 = controllable_DEQ & ~n38571;
  assign n38573 = ~n12697 & ~n38572;
  assign n38574 = ~i_FULL & ~n38573;
  assign n38575 = ~n38566 & ~n38574;
  assign n38576 = i_nEMPTY & ~n38575;
  assign n38577 = ~n9951 & ~n37768;
  assign n38578 = ~controllable_BtoR_REQ0 & ~n38577;
  assign n38579 = ~controllable_BtoR_REQ0 & ~n38578;
  assign n38580 = ~i_RtoB_ACK0 & ~n38579;
  assign n38581 = ~i_RtoB_ACK0 & ~n38580;
  assign n38582 = controllable_DEQ & ~n38581;
  assign n38583 = ~n12715 & ~n38582;
  assign n38584 = i_FULL & ~n38583;
  assign n38585 = ~n9973 & ~n37802;
  assign n38586 = ~controllable_BtoR_REQ0 & ~n38585;
  assign n38587 = ~controllable_BtoR_REQ0 & ~n38586;
  assign n38588 = ~i_RtoB_ACK0 & ~n38587;
  assign n38589 = ~i_RtoB_ACK0 & ~n38588;
  assign n38590 = controllable_DEQ & ~n38589;
  assign n38591 = ~n12731 & ~n38590;
  assign n38592 = ~i_FULL & ~n38591;
  assign n38593 = ~n38584 & ~n38592;
  assign n38594 = ~i_nEMPTY & ~n38593;
  assign n38595 = ~n38576 & ~n38594;
  assign n38596 = ~controllable_BtoS_ACK0 & ~n38595;
  assign n38597 = ~n38554 & ~n38596;
  assign n38598 = n4465 & ~n38597;
  assign n38599 = ~n12781 & ~n37894;
  assign n38600 = ~n4465 & ~n38599;
  assign n38601 = ~n38598 & ~n38600;
  assign n38602 = ~i_StoB_REQ10 & ~n38601;
  assign n38603 = ~n38512 & ~n38602;
  assign n38604 = ~controllable_BtoS_ACK10 & ~n38603;
  assign n38605 = ~n12355 & ~n38604;
  assign n38606 = n4464 & ~n38605;
  assign n38607 = ~n12865 & ~n12893;
  assign n38608 = ~controllable_BtoR_REQ0 & ~n38607;
  assign n38609 = ~controllable_BtoR_REQ0 & ~n38608;
  assign n38610 = ~i_RtoB_ACK0 & ~n38609;
  assign n38611 = ~n12863 & ~n38610;
  assign n38612 = controllable_DEQ & ~n38611;
  assign n38613 = ~n12887 & ~n38612;
  assign n38614 = i_FULL & ~n38613;
  assign n38615 = ~n12911 & ~n38614;
  assign n38616 = i_nEMPTY & ~n38615;
  assign n38617 = ~n12940 & ~n38616;
  assign n38618 = controllable_BtoS_ACK0 & ~n38617;
  assign n38619 = ~n12950 & ~n12978;
  assign n38620 = ~controllable_BtoR_REQ0 & ~n38619;
  assign n38621 = ~controllable_BtoR_REQ0 & ~n38620;
  assign n38622 = ~i_RtoB_ACK0 & ~n38621;
  assign n38623 = ~n12948 & ~n38622;
  assign n38624 = controllable_DEQ & ~n38623;
  assign n38625 = ~n12972 & ~n38624;
  assign n38626 = i_FULL & ~n38625;
  assign n38627 = ~n12996 & ~n38626;
  assign n38628 = i_nEMPTY & ~n38627;
  assign n38629 = ~n13025 & ~n38628;
  assign n38630 = ~controllable_BtoS_ACK0 & ~n38629;
  assign n38631 = ~n38618 & ~n38630;
  assign n38632 = n4465 & ~n38631;
  assign n38633 = ~n11059 & ~n38630;
  assign n38634 = ~n4465 & ~n38633;
  assign n38635 = ~n38632 & ~n38634;
  assign n38636 = i_StoB_REQ10 & ~n38635;
  assign n38637 = ~n10882 & ~n38150;
  assign n38638 = ~controllable_BtoR_REQ0 & ~n38637;
  assign n38639 = ~controllable_BtoR_REQ0 & ~n38638;
  assign n38640 = i_RtoB_ACK0 & ~n38639;
  assign n38641 = ~n10912 & ~n38156;
  assign n38642 = ~controllable_BtoR_REQ0 & ~n38641;
  assign n38643 = ~controllable_BtoR_REQ0 & ~n38642;
  assign n38644 = ~i_RtoB_ACK0 & ~n38643;
  assign n38645 = ~n38640 & ~n38644;
  assign n38646 = controllable_DEQ & ~n38645;
  assign n38647 = ~n13049 & ~n38646;
  assign n38648 = i_FULL & ~n38647;
  assign n38649 = ~n10912 & ~n38166;
  assign n38650 = ~controllable_BtoR_REQ0 & ~n38649;
  assign n38651 = ~controllable_BtoR_REQ0 & ~n38650;
  assign n38652 = ~i_RtoB_ACK0 & ~n38651;
  assign n38653 = ~n38640 & ~n38652;
  assign n38654 = controllable_DEQ & ~n38653;
  assign n38655 = ~n13059 & ~n38654;
  assign n38656 = ~i_FULL & ~n38655;
  assign n38657 = ~n38648 & ~n38656;
  assign n38658 = i_nEMPTY & ~n38657;
  assign n38659 = ~n10049 & ~n38178;
  assign n38660 = ~controllable_BtoR_REQ0 & ~n38659;
  assign n38661 = ~controllable_BtoR_REQ0 & ~n38660;
  assign n38662 = ~i_RtoB_ACK0 & ~n38661;
  assign n38663 = ~i_RtoB_ACK0 & ~n38662;
  assign n38664 = controllable_DEQ & ~n38663;
  assign n38665 = ~n13071 & ~n38664;
  assign n38666 = i_FULL & ~n38665;
  assign n38667 = ~n10061 & ~n38188;
  assign n38668 = ~controllable_BtoR_REQ0 & ~n38667;
  assign n38669 = ~controllable_BtoR_REQ0 & ~n38668;
  assign n38670 = ~i_RtoB_ACK0 & ~n38669;
  assign n38671 = ~i_RtoB_ACK0 & ~n38670;
  assign n38672 = controllable_DEQ & ~n38671;
  assign n38673 = ~n13081 & ~n38672;
  assign n38674 = ~i_FULL & ~n38673;
  assign n38675 = ~n38666 & ~n38674;
  assign n38676 = ~i_nEMPTY & ~n38675;
  assign n38677 = ~n38658 & ~n38676;
  assign n38678 = controllable_BtoS_ACK0 & ~n38677;
  assign n38679 = ~n10949 & ~n38202;
  assign n38680 = ~controllable_BtoR_REQ0 & ~n38679;
  assign n38681 = ~controllable_BtoR_REQ0 & ~n38680;
  assign n38682 = i_RtoB_ACK0 & ~n38681;
  assign n38683 = ~n10979 & ~n38208;
  assign n38684 = ~controllable_BtoR_REQ0 & ~n38683;
  assign n38685 = ~controllable_BtoR_REQ0 & ~n38684;
  assign n38686 = ~i_RtoB_ACK0 & ~n38685;
  assign n38687 = ~n38682 & ~n38686;
  assign n38688 = controllable_DEQ & ~n38687;
  assign n38689 = ~n13103 & ~n38688;
  assign n38690 = i_FULL & ~n38689;
  assign n38691 = ~n10979 & ~n38218;
  assign n38692 = ~controllable_BtoR_REQ0 & ~n38691;
  assign n38693 = ~controllable_BtoR_REQ0 & ~n38692;
  assign n38694 = ~i_RtoB_ACK0 & ~n38693;
  assign n38695 = ~n38682 & ~n38694;
  assign n38696 = controllable_DEQ & ~n38695;
  assign n38697 = ~n13113 & ~n38696;
  assign n38698 = ~i_FULL & ~n38697;
  assign n38699 = ~n38690 & ~n38698;
  assign n38700 = i_nEMPTY & ~n38699;
  assign n38701 = ~n9951 & ~n38230;
  assign n38702 = ~controllable_BtoR_REQ0 & ~n38701;
  assign n38703 = ~controllable_BtoR_REQ0 & ~n38702;
  assign n38704 = ~i_RtoB_ACK0 & ~n38703;
  assign n38705 = ~i_RtoB_ACK0 & ~n38704;
  assign n38706 = controllable_DEQ & ~n38705;
  assign n38707 = ~n13125 & ~n38706;
  assign n38708 = i_FULL & ~n38707;
  assign n38709 = ~n9973 & ~n38240;
  assign n38710 = ~controllable_BtoR_REQ0 & ~n38709;
  assign n38711 = ~controllable_BtoR_REQ0 & ~n38710;
  assign n38712 = ~i_RtoB_ACK0 & ~n38711;
  assign n38713 = ~i_RtoB_ACK0 & ~n38712;
  assign n38714 = controllable_DEQ & ~n38713;
  assign n38715 = ~n13135 & ~n38714;
  assign n38716 = ~i_FULL & ~n38715;
  assign n38717 = ~n38708 & ~n38716;
  assign n38718 = ~i_nEMPTY & ~n38717;
  assign n38719 = ~n38700 & ~n38718;
  assign n38720 = ~controllable_BtoS_ACK0 & ~n38719;
  assign n38721 = ~n38678 & ~n38720;
  assign n38722 = n4465 & ~n38721;
  assign n38723 = ~n38308 & ~n38722;
  assign n38724 = ~i_StoB_REQ10 & ~n38723;
  assign n38725 = ~n38636 & ~n38724;
  assign n38726 = ~controllable_BtoS_ACK10 & ~n38725;
  assign n38727 = ~n12857 & ~n38726;
  assign n38728 = ~n4464 & ~n38727;
  assign n38729 = ~n38606 & ~n38728;
  assign n38730 = ~n4463 & ~n38729;
  assign n38731 = ~n12155 & ~n38730;
  assign n38732 = ~n4462 & ~n38731;
  assign n38733 = ~n38482 & ~n38732;
  assign n38734 = n4461 & ~n38733;
  assign n38735 = ~n11172 & ~n36892;
  assign n38736 = ~controllable_DEQ & ~n38735;
  assign n38737 = ~n14081 & ~n38736;
  assign n38738 = i_nEMPTY & ~n38737;
  assign n38739 = ~n11149 & ~n36927;
  assign n38740 = ~controllable_DEQ & ~n38739;
  assign n38741 = ~n11194 & ~n38740;
  assign n38742 = i_FULL & ~n38741;
  assign n38743 = ~n14103 & ~n36933;
  assign n38744 = ~controllable_BtoR_REQ0 & ~n38743;
  assign n38745 = ~controllable_BtoR_REQ0 & ~n38744;
  assign n38746 = ~i_RtoB_ACK0 & ~n38745;
  assign n38747 = ~n11149 & ~n38746;
  assign n38748 = ~controllable_DEQ & ~n38747;
  assign n38749 = ~n11209 & ~n38748;
  assign n38750 = ~i_FULL & ~n38749;
  assign n38751 = ~n38742 & ~n38750;
  assign n38752 = ~i_nEMPTY & ~n38751;
  assign n38753 = ~n38738 & ~n38752;
  assign n38754 = controllable_BtoS_ACK0 & ~n38753;
  assign n38755 = ~n5365 & ~n37073;
  assign n38756 = ~controllable_DEQ & ~n38755;
  assign n38757 = ~n14124 & ~n38756;
  assign n38758 = i_nEMPTY & ~n38757;
  assign n38759 = ~n5342 & ~n37108;
  assign n38760 = ~controllable_DEQ & ~n38759;
  assign n38761 = ~n5387 & ~n38760;
  assign n38762 = i_FULL & ~n38761;
  assign n38763 = ~n13226 & ~n37114;
  assign n38764 = ~controllable_BtoR_REQ0 & ~n38763;
  assign n38765 = ~controllable_BtoR_REQ0 & ~n38764;
  assign n38766 = ~i_RtoB_ACK0 & ~n38765;
  assign n38767 = ~n5342 & ~n38766;
  assign n38768 = ~controllable_DEQ & ~n38767;
  assign n38769 = ~n5402 & ~n38768;
  assign n38770 = ~i_FULL & ~n38769;
  assign n38771 = ~n38762 & ~n38770;
  assign n38772 = ~i_nEMPTY & ~n38771;
  assign n38773 = ~n38758 & ~n38772;
  assign n38774 = ~controllable_BtoS_ACK0 & ~n38773;
  assign n38775 = ~n38754 & ~n38774;
  assign n38776 = n4465 & ~n38775;
  assign n38777 = ~n13240 & ~n38776;
  assign n38778 = i_StoB_REQ10 & ~n38777;
  assign n38779 = ~controllable_BtoS_ACK13 & ~n9275;
  assign n38780 = ~controllable_BtoS_ACK13 & ~n38779;
  assign n38781 = i_StoB_REQ13 & ~n38780;
  assign n38782 = i_StoB_REQ2 & ~n9153;
  assign n38783 = ~controllable_BtoS_ACK2 & ~n38782;
  assign n38784 = ~controllable_BtoS_ACK2 & ~n38783;
  assign n38785 = n4477 & ~n38784;
  assign n38786 = ~n5621 & ~n38785;
  assign n38787 = n4476 & ~n38786;
  assign n38788 = ~n36936 & ~n38787;
  assign n38789 = ~i_StoB_REQ3 & ~n38788;
  assign n38790 = ~i_StoB_REQ3 & ~n38789;
  assign n38791 = controllable_BtoS_ACK3 & ~n38790;
  assign n38792 = ~n9175 & ~n38789;
  assign n38793 = ~controllable_BtoS_ACK3 & ~n38792;
  assign n38794 = ~n38791 & ~n38793;
  assign n38795 = n4475 & ~n38794;
  assign n38796 = ~n36946 & ~n38795;
  assign n38797 = ~i_StoB_REQ4 & ~n38796;
  assign n38798 = ~i_StoB_REQ4 & ~n38797;
  assign n38799 = controllable_BtoS_ACK4 & ~n38798;
  assign n38800 = ~n9188 & ~n38797;
  assign n38801 = ~controllable_BtoS_ACK4 & ~n38800;
  assign n38802 = ~n38799 & ~n38801;
  assign n38803 = n4474 & ~n38802;
  assign n38804 = ~n36956 & ~n38803;
  assign n38805 = ~i_StoB_REQ5 & ~n38804;
  assign n38806 = ~i_StoB_REQ5 & ~n38805;
  assign n38807 = controllable_BtoS_ACK5 & ~n38806;
  assign n38808 = ~n9201 & ~n38805;
  assign n38809 = ~controllable_BtoS_ACK5 & ~n38808;
  assign n38810 = ~n38807 & ~n38809;
  assign n38811 = n4473 & ~n38810;
  assign n38812 = ~n36966 & ~n38811;
  assign n38813 = ~i_StoB_REQ8 & ~n38812;
  assign n38814 = ~i_StoB_REQ8 & ~n38813;
  assign n38815 = controllable_BtoS_ACK8 & ~n38814;
  assign n38816 = ~n9214 & ~n38813;
  assign n38817 = ~controllable_BtoS_ACK8 & ~n38816;
  assign n38818 = ~n38815 & ~n38817;
  assign n38819 = n4472 & ~n38818;
  assign n38820 = ~n36976 & ~n38819;
  assign n38821 = n4471 & ~n38820;
  assign n38822 = ~n4819 & ~n38821;
  assign n38823 = ~i_StoB_REQ6 & ~n38822;
  assign n38824 = ~i_StoB_REQ6 & ~n38823;
  assign n38825 = controllable_BtoS_ACK6 & ~n38824;
  assign n38826 = i_StoB_REQ6 & ~n9106;
  assign n38827 = ~n38823 & ~n38826;
  assign n38828 = ~controllable_BtoS_ACK6 & ~n38827;
  assign n38829 = ~n38825 & ~n38828;
  assign n38830 = ~i_StoB_REQ7 & ~n38829;
  assign n38831 = ~i_StoB_REQ7 & ~n38830;
  assign n38832 = controllable_BtoS_ACK7 & ~n38831;
  assign n38833 = ~n9235 & ~n38830;
  assign n38834 = ~controllable_BtoS_ACK7 & ~n38833;
  assign n38835 = ~n38832 & ~n38834;
  assign n38836 = n4470 & ~n38835;
  assign n38837 = ~n36995 & ~n38836;
  assign n38838 = n4469 & ~n38837;
  assign n38839 = ~n4876 & ~n38838;
  assign n38840 = ~i_StoB_REQ9 & ~n38839;
  assign n38841 = ~i_StoB_REQ9 & ~n38840;
  assign n38842 = controllable_BtoS_ACK9 & ~n38841;
  assign n38843 = i_StoB_REQ9 & ~n9123;
  assign n38844 = ~n38840 & ~n38843;
  assign n38845 = ~controllable_BtoS_ACK9 & ~n38844;
  assign n38846 = ~n38842 & ~n38845;
  assign n38847 = n4468 & ~n38846;
  assign n38848 = ~n4901 & ~n38847;
  assign n38849 = ~i_StoB_REQ11 & ~n38848;
  assign n38850 = ~i_StoB_REQ11 & ~n38849;
  assign n38851 = controllable_BtoS_ACK11 & ~n38850;
  assign n38852 = i_StoB_REQ11 & ~n9131;
  assign n38853 = ~n38849 & ~n38852;
  assign n38854 = ~controllable_BtoS_ACK11 & ~n38853;
  assign n38855 = ~n38851 & ~n38854;
  assign n38856 = n4467 & ~n38855;
  assign n38857 = ~n4931 & ~n38856;
  assign n38858 = ~i_StoB_REQ12 & ~n38857;
  assign n38859 = ~i_StoB_REQ12 & ~n38858;
  assign n38860 = controllable_BtoS_ACK12 & ~n38859;
  assign n38861 = i_StoB_REQ12 & ~n9269;
  assign n38862 = ~n38858 & ~n38861;
  assign n38863 = ~controllable_BtoS_ACK12 & ~n38862;
  assign n38864 = ~n38860 & ~n38863;
  assign n38865 = ~i_StoB_REQ13 & ~n38864;
  assign n38866 = ~n38781 & ~n38865;
  assign n38867 = n4466 & ~n38866;
  assign n38868 = ~n37027 & ~n38867;
  assign n38869 = ~i_StoB_REQ0 & ~n38868;
  assign n38870 = ~i_StoB_REQ0 & ~n38869;
  assign n38871 = ~i_StoB_REQ14 & ~n38870;
  assign n38872 = ~i_StoB_REQ14 & ~n38871;
  assign n38873 = controllable_BtoS_ACK14 & ~n38872;
  assign n38874 = ~n10454 & ~n38871;
  assign n38875 = ~controllable_BtoS_ACK14 & ~n38874;
  assign n38876 = ~n38873 & ~n38875;
  assign n38877 = ~controllable_ENQ & ~n38876;
  assign n38878 = ~n37246 & ~n38877;
  assign n38879 = i_RtoB_ACK1 & ~n38878;
  assign n38880 = ~n11660 & ~n38879;
  assign n38881 = controllable_BtoR_REQ1 & ~n38880;
  assign n38882 = ~n11668 & ~n38881;
  assign n38883 = ~controllable_BtoR_REQ0 & ~n38882;
  assign n38884 = ~controllable_BtoR_REQ0 & ~n38883;
  assign n38885 = ~i_RtoB_ACK0 & ~n38884;
  assign n38886 = ~n11654 & ~n38885;
  assign n38887 = controllable_DEQ & ~n38886;
  assign n38888 = i_RtoB_ACK1 & ~n37455;
  assign n38889 = ~n11429 & ~n38888;
  assign n38890 = controllable_BtoR_REQ1 & ~n38889;
  assign n38891 = ~n11686 & ~n38890;
  assign n38892 = ~controllable_BtoR_REQ0 & ~n38891;
  assign n38893 = ~controllable_BtoR_REQ0 & ~n38892;
  assign n38894 = ~i_RtoB_ACK0 & ~n38893;
  assign n38895 = ~n11683 & ~n38894;
  assign n38896 = ~controllable_DEQ & ~n38895;
  assign n38897 = ~n38887 & ~n38896;
  assign n38898 = i_FULL & ~n38897;
  assign n38899 = ~n11698 & ~n38879;
  assign n38900 = controllable_BtoR_REQ1 & ~n38899;
  assign n38901 = ~n11703 & ~n38900;
  assign n38902 = ~controllable_BtoR_REQ0 & ~n38901;
  assign n38903 = ~controllable_BtoR_REQ0 & ~n38902;
  assign n38904 = ~i_RtoB_ACK0 & ~n38903;
  assign n38905 = ~n11654 & ~n38904;
  assign n38906 = controllable_DEQ & ~n38905;
  assign n38907 = ~n11666 & ~n38888;
  assign n38908 = controllable_BtoR_REQ1 & ~n38907;
  assign n38909 = ~n11712 & ~n38908;
  assign n38910 = ~controllable_BtoR_REQ0 & ~n38909;
  assign n38911 = ~controllable_BtoR_REQ0 & ~n38910;
  assign n38912 = ~i_RtoB_ACK0 & ~n38911;
  assign n38913 = ~n11683 & ~n38912;
  assign n38914 = ~controllable_DEQ & ~n38913;
  assign n38915 = ~n38906 & ~n38914;
  assign n38916 = ~i_FULL & ~n38915;
  assign n38917 = ~n38898 & ~n38916;
  assign n38918 = i_nEMPTY & ~n38917;
  assign n38919 = ~controllable_ENQ & ~n38877;
  assign n38920 = i_RtoB_ACK1 & ~n38919;
  assign n38921 = ~n11726 & ~n38920;
  assign n38922 = controllable_BtoR_REQ1 & ~n38921;
  assign n38923 = ~n11732 & ~n38922;
  assign n38924 = ~controllable_BtoR_REQ0 & ~n38923;
  assign n38925 = ~controllable_BtoR_REQ0 & ~n38924;
  assign n38926 = ~i_RtoB_ACK0 & ~n38925;
  assign n38927 = ~i_RtoB_ACK0 & ~n38926;
  assign n38928 = controllable_DEQ & ~n38927;
  assign n38929 = i_RtoB_ACK1 & ~n37517;
  assign n38930 = ~n11479 & ~n38929;
  assign n38931 = controllable_BtoR_REQ1 & ~n38930;
  assign n38932 = ~n11740 & ~n38931;
  assign n38933 = ~controllable_BtoR_REQ0 & ~n38932;
  assign n38934 = ~controllable_BtoR_REQ0 & ~n38933;
  assign n38935 = ~i_RtoB_ACK0 & ~n38934;
  assign n38936 = ~n11654 & ~n38935;
  assign n38937 = ~controllable_DEQ & ~n38936;
  assign n38938 = ~n38928 & ~n38937;
  assign n38939 = i_FULL & ~n38938;
  assign n38940 = i_RtoB_ACK1 & ~n38876;
  assign n38941 = ~n11676 & ~n38940;
  assign n38942 = controllable_BtoR_REQ1 & ~n38941;
  assign n38943 = ~n11750 & ~n38942;
  assign n38944 = ~controllable_BtoR_REQ0 & ~n38943;
  assign n38945 = ~controllable_BtoR_REQ0 & ~n38944;
  assign n38946 = ~i_RtoB_ACK0 & ~n38945;
  assign n38947 = ~i_RtoB_ACK0 & ~n38946;
  assign n38948 = controllable_DEQ & ~n38947;
  assign n38949 = ~n11655 & ~n37516;
  assign n38950 = i_RtoB_ACK1 & ~n38949;
  assign n38951 = ~n11660 & ~n38950;
  assign n38952 = controllable_BtoR_REQ1 & ~n38951;
  assign n38953 = ~n11758 & ~n38952;
  assign n38954 = ~controllable_BtoR_REQ0 & ~n38953;
  assign n38955 = ~controllable_BtoR_REQ0 & ~n38954;
  assign n38956 = ~i_RtoB_ACK0 & ~n38955;
  assign n38957 = ~n11654 & ~n38956;
  assign n38958 = ~controllable_DEQ & ~n38957;
  assign n38959 = ~n38948 & ~n38958;
  assign n38960 = ~i_FULL & ~n38959;
  assign n38961 = ~n38939 & ~n38960;
  assign n38962 = ~i_nEMPTY & ~n38961;
  assign n38963 = ~n38918 & ~n38962;
  assign n38964 = controllable_BtoS_ACK0 & ~n38963;
  assign n38965 = ~n9771 & ~n38869;
  assign n38966 = ~i_StoB_REQ14 & ~n38965;
  assign n38967 = ~i_StoB_REQ14 & ~n38966;
  assign n38968 = controllable_BtoS_ACK14 & ~n38967;
  assign n38969 = ~n10584 & ~n38966;
  assign n38970 = ~controllable_BtoS_ACK14 & ~n38969;
  assign n38971 = ~n38968 & ~n38970;
  assign n38972 = ~controllable_ENQ & ~n38971;
  assign n38973 = ~n37688 & ~n38972;
  assign n38974 = i_RtoB_ACK1 & ~n38973;
  assign n38975 = ~n11807 & ~n38974;
  assign n38976 = controllable_BtoR_REQ1 & ~n38975;
  assign n38977 = ~n11815 & ~n38976;
  assign n38978 = ~controllable_BtoR_REQ0 & ~n38977;
  assign n38979 = ~controllable_BtoR_REQ0 & ~n38978;
  assign n38980 = ~i_RtoB_ACK0 & ~n38979;
  assign n38981 = ~n11801 & ~n38980;
  assign n38982 = controllable_DEQ & ~n38981;
  assign n38983 = i_RtoB_ACK1 & ~n37718;
  assign n38984 = ~n7288 & ~n38983;
  assign n38985 = controllable_BtoR_REQ1 & ~n38984;
  assign n38986 = ~n11833 & ~n38985;
  assign n38987 = ~controllable_BtoR_REQ0 & ~n38986;
  assign n38988 = ~controllable_BtoR_REQ0 & ~n38987;
  assign n38989 = ~i_RtoB_ACK0 & ~n38988;
  assign n38990 = ~n11830 & ~n38989;
  assign n38991 = ~controllable_DEQ & ~n38990;
  assign n38992 = ~n38982 & ~n38991;
  assign n38993 = i_FULL & ~n38992;
  assign n38994 = ~n11845 & ~n38974;
  assign n38995 = controllable_BtoR_REQ1 & ~n38994;
  assign n38996 = ~n11850 & ~n38995;
  assign n38997 = ~controllable_BtoR_REQ0 & ~n38996;
  assign n38998 = ~controllable_BtoR_REQ0 & ~n38997;
  assign n38999 = ~i_RtoB_ACK0 & ~n38998;
  assign n39000 = ~n11801 & ~n38999;
  assign n39001 = controllable_DEQ & ~n39000;
  assign n39002 = ~n11813 & ~n38983;
  assign n39003 = controllable_BtoR_REQ1 & ~n39002;
  assign n39004 = ~n11859 & ~n39003;
  assign n39005 = ~controllable_BtoR_REQ0 & ~n39004;
  assign n39006 = ~controllable_BtoR_REQ0 & ~n39005;
  assign n39007 = ~i_RtoB_ACK0 & ~n39006;
  assign n39008 = ~n11830 & ~n39007;
  assign n39009 = ~controllable_DEQ & ~n39008;
  assign n39010 = ~n39001 & ~n39009;
  assign n39011 = ~i_FULL & ~n39010;
  assign n39012 = ~n38993 & ~n39011;
  assign n39013 = i_nEMPTY & ~n39012;
  assign n39014 = ~controllable_ENQ & ~n38972;
  assign n39015 = i_RtoB_ACK1 & ~n39014;
  assign n39016 = ~n11873 & ~n39015;
  assign n39017 = controllable_BtoR_REQ1 & ~n39016;
  assign n39018 = ~n11879 & ~n39017;
  assign n39019 = ~controllable_BtoR_REQ0 & ~n39018;
  assign n39020 = ~controllable_BtoR_REQ0 & ~n39019;
  assign n39021 = ~i_RtoB_ACK0 & ~n39020;
  assign n39022 = ~i_RtoB_ACK0 & ~n39021;
  assign n39023 = controllable_DEQ & ~n39022;
  assign n39024 = i_RtoB_ACK1 & ~n37780;
  assign n39025 = ~n7345 & ~n39024;
  assign n39026 = controllable_BtoR_REQ1 & ~n39025;
  assign n39027 = ~n11887 & ~n39026;
  assign n39028 = ~controllable_BtoR_REQ0 & ~n39027;
  assign n39029 = ~controllable_BtoR_REQ0 & ~n39028;
  assign n39030 = ~i_RtoB_ACK0 & ~n39029;
  assign n39031 = ~n11801 & ~n39030;
  assign n39032 = ~controllable_DEQ & ~n39031;
  assign n39033 = ~n39023 & ~n39032;
  assign n39034 = i_FULL & ~n39033;
  assign n39035 = i_RtoB_ACK1 & ~n38971;
  assign n39036 = ~n11823 & ~n39035;
  assign n39037 = controllable_BtoR_REQ1 & ~n39036;
  assign n39038 = ~n11897 & ~n39037;
  assign n39039 = ~controllable_BtoR_REQ0 & ~n39038;
  assign n39040 = ~controllable_BtoR_REQ0 & ~n39039;
  assign n39041 = ~i_RtoB_ACK0 & ~n39040;
  assign n39042 = ~i_RtoB_ACK0 & ~n39041;
  assign n39043 = controllable_DEQ & ~n39042;
  assign n39044 = ~n11802 & ~n37779;
  assign n39045 = i_RtoB_ACK1 & ~n39044;
  assign n39046 = ~n11807 & ~n39045;
  assign n39047 = controllable_BtoR_REQ1 & ~n39046;
  assign n39048 = ~n11905 & ~n39047;
  assign n39049 = ~controllable_BtoR_REQ0 & ~n39048;
  assign n39050 = ~controllable_BtoR_REQ0 & ~n39049;
  assign n39051 = ~i_RtoB_ACK0 & ~n39050;
  assign n39052 = ~n11801 & ~n39051;
  assign n39053 = ~controllable_DEQ & ~n39052;
  assign n39054 = ~n39043 & ~n39053;
  assign n39055 = ~i_FULL & ~n39054;
  assign n39056 = ~n39034 & ~n39055;
  assign n39057 = ~i_nEMPTY & ~n39056;
  assign n39058 = ~n39013 & ~n39057;
  assign n39059 = ~controllable_BtoS_ACK0 & ~n39058;
  assign n39060 = ~n38964 & ~n39059;
  assign n39061 = n4465 & ~n39060;
  assign n39062 = ~n7270 & ~n37850;
  assign n39063 = ~controllable_BtoR_REQ0 & ~n39062;
  assign n39064 = ~controllable_BtoR_REQ0 & ~n39063;
  assign n39065 = ~i_RtoB_ACK0 & ~n39064;
  assign n39066 = ~n7246 & ~n39065;
  assign n39067 = controllable_DEQ & ~n39066;
  assign n39068 = ~n13428 & ~n39067;
  assign n39069 = i_FULL & ~n39068;
  assign n39070 = ~n7307 & ~n37860;
  assign n39071 = ~controllable_BtoR_REQ0 & ~n39070;
  assign n39072 = ~controllable_BtoR_REQ0 & ~n39071;
  assign n39073 = ~i_RtoB_ACK0 & ~n39072;
  assign n39074 = ~n7246 & ~n39073;
  assign n39075 = controllable_DEQ & ~n39074;
  assign n39076 = ~n13442 & ~n39075;
  assign n39077 = ~i_FULL & ~n39076;
  assign n39078 = ~n39069 & ~n39077;
  assign n39079 = i_nEMPTY & ~n39078;
  assign n39080 = ~n7336 & ~n37872;
  assign n39081 = ~controllable_BtoR_REQ0 & ~n39080;
  assign n39082 = ~controllable_BtoR_REQ0 & ~n39081;
  assign n39083 = ~i_RtoB_ACK0 & ~n39082;
  assign n39084 = ~i_RtoB_ACK0 & ~n39083;
  assign n39085 = controllable_DEQ & ~n39084;
  assign n39086 = ~n13452 & ~n39085;
  assign n39087 = i_FULL & ~n39086;
  assign n39088 = ~n7357 & ~n37882;
  assign n39089 = ~controllable_BtoR_REQ0 & ~n39088;
  assign n39090 = ~controllable_BtoR_REQ0 & ~n39089;
  assign n39091 = ~i_RtoB_ACK0 & ~n39090;
  assign n39092 = ~i_RtoB_ACK0 & ~n39091;
  assign n39093 = controllable_DEQ & ~n39092;
  assign n39094 = ~n13460 & ~n39093;
  assign n39095 = ~i_FULL & ~n39094;
  assign n39096 = ~n39087 & ~n39095;
  assign n39097 = ~i_nEMPTY & ~n39096;
  assign n39098 = ~n39079 & ~n39097;
  assign n39099 = ~controllable_BtoS_ACK0 & ~n39098;
  assign n39100 = ~n13416 & ~n39099;
  assign n39101 = ~n4465 & ~n39100;
  assign n39102 = ~n39061 & ~n39101;
  assign n39103 = ~i_StoB_REQ10 & ~n39102;
  assign n39104 = ~n38778 & ~n39103;
  assign n39105 = controllable_BtoS_ACK10 & ~n39104;
  assign n39106 = ~n9302 & ~n12173;
  assign n39107 = i_RtoB_ACK1 & ~n39106;
  assign n39108 = ~n11666 & ~n39107;
  assign n39109 = controllable_BtoR_REQ1 & ~n39108;
  assign n39110 = ~n11668 & ~n39109;
  assign n39111 = ~controllable_BtoR_REQ0 & ~n39110;
  assign n39112 = ~controllable_BtoR_REQ0 & ~n39111;
  assign n39113 = ~i_RtoB_ACK0 & ~n39112;
  assign n39114 = ~n36644 & ~n39113;
  assign n39115 = controllable_DEQ & ~n39114;
  assign n39116 = ~n11686 & ~n37470;
  assign n39117 = ~controllable_BtoR_REQ0 & ~n39116;
  assign n39118 = ~controllable_BtoR_REQ0 & ~n39117;
  assign n39119 = ~i_RtoB_ACK0 & ~n39118;
  assign n39120 = ~n36662 & ~n39119;
  assign n39121 = ~controllable_DEQ & ~n39120;
  assign n39122 = ~n39115 & ~n39121;
  assign n39123 = i_FULL & ~n39122;
  assign n39124 = ~n11701 & ~n39107;
  assign n39125 = controllable_BtoR_REQ1 & ~n39124;
  assign n39126 = ~n11703 & ~n39125;
  assign n39127 = ~controllable_BtoR_REQ0 & ~n39126;
  assign n39128 = ~controllable_BtoR_REQ0 & ~n39127;
  assign n39129 = ~i_RtoB_ACK0 & ~n39128;
  assign n39130 = ~n36644 & ~n39129;
  assign n39131 = controllable_DEQ & ~n39130;
  assign n39132 = ~n11712 & ~n37488;
  assign n39133 = ~controllable_BtoR_REQ0 & ~n39132;
  assign n39134 = ~controllable_BtoR_REQ0 & ~n39133;
  assign n39135 = ~i_RtoB_ACK0 & ~n39134;
  assign n39136 = ~n36662 & ~n39135;
  assign n39137 = ~controllable_DEQ & ~n39136;
  assign n39138 = ~n39131 & ~n39137;
  assign n39139 = ~i_FULL & ~n39138;
  assign n39140 = ~n39123 & ~n39139;
  assign n39141 = i_nEMPTY & ~n39140;
  assign n39142 = i_RtoB_ACK1 & ~n12204;
  assign n39143 = ~n11730 & ~n39142;
  assign n39144 = controllable_BtoR_REQ1 & ~n39143;
  assign n39145 = ~n11732 & ~n39144;
  assign n39146 = ~controllable_BtoR_REQ0 & ~n39145;
  assign n39147 = ~controllable_BtoR_REQ0 & ~n39146;
  assign n39148 = ~i_RtoB_ACK0 & ~n39147;
  assign n39149 = ~i_RtoB_ACK0 & ~n39148;
  assign n39150 = controllable_DEQ & ~n39149;
  assign n39151 = ~n11740 & ~n37529;
  assign n39152 = ~controllable_BtoR_REQ0 & ~n39151;
  assign n39153 = ~controllable_BtoR_REQ0 & ~n39152;
  assign n39154 = ~i_RtoB_ACK0 & ~n39153;
  assign n39155 = ~n36644 & ~n39154;
  assign n39156 = ~controllable_DEQ & ~n39155;
  assign n39157 = ~n39150 & ~n39156;
  assign n39158 = i_FULL & ~n39157;
  assign n39159 = ~n11701 & ~n14082;
  assign n39160 = controllable_BtoR_REQ1 & ~n39159;
  assign n39161 = ~n11750 & ~n39160;
  assign n39162 = ~controllable_BtoR_REQ0 & ~n39161;
  assign n39163 = ~controllable_BtoR_REQ0 & ~n39162;
  assign n39164 = ~i_RtoB_ACK0 & ~n39163;
  assign n39165 = ~i_RtoB_ACK0 & ~n39164;
  assign n39166 = controllable_DEQ & ~n39165;
  assign n39167 = ~n11668 & ~n37970;
  assign n39168 = ~controllable_BtoR_REQ0 & ~n39167;
  assign n39169 = ~controllable_BtoR_REQ0 & ~n39168;
  assign n39170 = ~i_RtoB_ACK0 & ~n39169;
  assign n39171 = ~n36644 & ~n39170;
  assign n39172 = ~controllable_DEQ & ~n39171;
  assign n39173 = ~n39166 & ~n39172;
  assign n39174 = ~i_FULL & ~n39173;
  assign n39175 = ~n39158 & ~n39174;
  assign n39176 = ~i_nEMPTY & ~n39175;
  assign n39177 = ~n39141 & ~n39176;
  assign n39178 = controllable_BtoS_ACK0 & ~n39177;
  assign n39179 = ~n9635 & ~n12264;
  assign n39180 = i_RtoB_ACK1 & ~n39179;
  assign n39181 = ~n11813 & ~n39180;
  assign n39182 = controllable_BtoR_REQ1 & ~n39181;
  assign n39183 = ~n11815 & ~n39182;
  assign n39184 = ~controllable_BtoR_REQ0 & ~n39183;
  assign n39185 = ~controllable_BtoR_REQ0 & ~n39184;
  assign n39186 = ~i_RtoB_ACK0 & ~n39185;
  assign n39187 = ~n36723 & ~n39186;
  assign n39188 = controllable_DEQ & ~n39187;
  assign n39189 = ~n11833 & ~n37733;
  assign n39190 = ~controllable_BtoR_REQ0 & ~n39189;
  assign n39191 = ~controllable_BtoR_REQ0 & ~n39190;
  assign n39192 = ~i_RtoB_ACK0 & ~n39191;
  assign n39193 = ~n36741 & ~n39192;
  assign n39194 = ~controllable_DEQ & ~n39193;
  assign n39195 = ~n39188 & ~n39194;
  assign n39196 = i_FULL & ~n39195;
  assign n39197 = ~n11848 & ~n39180;
  assign n39198 = controllable_BtoR_REQ1 & ~n39197;
  assign n39199 = ~n11850 & ~n39198;
  assign n39200 = ~controllable_BtoR_REQ0 & ~n39199;
  assign n39201 = ~controllable_BtoR_REQ0 & ~n39200;
  assign n39202 = ~i_RtoB_ACK0 & ~n39201;
  assign n39203 = ~n36723 & ~n39202;
  assign n39204 = controllable_DEQ & ~n39203;
  assign n39205 = ~n11859 & ~n37751;
  assign n39206 = ~controllable_BtoR_REQ0 & ~n39205;
  assign n39207 = ~controllable_BtoR_REQ0 & ~n39206;
  assign n39208 = ~i_RtoB_ACK0 & ~n39207;
  assign n39209 = ~n36741 & ~n39208;
  assign n39210 = ~controllable_DEQ & ~n39209;
  assign n39211 = ~n39204 & ~n39210;
  assign n39212 = ~i_FULL & ~n39211;
  assign n39213 = ~n39196 & ~n39212;
  assign n39214 = i_nEMPTY & ~n39213;
  assign n39215 = i_RtoB_ACK1 & ~n12290;
  assign n39216 = ~n11877 & ~n39215;
  assign n39217 = controllable_BtoR_REQ1 & ~n39216;
  assign n39218 = ~n11879 & ~n39217;
  assign n39219 = ~controllable_BtoR_REQ0 & ~n39218;
  assign n39220 = ~controllable_BtoR_REQ0 & ~n39219;
  assign n39221 = ~i_RtoB_ACK0 & ~n39220;
  assign n39222 = ~i_RtoB_ACK0 & ~n39221;
  assign n39223 = controllable_DEQ & ~n39222;
  assign n39224 = ~n11887 & ~n37792;
  assign n39225 = ~controllable_BtoR_REQ0 & ~n39224;
  assign n39226 = ~controllable_BtoR_REQ0 & ~n39225;
  assign n39227 = ~i_RtoB_ACK0 & ~n39226;
  assign n39228 = ~n36723 & ~n39227;
  assign n39229 = ~controllable_DEQ & ~n39228;
  assign n39230 = ~n39223 & ~n39229;
  assign n39231 = i_FULL & ~n39230;
  assign n39232 = ~n11848 & ~n14125;
  assign n39233 = controllable_BtoR_REQ1 & ~n39232;
  assign n39234 = ~n11897 & ~n39233;
  assign n39235 = ~controllable_BtoR_REQ0 & ~n39234;
  assign n39236 = ~controllable_BtoR_REQ0 & ~n39235;
  assign n39237 = ~i_RtoB_ACK0 & ~n39236;
  assign n39238 = ~i_RtoB_ACK0 & ~n39237;
  assign n39239 = controllable_DEQ & ~n39238;
  assign n39240 = ~n11815 & ~n38054;
  assign n39241 = ~controllable_BtoR_REQ0 & ~n39240;
  assign n39242 = ~controllable_BtoR_REQ0 & ~n39241;
  assign n39243 = ~i_RtoB_ACK0 & ~n39242;
  assign n39244 = ~n36723 & ~n39243;
  assign n39245 = ~controllable_DEQ & ~n39244;
  assign n39246 = ~n39239 & ~n39245;
  assign n39247 = ~i_FULL & ~n39246;
  assign n39248 = ~n39231 & ~n39247;
  assign n39249 = ~i_nEMPTY & ~n39248;
  assign n39250 = ~n39214 & ~n39249;
  assign n39251 = ~controllable_BtoS_ACK0 & ~n39250;
  assign n39252 = ~n39178 & ~n39251;
  assign n39253 = n4465 & ~n39252;
  assign n39254 = ~n7270 & ~n38078;
  assign n39255 = ~controllable_BtoR_REQ0 & ~n39254;
  assign n39256 = ~controllable_BtoR_REQ0 & ~n39255;
  assign n39257 = ~i_RtoB_ACK0 & ~n39256;
  assign n39258 = ~n7614 & ~n39257;
  assign n39259 = controllable_DEQ & ~n39258;
  assign n39260 = ~n13601 & ~n39259;
  assign n39261 = i_FULL & ~n39260;
  assign n39262 = ~n7307 & ~n38088;
  assign n39263 = ~controllable_BtoR_REQ0 & ~n39262;
  assign n39264 = ~controllable_BtoR_REQ0 & ~n39263;
  assign n39265 = ~i_RtoB_ACK0 & ~n39264;
  assign n39266 = ~n7614 & ~n39265;
  assign n39267 = controllable_DEQ & ~n39266;
  assign n39268 = ~n13611 & ~n39267;
  assign n39269 = ~i_FULL & ~n39268;
  assign n39270 = ~n39261 & ~n39269;
  assign n39271 = i_nEMPTY & ~n39270;
  assign n39272 = ~n7336 & ~n38100;
  assign n39273 = ~controllable_BtoR_REQ0 & ~n39272;
  assign n39274 = ~controllable_BtoR_REQ0 & ~n39273;
  assign n39275 = ~i_RtoB_ACK0 & ~n39274;
  assign n39276 = ~i_RtoB_ACK0 & ~n39275;
  assign n39277 = controllable_DEQ & ~n39276;
  assign n39278 = ~n13617 & ~n39277;
  assign n39279 = i_FULL & ~n39278;
  assign n39280 = ~n7357 & ~n38110;
  assign n39281 = ~controllable_BtoR_REQ0 & ~n39280;
  assign n39282 = ~controllable_BtoR_REQ0 & ~n39281;
  assign n39283 = ~i_RtoB_ACK0 & ~n39282;
  assign n39284 = ~i_RtoB_ACK0 & ~n39283;
  assign n39285 = controllable_DEQ & ~n39284;
  assign n39286 = ~n13620 & ~n39285;
  assign n39287 = ~i_FULL & ~n39286;
  assign n39288 = ~n39279 & ~n39287;
  assign n39289 = ~i_nEMPTY & ~n39288;
  assign n39290 = ~n39271 & ~n39289;
  assign n39291 = ~controllable_BtoS_ACK0 & ~n39290;
  assign n39292 = ~n13593 & ~n39291;
  assign n39293 = ~n4465 & ~n39292;
  assign n39294 = ~n39253 & ~n39293;
  assign n39295 = i_StoB_REQ10 & ~n39294;
  assign n39296 = ~n39103 & ~n39295;
  assign n39297 = ~controllable_BtoS_ACK10 & ~n39296;
  assign n39298 = ~n39105 & ~n39297;
  assign n39299 = n4464 & ~n39298;
  assign n39300 = ~n5238 & ~n10458;
  assign n39301 = i_RtoB_ACK1 & ~n39300;
  assign n39302 = ~n7932 & ~n39301;
  assign n39303 = controllable_BtoR_REQ1 & ~n39302;
  assign n39304 = ~n7940 & ~n39303;
  assign n39305 = ~controllable_BtoR_REQ0 & ~n39304;
  assign n39306 = ~controllable_BtoR_REQ0 & ~n39305;
  assign n39307 = ~i_RtoB_ACK0 & ~n39306;
  assign n39308 = ~n7921 & ~n39307;
  assign n39309 = controllable_DEQ & ~n39308;
  assign n39310 = ~n13713 & ~n39309;
  assign n39311 = i_FULL & ~n39310;
  assign n39312 = ~n7972 & ~n39301;
  assign n39313 = controllable_BtoR_REQ1 & ~n39312;
  assign n39314 = ~n7977 & ~n39313;
  assign n39315 = ~controllable_BtoR_REQ0 & ~n39314;
  assign n39316 = ~controllable_BtoR_REQ0 & ~n39315;
  assign n39317 = ~i_RtoB_ACK0 & ~n39316;
  assign n39318 = ~n7921 & ~n39317;
  assign n39319 = controllable_DEQ & ~n39318;
  assign n39320 = ~n13731 & ~n39319;
  assign n39321 = ~i_FULL & ~n39320;
  assign n39322 = ~n39311 & ~n39321;
  assign n39323 = i_nEMPTY & ~n39322;
  assign n39324 = ~n8006 & ~n38178;
  assign n39325 = ~controllable_BtoR_REQ0 & ~n39324;
  assign n39326 = ~controllable_BtoR_REQ0 & ~n39325;
  assign n39327 = ~i_RtoB_ACK0 & ~n39326;
  assign n39328 = ~i_RtoB_ACK0 & ~n39327;
  assign n39329 = controllable_DEQ & ~n39328;
  assign n39330 = ~n13744 & ~n39329;
  assign n39331 = i_FULL & ~n39330;
  assign n39332 = ~n8027 & ~n38188;
  assign n39333 = ~controllable_BtoR_REQ0 & ~n39332;
  assign n39334 = ~controllable_BtoR_REQ0 & ~n39333;
  assign n39335 = ~i_RtoB_ACK0 & ~n39334;
  assign n39336 = ~i_RtoB_ACK0 & ~n39335;
  assign n39337 = controllable_DEQ & ~n39336;
  assign n39338 = ~n13752 & ~n39337;
  assign n39339 = ~i_FULL & ~n39338;
  assign n39340 = ~n39331 & ~n39339;
  assign n39341 = ~i_nEMPTY & ~n39340;
  assign n39342 = ~n39323 & ~n39341;
  assign n39343 = controllable_BtoS_ACK0 & ~n39342;
  assign n39344 = ~n8946 & ~n10588;
  assign n39345 = i_RtoB_ACK1 & ~n39344;
  assign n39346 = ~n8096 & ~n39345;
  assign n39347 = controllable_BtoR_REQ1 & ~n39346;
  assign n39348 = ~n8104 & ~n39347;
  assign n39349 = ~controllable_BtoR_REQ0 & ~n39348;
  assign n39350 = ~controllable_BtoR_REQ0 & ~n39349;
  assign n39351 = ~i_RtoB_ACK0 & ~n39350;
  assign n39352 = ~n8088 & ~n39351;
  assign n39353 = controllable_DEQ & ~n39352;
  assign n39354 = ~n13777 & ~n39353;
  assign n39355 = i_FULL & ~n39354;
  assign n39356 = ~n8136 & ~n39345;
  assign n39357 = controllable_BtoR_REQ1 & ~n39356;
  assign n39358 = ~n8141 & ~n39357;
  assign n39359 = ~controllable_BtoR_REQ0 & ~n39358;
  assign n39360 = ~controllable_BtoR_REQ0 & ~n39359;
  assign n39361 = ~i_RtoB_ACK0 & ~n39360;
  assign n39362 = ~n8088 & ~n39361;
  assign n39363 = controllable_DEQ & ~n39362;
  assign n39364 = ~n13795 & ~n39363;
  assign n39365 = ~i_FULL & ~n39364;
  assign n39366 = ~n39355 & ~n39365;
  assign n39367 = i_nEMPTY & ~n39366;
  assign n39368 = ~n8170 & ~n38230;
  assign n39369 = ~controllable_BtoR_REQ0 & ~n39368;
  assign n39370 = ~controllable_BtoR_REQ0 & ~n39369;
  assign n39371 = ~i_RtoB_ACK0 & ~n39370;
  assign n39372 = ~i_RtoB_ACK0 & ~n39371;
  assign n39373 = controllable_DEQ & ~n39372;
  assign n39374 = ~n13808 & ~n39373;
  assign n39375 = i_FULL & ~n39374;
  assign n39376 = ~n8191 & ~n38240;
  assign n39377 = ~controllable_BtoR_REQ0 & ~n39376;
  assign n39378 = ~controllable_BtoR_REQ0 & ~n39377;
  assign n39379 = ~i_RtoB_ACK0 & ~n39378;
  assign n39380 = ~i_RtoB_ACK0 & ~n39379;
  assign n39381 = controllable_DEQ & ~n39380;
  assign n39382 = ~n13816 & ~n39381;
  assign n39383 = ~i_FULL & ~n39382;
  assign n39384 = ~n39375 & ~n39383;
  assign n39385 = ~i_nEMPTY & ~n39384;
  assign n39386 = ~n39367 & ~n39385;
  assign n39387 = ~controllable_BtoS_ACK0 & ~n39386;
  assign n39388 = ~n39343 & ~n39387;
  assign n39389 = n4465 & ~n39388;
  assign n39390 = ~n8345 & ~n38262;
  assign n39391 = ~controllable_BtoR_REQ0 & ~n39390;
  assign n39392 = ~controllable_BtoR_REQ0 & ~n39391;
  assign n39393 = ~i_RtoB_ACK0 & ~n39392;
  assign n39394 = ~n8331 & ~n39393;
  assign n39395 = controllable_DEQ & ~n39394;
  assign n39396 = ~n13870 & ~n39395;
  assign n39397 = i_FULL & ~n39396;
  assign n39398 = ~n8380 & ~n38272;
  assign n39399 = ~controllable_BtoR_REQ0 & ~n39398;
  assign n39400 = ~controllable_BtoR_REQ0 & ~n39399;
  assign n39401 = ~i_RtoB_ACK0 & ~n39400;
  assign n39402 = ~n8331 & ~n39401;
  assign n39403 = controllable_DEQ & ~n39402;
  assign n39404 = ~n13884 & ~n39403;
  assign n39405 = ~i_FULL & ~n39404;
  assign n39406 = ~n39397 & ~n39405;
  assign n39407 = i_nEMPTY & ~n39406;
  assign n39408 = ~n8409 & ~n38284;
  assign n39409 = ~controllable_BtoR_REQ0 & ~n39408;
  assign n39410 = ~controllable_BtoR_REQ0 & ~n39409;
  assign n39411 = ~i_RtoB_ACK0 & ~n39410;
  assign n39412 = ~i_RtoB_ACK0 & ~n39411;
  assign n39413 = controllable_DEQ & ~n39412;
  assign n39414 = ~n13894 & ~n39413;
  assign n39415 = i_FULL & ~n39414;
  assign n39416 = ~n8427 & ~n38294;
  assign n39417 = ~controllable_BtoR_REQ0 & ~n39416;
  assign n39418 = ~controllable_BtoR_REQ0 & ~n39417;
  assign n39419 = ~i_RtoB_ACK0 & ~n39418;
  assign n39420 = ~i_RtoB_ACK0 & ~n39419;
  assign n39421 = controllable_DEQ & ~n39420;
  assign n39422 = ~n13902 & ~n39421;
  assign n39423 = ~i_FULL & ~n39422;
  assign n39424 = ~n39415 & ~n39423;
  assign n39425 = ~i_nEMPTY & ~n39424;
  assign n39426 = ~n39407 & ~n39425;
  assign n39427 = ~controllable_BtoS_ACK0 & ~n39426;
  assign n39428 = ~n13858 & ~n39427;
  assign n39429 = ~n4465 & ~n39428;
  assign n39430 = ~n39389 & ~n39429;
  assign n39431 = ~i_StoB_REQ10 & ~n39430;
  assign n39432 = ~n13694 & ~n39431;
  assign n39433 = controllable_BtoS_ACK10 & ~n39432;
  assign n39434 = ~n7940 & ~n38320;
  assign n39435 = ~controllable_BtoR_REQ0 & ~n39434;
  assign n39436 = ~controllable_BtoR_REQ0 & ~n39435;
  assign n39437 = ~i_RtoB_ACK0 & ~n39436;
  assign n39438 = ~n8468 & ~n39437;
  assign n39439 = controllable_DEQ & ~n39438;
  assign n39440 = ~n13926 & ~n39439;
  assign n39441 = i_FULL & ~n39440;
  assign n39442 = ~n7977 & ~n38330;
  assign n39443 = ~controllable_BtoR_REQ0 & ~n39442;
  assign n39444 = ~controllable_BtoR_REQ0 & ~n39443;
  assign n39445 = ~i_RtoB_ACK0 & ~n39444;
  assign n39446 = ~n8468 & ~n39445;
  assign n39447 = controllable_DEQ & ~n39446;
  assign n39448 = ~n13940 & ~n39447;
  assign n39449 = ~i_FULL & ~n39448;
  assign n39450 = ~n39441 & ~n39449;
  assign n39451 = i_nEMPTY & ~n39450;
  assign n39452 = ~n8006 & ~n38342;
  assign n39453 = ~controllable_BtoR_REQ0 & ~n39452;
  assign n39454 = ~controllable_BtoR_REQ0 & ~n39453;
  assign n39455 = ~i_RtoB_ACK0 & ~n39454;
  assign n39456 = ~i_RtoB_ACK0 & ~n39455;
  assign n39457 = controllable_DEQ & ~n39456;
  assign n39458 = ~n13950 & ~n39457;
  assign n39459 = i_FULL & ~n39458;
  assign n39460 = ~n8027 & ~n38352;
  assign n39461 = ~controllable_BtoR_REQ0 & ~n39460;
  assign n39462 = ~controllable_BtoR_REQ0 & ~n39461;
  assign n39463 = ~i_RtoB_ACK0 & ~n39462;
  assign n39464 = ~i_RtoB_ACK0 & ~n39463;
  assign n39465 = controllable_DEQ & ~n39464;
  assign n39466 = ~n13953 & ~n39465;
  assign n39467 = ~i_FULL & ~n39466;
  assign n39468 = ~n39459 & ~n39467;
  assign n39469 = ~i_nEMPTY & ~n39468;
  assign n39470 = ~n39451 & ~n39469;
  assign n39471 = controllable_BtoS_ACK0 & ~n39470;
  assign n39472 = ~n8104 & ~n38372;
  assign n39473 = ~controllable_BtoR_REQ0 & ~n39472;
  assign n39474 = ~controllable_BtoR_REQ0 & ~n39473;
  assign n39475 = ~i_RtoB_ACK0 & ~n39474;
  assign n39476 = ~n8547 & ~n39475;
  assign n39477 = controllable_DEQ & ~n39476;
  assign n39478 = ~n13971 & ~n39477;
  assign n39479 = i_FULL & ~n39478;
  assign n39480 = ~n8141 & ~n38382;
  assign n39481 = ~controllable_BtoR_REQ0 & ~n39480;
  assign n39482 = ~controllable_BtoR_REQ0 & ~n39481;
  assign n39483 = ~i_RtoB_ACK0 & ~n39482;
  assign n39484 = ~n8547 & ~n39483;
  assign n39485 = controllable_DEQ & ~n39484;
  assign n39486 = ~n13985 & ~n39485;
  assign n39487 = ~i_FULL & ~n39486;
  assign n39488 = ~n39479 & ~n39487;
  assign n39489 = i_nEMPTY & ~n39488;
  assign n39490 = ~n8170 & ~n38394;
  assign n39491 = ~controllable_BtoR_REQ0 & ~n39490;
  assign n39492 = ~controllable_BtoR_REQ0 & ~n39491;
  assign n39493 = ~i_RtoB_ACK0 & ~n39492;
  assign n39494 = ~i_RtoB_ACK0 & ~n39493;
  assign n39495 = controllable_DEQ & ~n39494;
  assign n39496 = ~n13995 & ~n39495;
  assign n39497 = i_FULL & ~n39496;
  assign n39498 = ~n8191 & ~n38404;
  assign n39499 = ~controllable_BtoR_REQ0 & ~n39498;
  assign n39500 = ~controllable_BtoR_REQ0 & ~n39499;
  assign n39501 = ~i_RtoB_ACK0 & ~n39500;
  assign n39502 = ~i_RtoB_ACK0 & ~n39501;
  assign n39503 = controllable_DEQ & ~n39502;
  assign n39504 = ~n13998 & ~n39503;
  assign n39505 = ~i_FULL & ~n39504;
  assign n39506 = ~n39497 & ~n39505;
  assign n39507 = ~i_nEMPTY & ~n39506;
  assign n39508 = ~n39489 & ~n39507;
  assign n39509 = ~controllable_BtoS_ACK0 & ~n39508;
  assign n39510 = ~n39471 & ~n39509;
  assign n39511 = n4465 & ~n39510;
  assign n39512 = ~n8345 & ~n38426;
  assign n39513 = ~controllable_BtoR_REQ0 & ~n39512;
  assign n39514 = ~controllable_BtoR_REQ0 & ~n39513;
  assign n39515 = ~i_RtoB_ACK0 & ~n39514;
  assign n39516 = ~n8679 & ~n39515;
  assign n39517 = controllable_DEQ & ~n39516;
  assign n39518 = ~n14035 & ~n39517;
  assign n39519 = i_FULL & ~n39518;
  assign n39520 = ~n8380 & ~n38436;
  assign n39521 = ~controllable_BtoR_REQ0 & ~n39520;
  assign n39522 = ~controllable_BtoR_REQ0 & ~n39521;
  assign n39523 = ~i_RtoB_ACK0 & ~n39522;
  assign n39524 = ~n8679 & ~n39523;
  assign n39525 = controllable_DEQ & ~n39524;
  assign n39526 = ~n14045 & ~n39525;
  assign n39527 = ~i_FULL & ~n39526;
  assign n39528 = ~n39519 & ~n39527;
  assign n39529 = i_nEMPTY & ~n39528;
  assign n39530 = ~n8409 & ~n38448;
  assign n39531 = ~controllable_BtoR_REQ0 & ~n39530;
  assign n39532 = ~controllable_BtoR_REQ0 & ~n39531;
  assign n39533 = ~i_RtoB_ACK0 & ~n39532;
  assign n39534 = ~i_RtoB_ACK0 & ~n39533;
  assign n39535 = controllable_DEQ & ~n39534;
  assign n39536 = ~n14051 & ~n39535;
  assign n39537 = i_FULL & ~n39536;
  assign n39538 = ~n8427 & ~n38458;
  assign n39539 = ~controllable_BtoR_REQ0 & ~n39538;
  assign n39540 = ~controllable_BtoR_REQ0 & ~n39539;
  assign n39541 = ~i_RtoB_ACK0 & ~n39540;
  assign n39542 = ~i_RtoB_ACK0 & ~n39541;
  assign n39543 = controllable_DEQ & ~n39542;
  assign n39544 = ~n14054 & ~n39543;
  assign n39545 = ~i_FULL & ~n39544;
  assign n39546 = ~n39537 & ~n39545;
  assign n39547 = ~i_nEMPTY & ~n39546;
  assign n39548 = ~n39529 & ~n39547;
  assign n39549 = ~controllable_BtoS_ACK0 & ~n39548;
  assign n39550 = ~n14027 & ~n39549;
  assign n39551 = ~n4465 & ~n39550;
  assign n39552 = ~n39511 & ~n39551;
  assign n39553 = i_StoB_REQ10 & ~n39552;
  assign n39554 = ~n39431 & ~n39553;
  assign n39555 = ~controllable_BtoS_ACK10 & ~n39554;
  assign n39556 = ~n39433 & ~n39555;
  assign n39557 = ~n4464 & ~n39556;
  assign n39558 = ~n39299 & ~n39557;
  assign n39559 = n4463 & ~n39558;
  assign n39560 = ~n38480 & ~n39559;
  assign n39561 = n4462 & ~n39560;
  assign n39562 = ~n11668 & ~n37256;
  assign n39563 = ~controllable_BtoR_REQ0 & ~n39562;
  assign n39564 = ~controllable_BtoR_REQ0 & ~n39563;
  assign n39565 = ~i_RtoB_ACK0 & ~n39564;
  assign n39566 = ~n11654 & ~n39565;
  assign n39567 = controllable_DEQ & ~n39566;
  assign n39568 = ~n14271 & ~n39567;
  assign n39569 = i_FULL & ~n39568;
  assign n39570 = ~n11703 & ~n37480;
  assign n39571 = ~controllable_BtoR_REQ0 & ~n39570;
  assign n39572 = ~controllable_BtoR_REQ0 & ~n39571;
  assign n39573 = ~i_RtoB_ACK0 & ~n39572;
  assign n39574 = ~n11654 & ~n39573;
  assign n39575 = controllable_DEQ & ~n39574;
  assign n39576 = ~n14285 & ~n39575;
  assign n39577 = ~i_FULL & ~n39576;
  assign n39578 = ~n39569 & ~n39577;
  assign n39579 = i_nEMPTY & ~n39578;
  assign n39580 = ~n11732 & ~n37505;
  assign n39581 = ~controllable_BtoR_REQ0 & ~n39580;
  assign n39582 = ~controllable_BtoR_REQ0 & ~n39581;
  assign n39583 = ~i_RtoB_ACK0 & ~n39582;
  assign n39584 = ~i_RtoB_ACK0 & ~n39583;
  assign n39585 = controllable_DEQ & ~n39584;
  assign n39586 = ~n14295 & ~n39585;
  assign n39587 = i_FULL & ~n39586;
  assign n39588 = ~n11750 & ~n37539;
  assign n39589 = ~controllable_BtoR_REQ0 & ~n39588;
  assign n39590 = ~controllable_BtoR_REQ0 & ~n39589;
  assign n39591 = ~i_RtoB_ACK0 & ~n39590;
  assign n39592 = ~i_RtoB_ACK0 & ~n39591;
  assign n39593 = controllable_DEQ & ~n39592;
  assign n39594 = ~n14303 & ~n39593;
  assign n39595 = ~i_FULL & ~n39594;
  assign n39596 = ~n39587 & ~n39595;
  assign n39597 = ~i_nEMPTY & ~n39596;
  assign n39598 = ~n39579 & ~n39597;
  assign n39599 = controllable_BtoS_ACK0 & ~n39598;
  assign n39600 = ~n11815 & ~n37698;
  assign n39601 = ~controllable_BtoR_REQ0 & ~n39600;
  assign n39602 = ~controllable_BtoR_REQ0 & ~n39601;
  assign n39603 = ~i_RtoB_ACK0 & ~n39602;
  assign n39604 = ~n11801 & ~n39603;
  assign n39605 = controllable_DEQ & ~n39604;
  assign n39606 = ~n14321 & ~n39605;
  assign n39607 = i_FULL & ~n39606;
  assign n39608 = ~n11850 & ~n37743;
  assign n39609 = ~controllable_BtoR_REQ0 & ~n39608;
  assign n39610 = ~controllable_BtoR_REQ0 & ~n39609;
  assign n39611 = ~i_RtoB_ACK0 & ~n39610;
  assign n39612 = ~n11801 & ~n39611;
  assign n39613 = controllable_DEQ & ~n39612;
  assign n39614 = ~n14335 & ~n39613;
  assign n39615 = ~i_FULL & ~n39614;
  assign n39616 = ~n39607 & ~n39615;
  assign n39617 = i_nEMPTY & ~n39616;
  assign n39618 = ~n11879 & ~n37768;
  assign n39619 = ~controllable_BtoR_REQ0 & ~n39618;
  assign n39620 = ~controllable_BtoR_REQ0 & ~n39619;
  assign n39621 = ~i_RtoB_ACK0 & ~n39620;
  assign n39622 = ~i_RtoB_ACK0 & ~n39621;
  assign n39623 = controllable_DEQ & ~n39622;
  assign n39624 = ~n14345 & ~n39623;
  assign n39625 = i_FULL & ~n39624;
  assign n39626 = ~n11897 & ~n37802;
  assign n39627 = ~controllable_BtoR_REQ0 & ~n39626;
  assign n39628 = ~controllable_BtoR_REQ0 & ~n39627;
  assign n39629 = ~i_RtoB_ACK0 & ~n39628;
  assign n39630 = ~i_RtoB_ACK0 & ~n39629;
  assign n39631 = controllable_DEQ & ~n39630;
  assign n39632 = ~n14353 & ~n39631;
  assign n39633 = ~i_FULL & ~n39632;
  assign n39634 = ~n39625 & ~n39633;
  assign n39635 = ~i_nEMPTY & ~n39634;
  assign n39636 = ~n39617 & ~n39635;
  assign n39637 = ~controllable_BtoS_ACK0 & ~n39636;
  assign n39638 = ~n39599 & ~n39637;
  assign n39639 = n4465 & ~n39638;
  assign n39640 = ~n14387 & ~n39099;
  assign n39641 = ~n4465 & ~n39640;
  assign n39642 = ~n39639 & ~n39641;
  assign n39643 = ~i_StoB_REQ10 & ~n39642;
  assign n39644 = ~n14259 & ~n39643;
  assign n39645 = ~controllable_BtoS_ACK10 & ~n39644;
  assign n39646 = ~n14163 & ~n39645;
  assign n39647 = n4464 & ~n39646;
  assign n39648 = ~n7940 & ~n38156;
  assign n39649 = ~controllable_BtoR_REQ0 & ~n39648;
  assign n39650 = ~controllable_BtoR_REQ0 & ~n39649;
  assign n39651 = ~i_RtoB_ACK0 & ~n39650;
  assign n39652 = ~n7921 & ~n39651;
  assign n39653 = controllable_DEQ & ~n39652;
  assign n39654 = ~n14501 & ~n39653;
  assign n39655 = i_FULL & ~n39654;
  assign n39656 = ~n7977 & ~n38166;
  assign n39657 = ~controllable_BtoR_REQ0 & ~n39656;
  assign n39658 = ~controllable_BtoR_REQ0 & ~n39657;
  assign n39659 = ~i_RtoB_ACK0 & ~n39658;
  assign n39660 = ~n7921 & ~n39659;
  assign n39661 = controllable_DEQ & ~n39660;
  assign n39662 = ~n14511 & ~n39661;
  assign n39663 = ~i_FULL & ~n39662;
  assign n39664 = ~n39655 & ~n39663;
  assign n39665 = i_nEMPTY & ~n39664;
  assign n39666 = ~n14517 & ~n39329;
  assign n39667 = i_FULL & ~n39666;
  assign n39668 = ~n14525 & ~n39337;
  assign n39669 = ~i_FULL & ~n39668;
  assign n39670 = ~n39667 & ~n39669;
  assign n39671 = ~i_nEMPTY & ~n39670;
  assign n39672 = ~n39665 & ~n39671;
  assign n39673 = controllable_BtoS_ACK0 & ~n39672;
  assign n39674 = ~n8104 & ~n38208;
  assign n39675 = ~controllable_BtoR_REQ0 & ~n39674;
  assign n39676 = ~controllable_BtoR_REQ0 & ~n39675;
  assign n39677 = ~i_RtoB_ACK0 & ~n39676;
  assign n39678 = ~n8088 & ~n39677;
  assign n39679 = controllable_DEQ & ~n39678;
  assign n39680 = ~n14539 & ~n39679;
  assign n39681 = i_FULL & ~n39680;
  assign n39682 = ~n8141 & ~n38218;
  assign n39683 = ~controllable_BtoR_REQ0 & ~n39682;
  assign n39684 = ~controllable_BtoR_REQ0 & ~n39683;
  assign n39685 = ~i_RtoB_ACK0 & ~n39684;
  assign n39686 = ~n8088 & ~n39685;
  assign n39687 = controllable_DEQ & ~n39686;
  assign n39688 = ~n14549 & ~n39687;
  assign n39689 = ~i_FULL & ~n39688;
  assign n39690 = ~n39681 & ~n39689;
  assign n39691 = i_nEMPTY & ~n39690;
  assign n39692 = ~n14555 & ~n39373;
  assign n39693 = i_FULL & ~n39692;
  assign n39694 = ~n14563 & ~n39381;
  assign n39695 = ~i_FULL & ~n39694;
  assign n39696 = ~n39693 & ~n39695;
  assign n39697 = ~i_nEMPTY & ~n39696;
  assign n39698 = ~n39691 & ~n39697;
  assign n39699 = ~controllable_BtoS_ACK0 & ~n39698;
  assign n39700 = ~n39673 & ~n39699;
  assign n39701 = n4465 & ~n39700;
  assign n39702 = ~n39429 & ~n39701;
  assign n39703 = ~i_StoB_REQ10 & ~n39702;
  assign n39704 = ~n14493 & ~n39703;
  assign n39705 = ~controllable_BtoS_ACK10 & ~n39704;
  assign n39706 = ~n14397 & ~n39705;
  assign n39707 = ~n4464 & ~n39706;
  assign n39708 = ~n39647 & ~n39707;
  assign n39709 = n4463 & ~n39708;
  assign n39710 = ~n38730 & ~n39709;
  assign n39711 = ~n4462 & ~n39710;
  assign n39712 = ~n39561 & ~n39711;
  assign n39713 = ~n4461 & ~n39712;
  assign n39714 = ~n38734 & ~n39713;
  assign n39715 = ~n4459 & ~n39714;
  assign n39716 = ~n17611 & ~n18248;
  assign n39717 = controllable_BtoS_ACK10 & ~n39716;
  assign n39718 = ~i_RtoB_ACK1 & ~n36646;
  assign n39719 = ~n36637 & ~n39718;
  assign n39720 = ~controllable_BtoR_REQ1 & ~n39719;
  assign n39721 = ~controllable_BtoR_REQ1 & ~n39720;
  assign n39722 = controllable_BtoR_REQ0 & ~n39721;
  assign n39723 = ~n17967 & ~n39722;
  assign n39724 = i_RtoB_ACK0 & ~n39723;
  assign n39725 = ~i_RtoB_ACK0 & ~n17975;
  assign n39726 = ~n39724 & ~n39725;
  assign n39727 = controllable_DEQ & ~n39726;
  assign n39728 = ~n11429 & ~n36656;
  assign n39729 = ~controllable_BtoR_REQ1 & ~n39728;
  assign n39730 = ~controllable_BtoR_REQ1 & ~n39729;
  assign n39731 = controllable_BtoR_REQ0 & ~n39730;
  assign n39732 = ~n17986 & ~n39731;
  assign n39733 = i_RtoB_ACK0 & ~n39732;
  assign n39734 = ~i_RtoB_ACK0 & ~n17994;
  assign n39735 = ~n39733 & ~n39734;
  assign n39736 = ~controllable_DEQ & ~n39735;
  assign n39737 = ~n39727 & ~n39736;
  assign n39738 = i_FULL & ~n39737;
  assign n39739 = ~i_RtoB_ACK1 & ~n36667;
  assign n39740 = ~n36637 & ~n39739;
  assign n39741 = ~controllable_BtoR_REQ1 & ~n39740;
  assign n39742 = ~controllable_BtoR_REQ1 & ~n39741;
  assign n39743 = controllable_BtoR_REQ0 & ~n39742;
  assign n39744 = ~n17967 & ~n39743;
  assign n39745 = i_RtoB_ACK0 & ~n39744;
  assign n39746 = ~i_RtoB_ACK0 & ~n18013;
  assign n39747 = ~n39745 & ~n39746;
  assign n39748 = controllable_DEQ & ~n39747;
  assign n39749 = ~n11666 & ~n36656;
  assign n39750 = ~controllable_BtoR_REQ1 & ~n39749;
  assign n39751 = ~controllable_BtoR_REQ1 & ~n39750;
  assign n39752 = controllable_BtoR_REQ0 & ~n39751;
  assign n39753 = ~n17986 & ~n39752;
  assign n39754 = i_RtoB_ACK0 & ~n39753;
  assign n39755 = ~i_RtoB_ACK0 & ~n18029;
  assign n39756 = ~n39754 & ~n39755;
  assign n39757 = ~controllable_DEQ & ~n39756;
  assign n39758 = ~n39748 & ~n39757;
  assign n39759 = ~i_FULL & ~n39758;
  assign n39760 = ~n39738 & ~n39759;
  assign n39761 = i_nEMPTY & ~n39760;
  assign n39762 = ~i_RtoB_ACK1 & ~n36683;
  assign n39763 = ~i_RtoB_ACK1 & ~n39762;
  assign n39764 = ~controllable_BtoR_REQ1 & ~n39763;
  assign n39765 = ~controllable_BtoR_REQ1 & ~n39764;
  assign n39766 = controllable_BtoR_REQ0 & ~n39765;
  assign n39767 = controllable_BtoR_REQ0 & ~n39766;
  assign n39768 = i_RtoB_ACK0 & ~n39767;
  assign n39769 = ~i_RtoB_ACK0 & ~n18050;
  assign n39770 = ~n39768 & ~n39769;
  assign n39771 = controllable_DEQ & ~n39770;
  assign n39772 = ~n11479 & ~n36637;
  assign n39773 = ~controllable_BtoR_REQ1 & ~n39772;
  assign n39774 = ~controllable_BtoR_REQ1 & ~n39773;
  assign n39775 = controllable_BtoR_REQ0 & ~n39774;
  assign n39776 = ~n17967 & ~n39775;
  assign n39777 = i_RtoB_ACK0 & ~n39776;
  assign n39778 = ~i_RtoB_ACK0 & ~n18066;
  assign n39779 = ~n39777 & ~n39778;
  assign n39780 = ~controllable_DEQ & ~n39779;
  assign n39781 = ~n39771 & ~n39780;
  assign n39782 = i_FULL & ~n39781;
  assign n39783 = ~i_RtoB_ACK1 & ~n36634;
  assign n39784 = ~i_RtoB_ACK1 & ~n39783;
  assign n39785 = ~controllable_BtoR_REQ1 & ~n39784;
  assign n39786 = ~controllable_BtoR_REQ1 & ~n39785;
  assign n39787 = controllable_BtoR_REQ0 & ~n39786;
  assign n39788 = controllable_BtoR_REQ0 & ~n39787;
  assign n39789 = i_RtoB_ACK0 & ~n39788;
  assign n39790 = ~i_RtoB_ACK0 & ~n18085;
  assign n39791 = ~n39789 & ~n39790;
  assign n39792 = controllable_DEQ & ~n39791;
  assign n39793 = ~controllable_DEQ & ~n39726;
  assign n39794 = ~n39792 & ~n39793;
  assign n39795 = ~i_FULL & ~n39794;
  assign n39796 = ~n39782 & ~n39795;
  assign n39797 = ~i_nEMPTY & ~n39796;
  assign n39798 = ~n39761 & ~n39797;
  assign n39799 = controllable_BtoS_ACK0 & ~n39798;
  assign n39800 = ~i_RtoB_ACK1 & ~n36725;
  assign n39801 = ~n36716 & ~n39800;
  assign n39802 = ~controllable_BtoR_REQ1 & ~n39801;
  assign n39803 = ~controllable_BtoR_REQ1 & ~n39802;
  assign n39804 = controllable_BtoR_REQ0 & ~n39803;
  assign n39805 = ~n18109 & ~n39804;
  assign n39806 = i_RtoB_ACK0 & ~n39805;
  assign n39807 = ~i_RtoB_ACK0 & ~n18117;
  assign n39808 = ~n39806 & ~n39807;
  assign n39809 = controllable_DEQ & ~n39808;
  assign n39810 = ~n7288 & ~n36735;
  assign n39811 = ~controllable_BtoR_REQ1 & ~n39810;
  assign n39812 = ~controllable_BtoR_REQ1 & ~n39811;
  assign n39813 = controllable_BtoR_REQ0 & ~n39812;
  assign n39814 = ~n18128 & ~n39813;
  assign n39815 = i_RtoB_ACK0 & ~n39814;
  assign n39816 = ~i_RtoB_ACK0 & ~n18136;
  assign n39817 = ~n39815 & ~n39816;
  assign n39818 = ~controllable_DEQ & ~n39817;
  assign n39819 = ~n39809 & ~n39818;
  assign n39820 = i_FULL & ~n39819;
  assign n39821 = ~i_RtoB_ACK1 & ~n36746;
  assign n39822 = ~n36716 & ~n39821;
  assign n39823 = ~controllable_BtoR_REQ1 & ~n39822;
  assign n39824 = ~controllable_BtoR_REQ1 & ~n39823;
  assign n39825 = controllable_BtoR_REQ0 & ~n39824;
  assign n39826 = ~n18109 & ~n39825;
  assign n39827 = i_RtoB_ACK0 & ~n39826;
  assign n39828 = ~i_RtoB_ACK0 & ~n18155;
  assign n39829 = ~n39827 & ~n39828;
  assign n39830 = controllable_DEQ & ~n39829;
  assign n39831 = ~n11813 & ~n36735;
  assign n39832 = ~controllable_BtoR_REQ1 & ~n39831;
  assign n39833 = ~controllable_BtoR_REQ1 & ~n39832;
  assign n39834 = controllable_BtoR_REQ0 & ~n39833;
  assign n39835 = ~n18128 & ~n39834;
  assign n39836 = i_RtoB_ACK0 & ~n39835;
  assign n39837 = ~i_RtoB_ACK0 & ~n18171;
  assign n39838 = ~n39836 & ~n39837;
  assign n39839 = ~controllable_DEQ & ~n39838;
  assign n39840 = ~n39830 & ~n39839;
  assign n39841 = ~i_FULL & ~n39840;
  assign n39842 = ~n39820 & ~n39841;
  assign n39843 = i_nEMPTY & ~n39842;
  assign n39844 = ~i_RtoB_ACK1 & ~n36762;
  assign n39845 = ~i_RtoB_ACK1 & ~n39844;
  assign n39846 = ~controllable_BtoR_REQ1 & ~n39845;
  assign n39847 = ~controllable_BtoR_REQ1 & ~n39846;
  assign n39848 = controllable_BtoR_REQ0 & ~n39847;
  assign n39849 = controllable_BtoR_REQ0 & ~n39848;
  assign n39850 = i_RtoB_ACK0 & ~n39849;
  assign n39851 = ~i_RtoB_ACK0 & ~n18192;
  assign n39852 = ~n39850 & ~n39851;
  assign n39853 = controllable_DEQ & ~n39852;
  assign n39854 = ~n7345 & ~n36716;
  assign n39855 = ~controllable_BtoR_REQ1 & ~n39854;
  assign n39856 = ~controllable_BtoR_REQ1 & ~n39855;
  assign n39857 = controllable_BtoR_REQ0 & ~n39856;
  assign n39858 = ~n18109 & ~n39857;
  assign n39859 = i_RtoB_ACK0 & ~n39858;
  assign n39860 = ~i_RtoB_ACK0 & ~n18208;
  assign n39861 = ~n39859 & ~n39860;
  assign n39862 = ~controllable_DEQ & ~n39861;
  assign n39863 = ~n39853 & ~n39862;
  assign n39864 = i_FULL & ~n39863;
  assign n39865 = ~i_RtoB_ACK1 & ~n36713;
  assign n39866 = ~i_RtoB_ACK1 & ~n39865;
  assign n39867 = ~controllable_BtoR_REQ1 & ~n39866;
  assign n39868 = ~controllable_BtoR_REQ1 & ~n39867;
  assign n39869 = controllable_BtoR_REQ0 & ~n39868;
  assign n39870 = controllable_BtoR_REQ0 & ~n39869;
  assign n39871 = i_RtoB_ACK0 & ~n39870;
  assign n39872 = ~i_RtoB_ACK0 & ~n18227;
  assign n39873 = ~n39871 & ~n39872;
  assign n39874 = controllable_DEQ & ~n39873;
  assign n39875 = ~controllable_DEQ & ~n39808;
  assign n39876 = ~n39874 & ~n39875;
  assign n39877 = ~i_FULL & ~n39876;
  assign n39878 = ~n39864 & ~n39877;
  assign n39879 = ~i_nEMPTY & ~n39878;
  assign n39880 = ~n39843 & ~n39879;
  assign n39881 = ~controllable_BtoS_ACK0 & ~n39880;
  assign n39882 = ~n39799 & ~n39881;
  assign n39883 = n4465 & ~n39882;
  assign n39884 = ~n15713 & ~n39883;
  assign n39885 = i_StoB_REQ10 & ~n39884;
  assign n39886 = ~n18248 & ~n39885;
  assign n39887 = ~controllable_BtoS_ACK10 & ~n39886;
  assign n39888 = ~n39717 & ~n39887;
  assign n39889 = n4464 & ~n39888;
  assign n39890 = ~n16695 & ~n39889;
  assign n39891 = n4463 & ~n39890;
  assign n39892 = ~i_RtoB_ACK1 & ~n36879;
  assign n39893 = ~controllable_BtoR_REQ1 & ~n39892;
  assign n39894 = ~controllable_BtoR_REQ1 & ~n39893;
  assign n39895 = controllable_BtoR_REQ0 & ~n39894;
  assign n39896 = ~n17555 & ~n39895;
  assign n39897 = i_RtoB_ACK0 & ~n39896;
  assign n39898 = ~n17564 & ~n39897;
  assign n39899 = ~controllable_DEQ & ~n39898;
  assign n39900 = ~n18432 & ~n39899;
  assign n39901 = i_nEMPTY & ~n39900;
  assign n39902 = ~i_RtoB_ACK1 & ~n36914;
  assign n39903 = ~controllable_BtoR_REQ1 & ~n39902;
  assign n39904 = ~controllable_BtoR_REQ1 & ~n39903;
  assign n39905 = controllable_BtoR_REQ0 & ~n39904;
  assign n39906 = ~n17538 & ~n39905;
  assign n39907 = i_RtoB_ACK0 & ~n39906;
  assign n39908 = ~n17583 & ~n39907;
  assign n39909 = ~controllable_DEQ & ~n39908;
  assign n39910 = ~n17577 & ~n39909;
  assign n39911 = i_FULL & ~n39910;
  assign n39912 = ~n17599 & ~n39907;
  assign n39913 = ~controllable_DEQ & ~n39912;
  assign n39914 = ~n17595 & ~n39913;
  assign n39915 = ~i_FULL & ~n39914;
  assign n39916 = ~n39911 & ~n39915;
  assign n39917 = ~i_nEMPTY & ~n39916;
  assign n39918 = ~n39901 & ~n39917;
  assign n39919 = controllable_BtoS_ACK0 & ~n39918;
  assign n39920 = ~i_RtoB_ACK1 & ~n37060;
  assign n39921 = ~controllable_BtoR_REQ1 & ~n39920;
  assign n39922 = ~controllable_BtoR_REQ1 & ~n39921;
  assign n39923 = controllable_BtoR_REQ0 & ~n39922;
  assign n39924 = ~n14834 & ~n39923;
  assign n39925 = i_RtoB_ACK0 & ~n39924;
  assign n39926 = ~n14843 & ~n39925;
  assign n39927 = ~controllable_DEQ & ~n39926;
  assign n39928 = ~n18460 & ~n39927;
  assign n39929 = i_nEMPTY & ~n39928;
  assign n39930 = ~i_RtoB_ACK1 & ~n37095;
  assign n39931 = ~controllable_BtoR_REQ1 & ~n39930;
  assign n39932 = ~controllable_BtoR_REQ1 & ~n39931;
  assign n39933 = controllable_BtoR_REQ0 & ~n39932;
  assign n39934 = ~n14817 & ~n39933;
  assign n39935 = i_RtoB_ACK0 & ~n39934;
  assign n39936 = ~n14862 & ~n39935;
  assign n39937 = ~controllable_DEQ & ~n39936;
  assign n39938 = ~n14856 & ~n39937;
  assign n39939 = i_FULL & ~n39938;
  assign n39940 = ~n14878 & ~n39935;
  assign n39941 = ~controllable_DEQ & ~n39940;
  assign n39942 = ~n14874 & ~n39941;
  assign n39943 = ~i_FULL & ~n39942;
  assign n39944 = ~n39939 & ~n39943;
  assign n39945 = ~i_nEMPTY & ~n39944;
  assign n39946 = ~n39929 & ~n39945;
  assign n39947 = ~controllable_BtoS_ACK0 & ~n39946;
  assign n39948 = ~n39919 & ~n39947;
  assign n39949 = n4465 & ~n39948;
  assign n39950 = ~n16773 & ~n39949;
  assign n39951 = i_StoB_REQ10 & ~n39950;
  assign n39952 = ~i_RtoB_ACK1 & ~n38878;
  assign n39953 = ~n11632 & ~n39952;
  assign n39954 = ~controllable_BtoR_REQ1 & ~n39953;
  assign n39955 = ~controllable_BtoR_REQ1 & ~n39954;
  assign n39956 = controllable_BtoR_REQ0 & ~n39955;
  assign n39957 = ~n17967 & ~n39956;
  assign n39958 = i_RtoB_ACK0 & ~n39957;
  assign n39959 = ~n17978 & ~n39958;
  assign n39960 = controllable_DEQ & ~n39959;
  assign n39961 = ~n11675 & ~n37456;
  assign n39962 = ~controllable_BtoR_REQ1 & ~n39961;
  assign n39963 = ~controllable_BtoR_REQ1 & ~n39962;
  assign n39964 = controllable_BtoR_REQ0 & ~n39963;
  assign n39965 = ~n17986 & ~n39964;
  assign n39966 = i_RtoB_ACK0 & ~n39965;
  assign n39967 = ~n17997 & ~n39966;
  assign n39968 = ~controllable_DEQ & ~n39967;
  assign n39969 = ~n39960 & ~n39968;
  assign n39970 = i_FULL & ~n39969;
  assign n39971 = ~n18016 & ~n39958;
  assign n39972 = controllable_DEQ & ~n39971;
  assign n39973 = ~n18032 & ~n39966;
  assign n39974 = ~controllable_DEQ & ~n39973;
  assign n39975 = ~n39972 & ~n39974;
  assign n39976 = ~i_FULL & ~n39975;
  assign n39977 = ~n39970 & ~n39976;
  assign n39978 = i_nEMPTY & ~n39977;
  assign n39979 = ~i_RtoB_ACK1 & ~n38919;
  assign n39980 = ~i_RtoB_ACK1 & ~n39979;
  assign n39981 = ~controllable_BtoR_REQ1 & ~n39980;
  assign n39982 = ~controllable_BtoR_REQ1 & ~n39981;
  assign n39983 = controllable_BtoR_REQ0 & ~n39982;
  assign n39984 = controllable_BtoR_REQ0 & ~n39983;
  assign n39985 = i_RtoB_ACK0 & ~n39984;
  assign n39986 = ~n18053 & ~n39985;
  assign n39987 = controllable_DEQ & ~n39986;
  assign n39988 = ~n11632 & ~n37518;
  assign n39989 = ~controllable_BtoR_REQ1 & ~n39988;
  assign n39990 = ~controllable_BtoR_REQ1 & ~n39989;
  assign n39991 = controllable_BtoR_REQ0 & ~n39990;
  assign n39992 = ~n17967 & ~n39991;
  assign n39993 = i_RtoB_ACK0 & ~n39992;
  assign n39994 = ~n18069 & ~n39993;
  assign n39995 = ~controllable_DEQ & ~n39994;
  assign n39996 = ~n39987 & ~n39995;
  assign n39997 = i_FULL & ~n39996;
  assign n39998 = ~i_RtoB_ACK1 & ~n38876;
  assign n39999 = ~i_RtoB_ACK1 & ~n39998;
  assign n40000 = ~controllable_BtoR_REQ1 & ~n39999;
  assign n40001 = ~controllable_BtoR_REQ1 & ~n40000;
  assign n40002 = controllable_BtoR_REQ0 & ~n40001;
  assign n40003 = controllable_BtoR_REQ0 & ~n40002;
  assign n40004 = i_RtoB_ACK0 & ~n40003;
  assign n40005 = ~n18088 & ~n40004;
  assign n40006 = controllable_DEQ & ~n40005;
  assign n40007 = ~i_RtoB_ACK1 & ~n38949;
  assign n40008 = ~n11632 & ~n40007;
  assign n40009 = ~controllable_BtoR_REQ1 & ~n40008;
  assign n40010 = ~controllable_BtoR_REQ1 & ~n40009;
  assign n40011 = controllable_BtoR_REQ0 & ~n40010;
  assign n40012 = ~n17967 & ~n40011;
  assign n40013 = i_RtoB_ACK0 & ~n40012;
  assign n40014 = ~n18094 & ~n40013;
  assign n40015 = ~controllable_DEQ & ~n40014;
  assign n40016 = ~n40006 & ~n40015;
  assign n40017 = ~i_FULL & ~n40016;
  assign n40018 = ~n39997 & ~n40017;
  assign n40019 = ~i_nEMPTY & ~n40018;
  assign n40020 = ~n39978 & ~n40019;
  assign n40021 = controllable_BtoS_ACK0 & ~n40020;
  assign n40022 = ~i_RtoB_ACK1 & ~n38973;
  assign n40023 = ~n11779 & ~n40022;
  assign n40024 = ~controllable_BtoR_REQ1 & ~n40023;
  assign n40025 = ~controllable_BtoR_REQ1 & ~n40024;
  assign n40026 = controllable_BtoR_REQ0 & ~n40025;
  assign n40027 = ~n18109 & ~n40026;
  assign n40028 = i_RtoB_ACK0 & ~n40027;
  assign n40029 = ~n18120 & ~n40028;
  assign n40030 = controllable_DEQ & ~n40029;
  assign n40031 = ~n11822 & ~n37719;
  assign n40032 = ~controllable_BtoR_REQ1 & ~n40031;
  assign n40033 = ~controllable_BtoR_REQ1 & ~n40032;
  assign n40034 = controllable_BtoR_REQ0 & ~n40033;
  assign n40035 = ~n18128 & ~n40034;
  assign n40036 = i_RtoB_ACK0 & ~n40035;
  assign n40037 = ~n18139 & ~n40036;
  assign n40038 = ~controllable_DEQ & ~n40037;
  assign n40039 = ~n40030 & ~n40038;
  assign n40040 = i_FULL & ~n40039;
  assign n40041 = ~n18158 & ~n40028;
  assign n40042 = controllable_DEQ & ~n40041;
  assign n40043 = ~n18174 & ~n40036;
  assign n40044 = ~controllable_DEQ & ~n40043;
  assign n40045 = ~n40042 & ~n40044;
  assign n40046 = ~i_FULL & ~n40045;
  assign n40047 = ~n40040 & ~n40046;
  assign n40048 = i_nEMPTY & ~n40047;
  assign n40049 = ~i_RtoB_ACK1 & ~n39014;
  assign n40050 = ~i_RtoB_ACK1 & ~n40049;
  assign n40051 = ~controllable_BtoR_REQ1 & ~n40050;
  assign n40052 = ~controllable_BtoR_REQ1 & ~n40051;
  assign n40053 = controllable_BtoR_REQ0 & ~n40052;
  assign n40054 = controllable_BtoR_REQ0 & ~n40053;
  assign n40055 = i_RtoB_ACK0 & ~n40054;
  assign n40056 = ~n18195 & ~n40055;
  assign n40057 = controllable_DEQ & ~n40056;
  assign n40058 = ~n11779 & ~n37781;
  assign n40059 = ~controllable_BtoR_REQ1 & ~n40058;
  assign n40060 = ~controllable_BtoR_REQ1 & ~n40059;
  assign n40061 = controllable_BtoR_REQ0 & ~n40060;
  assign n40062 = ~n18109 & ~n40061;
  assign n40063 = i_RtoB_ACK0 & ~n40062;
  assign n40064 = ~n18211 & ~n40063;
  assign n40065 = ~controllable_DEQ & ~n40064;
  assign n40066 = ~n40057 & ~n40065;
  assign n40067 = i_FULL & ~n40066;
  assign n40068 = ~i_RtoB_ACK1 & ~n38971;
  assign n40069 = ~i_RtoB_ACK1 & ~n40068;
  assign n40070 = ~controllable_BtoR_REQ1 & ~n40069;
  assign n40071 = ~controllable_BtoR_REQ1 & ~n40070;
  assign n40072 = controllable_BtoR_REQ0 & ~n40071;
  assign n40073 = controllable_BtoR_REQ0 & ~n40072;
  assign n40074 = i_RtoB_ACK0 & ~n40073;
  assign n40075 = ~n18230 & ~n40074;
  assign n40076 = controllable_DEQ & ~n40075;
  assign n40077 = ~i_RtoB_ACK1 & ~n39044;
  assign n40078 = ~n11779 & ~n40077;
  assign n40079 = ~controllable_BtoR_REQ1 & ~n40078;
  assign n40080 = ~controllable_BtoR_REQ1 & ~n40079;
  assign n40081 = controllable_BtoR_REQ0 & ~n40080;
  assign n40082 = ~n18109 & ~n40081;
  assign n40083 = i_RtoB_ACK0 & ~n40082;
  assign n40084 = ~n18236 & ~n40083;
  assign n40085 = ~controllable_DEQ & ~n40084;
  assign n40086 = ~n40076 & ~n40085;
  assign n40087 = ~i_FULL & ~n40086;
  assign n40088 = ~n40067 & ~n40087;
  assign n40089 = ~i_nEMPTY & ~n40088;
  assign n40090 = ~n40048 & ~n40089;
  assign n40091 = ~controllable_BtoS_ACK0 & ~n40090;
  assign n40092 = ~n40021 & ~n40091;
  assign n40093 = n4465 & ~n40092;
  assign n40094 = ~n7196 & ~n17686;
  assign n40095 = ~controllable_BtoR_REQ1 & ~n40094;
  assign n40096 = ~controllable_BtoR_REQ1 & ~n40095;
  assign n40097 = controllable_BtoR_REQ0 & ~n40096;
  assign n40098 = ~n15274 & ~n40097;
  assign n40099 = i_RtoB_ACK0 & ~n40098;
  assign n40100 = ~n15285 & ~n40099;
  assign n40101 = controllable_DEQ & ~n40100;
  assign n40102 = ~n16921 & ~n40101;
  assign n40103 = i_FULL & ~n40102;
  assign n40104 = ~n15323 & ~n40099;
  assign n40105 = controllable_DEQ & ~n40104;
  assign n40106 = ~n16927 & ~n40105;
  assign n40107 = ~i_FULL & ~n40106;
  assign n40108 = ~n40103 & ~n40107;
  assign n40109 = i_nEMPTY & ~n40108;
  assign n40110 = ~n15360 & ~n17731;
  assign n40111 = controllable_DEQ & ~n40110;
  assign n40112 = ~n16939 & ~n40111;
  assign n40113 = i_FULL & ~n40112;
  assign n40114 = ~n15395 & ~n17764;
  assign n40115 = controllable_DEQ & ~n40114;
  assign n40116 = ~n16943 & ~n40115;
  assign n40117 = ~i_FULL & ~n40116;
  assign n40118 = ~n40113 & ~n40117;
  assign n40119 = ~i_nEMPTY & ~n40118;
  assign n40120 = ~n40109 & ~n40119;
  assign n40121 = ~controllable_BtoS_ACK0 & ~n40120;
  assign n40122 = ~n16904 & ~n40121;
  assign n40123 = ~n4465 & ~n40122;
  assign n40124 = ~n40093 & ~n40123;
  assign n40125 = ~i_StoB_REQ10 & ~n40124;
  assign n40126 = ~n39951 & ~n40125;
  assign n40127 = controllable_BtoS_ACK10 & ~n40126;
  assign n40128 = ~i_RtoB_ACK1 & ~n39106;
  assign n40129 = ~n36637 & ~n40128;
  assign n40130 = ~controllable_BtoR_REQ1 & ~n40129;
  assign n40131 = ~controllable_BtoR_REQ1 & ~n40130;
  assign n40132 = controllable_BtoR_REQ0 & ~n40131;
  assign n40133 = ~n17967 & ~n40132;
  assign n40134 = i_RtoB_ACK0 & ~n40133;
  assign n40135 = ~n39725 & ~n40134;
  assign n40136 = controllable_DEQ & ~n40135;
  assign n40137 = ~n36656 & ~n37915;
  assign n40138 = ~controllable_BtoR_REQ1 & ~n40137;
  assign n40139 = ~controllable_BtoR_REQ1 & ~n40138;
  assign n40140 = controllable_BtoR_REQ0 & ~n40139;
  assign n40141 = ~n17986 & ~n40140;
  assign n40142 = i_RtoB_ACK0 & ~n40141;
  assign n40143 = ~n39734 & ~n40142;
  assign n40144 = ~controllable_DEQ & ~n40143;
  assign n40145 = ~n40136 & ~n40144;
  assign n40146 = i_FULL & ~n40145;
  assign n40147 = ~n39746 & ~n40134;
  assign n40148 = controllable_DEQ & ~n40147;
  assign n40149 = ~n39755 & ~n40142;
  assign n40150 = ~controllable_DEQ & ~n40149;
  assign n40151 = ~n40148 & ~n40150;
  assign n40152 = ~i_FULL & ~n40151;
  assign n40153 = ~n40146 & ~n40152;
  assign n40154 = i_nEMPTY & ~n40153;
  assign n40155 = controllable_BtoR_REQ0 & ~n20238;
  assign n40156 = controllable_BtoR_REQ0 & ~n40155;
  assign n40157 = i_RtoB_ACK0 & ~n40156;
  assign n40158 = ~n39769 & ~n40157;
  assign n40159 = controllable_DEQ & ~n40158;
  assign n40160 = ~n36637 & ~n37948;
  assign n40161 = ~controllable_BtoR_REQ1 & ~n40160;
  assign n40162 = ~controllable_BtoR_REQ1 & ~n40161;
  assign n40163 = controllable_BtoR_REQ0 & ~n40162;
  assign n40164 = ~n17967 & ~n40163;
  assign n40165 = i_RtoB_ACK0 & ~n40164;
  assign n40166 = ~n39778 & ~n40165;
  assign n40167 = ~controllable_DEQ & ~n40166;
  assign n40168 = ~n40159 & ~n40167;
  assign n40169 = i_FULL & ~n40168;
  assign n40170 = controllable_BtoR_REQ0 & ~n18434;
  assign n40171 = i_RtoB_ACK0 & ~n40170;
  assign n40172 = ~n39790 & ~n40171;
  assign n40173 = controllable_DEQ & ~n40172;
  assign n40174 = ~i_RtoB_ACK1 & ~n37967;
  assign n40175 = ~n36637 & ~n40174;
  assign n40176 = ~controllable_BtoR_REQ1 & ~n40175;
  assign n40177 = ~controllable_BtoR_REQ1 & ~n40176;
  assign n40178 = controllable_BtoR_REQ0 & ~n40177;
  assign n40179 = ~n17967 & ~n40178;
  assign n40180 = i_RtoB_ACK0 & ~n40179;
  assign n40181 = ~n39725 & ~n40180;
  assign n40182 = ~controllable_DEQ & ~n40181;
  assign n40183 = ~n40173 & ~n40182;
  assign n40184 = ~i_FULL & ~n40183;
  assign n40185 = ~n40169 & ~n40184;
  assign n40186 = ~i_nEMPTY & ~n40185;
  assign n40187 = ~n40154 & ~n40186;
  assign n40188 = controllable_BtoS_ACK0 & ~n40187;
  assign n40189 = ~i_RtoB_ACK1 & ~n39179;
  assign n40190 = ~n36716 & ~n40189;
  assign n40191 = ~controllable_BtoR_REQ1 & ~n40190;
  assign n40192 = ~controllable_BtoR_REQ1 & ~n40191;
  assign n40193 = controllable_BtoR_REQ0 & ~n40192;
  assign n40194 = ~n18109 & ~n40193;
  assign n40195 = i_RtoB_ACK0 & ~n40194;
  assign n40196 = ~n39807 & ~n40195;
  assign n40197 = controllable_DEQ & ~n40196;
  assign n40198 = ~n36735 & ~n37999;
  assign n40199 = ~controllable_BtoR_REQ1 & ~n40198;
  assign n40200 = ~controllable_BtoR_REQ1 & ~n40199;
  assign n40201 = controllable_BtoR_REQ0 & ~n40200;
  assign n40202 = ~n18128 & ~n40201;
  assign n40203 = i_RtoB_ACK0 & ~n40202;
  assign n40204 = ~n39816 & ~n40203;
  assign n40205 = ~controllable_DEQ & ~n40204;
  assign n40206 = ~n40197 & ~n40205;
  assign n40207 = i_FULL & ~n40206;
  assign n40208 = ~n39828 & ~n40195;
  assign n40209 = controllable_DEQ & ~n40208;
  assign n40210 = ~n39837 & ~n40203;
  assign n40211 = ~controllable_DEQ & ~n40210;
  assign n40212 = ~n40209 & ~n40211;
  assign n40213 = ~i_FULL & ~n40212;
  assign n40214 = ~n40207 & ~n40213;
  assign n40215 = i_nEMPTY & ~n40214;
  assign n40216 = controllable_BtoR_REQ0 & ~n20291;
  assign n40217 = controllable_BtoR_REQ0 & ~n40216;
  assign n40218 = i_RtoB_ACK0 & ~n40217;
  assign n40219 = ~n39851 & ~n40218;
  assign n40220 = controllable_DEQ & ~n40219;
  assign n40221 = ~n36716 & ~n38032;
  assign n40222 = ~controllable_BtoR_REQ1 & ~n40221;
  assign n40223 = ~controllable_BtoR_REQ1 & ~n40222;
  assign n40224 = controllable_BtoR_REQ0 & ~n40223;
  assign n40225 = ~n18109 & ~n40224;
  assign n40226 = i_RtoB_ACK0 & ~n40225;
  assign n40227 = ~n39860 & ~n40226;
  assign n40228 = ~controllable_DEQ & ~n40227;
  assign n40229 = ~n40220 & ~n40228;
  assign n40230 = i_FULL & ~n40229;
  assign n40231 = controllable_BtoR_REQ0 & ~n18462;
  assign n40232 = i_RtoB_ACK0 & ~n40231;
  assign n40233 = ~n39872 & ~n40232;
  assign n40234 = controllable_DEQ & ~n40233;
  assign n40235 = ~i_RtoB_ACK1 & ~n38051;
  assign n40236 = ~n36716 & ~n40235;
  assign n40237 = ~controllable_BtoR_REQ1 & ~n40236;
  assign n40238 = ~controllable_BtoR_REQ1 & ~n40237;
  assign n40239 = controllable_BtoR_REQ0 & ~n40238;
  assign n40240 = ~n18109 & ~n40239;
  assign n40241 = i_RtoB_ACK0 & ~n40240;
  assign n40242 = ~n39807 & ~n40241;
  assign n40243 = ~controllable_DEQ & ~n40242;
  assign n40244 = ~n40234 & ~n40243;
  assign n40245 = ~i_FULL & ~n40244;
  assign n40246 = ~n40230 & ~n40245;
  assign n40247 = ~i_nEMPTY & ~n40246;
  assign n40248 = ~n40215 & ~n40247;
  assign n40249 = ~controllable_BtoS_ACK0 & ~n40248;
  assign n40250 = ~n40188 & ~n40249;
  assign n40251 = n4465 & ~n40250;
  assign n40252 = ~n7607 & ~n18518;
  assign n40253 = ~controllable_BtoR_REQ1 & ~n40252;
  assign n40254 = ~controllable_BtoR_REQ1 & ~n40253;
  assign n40255 = controllable_BtoR_REQ0 & ~n40254;
  assign n40256 = ~n15274 & ~n40255;
  assign n40257 = i_RtoB_ACK0 & ~n40256;
  assign n40258 = ~n15637 & ~n40257;
  assign n40259 = controllable_DEQ & ~n40258;
  assign n40260 = ~n17098 & ~n40259;
  assign n40261 = i_FULL & ~n40260;
  assign n40262 = ~n15658 & ~n40257;
  assign n40263 = controllable_DEQ & ~n40262;
  assign n40264 = ~n17104 & ~n40263;
  assign n40265 = ~i_FULL & ~n40264;
  assign n40266 = ~n40261 & ~n40265;
  assign n40267 = i_nEMPTY & ~n40266;
  assign n40268 = ~n15681 & ~n17925;
  assign n40269 = controllable_DEQ & ~n40268;
  assign n40270 = ~n17116 & ~n40269;
  assign n40271 = i_FULL & ~n40270;
  assign n40272 = ~n15702 & ~n17943;
  assign n40273 = controllable_DEQ & ~n40272;
  assign n40274 = ~n17119 & ~n40273;
  assign n40275 = ~i_FULL & ~n40274;
  assign n40276 = ~n40271 & ~n40275;
  assign n40277 = ~i_nEMPTY & ~n40276;
  assign n40278 = ~n40267 & ~n40277;
  assign n40279 = ~controllable_BtoS_ACK0 & ~n40278;
  assign n40280 = ~n17081 & ~n40279;
  assign n40281 = ~n4465 & ~n40280;
  assign n40282 = ~n40251 & ~n40281;
  assign n40283 = i_StoB_REQ10 & ~n40282;
  assign n40284 = ~n40125 & ~n40283;
  assign n40285 = ~controllable_BtoS_ACK10 & ~n40284;
  assign n40286 = ~n40127 & ~n40285;
  assign n40287 = n4464 & ~n40286;
  assign n40288 = ~i_RtoB_ACK1 & ~n39300;
  assign n40289 = ~n7886 & ~n40288;
  assign n40290 = ~controllable_BtoR_REQ1 & ~n40289;
  assign n40291 = ~controllable_BtoR_REQ1 & ~n40290;
  assign n40292 = controllable_BtoR_REQ0 & ~n40291;
  assign n40293 = ~n15882 & ~n40292;
  assign n40294 = i_RtoB_ACK0 & ~n40293;
  assign n40295 = ~n15893 & ~n40294;
  assign n40296 = controllable_DEQ & ~n40295;
  assign n40297 = ~n17200 & ~n40296;
  assign n40298 = i_FULL & ~n40297;
  assign n40299 = ~n15931 & ~n40294;
  assign n40300 = controllable_DEQ & ~n40299;
  assign n40301 = ~n17206 & ~n40300;
  assign n40302 = ~i_FULL & ~n40301;
  assign n40303 = ~n40298 & ~n40302;
  assign n40304 = i_nEMPTY & ~n40303;
  assign n40305 = ~n15217 & ~n15968;
  assign n40306 = controllable_DEQ & ~n40305;
  assign n40307 = ~n17218 & ~n40306;
  assign n40308 = i_FULL & ~n40307;
  assign n40309 = ~n15245 & ~n16003;
  assign n40310 = controllable_DEQ & ~n40309;
  assign n40311 = ~n17222 & ~n40310;
  assign n40312 = ~i_FULL & ~n40311;
  assign n40313 = ~n40308 & ~n40312;
  assign n40314 = ~i_nEMPTY & ~n40313;
  assign n40315 = ~n40304 & ~n40314;
  assign n40316 = controllable_BtoS_ACK0 & ~n40315;
  assign n40317 = ~i_RtoB_ACK1 & ~n39344;
  assign n40318 = ~n8057 & ~n40317;
  assign n40319 = ~controllable_BtoR_REQ1 & ~n40318;
  assign n40320 = ~controllable_BtoR_REQ1 & ~n40319;
  assign n40321 = controllable_BtoR_REQ0 & ~n40320;
  assign n40322 = ~n16024 & ~n40321;
  assign n40323 = i_RtoB_ACK0 & ~n40322;
  assign n40324 = ~n16035 & ~n40323;
  assign n40325 = controllable_DEQ & ~n40324;
  assign n40326 = ~n17245 & ~n40325;
  assign n40327 = i_FULL & ~n40326;
  assign n40328 = ~n16073 & ~n40323;
  assign n40329 = controllable_DEQ & ~n40328;
  assign n40330 = ~n17251 & ~n40329;
  assign n40331 = ~i_FULL & ~n40330;
  assign n40332 = ~n40327 & ~n40331;
  assign n40333 = i_nEMPTY & ~n40332;
  assign n40334 = ~n16110 & ~n17731;
  assign n40335 = controllable_DEQ & ~n40334;
  assign n40336 = ~n17263 & ~n40335;
  assign n40337 = i_FULL & ~n40336;
  assign n40338 = ~n16145 & ~n17764;
  assign n40339 = controllable_DEQ & ~n40338;
  assign n40340 = ~n17267 & ~n40339;
  assign n40341 = ~i_FULL & ~n40340;
  assign n40342 = ~n40337 & ~n40341;
  assign n40343 = ~i_nEMPTY & ~n40342;
  assign n40344 = ~n40333 & ~n40343;
  assign n40345 = ~controllable_BtoS_ACK0 & ~n40344;
  assign n40346 = ~n40316 & ~n40345;
  assign n40347 = n4465 & ~n40346;
  assign n40348 = ~n8313 & ~n17686;
  assign n40349 = ~controllable_BtoR_REQ1 & ~n40348;
  assign n40350 = ~controllable_BtoR_REQ1 & ~n40349;
  assign n40351 = controllable_BtoR_REQ0 & ~n40350;
  assign n40352 = ~n16255 & ~n40351;
  assign n40353 = i_RtoB_ACK0 & ~n40352;
  assign n40354 = ~n16266 & ~n40353;
  assign n40355 = controllable_DEQ & ~n40354;
  assign n40356 = ~n17329 & ~n40355;
  assign n40357 = i_FULL & ~n40356;
  assign n40358 = ~n16304 & ~n40353;
  assign n40359 = controllable_DEQ & ~n40358;
  assign n40360 = ~n17335 & ~n40359;
  assign n40361 = ~i_FULL & ~n40360;
  assign n40362 = ~n40357 & ~n40361;
  assign n40363 = i_nEMPTY & ~n40362;
  assign n40364 = ~n16341 & ~n17731;
  assign n40365 = controllable_DEQ & ~n40364;
  assign n40366 = ~n17347 & ~n40365;
  assign n40367 = i_FULL & ~n40366;
  assign n40368 = ~n16376 & ~n17764;
  assign n40369 = controllable_DEQ & ~n40368;
  assign n40370 = ~n17351 & ~n40369;
  assign n40371 = ~i_FULL & ~n40370;
  assign n40372 = ~n40367 & ~n40371;
  assign n40373 = ~i_nEMPTY & ~n40372;
  assign n40374 = ~n40363 & ~n40373;
  assign n40375 = ~controllable_BtoS_ACK0 & ~n40374;
  assign n40376 = ~n17312 & ~n40375;
  assign n40377 = ~n4465 & ~n40376;
  assign n40378 = ~n40347 & ~n40377;
  assign n40379 = ~i_StoB_REQ10 & ~n40378;
  assign n40380 = ~n17183 & ~n40379;
  assign n40381 = controllable_BtoS_ACK10 & ~n40380;
  assign n40382 = ~n8461 & ~n17046;
  assign n40383 = ~controllable_BtoR_REQ1 & ~n40382;
  assign n40384 = ~controllable_BtoR_REQ1 & ~n40383;
  assign n40385 = controllable_BtoR_REQ0 & ~n40384;
  assign n40386 = ~n15882 & ~n40385;
  assign n40387 = i_RtoB_ACK0 & ~n40386;
  assign n40388 = ~n16404 & ~n40387;
  assign n40389 = controllable_DEQ & ~n40388;
  assign n40390 = ~n17380 & ~n40389;
  assign n40391 = i_FULL & ~n40390;
  assign n40392 = ~n16425 & ~n40387;
  assign n40393 = controllable_DEQ & ~n40392;
  assign n40394 = ~n17386 & ~n40393;
  assign n40395 = ~i_FULL & ~n40394;
  assign n40396 = ~n40391 & ~n40395;
  assign n40397 = i_nEMPTY & ~n40396;
  assign n40398 = ~n15604 & ~n16448;
  assign n40399 = controllable_DEQ & ~n40398;
  assign n40400 = ~n17398 & ~n40399;
  assign n40401 = i_FULL & ~n40400;
  assign n40402 = ~n15619 & ~n16469;
  assign n40403 = controllable_DEQ & ~n40402;
  assign n40404 = ~n17401 & ~n40403;
  assign n40405 = ~i_FULL & ~n40404;
  assign n40406 = ~n40401 & ~n40405;
  assign n40407 = ~i_nEMPTY & ~n40406;
  assign n40408 = ~n40397 & ~n40407;
  assign n40409 = controllable_BtoS_ACK0 & ~n40408;
  assign n40410 = ~n8540 & ~n18518;
  assign n40411 = ~controllable_BtoR_REQ1 & ~n40410;
  assign n40412 = ~controllable_BtoR_REQ1 & ~n40411;
  assign n40413 = controllable_BtoR_REQ0 & ~n40412;
  assign n40414 = ~n16024 & ~n40413;
  assign n40415 = i_RtoB_ACK0 & ~n40414;
  assign n40416 = ~n16486 & ~n40415;
  assign n40417 = controllable_DEQ & ~n40416;
  assign n40418 = ~n17424 & ~n40417;
  assign n40419 = i_FULL & ~n40418;
  assign n40420 = ~n16507 & ~n40415;
  assign n40421 = controllable_DEQ & ~n40420;
  assign n40422 = ~n17430 & ~n40421;
  assign n40423 = ~i_FULL & ~n40422;
  assign n40424 = ~n40419 & ~n40423;
  assign n40425 = i_nEMPTY & ~n40424;
  assign n40426 = ~n16530 & ~n17925;
  assign n40427 = controllable_DEQ & ~n40426;
  assign n40428 = ~n17442 & ~n40427;
  assign n40429 = i_FULL & ~n40428;
  assign n40430 = ~n16551 & ~n17943;
  assign n40431 = controllable_DEQ & ~n40430;
  assign n40432 = ~n17445 & ~n40431;
  assign n40433 = ~i_FULL & ~n40432;
  assign n40434 = ~n40429 & ~n40433;
  assign n40435 = ~i_nEMPTY & ~n40434;
  assign n40436 = ~n40425 & ~n40435;
  assign n40437 = ~controllable_BtoS_ACK0 & ~n40436;
  assign n40438 = ~n40409 & ~n40437;
  assign n40439 = n4465 & ~n40438;
  assign n40440 = ~n8672 & ~n18518;
  assign n40441 = ~controllable_BtoR_REQ1 & ~n40440;
  assign n40442 = ~controllable_BtoR_REQ1 & ~n40441;
  assign n40443 = controllable_BtoR_REQ0 & ~n40442;
  assign n40444 = ~n16255 & ~n40443;
  assign n40445 = i_RtoB_ACK0 & ~n40444;
  assign n40446 = ~n16613 & ~n40445;
  assign n40447 = controllable_DEQ & ~n40446;
  assign n40448 = ~n17493 & ~n40447;
  assign n40449 = i_FULL & ~n40448;
  assign n40450 = ~n16634 & ~n40445;
  assign n40451 = controllable_DEQ & ~n40450;
  assign n40452 = ~n17499 & ~n40451;
  assign n40453 = ~i_FULL & ~n40452;
  assign n40454 = ~n40449 & ~n40453;
  assign n40455 = i_nEMPTY & ~n40454;
  assign n40456 = ~n16657 & ~n17925;
  assign n40457 = controllable_DEQ & ~n40456;
  assign n40458 = ~n17511 & ~n40457;
  assign n40459 = i_FULL & ~n40458;
  assign n40460 = ~n16678 & ~n17943;
  assign n40461 = controllable_DEQ & ~n40460;
  assign n40462 = ~n17514 & ~n40461;
  assign n40463 = ~i_FULL & ~n40462;
  assign n40464 = ~n40459 & ~n40463;
  assign n40465 = ~i_nEMPTY & ~n40464;
  assign n40466 = ~n40455 & ~n40465;
  assign n40467 = ~controllable_BtoS_ACK0 & ~n40466;
  assign n40468 = ~n17476 & ~n40467;
  assign n40469 = ~n4465 & ~n40468;
  assign n40470 = ~n40439 & ~n40469;
  assign n40471 = i_StoB_REQ10 & ~n40470;
  assign n40472 = ~n40379 & ~n40471;
  assign n40473 = ~controllable_BtoS_ACK10 & ~n40472;
  assign n40474 = ~n40381 & ~n40473;
  assign n40475 = ~n4464 & ~n40474;
  assign n40476 = ~n40287 & ~n40475;
  assign n40477 = ~n4463 & ~n40476;
  assign n40478 = ~n39891 & ~n40477;
  assign n40479 = n4462 & ~n40478;
  assign n40480 = ~n11632 & ~n17276;
  assign n40481 = ~controllable_BtoR_REQ1 & ~n40480;
  assign n40482 = ~controllable_BtoR_REQ1 & ~n40481;
  assign n40483 = controllable_BtoR_REQ0 & ~n40482;
  assign n40484 = ~n17967 & ~n40483;
  assign n40485 = i_RtoB_ACK0 & ~n40484;
  assign n40486 = ~n17978 & ~n40485;
  assign n40487 = controllable_DEQ & ~n40486;
  assign n40488 = ~n18584 & ~n40487;
  assign n40489 = i_FULL & ~n40488;
  assign n40490 = ~n18016 & ~n40485;
  assign n40491 = controllable_DEQ & ~n40490;
  assign n40492 = ~n18590 & ~n40491;
  assign n40493 = ~i_FULL & ~n40492;
  assign n40494 = ~n40489 & ~n40493;
  assign n40495 = i_nEMPTY & ~n40494;
  assign n40496 = ~n15217 & ~n18053;
  assign n40497 = controllable_DEQ & ~n40496;
  assign n40498 = ~n18602 & ~n40497;
  assign n40499 = i_FULL & ~n40498;
  assign n40500 = ~n15245 & ~n18088;
  assign n40501 = controllable_DEQ & ~n40500;
  assign n40502 = ~n18606 & ~n40501;
  assign n40503 = ~i_FULL & ~n40502;
  assign n40504 = ~n40499 & ~n40503;
  assign n40505 = ~i_nEMPTY & ~n40504;
  assign n40506 = ~n40495 & ~n40505;
  assign n40507 = controllable_BtoS_ACK0 & ~n40506;
  assign n40508 = ~n11779 & ~n17686;
  assign n40509 = ~controllable_BtoR_REQ1 & ~n40508;
  assign n40510 = ~controllable_BtoR_REQ1 & ~n40509;
  assign n40511 = controllable_BtoR_REQ0 & ~n40510;
  assign n40512 = ~n18109 & ~n40511;
  assign n40513 = i_RtoB_ACK0 & ~n40512;
  assign n40514 = ~n18120 & ~n40513;
  assign n40515 = controllable_DEQ & ~n40514;
  assign n40516 = ~n18629 & ~n40515;
  assign n40517 = i_FULL & ~n40516;
  assign n40518 = ~n18158 & ~n40513;
  assign n40519 = controllable_DEQ & ~n40518;
  assign n40520 = ~n18635 & ~n40519;
  assign n40521 = ~i_FULL & ~n40520;
  assign n40522 = ~n40517 & ~n40521;
  assign n40523 = i_nEMPTY & ~n40522;
  assign n40524 = ~n17731 & ~n18195;
  assign n40525 = controllable_DEQ & ~n40524;
  assign n40526 = ~n18647 & ~n40525;
  assign n40527 = i_FULL & ~n40526;
  assign n40528 = ~n17764 & ~n18230;
  assign n40529 = controllable_DEQ & ~n40528;
  assign n40530 = ~n18651 & ~n40529;
  assign n40531 = ~i_FULL & ~n40530;
  assign n40532 = ~n40527 & ~n40531;
  assign n40533 = ~i_nEMPTY & ~n40532;
  assign n40534 = ~n40523 & ~n40533;
  assign n40535 = ~controllable_BtoS_ACK0 & ~n40534;
  assign n40536 = ~n40507 & ~n40535;
  assign n40537 = n4465 & ~n40536;
  assign n40538 = ~n18683 & ~n40121;
  assign n40539 = ~n4465 & ~n40538;
  assign n40540 = ~n40537 & ~n40539;
  assign n40541 = ~i_StoB_REQ10 & ~n40540;
  assign n40542 = ~n18567 & ~n40541;
  assign n40543 = ~controllable_BtoS_ACK10 & ~n40542;
  assign n40544 = ~n18486 & ~n40543;
  assign n40545 = n4464 & ~n40544;
  assign n40546 = ~n7886 & ~n17276;
  assign n40547 = ~controllable_BtoR_REQ1 & ~n40546;
  assign n40548 = ~controllable_BtoR_REQ1 & ~n40547;
  assign n40549 = controllable_BtoR_REQ0 & ~n40548;
  assign n40550 = ~n15882 & ~n40549;
  assign n40551 = i_RtoB_ACK0 & ~n40550;
  assign n40552 = ~n15893 & ~n40551;
  assign n40553 = controllable_DEQ & ~n40552;
  assign n40554 = ~n18778 & ~n40553;
  assign n40555 = i_FULL & ~n40554;
  assign n40556 = ~n15931 & ~n40551;
  assign n40557 = controllable_DEQ & ~n40556;
  assign n40558 = ~n18784 & ~n40557;
  assign n40559 = ~i_FULL & ~n40558;
  assign n40560 = ~n40555 & ~n40559;
  assign n40561 = i_nEMPTY & ~n40560;
  assign n40562 = ~n18796 & ~n40306;
  assign n40563 = i_FULL & ~n40562;
  assign n40564 = ~n18800 & ~n40310;
  assign n40565 = ~i_FULL & ~n40564;
  assign n40566 = ~n40563 & ~n40565;
  assign n40567 = ~i_nEMPTY & ~n40566;
  assign n40568 = ~n40561 & ~n40567;
  assign n40569 = controllable_BtoS_ACK0 & ~n40568;
  assign n40570 = ~n8057 & ~n17686;
  assign n40571 = ~controllable_BtoR_REQ1 & ~n40570;
  assign n40572 = ~controllable_BtoR_REQ1 & ~n40571;
  assign n40573 = controllable_BtoR_REQ0 & ~n40572;
  assign n40574 = ~n16024 & ~n40573;
  assign n40575 = i_RtoB_ACK0 & ~n40574;
  assign n40576 = ~n16035 & ~n40575;
  assign n40577 = controllable_DEQ & ~n40576;
  assign n40578 = ~n18823 & ~n40577;
  assign n40579 = i_FULL & ~n40578;
  assign n40580 = ~n16073 & ~n40575;
  assign n40581 = controllable_DEQ & ~n40580;
  assign n40582 = ~n18829 & ~n40581;
  assign n40583 = ~i_FULL & ~n40582;
  assign n40584 = ~n40579 & ~n40583;
  assign n40585 = i_nEMPTY & ~n40584;
  assign n40586 = ~n18841 & ~n40335;
  assign n40587 = i_FULL & ~n40586;
  assign n40588 = ~n18845 & ~n40339;
  assign n40589 = ~i_FULL & ~n40588;
  assign n40590 = ~n40587 & ~n40589;
  assign n40591 = ~i_nEMPTY & ~n40590;
  assign n40592 = ~n40585 & ~n40591;
  assign n40593 = ~controllable_BtoS_ACK0 & ~n40592;
  assign n40594 = ~n40569 & ~n40593;
  assign n40595 = n4465 & ~n40594;
  assign n40596 = ~n40377 & ~n40595;
  assign n40597 = ~i_StoB_REQ10 & ~n40596;
  assign n40598 = ~n18761 & ~n40597;
  assign n40599 = ~controllable_BtoS_ACK10 & ~n40598;
  assign n40600 = ~n18693 & ~n40599;
  assign n40601 = ~n4464 & ~n40600;
  assign n40602 = ~n40545 & ~n40601;
  assign n40603 = ~n4463 & ~n40602;
  assign n40604 = ~n18424 & ~n40603;
  assign n40605 = ~n4462 & ~n40604;
  assign n40606 = ~n40479 & ~n40605;
  assign n40607 = n4461 & ~n40606;
  assign n40608 = ~controllable_BtoR_REQ1 & ~n36887;
  assign n40609 = ~controllable_BtoR_REQ1 & ~n40608;
  assign n40610 = ~controllable_BtoR_REQ0 & ~n40609;
  assign n40611 = ~n17562 & ~n40610;
  assign n40612 = ~i_RtoB_ACK0 & ~n40611;
  assign n40613 = ~n39897 & ~n40612;
  assign n40614 = ~controllable_DEQ & ~n40613;
  assign n40615 = ~n20225 & ~n40614;
  assign n40616 = i_FULL & ~n40615;
  assign n40617 = ~n36886 & ~n36899;
  assign n40618 = ~controllable_BtoR_REQ1 & ~n40617;
  assign n40619 = ~controllable_BtoR_REQ1 & ~n40618;
  assign n40620 = ~controllable_BtoR_REQ0 & ~n40619;
  assign n40621 = ~n17562 & ~n40620;
  assign n40622 = ~i_RtoB_ACK0 & ~n40621;
  assign n40623 = ~n39897 & ~n40622;
  assign n40624 = ~controllable_DEQ & ~n40623;
  assign n40625 = ~n20225 & ~n40624;
  assign n40626 = ~i_FULL & ~n40625;
  assign n40627 = ~n40616 & ~n40626;
  assign n40628 = i_nEMPTY & ~n40627;
  assign n40629 = ~controllable_BtoR_REQ1 & ~n36922;
  assign n40630 = ~controllable_BtoR_REQ1 & ~n40629;
  assign n40631 = ~controllable_BtoR_REQ0 & ~n40630;
  assign n40632 = ~n17581 & ~n40631;
  assign n40633 = ~i_RtoB_ACK0 & ~n40632;
  assign n40634 = ~n39907 & ~n40633;
  assign n40635 = ~controllable_DEQ & ~n40634;
  assign n40636 = ~n20243 & ~n40635;
  assign n40637 = i_FULL & ~n40636;
  assign n40638 = ~n36921 & ~n37040;
  assign n40639 = ~controllable_BtoR_REQ1 & ~n40638;
  assign n40640 = ~controllable_BtoR_REQ1 & ~n40639;
  assign n40641 = ~controllable_BtoR_REQ0 & ~n40640;
  assign n40642 = ~n17545 & ~n40641;
  assign n40643 = ~i_RtoB_ACK0 & ~n40642;
  assign n40644 = ~n39907 & ~n40643;
  assign n40645 = ~controllable_DEQ & ~n40644;
  assign n40646 = ~n20258 & ~n40645;
  assign n40647 = ~i_FULL & ~n40646;
  assign n40648 = ~n40637 & ~n40647;
  assign n40649 = ~i_nEMPTY & ~n40648;
  assign n40650 = ~n40628 & ~n40649;
  assign n40651 = controllable_BtoS_ACK0 & ~n40650;
  assign n40652 = ~controllable_BtoR_REQ1 & ~n37068;
  assign n40653 = ~controllable_BtoR_REQ1 & ~n40652;
  assign n40654 = ~controllable_BtoR_REQ0 & ~n40653;
  assign n40655 = ~n14841 & ~n40654;
  assign n40656 = ~i_RtoB_ACK0 & ~n40655;
  assign n40657 = ~n39925 & ~n40656;
  assign n40658 = ~controllable_DEQ & ~n40657;
  assign n40659 = ~n20280 & ~n40658;
  assign n40660 = i_FULL & ~n40659;
  assign n40661 = ~n37067 & ~n37080;
  assign n40662 = ~controllable_BtoR_REQ1 & ~n40661;
  assign n40663 = ~controllable_BtoR_REQ1 & ~n40662;
  assign n40664 = ~controllable_BtoR_REQ0 & ~n40663;
  assign n40665 = ~n14841 & ~n40664;
  assign n40666 = ~i_RtoB_ACK0 & ~n40665;
  assign n40667 = ~n39925 & ~n40666;
  assign n40668 = ~controllable_DEQ & ~n40667;
  assign n40669 = ~n20280 & ~n40668;
  assign n40670 = ~i_FULL & ~n40669;
  assign n40671 = ~n40660 & ~n40670;
  assign n40672 = i_nEMPTY & ~n40671;
  assign n40673 = ~controllable_BtoR_REQ1 & ~n37103;
  assign n40674 = ~controllable_BtoR_REQ1 & ~n40673;
  assign n40675 = ~controllable_BtoR_REQ0 & ~n40674;
  assign n40676 = ~n14860 & ~n40675;
  assign n40677 = ~i_RtoB_ACK0 & ~n40676;
  assign n40678 = ~n39935 & ~n40677;
  assign n40679 = ~controllable_DEQ & ~n40678;
  assign n40680 = ~n20296 & ~n40679;
  assign n40681 = i_FULL & ~n40680;
  assign n40682 = ~n37102 & ~n37126;
  assign n40683 = ~controllable_BtoR_REQ1 & ~n40682;
  assign n40684 = ~controllable_BtoR_REQ1 & ~n40683;
  assign n40685 = ~controllable_BtoR_REQ0 & ~n40684;
  assign n40686 = ~n14824 & ~n40685;
  assign n40687 = ~i_RtoB_ACK0 & ~n40686;
  assign n40688 = ~n39935 & ~n40687;
  assign n40689 = ~controllable_DEQ & ~n40688;
  assign n40690 = ~n20311 & ~n40689;
  assign n40691 = ~i_FULL & ~n40690;
  assign n40692 = ~n40681 & ~n40691;
  assign n40693 = ~i_nEMPTY & ~n40692;
  assign n40694 = ~n40672 & ~n40693;
  assign n40695 = ~controllable_BtoS_ACK0 & ~n40694;
  assign n40696 = ~n40651 & ~n40695;
  assign n40697 = n4465 & ~n40696;
  assign n40698 = ~n19016 & ~n19022;
  assign n40699 = i_FULL & ~n40698;
  assign n40700 = ~n19032 & ~n40699;
  assign n40701 = i_nEMPTY & ~n40700;
  assign n40702 = ~n19063 & ~n40701;
  assign n40703 = ~controllable_BtoS_ACK0 & ~n40702;
  assign n40704 = ~n14811 & ~n40703;
  assign n40705 = ~n4465 & ~n40704;
  assign n40706 = ~n40697 & ~n40705;
  assign n40707 = i_StoB_REQ10 & ~n40706;
  assign n40708 = ~n17280 & ~n17967;
  assign n40709 = i_RtoB_ACK0 & ~n40708;
  assign n40710 = i_RtoB_ACK1 & ~n37247;
  assign n40711 = ~n37259 & ~n40710;
  assign n40712 = ~controllable_BtoR_REQ1 & ~n40711;
  assign n40713 = ~controllable_BtoR_REQ1 & ~n40712;
  assign n40714 = ~controllable_BtoR_REQ0 & ~n40713;
  assign n40715 = ~n17974 & ~n40714;
  assign n40716 = ~i_RtoB_ACK0 & ~n40715;
  assign n40717 = ~n40709 & ~n40716;
  assign n40718 = controllable_DEQ & ~n40717;
  assign n40719 = ~n11675 & ~n37915;
  assign n40720 = ~controllable_BtoR_REQ1 & ~n40719;
  assign n40721 = ~controllable_BtoR_REQ1 & ~n40720;
  assign n40722 = controllable_BtoR_REQ0 & ~n40721;
  assign n40723 = ~n17986 & ~n40722;
  assign n40724 = i_RtoB_ACK0 & ~n40723;
  assign n40725 = ~n12387 & ~n38888;
  assign n40726 = ~controllable_BtoR_REQ1 & ~n40725;
  assign n40727 = ~controllable_BtoR_REQ1 & ~n40726;
  assign n40728 = ~controllable_BtoR_REQ0 & ~n40727;
  assign n40729 = ~n17993 & ~n40728;
  assign n40730 = ~i_RtoB_ACK0 & ~n40729;
  assign n40731 = ~n40724 & ~n40730;
  assign n40732 = ~controllable_DEQ & ~n40731;
  assign n40733 = ~n40718 & ~n40732;
  assign n40734 = i_FULL & ~n40733;
  assign n40735 = ~n18012 & ~n40714;
  assign n40736 = ~i_RtoB_ACK0 & ~n40735;
  assign n40737 = ~n40709 & ~n40736;
  assign n40738 = controllable_DEQ & ~n40737;
  assign n40739 = ~n37491 & ~n38888;
  assign n40740 = ~controllable_BtoR_REQ1 & ~n40739;
  assign n40741 = ~controllable_BtoR_REQ1 & ~n40740;
  assign n40742 = ~controllable_BtoR_REQ0 & ~n40741;
  assign n40743 = ~n18028 & ~n40742;
  assign n40744 = ~i_RtoB_ACK0 & ~n40743;
  assign n40745 = ~n40724 & ~n40744;
  assign n40746 = ~controllable_DEQ & ~n40745;
  assign n40747 = ~n40738 & ~n40746;
  assign n40748 = ~i_FULL & ~n40747;
  assign n40749 = ~n40734 & ~n40748;
  assign n40750 = i_nEMPTY & ~n40749;
  assign n40751 = ~controllable_BtoR_REQ1 & ~n37509;
  assign n40752 = ~controllable_BtoR_REQ0 & ~n40751;
  assign n40753 = ~n18049 & ~n40752;
  assign n40754 = ~i_RtoB_ACK0 & ~n40753;
  assign n40755 = ~n15217 & ~n40754;
  assign n40756 = controllable_DEQ & ~n40755;
  assign n40757 = ~n11632 & ~n37948;
  assign n40758 = ~controllable_BtoR_REQ1 & ~n40757;
  assign n40759 = ~controllable_BtoR_REQ1 & ~n40758;
  assign n40760 = controllable_BtoR_REQ0 & ~n40759;
  assign n40761 = ~n17967 & ~n40760;
  assign n40762 = i_RtoB_ACK0 & ~n40761;
  assign n40763 = ~n12431 & ~n38929;
  assign n40764 = ~controllable_BtoR_REQ1 & ~n40763;
  assign n40765 = ~controllable_BtoR_REQ1 & ~n40764;
  assign n40766 = ~controllable_BtoR_REQ0 & ~n40765;
  assign n40767 = ~n18065 & ~n40766;
  assign n40768 = ~i_RtoB_ACK0 & ~n40767;
  assign n40769 = ~n40762 & ~n40768;
  assign n40770 = ~controllable_DEQ & ~n40769;
  assign n40771 = ~n40756 & ~n40770;
  assign n40772 = i_FULL & ~n40771;
  assign n40773 = ~controllable_BtoR_REQ1 & ~n37542;
  assign n40774 = ~controllable_BtoR_REQ0 & ~n40773;
  assign n40775 = ~n18084 & ~n40774;
  assign n40776 = ~i_RtoB_ACK0 & ~n40775;
  assign n40777 = ~n15245 & ~n40776;
  assign n40778 = controllable_DEQ & ~n40777;
  assign n40779 = ~i_RtoB_ACK1 & ~n37549;
  assign n40780 = ~n11632 & ~n40779;
  assign n40781 = ~controllable_BtoR_REQ1 & ~n40780;
  assign n40782 = ~controllable_BtoR_REQ1 & ~n40781;
  assign n40783 = controllable_BtoR_REQ0 & ~n40782;
  assign n40784 = ~n17967 & ~n40783;
  assign n40785 = i_RtoB_ACK0 & ~n40784;
  assign n40786 = ~n37664 & ~n38929;
  assign n40787 = ~controllable_BtoR_REQ1 & ~n40786;
  assign n40788 = ~controllable_BtoR_REQ1 & ~n40787;
  assign n40789 = ~controllable_BtoR_REQ0 & ~n40788;
  assign n40790 = ~n17974 & ~n40789;
  assign n40791 = ~i_RtoB_ACK0 & ~n40790;
  assign n40792 = ~n40785 & ~n40791;
  assign n40793 = ~controllable_DEQ & ~n40792;
  assign n40794 = ~n40778 & ~n40793;
  assign n40795 = ~i_FULL & ~n40794;
  assign n40796 = ~n40772 & ~n40795;
  assign n40797 = ~i_nEMPTY & ~n40796;
  assign n40798 = ~n40750 & ~n40797;
  assign n40799 = controllable_BtoS_ACK0 & ~n40798;
  assign n40800 = ~n17690 & ~n18109;
  assign n40801 = i_RtoB_ACK0 & ~n40800;
  assign n40802 = i_RtoB_ACK1 & ~n37689;
  assign n40803 = ~n37701 & ~n40802;
  assign n40804 = ~controllable_BtoR_REQ1 & ~n40803;
  assign n40805 = ~controllable_BtoR_REQ1 & ~n40804;
  assign n40806 = ~controllable_BtoR_REQ0 & ~n40805;
  assign n40807 = ~n18116 & ~n40806;
  assign n40808 = ~i_RtoB_ACK0 & ~n40807;
  assign n40809 = ~n40801 & ~n40808;
  assign n40810 = controllable_DEQ & ~n40809;
  assign n40811 = ~n11822 & ~n37999;
  assign n40812 = ~controllable_BtoR_REQ1 & ~n40811;
  assign n40813 = ~controllable_BtoR_REQ1 & ~n40812;
  assign n40814 = controllable_BtoR_REQ0 & ~n40813;
  assign n40815 = ~n18128 & ~n40814;
  assign n40816 = i_RtoB_ACK0 & ~n40815;
  assign n40817 = ~n9913 & ~n38983;
  assign n40818 = ~controllable_BtoR_REQ1 & ~n40817;
  assign n40819 = ~controllable_BtoR_REQ1 & ~n40818;
  assign n40820 = ~controllable_BtoR_REQ0 & ~n40819;
  assign n40821 = ~n18135 & ~n40820;
  assign n40822 = ~i_RtoB_ACK0 & ~n40821;
  assign n40823 = ~n40816 & ~n40822;
  assign n40824 = ~controllable_DEQ & ~n40823;
  assign n40825 = ~n40810 & ~n40824;
  assign n40826 = i_FULL & ~n40825;
  assign n40827 = ~n18154 & ~n40806;
  assign n40828 = ~i_RtoB_ACK0 & ~n40827;
  assign n40829 = ~n40801 & ~n40828;
  assign n40830 = controllable_DEQ & ~n40829;
  assign n40831 = ~n37754 & ~n38983;
  assign n40832 = ~controllable_BtoR_REQ1 & ~n40831;
  assign n40833 = ~controllable_BtoR_REQ1 & ~n40832;
  assign n40834 = ~controllable_BtoR_REQ0 & ~n40833;
  assign n40835 = ~n18170 & ~n40834;
  assign n40836 = ~i_RtoB_ACK0 & ~n40835;
  assign n40837 = ~n40816 & ~n40836;
  assign n40838 = ~controllable_DEQ & ~n40837;
  assign n40839 = ~n40830 & ~n40838;
  assign n40840 = ~i_FULL & ~n40839;
  assign n40841 = ~n40826 & ~n40840;
  assign n40842 = i_nEMPTY & ~n40841;
  assign n40843 = ~controllable_BtoR_REQ1 & ~n37772;
  assign n40844 = ~controllable_BtoR_REQ0 & ~n40843;
  assign n40845 = ~n18191 & ~n40844;
  assign n40846 = ~i_RtoB_ACK0 & ~n40845;
  assign n40847 = ~n17731 & ~n40846;
  assign n40848 = controllable_DEQ & ~n40847;
  assign n40849 = ~n11779 & ~n38032;
  assign n40850 = ~controllable_BtoR_REQ1 & ~n40849;
  assign n40851 = ~controllable_BtoR_REQ1 & ~n40850;
  assign n40852 = controllable_BtoR_REQ0 & ~n40851;
  assign n40853 = ~n18109 & ~n40852;
  assign n40854 = i_RtoB_ACK0 & ~n40853;
  assign n40855 = ~n9961 & ~n39024;
  assign n40856 = ~controllable_BtoR_REQ1 & ~n40855;
  assign n40857 = ~controllable_BtoR_REQ1 & ~n40856;
  assign n40858 = ~controllable_BtoR_REQ0 & ~n40857;
  assign n40859 = ~n18207 & ~n40858;
  assign n40860 = ~i_RtoB_ACK0 & ~n40859;
  assign n40861 = ~n40854 & ~n40860;
  assign n40862 = ~controllable_DEQ & ~n40861;
  assign n40863 = ~n40848 & ~n40862;
  assign n40864 = i_FULL & ~n40863;
  assign n40865 = ~controllable_BtoR_REQ1 & ~n37805;
  assign n40866 = ~controllable_BtoR_REQ0 & ~n40865;
  assign n40867 = ~n18226 & ~n40866;
  assign n40868 = ~i_RtoB_ACK0 & ~n40867;
  assign n40869 = ~n17764 & ~n40868;
  assign n40870 = controllable_DEQ & ~n40869;
  assign n40871 = ~i_RtoB_ACK1 & ~n37812;
  assign n40872 = ~n11779 & ~n40871;
  assign n40873 = ~controllable_BtoR_REQ1 & ~n40872;
  assign n40874 = ~controllable_BtoR_REQ1 & ~n40873;
  assign n40875 = controllable_BtoR_REQ0 & ~n40874;
  assign n40876 = ~n18109 & ~n40875;
  assign n40877 = i_RtoB_ACK0 & ~n40876;
  assign n40878 = ~n37826 & ~n39024;
  assign n40879 = ~controllable_BtoR_REQ1 & ~n40878;
  assign n40880 = ~controllable_BtoR_REQ1 & ~n40879;
  assign n40881 = ~controllable_BtoR_REQ0 & ~n40880;
  assign n40882 = ~n18116 & ~n40881;
  assign n40883 = ~i_RtoB_ACK0 & ~n40882;
  assign n40884 = ~n40877 & ~n40883;
  assign n40885 = ~controllable_DEQ & ~n40884;
  assign n40886 = ~n40870 & ~n40885;
  assign n40887 = ~i_FULL & ~n40886;
  assign n40888 = ~n40864 & ~n40887;
  assign n40889 = ~i_nEMPTY & ~n40888;
  assign n40890 = ~n40842 & ~n40889;
  assign n40891 = ~controllable_BtoS_ACK0 & ~n40890;
  assign n40892 = ~n40799 & ~n40891;
  assign n40893 = n4465 & ~n40892;
  assign n40894 = ~n15274 & ~n17690;
  assign n40895 = i_RtoB_ACK0 & ~n40894;
  assign n40896 = ~n15281 & ~n17701;
  assign n40897 = ~i_RtoB_ACK0 & ~n40896;
  assign n40898 = ~n40895 & ~n40897;
  assign n40899 = controllable_DEQ & ~n40898;
  assign n40900 = ~n19327 & ~n40899;
  assign n40901 = i_FULL & ~n40900;
  assign n40902 = ~n19331 & ~n40895;
  assign n40903 = controllable_DEQ & ~n40902;
  assign n40904 = ~n19341 & ~n40903;
  assign n40905 = ~i_FULL & ~n40904;
  assign n40906 = ~n40901 & ~n40905;
  assign n40907 = i_nEMPTY & ~n40906;
  assign n40908 = ~n17731 & ~n19347;
  assign n40909 = controllable_DEQ & ~n40908;
  assign n40910 = ~n19357 & ~n40909;
  assign n40911 = i_FULL & ~n40910;
  assign n40912 = ~n17764 & ~n19361;
  assign n40913 = controllable_DEQ & ~n40912;
  assign n40914 = ~n19371 & ~n40913;
  assign n40915 = ~i_FULL & ~n40914;
  assign n40916 = ~n40911 & ~n40915;
  assign n40917 = ~i_nEMPTY & ~n40916;
  assign n40918 = ~n40907 & ~n40917;
  assign n40919 = ~controllable_BtoS_ACK0 & ~n40918;
  assign n40920 = ~n19311 & ~n40919;
  assign n40921 = ~n4465 & ~n40920;
  assign n40922 = ~n40893 & ~n40921;
  assign n40923 = ~i_StoB_REQ10 & ~n40922;
  assign n40924 = ~n40707 & ~n40923;
  assign n40925 = controllable_BtoS_ACK10 & ~n40924;
  assign n40926 = ~n17050 & ~n17967;
  assign n40927 = i_RtoB_ACK0 & ~n40926;
  assign n40928 = controllable_BtoR_REQ0 & ~n17975;
  assign n40929 = ~n17622 & ~n40928;
  assign n40930 = ~i_RtoB_ACK0 & ~n40929;
  assign n40931 = ~n40927 & ~n40930;
  assign n40932 = controllable_DEQ & ~n40931;
  assign n40933 = controllable_BtoR_REQ0 & ~n17994;
  assign n40934 = ~n12387 & ~n37468;
  assign n40935 = ~controllable_BtoR_REQ1 & ~n40934;
  assign n40936 = ~controllable_BtoR_REQ1 & ~n40935;
  assign n40937 = ~controllable_BtoR_REQ0 & ~n40936;
  assign n40938 = ~n40933 & ~n40937;
  assign n40939 = ~i_RtoB_ACK0 & ~n40938;
  assign n40940 = ~n40142 & ~n40939;
  assign n40941 = ~controllable_DEQ & ~n40940;
  assign n40942 = ~n40932 & ~n40941;
  assign n40943 = i_FULL & ~n40942;
  assign n40944 = controllable_BtoR_REQ0 & ~n18013;
  assign n40945 = ~n17622 & ~n40944;
  assign n40946 = ~i_RtoB_ACK0 & ~n40945;
  assign n40947 = ~n40927 & ~n40946;
  assign n40948 = controllable_DEQ & ~n40947;
  assign n40949 = controllable_BtoR_REQ0 & ~n18029;
  assign n40950 = ~n37468 & ~n37491;
  assign n40951 = ~controllable_BtoR_REQ1 & ~n40950;
  assign n40952 = ~controllable_BtoR_REQ1 & ~n40951;
  assign n40953 = ~controllable_BtoR_REQ0 & ~n40952;
  assign n40954 = ~n40949 & ~n40953;
  assign n40955 = ~i_RtoB_ACK0 & ~n40954;
  assign n40956 = ~n40142 & ~n40955;
  assign n40957 = ~controllable_DEQ & ~n40956;
  assign n40958 = ~n40948 & ~n40957;
  assign n40959 = ~i_FULL & ~n40958;
  assign n40960 = ~n40943 & ~n40959;
  assign n40961 = i_nEMPTY & ~n40960;
  assign n40962 = controllable_BtoR_REQ0 & ~n18050;
  assign n40963 = ~n17647 & ~n40962;
  assign n40964 = ~i_RtoB_ACK0 & ~n40963;
  assign n40965 = ~n15604 & ~n40964;
  assign n40966 = controllable_DEQ & ~n40965;
  assign n40967 = controllable_BtoR_REQ0 & ~n18066;
  assign n40968 = ~n12431 & ~n37527;
  assign n40969 = ~controllable_BtoR_REQ1 & ~n40968;
  assign n40970 = ~controllable_BtoR_REQ1 & ~n40969;
  assign n40971 = ~controllable_BtoR_REQ0 & ~n40970;
  assign n40972 = ~n40967 & ~n40971;
  assign n40973 = ~i_RtoB_ACK0 & ~n40972;
  assign n40974 = ~n40165 & ~n40973;
  assign n40975 = ~controllable_DEQ & ~n40974;
  assign n40976 = ~n40966 & ~n40975;
  assign n40977 = i_FULL & ~n40976;
  assign n40978 = controllable_BtoR_REQ0 & ~n18085;
  assign n40979 = ~n17669 & ~n40978;
  assign n40980 = ~i_RtoB_ACK0 & ~n40979;
  assign n40981 = ~n15619 & ~n40980;
  assign n40982 = controllable_DEQ & ~n40981;
  assign n40983 = ~n37491 & ~n37527;
  assign n40984 = ~controllable_BtoR_REQ1 & ~n40983;
  assign n40985 = ~controllable_BtoR_REQ1 & ~n40984;
  assign n40986 = ~controllable_BtoR_REQ0 & ~n40985;
  assign n40987 = ~n40928 & ~n40986;
  assign n40988 = ~i_RtoB_ACK0 & ~n40987;
  assign n40989 = ~n40180 & ~n40988;
  assign n40990 = ~controllable_DEQ & ~n40989;
  assign n40991 = ~n40982 & ~n40990;
  assign n40992 = ~i_FULL & ~n40991;
  assign n40993 = ~n40977 & ~n40992;
  assign n40994 = ~i_nEMPTY & ~n40993;
  assign n40995 = ~n40961 & ~n40994;
  assign n40996 = controllable_BtoS_ACK0 & ~n40995;
  assign n40997 = ~n18109 & ~n18522;
  assign n40998 = i_RtoB_ACK0 & ~n40997;
  assign n40999 = controllable_BtoR_REQ0 & ~n18117;
  assign n41000 = ~n17701 & ~n40999;
  assign n41001 = ~i_RtoB_ACK0 & ~n41000;
  assign n41002 = ~n40998 & ~n41001;
  assign n41003 = controllable_DEQ & ~n41002;
  assign n41004 = controllable_BtoR_REQ0 & ~n18136;
  assign n41005 = ~n9913 & ~n37731;
  assign n41006 = ~controllable_BtoR_REQ1 & ~n41005;
  assign n41007 = ~controllable_BtoR_REQ1 & ~n41006;
  assign n41008 = ~controllable_BtoR_REQ0 & ~n41007;
  assign n41009 = ~n41004 & ~n41008;
  assign n41010 = ~i_RtoB_ACK0 & ~n41009;
  assign n41011 = ~n40203 & ~n41010;
  assign n41012 = ~controllable_DEQ & ~n41011;
  assign n41013 = ~n41003 & ~n41012;
  assign n41014 = i_FULL & ~n41013;
  assign n41015 = controllable_BtoR_REQ0 & ~n18155;
  assign n41016 = ~n17701 & ~n41015;
  assign n41017 = ~i_RtoB_ACK0 & ~n41016;
  assign n41018 = ~n40998 & ~n41017;
  assign n41019 = controllable_DEQ & ~n41018;
  assign n41020 = controllable_BtoR_REQ0 & ~n18171;
  assign n41021 = ~n37731 & ~n37754;
  assign n41022 = ~controllable_BtoR_REQ1 & ~n41021;
  assign n41023 = ~controllable_BtoR_REQ1 & ~n41022;
  assign n41024 = ~controllable_BtoR_REQ0 & ~n41023;
  assign n41025 = ~n41020 & ~n41024;
  assign n41026 = ~i_RtoB_ACK0 & ~n41025;
  assign n41027 = ~n40203 & ~n41026;
  assign n41028 = ~controllable_DEQ & ~n41027;
  assign n41029 = ~n41019 & ~n41028;
  assign n41030 = ~i_FULL & ~n41029;
  assign n41031 = ~n41014 & ~n41030;
  assign n41032 = i_nEMPTY & ~n41031;
  assign n41033 = controllable_BtoR_REQ0 & ~n18192;
  assign n41034 = ~n17737 & ~n41033;
  assign n41035 = ~i_RtoB_ACK0 & ~n41034;
  assign n41036 = ~n17925 & ~n41035;
  assign n41037 = controllable_DEQ & ~n41036;
  assign n41038 = controllable_BtoR_REQ0 & ~n18208;
  assign n41039 = ~n9961 & ~n37790;
  assign n41040 = ~controllable_BtoR_REQ1 & ~n41039;
  assign n41041 = ~controllable_BtoR_REQ1 & ~n41040;
  assign n41042 = ~controllable_BtoR_REQ0 & ~n41041;
  assign n41043 = ~n41038 & ~n41042;
  assign n41044 = ~i_RtoB_ACK0 & ~n41043;
  assign n41045 = ~n40226 & ~n41044;
  assign n41046 = ~controllable_DEQ & ~n41045;
  assign n41047 = ~n41037 & ~n41046;
  assign n41048 = i_FULL & ~n41047;
  assign n41049 = controllable_BtoR_REQ0 & ~n18227;
  assign n41050 = ~n17770 & ~n41049;
  assign n41051 = ~i_RtoB_ACK0 & ~n41050;
  assign n41052 = ~n17943 & ~n41051;
  assign n41053 = controllable_DEQ & ~n41052;
  assign n41054 = ~n37754 & ~n37790;
  assign n41055 = ~controllable_BtoR_REQ1 & ~n41054;
  assign n41056 = ~controllable_BtoR_REQ1 & ~n41055;
  assign n41057 = ~controllable_BtoR_REQ0 & ~n41056;
  assign n41058 = ~n40999 & ~n41057;
  assign n41059 = ~i_RtoB_ACK0 & ~n41058;
  assign n41060 = ~n40241 & ~n41059;
  assign n41061 = ~controllable_DEQ & ~n41060;
  assign n41062 = ~n41053 & ~n41061;
  assign n41063 = ~i_FULL & ~n41062;
  assign n41064 = ~n41048 & ~n41063;
  assign n41065 = ~i_nEMPTY & ~n41064;
  assign n41066 = ~n41032 & ~n41065;
  assign n41067 = ~controllable_BtoS_ACK0 & ~n41066;
  assign n41068 = ~n40996 & ~n41067;
  assign n41069 = n4465 & ~n41068;
  assign n41070 = ~n15274 & ~n18522;
  assign n41071 = i_RtoB_ACK0 & ~n41070;
  assign n41072 = ~n17701 & ~n19554;
  assign n41073 = ~i_RtoB_ACK0 & ~n41072;
  assign n41074 = ~n41071 & ~n41073;
  assign n41075 = controllable_DEQ & ~n41074;
  assign n41076 = ~n19563 & ~n41075;
  assign n41077 = i_FULL & ~n41076;
  assign n41078 = ~n19568 & ~n41071;
  assign n41079 = controllable_DEQ & ~n41078;
  assign n41080 = ~n19575 & ~n41079;
  assign n41081 = ~i_FULL & ~n41080;
  assign n41082 = ~n41077 & ~n41081;
  assign n41083 = i_nEMPTY & ~n41082;
  assign n41084 = ~n17925 & ~n19582;
  assign n41085 = controllable_DEQ & ~n41084;
  assign n41086 = ~n19589 & ~n41085;
  assign n41087 = i_FULL & ~n41086;
  assign n41088 = ~n17943 & ~n19594;
  assign n41089 = controllable_DEQ & ~n41088;
  assign n41090 = ~n19597 & ~n41089;
  assign n41091 = ~i_FULL & ~n41090;
  assign n41092 = ~n41087 & ~n41091;
  assign n41093 = ~i_nEMPTY & ~n41092;
  assign n41094 = ~n41083 & ~n41093;
  assign n41095 = ~controllable_BtoS_ACK0 & ~n41094;
  assign n41096 = ~n19553 & ~n41095;
  assign n41097 = ~n4465 & ~n41096;
  assign n41098 = ~n41069 & ~n41097;
  assign n41099 = i_StoB_REQ10 & ~n41098;
  assign n41100 = ~n40923 & ~n41099;
  assign n41101 = ~controllable_BtoS_ACK10 & ~n41100;
  assign n41102 = ~n40925 & ~n41101;
  assign n41103 = n4464 & ~n41102;
  assign n41104 = ~n19626 & ~n19632;
  assign n41105 = i_FULL & ~n41104;
  assign n41106 = ~n19642 & ~n41105;
  assign n41107 = i_nEMPTY & ~n41106;
  assign n41108 = ~n19673 & ~n41107;
  assign n41109 = controllable_BtoS_ACK0 & ~n41108;
  assign n41110 = ~n19690 & ~n19696;
  assign n41111 = i_FULL & ~n41110;
  assign n41112 = ~n19706 & ~n41111;
  assign n41113 = i_nEMPTY & ~n41112;
  assign n41114 = ~n19737 & ~n41113;
  assign n41115 = ~controllable_BtoS_ACK0 & ~n41114;
  assign n41116 = ~n41109 & ~n41115;
  assign n41117 = n4465 & ~n41116;
  assign n41118 = ~n14811 & ~n41115;
  assign n41119 = ~n4465 & ~n41118;
  assign n41120 = ~n41117 & ~n41119;
  assign n41121 = i_StoB_REQ10 & ~n41120;
  assign n41122 = ~n15882 & ~n17280;
  assign n41123 = i_RtoB_ACK0 & ~n41122;
  assign n41124 = ~n15889 & ~n19767;
  assign n41125 = ~i_RtoB_ACK0 & ~n41124;
  assign n41126 = ~n41123 & ~n41125;
  assign n41127 = controllable_DEQ & ~n41126;
  assign n41128 = ~n19761 & ~n41127;
  assign n41129 = i_FULL & ~n41128;
  assign n41130 = ~n19769 & ~n41123;
  assign n41131 = controllable_DEQ & ~n41130;
  assign n41132 = ~n19779 & ~n41131;
  assign n41133 = ~i_FULL & ~n41132;
  assign n41134 = ~n41129 & ~n41133;
  assign n41135 = i_nEMPTY & ~n41134;
  assign n41136 = ~n15217 & ~n19787;
  assign n41137 = controllable_DEQ & ~n41136;
  assign n41138 = ~n19797 & ~n41137;
  assign n41139 = i_FULL & ~n41138;
  assign n41140 = ~n15245 & ~n19803;
  assign n41141 = controllable_DEQ & ~n41140;
  assign n41142 = ~n19813 & ~n41141;
  assign n41143 = ~i_FULL & ~n41142;
  assign n41144 = ~n41139 & ~n41143;
  assign n41145 = ~i_nEMPTY & ~n41144;
  assign n41146 = ~n41135 & ~n41145;
  assign n41147 = controllable_BtoS_ACK0 & ~n41146;
  assign n41148 = ~n16024 & ~n17690;
  assign n41149 = i_RtoB_ACK0 & ~n41148;
  assign n41150 = ~n16031 & ~n19841;
  assign n41151 = ~i_RtoB_ACK0 & ~n41150;
  assign n41152 = ~n41149 & ~n41151;
  assign n41153 = controllable_DEQ & ~n41152;
  assign n41154 = ~n19835 & ~n41153;
  assign n41155 = i_FULL & ~n41154;
  assign n41156 = ~n19843 & ~n41149;
  assign n41157 = controllable_DEQ & ~n41156;
  assign n41158 = ~n19853 & ~n41157;
  assign n41159 = ~i_FULL & ~n41158;
  assign n41160 = ~n41155 & ~n41159;
  assign n41161 = i_nEMPTY & ~n41160;
  assign n41162 = ~n17731 & ~n19861;
  assign n41163 = controllable_DEQ & ~n41162;
  assign n41164 = ~n19871 & ~n41163;
  assign n41165 = i_FULL & ~n41164;
  assign n41166 = ~n17764 & ~n19877;
  assign n41167 = controllable_DEQ & ~n41166;
  assign n41168 = ~n19887 & ~n41167;
  assign n41169 = ~i_FULL & ~n41168;
  assign n41170 = ~n41165 & ~n41169;
  assign n41171 = ~i_nEMPTY & ~n41170;
  assign n41172 = ~n41161 & ~n41171;
  assign n41173 = ~controllable_BtoS_ACK0 & ~n41172;
  assign n41174 = ~n41147 & ~n41173;
  assign n41175 = n4465 & ~n41174;
  assign n41176 = ~n16255 & ~n17690;
  assign n41177 = i_RtoB_ACK0 & ~n41176;
  assign n41178 = ~n16262 & ~n17701;
  assign n41179 = ~i_RtoB_ACK0 & ~n41178;
  assign n41180 = ~n41177 & ~n41179;
  assign n41181 = controllable_DEQ & ~n41180;
  assign n41182 = ~n19945 & ~n41181;
  assign n41183 = i_FULL & ~n41182;
  assign n41184 = ~n19949 & ~n41177;
  assign n41185 = controllable_DEQ & ~n41184;
  assign n41186 = ~n19959 & ~n41185;
  assign n41187 = ~i_FULL & ~n41186;
  assign n41188 = ~n41183 & ~n41187;
  assign n41189 = i_nEMPTY & ~n41188;
  assign n41190 = ~n17731 & ~n19965;
  assign n41191 = controllable_DEQ & ~n41190;
  assign n41192 = ~n19975 & ~n41191;
  assign n41193 = i_FULL & ~n41192;
  assign n41194 = ~n17764 & ~n19979;
  assign n41195 = controllable_DEQ & ~n41194;
  assign n41196 = ~n19989 & ~n41195;
  assign n41197 = ~i_FULL & ~n41196;
  assign n41198 = ~n41193 & ~n41197;
  assign n41199 = ~i_nEMPTY & ~n41198;
  assign n41200 = ~n41189 & ~n41199;
  assign n41201 = ~controllable_BtoS_ACK0 & ~n41200;
  assign n41202 = ~n19929 & ~n41201;
  assign n41203 = ~n4465 & ~n41202;
  assign n41204 = ~n41175 & ~n41203;
  assign n41205 = ~i_StoB_REQ10 & ~n41204;
  assign n41206 = ~n41121 & ~n41205;
  assign n41207 = controllable_BtoS_ACK10 & ~n41206;
  assign n41208 = ~n15882 & ~n17050;
  assign n41209 = i_RtoB_ACK0 & ~n41208;
  assign n41210 = ~n17622 & ~n20002;
  assign n41211 = ~i_RtoB_ACK0 & ~n41210;
  assign n41212 = ~n41209 & ~n41211;
  assign n41213 = controllable_DEQ & ~n41212;
  assign n41214 = ~n20019 & ~n41213;
  assign n41215 = i_FULL & ~n41214;
  assign n41216 = ~n20024 & ~n41209;
  assign n41217 = controllable_DEQ & ~n41216;
  assign n41218 = ~n20035 & ~n41217;
  assign n41219 = ~i_FULL & ~n41218;
  assign n41220 = ~n41215 & ~n41219;
  assign n41221 = i_nEMPTY & ~n41220;
  assign n41222 = ~n15604 & ~n20042;
  assign n41223 = controllable_DEQ & ~n41222;
  assign n41224 = ~n20053 & ~n41223;
  assign n41225 = i_FULL & ~n41224;
  assign n41226 = ~n15619 & ~n20058;
  assign n41227 = controllable_DEQ & ~n41226;
  assign n41228 = ~n20061 & ~n41227;
  assign n41229 = ~i_FULL & ~n41228;
  assign n41230 = ~n41225 & ~n41229;
  assign n41231 = ~i_nEMPTY & ~n41230;
  assign n41232 = ~n41221 & ~n41231;
  assign n41233 = controllable_BtoS_ACK0 & ~n41232;
  assign n41234 = ~n16024 & ~n18522;
  assign n41235 = i_RtoB_ACK0 & ~n41234;
  assign n41236 = ~n17701 & ~n20068;
  assign n41237 = ~i_RtoB_ACK0 & ~n41236;
  assign n41238 = ~n41235 & ~n41237;
  assign n41239 = controllable_DEQ & ~n41238;
  assign n41240 = ~n20077 & ~n41239;
  assign n41241 = i_FULL & ~n41240;
  assign n41242 = ~n20082 & ~n41235;
  assign n41243 = controllable_DEQ & ~n41242;
  assign n41244 = ~n20089 & ~n41243;
  assign n41245 = ~i_FULL & ~n41244;
  assign n41246 = ~n41241 & ~n41245;
  assign n41247 = i_nEMPTY & ~n41246;
  assign n41248 = ~n17925 & ~n20096;
  assign n41249 = controllable_DEQ & ~n41248;
  assign n41250 = ~n20103 & ~n41249;
  assign n41251 = i_FULL & ~n41250;
  assign n41252 = ~n17943 & ~n20108;
  assign n41253 = controllable_DEQ & ~n41252;
  assign n41254 = ~n20111 & ~n41253;
  assign n41255 = ~i_FULL & ~n41254;
  assign n41256 = ~n41251 & ~n41255;
  assign n41257 = ~i_nEMPTY & ~n41256;
  assign n41258 = ~n41247 & ~n41257;
  assign n41259 = ~controllable_BtoS_ACK0 & ~n41258;
  assign n41260 = ~n41233 & ~n41259;
  assign n41261 = n4465 & ~n41260;
  assign n41262 = ~n16255 & ~n18522;
  assign n41263 = i_RtoB_ACK0 & ~n41262;
  assign n41264 = ~n17701 & ~n20156;
  assign n41265 = ~i_RtoB_ACK0 & ~n41264;
  assign n41266 = ~n41263 & ~n41265;
  assign n41267 = controllable_DEQ & ~n41266;
  assign n41268 = ~n20165 & ~n41267;
  assign n41269 = i_FULL & ~n41268;
  assign n41270 = ~n20170 & ~n41263;
  assign n41271 = controllable_DEQ & ~n41270;
  assign n41272 = ~n20177 & ~n41271;
  assign n41273 = ~i_FULL & ~n41272;
  assign n41274 = ~n41269 & ~n41273;
  assign n41275 = i_nEMPTY & ~n41274;
  assign n41276 = ~n17925 & ~n20184;
  assign n41277 = controllable_DEQ & ~n41276;
  assign n41278 = ~n20191 & ~n41277;
  assign n41279 = i_FULL & ~n41278;
  assign n41280 = ~n17943 & ~n20196;
  assign n41281 = controllable_DEQ & ~n41280;
  assign n41282 = ~n20199 & ~n41281;
  assign n41283 = ~i_FULL & ~n41282;
  assign n41284 = ~n41279 & ~n41283;
  assign n41285 = ~i_nEMPTY & ~n41284;
  assign n41286 = ~n41275 & ~n41285;
  assign n41287 = ~controllable_BtoS_ACK0 & ~n41286;
  assign n41288 = ~n20155 & ~n41287;
  assign n41289 = ~n4465 & ~n41288;
  assign n41290 = ~n41261 & ~n41289;
  assign n41291 = i_StoB_REQ10 & ~n41290;
  assign n41292 = ~n41205 & ~n41291;
  assign n41293 = ~controllable_BtoS_ACK10 & ~n41292;
  assign n41294 = ~n41207 & ~n41293;
  assign n41295 = ~n4464 & ~n41294;
  assign n41296 = ~n41103 & ~n41295;
  assign n41297 = n4462 & ~n41296;
  assign n41298 = ~n17622 & ~n20366;
  assign n41299 = ~i_RtoB_ACK0 & ~n41298;
  assign n41300 = ~n18488 & ~n41299;
  assign n41301 = controllable_DEQ & ~n41300;
  assign n41302 = ~n20383 & ~n41301;
  assign n41303 = i_FULL & ~n41302;
  assign n41304 = ~n20401 & ~n41303;
  assign n41305 = i_nEMPTY & ~n41304;
  assign n41306 = ~n20429 & ~n41305;
  assign n41307 = controllable_BtoS_ACK0 & ~n41306;
  assign n41308 = ~n17701 & ~n20432;
  assign n41309 = ~i_RtoB_ACK0 & ~n41308;
  assign n41310 = ~n18524 & ~n41309;
  assign n41311 = controllable_DEQ & ~n41310;
  assign n41312 = ~n20441 & ~n41311;
  assign n41313 = i_FULL & ~n41312;
  assign n41314 = ~n20455 & ~n41313;
  assign n41315 = i_nEMPTY & ~n41314;
  assign n41316 = ~n20479 & ~n41315;
  assign n41317 = ~controllable_BtoS_ACK0 & ~n41316;
  assign n41318 = ~n41307 & ~n41317;
  assign n41319 = n4465 & ~n41318;
  assign n41320 = ~n19553 & ~n41317;
  assign n41321 = ~n4465 & ~n41320;
  assign n41322 = ~n41319 & ~n41321;
  assign n41323 = i_StoB_REQ10 & ~n41322;
  assign n41324 = ~n17622 & ~n17974;
  assign n41325 = ~i_RtoB_ACK0 & ~n41324;
  assign n41326 = ~n40709 & ~n41325;
  assign n41327 = controllable_DEQ & ~n41326;
  assign n41328 = ~n20495 & ~n41327;
  assign n41329 = i_FULL & ~n41328;
  assign n41330 = ~n20499 & ~n40709;
  assign n41331 = controllable_DEQ & ~n41330;
  assign n41332 = ~n20505 & ~n41331;
  assign n41333 = ~i_FULL & ~n41332;
  assign n41334 = ~n41329 & ~n41333;
  assign n41335 = i_nEMPTY & ~n41334;
  assign n41336 = ~n15217 & ~n20511;
  assign n41337 = controllable_DEQ & ~n41336;
  assign n41338 = ~n20517 & ~n41337;
  assign n41339 = i_FULL & ~n41338;
  assign n41340 = ~n15245 & ~n20521;
  assign n41341 = controllable_DEQ & ~n41340;
  assign n41342 = ~n20531 & ~n41341;
  assign n41343 = ~i_FULL & ~n41342;
  assign n41344 = ~n41339 & ~n41343;
  assign n41345 = ~i_nEMPTY & ~n41344;
  assign n41346 = ~n41335 & ~n41345;
  assign n41347 = controllable_BtoS_ACK0 & ~n41346;
  assign n41348 = ~n17701 & ~n18116;
  assign n41349 = ~i_RtoB_ACK0 & ~n41348;
  assign n41350 = ~n40801 & ~n41349;
  assign n41351 = controllable_DEQ & ~n41350;
  assign n41352 = ~n20545 & ~n41351;
  assign n41353 = i_FULL & ~n41352;
  assign n41354 = ~n20549 & ~n40801;
  assign n41355 = controllable_DEQ & ~n41354;
  assign n41356 = ~n20555 & ~n41355;
  assign n41357 = ~i_FULL & ~n41356;
  assign n41358 = ~n41353 & ~n41357;
  assign n41359 = i_nEMPTY & ~n41358;
  assign n41360 = ~n17731 & ~n20561;
  assign n41361 = controllable_DEQ & ~n41360;
  assign n41362 = ~n20567 & ~n41361;
  assign n41363 = i_FULL & ~n41362;
  assign n41364 = ~n17764 & ~n20571;
  assign n41365 = controllable_DEQ & ~n41364;
  assign n41366 = ~n20577 & ~n41365;
  assign n41367 = ~i_FULL & ~n41366;
  assign n41368 = ~n41363 & ~n41367;
  assign n41369 = ~i_nEMPTY & ~n41368;
  assign n41370 = ~n41359 & ~n41369;
  assign n41371 = ~controllable_BtoS_ACK0 & ~n41370;
  assign n41372 = ~n41347 & ~n41371;
  assign n41373 = n4465 & ~n41372;
  assign n41374 = ~n20619 & ~n40919;
  assign n41375 = ~n4465 & ~n41374;
  assign n41376 = ~n41373 & ~n41375;
  assign n41377 = ~i_StoB_REQ10 & ~n41376;
  assign n41378 = ~n41323 & ~n41377;
  assign n41379 = ~controllable_BtoS_ACK10 & ~n41378;
  assign n41380 = ~n20365 & ~n41379;
  assign n41381 = n4464 & ~n41380;
  assign n41382 = ~n17622 & ~n20680;
  assign n41383 = ~i_RtoB_ACK0 & ~n41382;
  assign n41384 = ~n18695 & ~n41383;
  assign n41385 = controllable_DEQ & ~n41384;
  assign n41386 = ~n20689 & ~n41385;
  assign n41387 = i_FULL & ~n41386;
  assign n41388 = ~n20703 & ~n41387;
  assign n41389 = i_nEMPTY & ~n41388;
  assign n41390 = ~n20727 & ~n41389;
  assign n41391 = controllable_BtoS_ACK0 & ~n41390;
  assign n41392 = ~n17701 & ~n20730;
  assign n41393 = ~i_RtoB_ACK0 & ~n41392;
  assign n41394 = ~n18726 & ~n41393;
  assign n41395 = controllable_DEQ & ~n41394;
  assign n41396 = ~n20739 & ~n41395;
  assign n41397 = i_FULL & ~n41396;
  assign n41398 = ~n20753 & ~n41397;
  assign n41399 = i_nEMPTY & ~n41398;
  assign n41400 = ~n20777 & ~n41399;
  assign n41401 = ~controllable_BtoS_ACK0 & ~n41400;
  assign n41402 = ~n41391 & ~n41401;
  assign n41403 = n4465 & ~n41402;
  assign n41404 = ~n20155 & ~n41401;
  assign n41405 = ~n4465 & ~n41404;
  assign n41406 = ~n41403 & ~n41405;
  assign n41407 = i_StoB_REQ10 & ~n41406;
  assign n41408 = ~n15889 & ~n17622;
  assign n41409 = ~i_RtoB_ACK0 & ~n41408;
  assign n41410 = ~n41123 & ~n41409;
  assign n41411 = controllable_DEQ & ~n41410;
  assign n41412 = ~n20793 & ~n41411;
  assign n41413 = i_FULL & ~n41412;
  assign n41414 = ~n20797 & ~n41123;
  assign n41415 = controllable_DEQ & ~n41414;
  assign n41416 = ~n20803 & ~n41415;
  assign n41417 = ~i_FULL & ~n41416;
  assign n41418 = ~n41413 & ~n41417;
  assign n41419 = i_nEMPTY & ~n41418;
  assign n41420 = ~n15217 & ~n20809;
  assign n41421 = controllable_DEQ & ~n41420;
  assign n41422 = ~n20815 & ~n41421;
  assign n41423 = i_FULL & ~n41422;
  assign n41424 = ~n15245 & ~n20819;
  assign n41425 = controllable_DEQ & ~n41424;
  assign n41426 = ~n20829 & ~n41425;
  assign n41427 = ~i_FULL & ~n41426;
  assign n41428 = ~n41423 & ~n41427;
  assign n41429 = ~i_nEMPTY & ~n41428;
  assign n41430 = ~n41419 & ~n41429;
  assign n41431 = controllable_BtoS_ACK0 & ~n41430;
  assign n41432 = ~n16031 & ~n17701;
  assign n41433 = ~i_RtoB_ACK0 & ~n41432;
  assign n41434 = ~n41149 & ~n41433;
  assign n41435 = controllable_DEQ & ~n41434;
  assign n41436 = ~n20843 & ~n41435;
  assign n41437 = i_FULL & ~n41436;
  assign n41438 = ~n20847 & ~n41149;
  assign n41439 = controllable_DEQ & ~n41438;
  assign n41440 = ~n20853 & ~n41439;
  assign n41441 = ~i_FULL & ~n41440;
  assign n41442 = ~n41437 & ~n41441;
  assign n41443 = i_nEMPTY & ~n41442;
  assign n41444 = ~n17731 & ~n20859;
  assign n41445 = controllable_DEQ & ~n41444;
  assign n41446 = ~n20865 & ~n41445;
  assign n41447 = i_FULL & ~n41446;
  assign n41448 = ~n17764 & ~n20869;
  assign n41449 = controllable_DEQ & ~n41448;
  assign n41450 = ~n20875 & ~n41449;
  assign n41451 = ~i_FULL & ~n41450;
  assign n41452 = ~n41447 & ~n41451;
  assign n41453 = ~i_nEMPTY & ~n41452;
  assign n41454 = ~n41443 & ~n41453;
  assign n41455 = ~controllable_BtoS_ACK0 & ~n41454;
  assign n41456 = ~n41431 & ~n41455;
  assign n41457 = n4465 & ~n41456;
  assign n41458 = ~n41203 & ~n41457;
  assign n41459 = ~i_StoB_REQ10 & ~n41458;
  assign n41460 = ~n41407 & ~n41459;
  assign n41461 = ~controllable_BtoS_ACK10 & ~n41460;
  assign n41462 = ~n20679 & ~n41461;
  assign n41463 = ~n4464 & ~n41462;
  assign n41464 = ~n41381 & ~n41463;
  assign n41465 = ~n4462 & ~n41464;
  assign n41466 = ~n41297 & ~n41465;
  assign n41467 = ~n4461 & ~n41466;
  assign n41468 = ~n40607 & ~n41467;
  assign n41469 = n4459 & ~n41468;
  assign n41470 = ~n39715 & ~n41469;
  assign n41471 = n4455 & ~n41470;
  assign n41472 = ~n23087 & ~n23399;
  assign n41473 = controllable_BtoS_ACK10 & ~n41472;
  assign n41474 = ~n36642 & ~n39722;
  assign n41475 = i_RtoB_ACK0 & ~n41474;
  assign n41476 = ~n36651 & ~n40928;
  assign n41477 = ~i_RtoB_ACK0 & ~n41476;
  assign n41478 = ~n41475 & ~n41477;
  assign n41479 = controllable_DEQ & ~n41478;
  assign n41480 = ~n36660 & ~n39731;
  assign n41481 = i_RtoB_ACK0 & ~n41480;
  assign n41482 = ~n11688 & ~n40933;
  assign n41483 = ~i_RtoB_ACK0 & ~n41482;
  assign n41484 = ~n41481 & ~n41483;
  assign n41485 = ~controllable_DEQ & ~n41484;
  assign n41486 = ~n41479 & ~n41485;
  assign n41487 = i_FULL & ~n41486;
  assign n41488 = ~n36642 & ~n39743;
  assign n41489 = i_RtoB_ACK0 & ~n41488;
  assign n41490 = ~n36672 & ~n40944;
  assign n41491 = ~i_RtoB_ACK0 & ~n41490;
  assign n41492 = ~n41489 & ~n41491;
  assign n41493 = controllable_DEQ & ~n41492;
  assign n41494 = ~n36660 & ~n39752;
  assign n41495 = i_RtoB_ACK0 & ~n41494;
  assign n41496 = ~n11714 & ~n40949;
  assign n41497 = ~i_RtoB_ACK0 & ~n41496;
  assign n41498 = ~n41495 & ~n41497;
  assign n41499 = ~controllable_DEQ & ~n41498;
  assign n41500 = ~n41493 & ~n41499;
  assign n41501 = ~i_FULL & ~n41500;
  assign n41502 = ~n41487 & ~n41501;
  assign n41503 = i_nEMPTY & ~n41502;
  assign n41504 = ~n36688 & ~n40962;
  assign n41505 = ~i_RtoB_ACK0 & ~n41504;
  assign n41506 = ~n39768 & ~n41505;
  assign n41507 = controllable_DEQ & ~n41506;
  assign n41508 = ~n36642 & ~n39775;
  assign n41509 = i_RtoB_ACK0 & ~n41508;
  assign n41510 = ~n11742 & ~n40967;
  assign n41511 = ~i_RtoB_ACK0 & ~n41510;
  assign n41512 = ~n41509 & ~n41511;
  assign n41513 = ~controllable_DEQ & ~n41512;
  assign n41514 = ~n41507 & ~n41513;
  assign n41515 = i_FULL & ~n41514;
  assign n41516 = ~n36698 & ~n40978;
  assign n41517 = ~i_RtoB_ACK0 & ~n41516;
  assign n41518 = ~n39789 & ~n41517;
  assign n41519 = controllable_DEQ & ~n41518;
  assign n41520 = ~controllable_DEQ & ~n41478;
  assign n41521 = ~n41519 & ~n41520;
  assign n41522 = ~i_FULL & ~n41521;
  assign n41523 = ~n41515 & ~n41522;
  assign n41524 = ~i_nEMPTY & ~n41523;
  assign n41525 = ~n41503 & ~n41524;
  assign n41526 = controllable_BtoS_ACK0 & ~n41525;
  assign n41527 = ~n36721 & ~n39804;
  assign n41528 = i_RtoB_ACK0 & ~n41527;
  assign n41529 = ~n36730 & ~n40999;
  assign n41530 = ~i_RtoB_ACK0 & ~n41529;
  assign n41531 = ~n41528 & ~n41530;
  assign n41532 = controllable_DEQ & ~n41531;
  assign n41533 = ~n36739 & ~n39813;
  assign n41534 = i_RtoB_ACK0 & ~n41533;
  assign n41535 = ~n11835 & ~n41004;
  assign n41536 = ~i_RtoB_ACK0 & ~n41535;
  assign n41537 = ~n41534 & ~n41536;
  assign n41538 = ~controllable_DEQ & ~n41537;
  assign n41539 = ~n41532 & ~n41538;
  assign n41540 = i_FULL & ~n41539;
  assign n41541 = ~n36721 & ~n39825;
  assign n41542 = i_RtoB_ACK0 & ~n41541;
  assign n41543 = ~n36751 & ~n41015;
  assign n41544 = ~i_RtoB_ACK0 & ~n41543;
  assign n41545 = ~n41542 & ~n41544;
  assign n41546 = controllable_DEQ & ~n41545;
  assign n41547 = ~n36739 & ~n39834;
  assign n41548 = i_RtoB_ACK0 & ~n41547;
  assign n41549 = ~n11861 & ~n41020;
  assign n41550 = ~i_RtoB_ACK0 & ~n41549;
  assign n41551 = ~n41548 & ~n41550;
  assign n41552 = ~controllable_DEQ & ~n41551;
  assign n41553 = ~n41546 & ~n41552;
  assign n41554 = ~i_FULL & ~n41553;
  assign n41555 = ~n41540 & ~n41554;
  assign n41556 = i_nEMPTY & ~n41555;
  assign n41557 = ~n36767 & ~n41033;
  assign n41558 = ~i_RtoB_ACK0 & ~n41557;
  assign n41559 = ~n39850 & ~n41558;
  assign n41560 = controllable_DEQ & ~n41559;
  assign n41561 = ~n36721 & ~n39857;
  assign n41562 = i_RtoB_ACK0 & ~n41561;
  assign n41563 = ~n11889 & ~n41038;
  assign n41564 = ~i_RtoB_ACK0 & ~n41563;
  assign n41565 = ~n41562 & ~n41564;
  assign n41566 = ~controllable_DEQ & ~n41565;
  assign n41567 = ~n41560 & ~n41566;
  assign n41568 = i_FULL & ~n41567;
  assign n41569 = ~n36777 & ~n41049;
  assign n41570 = ~i_RtoB_ACK0 & ~n41569;
  assign n41571 = ~n39871 & ~n41570;
  assign n41572 = controllable_DEQ & ~n41571;
  assign n41573 = ~controllable_DEQ & ~n41531;
  assign n41574 = ~n41572 & ~n41573;
  assign n41575 = ~i_FULL & ~n41574;
  assign n41576 = ~n41568 & ~n41575;
  assign n41577 = ~i_nEMPTY & ~n41576;
  assign n41578 = ~n41556 & ~n41577;
  assign n41579 = ~controllable_BtoS_ACK0 & ~n41578;
  assign n41580 = ~n41526 & ~n41579;
  assign n41581 = n4465 & ~n41580;
  assign n41582 = ~n21471 & ~n41581;
  assign n41583 = i_StoB_REQ10 & ~n41582;
  assign n41584 = ~n23399 & ~n41583;
  assign n41585 = ~controllable_BtoS_ACK10 & ~n41584;
  assign n41586 = ~n41473 & ~n41585;
  assign n41587 = n4464 & ~n41586;
  assign n41588 = ~n21981 & ~n41587;
  assign n41589 = n4463 & ~n41588;
  assign n41590 = ~n36883 & ~n39895;
  assign n41591 = i_RtoB_ACK0 & ~n41590;
  assign n41592 = ~n17562 & ~n36890;
  assign n41593 = ~i_RtoB_ACK0 & ~n41592;
  assign n41594 = ~n41591 & ~n41593;
  assign n41595 = ~controllable_DEQ & ~n41594;
  assign n41596 = ~n23529 & ~n41595;
  assign n41597 = i_FULL & ~n41596;
  assign n41598 = ~n17562 & ~n36903;
  assign n41599 = ~i_RtoB_ACK0 & ~n41598;
  assign n41600 = ~n41591 & ~n41599;
  assign n41601 = ~controllable_DEQ & ~n41600;
  assign n41602 = ~n23529 & ~n41601;
  assign n41603 = ~i_FULL & ~n41602;
  assign n41604 = ~n41597 & ~n41603;
  assign n41605 = i_nEMPTY & ~n41604;
  assign n41606 = ~n36918 & ~n39905;
  assign n41607 = i_RtoB_ACK0 & ~n41606;
  assign n41608 = ~n17581 & ~n36925;
  assign n41609 = ~i_RtoB_ACK0 & ~n41608;
  assign n41610 = ~n41607 & ~n41609;
  assign n41611 = ~controllable_DEQ & ~n41610;
  assign n41612 = ~n23541 & ~n41611;
  assign n41613 = i_FULL & ~n41612;
  assign n41614 = ~n17545 & ~n37044;
  assign n41615 = ~i_RtoB_ACK0 & ~n41614;
  assign n41616 = ~n41607 & ~n41615;
  assign n41617 = ~controllable_DEQ & ~n41616;
  assign n41618 = ~n23551 & ~n41617;
  assign n41619 = ~i_FULL & ~n41618;
  assign n41620 = ~n41613 & ~n41619;
  assign n41621 = ~i_nEMPTY & ~n41620;
  assign n41622 = ~n41605 & ~n41621;
  assign n41623 = controllable_BtoS_ACK0 & ~n41622;
  assign n41624 = ~n37064 & ~n39923;
  assign n41625 = i_RtoB_ACK0 & ~n41624;
  assign n41626 = ~n14841 & ~n37071;
  assign n41627 = ~i_RtoB_ACK0 & ~n41626;
  assign n41628 = ~n41625 & ~n41627;
  assign n41629 = ~controllable_DEQ & ~n41628;
  assign n41630 = ~n23567 & ~n41629;
  assign n41631 = i_FULL & ~n41630;
  assign n41632 = ~n14841 & ~n37084;
  assign n41633 = ~i_RtoB_ACK0 & ~n41632;
  assign n41634 = ~n41625 & ~n41633;
  assign n41635 = ~controllable_DEQ & ~n41634;
  assign n41636 = ~n23567 & ~n41635;
  assign n41637 = ~i_FULL & ~n41636;
  assign n41638 = ~n41631 & ~n41637;
  assign n41639 = i_nEMPTY & ~n41638;
  assign n41640 = ~n37099 & ~n39933;
  assign n41641 = i_RtoB_ACK0 & ~n41640;
  assign n41642 = ~n14860 & ~n37106;
  assign n41643 = ~i_RtoB_ACK0 & ~n41642;
  assign n41644 = ~n41641 & ~n41643;
  assign n41645 = ~controllable_DEQ & ~n41644;
  assign n41646 = ~n23579 & ~n41645;
  assign n41647 = i_FULL & ~n41646;
  assign n41648 = ~n14824 & ~n37130;
  assign n41649 = ~i_RtoB_ACK0 & ~n41648;
  assign n41650 = ~n41641 & ~n41649;
  assign n41651 = ~controllable_DEQ & ~n41650;
  assign n41652 = ~n23589 & ~n41651;
  assign n41653 = ~i_FULL & ~n41652;
  assign n41654 = ~n41647 & ~n41653;
  assign n41655 = ~i_nEMPTY & ~n41654;
  assign n41656 = ~n41639 & ~n41655;
  assign n41657 = ~controllable_BtoS_ACK0 & ~n41656;
  assign n41658 = ~n41623 & ~n41657;
  assign n41659 = n4465 & ~n41658;
  assign n41660 = ~n22097 & ~n22103;
  assign n41661 = i_FULL & ~n41660;
  assign n41662 = ~n22109 & ~n41661;
  assign n41663 = i_nEMPTY & ~n41662;
  assign n41664 = ~n22133 & ~n41663;
  assign n41665 = ~controllable_BtoS_ACK0 & ~n41664;
  assign n41666 = ~n21013 & ~n41665;
  assign n41667 = ~n4465 & ~n41666;
  assign n41668 = ~n41659 & ~n41667;
  assign n41669 = i_StoB_REQ10 & ~n41668;
  assign n41670 = ~n37252 & ~n39956;
  assign n41671 = i_RtoB_ACK0 & ~n41670;
  assign n41672 = ~n17974 & ~n37263;
  assign n41673 = ~i_RtoB_ACK0 & ~n41672;
  assign n41674 = ~n41671 & ~n41673;
  assign n41675 = controllable_DEQ & ~n41674;
  assign n41676 = ~n37460 & ~n39964;
  assign n41677 = i_RtoB_ACK0 & ~n41676;
  assign n41678 = ~n17993 & ~n37472;
  assign n41679 = ~i_RtoB_ACK0 & ~n41678;
  assign n41680 = ~n41677 & ~n41679;
  assign n41681 = ~controllable_DEQ & ~n41680;
  assign n41682 = ~n41675 & ~n41681;
  assign n41683 = i_FULL & ~n41682;
  assign n41684 = ~n18012 & ~n37482;
  assign n41685 = ~i_RtoB_ACK0 & ~n41684;
  assign n41686 = ~n41671 & ~n41685;
  assign n41687 = controllable_DEQ & ~n41686;
  assign n41688 = ~n18028 & ~n37495;
  assign n41689 = ~i_RtoB_ACK0 & ~n41688;
  assign n41690 = ~n41677 & ~n41689;
  assign n41691 = ~controllable_DEQ & ~n41690;
  assign n41692 = ~n41687 & ~n41691;
  assign n41693 = ~i_FULL & ~n41692;
  assign n41694 = ~n41683 & ~n41693;
  assign n41695 = i_nEMPTY & ~n41694;
  assign n41696 = ~n18049 & ~n37511;
  assign n41697 = ~i_RtoB_ACK0 & ~n41696;
  assign n41698 = ~n39985 & ~n41697;
  assign n41699 = controllable_DEQ & ~n41698;
  assign n41700 = ~n37522 & ~n39991;
  assign n41701 = i_RtoB_ACK0 & ~n41700;
  assign n41702 = ~n18065 & ~n37531;
  assign n41703 = ~i_RtoB_ACK0 & ~n41702;
  assign n41704 = ~n41701 & ~n41703;
  assign n41705 = ~controllable_DEQ & ~n41704;
  assign n41706 = ~n41699 & ~n41705;
  assign n41707 = i_FULL & ~n41706;
  assign n41708 = ~n18084 & ~n37544;
  assign n41709 = ~i_RtoB_ACK0 & ~n41708;
  assign n41710 = ~n40004 & ~n41709;
  assign n41711 = controllable_DEQ & ~n41710;
  assign n41712 = ~n37522 & ~n40011;
  assign n41713 = i_RtoB_ACK0 & ~n41712;
  assign n41714 = ~n17974 & ~n37668;
  assign n41715 = ~i_RtoB_ACK0 & ~n41714;
  assign n41716 = ~n41713 & ~n41715;
  assign n41717 = ~controllable_DEQ & ~n41716;
  assign n41718 = ~n41711 & ~n41717;
  assign n41719 = ~i_FULL & ~n41718;
  assign n41720 = ~n41707 & ~n41719;
  assign n41721 = ~i_nEMPTY & ~n41720;
  assign n41722 = ~n41695 & ~n41721;
  assign n41723 = controllable_BtoS_ACK0 & ~n41722;
  assign n41724 = ~n37694 & ~n40026;
  assign n41725 = i_RtoB_ACK0 & ~n41724;
  assign n41726 = ~n18116 & ~n37705;
  assign n41727 = ~i_RtoB_ACK0 & ~n41726;
  assign n41728 = ~n41725 & ~n41727;
  assign n41729 = controllable_DEQ & ~n41728;
  assign n41730 = ~n37723 & ~n40034;
  assign n41731 = i_RtoB_ACK0 & ~n41730;
  assign n41732 = ~n18135 & ~n37735;
  assign n41733 = ~i_RtoB_ACK0 & ~n41732;
  assign n41734 = ~n41731 & ~n41733;
  assign n41735 = ~controllable_DEQ & ~n41734;
  assign n41736 = ~n41729 & ~n41735;
  assign n41737 = i_FULL & ~n41736;
  assign n41738 = ~n18154 & ~n37745;
  assign n41739 = ~i_RtoB_ACK0 & ~n41738;
  assign n41740 = ~n41725 & ~n41739;
  assign n41741 = controllable_DEQ & ~n41740;
  assign n41742 = ~n18170 & ~n37758;
  assign n41743 = ~i_RtoB_ACK0 & ~n41742;
  assign n41744 = ~n41731 & ~n41743;
  assign n41745 = ~controllable_DEQ & ~n41744;
  assign n41746 = ~n41741 & ~n41745;
  assign n41747 = ~i_FULL & ~n41746;
  assign n41748 = ~n41737 & ~n41747;
  assign n41749 = i_nEMPTY & ~n41748;
  assign n41750 = ~n18191 & ~n37774;
  assign n41751 = ~i_RtoB_ACK0 & ~n41750;
  assign n41752 = ~n40055 & ~n41751;
  assign n41753 = controllable_DEQ & ~n41752;
  assign n41754 = ~n37785 & ~n40061;
  assign n41755 = i_RtoB_ACK0 & ~n41754;
  assign n41756 = ~n18207 & ~n37794;
  assign n41757 = ~i_RtoB_ACK0 & ~n41756;
  assign n41758 = ~n41755 & ~n41757;
  assign n41759 = ~controllable_DEQ & ~n41758;
  assign n41760 = ~n41753 & ~n41759;
  assign n41761 = i_FULL & ~n41760;
  assign n41762 = ~n18226 & ~n37807;
  assign n41763 = ~i_RtoB_ACK0 & ~n41762;
  assign n41764 = ~n40074 & ~n41763;
  assign n41765 = controllable_DEQ & ~n41764;
  assign n41766 = ~n37785 & ~n40081;
  assign n41767 = i_RtoB_ACK0 & ~n41766;
  assign n41768 = ~n18116 & ~n37830;
  assign n41769 = ~i_RtoB_ACK0 & ~n41768;
  assign n41770 = ~n41767 & ~n41769;
  assign n41771 = ~controllable_DEQ & ~n41770;
  assign n41772 = ~n41765 & ~n41771;
  assign n41773 = ~i_FULL & ~n41772;
  assign n41774 = ~n41761 & ~n41773;
  assign n41775 = ~i_nEMPTY & ~n41774;
  assign n41776 = ~n41749 & ~n41775;
  assign n41777 = ~controllable_BtoS_ACK0 & ~n41776;
  assign n41778 = ~n41723 & ~n41777;
  assign n41779 = n4465 & ~n41778;
  assign n41780 = ~n37846 & ~n40097;
  assign n41781 = i_RtoB_ACK0 & ~n41780;
  assign n41782 = ~n15281 & ~n37852;
  assign n41783 = ~i_RtoB_ACK0 & ~n41782;
  assign n41784 = ~n41781 & ~n41783;
  assign n41785 = controllable_DEQ & ~n41784;
  assign n41786 = ~n22297 & ~n41785;
  assign n41787 = i_FULL & ~n41786;
  assign n41788 = ~n15319 & ~n37862;
  assign n41789 = ~i_RtoB_ACK0 & ~n41788;
  assign n41790 = ~n41781 & ~n41789;
  assign n41791 = controllable_DEQ & ~n41790;
  assign n41792 = ~n22307 & ~n41791;
  assign n41793 = ~i_FULL & ~n41792;
  assign n41794 = ~n41787 & ~n41793;
  assign n41795 = i_nEMPTY & ~n41794;
  assign n41796 = ~n15356 & ~n37874;
  assign n41797 = ~i_RtoB_ACK0 & ~n41796;
  assign n41798 = ~n17731 & ~n41797;
  assign n41799 = controllable_DEQ & ~n41798;
  assign n41800 = ~n22321 & ~n41799;
  assign n41801 = i_FULL & ~n41800;
  assign n41802 = ~n15391 & ~n37884;
  assign n41803 = ~i_RtoB_ACK0 & ~n41802;
  assign n41804 = ~n17764 & ~n41803;
  assign n41805 = controllable_DEQ & ~n41804;
  assign n41806 = ~n22331 & ~n41805;
  assign n41807 = ~i_FULL & ~n41806;
  assign n41808 = ~n41801 & ~n41807;
  assign n41809 = ~i_nEMPTY & ~n41808;
  assign n41810 = ~n41795 & ~n41809;
  assign n41811 = ~controllable_BtoS_ACK0 & ~n41810;
  assign n41812 = ~n22285 & ~n41811;
  assign n41813 = ~n4465 & ~n41812;
  assign n41814 = ~n41779 & ~n41813;
  assign n41815 = ~i_StoB_REQ10 & ~n41814;
  assign n41816 = ~n41669 & ~n41815;
  assign n41817 = controllable_BtoS_ACK10 & ~n41816;
  assign n41818 = ~n37904 & ~n40132;
  assign n41819 = i_RtoB_ACK0 & ~n41818;
  assign n41820 = ~n37910 & ~n40928;
  assign n41821 = ~i_RtoB_ACK0 & ~n41820;
  assign n41822 = ~n41819 & ~n41821;
  assign n41823 = controllable_DEQ & ~n41822;
  assign n41824 = ~n37919 & ~n40140;
  assign n41825 = i_RtoB_ACK0 & ~n41824;
  assign n41826 = ~n37472 & ~n40933;
  assign n41827 = ~i_RtoB_ACK0 & ~n41826;
  assign n41828 = ~n41825 & ~n41827;
  assign n41829 = ~controllable_DEQ & ~n41828;
  assign n41830 = ~n41823 & ~n41829;
  assign n41831 = i_FULL & ~n41830;
  assign n41832 = ~n37929 & ~n40944;
  assign n41833 = ~i_RtoB_ACK0 & ~n41832;
  assign n41834 = ~n41819 & ~n41833;
  assign n41835 = controllable_DEQ & ~n41834;
  assign n41836 = ~n37495 & ~n40949;
  assign n41837 = ~i_RtoB_ACK0 & ~n41836;
  assign n41838 = ~n41825 & ~n41837;
  assign n41839 = ~controllable_DEQ & ~n41838;
  assign n41840 = ~n41835 & ~n41839;
  assign n41841 = ~i_FULL & ~n41840;
  assign n41842 = ~n41831 & ~n41841;
  assign n41843 = i_nEMPTY & ~n41842;
  assign n41844 = ~n37943 & ~n40962;
  assign n41845 = ~i_RtoB_ACK0 & ~n41844;
  assign n41846 = ~n40157 & ~n41845;
  assign n41847 = controllable_DEQ & ~n41846;
  assign n41848 = ~n37952 & ~n40163;
  assign n41849 = i_RtoB_ACK0 & ~n41848;
  assign n41850 = ~n37531 & ~n40967;
  assign n41851 = ~i_RtoB_ACK0 & ~n41850;
  assign n41852 = ~n41849 & ~n41851;
  assign n41853 = ~controllable_DEQ & ~n41852;
  assign n41854 = ~n41847 & ~n41853;
  assign n41855 = i_FULL & ~n41854;
  assign n41856 = ~n37962 & ~n40978;
  assign n41857 = ~i_RtoB_ACK0 & ~n41856;
  assign n41858 = ~n40171 & ~n41857;
  assign n41859 = controllable_DEQ & ~n41858;
  assign n41860 = ~n37952 & ~n40178;
  assign n41861 = i_RtoB_ACK0 & ~n41860;
  assign n41862 = ~n37974 & ~n40928;
  assign n41863 = ~i_RtoB_ACK0 & ~n41862;
  assign n41864 = ~n41861 & ~n41863;
  assign n41865 = ~controllable_DEQ & ~n41864;
  assign n41866 = ~n41859 & ~n41865;
  assign n41867 = ~i_FULL & ~n41866;
  assign n41868 = ~n41855 & ~n41867;
  assign n41869 = ~i_nEMPTY & ~n41868;
  assign n41870 = ~n41843 & ~n41869;
  assign n41871 = controllable_BtoS_ACK0 & ~n41870;
  assign n41872 = ~n37988 & ~n40193;
  assign n41873 = i_RtoB_ACK0 & ~n41872;
  assign n41874 = ~n37994 & ~n40999;
  assign n41875 = ~i_RtoB_ACK0 & ~n41874;
  assign n41876 = ~n41873 & ~n41875;
  assign n41877 = controllable_DEQ & ~n41876;
  assign n41878 = ~n38003 & ~n40201;
  assign n41879 = i_RtoB_ACK0 & ~n41878;
  assign n41880 = ~n37735 & ~n41004;
  assign n41881 = ~i_RtoB_ACK0 & ~n41880;
  assign n41882 = ~n41879 & ~n41881;
  assign n41883 = ~controllable_DEQ & ~n41882;
  assign n41884 = ~n41877 & ~n41883;
  assign n41885 = i_FULL & ~n41884;
  assign n41886 = ~n38013 & ~n41015;
  assign n41887 = ~i_RtoB_ACK0 & ~n41886;
  assign n41888 = ~n41873 & ~n41887;
  assign n41889 = controllable_DEQ & ~n41888;
  assign n41890 = ~n37758 & ~n41020;
  assign n41891 = ~i_RtoB_ACK0 & ~n41890;
  assign n41892 = ~n41879 & ~n41891;
  assign n41893 = ~controllable_DEQ & ~n41892;
  assign n41894 = ~n41889 & ~n41893;
  assign n41895 = ~i_FULL & ~n41894;
  assign n41896 = ~n41885 & ~n41895;
  assign n41897 = i_nEMPTY & ~n41896;
  assign n41898 = ~n38027 & ~n41033;
  assign n41899 = ~i_RtoB_ACK0 & ~n41898;
  assign n41900 = ~n40218 & ~n41899;
  assign n41901 = controllable_DEQ & ~n41900;
  assign n41902 = ~n38036 & ~n40224;
  assign n41903 = i_RtoB_ACK0 & ~n41902;
  assign n41904 = ~n37794 & ~n41038;
  assign n41905 = ~i_RtoB_ACK0 & ~n41904;
  assign n41906 = ~n41903 & ~n41905;
  assign n41907 = ~controllable_DEQ & ~n41906;
  assign n41908 = ~n41901 & ~n41907;
  assign n41909 = i_FULL & ~n41908;
  assign n41910 = ~n38046 & ~n41049;
  assign n41911 = ~i_RtoB_ACK0 & ~n41910;
  assign n41912 = ~n40232 & ~n41911;
  assign n41913 = controllable_DEQ & ~n41912;
  assign n41914 = ~n38036 & ~n40239;
  assign n41915 = i_RtoB_ACK0 & ~n41914;
  assign n41916 = ~n38058 & ~n40999;
  assign n41917 = ~i_RtoB_ACK0 & ~n41916;
  assign n41918 = ~n41915 & ~n41917;
  assign n41919 = ~controllable_DEQ & ~n41918;
  assign n41920 = ~n41913 & ~n41919;
  assign n41921 = ~i_FULL & ~n41920;
  assign n41922 = ~n41909 & ~n41921;
  assign n41923 = ~i_nEMPTY & ~n41922;
  assign n41924 = ~n41897 & ~n41923;
  assign n41925 = ~controllable_BtoS_ACK0 & ~n41924;
  assign n41926 = ~n41871 & ~n41925;
  assign n41927 = n4465 & ~n41926;
  assign n41928 = ~n38074 & ~n40255;
  assign n41929 = i_RtoB_ACK0 & ~n41928;
  assign n41930 = ~n19554 & ~n38080;
  assign n41931 = ~i_RtoB_ACK0 & ~n41930;
  assign n41932 = ~n41929 & ~n41931;
  assign n41933 = controllable_DEQ & ~n41932;
  assign n41934 = ~n22492 & ~n41933;
  assign n41935 = i_FULL & ~n41934;
  assign n41936 = ~n19566 & ~n38090;
  assign n41937 = ~i_RtoB_ACK0 & ~n41936;
  assign n41938 = ~n41929 & ~n41937;
  assign n41939 = controllable_DEQ & ~n41938;
  assign n41940 = ~n22502 & ~n41939;
  assign n41941 = ~i_FULL & ~n41940;
  assign n41942 = ~n41935 & ~n41941;
  assign n41943 = i_nEMPTY & ~n41942;
  assign n41944 = ~n19580 & ~n38102;
  assign n41945 = ~i_RtoB_ACK0 & ~n41944;
  assign n41946 = ~n17925 & ~n41945;
  assign n41947 = controllable_DEQ & ~n41946;
  assign n41948 = ~n22516 & ~n41947;
  assign n41949 = i_FULL & ~n41948;
  assign n41950 = ~n19592 & ~n38112;
  assign n41951 = ~i_RtoB_ACK0 & ~n41950;
  assign n41952 = ~n17943 & ~n41951;
  assign n41953 = controllable_DEQ & ~n41952;
  assign n41954 = ~n22523 & ~n41953;
  assign n41955 = ~i_FULL & ~n41954;
  assign n41956 = ~n41949 & ~n41955;
  assign n41957 = ~i_nEMPTY & ~n41956;
  assign n41958 = ~n41943 & ~n41957;
  assign n41959 = ~controllable_BtoS_ACK0 & ~n41958;
  assign n41960 = ~n22480 & ~n41959;
  assign n41961 = ~n4465 & ~n41960;
  assign n41962 = ~n41927 & ~n41961;
  assign n41963 = i_StoB_REQ10 & ~n41962;
  assign n41964 = ~n41815 & ~n41963;
  assign n41965 = ~controllable_BtoS_ACK10 & ~n41964;
  assign n41966 = ~n41817 & ~n41965;
  assign n41967 = n4464 & ~n41966;
  assign n41968 = ~n22549 & ~n22555;
  assign n41969 = i_FULL & ~n41968;
  assign n41970 = ~n22561 & ~n41969;
  assign n41971 = i_nEMPTY & ~n41970;
  assign n41972 = ~n22585 & ~n41971;
  assign n41973 = controllable_BtoS_ACK0 & ~n41972;
  assign n41974 = ~n22599 & ~n22605;
  assign n41975 = i_FULL & ~n41974;
  assign n41976 = ~n22611 & ~n41975;
  assign n41977 = i_nEMPTY & ~n41976;
  assign n41978 = ~n22635 & ~n41977;
  assign n41979 = ~controllable_BtoS_ACK0 & ~n41978;
  assign n41980 = ~n41973 & ~n41979;
  assign n41981 = n4465 & ~n41980;
  assign n41982 = ~n21013 & ~n41979;
  assign n41983 = ~n4465 & ~n41982;
  assign n41984 = ~n41981 & ~n41983;
  assign n41985 = i_StoB_REQ10 & ~n41984;
  assign n41986 = ~n38152 & ~n40292;
  assign n41987 = i_RtoB_ACK0 & ~n41986;
  assign n41988 = ~n15889 & ~n38158;
  assign n41989 = ~i_RtoB_ACK0 & ~n41988;
  assign n41990 = ~n41987 & ~n41989;
  assign n41991 = controllable_DEQ & ~n41990;
  assign n41992 = ~n22655 & ~n41991;
  assign n41993 = i_FULL & ~n41992;
  assign n41994 = ~n15927 & ~n38168;
  assign n41995 = ~i_RtoB_ACK0 & ~n41994;
  assign n41996 = ~n41987 & ~n41995;
  assign n41997 = controllable_DEQ & ~n41996;
  assign n41998 = ~n22665 & ~n41997;
  assign n41999 = ~i_FULL & ~n41998;
  assign n42000 = ~n41993 & ~n41999;
  assign n42001 = i_nEMPTY & ~n42000;
  assign n42002 = ~n15964 & ~n38180;
  assign n42003 = ~i_RtoB_ACK0 & ~n42002;
  assign n42004 = ~n15217 & ~n42003;
  assign n42005 = controllable_DEQ & ~n42004;
  assign n42006 = ~n22679 & ~n42005;
  assign n42007 = i_FULL & ~n42006;
  assign n42008 = ~n15999 & ~n38190;
  assign n42009 = ~i_RtoB_ACK0 & ~n42008;
  assign n42010 = ~n15245 & ~n42009;
  assign n42011 = controllable_DEQ & ~n42010;
  assign n42012 = ~n22689 & ~n42011;
  assign n42013 = ~i_FULL & ~n42012;
  assign n42014 = ~n42007 & ~n42013;
  assign n42015 = ~i_nEMPTY & ~n42014;
  assign n42016 = ~n42001 & ~n42015;
  assign n42017 = controllable_BtoS_ACK0 & ~n42016;
  assign n42018 = ~n38204 & ~n40321;
  assign n42019 = i_RtoB_ACK0 & ~n42018;
  assign n42020 = ~n16031 & ~n38210;
  assign n42021 = ~i_RtoB_ACK0 & ~n42020;
  assign n42022 = ~n42019 & ~n42021;
  assign n42023 = controllable_DEQ & ~n42022;
  assign n42024 = ~n22707 & ~n42023;
  assign n42025 = i_FULL & ~n42024;
  assign n42026 = ~n16069 & ~n38220;
  assign n42027 = ~i_RtoB_ACK0 & ~n42026;
  assign n42028 = ~n42019 & ~n42027;
  assign n42029 = controllable_DEQ & ~n42028;
  assign n42030 = ~n22717 & ~n42029;
  assign n42031 = ~i_FULL & ~n42030;
  assign n42032 = ~n42025 & ~n42031;
  assign n42033 = i_nEMPTY & ~n42032;
  assign n42034 = ~n16106 & ~n38232;
  assign n42035 = ~i_RtoB_ACK0 & ~n42034;
  assign n42036 = ~n17731 & ~n42035;
  assign n42037 = controllable_DEQ & ~n42036;
  assign n42038 = ~n22731 & ~n42037;
  assign n42039 = i_FULL & ~n42038;
  assign n42040 = ~n16141 & ~n38242;
  assign n42041 = ~i_RtoB_ACK0 & ~n42040;
  assign n42042 = ~n17764 & ~n42041;
  assign n42043 = controllable_DEQ & ~n42042;
  assign n42044 = ~n22741 & ~n42043;
  assign n42045 = ~i_FULL & ~n42044;
  assign n42046 = ~n42039 & ~n42045;
  assign n42047 = ~i_nEMPTY & ~n42046;
  assign n42048 = ~n42033 & ~n42047;
  assign n42049 = ~controllable_BtoS_ACK0 & ~n42048;
  assign n42050 = ~n42017 & ~n42049;
  assign n42051 = n4465 & ~n42050;
  assign n42052 = ~n38258 & ~n40351;
  assign n42053 = i_RtoB_ACK0 & ~n42052;
  assign n42054 = ~n16262 & ~n38264;
  assign n42055 = ~i_RtoB_ACK0 & ~n42054;
  assign n42056 = ~n42053 & ~n42055;
  assign n42057 = controllable_DEQ & ~n42056;
  assign n42058 = ~n22801 & ~n42057;
  assign n42059 = i_FULL & ~n42058;
  assign n42060 = ~n16300 & ~n38274;
  assign n42061 = ~i_RtoB_ACK0 & ~n42060;
  assign n42062 = ~n42053 & ~n42061;
  assign n42063 = controllable_DEQ & ~n42062;
  assign n42064 = ~n22811 & ~n42063;
  assign n42065 = ~i_FULL & ~n42064;
  assign n42066 = ~n42059 & ~n42065;
  assign n42067 = i_nEMPTY & ~n42066;
  assign n42068 = ~n16337 & ~n38286;
  assign n42069 = ~i_RtoB_ACK0 & ~n42068;
  assign n42070 = ~n17731 & ~n42069;
  assign n42071 = controllable_DEQ & ~n42070;
  assign n42072 = ~n22825 & ~n42071;
  assign n42073 = i_FULL & ~n42072;
  assign n42074 = ~n16372 & ~n38296;
  assign n42075 = ~i_RtoB_ACK0 & ~n42074;
  assign n42076 = ~n17764 & ~n42075;
  assign n42077 = controllable_DEQ & ~n42076;
  assign n42078 = ~n22835 & ~n42077;
  assign n42079 = ~i_FULL & ~n42078;
  assign n42080 = ~n42073 & ~n42079;
  assign n42081 = ~i_nEMPTY & ~n42080;
  assign n42082 = ~n42067 & ~n42081;
  assign n42083 = ~controllable_BtoS_ACK0 & ~n42082;
  assign n42084 = ~n22789 & ~n42083;
  assign n42085 = ~n4465 & ~n42084;
  assign n42086 = ~n42051 & ~n42085;
  assign n42087 = ~i_StoB_REQ10 & ~n42086;
  assign n42088 = ~n41985 & ~n42087;
  assign n42089 = controllable_BtoS_ACK10 & ~n42088;
  assign n42090 = ~n38316 & ~n40385;
  assign n42091 = i_RtoB_ACK0 & ~n42090;
  assign n42092 = ~n20002 & ~n38322;
  assign n42093 = ~i_RtoB_ACK0 & ~n42092;
  assign n42094 = ~n42091 & ~n42093;
  assign n42095 = controllable_DEQ & ~n42094;
  assign n42096 = ~n22859 & ~n42095;
  assign n42097 = i_FULL & ~n42096;
  assign n42098 = ~n20022 & ~n38332;
  assign n42099 = ~i_RtoB_ACK0 & ~n42098;
  assign n42100 = ~n42091 & ~n42099;
  assign n42101 = controllable_DEQ & ~n42100;
  assign n42102 = ~n22869 & ~n42101;
  assign n42103 = ~i_FULL & ~n42102;
  assign n42104 = ~n42097 & ~n42103;
  assign n42105 = i_nEMPTY & ~n42104;
  assign n42106 = ~n20040 & ~n38344;
  assign n42107 = ~i_RtoB_ACK0 & ~n42106;
  assign n42108 = ~n15604 & ~n42107;
  assign n42109 = controllable_DEQ & ~n42108;
  assign n42110 = ~n22883 & ~n42109;
  assign n42111 = i_FULL & ~n42110;
  assign n42112 = ~n20056 & ~n38354;
  assign n42113 = ~i_RtoB_ACK0 & ~n42112;
  assign n42114 = ~n15619 & ~n42113;
  assign n42115 = controllable_DEQ & ~n42114;
  assign n42116 = ~n22890 & ~n42115;
  assign n42117 = ~i_FULL & ~n42116;
  assign n42118 = ~n42111 & ~n42117;
  assign n42119 = ~i_nEMPTY & ~n42118;
  assign n42120 = ~n42105 & ~n42119;
  assign n42121 = controllable_BtoS_ACK0 & ~n42120;
  assign n42122 = ~n38368 & ~n40413;
  assign n42123 = i_RtoB_ACK0 & ~n42122;
  assign n42124 = ~n20068 & ~n38374;
  assign n42125 = ~i_RtoB_ACK0 & ~n42124;
  assign n42126 = ~n42123 & ~n42125;
  assign n42127 = controllable_DEQ & ~n42126;
  assign n42128 = ~n22908 & ~n42127;
  assign n42129 = i_FULL & ~n42128;
  assign n42130 = ~n20080 & ~n38384;
  assign n42131 = ~i_RtoB_ACK0 & ~n42130;
  assign n42132 = ~n42123 & ~n42131;
  assign n42133 = controllable_DEQ & ~n42132;
  assign n42134 = ~n22918 & ~n42133;
  assign n42135 = ~i_FULL & ~n42134;
  assign n42136 = ~n42129 & ~n42135;
  assign n42137 = i_nEMPTY & ~n42136;
  assign n42138 = ~n20094 & ~n38396;
  assign n42139 = ~i_RtoB_ACK0 & ~n42138;
  assign n42140 = ~n17925 & ~n42139;
  assign n42141 = controllable_DEQ & ~n42140;
  assign n42142 = ~n22932 & ~n42141;
  assign n42143 = i_FULL & ~n42142;
  assign n42144 = ~n20106 & ~n38406;
  assign n42145 = ~i_RtoB_ACK0 & ~n42144;
  assign n42146 = ~n17943 & ~n42145;
  assign n42147 = controllable_DEQ & ~n42146;
  assign n42148 = ~n22939 & ~n42147;
  assign n42149 = ~i_FULL & ~n42148;
  assign n42150 = ~n42143 & ~n42149;
  assign n42151 = ~i_nEMPTY & ~n42150;
  assign n42152 = ~n42137 & ~n42151;
  assign n42153 = ~controllable_BtoS_ACK0 & ~n42152;
  assign n42154 = ~n42121 & ~n42153;
  assign n42155 = n4465 & ~n42154;
  assign n42156 = ~n38422 & ~n40443;
  assign n42157 = i_RtoB_ACK0 & ~n42156;
  assign n42158 = ~n20156 & ~n38428;
  assign n42159 = ~i_RtoB_ACK0 & ~n42158;
  assign n42160 = ~n42157 & ~n42159;
  assign n42161 = controllable_DEQ & ~n42160;
  assign n42162 = ~n22996 & ~n42161;
  assign n42163 = i_FULL & ~n42162;
  assign n42164 = ~n20168 & ~n38438;
  assign n42165 = ~i_RtoB_ACK0 & ~n42164;
  assign n42166 = ~n42157 & ~n42165;
  assign n42167 = controllable_DEQ & ~n42166;
  assign n42168 = ~n23006 & ~n42167;
  assign n42169 = ~i_FULL & ~n42168;
  assign n42170 = ~n42163 & ~n42169;
  assign n42171 = i_nEMPTY & ~n42170;
  assign n42172 = ~n20182 & ~n38450;
  assign n42173 = ~i_RtoB_ACK0 & ~n42172;
  assign n42174 = ~n17925 & ~n42173;
  assign n42175 = controllable_DEQ & ~n42174;
  assign n42176 = ~n23020 & ~n42175;
  assign n42177 = i_FULL & ~n42176;
  assign n42178 = ~n20194 & ~n38460;
  assign n42179 = ~i_RtoB_ACK0 & ~n42178;
  assign n42180 = ~n17943 & ~n42179;
  assign n42181 = controllable_DEQ & ~n42180;
  assign n42182 = ~n23027 & ~n42181;
  assign n42183 = ~i_FULL & ~n42182;
  assign n42184 = ~n42177 & ~n42183;
  assign n42185 = ~i_nEMPTY & ~n42184;
  assign n42186 = ~n42171 & ~n42185;
  assign n42187 = ~controllable_BtoS_ACK0 & ~n42186;
  assign n42188 = ~n22984 & ~n42187;
  assign n42189 = ~n4465 & ~n42188;
  assign n42190 = ~n42155 & ~n42189;
  assign n42191 = i_StoB_REQ10 & ~n42190;
  assign n42192 = ~n42087 & ~n42191;
  assign n42193 = ~controllable_BtoS_ACK10 & ~n42192;
  assign n42194 = ~n42089 & ~n42193;
  assign n42195 = ~n4464 & ~n42194;
  assign n42196 = ~n41967 & ~n42195;
  assign n42197 = ~n4463 & ~n42196;
  assign n42198 = ~n41589 & ~n42197;
  assign n42199 = n4462 & ~n42198;
  assign n42200 = ~n20366 & ~n38484;
  assign n42201 = ~i_RtoB_ACK0 & ~n42200;
  assign n42202 = ~n23625 & ~n42201;
  assign n42203 = controllable_DEQ & ~n42202;
  assign n42204 = ~n23635 & ~n42203;
  assign n42205 = i_FULL & ~n42204;
  assign n42206 = ~n23647 & ~n42205;
  assign n42207 = i_nEMPTY & ~n42206;
  assign n42208 = ~n23670 & ~n42207;
  assign n42209 = controllable_BtoS_ACK0 & ~n42208;
  assign n42210 = ~n20432 & ~n38496;
  assign n42211 = ~i_RtoB_ACK0 & ~n42210;
  assign n42212 = ~n23674 & ~n42211;
  assign n42213 = controllable_DEQ & ~n42212;
  assign n42214 = ~n23684 & ~n42213;
  assign n42215 = i_FULL & ~n42214;
  assign n42216 = ~n23696 & ~n42215;
  assign n42217 = i_nEMPTY & ~n42216;
  assign n42218 = ~n23719 & ~n42217;
  assign n42219 = ~controllable_BtoS_ACK0 & ~n42218;
  assign n42220 = ~n42209 & ~n42219;
  assign n42221 = n4465 & ~n42220;
  assign n42222 = ~n22480 & ~n42219;
  assign n42223 = ~n4465 & ~n42222;
  assign n42224 = ~n42221 & ~n42223;
  assign n42225 = i_StoB_REQ10 & ~n42224;
  assign n42226 = ~n38514 & ~n40483;
  assign n42227 = i_RtoB_ACK0 & ~n42226;
  assign n42228 = ~n17974 & ~n38518;
  assign n42229 = ~i_RtoB_ACK0 & ~n42228;
  assign n42230 = ~n42227 & ~n42229;
  assign n42231 = controllable_DEQ & ~n42230;
  assign n42232 = ~n23739 & ~n42231;
  assign n42233 = i_FULL & ~n42232;
  assign n42234 = ~n18012 & ~n38526;
  assign n42235 = ~i_RtoB_ACK0 & ~n42234;
  assign n42236 = ~n42227 & ~n42235;
  assign n42237 = controllable_DEQ & ~n42236;
  assign n42238 = ~n23749 & ~n42237;
  assign n42239 = ~i_FULL & ~n42238;
  assign n42240 = ~n42233 & ~n42239;
  assign n42241 = i_nEMPTY & ~n42240;
  assign n42242 = ~n18049 & ~n38536;
  assign n42243 = ~i_RtoB_ACK0 & ~n42242;
  assign n42244 = ~n15217 & ~n42243;
  assign n42245 = controllable_DEQ & ~n42244;
  assign n42246 = ~n23763 & ~n42245;
  assign n42247 = i_FULL & ~n42246;
  assign n42248 = ~n18084 & ~n38544;
  assign n42249 = ~i_RtoB_ACK0 & ~n42248;
  assign n42250 = ~n15245 & ~n42249;
  assign n42251 = controllable_DEQ & ~n42250;
  assign n42252 = ~n23773 & ~n42251;
  assign n42253 = ~i_FULL & ~n42252;
  assign n42254 = ~n42247 & ~n42253;
  assign n42255 = ~i_nEMPTY & ~n42254;
  assign n42256 = ~n42241 & ~n42255;
  assign n42257 = controllable_BtoS_ACK0 & ~n42256;
  assign n42258 = ~n38556 & ~n40511;
  assign n42259 = i_RtoB_ACK0 & ~n42258;
  assign n42260 = ~n18116 & ~n38560;
  assign n42261 = ~i_RtoB_ACK0 & ~n42260;
  assign n42262 = ~n42259 & ~n42261;
  assign n42263 = controllable_DEQ & ~n42262;
  assign n42264 = ~n23791 & ~n42263;
  assign n42265 = i_FULL & ~n42264;
  assign n42266 = ~n18154 & ~n38568;
  assign n42267 = ~i_RtoB_ACK0 & ~n42266;
  assign n42268 = ~n42259 & ~n42267;
  assign n42269 = controllable_DEQ & ~n42268;
  assign n42270 = ~n23801 & ~n42269;
  assign n42271 = ~i_FULL & ~n42270;
  assign n42272 = ~n42265 & ~n42271;
  assign n42273 = i_nEMPTY & ~n42272;
  assign n42274 = ~n18191 & ~n38578;
  assign n42275 = ~i_RtoB_ACK0 & ~n42274;
  assign n42276 = ~n17731 & ~n42275;
  assign n42277 = controllable_DEQ & ~n42276;
  assign n42278 = ~n23815 & ~n42277;
  assign n42279 = i_FULL & ~n42278;
  assign n42280 = ~n18226 & ~n38586;
  assign n42281 = ~i_RtoB_ACK0 & ~n42280;
  assign n42282 = ~n17764 & ~n42281;
  assign n42283 = controllable_DEQ & ~n42282;
  assign n42284 = ~n23825 & ~n42283;
  assign n42285 = ~i_FULL & ~n42284;
  assign n42286 = ~n42279 & ~n42285;
  assign n42287 = ~i_nEMPTY & ~n42286;
  assign n42288 = ~n42273 & ~n42287;
  assign n42289 = ~controllable_BtoS_ACK0 & ~n42288;
  assign n42290 = ~n42257 & ~n42289;
  assign n42291 = n4465 & ~n42290;
  assign n42292 = ~n23867 & ~n41811;
  assign n42293 = ~n4465 & ~n42292;
  assign n42294 = ~n42291 & ~n42293;
  assign n42295 = ~i_StoB_REQ10 & ~n42294;
  assign n42296 = ~n42225 & ~n42295;
  assign n42297 = ~controllable_BtoS_ACK10 & ~n42296;
  assign n42298 = ~n23623 & ~n42297;
  assign n42299 = n4464 & ~n42298;
  assign n42300 = ~n20680 & ~n38608;
  assign n42301 = ~i_RtoB_ACK0 & ~n42300;
  assign n42302 = ~n23929 & ~n42301;
  assign n42303 = controllable_DEQ & ~n42302;
  assign n42304 = ~n23939 & ~n42303;
  assign n42305 = i_FULL & ~n42304;
  assign n42306 = ~n23951 & ~n42305;
  assign n42307 = i_nEMPTY & ~n42306;
  assign n42308 = ~n23974 & ~n42307;
  assign n42309 = controllable_BtoS_ACK0 & ~n42308;
  assign n42310 = ~n20730 & ~n38620;
  assign n42311 = ~i_RtoB_ACK0 & ~n42310;
  assign n42312 = ~n23978 & ~n42311;
  assign n42313 = controllable_DEQ & ~n42312;
  assign n42314 = ~n23988 & ~n42313;
  assign n42315 = i_FULL & ~n42314;
  assign n42316 = ~n24000 & ~n42315;
  assign n42317 = i_nEMPTY & ~n42316;
  assign n42318 = ~n24023 & ~n42317;
  assign n42319 = ~controllable_BtoS_ACK0 & ~n42318;
  assign n42320 = ~n42309 & ~n42319;
  assign n42321 = n4465 & ~n42320;
  assign n42322 = ~n22984 & ~n42319;
  assign n42323 = ~n4465 & ~n42322;
  assign n42324 = ~n42321 & ~n42323;
  assign n42325 = i_StoB_REQ10 & ~n42324;
  assign n42326 = ~n38638 & ~n40549;
  assign n42327 = i_RtoB_ACK0 & ~n42326;
  assign n42328 = ~n15889 & ~n38642;
  assign n42329 = ~i_RtoB_ACK0 & ~n42328;
  assign n42330 = ~n42327 & ~n42329;
  assign n42331 = controllable_DEQ & ~n42330;
  assign n42332 = ~n24041 & ~n42331;
  assign n42333 = i_FULL & ~n42332;
  assign n42334 = ~n15927 & ~n38650;
  assign n42335 = ~i_RtoB_ACK0 & ~n42334;
  assign n42336 = ~n42327 & ~n42335;
  assign n42337 = controllable_DEQ & ~n42336;
  assign n42338 = ~n24049 & ~n42337;
  assign n42339 = ~i_FULL & ~n42338;
  assign n42340 = ~n42333 & ~n42339;
  assign n42341 = i_nEMPTY & ~n42340;
  assign n42342 = ~n15964 & ~n38660;
  assign n42343 = ~i_RtoB_ACK0 & ~n42342;
  assign n42344 = ~n15217 & ~n42343;
  assign n42345 = controllable_DEQ & ~n42344;
  assign n42346 = ~n24061 & ~n42345;
  assign n42347 = i_FULL & ~n42346;
  assign n42348 = ~n15999 & ~n38668;
  assign n42349 = ~i_RtoB_ACK0 & ~n42348;
  assign n42350 = ~n15245 & ~n42349;
  assign n42351 = controllable_DEQ & ~n42350;
  assign n42352 = ~n24069 & ~n42351;
  assign n42353 = ~i_FULL & ~n42352;
  assign n42354 = ~n42347 & ~n42353;
  assign n42355 = ~i_nEMPTY & ~n42354;
  assign n42356 = ~n42341 & ~n42355;
  assign n42357 = controllable_BtoS_ACK0 & ~n42356;
  assign n42358 = ~n38680 & ~n40573;
  assign n42359 = i_RtoB_ACK0 & ~n42358;
  assign n42360 = ~n16031 & ~n38684;
  assign n42361 = ~i_RtoB_ACK0 & ~n42360;
  assign n42362 = ~n42359 & ~n42361;
  assign n42363 = controllable_DEQ & ~n42362;
  assign n42364 = ~n24085 & ~n42363;
  assign n42365 = i_FULL & ~n42364;
  assign n42366 = ~n16069 & ~n38692;
  assign n42367 = ~i_RtoB_ACK0 & ~n42366;
  assign n42368 = ~n42359 & ~n42367;
  assign n42369 = controllable_DEQ & ~n42368;
  assign n42370 = ~n24093 & ~n42369;
  assign n42371 = ~i_FULL & ~n42370;
  assign n42372 = ~n42365 & ~n42371;
  assign n42373 = i_nEMPTY & ~n42372;
  assign n42374 = ~n16106 & ~n38702;
  assign n42375 = ~i_RtoB_ACK0 & ~n42374;
  assign n42376 = ~n17731 & ~n42375;
  assign n42377 = controllable_DEQ & ~n42376;
  assign n42378 = ~n24105 & ~n42377;
  assign n42379 = i_FULL & ~n42378;
  assign n42380 = ~n16141 & ~n38710;
  assign n42381 = ~i_RtoB_ACK0 & ~n42380;
  assign n42382 = ~n17764 & ~n42381;
  assign n42383 = controllable_DEQ & ~n42382;
  assign n42384 = ~n24113 & ~n42383;
  assign n42385 = ~i_FULL & ~n42384;
  assign n42386 = ~n42379 & ~n42385;
  assign n42387 = ~i_nEMPTY & ~n42386;
  assign n42388 = ~n42373 & ~n42387;
  assign n42389 = ~controllable_BtoS_ACK0 & ~n42388;
  assign n42390 = ~n42357 & ~n42389;
  assign n42391 = n4465 & ~n42390;
  assign n42392 = ~n42085 & ~n42391;
  assign n42393 = ~i_StoB_REQ10 & ~n42392;
  assign n42394 = ~n42325 & ~n42393;
  assign n42395 = ~controllable_BtoS_ACK10 & ~n42394;
  assign n42396 = ~n23927 & ~n42395;
  assign n42397 = ~n4464 & ~n42396;
  assign n42398 = ~n42299 & ~n42397;
  assign n42399 = ~n4463 & ~n42398;
  assign n42400 = ~n23523 & ~n42399;
  assign n42401 = ~n4462 & ~n42400;
  assign n42402 = ~n42199 & ~n42401;
  assign n42403 = n4461 & ~n42402;
  assign n42404 = ~n11170 & ~n39895;
  assign n42405 = i_RtoB_ACK0 & ~n42404;
  assign n42406 = ~n41593 & ~n42405;
  assign n42407 = ~controllable_DEQ & ~n42406;
  assign n42408 = ~n25129 & ~n42407;
  assign n42409 = i_nEMPTY & ~n42408;
  assign n42410 = ~n11147 & ~n39905;
  assign n42411 = i_RtoB_ACK0 & ~n42410;
  assign n42412 = ~n41609 & ~n42411;
  assign n42413 = ~controllable_DEQ & ~n42412;
  assign n42414 = ~n23063 & ~n42413;
  assign n42415 = i_FULL & ~n42414;
  assign n42416 = ~n17545 & ~n38744;
  assign n42417 = ~i_RtoB_ACK0 & ~n42416;
  assign n42418 = ~n42411 & ~n42417;
  assign n42419 = ~controllable_DEQ & ~n42418;
  assign n42420 = ~n23073 & ~n42419;
  assign n42421 = ~i_FULL & ~n42420;
  assign n42422 = ~n42415 & ~n42421;
  assign n42423 = ~i_nEMPTY & ~n42422;
  assign n42424 = ~n42409 & ~n42423;
  assign n42425 = controllable_BtoS_ACK0 & ~n42424;
  assign n42426 = ~n5363 & ~n39923;
  assign n42427 = i_RtoB_ACK0 & ~n42426;
  assign n42428 = ~n41627 & ~n42427;
  assign n42429 = ~controllable_DEQ & ~n42428;
  assign n42430 = ~n25157 & ~n42429;
  assign n42431 = i_nEMPTY & ~n42430;
  assign n42432 = ~n5340 & ~n39933;
  assign n42433 = i_RtoB_ACK0 & ~n42432;
  assign n42434 = ~n41643 & ~n42433;
  assign n42435 = ~controllable_DEQ & ~n42434;
  assign n42436 = ~n21031 & ~n42435;
  assign n42437 = i_FULL & ~n42436;
  assign n42438 = ~n14824 & ~n38764;
  assign n42439 = ~i_RtoB_ACK0 & ~n42438;
  assign n42440 = ~n42433 & ~n42439;
  assign n42441 = ~controllable_DEQ & ~n42440;
  assign n42442 = ~n21041 & ~n42441;
  assign n42443 = ~i_FULL & ~n42442;
  assign n42444 = ~n42437 & ~n42443;
  assign n42445 = ~i_nEMPTY & ~n42444;
  assign n42446 = ~n42431 & ~n42445;
  assign n42447 = ~controllable_BtoS_ACK0 & ~n42446;
  assign n42448 = ~n42425 & ~n42447;
  assign n42449 = n4465 & ~n42448;
  assign n42450 = ~n24215 & ~n42449;
  assign n42451 = i_StoB_REQ10 & ~n42450;
  assign n42452 = ~n11652 & ~n17280;
  assign n42453 = i_RtoB_ACK0 & ~n42452;
  assign n42454 = ~n17974 & ~n38883;
  assign n42455 = ~i_RtoB_ACK0 & ~n42454;
  assign n42456 = ~n42453 & ~n42455;
  assign n42457 = controllable_DEQ & ~n42456;
  assign n42458 = ~n11681 & ~n40722;
  assign n42459 = i_RtoB_ACK0 & ~n42458;
  assign n42460 = ~n17993 & ~n38892;
  assign n42461 = ~i_RtoB_ACK0 & ~n42460;
  assign n42462 = ~n42459 & ~n42461;
  assign n42463 = ~controllable_DEQ & ~n42462;
  assign n42464 = ~n42457 & ~n42463;
  assign n42465 = i_FULL & ~n42464;
  assign n42466 = ~n18012 & ~n38902;
  assign n42467 = ~i_RtoB_ACK0 & ~n42466;
  assign n42468 = ~n42453 & ~n42467;
  assign n42469 = controllable_DEQ & ~n42468;
  assign n42470 = ~n18028 & ~n38910;
  assign n42471 = ~i_RtoB_ACK0 & ~n42470;
  assign n42472 = ~n42459 & ~n42471;
  assign n42473 = ~controllable_DEQ & ~n42472;
  assign n42474 = ~n42469 & ~n42473;
  assign n42475 = ~i_FULL & ~n42474;
  assign n42476 = ~n42465 & ~n42475;
  assign n42477 = i_nEMPTY & ~n42476;
  assign n42478 = ~n18049 & ~n38924;
  assign n42479 = ~i_RtoB_ACK0 & ~n42478;
  assign n42480 = ~n15217 & ~n42479;
  assign n42481 = controllable_DEQ & ~n42480;
  assign n42482 = ~n11652 & ~n40760;
  assign n42483 = i_RtoB_ACK0 & ~n42482;
  assign n42484 = ~n18065 & ~n38933;
  assign n42485 = ~i_RtoB_ACK0 & ~n42484;
  assign n42486 = ~n42483 & ~n42485;
  assign n42487 = ~controllable_DEQ & ~n42486;
  assign n42488 = ~n42481 & ~n42487;
  assign n42489 = i_FULL & ~n42488;
  assign n42490 = ~n18084 & ~n38944;
  assign n42491 = ~i_RtoB_ACK0 & ~n42490;
  assign n42492 = ~n15245 & ~n42491;
  assign n42493 = controllable_DEQ & ~n42492;
  assign n42494 = ~n11652 & ~n40783;
  assign n42495 = i_RtoB_ACK0 & ~n42494;
  assign n42496 = ~n17974 & ~n38954;
  assign n42497 = ~i_RtoB_ACK0 & ~n42496;
  assign n42498 = ~n42495 & ~n42497;
  assign n42499 = ~controllable_DEQ & ~n42498;
  assign n42500 = ~n42493 & ~n42499;
  assign n42501 = ~i_FULL & ~n42500;
  assign n42502 = ~n42489 & ~n42501;
  assign n42503 = ~i_nEMPTY & ~n42502;
  assign n42504 = ~n42477 & ~n42503;
  assign n42505 = controllable_BtoS_ACK0 & ~n42504;
  assign n42506 = ~n11799 & ~n17690;
  assign n42507 = i_RtoB_ACK0 & ~n42506;
  assign n42508 = ~n18116 & ~n38978;
  assign n42509 = ~i_RtoB_ACK0 & ~n42508;
  assign n42510 = ~n42507 & ~n42509;
  assign n42511 = controllable_DEQ & ~n42510;
  assign n42512 = ~n11828 & ~n40814;
  assign n42513 = i_RtoB_ACK0 & ~n42512;
  assign n42514 = ~n18135 & ~n38987;
  assign n42515 = ~i_RtoB_ACK0 & ~n42514;
  assign n42516 = ~n42513 & ~n42515;
  assign n42517 = ~controllable_DEQ & ~n42516;
  assign n42518 = ~n42511 & ~n42517;
  assign n42519 = i_FULL & ~n42518;
  assign n42520 = ~n18154 & ~n38997;
  assign n42521 = ~i_RtoB_ACK0 & ~n42520;
  assign n42522 = ~n42507 & ~n42521;
  assign n42523 = controllable_DEQ & ~n42522;
  assign n42524 = ~n18170 & ~n39005;
  assign n42525 = ~i_RtoB_ACK0 & ~n42524;
  assign n42526 = ~n42513 & ~n42525;
  assign n42527 = ~controllable_DEQ & ~n42526;
  assign n42528 = ~n42523 & ~n42527;
  assign n42529 = ~i_FULL & ~n42528;
  assign n42530 = ~n42519 & ~n42529;
  assign n42531 = i_nEMPTY & ~n42530;
  assign n42532 = ~n18191 & ~n39019;
  assign n42533 = ~i_RtoB_ACK0 & ~n42532;
  assign n42534 = ~n17731 & ~n42533;
  assign n42535 = controllable_DEQ & ~n42534;
  assign n42536 = ~n11799 & ~n40852;
  assign n42537 = i_RtoB_ACK0 & ~n42536;
  assign n42538 = ~n18207 & ~n39028;
  assign n42539 = ~i_RtoB_ACK0 & ~n42538;
  assign n42540 = ~n42537 & ~n42539;
  assign n42541 = ~controllable_DEQ & ~n42540;
  assign n42542 = ~n42535 & ~n42541;
  assign n42543 = i_FULL & ~n42542;
  assign n42544 = ~n18226 & ~n39039;
  assign n42545 = ~i_RtoB_ACK0 & ~n42544;
  assign n42546 = ~n17764 & ~n42545;
  assign n42547 = controllable_DEQ & ~n42546;
  assign n42548 = ~n11799 & ~n40875;
  assign n42549 = i_RtoB_ACK0 & ~n42548;
  assign n42550 = ~n18116 & ~n39049;
  assign n42551 = ~i_RtoB_ACK0 & ~n42550;
  assign n42552 = ~n42549 & ~n42551;
  assign n42553 = ~controllable_DEQ & ~n42552;
  assign n42554 = ~n42547 & ~n42553;
  assign n42555 = ~i_FULL & ~n42554;
  assign n42556 = ~n42543 & ~n42555;
  assign n42557 = ~i_nEMPTY & ~n42556;
  assign n42558 = ~n42531 & ~n42557;
  assign n42559 = ~controllable_BtoS_ACK0 & ~n42558;
  assign n42560 = ~n42505 & ~n42559;
  assign n42561 = n4465 & ~n42560;
  assign n42562 = ~n7244 & ~n17690;
  assign n42563 = i_RtoB_ACK0 & ~n42562;
  assign n42564 = ~n15281 & ~n39063;
  assign n42565 = ~i_RtoB_ACK0 & ~n42564;
  assign n42566 = ~n42563 & ~n42565;
  assign n42567 = controllable_DEQ & ~n42566;
  assign n42568 = ~n24351 & ~n42567;
  assign n42569 = i_FULL & ~n42568;
  assign n42570 = ~n15319 & ~n39071;
  assign n42571 = ~i_RtoB_ACK0 & ~n42570;
  assign n42572 = ~n42563 & ~n42571;
  assign n42573 = controllable_DEQ & ~n42572;
  assign n42574 = ~n24361 & ~n42573;
  assign n42575 = ~i_FULL & ~n42574;
  assign n42576 = ~n42569 & ~n42575;
  assign n42577 = i_nEMPTY & ~n42576;
  assign n42578 = ~n15356 & ~n39081;
  assign n42579 = ~i_RtoB_ACK0 & ~n42578;
  assign n42580 = ~n17731 & ~n42579;
  assign n42581 = controllable_DEQ & ~n42580;
  assign n42582 = ~n24371 & ~n42581;
  assign n42583 = i_FULL & ~n42582;
  assign n42584 = ~n15391 & ~n39089;
  assign n42585 = ~i_RtoB_ACK0 & ~n42584;
  assign n42586 = ~n17764 & ~n42585;
  assign n42587 = controllable_DEQ & ~n42586;
  assign n42588 = ~n24377 & ~n42587;
  assign n42589 = ~i_FULL & ~n42588;
  assign n42590 = ~n42583 & ~n42589;
  assign n42591 = ~i_nEMPTY & ~n42590;
  assign n42592 = ~n42577 & ~n42591;
  assign n42593 = ~controllable_BtoS_ACK0 & ~n42592;
  assign n42594 = ~n24339 & ~n42593;
  assign n42595 = ~n4465 & ~n42594;
  assign n42596 = ~n42561 & ~n42595;
  assign n42597 = ~i_StoB_REQ10 & ~n42596;
  assign n42598 = ~n42451 & ~n42597;
  assign n42599 = controllable_BtoS_ACK10 & ~n42598;
  assign n42600 = ~n17050 & ~n36642;
  assign n42601 = i_RtoB_ACK0 & ~n42600;
  assign n42602 = ~n39111 & ~n40928;
  assign n42603 = ~i_RtoB_ACK0 & ~n42602;
  assign n42604 = ~n42601 & ~n42603;
  assign n42605 = controllable_DEQ & ~n42604;
  assign n42606 = ~n36660 & ~n40140;
  assign n42607 = i_RtoB_ACK0 & ~n42606;
  assign n42608 = ~n39117 & ~n40933;
  assign n42609 = ~i_RtoB_ACK0 & ~n42608;
  assign n42610 = ~n42607 & ~n42609;
  assign n42611 = ~controllable_DEQ & ~n42610;
  assign n42612 = ~n42605 & ~n42611;
  assign n42613 = i_FULL & ~n42612;
  assign n42614 = ~n39127 & ~n40944;
  assign n42615 = ~i_RtoB_ACK0 & ~n42614;
  assign n42616 = ~n42601 & ~n42615;
  assign n42617 = controllable_DEQ & ~n42616;
  assign n42618 = ~n39133 & ~n40949;
  assign n42619 = ~i_RtoB_ACK0 & ~n42618;
  assign n42620 = ~n42607 & ~n42619;
  assign n42621 = ~controllable_DEQ & ~n42620;
  assign n42622 = ~n42617 & ~n42621;
  assign n42623 = ~i_FULL & ~n42622;
  assign n42624 = ~n42613 & ~n42623;
  assign n42625 = i_nEMPTY & ~n42624;
  assign n42626 = ~n39146 & ~n40962;
  assign n42627 = ~i_RtoB_ACK0 & ~n42626;
  assign n42628 = ~n15604 & ~n42627;
  assign n42629 = controllable_DEQ & ~n42628;
  assign n42630 = ~n36642 & ~n40163;
  assign n42631 = i_RtoB_ACK0 & ~n42630;
  assign n42632 = ~n39152 & ~n40967;
  assign n42633 = ~i_RtoB_ACK0 & ~n42632;
  assign n42634 = ~n42631 & ~n42633;
  assign n42635 = ~controllable_DEQ & ~n42634;
  assign n42636 = ~n42629 & ~n42635;
  assign n42637 = i_FULL & ~n42636;
  assign n42638 = ~n39162 & ~n40978;
  assign n42639 = ~i_RtoB_ACK0 & ~n42638;
  assign n42640 = ~n15619 & ~n42639;
  assign n42641 = controllable_DEQ & ~n42640;
  assign n42642 = ~n36642 & ~n40178;
  assign n42643 = i_RtoB_ACK0 & ~n42642;
  assign n42644 = ~n39168 & ~n40928;
  assign n42645 = ~i_RtoB_ACK0 & ~n42644;
  assign n42646 = ~n42643 & ~n42645;
  assign n42647 = ~controllable_DEQ & ~n42646;
  assign n42648 = ~n42641 & ~n42647;
  assign n42649 = ~i_FULL & ~n42648;
  assign n42650 = ~n42637 & ~n42649;
  assign n42651 = ~i_nEMPTY & ~n42650;
  assign n42652 = ~n42625 & ~n42651;
  assign n42653 = controllable_BtoS_ACK0 & ~n42652;
  assign n42654 = ~n18522 & ~n36721;
  assign n42655 = i_RtoB_ACK0 & ~n42654;
  assign n42656 = ~n39184 & ~n40999;
  assign n42657 = ~i_RtoB_ACK0 & ~n42656;
  assign n42658 = ~n42655 & ~n42657;
  assign n42659 = controllable_DEQ & ~n42658;
  assign n42660 = ~n36739 & ~n40201;
  assign n42661 = i_RtoB_ACK0 & ~n42660;
  assign n42662 = ~n39190 & ~n41004;
  assign n42663 = ~i_RtoB_ACK0 & ~n42662;
  assign n42664 = ~n42661 & ~n42663;
  assign n42665 = ~controllable_DEQ & ~n42664;
  assign n42666 = ~n42659 & ~n42665;
  assign n42667 = i_FULL & ~n42666;
  assign n42668 = ~n39200 & ~n41015;
  assign n42669 = ~i_RtoB_ACK0 & ~n42668;
  assign n42670 = ~n42655 & ~n42669;
  assign n42671 = controllable_DEQ & ~n42670;
  assign n42672 = ~n39206 & ~n41020;
  assign n42673 = ~i_RtoB_ACK0 & ~n42672;
  assign n42674 = ~n42661 & ~n42673;
  assign n42675 = ~controllable_DEQ & ~n42674;
  assign n42676 = ~n42671 & ~n42675;
  assign n42677 = ~i_FULL & ~n42676;
  assign n42678 = ~n42667 & ~n42677;
  assign n42679 = i_nEMPTY & ~n42678;
  assign n42680 = ~n39219 & ~n41033;
  assign n42681 = ~i_RtoB_ACK0 & ~n42680;
  assign n42682 = ~n17925 & ~n42681;
  assign n42683 = controllable_DEQ & ~n42682;
  assign n42684 = ~n36721 & ~n40224;
  assign n42685 = i_RtoB_ACK0 & ~n42684;
  assign n42686 = ~n39225 & ~n41038;
  assign n42687 = ~i_RtoB_ACK0 & ~n42686;
  assign n42688 = ~n42685 & ~n42687;
  assign n42689 = ~controllable_DEQ & ~n42688;
  assign n42690 = ~n42683 & ~n42689;
  assign n42691 = i_FULL & ~n42690;
  assign n42692 = ~n39235 & ~n41049;
  assign n42693 = ~i_RtoB_ACK0 & ~n42692;
  assign n42694 = ~n17943 & ~n42693;
  assign n42695 = controllable_DEQ & ~n42694;
  assign n42696 = ~n36721 & ~n40239;
  assign n42697 = i_RtoB_ACK0 & ~n42696;
  assign n42698 = ~n39241 & ~n40999;
  assign n42699 = ~i_RtoB_ACK0 & ~n42698;
  assign n42700 = ~n42697 & ~n42699;
  assign n42701 = ~controllable_DEQ & ~n42700;
  assign n42702 = ~n42695 & ~n42701;
  assign n42703 = ~i_FULL & ~n42702;
  assign n42704 = ~n42691 & ~n42703;
  assign n42705 = ~i_nEMPTY & ~n42704;
  assign n42706 = ~n42679 & ~n42705;
  assign n42707 = ~controllable_BtoS_ACK0 & ~n42706;
  assign n42708 = ~n42653 & ~n42707;
  assign n42709 = n4465 & ~n42708;
  assign n42710 = ~n7612 & ~n18522;
  assign n42711 = i_RtoB_ACK0 & ~n42710;
  assign n42712 = ~n19554 & ~n39255;
  assign n42713 = ~i_RtoB_ACK0 & ~n42712;
  assign n42714 = ~n42711 & ~n42713;
  assign n42715 = controllable_DEQ & ~n42714;
  assign n42716 = ~n24514 & ~n42715;
  assign n42717 = i_FULL & ~n42716;
  assign n42718 = ~n19566 & ~n39263;
  assign n42719 = ~i_RtoB_ACK0 & ~n42718;
  assign n42720 = ~n42711 & ~n42719;
  assign n42721 = controllable_DEQ & ~n42720;
  assign n42722 = ~n24524 & ~n42721;
  assign n42723 = ~i_FULL & ~n42722;
  assign n42724 = ~n42717 & ~n42723;
  assign n42725 = i_nEMPTY & ~n42724;
  assign n42726 = ~n19580 & ~n39273;
  assign n42727 = ~i_RtoB_ACK0 & ~n42726;
  assign n42728 = ~n17925 & ~n42727;
  assign n42729 = controllable_DEQ & ~n42728;
  assign n42730 = ~n24534 & ~n42729;
  assign n42731 = i_FULL & ~n42730;
  assign n42732 = ~n19592 & ~n39281;
  assign n42733 = ~i_RtoB_ACK0 & ~n42732;
  assign n42734 = ~n17943 & ~n42733;
  assign n42735 = controllable_DEQ & ~n42734;
  assign n42736 = ~n24537 & ~n42735;
  assign n42737 = ~i_FULL & ~n42736;
  assign n42738 = ~n42731 & ~n42737;
  assign n42739 = ~i_nEMPTY & ~n42738;
  assign n42740 = ~n42725 & ~n42739;
  assign n42741 = ~controllable_BtoS_ACK0 & ~n42740;
  assign n42742 = ~n24502 & ~n42741;
  assign n42743 = ~n4465 & ~n42742;
  assign n42744 = ~n42709 & ~n42743;
  assign n42745 = i_StoB_REQ10 & ~n42744;
  assign n42746 = ~n42597 & ~n42745;
  assign n42747 = ~controllable_BtoS_ACK10 & ~n42746;
  assign n42748 = ~n42599 & ~n42747;
  assign n42749 = n4464 & ~n42748;
  assign n42750 = ~n7919 & ~n17280;
  assign n42751 = i_RtoB_ACK0 & ~n42750;
  assign n42752 = ~n15889 & ~n39305;
  assign n42753 = ~i_RtoB_ACK0 & ~n42752;
  assign n42754 = ~n42751 & ~n42753;
  assign n42755 = controllable_DEQ & ~n42754;
  assign n42756 = ~n24621 & ~n42755;
  assign n42757 = i_FULL & ~n42756;
  assign n42758 = ~n15927 & ~n39315;
  assign n42759 = ~i_RtoB_ACK0 & ~n42758;
  assign n42760 = ~n42751 & ~n42759;
  assign n42761 = controllable_DEQ & ~n42760;
  assign n42762 = ~n24631 & ~n42761;
  assign n42763 = ~i_FULL & ~n42762;
  assign n42764 = ~n42757 & ~n42763;
  assign n42765 = i_nEMPTY & ~n42764;
  assign n42766 = ~n15964 & ~n39325;
  assign n42767 = ~i_RtoB_ACK0 & ~n42766;
  assign n42768 = ~n15217 & ~n42767;
  assign n42769 = controllable_DEQ & ~n42768;
  assign n42770 = ~n24641 & ~n42769;
  assign n42771 = i_FULL & ~n42770;
  assign n42772 = ~n15999 & ~n39333;
  assign n42773 = ~i_RtoB_ACK0 & ~n42772;
  assign n42774 = ~n15245 & ~n42773;
  assign n42775 = controllable_DEQ & ~n42774;
  assign n42776 = ~n24647 & ~n42775;
  assign n42777 = ~i_FULL & ~n42776;
  assign n42778 = ~n42771 & ~n42777;
  assign n42779 = ~i_nEMPTY & ~n42778;
  assign n42780 = ~n42765 & ~n42779;
  assign n42781 = controllable_BtoS_ACK0 & ~n42780;
  assign n42782 = ~n8086 & ~n17690;
  assign n42783 = i_RtoB_ACK0 & ~n42782;
  assign n42784 = ~n16031 & ~n39349;
  assign n42785 = ~i_RtoB_ACK0 & ~n42784;
  assign n42786 = ~n42783 & ~n42785;
  assign n42787 = controllable_DEQ & ~n42786;
  assign n42788 = ~n24665 & ~n42787;
  assign n42789 = i_FULL & ~n42788;
  assign n42790 = ~n16069 & ~n39359;
  assign n42791 = ~i_RtoB_ACK0 & ~n42790;
  assign n42792 = ~n42783 & ~n42791;
  assign n42793 = controllable_DEQ & ~n42792;
  assign n42794 = ~n24675 & ~n42793;
  assign n42795 = ~i_FULL & ~n42794;
  assign n42796 = ~n42789 & ~n42795;
  assign n42797 = i_nEMPTY & ~n42796;
  assign n42798 = ~n16106 & ~n39369;
  assign n42799 = ~i_RtoB_ACK0 & ~n42798;
  assign n42800 = ~n17731 & ~n42799;
  assign n42801 = controllable_DEQ & ~n42800;
  assign n42802 = ~n24685 & ~n42801;
  assign n42803 = i_FULL & ~n42802;
  assign n42804 = ~n16141 & ~n39377;
  assign n42805 = ~i_RtoB_ACK0 & ~n42804;
  assign n42806 = ~n17764 & ~n42805;
  assign n42807 = controllable_DEQ & ~n42806;
  assign n42808 = ~n24691 & ~n42807;
  assign n42809 = ~i_FULL & ~n42808;
  assign n42810 = ~n42803 & ~n42809;
  assign n42811 = ~i_nEMPTY & ~n42810;
  assign n42812 = ~n42797 & ~n42811;
  assign n42813 = ~controllable_BtoS_ACK0 & ~n42812;
  assign n42814 = ~n42781 & ~n42813;
  assign n42815 = n4465 & ~n42814;
  assign n42816 = ~n8329 & ~n17690;
  assign n42817 = i_RtoB_ACK0 & ~n42816;
  assign n42818 = ~n16262 & ~n39391;
  assign n42819 = ~i_RtoB_ACK0 & ~n42818;
  assign n42820 = ~n42817 & ~n42819;
  assign n42821 = controllable_DEQ & ~n42820;
  assign n42822 = ~n24743 & ~n42821;
  assign n42823 = i_FULL & ~n42822;
  assign n42824 = ~n16300 & ~n39399;
  assign n42825 = ~i_RtoB_ACK0 & ~n42824;
  assign n42826 = ~n42817 & ~n42825;
  assign n42827 = controllable_DEQ & ~n42826;
  assign n42828 = ~n24753 & ~n42827;
  assign n42829 = ~i_FULL & ~n42828;
  assign n42830 = ~n42823 & ~n42829;
  assign n42831 = i_nEMPTY & ~n42830;
  assign n42832 = ~n16337 & ~n39409;
  assign n42833 = ~i_RtoB_ACK0 & ~n42832;
  assign n42834 = ~n17731 & ~n42833;
  assign n42835 = controllable_DEQ & ~n42834;
  assign n42836 = ~n24763 & ~n42835;
  assign n42837 = i_FULL & ~n42836;
  assign n42838 = ~n16372 & ~n39417;
  assign n42839 = ~i_RtoB_ACK0 & ~n42838;
  assign n42840 = ~n17764 & ~n42839;
  assign n42841 = controllable_DEQ & ~n42840;
  assign n42842 = ~n24769 & ~n42841;
  assign n42843 = ~i_FULL & ~n42842;
  assign n42844 = ~n42837 & ~n42843;
  assign n42845 = ~i_nEMPTY & ~n42844;
  assign n42846 = ~n42831 & ~n42845;
  assign n42847 = ~controllable_BtoS_ACK0 & ~n42846;
  assign n42848 = ~n24731 & ~n42847;
  assign n42849 = ~n4465 & ~n42848;
  assign n42850 = ~n42815 & ~n42849;
  assign n42851 = ~i_StoB_REQ10 & ~n42850;
  assign n42852 = ~n24609 & ~n42851;
  assign n42853 = controllable_BtoS_ACK10 & ~n42852;
  assign n42854 = ~n8466 & ~n17050;
  assign n42855 = i_RtoB_ACK0 & ~n42854;
  assign n42856 = ~n20002 & ~n39435;
  assign n42857 = ~i_RtoB_ACK0 & ~n42856;
  assign n42858 = ~n42855 & ~n42857;
  assign n42859 = controllable_DEQ & ~n42858;
  assign n42860 = ~n24793 & ~n42859;
  assign n42861 = i_FULL & ~n42860;
  assign n42862 = ~n20022 & ~n39443;
  assign n42863 = ~i_RtoB_ACK0 & ~n42862;
  assign n42864 = ~n42855 & ~n42863;
  assign n42865 = controllable_DEQ & ~n42864;
  assign n42866 = ~n24803 & ~n42865;
  assign n42867 = ~i_FULL & ~n42866;
  assign n42868 = ~n42861 & ~n42867;
  assign n42869 = i_nEMPTY & ~n42868;
  assign n42870 = ~n20040 & ~n39453;
  assign n42871 = ~i_RtoB_ACK0 & ~n42870;
  assign n42872 = ~n15604 & ~n42871;
  assign n42873 = controllable_DEQ & ~n42872;
  assign n42874 = ~n24813 & ~n42873;
  assign n42875 = i_FULL & ~n42874;
  assign n42876 = ~n20056 & ~n39461;
  assign n42877 = ~i_RtoB_ACK0 & ~n42876;
  assign n42878 = ~n15619 & ~n42877;
  assign n42879 = controllable_DEQ & ~n42878;
  assign n42880 = ~n24816 & ~n42879;
  assign n42881 = ~i_FULL & ~n42880;
  assign n42882 = ~n42875 & ~n42881;
  assign n42883 = ~i_nEMPTY & ~n42882;
  assign n42884 = ~n42869 & ~n42883;
  assign n42885 = controllable_BtoS_ACK0 & ~n42884;
  assign n42886 = ~n8545 & ~n18522;
  assign n42887 = i_RtoB_ACK0 & ~n42886;
  assign n42888 = ~n20068 & ~n39473;
  assign n42889 = ~i_RtoB_ACK0 & ~n42888;
  assign n42890 = ~n42887 & ~n42889;
  assign n42891 = controllable_DEQ & ~n42890;
  assign n42892 = ~n24834 & ~n42891;
  assign n42893 = i_FULL & ~n42892;
  assign n42894 = ~n20080 & ~n39481;
  assign n42895 = ~i_RtoB_ACK0 & ~n42894;
  assign n42896 = ~n42887 & ~n42895;
  assign n42897 = controllable_DEQ & ~n42896;
  assign n42898 = ~n24844 & ~n42897;
  assign n42899 = ~i_FULL & ~n42898;
  assign n42900 = ~n42893 & ~n42899;
  assign n42901 = i_nEMPTY & ~n42900;
  assign n42902 = ~n20094 & ~n39491;
  assign n42903 = ~i_RtoB_ACK0 & ~n42902;
  assign n42904 = ~n17925 & ~n42903;
  assign n42905 = controllable_DEQ & ~n42904;
  assign n42906 = ~n24854 & ~n42905;
  assign n42907 = i_FULL & ~n42906;
  assign n42908 = ~n20106 & ~n39499;
  assign n42909 = ~i_RtoB_ACK0 & ~n42908;
  assign n42910 = ~n17943 & ~n42909;
  assign n42911 = controllable_DEQ & ~n42910;
  assign n42912 = ~n24857 & ~n42911;
  assign n42913 = ~i_FULL & ~n42912;
  assign n42914 = ~n42907 & ~n42913;
  assign n42915 = ~i_nEMPTY & ~n42914;
  assign n42916 = ~n42901 & ~n42915;
  assign n42917 = ~controllable_BtoS_ACK0 & ~n42916;
  assign n42918 = ~n42885 & ~n42917;
  assign n42919 = n4465 & ~n42918;
  assign n42920 = ~n8677 & ~n18522;
  assign n42921 = i_RtoB_ACK0 & ~n42920;
  assign n42922 = ~n20156 & ~n39513;
  assign n42923 = ~i_RtoB_ACK0 & ~n42922;
  assign n42924 = ~n42921 & ~n42923;
  assign n42925 = controllable_DEQ & ~n42924;
  assign n42926 = ~n24906 & ~n42925;
  assign n42927 = i_FULL & ~n42926;
  assign n42928 = ~n20168 & ~n39521;
  assign n42929 = ~i_RtoB_ACK0 & ~n42928;
  assign n42930 = ~n42921 & ~n42929;
  assign n42931 = controllable_DEQ & ~n42930;
  assign n42932 = ~n24916 & ~n42931;
  assign n42933 = ~i_FULL & ~n42932;
  assign n42934 = ~n42927 & ~n42933;
  assign n42935 = i_nEMPTY & ~n42934;
  assign n42936 = ~n20182 & ~n39531;
  assign n42937 = ~i_RtoB_ACK0 & ~n42936;
  assign n42938 = ~n17925 & ~n42937;
  assign n42939 = controllable_DEQ & ~n42938;
  assign n42940 = ~n24926 & ~n42939;
  assign n42941 = i_FULL & ~n42940;
  assign n42942 = ~n20194 & ~n39539;
  assign n42943 = ~i_RtoB_ACK0 & ~n42942;
  assign n42944 = ~n17943 & ~n42943;
  assign n42945 = controllable_DEQ & ~n42944;
  assign n42946 = ~n24929 & ~n42945;
  assign n42947 = ~i_FULL & ~n42946;
  assign n42948 = ~n42941 & ~n42947;
  assign n42949 = ~i_nEMPTY & ~n42948;
  assign n42950 = ~n42935 & ~n42949;
  assign n42951 = ~controllable_BtoS_ACK0 & ~n42950;
  assign n42952 = ~n24894 & ~n42951;
  assign n42953 = ~n4465 & ~n42952;
  assign n42954 = ~n42919 & ~n42953;
  assign n42955 = i_StoB_REQ10 & ~n42954;
  assign n42956 = ~n42851 & ~n42955;
  assign n42957 = ~controllable_BtoS_ACK10 & ~n42956;
  assign n42958 = ~n42853 & ~n42957;
  assign n42959 = ~n4464 & ~n42958;
  assign n42960 = ~n42749 & ~n42959;
  assign n42961 = n4463 & ~n42960;
  assign n42962 = ~n25577 & ~n41595;
  assign n42963 = i_FULL & ~n42962;
  assign n42964 = ~n25577 & ~n41601;
  assign n42965 = ~i_FULL & ~n42964;
  assign n42966 = ~n42963 & ~n42965;
  assign n42967 = i_nEMPTY & ~n42966;
  assign n42968 = ~n41621 & ~n42967;
  assign n42969 = controllable_BtoS_ACK0 & ~n42968;
  assign n42970 = ~n25599 & ~n41629;
  assign n42971 = i_FULL & ~n42970;
  assign n42972 = ~n25599 & ~n41635;
  assign n42973 = ~i_FULL & ~n42972;
  assign n42974 = ~n42971 & ~n42973;
  assign n42975 = i_nEMPTY & ~n42974;
  assign n42976 = ~n41655 & ~n42975;
  assign n42977 = ~controllable_BtoS_ACK0 & ~n42976;
  assign n42978 = ~n42969 & ~n42977;
  assign n42979 = n4465 & ~n42978;
  assign n42980 = ~n41667 & ~n42979;
  assign n42981 = i_StoB_REQ10 & ~n42980;
  assign n42982 = ~n17280 & ~n37252;
  assign n42983 = i_RtoB_ACK0 & ~n42982;
  assign n42984 = ~n41673 & ~n42983;
  assign n42985 = controllable_DEQ & ~n42984;
  assign n42986 = ~n37460 & ~n40722;
  assign n42987 = i_RtoB_ACK0 & ~n42986;
  assign n42988 = ~n41679 & ~n42987;
  assign n42989 = ~controllable_DEQ & ~n42988;
  assign n42990 = ~n42985 & ~n42989;
  assign n42991 = i_FULL & ~n42990;
  assign n42992 = ~n41685 & ~n42983;
  assign n42993 = controllable_DEQ & ~n42992;
  assign n42994 = ~n41689 & ~n42987;
  assign n42995 = ~controllable_DEQ & ~n42994;
  assign n42996 = ~n42993 & ~n42995;
  assign n42997 = ~i_FULL & ~n42996;
  assign n42998 = ~n42991 & ~n42997;
  assign n42999 = i_nEMPTY & ~n42998;
  assign n43000 = ~n15217 & ~n41697;
  assign n43001 = controllable_DEQ & ~n43000;
  assign n43002 = ~n37522 & ~n40760;
  assign n43003 = i_RtoB_ACK0 & ~n43002;
  assign n43004 = ~n41703 & ~n43003;
  assign n43005 = ~controllable_DEQ & ~n43004;
  assign n43006 = ~n43001 & ~n43005;
  assign n43007 = i_FULL & ~n43006;
  assign n43008 = ~n15245 & ~n41709;
  assign n43009 = controllable_DEQ & ~n43008;
  assign n43010 = ~n37522 & ~n40783;
  assign n43011 = i_RtoB_ACK0 & ~n43010;
  assign n43012 = ~n41715 & ~n43011;
  assign n43013 = ~controllable_DEQ & ~n43012;
  assign n43014 = ~n43009 & ~n43013;
  assign n43015 = ~i_FULL & ~n43014;
  assign n43016 = ~n43007 & ~n43015;
  assign n43017 = ~i_nEMPTY & ~n43016;
  assign n43018 = ~n42999 & ~n43017;
  assign n43019 = controllable_BtoS_ACK0 & ~n43018;
  assign n43020 = ~n17690 & ~n37694;
  assign n43021 = i_RtoB_ACK0 & ~n43020;
  assign n43022 = ~n41727 & ~n43021;
  assign n43023 = controllable_DEQ & ~n43022;
  assign n43024 = ~n37723 & ~n40814;
  assign n43025 = i_RtoB_ACK0 & ~n43024;
  assign n43026 = ~n41733 & ~n43025;
  assign n43027 = ~controllable_DEQ & ~n43026;
  assign n43028 = ~n43023 & ~n43027;
  assign n43029 = i_FULL & ~n43028;
  assign n43030 = ~n41739 & ~n43021;
  assign n43031 = controllable_DEQ & ~n43030;
  assign n43032 = ~n41743 & ~n43025;
  assign n43033 = ~controllable_DEQ & ~n43032;
  assign n43034 = ~n43031 & ~n43033;
  assign n43035 = ~i_FULL & ~n43034;
  assign n43036 = ~n43029 & ~n43035;
  assign n43037 = i_nEMPTY & ~n43036;
  assign n43038 = ~n17731 & ~n41751;
  assign n43039 = controllable_DEQ & ~n43038;
  assign n43040 = ~n37785 & ~n40852;
  assign n43041 = i_RtoB_ACK0 & ~n43040;
  assign n43042 = ~n41757 & ~n43041;
  assign n43043 = ~controllable_DEQ & ~n43042;
  assign n43044 = ~n43039 & ~n43043;
  assign n43045 = i_FULL & ~n43044;
  assign n43046 = ~n17764 & ~n41763;
  assign n43047 = controllable_DEQ & ~n43046;
  assign n43048 = ~n37785 & ~n40875;
  assign n43049 = i_RtoB_ACK0 & ~n43048;
  assign n43050 = ~n41769 & ~n43049;
  assign n43051 = ~controllable_DEQ & ~n43050;
  assign n43052 = ~n43047 & ~n43051;
  assign n43053 = ~i_FULL & ~n43052;
  assign n43054 = ~n43045 & ~n43053;
  assign n43055 = ~i_nEMPTY & ~n43054;
  assign n43056 = ~n43037 & ~n43055;
  assign n43057 = ~controllable_BtoS_ACK0 & ~n43056;
  assign n43058 = ~n43019 & ~n43057;
  assign n43059 = n4465 & ~n43058;
  assign n43060 = ~n17690 & ~n37846;
  assign n43061 = i_RtoB_ACK0 & ~n43060;
  assign n43062 = ~n41783 & ~n43061;
  assign n43063 = controllable_DEQ & ~n43062;
  assign n43064 = ~n22297 & ~n43063;
  assign n43065 = i_FULL & ~n43064;
  assign n43066 = ~n41789 & ~n43061;
  assign n43067 = controllable_DEQ & ~n43066;
  assign n43068 = ~n22307 & ~n43067;
  assign n43069 = ~i_FULL & ~n43068;
  assign n43070 = ~n43065 & ~n43069;
  assign n43071 = i_nEMPTY & ~n43070;
  assign n43072 = ~n41809 & ~n43071;
  assign n43073 = ~controllable_BtoS_ACK0 & ~n43072;
  assign n43074 = ~n25035 & ~n43073;
  assign n43075 = ~n4465 & ~n43074;
  assign n43076 = ~n43059 & ~n43075;
  assign n43077 = ~i_StoB_REQ10 & ~n43076;
  assign n43078 = ~n42981 & ~n43077;
  assign n43079 = controllable_BtoS_ACK10 & ~n43078;
  assign n43080 = ~n17050 & ~n37904;
  assign n43081 = i_RtoB_ACK0 & ~n43080;
  assign n43082 = ~n41821 & ~n43081;
  assign n43083 = controllable_DEQ & ~n43082;
  assign n43084 = ~n41829 & ~n43083;
  assign n43085 = i_FULL & ~n43084;
  assign n43086 = ~n41833 & ~n43081;
  assign n43087 = controllable_DEQ & ~n43086;
  assign n43088 = ~n41839 & ~n43087;
  assign n43089 = ~i_FULL & ~n43088;
  assign n43090 = ~n43085 & ~n43089;
  assign n43091 = i_nEMPTY & ~n43090;
  assign n43092 = ~n15604 & ~n41845;
  assign n43093 = controllable_DEQ & ~n43092;
  assign n43094 = ~n41853 & ~n43093;
  assign n43095 = i_FULL & ~n43094;
  assign n43096 = ~n15619 & ~n41857;
  assign n43097 = controllable_DEQ & ~n43096;
  assign n43098 = ~n41865 & ~n43097;
  assign n43099 = ~i_FULL & ~n43098;
  assign n43100 = ~n43095 & ~n43099;
  assign n43101 = ~i_nEMPTY & ~n43100;
  assign n43102 = ~n43091 & ~n43101;
  assign n43103 = controllable_BtoS_ACK0 & ~n43102;
  assign n43104 = ~n18522 & ~n37988;
  assign n43105 = i_RtoB_ACK0 & ~n43104;
  assign n43106 = ~n41875 & ~n43105;
  assign n43107 = controllable_DEQ & ~n43106;
  assign n43108 = ~n41883 & ~n43107;
  assign n43109 = i_FULL & ~n43108;
  assign n43110 = ~n41887 & ~n43105;
  assign n43111 = controllable_DEQ & ~n43110;
  assign n43112 = ~n41893 & ~n43111;
  assign n43113 = ~i_FULL & ~n43112;
  assign n43114 = ~n43109 & ~n43113;
  assign n43115 = i_nEMPTY & ~n43114;
  assign n43116 = ~n17925 & ~n41899;
  assign n43117 = controllable_DEQ & ~n43116;
  assign n43118 = ~n41907 & ~n43117;
  assign n43119 = i_FULL & ~n43118;
  assign n43120 = ~n17943 & ~n41911;
  assign n43121 = controllable_DEQ & ~n43120;
  assign n43122 = ~n41919 & ~n43121;
  assign n43123 = ~i_FULL & ~n43122;
  assign n43124 = ~n43119 & ~n43123;
  assign n43125 = ~i_nEMPTY & ~n43124;
  assign n43126 = ~n43115 & ~n43125;
  assign n43127 = ~controllable_BtoS_ACK0 & ~n43126;
  assign n43128 = ~n43103 & ~n43127;
  assign n43129 = n4465 & ~n43128;
  assign n43130 = ~n18522 & ~n38074;
  assign n43131 = i_RtoB_ACK0 & ~n43130;
  assign n43132 = ~n41931 & ~n43131;
  assign n43133 = controllable_DEQ & ~n43132;
  assign n43134 = ~n22492 & ~n43133;
  assign n43135 = i_FULL & ~n43134;
  assign n43136 = ~n41937 & ~n43131;
  assign n43137 = controllable_DEQ & ~n43136;
  assign n43138 = ~n22502 & ~n43137;
  assign n43139 = ~i_FULL & ~n43138;
  assign n43140 = ~n43135 & ~n43139;
  assign n43141 = i_nEMPTY & ~n43140;
  assign n43142 = ~n41957 & ~n43141;
  assign n43143 = ~controllable_BtoS_ACK0 & ~n43142;
  assign n43144 = ~n22480 & ~n43143;
  assign n43145 = ~n4465 & ~n43144;
  assign n43146 = ~n43129 & ~n43145;
  assign n43147 = i_StoB_REQ10 & ~n43146;
  assign n43148 = ~n43077 & ~n43147;
  assign n43149 = ~controllable_BtoS_ACK10 & ~n43148;
  assign n43150 = ~n43079 & ~n43149;
  assign n43151 = n4464 & ~n43150;
  assign n43152 = ~n17280 & ~n38152;
  assign n43153 = i_RtoB_ACK0 & ~n43152;
  assign n43154 = ~n41989 & ~n43153;
  assign n43155 = controllable_DEQ & ~n43154;
  assign n43156 = ~n25053 & ~n43155;
  assign n43157 = i_FULL & ~n43156;
  assign n43158 = ~n41995 & ~n43153;
  assign n43159 = controllable_DEQ & ~n43158;
  assign n43160 = ~n25059 & ~n43159;
  assign n43161 = ~i_FULL & ~n43160;
  assign n43162 = ~n43157 & ~n43161;
  assign n43163 = i_nEMPTY & ~n43162;
  assign n43164 = ~n25067 & ~n42005;
  assign n43165 = i_FULL & ~n43164;
  assign n43166 = ~n25071 & ~n42011;
  assign n43167 = ~i_FULL & ~n43166;
  assign n43168 = ~n43165 & ~n43167;
  assign n43169 = ~i_nEMPTY & ~n43168;
  assign n43170 = ~n43163 & ~n43169;
  assign n43171 = controllable_BtoS_ACK0 & ~n43170;
  assign n43172 = ~n17690 & ~n38204;
  assign n43173 = i_RtoB_ACK0 & ~n43172;
  assign n43174 = ~n42021 & ~n43173;
  assign n43175 = controllable_DEQ & ~n43174;
  assign n43176 = ~n25085 & ~n43175;
  assign n43177 = i_FULL & ~n43176;
  assign n43178 = ~n42027 & ~n43173;
  assign n43179 = controllable_DEQ & ~n43178;
  assign n43180 = ~n25091 & ~n43179;
  assign n43181 = ~i_FULL & ~n43180;
  assign n43182 = ~n43177 & ~n43181;
  assign n43183 = i_nEMPTY & ~n43182;
  assign n43184 = ~n25099 & ~n42037;
  assign n43185 = i_FULL & ~n43184;
  assign n43186 = ~n25103 & ~n42043;
  assign n43187 = ~i_FULL & ~n43186;
  assign n43188 = ~n43185 & ~n43187;
  assign n43189 = ~i_nEMPTY & ~n43188;
  assign n43190 = ~n43183 & ~n43189;
  assign n43191 = ~controllable_BtoS_ACK0 & ~n43190;
  assign n43192 = ~n43171 & ~n43191;
  assign n43193 = n4465 & ~n43192;
  assign n43194 = ~n17690 & ~n38258;
  assign n43195 = i_RtoB_ACK0 & ~n43194;
  assign n43196 = ~n42055 & ~n43195;
  assign n43197 = controllable_DEQ & ~n43196;
  assign n43198 = ~n22801 & ~n43197;
  assign n43199 = i_FULL & ~n43198;
  assign n43200 = ~n42061 & ~n43195;
  assign n43201 = controllable_DEQ & ~n43200;
  assign n43202 = ~n22811 & ~n43201;
  assign n43203 = ~i_FULL & ~n43202;
  assign n43204 = ~n43199 & ~n43203;
  assign n43205 = i_nEMPTY & ~n43204;
  assign n43206 = ~n42081 & ~n43205;
  assign n43207 = ~controllable_BtoS_ACK0 & ~n43206;
  assign n43208 = ~n22789 & ~n43207;
  assign n43209 = ~n4465 & ~n43208;
  assign n43210 = ~n43193 & ~n43209;
  assign n43211 = ~i_StoB_REQ10 & ~n43210;
  assign n43212 = ~n41985 & ~n43211;
  assign n43213 = controllable_BtoS_ACK10 & ~n43212;
  assign n43214 = ~n17050 & ~n38316;
  assign n43215 = i_RtoB_ACK0 & ~n43214;
  assign n43216 = ~n42093 & ~n43215;
  assign n43217 = controllable_DEQ & ~n43216;
  assign n43218 = ~n22859 & ~n43217;
  assign n43219 = i_FULL & ~n43218;
  assign n43220 = ~n42099 & ~n43215;
  assign n43221 = controllable_DEQ & ~n43220;
  assign n43222 = ~n22869 & ~n43221;
  assign n43223 = ~i_FULL & ~n43222;
  assign n43224 = ~n43219 & ~n43223;
  assign n43225 = i_nEMPTY & ~n43224;
  assign n43226 = ~n42119 & ~n43225;
  assign n43227 = controllable_BtoS_ACK0 & ~n43226;
  assign n43228 = ~n18522 & ~n38368;
  assign n43229 = i_RtoB_ACK0 & ~n43228;
  assign n43230 = ~n42125 & ~n43229;
  assign n43231 = controllable_DEQ & ~n43230;
  assign n43232 = ~n22908 & ~n43231;
  assign n43233 = i_FULL & ~n43232;
  assign n43234 = ~n42131 & ~n43229;
  assign n43235 = controllable_DEQ & ~n43234;
  assign n43236 = ~n22918 & ~n43235;
  assign n43237 = ~i_FULL & ~n43236;
  assign n43238 = ~n43233 & ~n43237;
  assign n43239 = i_nEMPTY & ~n43238;
  assign n43240 = ~n42151 & ~n43239;
  assign n43241 = ~controllable_BtoS_ACK0 & ~n43240;
  assign n43242 = ~n43227 & ~n43241;
  assign n43243 = n4465 & ~n43242;
  assign n43244 = ~n18522 & ~n38422;
  assign n43245 = i_RtoB_ACK0 & ~n43244;
  assign n43246 = ~n42159 & ~n43245;
  assign n43247 = controllable_DEQ & ~n43246;
  assign n43248 = ~n22996 & ~n43247;
  assign n43249 = i_FULL & ~n43248;
  assign n43250 = ~n42165 & ~n43245;
  assign n43251 = controllable_DEQ & ~n43250;
  assign n43252 = ~n23006 & ~n43251;
  assign n43253 = ~i_FULL & ~n43252;
  assign n43254 = ~n43249 & ~n43253;
  assign n43255 = i_nEMPTY & ~n43254;
  assign n43256 = ~n42185 & ~n43255;
  assign n43257 = ~controllable_BtoS_ACK0 & ~n43256;
  assign n43258 = ~n22984 & ~n43257;
  assign n43259 = ~n4465 & ~n43258;
  assign n43260 = ~n43243 & ~n43259;
  assign n43261 = i_StoB_REQ10 & ~n43260;
  assign n43262 = ~n43211 & ~n43261;
  assign n43263 = ~controllable_BtoS_ACK10 & ~n43262;
  assign n43264 = ~n43213 & ~n43263;
  assign n43265 = ~n4464 & ~n43264;
  assign n43266 = ~n43151 & ~n43265;
  assign n43267 = ~n4463 & ~n43266;
  assign n43268 = ~n42961 & ~n43267;
  assign n43269 = n4462 & ~n43268;
  assign n43270 = ~n17974 & ~n39563;
  assign n43271 = ~i_RtoB_ACK0 & ~n43270;
  assign n43272 = ~n42453 & ~n43271;
  assign n43273 = controllable_DEQ & ~n43272;
  assign n43274 = ~n25285 & ~n43273;
  assign n43275 = i_FULL & ~n43274;
  assign n43276 = ~n18012 & ~n39571;
  assign n43277 = ~i_RtoB_ACK0 & ~n43276;
  assign n43278 = ~n42453 & ~n43277;
  assign n43279 = controllable_DEQ & ~n43278;
  assign n43280 = ~n25295 & ~n43279;
  assign n43281 = ~i_FULL & ~n43280;
  assign n43282 = ~n43275 & ~n43281;
  assign n43283 = i_nEMPTY & ~n43282;
  assign n43284 = ~n18049 & ~n39581;
  assign n43285 = ~i_RtoB_ACK0 & ~n43284;
  assign n43286 = ~n15217 & ~n43285;
  assign n43287 = controllable_DEQ & ~n43286;
  assign n43288 = ~n25305 & ~n43287;
  assign n43289 = i_FULL & ~n43288;
  assign n43290 = ~n18084 & ~n39589;
  assign n43291 = ~i_RtoB_ACK0 & ~n43290;
  assign n43292 = ~n15245 & ~n43291;
  assign n43293 = controllable_DEQ & ~n43292;
  assign n43294 = ~n25311 & ~n43293;
  assign n43295 = ~i_FULL & ~n43294;
  assign n43296 = ~n43289 & ~n43295;
  assign n43297 = ~i_nEMPTY & ~n43296;
  assign n43298 = ~n43283 & ~n43297;
  assign n43299 = controllable_BtoS_ACK0 & ~n43298;
  assign n43300 = ~n18116 & ~n39601;
  assign n43301 = ~i_RtoB_ACK0 & ~n43300;
  assign n43302 = ~n42507 & ~n43301;
  assign n43303 = controllable_DEQ & ~n43302;
  assign n43304 = ~n25329 & ~n43303;
  assign n43305 = i_FULL & ~n43304;
  assign n43306 = ~n18154 & ~n39609;
  assign n43307 = ~i_RtoB_ACK0 & ~n43306;
  assign n43308 = ~n42507 & ~n43307;
  assign n43309 = controllable_DEQ & ~n43308;
  assign n43310 = ~n25339 & ~n43309;
  assign n43311 = ~i_FULL & ~n43310;
  assign n43312 = ~n43305 & ~n43311;
  assign n43313 = i_nEMPTY & ~n43312;
  assign n43314 = ~n18191 & ~n39619;
  assign n43315 = ~i_RtoB_ACK0 & ~n43314;
  assign n43316 = ~n17731 & ~n43315;
  assign n43317 = controllable_DEQ & ~n43316;
  assign n43318 = ~n25349 & ~n43317;
  assign n43319 = i_FULL & ~n43318;
  assign n43320 = ~n18226 & ~n39627;
  assign n43321 = ~i_RtoB_ACK0 & ~n43320;
  assign n43322 = ~n17764 & ~n43321;
  assign n43323 = controllable_DEQ & ~n43322;
  assign n43324 = ~n25355 & ~n43323;
  assign n43325 = ~i_FULL & ~n43324;
  assign n43326 = ~n43319 & ~n43325;
  assign n43327 = ~i_nEMPTY & ~n43326;
  assign n43328 = ~n43313 & ~n43327;
  assign n43329 = ~controllable_BtoS_ACK0 & ~n43328;
  assign n43330 = ~n43299 & ~n43329;
  assign n43331 = n4465 & ~n43330;
  assign n43332 = ~n25389 & ~n42593;
  assign n43333 = ~n4465 & ~n43332;
  assign n43334 = ~n43331 & ~n43333;
  assign n43335 = ~i_StoB_REQ10 & ~n43334;
  assign n43336 = ~n25273 & ~n43335;
  assign n43337 = ~controllable_BtoS_ACK10 & ~n43336;
  assign n43338 = ~n25185 & ~n43337;
  assign n43339 = n4464 & ~n43338;
  assign n43340 = ~n15889 & ~n39649;
  assign n43341 = ~i_RtoB_ACK0 & ~n43340;
  assign n43342 = ~n42751 & ~n43341;
  assign n43343 = controllable_DEQ & ~n43342;
  assign n43344 = ~n25495 & ~n43343;
  assign n43345 = i_FULL & ~n43344;
  assign n43346 = ~n15927 & ~n39657;
  assign n43347 = ~i_RtoB_ACK0 & ~n43346;
  assign n43348 = ~n42751 & ~n43347;
  assign n43349 = controllable_DEQ & ~n43348;
  assign n43350 = ~n25505 & ~n43349;
  assign n43351 = ~i_FULL & ~n43350;
  assign n43352 = ~n43345 & ~n43351;
  assign n43353 = i_nEMPTY & ~n43352;
  assign n43354 = ~n25513 & ~n42769;
  assign n43355 = i_FULL & ~n43354;
  assign n43356 = ~n25519 & ~n42775;
  assign n43357 = ~i_FULL & ~n43356;
  assign n43358 = ~n43355 & ~n43357;
  assign n43359 = ~i_nEMPTY & ~n43358;
  assign n43360 = ~n43353 & ~n43359;
  assign n43361 = controllable_BtoS_ACK0 & ~n43360;
  assign n43362 = ~n16031 & ~n39675;
  assign n43363 = ~i_RtoB_ACK0 & ~n43362;
  assign n43364 = ~n42783 & ~n43363;
  assign n43365 = controllable_DEQ & ~n43364;
  assign n43366 = ~n25533 & ~n43365;
  assign n43367 = i_FULL & ~n43366;
  assign n43368 = ~n16069 & ~n39683;
  assign n43369 = ~i_RtoB_ACK0 & ~n43368;
  assign n43370 = ~n42783 & ~n43369;
  assign n43371 = controllable_DEQ & ~n43370;
  assign n43372 = ~n25543 & ~n43371;
  assign n43373 = ~i_FULL & ~n43372;
  assign n43374 = ~n43367 & ~n43373;
  assign n43375 = i_nEMPTY & ~n43374;
  assign n43376 = ~n25551 & ~n42801;
  assign n43377 = i_FULL & ~n43376;
  assign n43378 = ~n25557 & ~n42807;
  assign n43379 = ~i_FULL & ~n43378;
  assign n43380 = ~n43377 & ~n43379;
  assign n43381 = ~i_nEMPTY & ~n43380;
  assign n43382 = ~n43375 & ~n43381;
  assign n43383 = ~controllable_BtoS_ACK0 & ~n43382;
  assign n43384 = ~n43361 & ~n43383;
  assign n43385 = n4465 & ~n43384;
  assign n43386 = ~n42849 & ~n43385;
  assign n43387 = ~i_StoB_REQ10 & ~n43386;
  assign n43388 = ~n25487 & ~n43387;
  assign n43389 = ~controllable_BtoS_ACK10 & ~n43388;
  assign n43390 = ~n25399 & ~n43389;
  assign n43391 = ~n4464 & ~n43390;
  assign n43392 = ~n43339 & ~n43391;
  assign n43393 = n4463 & ~n43392;
  assign n43394 = ~n17280 & ~n38514;
  assign n43395 = i_RtoB_ACK0 & ~n43394;
  assign n43396 = ~n42229 & ~n43395;
  assign n43397 = controllable_DEQ & ~n43396;
  assign n43398 = ~n23739 & ~n43397;
  assign n43399 = i_FULL & ~n43398;
  assign n43400 = ~n42235 & ~n43395;
  assign n43401 = controllable_DEQ & ~n43400;
  assign n43402 = ~n23749 & ~n43401;
  assign n43403 = ~i_FULL & ~n43402;
  assign n43404 = ~n43399 & ~n43403;
  assign n43405 = i_nEMPTY & ~n43404;
  assign n43406 = ~n42255 & ~n43405;
  assign n43407 = controllable_BtoS_ACK0 & ~n43406;
  assign n43408 = ~n17690 & ~n38556;
  assign n43409 = i_RtoB_ACK0 & ~n43408;
  assign n43410 = ~n42261 & ~n43409;
  assign n43411 = controllable_DEQ & ~n43410;
  assign n43412 = ~n23791 & ~n43411;
  assign n43413 = i_FULL & ~n43412;
  assign n43414 = ~n42267 & ~n43409;
  assign n43415 = controllable_DEQ & ~n43414;
  assign n43416 = ~n23801 & ~n43415;
  assign n43417 = ~i_FULL & ~n43416;
  assign n43418 = ~n43413 & ~n43417;
  assign n43419 = i_nEMPTY & ~n43418;
  assign n43420 = ~n42287 & ~n43419;
  assign n43421 = ~controllable_BtoS_ACK0 & ~n43420;
  assign n43422 = ~n43407 & ~n43421;
  assign n43423 = n4465 & ~n43422;
  assign n43424 = ~n23867 & ~n43073;
  assign n43425 = ~n4465 & ~n43424;
  assign n43426 = ~n43423 & ~n43425;
  assign n43427 = ~i_StoB_REQ10 & ~n43426;
  assign n43428 = ~n42225 & ~n43427;
  assign n43429 = ~controllable_BtoS_ACK10 & ~n43428;
  assign n43430 = ~n25623 & ~n43429;
  assign n43431 = n4464 & ~n43430;
  assign n43432 = ~n17280 & ~n38638;
  assign n43433 = i_RtoB_ACK0 & ~n43432;
  assign n43434 = ~n42329 & ~n43433;
  assign n43435 = controllable_DEQ & ~n43434;
  assign n43436 = ~n24041 & ~n43435;
  assign n43437 = i_FULL & ~n43436;
  assign n43438 = ~n42335 & ~n43433;
  assign n43439 = controllable_DEQ & ~n43438;
  assign n43440 = ~n24049 & ~n43439;
  assign n43441 = ~i_FULL & ~n43440;
  assign n43442 = ~n43437 & ~n43441;
  assign n43443 = i_nEMPTY & ~n43442;
  assign n43444 = ~n42355 & ~n43443;
  assign n43445 = controllable_BtoS_ACK0 & ~n43444;
  assign n43446 = ~n17690 & ~n38680;
  assign n43447 = i_RtoB_ACK0 & ~n43446;
  assign n43448 = ~n42361 & ~n43447;
  assign n43449 = controllable_DEQ & ~n43448;
  assign n43450 = ~n24085 & ~n43449;
  assign n43451 = i_FULL & ~n43450;
  assign n43452 = ~n42367 & ~n43447;
  assign n43453 = controllable_DEQ & ~n43452;
  assign n43454 = ~n24093 & ~n43453;
  assign n43455 = ~i_FULL & ~n43454;
  assign n43456 = ~n43451 & ~n43455;
  assign n43457 = i_nEMPTY & ~n43456;
  assign n43458 = ~n42387 & ~n43457;
  assign n43459 = ~controllable_BtoS_ACK0 & ~n43458;
  assign n43460 = ~n43445 & ~n43459;
  assign n43461 = n4465 & ~n43460;
  assign n43462 = ~n43209 & ~n43461;
  assign n43463 = ~i_StoB_REQ10 & ~n43462;
  assign n43464 = ~n42325 & ~n43463;
  assign n43465 = ~controllable_BtoS_ACK10 & ~n43464;
  assign n43466 = ~n23927 & ~n43465;
  assign n43467 = ~n4464 & ~n43466;
  assign n43468 = ~n43431 & ~n43467;
  assign n43469 = ~n4463 & ~n43468;
  assign n43470 = ~n43393 & ~n43469;
  assign n43471 = ~n4462 & ~n43470;
  assign n43472 = ~n43269 & ~n43471;
  assign n43473 = ~n4461 & ~n43472;
  assign n43474 = ~n42403 & ~n43473;
  assign n43475 = ~n4459 & ~n43474;
  assign n43476 = ~n25855 & ~n42407;
  assign n43477 = i_nEMPTY & ~n43476;
  assign n43478 = ~n42423 & ~n43477;
  assign n43479 = controllable_BtoS_ACK0 & ~n43478;
  assign n43480 = ~n25889 & ~n42429;
  assign n43481 = i_nEMPTY & ~n43480;
  assign n43482 = ~n42445 & ~n43481;
  assign n43483 = ~controllable_BtoS_ACK0 & ~n43482;
  assign n43484 = ~n43479 & ~n43483;
  assign n43485 = n4465 & ~n43484;
  assign n43486 = ~n24215 & ~n43485;
  assign n43487 = i_StoB_REQ10 & ~n43486;
  assign n43488 = ~n11650 & ~n37154;
  assign n43489 = ~controllable_BtoR_REQ0 & ~n43488;
  assign n43490 = ~n39956 & ~n43489;
  assign n43491 = i_RtoB_ACK0 & ~n43490;
  assign n43492 = ~n43271 & ~n43491;
  assign n43493 = controllable_DEQ & ~n43492;
  assign n43494 = ~n11681 & ~n39964;
  assign n43495 = i_RtoB_ACK0 & ~n43494;
  assign n43496 = ~n17993 & ~n39117;
  assign n43497 = ~i_RtoB_ACK0 & ~n43496;
  assign n43498 = ~n43495 & ~n43497;
  assign n43499 = ~controllable_DEQ & ~n43498;
  assign n43500 = ~n43493 & ~n43499;
  assign n43501 = i_FULL & ~n43500;
  assign n43502 = ~n43277 & ~n43491;
  assign n43503 = controllable_DEQ & ~n43502;
  assign n43504 = ~n18028 & ~n39133;
  assign n43505 = ~i_RtoB_ACK0 & ~n43504;
  assign n43506 = ~n43495 & ~n43505;
  assign n43507 = ~controllable_DEQ & ~n43506;
  assign n43508 = ~n43503 & ~n43507;
  assign n43509 = ~i_FULL & ~n43508;
  assign n43510 = ~n43501 & ~n43509;
  assign n43511 = i_nEMPTY & ~n43510;
  assign n43512 = ~n39985 & ~n43285;
  assign n43513 = controllable_DEQ & ~n43512;
  assign n43514 = ~n11652 & ~n39991;
  assign n43515 = i_RtoB_ACK0 & ~n43514;
  assign n43516 = ~n18065 & ~n39152;
  assign n43517 = ~i_RtoB_ACK0 & ~n43516;
  assign n43518 = ~n43515 & ~n43517;
  assign n43519 = ~controllable_DEQ & ~n43518;
  assign n43520 = ~n43513 & ~n43519;
  assign n43521 = i_FULL & ~n43520;
  assign n43522 = ~n40004 & ~n43291;
  assign n43523 = controllable_DEQ & ~n43522;
  assign n43524 = ~n11652 & ~n40011;
  assign n43525 = i_RtoB_ACK0 & ~n43524;
  assign n43526 = ~n11758 & ~n37552;
  assign n43527 = ~controllable_BtoR_REQ0 & ~n43526;
  assign n43528 = ~n17974 & ~n43527;
  assign n43529 = ~i_RtoB_ACK0 & ~n43528;
  assign n43530 = ~n43525 & ~n43529;
  assign n43531 = ~controllable_DEQ & ~n43530;
  assign n43532 = ~n43523 & ~n43531;
  assign n43533 = ~i_FULL & ~n43532;
  assign n43534 = ~n43521 & ~n43533;
  assign n43535 = ~i_nEMPTY & ~n43534;
  assign n43536 = ~n43511 & ~n43535;
  assign n43537 = controllable_BtoS_ACK0 & ~n43536;
  assign n43538 = ~n11797 & ~n37680;
  assign n43539 = ~controllable_BtoR_REQ0 & ~n43538;
  assign n43540 = ~n40026 & ~n43539;
  assign n43541 = i_RtoB_ACK0 & ~n43540;
  assign n43542 = ~n43301 & ~n43541;
  assign n43543 = controllable_DEQ & ~n43542;
  assign n43544 = ~n11828 & ~n40034;
  assign n43545 = i_RtoB_ACK0 & ~n43544;
  assign n43546 = ~n18135 & ~n39190;
  assign n43547 = ~i_RtoB_ACK0 & ~n43546;
  assign n43548 = ~n43545 & ~n43547;
  assign n43549 = ~controllable_DEQ & ~n43548;
  assign n43550 = ~n43543 & ~n43549;
  assign n43551 = i_FULL & ~n43550;
  assign n43552 = ~n43307 & ~n43541;
  assign n43553 = controllable_DEQ & ~n43552;
  assign n43554 = ~n18170 & ~n39206;
  assign n43555 = ~i_RtoB_ACK0 & ~n43554;
  assign n43556 = ~n43545 & ~n43555;
  assign n43557 = ~controllable_DEQ & ~n43556;
  assign n43558 = ~n43553 & ~n43557;
  assign n43559 = ~i_FULL & ~n43558;
  assign n43560 = ~n43551 & ~n43559;
  assign n43561 = i_nEMPTY & ~n43560;
  assign n43562 = ~n40055 & ~n43315;
  assign n43563 = controllable_DEQ & ~n43562;
  assign n43564 = ~n11799 & ~n40061;
  assign n43565 = i_RtoB_ACK0 & ~n43564;
  assign n43566 = ~n18207 & ~n39225;
  assign n43567 = ~i_RtoB_ACK0 & ~n43566;
  assign n43568 = ~n43565 & ~n43567;
  assign n43569 = ~controllable_DEQ & ~n43568;
  assign n43570 = ~n43563 & ~n43569;
  assign n43571 = i_FULL & ~n43570;
  assign n43572 = ~n40074 & ~n43321;
  assign n43573 = controllable_DEQ & ~n43572;
  assign n43574 = ~n11799 & ~n40081;
  assign n43575 = i_RtoB_ACK0 & ~n43574;
  assign n43576 = ~n11905 & ~n37815;
  assign n43577 = ~controllable_BtoR_REQ0 & ~n43576;
  assign n43578 = ~n18116 & ~n43577;
  assign n43579 = ~i_RtoB_ACK0 & ~n43578;
  assign n43580 = ~n43575 & ~n43579;
  assign n43581 = ~controllable_DEQ & ~n43580;
  assign n43582 = ~n43573 & ~n43581;
  assign n43583 = ~i_FULL & ~n43582;
  assign n43584 = ~n43571 & ~n43583;
  assign n43585 = ~i_nEMPTY & ~n43584;
  assign n43586 = ~n43561 & ~n43585;
  assign n43587 = ~controllable_BtoS_ACK0 & ~n43586;
  assign n43588 = ~n43537 & ~n43587;
  assign n43589 = n4465 & ~n43588;
  assign n43590 = ~n7242 & ~n37844;
  assign n43591 = ~controllable_BtoR_REQ0 & ~n43590;
  assign n43592 = ~n40097 & ~n43591;
  assign n43593 = i_RtoB_ACK0 & ~n43592;
  assign n43594 = ~n42565 & ~n43593;
  assign n43595 = controllable_DEQ & ~n43594;
  assign n43596 = ~n24351 & ~n43595;
  assign n43597 = i_FULL & ~n43596;
  assign n43598 = ~n42571 & ~n43593;
  assign n43599 = controllable_DEQ & ~n43598;
  assign n43600 = ~n24361 & ~n43599;
  assign n43601 = ~i_FULL & ~n43600;
  assign n43602 = ~n43597 & ~n43601;
  assign n43603 = i_nEMPTY & ~n43602;
  assign n43604 = ~n42591 & ~n43603;
  assign n43605 = ~controllable_BtoS_ACK0 & ~n43604;
  assign n43606 = ~n25759 & ~n43605;
  assign n43607 = ~n4465 & ~n43606;
  assign n43608 = ~n43589 & ~n43607;
  assign n43609 = ~i_StoB_REQ10 & ~n43608;
  assign n43610 = ~n43487 & ~n43609;
  assign n43611 = controllable_BtoS_ACK10 & ~n43610;
  assign n43612 = ~n11650 & ~n37902;
  assign n43613 = ~controllable_BtoR_REQ0 & ~n43612;
  assign n43614 = ~n40132 & ~n43613;
  assign n43615 = i_RtoB_ACK0 & ~n43614;
  assign n43616 = ~n11668 & ~n37908;
  assign n43617 = ~controllable_BtoR_REQ0 & ~n43616;
  assign n43618 = ~n40928 & ~n43617;
  assign n43619 = ~i_RtoB_ACK0 & ~n43618;
  assign n43620 = ~n43615 & ~n43619;
  assign n43621 = controllable_DEQ & ~n43620;
  assign n43622 = ~n42611 & ~n43621;
  assign n43623 = i_FULL & ~n43622;
  assign n43624 = ~n11703 & ~n37927;
  assign n43625 = ~controllable_BtoR_REQ0 & ~n43624;
  assign n43626 = ~n40944 & ~n43625;
  assign n43627 = ~i_RtoB_ACK0 & ~n43626;
  assign n43628 = ~n43615 & ~n43627;
  assign n43629 = controllable_DEQ & ~n43628;
  assign n43630 = ~n42621 & ~n43629;
  assign n43631 = ~i_FULL & ~n43630;
  assign n43632 = ~n43623 & ~n43631;
  assign n43633 = i_nEMPTY & ~n43632;
  assign n43634 = ~n11732 & ~n37941;
  assign n43635 = ~controllable_BtoR_REQ0 & ~n43634;
  assign n43636 = ~n40962 & ~n43635;
  assign n43637 = ~i_RtoB_ACK0 & ~n43636;
  assign n43638 = ~n40157 & ~n43637;
  assign n43639 = controllable_DEQ & ~n43638;
  assign n43640 = ~n42635 & ~n43639;
  assign n43641 = i_FULL & ~n43640;
  assign n43642 = ~n11750 & ~n37960;
  assign n43643 = ~controllable_BtoR_REQ0 & ~n43642;
  assign n43644 = ~n40978 & ~n43643;
  assign n43645 = ~i_RtoB_ACK0 & ~n43644;
  assign n43646 = ~n40171 & ~n43645;
  assign n43647 = controllable_DEQ & ~n43646;
  assign n43648 = ~n42647 & ~n43647;
  assign n43649 = ~i_FULL & ~n43648;
  assign n43650 = ~n43641 & ~n43649;
  assign n43651 = ~i_nEMPTY & ~n43650;
  assign n43652 = ~n43633 & ~n43651;
  assign n43653 = controllable_BtoS_ACK0 & ~n43652;
  assign n43654 = ~n11797 & ~n37986;
  assign n43655 = ~controllable_BtoR_REQ0 & ~n43654;
  assign n43656 = ~n40193 & ~n43655;
  assign n43657 = i_RtoB_ACK0 & ~n43656;
  assign n43658 = ~n11815 & ~n37992;
  assign n43659 = ~controllable_BtoR_REQ0 & ~n43658;
  assign n43660 = ~n40999 & ~n43659;
  assign n43661 = ~i_RtoB_ACK0 & ~n43660;
  assign n43662 = ~n43657 & ~n43661;
  assign n43663 = controllable_DEQ & ~n43662;
  assign n43664 = ~n42665 & ~n43663;
  assign n43665 = i_FULL & ~n43664;
  assign n43666 = ~n11850 & ~n38011;
  assign n43667 = ~controllable_BtoR_REQ0 & ~n43666;
  assign n43668 = ~n41015 & ~n43667;
  assign n43669 = ~i_RtoB_ACK0 & ~n43668;
  assign n43670 = ~n43657 & ~n43669;
  assign n43671 = controllable_DEQ & ~n43670;
  assign n43672 = ~n42675 & ~n43671;
  assign n43673 = ~i_FULL & ~n43672;
  assign n43674 = ~n43665 & ~n43673;
  assign n43675 = i_nEMPTY & ~n43674;
  assign n43676 = ~n11879 & ~n38025;
  assign n43677 = ~controllable_BtoR_REQ0 & ~n43676;
  assign n43678 = ~n41033 & ~n43677;
  assign n43679 = ~i_RtoB_ACK0 & ~n43678;
  assign n43680 = ~n40218 & ~n43679;
  assign n43681 = controllable_DEQ & ~n43680;
  assign n43682 = ~n42689 & ~n43681;
  assign n43683 = i_FULL & ~n43682;
  assign n43684 = ~n11897 & ~n38044;
  assign n43685 = ~controllable_BtoR_REQ0 & ~n43684;
  assign n43686 = ~n41049 & ~n43685;
  assign n43687 = ~i_RtoB_ACK0 & ~n43686;
  assign n43688 = ~n40232 & ~n43687;
  assign n43689 = controllable_DEQ & ~n43688;
  assign n43690 = ~n42701 & ~n43689;
  assign n43691 = ~i_FULL & ~n43690;
  assign n43692 = ~n43683 & ~n43691;
  assign n43693 = ~i_nEMPTY & ~n43692;
  assign n43694 = ~n43675 & ~n43693;
  assign n43695 = ~controllable_BtoS_ACK0 & ~n43694;
  assign n43696 = ~n43653 & ~n43695;
  assign n43697 = n4465 & ~n43696;
  assign n43698 = ~n7242 & ~n38072;
  assign n43699 = ~controllable_BtoR_REQ0 & ~n43698;
  assign n43700 = ~n40255 & ~n43699;
  assign n43701 = i_RtoB_ACK0 & ~n43700;
  assign n43702 = ~n42713 & ~n43701;
  assign n43703 = controllable_DEQ & ~n43702;
  assign n43704 = ~n24514 & ~n43703;
  assign n43705 = i_FULL & ~n43704;
  assign n43706 = ~n42719 & ~n43701;
  assign n43707 = controllable_DEQ & ~n43706;
  assign n43708 = ~n24524 & ~n43707;
  assign n43709 = ~i_FULL & ~n43708;
  assign n43710 = ~n43705 & ~n43709;
  assign n43711 = i_nEMPTY & ~n43710;
  assign n43712 = ~n42739 & ~n43711;
  assign n43713 = ~controllable_BtoS_ACK0 & ~n43712;
  assign n43714 = ~n24502 & ~n43713;
  assign n43715 = ~n4465 & ~n43714;
  assign n43716 = ~n43697 & ~n43715;
  assign n43717 = i_StoB_REQ10 & ~n43716;
  assign n43718 = ~n43609 & ~n43717;
  assign n43719 = ~controllable_BtoS_ACK10 & ~n43718;
  assign n43720 = ~n43611 & ~n43719;
  assign n43721 = n4464 & ~n43720;
  assign n43722 = ~n7917 & ~n38150;
  assign n43723 = ~controllable_BtoR_REQ0 & ~n43722;
  assign n43724 = ~n40292 & ~n43723;
  assign n43725 = i_RtoB_ACK0 & ~n43724;
  assign n43726 = ~n43341 & ~n43725;
  assign n43727 = controllable_DEQ & ~n43726;
  assign n43728 = ~n25777 & ~n43727;
  assign n43729 = i_FULL & ~n43728;
  assign n43730 = ~n43347 & ~n43725;
  assign n43731 = controllable_DEQ & ~n43730;
  assign n43732 = ~n25783 & ~n43731;
  assign n43733 = ~i_FULL & ~n43732;
  assign n43734 = ~n43729 & ~n43733;
  assign n43735 = i_nEMPTY & ~n43734;
  assign n43736 = ~n25791 & ~n42769;
  assign n43737 = i_FULL & ~n43736;
  assign n43738 = ~n25795 & ~n42775;
  assign n43739 = ~i_FULL & ~n43738;
  assign n43740 = ~n43737 & ~n43739;
  assign n43741 = ~i_nEMPTY & ~n43740;
  assign n43742 = ~n43735 & ~n43741;
  assign n43743 = controllable_BtoS_ACK0 & ~n43742;
  assign n43744 = ~n8084 & ~n38202;
  assign n43745 = ~controllable_BtoR_REQ0 & ~n43744;
  assign n43746 = ~n40321 & ~n43745;
  assign n43747 = i_RtoB_ACK0 & ~n43746;
  assign n43748 = ~n43363 & ~n43747;
  assign n43749 = controllable_DEQ & ~n43748;
  assign n43750 = ~n25809 & ~n43749;
  assign n43751 = i_FULL & ~n43750;
  assign n43752 = ~n43369 & ~n43747;
  assign n43753 = controllable_DEQ & ~n43752;
  assign n43754 = ~n25815 & ~n43753;
  assign n43755 = ~i_FULL & ~n43754;
  assign n43756 = ~n43751 & ~n43755;
  assign n43757 = i_nEMPTY & ~n43756;
  assign n43758 = ~n25823 & ~n42801;
  assign n43759 = i_FULL & ~n43758;
  assign n43760 = ~n25827 & ~n42807;
  assign n43761 = ~i_FULL & ~n43760;
  assign n43762 = ~n43759 & ~n43761;
  assign n43763 = ~i_nEMPTY & ~n43762;
  assign n43764 = ~n43757 & ~n43763;
  assign n43765 = ~controllable_BtoS_ACK0 & ~n43764;
  assign n43766 = ~n43743 & ~n43765;
  assign n43767 = n4465 & ~n43766;
  assign n43768 = ~n8327 & ~n38256;
  assign n43769 = ~controllable_BtoR_REQ0 & ~n43768;
  assign n43770 = ~n40351 & ~n43769;
  assign n43771 = i_RtoB_ACK0 & ~n43770;
  assign n43772 = ~n42819 & ~n43771;
  assign n43773 = controllable_DEQ & ~n43772;
  assign n43774 = ~n24743 & ~n43773;
  assign n43775 = i_FULL & ~n43774;
  assign n43776 = ~n42825 & ~n43771;
  assign n43777 = controllable_DEQ & ~n43776;
  assign n43778 = ~n24753 & ~n43777;
  assign n43779 = ~i_FULL & ~n43778;
  assign n43780 = ~n43775 & ~n43779;
  assign n43781 = i_nEMPTY & ~n43780;
  assign n43782 = ~n42845 & ~n43781;
  assign n43783 = ~controllable_BtoS_ACK0 & ~n43782;
  assign n43784 = ~n24731 & ~n43783;
  assign n43785 = ~n4465 & ~n43784;
  assign n43786 = ~n43767 & ~n43785;
  assign n43787 = ~i_StoB_REQ10 & ~n43786;
  assign n43788 = ~n24609 & ~n43787;
  assign n43789 = controllable_BtoS_ACK10 & ~n43788;
  assign n43790 = ~n7917 & ~n38314;
  assign n43791 = ~controllable_BtoR_REQ0 & ~n43790;
  assign n43792 = ~n40385 & ~n43791;
  assign n43793 = i_RtoB_ACK0 & ~n43792;
  assign n43794 = ~n42857 & ~n43793;
  assign n43795 = controllable_DEQ & ~n43794;
  assign n43796 = ~n24793 & ~n43795;
  assign n43797 = i_FULL & ~n43796;
  assign n43798 = ~n42863 & ~n43793;
  assign n43799 = controllable_DEQ & ~n43798;
  assign n43800 = ~n24803 & ~n43799;
  assign n43801 = ~i_FULL & ~n43800;
  assign n43802 = ~n43797 & ~n43801;
  assign n43803 = i_nEMPTY & ~n43802;
  assign n43804 = ~n42883 & ~n43803;
  assign n43805 = controllable_BtoS_ACK0 & ~n43804;
  assign n43806 = ~n8084 & ~n38366;
  assign n43807 = ~controllable_BtoR_REQ0 & ~n43806;
  assign n43808 = ~n40413 & ~n43807;
  assign n43809 = i_RtoB_ACK0 & ~n43808;
  assign n43810 = ~n42889 & ~n43809;
  assign n43811 = controllable_DEQ & ~n43810;
  assign n43812 = ~n24834 & ~n43811;
  assign n43813 = i_FULL & ~n43812;
  assign n43814 = ~n42895 & ~n43809;
  assign n43815 = controllable_DEQ & ~n43814;
  assign n43816 = ~n24844 & ~n43815;
  assign n43817 = ~i_FULL & ~n43816;
  assign n43818 = ~n43813 & ~n43817;
  assign n43819 = i_nEMPTY & ~n43818;
  assign n43820 = ~n42915 & ~n43819;
  assign n43821 = ~controllable_BtoS_ACK0 & ~n43820;
  assign n43822 = ~n43805 & ~n43821;
  assign n43823 = n4465 & ~n43822;
  assign n43824 = ~n8327 & ~n38420;
  assign n43825 = ~controllable_BtoR_REQ0 & ~n43824;
  assign n43826 = ~n40443 & ~n43825;
  assign n43827 = i_RtoB_ACK0 & ~n43826;
  assign n43828 = ~n42923 & ~n43827;
  assign n43829 = controllable_DEQ & ~n43828;
  assign n43830 = ~n24906 & ~n43829;
  assign n43831 = i_FULL & ~n43830;
  assign n43832 = ~n42929 & ~n43827;
  assign n43833 = controllable_DEQ & ~n43832;
  assign n43834 = ~n24916 & ~n43833;
  assign n43835 = ~i_FULL & ~n43834;
  assign n43836 = ~n43831 & ~n43835;
  assign n43837 = i_nEMPTY & ~n43836;
  assign n43838 = ~n42949 & ~n43837;
  assign n43839 = ~controllable_BtoS_ACK0 & ~n43838;
  assign n43840 = ~n24894 & ~n43839;
  assign n43841 = ~n4465 & ~n43840;
  assign n43842 = ~n43823 & ~n43841;
  assign n43843 = i_StoB_REQ10 & ~n43842;
  assign n43844 = ~n43787 & ~n43843;
  assign n43845 = ~controllable_BtoS_ACK10 & ~n43844;
  assign n43846 = ~n43789 & ~n43845;
  assign n43847 = ~n4464 & ~n43846;
  assign n43848 = ~n43721 & ~n43847;
  assign n43849 = ~n4463 & ~n43848;
  assign n43850 = ~n41589 & ~n43849;
  assign n43851 = n4462 & ~n43850;
  assign n43852 = ~n40483 & ~n43489;
  assign n43853 = i_RtoB_ACK0 & ~n43852;
  assign n43854 = ~n43271 & ~n43853;
  assign n43855 = controllable_DEQ & ~n43854;
  assign n43856 = ~n25285 & ~n43855;
  assign n43857 = i_FULL & ~n43856;
  assign n43858 = ~n43277 & ~n43853;
  assign n43859 = controllable_DEQ & ~n43858;
  assign n43860 = ~n25295 & ~n43859;
  assign n43861 = ~i_FULL & ~n43860;
  assign n43862 = ~n43857 & ~n43861;
  assign n43863 = i_nEMPTY & ~n43862;
  assign n43864 = ~n43297 & ~n43863;
  assign n43865 = controllable_BtoS_ACK0 & ~n43864;
  assign n43866 = ~n40511 & ~n43539;
  assign n43867 = i_RtoB_ACK0 & ~n43866;
  assign n43868 = ~n43301 & ~n43867;
  assign n43869 = controllable_DEQ & ~n43868;
  assign n43870 = ~n25329 & ~n43869;
  assign n43871 = i_FULL & ~n43870;
  assign n43872 = ~n43307 & ~n43867;
  assign n43873 = controllable_DEQ & ~n43872;
  assign n43874 = ~n25339 & ~n43873;
  assign n43875 = ~i_FULL & ~n43874;
  assign n43876 = ~n43871 & ~n43875;
  assign n43877 = i_nEMPTY & ~n43876;
  assign n43878 = ~n43327 & ~n43877;
  assign n43879 = ~controllable_BtoS_ACK0 & ~n43878;
  assign n43880 = ~n43865 & ~n43879;
  assign n43881 = n4465 & ~n43880;
  assign n43882 = ~n25389 & ~n43605;
  assign n43883 = ~n4465 & ~n43882;
  assign n43884 = ~n43881 & ~n43883;
  assign n43885 = ~i_StoB_REQ10 & ~n43884;
  assign n43886 = ~n25273 & ~n43885;
  assign n43887 = ~controllable_BtoS_ACK10 & ~n43886;
  assign n43888 = ~n25913 & ~n43887;
  assign n43889 = n4464 & ~n43888;
  assign n43890 = ~n40549 & ~n43723;
  assign n43891 = i_RtoB_ACK0 & ~n43890;
  assign n43892 = ~n43341 & ~n43891;
  assign n43893 = controllable_DEQ & ~n43892;
  assign n43894 = ~n25495 & ~n43893;
  assign n43895 = i_FULL & ~n43894;
  assign n43896 = ~n43347 & ~n43891;
  assign n43897 = controllable_DEQ & ~n43896;
  assign n43898 = ~n25505 & ~n43897;
  assign n43899 = ~i_FULL & ~n43898;
  assign n43900 = ~n43895 & ~n43899;
  assign n43901 = i_nEMPTY & ~n43900;
  assign n43902 = ~n43359 & ~n43901;
  assign n43903 = controllable_BtoS_ACK0 & ~n43902;
  assign n43904 = ~n40573 & ~n43745;
  assign n43905 = i_RtoB_ACK0 & ~n43904;
  assign n43906 = ~n43363 & ~n43905;
  assign n43907 = controllable_DEQ & ~n43906;
  assign n43908 = ~n25533 & ~n43907;
  assign n43909 = i_FULL & ~n43908;
  assign n43910 = ~n43369 & ~n43905;
  assign n43911 = controllable_DEQ & ~n43910;
  assign n43912 = ~n25543 & ~n43911;
  assign n43913 = ~i_FULL & ~n43912;
  assign n43914 = ~n43909 & ~n43913;
  assign n43915 = i_nEMPTY & ~n43914;
  assign n43916 = ~n43381 & ~n43915;
  assign n43917 = ~controllable_BtoS_ACK0 & ~n43916;
  assign n43918 = ~n43903 & ~n43917;
  assign n43919 = n4465 & ~n43918;
  assign n43920 = ~n43785 & ~n43919;
  assign n43921 = ~i_StoB_REQ10 & ~n43920;
  assign n43922 = ~n25487 & ~n43921;
  assign n43923 = ~controllable_BtoS_ACK10 & ~n43922;
  assign n43924 = ~n25399 & ~n43923;
  assign n43925 = ~n4464 & ~n43924;
  assign n43926 = ~n43889 & ~n43925;
  assign n43927 = ~n4463 & ~n43926;
  assign n43928 = ~n23523 & ~n43927;
  assign n43929 = ~n4462 & ~n43928;
  assign n43930 = ~n43851 & ~n43929;
  assign n43931 = n4461 & ~n43930;
  assign n43932 = ~controllable_BtoR_REQ0 & ~n36887;
  assign n43933 = ~n17562 & ~n43932;
  assign n43934 = ~i_RtoB_ACK0 & ~n43933;
  assign n43935 = ~n42405 & ~n43934;
  assign n43936 = ~controllable_DEQ & ~n43935;
  assign n43937 = ~n27153 & ~n43936;
  assign n43938 = i_FULL & ~n43937;
  assign n43939 = ~n36888 & ~n40618;
  assign n43940 = ~controllable_BtoR_REQ0 & ~n43939;
  assign n43941 = ~n17562 & ~n43940;
  assign n43942 = ~i_RtoB_ACK0 & ~n43941;
  assign n43943 = ~n42405 & ~n43942;
  assign n43944 = ~controllable_DEQ & ~n43943;
  assign n43945 = ~n27153 & ~n43944;
  assign n43946 = ~i_FULL & ~n43945;
  assign n43947 = ~n43938 & ~n43946;
  assign n43948 = i_nEMPTY & ~n43947;
  assign n43949 = ~controllable_BtoR_REQ0 & ~n36922;
  assign n43950 = ~n17581 & ~n43949;
  assign n43951 = ~i_RtoB_ACK0 & ~n43950;
  assign n43952 = ~n42411 & ~n43951;
  assign n43953 = ~controllable_DEQ & ~n43952;
  assign n43954 = ~n23541 & ~n43953;
  assign n43955 = i_FULL & ~n43954;
  assign n43956 = ~n36933 & ~n40639;
  assign n43957 = ~controllable_BtoR_REQ0 & ~n43956;
  assign n43958 = ~n17545 & ~n43957;
  assign n43959 = ~i_RtoB_ACK0 & ~n43958;
  assign n43960 = ~n42411 & ~n43959;
  assign n43961 = ~controllable_DEQ & ~n43960;
  assign n43962 = ~n23551 & ~n43961;
  assign n43963 = ~i_FULL & ~n43962;
  assign n43964 = ~n43955 & ~n43963;
  assign n43965 = ~i_nEMPTY & ~n43964;
  assign n43966 = ~n43948 & ~n43965;
  assign n43967 = controllable_BtoS_ACK0 & ~n43966;
  assign n43968 = ~controllable_BtoR_REQ0 & ~n37068;
  assign n43969 = ~n14841 & ~n43968;
  assign n43970 = ~i_RtoB_ACK0 & ~n43969;
  assign n43971 = ~n42427 & ~n43970;
  assign n43972 = ~controllable_DEQ & ~n43971;
  assign n43973 = ~n27187 & ~n43972;
  assign n43974 = i_FULL & ~n43973;
  assign n43975 = ~n37069 & ~n40662;
  assign n43976 = ~controllable_BtoR_REQ0 & ~n43975;
  assign n43977 = ~n14841 & ~n43976;
  assign n43978 = ~i_RtoB_ACK0 & ~n43977;
  assign n43979 = ~n42427 & ~n43978;
  assign n43980 = ~controllable_DEQ & ~n43979;
  assign n43981 = ~n27187 & ~n43980;
  assign n43982 = ~i_FULL & ~n43981;
  assign n43983 = ~n43974 & ~n43982;
  assign n43984 = i_nEMPTY & ~n43983;
  assign n43985 = ~controllable_BtoR_REQ0 & ~n37103;
  assign n43986 = ~n14860 & ~n43985;
  assign n43987 = ~i_RtoB_ACK0 & ~n43986;
  assign n43988 = ~n42433 & ~n43987;
  assign n43989 = ~controllable_DEQ & ~n43988;
  assign n43990 = ~n23579 & ~n43989;
  assign n43991 = i_FULL & ~n43990;
  assign n43992 = ~n37114 & ~n40683;
  assign n43993 = ~controllable_BtoR_REQ0 & ~n43992;
  assign n43994 = ~n14824 & ~n43993;
  assign n43995 = ~i_RtoB_ACK0 & ~n43994;
  assign n43996 = ~n42433 & ~n43995;
  assign n43997 = ~controllable_DEQ & ~n43996;
  assign n43998 = ~n23589 & ~n43997;
  assign n43999 = ~i_FULL & ~n43998;
  assign n44000 = ~n43991 & ~n43999;
  assign n44001 = ~i_nEMPTY & ~n44000;
  assign n44002 = ~n43984 & ~n44001;
  assign n44003 = ~controllable_BtoS_ACK0 & ~n44002;
  assign n44004 = ~n43967 & ~n44003;
  assign n44005 = n4465 & ~n44004;
  assign n44006 = ~n26030 & ~n26038;
  assign n44007 = i_FULL & ~n44006;
  assign n44008 = ~n26046 & ~n44007;
  assign n44009 = i_nEMPTY & ~n44008;
  assign n44010 = ~n26065 & ~n44009;
  assign n44011 = ~controllable_BtoS_ACK0 & ~n44010;
  assign n44012 = ~n21013 & ~n44011;
  assign n44013 = ~n4465 & ~n44012;
  assign n44014 = ~n44005 & ~n44013;
  assign n44015 = i_StoB_REQ10 & ~n44014;
  assign n44016 = ~n38881 & ~n40712;
  assign n44017 = ~controllable_BtoR_REQ0 & ~n44016;
  assign n44018 = ~n17974 & ~n44017;
  assign n44019 = ~i_RtoB_ACK0 & ~n44018;
  assign n44020 = ~n42453 & ~n44019;
  assign n44021 = controllable_DEQ & ~n44020;
  assign n44022 = ~n38890 & ~n40726;
  assign n44023 = ~controllable_BtoR_REQ0 & ~n44022;
  assign n44024 = ~n17993 & ~n44023;
  assign n44025 = ~i_RtoB_ACK0 & ~n44024;
  assign n44026 = ~n42459 & ~n44025;
  assign n44027 = ~controllable_DEQ & ~n44026;
  assign n44028 = ~n44021 & ~n44027;
  assign n44029 = i_FULL & ~n44028;
  assign n44030 = ~n38900 & ~n40712;
  assign n44031 = ~controllable_BtoR_REQ0 & ~n44030;
  assign n44032 = ~n18012 & ~n44031;
  assign n44033 = ~i_RtoB_ACK0 & ~n44032;
  assign n44034 = ~n42453 & ~n44033;
  assign n44035 = controllable_DEQ & ~n44034;
  assign n44036 = ~n38908 & ~n40740;
  assign n44037 = ~controllable_BtoR_REQ0 & ~n44036;
  assign n44038 = ~n18028 & ~n44037;
  assign n44039 = ~i_RtoB_ACK0 & ~n44038;
  assign n44040 = ~n42459 & ~n44039;
  assign n44041 = ~controllable_DEQ & ~n44040;
  assign n44042 = ~n44035 & ~n44041;
  assign n44043 = ~i_FULL & ~n44042;
  assign n44044 = ~n44029 & ~n44043;
  assign n44045 = i_nEMPTY & ~n44044;
  assign n44046 = ~n37509 & ~n38922;
  assign n44047 = ~controllable_BtoR_REQ0 & ~n44046;
  assign n44048 = ~n18049 & ~n44047;
  assign n44049 = ~i_RtoB_ACK0 & ~n44048;
  assign n44050 = ~n15217 & ~n44049;
  assign n44051 = controllable_DEQ & ~n44050;
  assign n44052 = ~n38931 & ~n40764;
  assign n44053 = ~controllable_BtoR_REQ0 & ~n44052;
  assign n44054 = ~n18065 & ~n44053;
  assign n44055 = ~i_RtoB_ACK0 & ~n44054;
  assign n44056 = ~n42483 & ~n44055;
  assign n44057 = ~controllable_DEQ & ~n44056;
  assign n44058 = ~n44051 & ~n44057;
  assign n44059 = i_FULL & ~n44058;
  assign n44060 = ~n37542 & ~n38942;
  assign n44061 = ~controllable_BtoR_REQ0 & ~n44060;
  assign n44062 = ~n18084 & ~n44061;
  assign n44063 = ~i_RtoB_ACK0 & ~n44062;
  assign n44064 = ~n15245 & ~n44063;
  assign n44065 = controllable_DEQ & ~n44064;
  assign n44066 = ~n38952 & ~n40787;
  assign n44067 = ~controllable_BtoR_REQ0 & ~n44066;
  assign n44068 = ~n17974 & ~n44067;
  assign n44069 = ~i_RtoB_ACK0 & ~n44068;
  assign n44070 = ~n42495 & ~n44069;
  assign n44071 = ~controllable_DEQ & ~n44070;
  assign n44072 = ~n44065 & ~n44071;
  assign n44073 = ~i_FULL & ~n44072;
  assign n44074 = ~n44059 & ~n44073;
  assign n44075 = ~i_nEMPTY & ~n44074;
  assign n44076 = ~n44045 & ~n44075;
  assign n44077 = controllable_BtoS_ACK0 & ~n44076;
  assign n44078 = ~n38976 & ~n40804;
  assign n44079 = ~controllable_BtoR_REQ0 & ~n44078;
  assign n44080 = ~n18116 & ~n44079;
  assign n44081 = ~i_RtoB_ACK0 & ~n44080;
  assign n44082 = ~n42507 & ~n44081;
  assign n44083 = controllable_DEQ & ~n44082;
  assign n44084 = ~n38985 & ~n40818;
  assign n44085 = ~controllable_BtoR_REQ0 & ~n44084;
  assign n44086 = ~n18135 & ~n44085;
  assign n44087 = ~i_RtoB_ACK0 & ~n44086;
  assign n44088 = ~n42513 & ~n44087;
  assign n44089 = ~controllable_DEQ & ~n44088;
  assign n44090 = ~n44083 & ~n44089;
  assign n44091 = i_FULL & ~n44090;
  assign n44092 = ~n38995 & ~n40804;
  assign n44093 = ~controllable_BtoR_REQ0 & ~n44092;
  assign n44094 = ~n18154 & ~n44093;
  assign n44095 = ~i_RtoB_ACK0 & ~n44094;
  assign n44096 = ~n42507 & ~n44095;
  assign n44097 = controllable_DEQ & ~n44096;
  assign n44098 = ~n39003 & ~n40832;
  assign n44099 = ~controllable_BtoR_REQ0 & ~n44098;
  assign n44100 = ~n18170 & ~n44099;
  assign n44101 = ~i_RtoB_ACK0 & ~n44100;
  assign n44102 = ~n42513 & ~n44101;
  assign n44103 = ~controllable_DEQ & ~n44102;
  assign n44104 = ~n44097 & ~n44103;
  assign n44105 = ~i_FULL & ~n44104;
  assign n44106 = ~n44091 & ~n44105;
  assign n44107 = i_nEMPTY & ~n44106;
  assign n44108 = ~n37772 & ~n39017;
  assign n44109 = ~controllable_BtoR_REQ0 & ~n44108;
  assign n44110 = ~n18191 & ~n44109;
  assign n44111 = ~i_RtoB_ACK0 & ~n44110;
  assign n44112 = ~n17731 & ~n44111;
  assign n44113 = controllable_DEQ & ~n44112;
  assign n44114 = ~n39026 & ~n40856;
  assign n44115 = ~controllable_BtoR_REQ0 & ~n44114;
  assign n44116 = ~n18207 & ~n44115;
  assign n44117 = ~i_RtoB_ACK0 & ~n44116;
  assign n44118 = ~n42537 & ~n44117;
  assign n44119 = ~controllable_DEQ & ~n44118;
  assign n44120 = ~n44113 & ~n44119;
  assign n44121 = i_FULL & ~n44120;
  assign n44122 = ~n37805 & ~n39037;
  assign n44123 = ~controllable_BtoR_REQ0 & ~n44122;
  assign n44124 = ~n18226 & ~n44123;
  assign n44125 = ~i_RtoB_ACK0 & ~n44124;
  assign n44126 = ~n17764 & ~n44125;
  assign n44127 = controllable_DEQ & ~n44126;
  assign n44128 = ~n39047 & ~n40879;
  assign n44129 = ~controllable_BtoR_REQ0 & ~n44128;
  assign n44130 = ~n18116 & ~n44129;
  assign n44131 = ~i_RtoB_ACK0 & ~n44130;
  assign n44132 = ~n42549 & ~n44131;
  assign n44133 = ~controllable_DEQ & ~n44132;
  assign n44134 = ~n44127 & ~n44133;
  assign n44135 = ~i_FULL & ~n44134;
  assign n44136 = ~n44121 & ~n44135;
  assign n44137 = ~i_nEMPTY & ~n44136;
  assign n44138 = ~n44107 & ~n44137;
  assign n44139 = ~controllable_BtoS_ACK0 & ~n44138;
  assign n44140 = ~n44077 & ~n44139;
  assign n44141 = n4465 & ~n44140;
  assign n44142 = ~n11317 & ~n37850;
  assign n44143 = ~controllable_BtoR_REQ0 & ~n44142;
  assign n44144 = ~n15281 & ~n44143;
  assign n44145 = ~i_RtoB_ACK0 & ~n44144;
  assign n44146 = ~n42563 & ~n44145;
  assign n44147 = controllable_DEQ & ~n44146;
  assign n44148 = ~n26219 & ~n44147;
  assign n44149 = i_FULL & ~n44148;
  assign n44150 = ~n11317 & ~n37860;
  assign n44151 = ~controllable_BtoR_REQ0 & ~n44150;
  assign n44152 = ~n15319 & ~n44151;
  assign n44153 = ~i_RtoB_ACK0 & ~n44152;
  assign n44154 = ~n42563 & ~n44153;
  assign n44155 = controllable_DEQ & ~n44154;
  assign n44156 = ~n26233 & ~n44155;
  assign n44157 = ~i_FULL & ~n44156;
  assign n44158 = ~n44149 & ~n44157;
  assign n44159 = i_nEMPTY & ~n44158;
  assign n44160 = ~n26243 & ~n41799;
  assign n44161 = i_FULL & ~n44160;
  assign n44162 = ~n26251 & ~n41805;
  assign n44163 = ~i_FULL & ~n44162;
  assign n44164 = ~n44161 & ~n44163;
  assign n44165 = ~i_nEMPTY & ~n44164;
  assign n44166 = ~n44159 & ~n44165;
  assign n44167 = ~controllable_BtoS_ACK0 & ~n44166;
  assign n44168 = ~n26207 & ~n44167;
  assign n44169 = ~n4465 & ~n44168;
  assign n44170 = ~n44141 & ~n44169;
  assign n44171 = ~i_StoB_REQ10 & ~n44170;
  assign n44172 = ~n44015 & ~n44171;
  assign n44173 = controllable_BtoS_ACK10 & ~n44172;
  assign n44174 = ~n11238 & ~n39109;
  assign n44175 = ~controllable_BtoR_REQ0 & ~n44174;
  assign n44176 = ~n40928 & ~n44175;
  assign n44177 = ~i_RtoB_ACK0 & ~n44176;
  assign n44178 = ~n42601 & ~n44177;
  assign n44179 = controllable_DEQ & ~n44178;
  assign n44180 = ~n37470 & ~n40935;
  assign n44181 = ~controllable_BtoR_REQ0 & ~n44180;
  assign n44182 = ~n40933 & ~n44181;
  assign n44183 = ~i_RtoB_ACK0 & ~n44182;
  assign n44184 = ~n42607 & ~n44183;
  assign n44185 = ~controllable_DEQ & ~n44184;
  assign n44186 = ~n44179 & ~n44185;
  assign n44187 = i_FULL & ~n44186;
  assign n44188 = ~n11238 & ~n39125;
  assign n44189 = ~controllable_BtoR_REQ0 & ~n44188;
  assign n44190 = ~n40944 & ~n44189;
  assign n44191 = ~i_RtoB_ACK0 & ~n44190;
  assign n44192 = ~n42601 & ~n44191;
  assign n44193 = controllable_DEQ & ~n44192;
  assign n44194 = ~n37488 & ~n40951;
  assign n44195 = ~controllable_BtoR_REQ0 & ~n44194;
  assign n44196 = ~n40949 & ~n44195;
  assign n44197 = ~i_RtoB_ACK0 & ~n44196;
  assign n44198 = ~n42607 & ~n44197;
  assign n44199 = ~controllable_DEQ & ~n44198;
  assign n44200 = ~n44193 & ~n44199;
  assign n44201 = ~i_FULL & ~n44200;
  assign n44202 = ~n44187 & ~n44201;
  assign n44203 = i_nEMPTY & ~n44202;
  assign n44204 = ~n10049 & ~n39144;
  assign n44205 = ~controllable_BtoR_REQ0 & ~n44204;
  assign n44206 = ~n40962 & ~n44205;
  assign n44207 = ~i_RtoB_ACK0 & ~n44206;
  assign n44208 = ~n15604 & ~n44207;
  assign n44209 = controllable_DEQ & ~n44208;
  assign n44210 = ~n37529 & ~n40969;
  assign n44211 = ~controllable_BtoR_REQ0 & ~n44210;
  assign n44212 = ~n40967 & ~n44211;
  assign n44213 = ~i_RtoB_ACK0 & ~n44212;
  assign n44214 = ~n42631 & ~n44213;
  assign n44215 = ~controllable_DEQ & ~n44214;
  assign n44216 = ~n44209 & ~n44215;
  assign n44217 = i_FULL & ~n44216;
  assign n44218 = ~n10061 & ~n39160;
  assign n44219 = ~controllable_BtoR_REQ0 & ~n44218;
  assign n44220 = ~n40978 & ~n44219;
  assign n44221 = ~i_RtoB_ACK0 & ~n44220;
  assign n44222 = ~n15619 & ~n44221;
  assign n44223 = controllable_DEQ & ~n44222;
  assign n44224 = ~n37970 & ~n40984;
  assign n44225 = ~controllable_BtoR_REQ0 & ~n44224;
  assign n44226 = ~n40928 & ~n44225;
  assign n44227 = ~i_RtoB_ACK0 & ~n44226;
  assign n44228 = ~n42643 & ~n44227;
  assign n44229 = ~controllable_DEQ & ~n44228;
  assign n44230 = ~n44223 & ~n44229;
  assign n44231 = ~i_FULL & ~n44230;
  assign n44232 = ~n44217 & ~n44231;
  assign n44233 = ~i_nEMPTY & ~n44232;
  assign n44234 = ~n44203 & ~n44233;
  assign n44235 = controllable_BtoS_ACK0 & ~n44234;
  assign n44236 = ~n11317 & ~n39182;
  assign n44237 = ~controllable_BtoR_REQ0 & ~n44236;
  assign n44238 = ~n40999 & ~n44237;
  assign n44239 = ~i_RtoB_ACK0 & ~n44238;
  assign n44240 = ~n42655 & ~n44239;
  assign n44241 = controllable_DEQ & ~n44240;
  assign n44242 = ~n37733 & ~n41006;
  assign n44243 = ~controllable_BtoR_REQ0 & ~n44242;
  assign n44244 = ~n41004 & ~n44243;
  assign n44245 = ~i_RtoB_ACK0 & ~n44244;
  assign n44246 = ~n42661 & ~n44245;
  assign n44247 = ~controllable_DEQ & ~n44246;
  assign n44248 = ~n44241 & ~n44247;
  assign n44249 = i_FULL & ~n44248;
  assign n44250 = ~n11317 & ~n39198;
  assign n44251 = ~controllable_BtoR_REQ0 & ~n44250;
  assign n44252 = ~n41015 & ~n44251;
  assign n44253 = ~i_RtoB_ACK0 & ~n44252;
  assign n44254 = ~n42655 & ~n44253;
  assign n44255 = controllable_DEQ & ~n44254;
  assign n44256 = ~n37751 & ~n41022;
  assign n44257 = ~controllable_BtoR_REQ0 & ~n44256;
  assign n44258 = ~n41020 & ~n44257;
  assign n44259 = ~i_RtoB_ACK0 & ~n44258;
  assign n44260 = ~n42661 & ~n44259;
  assign n44261 = ~controllable_DEQ & ~n44260;
  assign n44262 = ~n44255 & ~n44261;
  assign n44263 = ~i_FULL & ~n44262;
  assign n44264 = ~n44249 & ~n44263;
  assign n44265 = i_nEMPTY & ~n44264;
  assign n44266 = ~n9951 & ~n39217;
  assign n44267 = ~controllable_BtoR_REQ0 & ~n44266;
  assign n44268 = ~n41033 & ~n44267;
  assign n44269 = ~i_RtoB_ACK0 & ~n44268;
  assign n44270 = ~n17925 & ~n44269;
  assign n44271 = controllable_DEQ & ~n44270;
  assign n44272 = ~n37792 & ~n41040;
  assign n44273 = ~controllable_BtoR_REQ0 & ~n44272;
  assign n44274 = ~n41038 & ~n44273;
  assign n44275 = ~i_RtoB_ACK0 & ~n44274;
  assign n44276 = ~n42685 & ~n44275;
  assign n44277 = ~controllable_DEQ & ~n44276;
  assign n44278 = ~n44271 & ~n44277;
  assign n44279 = i_FULL & ~n44278;
  assign n44280 = ~n9973 & ~n39233;
  assign n44281 = ~controllable_BtoR_REQ0 & ~n44280;
  assign n44282 = ~n41049 & ~n44281;
  assign n44283 = ~i_RtoB_ACK0 & ~n44282;
  assign n44284 = ~n17943 & ~n44283;
  assign n44285 = controllable_DEQ & ~n44284;
  assign n44286 = ~n38054 & ~n41055;
  assign n44287 = ~controllable_BtoR_REQ0 & ~n44286;
  assign n44288 = ~n40999 & ~n44287;
  assign n44289 = ~i_RtoB_ACK0 & ~n44288;
  assign n44290 = ~n42697 & ~n44289;
  assign n44291 = ~controllable_DEQ & ~n44290;
  assign n44292 = ~n44285 & ~n44291;
  assign n44293 = ~i_FULL & ~n44292;
  assign n44294 = ~n44279 & ~n44293;
  assign n44295 = ~i_nEMPTY & ~n44294;
  assign n44296 = ~n44265 & ~n44295;
  assign n44297 = ~controllable_BtoS_ACK0 & ~n44296;
  assign n44298 = ~n44235 & ~n44297;
  assign n44299 = n4465 & ~n44298;
  assign n44300 = ~n11317 & ~n38078;
  assign n44301 = ~controllable_BtoR_REQ0 & ~n44300;
  assign n44302 = ~n19554 & ~n44301;
  assign n44303 = ~i_RtoB_ACK0 & ~n44302;
  assign n44304 = ~n42711 & ~n44303;
  assign n44305 = controllable_DEQ & ~n44304;
  assign n44306 = ~n26394 & ~n44305;
  assign n44307 = i_FULL & ~n44306;
  assign n44308 = ~n11317 & ~n38088;
  assign n44309 = ~controllable_BtoR_REQ0 & ~n44308;
  assign n44310 = ~n19566 & ~n44309;
  assign n44311 = ~i_RtoB_ACK0 & ~n44310;
  assign n44312 = ~n42711 & ~n44311;
  assign n44313 = controllable_DEQ & ~n44312;
  assign n44314 = ~n26406 & ~n44313;
  assign n44315 = ~i_FULL & ~n44314;
  assign n44316 = ~n44307 & ~n44315;
  assign n44317 = i_nEMPTY & ~n44316;
  assign n44318 = ~n26414 & ~n41947;
  assign n44319 = i_FULL & ~n44318;
  assign n44320 = ~n26417 & ~n41953;
  assign n44321 = ~i_FULL & ~n44320;
  assign n44322 = ~n44319 & ~n44321;
  assign n44323 = ~i_nEMPTY & ~n44322;
  assign n44324 = ~n44317 & ~n44323;
  assign n44325 = ~controllable_BtoS_ACK0 & ~n44324;
  assign n44326 = ~n26384 & ~n44325;
  assign n44327 = ~n4465 & ~n44326;
  assign n44328 = ~n44299 & ~n44327;
  assign n44329 = i_StoB_REQ10 & ~n44328;
  assign n44330 = ~n44171 & ~n44329;
  assign n44331 = ~controllable_BtoS_ACK10 & ~n44330;
  assign n44332 = ~n44173 & ~n44331;
  assign n44333 = n4464 & ~n44332;
  assign n44334 = ~n26442 & ~n26450;
  assign n44335 = i_FULL & ~n44334;
  assign n44336 = ~n26458 & ~n44335;
  assign n44337 = i_nEMPTY & ~n44336;
  assign n44338 = ~n26477 & ~n44337;
  assign n44339 = controllable_BtoS_ACK0 & ~n44338;
  assign n44340 = ~n26490 & ~n26498;
  assign n44341 = i_FULL & ~n44340;
  assign n44342 = ~n26506 & ~n44341;
  assign n44343 = i_nEMPTY & ~n44342;
  assign n44344 = ~n26525 & ~n44343;
  assign n44345 = ~controllable_BtoS_ACK0 & ~n44344;
  assign n44346 = ~n44339 & ~n44345;
  assign n44347 = n4465 & ~n44346;
  assign n44348 = ~n21013 & ~n44345;
  assign n44349 = ~n4465 & ~n44348;
  assign n44350 = ~n44347 & ~n44349;
  assign n44351 = i_StoB_REQ10 & ~n44350;
  assign n44352 = ~n19765 & ~n39303;
  assign n44353 = ~controllable_BtoR_REQ0 & ~n44352;
  assign n44354 = ~n15889 & ~n44353;
  assign n44355 = ~i_RtoB_ACK0 & ~n44354;
  assign n44356 = ~n42751 & ~n44355;
  assign n44357 = controllable_DEQ & ~n44356;
  assign n44358 = ~n26545 & ~n44357;
  assign n44359 = i_FULL & ~n44358;
  assign n44360 = ~n19765 & ~n39313;
  assign n44361 = ~controllable_BtoR_REQ0 & ~n44360;
  assign n44362 = ~n15927 & ~n44361;
  assign n44363 = ~i_RtoB_ACK0 & ~n44362;
  assign n44364 = ~n42751 & ~n44363;
  assign n44365 = controllable_DEQ & ~n44364;
  assign n44366 = ~n26559 & ~n44365;
  assign n44367 = ~i_FULL & ~n44366;
  assign n44368 = ~n44359 & ~n44367;
  assign n44369 = i_nEMPTY & ~n44368;
  assign n44370 = ~n26569 & ~n42005;
  assign n44371 = i_FULL & ~n44370;
  assign n44372 = ~n26577 & ~n42011;
  assign n44373 = ~i_FULL & ~n44372;
  assign n44374 = ~n44371 & ~n44373;
  assign n44375 = ~i_nEMPTY & ~n44374;
  assign n44376 = ~n44369 & ~n44375;
  assign n44377 = controllable_BtoS_ACK0 & ~n44376;
  assign n44378 = ~n19839 & ~n39347;
  assign n44379 = ~controllable_BtoR_REQ0 & ~n44378;
  assign n44380 = ~n16031 & ~n44379;
  assign n44381 = ~i_RtoB_ACK0 & ~n44380;
  assign n44382 = ~n42783 & ~n44381;
  assign n44383 = controllable_DEQ & ~n44382;
  assign n44384 = ~n26595 & ~n44383;
  assign n44385 = i_FULL & ~n44384;
  assign n44386 = ~n19839 & ~n39357;
  assign n44387 = ~controllable_BtoR_REQ0 & ~n44386;
  assign n44388 = ~n16069 & ~n44387;
  assign n44389 = ~i_RtoB_ACK0 & ~n44388;
  assign n44390 = ~n42783 & ~n44389;
  assign n44391 = controllable_DEQ & ~n44390;
  assign n44392 = ~n26609 & ~n44391;
  assign n44393 = ~i_FULL & ~n44392;
  assign n44394 = ~n44385 & ~n44393;
  assign n44395 = i_nEMPTY & ~n44394;
  assign n44396 = ~n26619 & ~n42037;
  assign n44397 = i_FULL & ~n44396;
  assign n44398 = ~n26627 & ~n42043;
  assign n44399 = ~i_FULL & ~n44398;
  assign n44400 = ~n44397 & ~n44399;
  assign n44401 = ~i_nEMPTY & ~n44400;
  assign n44402 = ~n44395 & ~n44401;
  assign n44403 = ~controllable_BtoS_ACK0 & ~n44402;
  assign n44404 = ~n44377 & ~n44403;
  assign n44405 = n4465 & ~n44404;
  assign n44406 = ~n11317 & ~n38262;
  assign n44407 = ~controllable_BtoR_REQ0 & ~n44406;
  assign n44408 = ~n16262 & ~n44407;
  assign n44409 = ~i_RtoB_ACK0 & ~n44408;
  assign n44410 = ~n42817 & ~n44409;
  assign n44411 = controllable_DEQ & ~n44410;
  assign n44412 = ~n26681 & ~n44411;
  assign n44413 = i_FULL & ~n44412;
  assign n44414 = ~n11317 & ~n38272;
  assign n44415 = ~controllable_BtoR_REQ0 & ~n44414;
  assign n44416 = ~n16300 & ~n44415;
  assign n44417 = ~i_RtoB_ACK0 & ~n44416;
  assign n44418 = ~n42817 & ~n44417;
  assign n44419 = controllable_DEQ & ~n44418;
  assign n44420 = ~n26695 & ~n44419;
  assign n44421 = ~i_FULL & ~n44420;
  assign n44422 = ~n44413 & ~n44421;
  assign n44423 = i_nEMPTY & ~n44422;
  assign n44424 = ~n26705 & ~n42071;
  assign n44425 = i_FULL & ~n44424;
  assign n44426 = ~n26713 & ~n42077;
  assign n44427 = ~i_FULL & ~n44426;
  assign n44428 = ~n44425 & ~n44427;
  assign n44429 = ~i_nEMPTY & ~n44428;
  assign n44430 = ~n44423 & ~n44429;
  assign n44431 = ~controllable_BtoS_ACK0 & ~n44430;
  assign n44432 = ~n26669 & ~n44431;
  assign n44433 = ~n4465 & ~n44432;
  assign n44434 = ~n44405 & ~n44433;
  assign n44435 = ~i_StoB_REQ10 & ~n44434;
  assign n44436 = ~n44351 & ~n44435;
  assign n44437 = controllable_BtoS_ACK10 & ~n44436;
  assign n44438 = ~n11238 & ~n38320;
  assign n44439 = ~controllable_BtoR_REQ0 & ~n44438;
  assign n44440 = ~n20002 & ~n44439;
  assign n44441 = ~i_RtoB_ACK0 & ~n44440;
  assign n44442 = ~n42855 & ~n44441;
  assign n44443 = controllable_DEQ & ~n44442;
  assign n44444 = ~n26737 & ~n44443;
  assign n44445 = i_FULL & ~n44444;
  assign n44446 = ~n11238 & ~n38330;
  assign n44447 = ~controllable_BtoR_REQ0 & ~n44446;
  assign n44448 = ~n20022 & ~n44447;
  assign n44449 = ~i_RtoB_ACK0 & ~n44448;
  assign n44450 = ~n42855 & ~n44449;
  assign n44451 = controllable_DEQ & ~n44450;
  assign n44452 = ~n26751 & ~n44451;
  assign n44453 = ~i_FULL & ~n44452;
  assign n44454 = ~n44445 & ~n44453;
  assign n44455 = i_nEMPTY & ~n44454;
  assign n44456 = ~n26761 & ~n42109;
  assign n44457 = i_FULL & ~n44456;
  assign n44458 = ~n26764 & ~n42115;
  assign n44459 = ~i_FULL & ~n44458;
  assign n44460 = ~n44457 & ~n44459;
  assign n44461 = ~i_nEMPTY & ~n44460;
  assign n44462 = ~n44455 & ~n44461;
  assign n44463 = controllable_BtoS_ACK0 & ~n44462;
  assign n44464 = ~n11317 & ~n38372;
  assign n44465 = ~controllable_BtoR_REQ0 & ~n44464;
  assign n44466 = ~n20068 & ~n44465;
  assign n44467 = ~i_RtoB_ACK0 & ~n44466;
  assign n44468 = ~n42887 & ~n44467;
  assign n44469 = controllable_DEQ & ~n44468;
  assign n44470 = ~n26780 & ~n44469;
  assign n44471 = i_FULL & ~n44470;
  assign n44472 = ~n11317 & ~n38382;
  assign n44473 = ~controllable_BtoR_REQ0 & ~n44472;
  assign n44474 = ~n20080 & ~n44473;
  assign n44475 = ~i_RtoB_ACK0 & ~n44474;
  assign n44476 = ~n42887 & ~n44475;
  assign n44477 = controllable_DEQ & ~n44476;
  assign n44478 = ~n26794 & ~n44477;
  assign n44479 = ~i_FULL & ~n44478;
  assign n44480 = ~n44471 & ~n44479;
  assign n44481 = i_nEMPTY & ~n44480;
  assign n44482 = ~n26802 & ~n42141;
  assign n44483 = i_FULL & ~n44482;
  assign n44484 = ~n26805 & ~n42147;
  assign n44485 = ~i_FULL & ~n44484;
  assign n44486 = ~n44483 & ~n44485;
  assign n44487 = ~i_nEMPTY & ~n44486;
  assign n44488 = ~n44481 & ~n44487;
  assign n44489 = ~controllable_BtoS_ACK0 & ~n44488;
  assign n44490 = ~n44463 & ~n44489;
  assign n44491 = n4465 & ~n44490;
  assign n44492 = ~n11317 & ~n38426;
  assign n44493 = ~controllable_BtoR_REQ0 & ~n44492;
  assign n44494 = ~n20156 & ~n44493;
  assign n44495 = ~i_RtoB_ACK0 & ~n44494;
  assign n44496 = ~n42921 & ~n44495;
  assign n44497 = controllable_DEQ & ~n44496;
  assign n44498 = ~n26848 & ~n44497;
  assign n44499 = i_FULL & ~n44498;
  assign n44500 = ~n11317 & ~n38436;
  assign n44501 = ~controllable_BtoR_REQ0 & ~n44500;
  assign n44502 = ~n20168 & ~n44501;
  assign n44503 = ~i_RtoB_ACK0 & ~n44502;
  assign n44504 = ~n42921 & ~n44503;
  assign n44505 = controllable_DEQ & ~n44504;
  assign n44506 = ~n26860 & ~n44505;
  assign n44507 = ~i_FULL & ~n44506;
  assign n44508 = ~n44499 & ~n44507;
  assign n44509 = i_nEMPTY & ~n44508;
  assign n44510 = ~n26868 & ~n42175;
  assign n44511 = i_FULL & ~n44510;
  assign n44512 = ~n26871 & ~n42181;
  assign n44513 = ~i_FULL & ~n44512;
  assign n44514 = ~n44511 & ~n44513;
  assign n44515 = ~i_nEMPTY & ~n44514;
  assign n44516 = ~n44509 & ~n44515;
  assign n44517 = ~controllable_BtoS_ACK0 & ~n44516;
  assign n44518 = ~n26838 & ~n44517;
  assign n44519 = ~n4465 & ~n44518;
  assign n44520 = ~n44491 & ~n44519;
  assign n44521 = i_StoB_REQ10 & ~n44520;
  assign n44522 = ~n44435 & ~n44521;
  assign n44523 = ~controllable_BtoS_ACK10 & ~n44522;
  assign n44524 = ~n44437 & ~n44523;
  assign n44525 = ~n4464 & ~n44524;
  assign n44526 = ~n44333 & ~n44525;
  assign n44527 = n4463 & ~n44526;
  assign n44528 = ~n27731 & ~n43936;
  assign n44529 = i_FULL & ~n44528;
  assign n44530 = ~n27731 & ~n43944;
  assign n44531 = ~i_FULL & ~n44530;
  assign n44532 = ~n44529 & ~n44531;
  assign n44533 = i_nEMPTY & ~n44532;
  assign n44534 = ~n43965 & ~n44533;
  assign n44535 = controllable_BtoS_ACK0 & ~n44534;
  assign n44536 = ~n27765 & ~n43972;
  assign n44537 = i_FULL & ~n44536;
  assign n44538 = ~n27765 & ~n43980;
  assign n44539 = ~i_FULL & ~n44538;
  assign n44540 = ~n44537 & ~n44539;
  assign n44541 = i_nEMPTY & ~n44540;
  assign n44542 = ~n44001 & ~n44541;
  assign n44543 = ~controllable_BtoS_ACK0 & ~n44542;
  assign n44544 = ~n44535 & ~n44543;
  assign n44545 = n4465 & ~n44544;
  assign n44546 = ~n44013 & ~n44545;
  assign n44547 = i_StoB_REQ10 & ~n44546;
  assign n44548 = ~n17280 & ~n43489;
  assign n44549 = i_RtoB_ACK0 & ~n44548;
  assign n44550 = ~n37256 & ~n40712;
  assign n44551 = ~controllable_BtoR_REQ0 & ~n44550;
  assign n44552 = ~n17974 & ~n44551;
  assign n44553 = ~i_RtoB_ACK0 & ~n44552;
  assign n44554 = ~n44549 & ~n44553;
  assign n44555 = controllable_DEQ & ~n44554;
  assign n44556 = ~n37470 & ~n40726;
  assign n44557 = ~controllable_BtoR_REQ0 & ~n44556;
  assign n44558 = ~n17993 & ~n44557;
  assign n44559 = ~i_RtoB_ACK0 & ~n44558;
  assign n44560 = ~n42459 & ~n44559;
  assign n44561 = ~controllable_DEQ & ~n44560;
  assign n44562 = ~n44555 & ~n44561;
  assign n44563 = i_FULL & ~n44562;
  assign n44564 = ~n37480 & ~n40712;
  assign n44565 = ~controllable_BtoR_REQ0 & ~n44564;
  assign n44566 = ~n18012 & ~n44565;
  assign n44567 = ~i_RtoB_ACK0 & ~n44566;
  assign n44568 = ~n44549 & ~n44567;
  assign n44569 = controllable_DEQ & ~n44568;
  assign n44570 = ~n37488 & ~n40740;
  assign n44571 = ~controllable_BtoR_REQ0 & ~n44570;
  assign n44572 = ~n18028 & ~n44571;
  assign n44573 = ~i_RtoB_ACK0 & ~n44572;
  assign n44574 = ~n42459 & ~n44573;
  assign n44575 = ~controllable_DEQ & ~n44574;
  assign n44576 = ~n44569 & ~n44575;
  assign n44577 = ~i_FULL & ~n44576;
  assign n44578 = ~n44563 & ~n44577;
  assign n44579 = i_nEMPTY & ~n44578;
  assign n44580 = ~n37529 & ~n40764;
  assign n44581 = ~controllable_BtoR_REQ0 & ~n44580;
  assign n44582 = ~n18065 & ~n44581;
  assign n44583 = ~i_RtoB_ACK0 & ~n44582;
  assign n44584 = ~n42483 & ~n44583;
  assign n44585 = ~controllable_DEQ & ~n44584;
  assign n44586 = ~n43001 & ~n44585;
  assign n44587 = i_FULL & ~n44586;
  assign n44588 = ~n37552 & ~n40787;
  assign n44589 = ~controllable_BtoR_REQ0 & ~n44588;
  assign n44590 = ~n17974 & ~n44589;
  assign n44591 = ~i_RtoB_ACK0 & ~n44590;
  assign n44592 = ~n42495 & ~n44591;
  assign n44593 = ~controllable_DEQ & ~n44592;
  assign n44594 = ~n43009 & ~n44593;
  assign n44595 = ~i_FULL & ~n44594;
  assign n44596 = ~n44587 & ~n44595;
  assign n44597 = ~i_nEMPTY & ~n44596;
  assign n44598 = ~n44579 & ~n44597;
  assign n44599 = controllable_BtoS_ACK0 & ~n44598;
  assign n44600 = ~n17690 & ~n43539;
  assign n44601 = i_RtoB_ACK0 & ~n44600;
  assign n44602 = ~n37698 & ~n40804;
  assign n44603 = ~controllable_BtoR_REQ0 & ~n44602;
  assign n44604 = ~n18116 & ~n44603;
  assign n44605 = ~i_RtoB_ACK0 & ~n44604;
  assign n44606 = ~n44601 & ~n44605;
  assign n44607 = controllable_DEQ & ~n44606;
  assign n44608 = ~n37733 & ~n40818;
  assign n44609 = ~controllable_BtoR_REQ0 & ~n44608;
  assign n44610 = ~n18135 & ~n44609;
  assign n44611 = ~i_RtoB_ACK0 & ~n44610;
  assign n44612 = ~n42513 & ~n44611;
  assign n44613 = ~controllable_DEQ & ~n44612;
  assign n44614 = ~n44607 & ~n44613;
  assign n44615 = i_FULL & ~n44614;
  assign n44616 = ~n37743 & ~n40804;
  assign n44617 = ~controllable_BtoR_REQ0 & ~n44616;
  assign n44618 = ~n18154 & ~n44617;
  assign n44619 = ~i_RtoB_ACK0 & ~n44618;
  assign n44620 = ~n44601 & ~n44619;
  assign n44621 = controllable_DEQ & ~n44620;
  assign n44622 = ~n37751 & ~n40832;
  assign n44623 = ~controllable_BtoR_REQ0 & ~n44622;
  assign n44624 = ~n18170 & ~n44623;
  assign n44625 = ~i_RtoB_ACK0 & ~n44624;
  assign n44626 = ~n42513 & ~n44625;
  assign n44627 = ~controllable_DEQ & ~n44626;
  assign n44628 = ~n44621 & ~n44627;
  assign n44629 = ~i_FULL & ~n44628;
  assign n44630 = ~n44615 & ~n44629;
  assign n44631 = i_nEMPTY & ~n44630;
  assign n44632 = ~n37792 & ~n40856;
  assign n44633 = ~controllable_BtoR_REQ0 & ~n44632;
  assign n44634 = ~n18207 & ~n44633;
  assign n44635 = ~i_RtoB_ACK0 & ~n44634;
  assign n44636 = ~n42537 & ~n44635;
  assign n44637 = ~controllable_DEQ & ~n44636;
  assign n44638 = ~n43039 & ~n44637;
  assign n44639 = i_FULL & ~n44638;
  assign n44640 = ~n37815 & ~n40879;
  assign n44641 = ~controllable_BtoR_REQ0 & ~n44640;
  assign n44642 = ~n18116 & ~n44641;
  assign n44643 = ~i_RtoB_ACK0 & ~n44642;
  assign n44644 = ~n42549 & ~n44643;
  assign n44645 = ~controllable_DEQ & ~n44644;
  assign n44646 = ~n43047 & ~n44645;
  assign n44647 = ~i_FULL & ~n44646;
  assign n44648 = ~n44639 & ~n44647;
  assign n44649 = ~i_nEMPTY & ~n44648;
  assign n44650 = ~n44631 & ~n44649;
  assign n44651 = ~controllable_BtoS_ACK0 & ~n44650;
  assign n44652 = ~n44599 & ~n44651;
  assign n44653 = n4465 & ~n44652;
  assign n44654 = ~n17690 & ~n43591;
  assign n44655 = i_RtoB_ACK0 & ~n44654;
  assign n44656 = ~n44145 & ~n44655;
  assign n44657 = controllable_DEQ & ~n44656;
  assign n44658 = ~n26219 & ~n44657;
  assign n44659 = i_FULL & ~n44658;
  assign n44660 = ~n44153 & ~n44655;
  assign n44661 = controllable_DEQ & ~n44660;
  assign n44662 = ~n26233 & ~n44661;
  assign n44663 = ~i_FULL & ~n44662;
  assign n44664 = ~n44659 & ~n44663;
  assign n44665 = i_nEMPTY & ~n44664;
  assign n44666 = ~n44165 & ~n44665;
  assign n44667 = ~controllable_BtoS_ACK0 & ~n44666;
  assign n44668 = ~n27023 & ~n44667;
  assign n44669 = ~n4465 & ~n44668;
  assign n44670 = ~n44653 & ~n44669;
  assign n44671 = ~i_StoB_REQ10 & ~n44670;
  assign n44672 = ~n44547 & ~n44671;
  assign n44673 = controllable_BtoS_ACK10 & ~n44672;
  assign n44674 = ~n17050 & ~n43613;
  assign n44675 = i_RtoB_ACK0 & ~n44674;
  assign n44676 = ~n11238 & ~n37908;
  assign n44677 = ~controllable_BtoR_REQ0 & ~n44676;
  assign n44678 = ~n40928 & ~n44677;
  assign n44679 = ~i_RtoB_ACK0 & ~n44678;
  assign n44680 = ~n44675 & ~n44679;
  assign n44681 = controllable_DEQ & ~n44680;
  assign n44682 = ~n44185 & ~n44681;
  assign n44683 = i_FULL & ~n44682;
  assign n44684 = ~n11238 & ~n37927;
  assign n44685 = ~controllable_BtoR_REQ0 & ~n44684;
  assign n44686 = ~n40944 & ~n44685;
  assign n44687 = ~i_RtoB_ACK0 & ~n44686;
  assign n44688 = ~n44675 & ~n44687;
  assign n44689 = controllable_DEQ & ~n44688;
  assign n44690 = ~n44199 & ~n44689;
  assign n44691 = ~i_FULL & ~n44690;
  assign n44692 = ~n44683 & ~n44691;
  assign n44693 = i_nEMPTY & ~n44692;
  assign n44694 = ~n43093 & ~n44215;
  assign n44695 = i_FULL & ~n44694;
  assign n44696 = ~n43097 & ~n44229;
  assign n44697 = ~i_FULL & ~n44696;
  assign n44698 = ~n44695 & ~n44697;
  assign n44699 = ~i_nEMPTY & ~n44698;
  assign n44700 = ~n44693 & ~n44699;
  assign n44701 = controllable_BtoS_ACK0 & ~n44700;
  assign n44702 = ~n18522 & ~n43655;
  assign n44703 = i_RtoB_ACK0 & ~n44702;
  assign n44704 = ~n11317 & ~n37992;
  assign n44705 = ~controllable_BtoR_REQ0 & ~n44704;
  assign n44706 = ~n40999 & ~n44705;
  assign n44707 = ~i_RtoB_ACK0 & ~n44706;
  assign n44708 = ~n44703 & ~n44707;
  assign n44709 = controllable_DEQ & ~n44708;
  assign n44710 = ~n44247 & ~n44709;
  assign n44711 = i_FULL & ~n44710;
  assign n44712 = ~n11317 & ~n38011;
  assign n44713 = ~controllable_BtoR_REQ0 & ~n44712;
  assign n44714 = ~n41015 & ~n44713;
  assign n44715 = ~i_RtoB_ACK0 & ~n44714;
  assign n44716 = ~n44703 & ~n44715;
  assign n44717 = controllable_DEQ & ~n44716;
  assign n44718 = ~n44261 & ~n44717;
  assign n44719 = ~i_FULL & ~n44718;
  assign n44720 = ~n44711 & ~n44719;
  assign n44721 = i_nEMPTY & ~n44720;
  assign n44722 = ~n43117 & ~n44277;
  assign n44723 = i_FULL & ~n44722;
  assign n44724 = ~n43121 & ~n44291;
  assign n44725 = ~i_FULL & ~n44724;
  assign n44726 = ~n44723 & ~n44725;
  assign n44727 = ~i_nEMPTY & ~n44726;
  assign n44728 = ~n44721 & ~n44727;
  assign n44729 = ~controllable_BtoS_ACK0 & ~n44728;
  assign n44730 = ~n44701 & ~n44729;
  assign n44731 = n4465 & ~n44730;
  assign n44732 = ~n18522 & ~n43699;
  assign n44733 = i_RtoB_ACK0 & ~n44732;
  assign n44734 = ~n44303 & ~n44733;
  assign n44735 = controllable_DEQ & ~n44734;
  assign n44736 = ~n26394 & ~n44735;
  assign n44737 = i_FULL & ~n44736;
  assign n44738 = ~n44311 & ~n44733;
  assign n44739 = controllable_DEQ & ~n44738;
  assign n44740 = ~n26406 & ~n44739;
  assign n44741 = ~i_FULL & ~n44740;
  assign n44742 = ~n44737 & ~n44741;
  assign n44743 = i_nEMPTY & ~n44742;
  assign n44744 = ~n44323 & ~n44743;
  assign n44745 = ~controllable_BtoS_ACK0 & ~n44744;
  assign n44746 = ~n26384 & ~n44745;
  assign n44747 = ~n4465 & ~n44746;
  assign n44748 = ~n44731 & ~n44747;
  assign n44749 = i_StoB_REQ10 & ~n44748;
  assign n44750 = ~n44671 & ~n44749;
  assign n44751 = ~controllable_BtoS_ACK10 & ~n44750;
  assign n44752 = ~n44673 & ~n44751;
  assign n44753 = n4464 & ~n44752;
  assign n44754 = ~n17280 & ~n43723;
  assign n44755 = i_RtoB_ACK0 & ~n44754;
  assign n44756 = ~n19765 & ~n38156;
  assign n44757 = ~controllable_BtoR_REQ0 & ~n44756;
  assign n44758 = ~n15889 & ~n44757;
  assign n44759 = ~i_RtoB_ACK0 & ~n44758;
  assign n44760 = ~n44755 & ~n44759;
  assign n44761 = controllable_DEQ & ~n44760;
  assign n44762 = ~n27045 & ~n44761;
  assign n44763 = i_FULL & ~n44762;
  assign n44764 = ~n19765 & ~n38166;
  assign n44765 = ~controllable_BtoR_REQ0 & ~n44764;
  assign n44766 = ~n15927 & ~n44765;
  assign n44767 = ~i_RtoB_ACK0 & ~n44766;
  assign n44768 = ~n44755 & ~n44767;
  assign n44769 = controllable_DEQ & ~n44768;
  assign n44770 = ~n27059 & ~n44769;
  assign n44771 = ~i_FULL & ~n44770;
  assign n44772 = ~n44763 & ~n44771;
  assign n44773 = i_nEMPTY & ~n44772;
  assign n44774 = ~n27069 & ~n42005;
  assign n44775 = i_FULL & ~n44774;
  assign n44776 = ~n27077 & ~n42011;
  assign n44777 = ~i_FULL & ~n44776;
  assign n44778 = ~n44775 & ~n44777;
  assign n44779 = ~i_nEMPTY & ~n44778;
  assign n44780 = ~n44773 & ~n44779;
  assign n44781 = controllable_BtoS_ACK0 & ~n44780;
  assign n44782 = ~n17690 & ~n43745;
  assign n44783 = i_RtoB_ACK0 & ~n44782;
  assign n44784 = ~n19839 & ~n38208;
  assign n44785 = ~controllable_BtoR_REQ0 & ~n44784;
  assign n44786 = ~n16031 & ~n44785;
  assign n44787 = ~i_RtoB_ACK0 & ~n44786;
  assign n44788 = ~n44783 & ~n44787;
  assign n44789 = controllable_DEQ & ~n44788;
  assign n44790 = ~n27095 & ~n44789;
  assign n44791 = i_FULL & ~n44790;
  assign n44792 = ~n19839 & ~n38218;
  assign n44793 = ~controllable_BtoR_REQ0 & ~n44792;
  assign n44794 = ~n16069 & ~n44793;
  assign n44795 = ~i_RtoB_ACK0 & ~n44794;
  assign n44796 = ~n44783 & ~n44795;
  assign n44797 = controllable_DEQ & ~n44796;
  assign n44798 = ~n27109 & ~n44797;
  assign n44799 = ~i_FULL & ~n44798;
  assign n44800 = ~n44791 & ~n44799;
  assign n44801 = i_nEMPTY & ~n44800;
  assign n44802 = ~n27119 & ~n42037;
  assign n44803 = i_FULL & ~n44802;
  assign n44804 = ~n27127 & ~n42043;
  assign n44805 = ~i_FULL & ~n44804;
  assign n44806 = ~n44803 & ~n44805;
  assign n44807 = ~i_nEMPTY & ~n44806;
  assign n44808 = ~n44801 & ~n44807;
  assign n44809 = ~controllable_BtoS_ACK0 & ~n44808;
  assign n44810 = ~n44781 & ~n44809;
  assign n44811 = n4465 & ~n44810;
  assign n44812 = ~n17690 & ~n43769;
  assign n44813 = i_RtoB_ACK0 & ~n44812;
  assign n44814 = ~n44409 & ~n44813;
  assign n44815 = controllable_DEQ & ~n44814;
  assign n44816 = ~n26681 & ~n44815;
  assign n44817 = i_FULL & ~n44816;
  assign n44818 = ~n44417 & ~n44813;
  assign n44819 = controllable_DEQ & ~n44818;
  assign n44820 = ~n26695 & ~n44819;
  assign n44821 = ~i_FULL & ~n44820;
  assign n44822 = ~n44817 & ~n44821;
  assign n44823 = i_nEMPTY & ~n44822;
  assign n44824 = ~n44429 & ~n44823;
  assign n44825 = ~controllable_BtoS_ACK0 & ~n44824;
  assign n44826 = ~n26669 & ~n44825;
  assign n44827 = ~n4465 & ~n44826;
  assign n44828 = ~n44811 & ~n44827;
  assign n44829 = ~i_StoB_REQ10 & ~n44828;
  assign n44830 = ~n44351 & ~n44829;
  assign n44831 = controllable_BtoS_ACK10 & ~n44830;
  assign n44832 = ~n17050 & ~n43791;
  assign n44833 = i_RtoB_ACK0 & ~n44832;
  assign n44834 = ~n44441 & ~n44833;
  assign n44835 = controllable_DEQ & ~n44834;
  assign n44836 = ~n26737 & ~n44835;
  assign n44837 = i_FULL & ~n44836;
  assign n44838 = ~n44449 & ~n44833;
  assign n44839 = controllable_DEQ & ~n44838;
  assign n44840 = ~n26751 & ~n44839;
  assign n44841 = ~i_FULL & ~n44840;
  assign n44842 = ~n44837 & ~n44841;
  assign n44843 = i_nEMPTY & ~n44842;
  assign n44844 = ~n44461 & ~n44843;
  assign n44845 = controllable_BtoS_ACK0 & ~n44844;
  assign n44846 = ~n18522 & ~n43807;
  assign n44847 = i_RtoB_ACK0 & ~n44846;
  assign n44848 = ~n44467 & ~n44847;
  assign n44849 = controllable_DEQ & ~n44848;
  assign n44850 = ~n26780 & ~n44849;
  assign n44851 = i_FULL & ~n44850;
  assign n44852 = ~n44475 & ~n44847;
  assign n44853 = controllable_DEQ & ~n44852;
  assign n44854 = ~n26794 & ~n44853;
  assign n44855 = ~i_FULL & ~n44854;
  assign n44856 = ~n44851 & ~n44855;
  assign n44857 = i_nEMPTY & ~n44856;
  assign n44858 = ~n44487 & ~n44857;
  assign n44859 = ~controllable_BtoS_ACK0 & ~n44858;
  assign n44860 = ~n44845 & ~n44859;
  assign n44861 = n4465 & ~n44860;
  assign n44862 = ~n18522 & ~n43825;
  assign n44863 = i_RtoB_ACK0 & ~n44862;
  assign n44864 = ~n44495 & ~n44863;
  assign n44865 = controllable_DEQ & ~n44864;
  assign n44866 = ~n26848 & ~n44865;
  assign n44867 = i_FULL & ~n44866;
  assign n44868 = ~n44503 & ~n44863;
  assign n44869 = controllable_DEQ & ~n44868;
  assign n44870 = ~n26860 & ~n44869;
  assign n44871 = ~i_FULL & ~n44870;
  assign n44872 = ~n44867 & ~n44871;
  assign n44873 = i_nEMPTY & ~n44872;
  assign n44874 = ~n44515 & ~n44873;
  assign n44875 = ~controllable_BtoS_ACK0 & ~n44874;
  assign n44876 = ~n26838 & ~n44875;
  assign n44877 = ~n4465 & ~n44876;
  assign n44878 = ~n44861 & ~n44877;
  assign n44879 = i_StoB_REQ10 & ~n44878;
  assign n44880 = ~n44829 & ~n44879;
  assign n44881 = ~controllable_BtoS_ACK10 & ~n44880;
  assign n44882 = ~n44831 & ~n44881;
  assign n44883 = ~n4464 & ~n44882;
  assign n44884 = ~n44753 & ~n44883;
  assign n44885 = ~n4463 & ~n44884;
  assign n44886 = ~n44527 & ~n44885;
  assign n44887 = n4462 & ~n44886;
  assign n44888 = ~n11238 & ~n12363;
  assign n44889 = ~controllable_BtoR_REQ0 & ~n44888;
  assign n44890 = ~n20366 & ~n44889;
  assign n44891 = ~i_RtoB_ACK0 & ~n44890;
  assign n44892 = ~n25187 & ~n44891;
  assign n44893 = controllable_DEQ & ~n44892;
  assign n44894 = ~n27263 & ~n44893;
  assign n44895 = i_FULL & ~n44894;
  assign n44896 = ~n27279 & ~n44895;
  assign n44897 = i_nEMPTY & ~n44896;
  assign n44898 = ~n27294 & ~n44897;
  assign n44899 = controllable_BtoS_ACK0 & ~n44898;
  assign n44900 = ~n11317 & ~n12464;
  assign n44901 = ~controllable_BtoR_REQ0 & ~n44900;
  assign n44902 = ~n20432 & ~n44901;
  assign n44903 = ~i_RtoB_ACK0 & ~n44902;
  assign n44904 = ~n25228 & ~n44903;
  assign n44905 = controllable_DEQ & ~n44904;
  assign n44906 = ~n27306 & ~n44905;
  assign n44907 = i_FULL & ~n44906;
  assign n44908 = ~n27322 & ~n44907;
  assign n44909 = i_nEMPTY & ~n44908;
  assign n44910 = ~n27335 & ~n44909;
  assign n44911 = ~controllable_BtoS_ACK0 & ~n44910;
  assign n44912 = ~n44899 & ~n44911;
  assign n44913 = n4465 & ~n44912;
  assign n44914 = ~n26384 & ~n44911;
  assign n44915 = ~n4465 & ~n44914;
  assign n44916 = ~n44913 & ~n44915;
  assign n44917 = i_StoB_REQ10 & ~n44916;
  assign n44918 = ~n11238 & ~n37256;
  assign n44919 = ~controllable_BtoR_REQ0 & ~n44918;
  assign n44920 = ~n17974 & ~n44919;
  assign n44921 = ~i_RtoB_ACK0 & ~n44920;
  assign n44922 = ~n42453 & ~n44921;
  assign n44923 = controllable_DEQ & ~n44922;
  assign n44924 = ~n27353 & ~n44923;
  assign n44925 = i_FULL & ~n44924;
  assign n44926 = ~n11238 & ~n37480;
  assign n44927 = ~controllable_BtoR_REQ0 & ~n44926;
  assign n44928 = ~n18012 & ~n44927;
  assign n44929 = ~i_RtoB_ACK0 & ~n44928;
  assign n44930 = ~n42453 & ~n44929;
  assign n44931 = controllable_DEQ & ~n44930;
  assign n44932 = ~n27367 & ~n44931;
  assign n44933 = ~i_FULL & ~n44932;
  assign n44934 = ~n44925 & ~n44933;
  assign n44935 = i_nEMPTY & ~n44934;
  assign n44936 = ~n27375 & ~n42245;
  assign n44937 = i_FULL & ~n44936;
  assign n44938 = ~n27383 & ~n42251;
  assign n44939 = ~i_FULL & ~n44938;
  assign n44940 = ~n44937 & ~n44939;
  assign n44941 = ~i_nEMPTY & ~n44940;
  assign n44942 = ~n44935 & ~n44941;
  assign n44943 = controllable_BtoS_ACK0 & ~n44942;
  assign n44944 = ~n11317 & ~n37698;
  assign n44945 = ~controllable_BtoR_REQ0 & ~n44944;
  assign n44946 = ~n18116 & ~n44945;
  assign n44947 = ~i_RtoB_ACK0 & ~n44946;
  assign n44948 = ~n42507 & ~n44947;
  assign n44949 = controllable_DEQ & ~n44948;
  assign n44950 = ~n27399 & ~n44949;
  assign n44951 = i_FULL & ~n44950;
  assign n44952 = ~n11317 & ~n37743;
  assign n44953 = ~controllable_BtoR_REQ0 & ~n44952;
  assign n44954 = ~n18154 & ~n44953;
  assign n44955 = ~i_RtoB_ACK0 & ~n44954;
  assign n44956 = ~n42507 & ~n44955;
  assign n44957 = controllable_DEQ & ~n44956;
  assign n44958 = ~n27413 & ~n44957;
  assign n44959 = ~i_FULL & ~n44958;
  assign n44960 = ~n44951 & ~n44959;
  assign n44961 = i_nEMPTY & ~n44960;
  assign n44962 = ~n27421 & ~n42277;
  assign n44963 = i_FULL & ~n44962;
  assign n44964 = ~n27429 & ~n42283;
  assign n44965 = ~i_FULL & ~n44964;
  assign n44966 = ~n44963 & ~n44965;
  assign n44967 = ~i_nEMPTY & ~n44966;
  assign n44968 = ~n44961 & ~n44967;
  assign n44969 = ~controllable_BtoS_ACK0 & ~n44968;
  assign n44970 = ~n44943 & ~n44969;
  assign n44971 = n4465 & ~n44970;
  assign n44972 = ~n27467 & ~n44167;
  assign n44973 = ~n4465 & ~n44972;
  assign n44974 = ~n44971 & ~n44973;
  assign n44975 = ~i_StoB_REQ10 & ~n44974;
  assign n44976 = ~n44917 & ~n44975;
  assign n44977 = ~controllable_BtoS_ACK10 & ~n44976;
  assign n44978 = ~n27251 & ~n44977;
  assign n44979 = n4464 & ~n44978;
  assign n44980 = ~n11238 & ~n12865;
  assign n44981 = ~controllable_BtoR_REQ0 & ~n44980;
  assign n44982 = ~n20680 & ~n44981;
  assign n44983 = ~i_RtoB_ACK0 & ~n44982;
  assign n44984 = ~n25401 & ~n44983;
  assign n44985 = controllable_DEQ & ~n44984;
  assign n44986 = ~n27549 & ~n44985;
  assign n44987 = i_FULL & ~n44986;
  assign n44988 = ~n27565 & ~n44987;
  assign n44989 = i_nEMPTY & ~n44988;
  assign n44990 = ~n27578 & ~n44989;
  assign n44991 = controllable_BtoS_ACK0 & ~n44990;
  assign n44992 = ~n11317 & ~n12950;
  assign n44993 = ~controllable_BtoR_REQ0 & ~n44992;
  assign n44994 = ~n20730 & ~n44993;
  assign n44995 = ~i_RtoB_ACK0 & ~n44994;
  assign n44996 = ~n25442 & ~n44995;
  assign n44997 = controllable_DEQ & ~n44996;
  assign n44998 = ~n27590 & ~n44997;
  assign n44999 = i_FULL & ~n44998;
  assign n45000 = ~n27606 & ~n44999;
  assign n45001 = i_nEMPTY & ~n45000;
  assign n45002 = ~n27619 & ~n45001;
  assign n45003 = ~controllable_BtoS_ACK0 & ~n45002;
  assign n45004 = ~n44991 & ~n45003;
  assign n45005 = n4465 & ~n45004;
  assign n45006 = ~n26838 & ~n45003;
  assign n45007 = ~n4465 & ~n45006;
  assign n45008 = ~n45005 & ~n45007;
  assign n45009 = i_StoB_REQ10 & ~n45008;
  assign n45010 = ~n11238 & ~n38156;
  assign n45011 = ~controllable_BtoR_REQ0 & ~n45010;
  assign n45012 = ~n15889 & ~n45011;
  assign n45013 = ~i_RtoB_ACK0 & ~n45012;
  assign n45014 = ~n42751 & ~n45013;
  assign n45015 = controllable_DEQ & ~n45014;
  assign n45016 = ~n27637 & ~n45015;
  assign n45017 = i_FULL & ~n45016;
  assign n45018 = ~n11238 & ~n38166;
  assign n45019 = ~controllable_BtoR_REQ0 & ~n45018;
  assign n45020 = ~n15927 & ~n45019;
  assign n45021 = ~i_RtoB_ACK0 & ~n45020;
  assign n45022 = ~n42751 & ~n45021;
  assign n45023 = controllable_DEQ & ~n45022;
  assign n45024 = ~n27649 & ~n45023;
  assign n45025 = ~i_FULL & ~n45024;
  assign n45026 = ~n45017 & ~n45025;
  assign n45027 = i_nEMPTY & ~n45026;
  assign n45028 = ~n27657 & ~n42345;
  assign n45029 = i_FULL & ~n45028;
  assign n45030 = ~n27665 & ~n42351;
  assign n45031 = ~i_FULL & ~n45030;
  assign n45032 = ~n45029 & ~n45031;
  assign n45033 = ~i_nEMPTY & ~n45032;
  assign n45034 = ~n45027 & ~n45033;
  assign n45035 = controllable_BtoS_ACK0 & ~n45034;
  assign n45036 = ~n11317 & ~n38208;
  assign n45037 = ~controllable_BtoR_REQ0 & ~n45036;
  assign n45038 = ~n16031 & ~n45037;
  assign n45039 = ~i_RtoB_ACK0 & ~n45038;
  assign n45040 = ~n42783 & ~n45039;
  assign n45041 = controllable_DEQ & ~n45040;
  assign n45042 = ~n27681 & ~n45041;
  assign n45043 = i_FULL & ~n45042;
  assign n45044 = ~n11317 & ~n38218;
  assign n45045 = ~controllable_BtoR_REQ0 & ~n45044;
  assign n45046 = ~n16069 & ~n45045;
  assign n45047 = ~i_RtoB_ACK0 & ~n45046;
  assign n45048 = ~n42783 & ~n45047;
  assign n45049 = controllable_DEQ & ~n45048;
  assign n45050 = ~n27693 & ~n45049;
  assign n45051 = ~i_FULL & ~n45050;
  assign n45052 = ~n45043 & ~n45051;
  assign n45053 = i_nEMPTY & ~n45052;
  assign n45054 = ~n27701 & ~n42377;
  assign n45055 = i_FULL & ~n45054;
  assign n45056 = ~n27709 & ~n42383;
  assign n45057 = ~i_FULL & ~n45056;
  assign n45058 = ~n45055 & ~n45057;
  assign n45059 = ~i_nEMPTY & ~n45058;
  assign n45060 = ~n45053 & ~n45059;
  assign n45061 = ~controllable_BtoS_ACK0 & ~n45060;
  assign n45062 = ~n45035 & ~n45061;
  assign n45063 = n4465 & ~n45062;
  assign n45064 = ~n44433 & ~n45063;
  assign n45065 = ~i_StoB_REQ10 & ~n45064;
  assign n45066 = ~n45009 & ~n45065;
  assign n45067 = ~controllable_BtoS_ACK10 & ~n45066;
  assign n45068 = ~n27539 & ~n45067;
  assign n45069 = ~n4464 & ~n45068;
  assign n45070 = ~n44979 & ~n45069;
  assign n45071 = n4463 & ~n45070;
  assign n45072 = ~n44549 & ~n44921;
  assign n45073 = controllable_DEQ & ~n45072;
  assign n45074 = ~n27353 & ~n45073;
  assign n45075 = i_FULL & ~n45074;
  assign n45076 = ~n44549 & ~n44929;
  assign n45077 = controllable_DEQ & ~n45076;
  assign n45078 = ~n27367 & ~n45077;
  assign n45079 = ~i_FULL & ~n45078;
  assign n45080 = ~n45075 & ~n45079;
  assign n45081 = i_nEMPTY & ~n45080;
  assign n45082 = ~n44941 & ~n45081;
  assign n45083 = controllable_BtoS_ACK0 & ~n45082;
  assign n45084 = ~n44601 & ~n44947;
  assign n45085 = controllable_DEQ & ~n45084;
  assign n45086 = ~n27399 & ~n45085;
  assign n45087 = i_FULL & ~n45086;
  assign n45088 = ~n44601 & ~n44955;
  assign n45089 = controllable_DEQ & ~n45088;
  assign n45090 = ~n27413 & ~n45089;
  assign n45091 = ~i_FULL & ~n45090;
  assign n45092 = ~n45087 & ~n45091;
  assign n45093 = i_nEMPTY & ~n45092;
  assign n45094 = ~n44967 & ~n45093;
  assign n45095 = ~controllable_BtoS_ACK0 & ~n45094;
  assign n45096 = ~n45083 & ~n45095;
  assign n45097 = n4465 & ~n45096;
  assign n45098 = ~n27467 & ~n44667;
  assign n45099 = ~n4465 & ~n45098;
  assign n45100 = ~n45097 & ~n45099;
  assign n45101 = ~i_StoB_REQ10 & ~n45100;
  assign n45102 = ~n44917 & ~n45101;
  assign n45103 = ~controllable_BtoS_ACK10 & ~n45102;
  assign n45104 = ~n27799 & ~n45103;
  assign n45105 = n4464 & ~n45104;
  assign n45106 = ~n44755 & ~n45013;
  assign n45107 = controllable_DEQ & ~n45106;
  assign n45108 = ~n27637 & ~n45107;
  assign n45109 = i_FULL & ~n45108;
  assign n45110 = ~n44755 & ~n45021;
  assign n45111 = controllable_DEQ & ~n45110;
  assign n45112 = ~n27649 & ~n45111;
  assign n45113 = ~i_FULL & ~n45112;
  assign n45114 = ~n45109 & ~n45113;
  assign n45115 = i_nEMPTY & ~n45114;
  assign n45116 = ~n45033 & ~n45115;
  assign n45117 = controllable_BtoS_ACK0 & ~n45116;
  assign n45118 = ~n44783 & ~n45039;
  assign n45119 = controllable_DEQ & ~n45118;
  assign n45120 = ~n27681 & ~n45119;
  assign n45121 = i_FULL & ~n45120;
  assign n45122 = ~n44783 & ~n45047;
  assign n45123 = controllable_DEQ & ~n45122;
  assign n45124 = ~n27693 & ~n45123;
  assign n45125 = ~i_FULL & ~n45124;
  assign n45126 = ~n45121 & ~n45125;
  assign n45127 = i_nEMPTY & ~n45126;
  assign n45128 = ~n45059 & ~n45127;
  assign n45129 = ~controllable_BtoS_ACK0 & ~n45128;
  assign n45130 = ~n45117 & ~n45129;
  assign n45131 = n4465 & ~n45130;
  assign n45132 = ~n44827 & ~n45131;
  assign n45133 = ~i_StoB_REQ10 & ~n45132;
  assign n45134 = ~n45009 & ~n45133;
  assign n45135 = ~controllable_BtoS_ACK10 & ~n45134;
  assign n45136 = ~n27539 & ~n45135;
  assign n45137 = ~n4464 & ~n45136;
  assign n45138 = ~n45105 & ~n45137;
  assign n45139 = ~n4463 & ~n45138;
  assign n45140 = ~n45071 & ~n45139;
  assign n45141 = ~n4462 & ~n45140;
  assign n45142 = ~n44887 & ~n45141;
  assign n45143 = ~n4461 & ~n45142;
  assign n45144 = ~n43931 & ~n45143;
  assign n45145 = n4459 & ~n45144;
  assign n45146 = ~n43475 & ~n45145;
  assign n45147 = ~n4455 & ~n45146;
  assign n45148 = ~n41471 & ~n45147;
  assign n45149 = n4445 & ~n45148;
  assign n45150 = ~i_RtoB_ACK1 & ~n37037;
  assign n45151 = ~i_RtoB_ACK1 & ~n45150;
  assign n45152 = controllable_BtoR_REQ1 & ~n45151;
  assign n45153 = ~controllable_BtoR_REQ1 & ~n12161;
  assign n45154 = ~n45152 & ~n45153;
  assign n45155 = ~controllable_BtoR_REQ0 & ~n45154;
  assign n45156 = ~controllable_BtoR_REQ0 & ~n45155;
  assign n45157 = i_RtoB_ACK0 & ~n45156;
  assign n45158 = ~controllable_BtoR_REQ1 & ~n14083;
  assign n45159 = ~n36888 & ~n45158;
  assign n45160 = ~controllable_BtoR_REQ0 & ~n45159;
  assign n45161 = ~controllable_BtoR_REQ0 & ~n45160;
  assign n45162 = ~i_RtoB_ACK0 & ~n45161;
  assign n45163 = ~n45157 & ~n45162;
  assign n45164 = ~controllable_DEQ & ~n45163;
  assign n45165 = ~n5251 & ~n45164;
  assign n45166 = i_FULL & ~n45165;
  assign n45167 = controllable_BtoR_REQ1 & ~n40617;
  assign n45168 = ~n14082 & ~n36899;
  assign n45169 = ~controllable_BtoR_REQ1 & ~n45168;
  assign n45170 = ~n45167 & ~n45169;
  assign n45171 = ~controllable_BtoR_REQ0 & ~n45170;
  assign n45172 = ~controllable_BtoR_REQ0 & ~n45171;
  assign n45173 = ~i_RtoB_ACK0 & ~n45172;
  assign n45174 = ~n45157 & ~n45173;
  assign n45175 = ~controllable_DEQ & ~n45174;
  assign n45176 = ~n5251 & ~n45175;
  assign n45177 = ~i_FULL & ~n45176;
  assign n45178 = ~n45166 & ~n45177;
  assign n45179 = i_nEMPTY & ~n45178;
  assign n45180 = controllable_ENQ & ~n37037;
  assign n45181 = controllable_ENQ & ~n45180;
  assign n45182 = ~i_RtoB_ACK1 & ~n45181;
  assign n45183 = ~i_RtoB_ACK1 & ~n45182;
  assign n45184 = controllable_BtoR_REQ1 & ~n45183;
  assign n45185 = ~controllable_BtoR_REQ1 & ~n12163;
  assign n45186 = ~n45184 & ~n45185;
  assign n45187 = ~controllable_BtoR_REQ0 & ~n45186;
  assign n45188 = ~controllable_BtoR_REQ0 & ~n45187;
  assign n45189 = i_RtoB_ACK0 & ~n45188;
  assign n45190 = ~controllable_BtoR_REQ1 & ~n14093;
  assign n45191 = ~n36923 & ~n45190;
  assign n45192 = ~controllable_BtoR_REQ0 & ~n45191;
  assign n45193 = ~controllable_BtoR_REQ0 & ~n45192;
  assign n45194 = ~i_RtoB_ACK0 & ~n45193;
  assign n45195 = ~n45189 & ~n45194;
  assign n45196 = ~controllable_DEQ & ~n45195;
  assign n45197 = ~n5281 & ~n45196;
  assign n45198 = i_FULL & ~n45197;
  assign n45199 = controllable_BtoR_REQ1 & ~n40638;
  assign n45200 = ~n14073 & ~n37040;
  assign n45201 = ~controllable_BtoR_REQ1 & ~n45200;
  assign n45202 = ~n45199 & ~n45201;
  assign n45203 = ~controllable_BtoR_REQ0 & ~n45202;
  assign n45204 = ~controllable_BtoR_REQ0 & ~n45203;
  assign n45205 = ~i_RtoB_ACK0 & ~n45204;
  assign n45206 = ~n45189 & ~n45205;
  assign n45207 = ~controllable_DEQ & ~n45206;
  assign n45208 = ~n5296 & ~n45207;
  assign n45209 = ~i_FULL & ~n45208;
  assign n45210 = ~n45198 & ~n45209;
  assign n45211 = ~i_nEMPTY & ~n45210;
  assign n45212 = ~n45179 & ~n45211;
  assign n45213 = controllable_BtoS_ACK0 & ~n45212;
  assign n45214 = ~i_RtoB_ACK1 & ~n37123;
  assign n45215 = ~i_RtoB_ACK1 & ~n45214;
  assign n45216 = controllable_BtoR_REQ1 & ~n45215;
  assign n45217 = ~controllable_BtoR_REQ1 & ~n12254;
  assign n45218 = ~n45216 & ~n45217;
  assign n45219 = ~controllable_BtoR_REQ0 & ~n45218;
  assign n45220 = ~controllable_BtoR_REQ0 & ~n45219;
  assign n45221 = i_RtoB_ACK0 & ~n45220;
  assign n45222 = ~controllable_BtoR_REQ1 & ~n14126;
  assign n45223 = ~n37069 & ~n45222;
  assign n45224 = ~controllable_BtoR_REQ0 & ~n45223;
  assign n45225 = ~controllable_BtoR_REQ0 & ~n45224;
  assign n45226 = ~i_RtoB_ACK0 & ~n45225;
  assign n45227 = ~n45221 & ~n45226;
  assign n45228 = ~controllable_DEQ & ~n45227;
  assign n45229 = ~n27884 & ~n45228;
  assign n45230 = i_FULL & ~n45229;
  assign n45231 = controllable_BtoR_REQ1 & ~n40661;
  assign n45232 = ~n14125 & ~n37080;
  assign n45233 = ~controllable_BtoR_REQ1 & ~n45232;
  assign n45234 = ~n45231 & ~n45233;
  assign n45235 = ~controllable_BtoR_REQ0 & ~n45234;
  assign n45236 = ~controllable_BtoR_REQ0 & ~n45235;
  assign n45237 = ~i_RtoB_ACK0 & ~n45236;
  assign n45238 = ~n45221 & ~n45237;
  assign n45239 = ~controllable_DEQ & ~n45238;
  assign n45240 = ~n27884 & ~n45239;
  assign n45241 = ~i_FULL & ~n45240;
  assign n45242 = ~n45230 & ~n45241;
  assign n45243 = i_nEMPTY & ~n45242;
  assign n45244 = controllable_ENQ & ~n37123;
  assign n45245 = controllable_ENQ & ~n45244;
  assign n45246 = ~i_RtoB_ACK1 & ~n45245;
  assign n45247 = ~i_RtoB_ACK1 & ~n45246;
  assign n45248 = controllable_BtoR_REQ1 & ~n45247;
  assign n45249 = ~controllable_BtoR_REQ1 & ~n12256;
  assign n45250 = ~n45248 & ~n45249;
  assign n45251 = ~controllable_BtoR_REQ0 & ~n45250;
  assign n45252 = ~controllable_BtoR_REQ0 & ~n45251;
  assign n45253 = i_RtoB_ACK0 & ~n45252;
  assign n45254 = ~controllable_BtoR_REQ1 & ~n14136;
  assign n45255 = ~n37104 & ~n45254;
  assign n45256 = ~controllable_BtoR_REQ0 & ~n45255;
  assign n45257 = ~controllable_BtoR_REQ0 & ~n45256;
  assign n45258 = ~i_RtoB_ACK0 & ~n45257;
  assign n45259 = ~n45253 & ~n45258;
  assign n45260 = ~controllable_DEQ & ~n45259;
  assign n45261 = ~n27900 & ~n45260;
  assign n45262 = i_FULL & ~n45261;
  assign n45263 = controllable_BtoR_REQ1 & ~n40682;
  assign n45264 = ~n14116 & ~n37126;
  assign n45265 = ~controllable_BtoR_REQ1 & ~n45264;
  assign n45266 = ~n45263 & ~n45265;
  assign n45267 = ~controllable_BtoR_REQ0 & ~n45266;
  assign n45268 = ~controllable_BtoR_REQ0 & ~n45267;
  assign n45269 = ~i_RtoB_ACK0 & ~n45268;
  assign n45270 = ~n45253 & ~n45269;
  assign n45271 = ~controllable_DEQ & ~n45270;
  assign n45272 = ~n27912 & ~n45271;
  assign n45273 = ~i_FULL & ~n45272;
  assign n45274 = ~n45262 & ~n45273;
  assign n45275 = ~i_nEMPTY & ~n45274;
  assign n45276 = ~n45243 & ~n45275;
  assign n45277 = ~controllable_BtoS_ACK0 & ~n45276;
  assign n45278 = ~n45213 & ~n45277;
  assign n45279 = n4465 & ~n45278;
  assign n45280 = ~n27884 & ~n27936;
  assign n45281 = i_FULL & ~n45280;
  assign n45282 = ~n27945 & ~n45281;
  assign n45283 = i_nEMPTY & ~n45282;
  assign n45284 = ~n27962 & ~n45283;
  assign n45285 = ~controllable_BtoS_ACK0 & ~n45284;
  assign n45286 = ~n5307 & ~n45285;
  assign n45287 = ~n4465 & ~n45286;
  assign n45288 = ~n45279 & ~n45287;
  assign n45289 = i_StoB_REQ10 & ~n45288;
  assign n45290 = ~i_RtoB_ACK1 & ~n37661;
  assign n45291 = ~n38940 & ~n45290;
  assign n45292 = controllable_BtoR_REQ1 & ~n45291;
  assign n45293 = ~n6217 & ~n9164;
  assign n45294 = n4476 & ~n45293;
  assign n45295 = ~n37271 & ~n45294;
  assign n45296 = ~i_StoB_REQ3 & ~n45295;
  assign n45297 = ~n9175 & ~n45296;
  assign n45298 = controllable_BtoS_ACK3 & ~n45297;
  assign n45299 = ~n6250 & ~n45296;
  assign n45300 = ~controllable_BtoS_ACK3 & ~n45299;
  assign n45301 = ~n45298 & ~n45300;
  assign n45302 = n4475 & ~n45301;
  assign n45303 = ~n37279 & ~n45302;
  assign n45304 = ~i_StoB_REQ4 & ~n45303;
  assign n45305 = ~n9188 & ~n45304;
  assign n45306 = controllable_BtoS_ACK4 & ~n45305;
  assign n45307 = ~n6283 & ~n45304;
  assign n45308 = ~controllable_BtoS_ACK4 & ~n45307;
  assign n45309 = ~n45306 & ~n45308;
  assign n45310 = n4474 & ~n45309;
  assign n45311 = ~n37287 & ~n45310;
  assign n45312 = ~i_StoB_REQ5 & ~n45311;
  assign n45313 = ~n9201 & ~n45312;
  assign n45314 = controllable_BtoS_ACK5 & ~n45313;
  assign n45315 = ~n6316 & ~n45312;
  assign n45316 = ~controllable_BtoS_ACK5 & ~n45315;
  assign n45317 = ~n45314 & ~n45316;
  assign n45318 = n4473 & ~n45317;
  assign n45319 = ~n37295 & ~n45318;
  assign n45320 = ~i_StoB_REQ8 & ~n45319;
  assign n45321 = ~n9214 & ~n45320;
  assign n45322 = controllable_BtoS_ACK8 & ~n45321;
  assign n45323 = ~n6341 & ~n45320;
  assign n45324 = ~controllable_BtoS_ACK8 & ~n45323;
  assign n45325 = ~n45322 & ~n45324;
  assign n45326 = n4472 & ~n45325;
  assign n45327 = ~n37303 & ~n45326;
  assign n45328 = n4471 & ~n45327;
  assign n45329 = ~n6022 & ~n45328;
  assign n45330 = ~i_StoB_REQ6 & ~n45329;
  assign n45331 = ~n38826 & ~n45330;
  assign n45332 = controllable_BtoS_ACK6 & ~n45331;
  assign n45333 = ~n6377 & ~n45330;
  assign n45334 = ~controllable_BtoS_ACK6 & ~n45333;
  assign n45335 = ~n45332 & ~n45334;
  assign n45336 = ~i_StoB_REQ7 & ~n45335;
  assign n45337 = ~n9235 & ~n45336;
  assign n45338 = controllable_BtoS_ACK7 & ~n45337;
  assign n45339 = ~n6404 & ~n45336;
  assign n45340 = ~controllable_BtoS_ACK7 & ~n45339;
  assign n45341 = ~n45338 & ~n45340;
  assign n45342 = n4470 & ~n45341;
  assign n45343 = ~n37318 & ~n45342;
  assign n45344 = n4469 & ~n45343;
  assign n45345 = ~n6095 & ~n45344;
  assign n45346 = ~i_StoB_REQ9 & ~n45345;
  assign n45347 = ~n38843 & ~n45346;
  assign n45348 = controllable_BtoS_ACK9 & ~n45347;
  assign n45349 = ~n6432 & ~n45346;
  assign n45350 = ~controllable_BtoS_ACK9 & ~n45349;
  assign n45351 = ~n45348 & ~n45350;
  assign n45352 = n4468 & ~n45351;
  assign n45353 = ~n6130 & ~n45352;
  assign n45354 = ~i_StoB_REQ11 & ~n45353;
  assign n45355 = ~n38852 & ~n45354;
  assign n45356 = controllable_BtoS_ACK11 & ~n45355;
  assign n45357 = ~n6462 & ~n45354;
  assign n45358 = ~controllable_BtoS_ACK11 & ~n45357;
  assign n45359 = ~n45356 & ~n45358;
  assign n45360 = n4467 & ~n45359;
  assign n45361 = ~n6168 & ~n45360;
  assign n45362 = ~i_StoB_REQ12 & ~n45361;
  assign n45363 = ~n38861 & ~n45362;
  assign n45364 = controllable_BtoS_ACK12 & ~n45363;
  assign n45365 = ~n6505 & ~n45362;
  assign n45366 = ~controllable_BtoS_ACK12 & ~n45365;
  assign n45367 = ~n45364 & ~n45366;
  assign n45368 = ~i_StoB_REQ13 & ~n45367;
  assign n45369 = ~n9278 & ~n45368;
  assign n45370 = n4466 & ~n45369;
  assign n45371 = ~n37448 & ~n45370;
  assign n45372 = ~i_StoB_REQ0 & ~n45371;
  assign n45373 = ~n9771 & ~n45372;
  assign n45374 = ~i_StoB_REQ14 & ~n45373;
  assign n45375 = ~n10454 & ~n45374;
  assign n45376 = controllable_BtoS_ACK14 & ~n45375;
  assign n45377 = ~n9287 & ~n45374;
  assign n45378 = ~controllable_BtoS_ACK14 & ~n45377;
  assign n45379 = ~n45376 & ~n45378;
  assign n45380 = ~controllable_BtoR_REQ1 & ~n45379;
  assign n45381 = ~n45292 & ~n45380;
  assign n45382 = ~controllable_BtoR_REQ0 & ~n45381;
  assign n45383 = ~controllable_BtoR_REQ0 & ~n45382;
  assign n45384 = i_RtoB_ACK0 & ~n45383;
  assign n45385 = controllable_BtoR_REQ1 & ~n40934;
  assign n45386 = i_RtoB_ACK1 & ~n45379;
  assign n45387 = ~n12387 & ~n45386;
  assign n45388 = ~controllable_BtoR_REQ1 & ~n45387;
  assign n45389 = ~n45385 & ~n45388;
  assign n45390 = ~controllable_BtoR_REQ0 & ~n45389;
  assign n45391 = ~controllable_BtoR_REQ0 & ~n45390;
  assign n45392 = ~i_RtoB_ACK0 & ~n45391;
  assign n45393 = ~n45384 & ~n45392;
  assign n45394 = ~controllable_DEQ & ~n45393;
  assign n45395 = ~n11244 & ~n45394;
  assign n45396 = i_FULL & ~n45395;
  assign n45397 = controllable_BtoR_REQ1 & ~n40950;
  assign n45398 = ~n37491 & ~n45386;
  assign n45399 = ~controllable_BtoR_REQ1 & ~n45398;
  assign n45400 = ~n45397 & ~n45399;
  assign n45401 = ~controllable_BtoR_REQ0 & ~n45400;
  assign n45402 = ~controllable_BtoR_REQ0 & ~n45401;
  assign n45403 = ~i_RtoB_ACK0 & ~n45402;
  assign n45404 = ~n45384 & ~n45403;
  assign n45405 = ~controllable_DEQ & ~n45404;
  assign n45406 = ~n11244 & ~n45405;
  assign n45407 = ~i_FULL & ~n45406;
  assign n45408 = ~n45396 & ~n45407;
  assign n45409 = i_nEMPTY & ~n45408;
  assign n45410 = controllable_ENQ & ~n38876;
  assign n45411 = controllable_ENQ & ~n45410;
  assign n45412 = i_RtoB_ACK1 & ~n45411;
  assign n45413 = controllable_ENQ & ~n37661;
  assign n45414 = controllable_ENQ & ~n45413;
  assign n45415 = ~i_RtoB_ACK1 & ~n45414;
  assign n45416 = ~n45412 & ~n45415;
  assign n45417 = controllable_BtoR_REQ1 & ~n45416;
  assign n45418 = controllable_ENQ & ~n45379;
  assign n45419 = controllable_ENQ & ~n45418;
  assign n45420 = ~controllable_BtoR_REQ1 & ~n45419;
  assign n45421 = ~n45417 & ~n45420;
  assign n45422 = ~controllable_BtoR_REQ0 & ~n45421;
  assign n45423 = ~controllable_BtoR_REQ0 & ~n45422;
  assign n45424 = i_RtoB_ACK0 & ~n45423;
  assign n45425 = controllable_BtoR_REQ1 & ~n40968;
  assign n45426 = i_RtoB_ACK1 & ~n45419;
  assign n45427 = ~n12431 & ~n45426;
  assign n45428 = ~controllable_BtoR_REQ1 & ~n45427;
  assign n45429 = ~n45425 & ~n45428;
  assign n45430 = ~controllable_BtoR_REQ0 & ~n45429;
  assign n45431 = ~controllable_BtoR_REQ0 & ~n45430;
  assign n45432 = ~i_RtoB_ACK0 & ~n45431;
  assign n45433 = ~n45424 & ~n45432;
  assign n45434 = ~controllable_DEQ & ~n45433;
  assign n45435 = ~n11269 & ~n45434;
  assign n45436 = i_FULL & ~n45435;
  assign n45437 = ~n37038 & ~n37525;
  assign n45438 = i_RtoB_ACK1 & ~n45437;
  assign n45439 = ~n37664 & ~n45438;
  assign n45440 = controllable_BtoR_REQ1 & ~n45439;
  assign n45441 = ~n37664 & ~n45426;
  assign n45442 = ~controllable_BtoR_REQ1 & ~n45441;
  assign n45443 = ~n45440 & ~n45442;
  assign n45444 = ~controllable_BtoR_REQ0 & ~n45443;
  assign n45445 = ~controllable_BtoR_REQ0 & ~n45444;
  assign n45446 = ~i_RtoB_ACK0 & ~n45445;
  assign n45447 = ~n45424 & ~n45446;
  assign n45448 = ~controllable_DEQ & ~n45447;
  assign n45449 = ~n11282 & ~n45448;
  assign n45450 = ~i_FULL & ~n45449;
  assign n45451 = ~n45436 & ~n45450;
  assign n45452 = ~i_nEMPTY & ~n45451;
  assign n45453 = ~n45409 & ~n45452;
  assign n45454 = controllable_BtoS_ACK0 & ~n45453;
  assign n45455 = ~i_RtoB_ACK1 & ~n37823;
  assign n45456 = ~n39035 & ~n45455;
  assign n45457 = controllable_BtoR_REQ1 & ~n45456;
  assign n45458 = ~n8058 & ~n45372;
  assign n45459 = ~i_StoB_REQ14 & ~n45458;
  assign n45460 = ~n10584 & ~n45459;
  assign n45461 = controllable_BtoS_ACK14 & ~n45460;
  assign n45462 = ~n9618 & ~n45459;
  assign n45463 = ~controllable_BtoS_ACK14 & ~n45462;
  assign n45464 = ~n45461 & ~n45463;
  assign n45465 = ~controllable_BtoR_REQ1 & ~n45464;
  assign n45466 = ~n45457 & ~n45465;
  assign n45467 = ~controllable_BtoR_REQ0 & ~n45466;
  assign n45468 = ~controllable_BtoR_REQ0 & ~n45467;
  assign n45469 = i_RtoB_ACK0 & ~n45468;
  assign n45470 = controllable_BtoR_REQ1 & ~n41005;
  assign n45471 = i_RtoB_ACK1 & ~n45464;
  assign n45472 = ~n9913 & ~n45471;
  assign n45473 = ~controllable_BtoR_REQ1 & ~n45472;
  assign n45474 = ~n45470 & ~n45473;
  assign n45475 = ~controllable_BtoR_REQ0 & ~n45474;
  assign n45476 = ~controllable_BtoR_REQ0 & ~n45475;
  assign n45477 = ~i_RtoB_ACK0 & ~n45476;
  assign n45478 = ~n45469 & ~n45477;
  assign n45479 = ~controllable_DEQ & ~n45478;
  assign n45480 = ~n11323 & ~n45479;
  assign n45481 = i_FULL & ~n45480;
  assign n45482 = controllable_BtoR_REQ1 & ~n41021;
  assign n45483 = ~n37754 & ~n45471;
  assign n45484 = ~controllable_BtoR_REQ1 & ~n45483;
  assign n45485 = ~n45482 & ~n45484;
  assign n45486 = ~controllable_BtoR_REQ0 & ~n45485;
  assign n45487 = ~controllable_BtoR_REQ0 & ~n45486;
  assign n45488 = ~i_RtoB_ACK0 & ~n45487;
  assign n45489 = ~n45469 & ~n45488;
  assign n45490 = ~controllable_DEQ & ~n45489;
  assign n45491 = ~n11323 & ~n45490;
  assign n45492 = ~i_FULL & ~n45491;
  assign n45493 = ~n45481 & ~n45492;
  assign n45494 = i_nEMPTY & ~n45493;
  assign n45495 = controllable_ENQ & ~n38971;
  assign n45496 = controllable_ENQ & ~n45495;
  assign n45497 = i_RtoB_ACK1 & ~n45496;
  assign n45498 = controllable_ENQ & ~n37823;
  assign n45499 = controllable_ENQ & ~n45498;
  assign n45500 = ~i_RtoB_ACK1 & ~n45499;
  assign n45501 = ~n45497 & ~n45500;
  assign n45502 = controllable_BtoR_REQ1 & ~n45501;
  assign n45503 = controllable_ENQ & ~n45464;
  assign n45504 = controllable_ENQ & ~n45503;
  assign n45505 = ~controllable_BtoR_REQ1 & ~n45504;
  assign n45506 = ~n45502 & ~n45505;
  assign n45507 = ~controllable_BtoR_REQ0 & ~n45506;
  assign n45508 = ~controllable_BtoR_REQ0 & ~n45507;
  assign n45509 = i_RtoB_ACK0 & ~n45508;
  assign n45510 = controllable_BtoR_REQ1 & ~n41039;
  assign n45511 = i_RtoB_ACK1 & ~n45504;
  assign n45512 = ~n9961 & ~n45511;
  assign n45513 = ~controllable_BtoR_REQ1 & ~n45512;
  assign n45514 = ~n45510 & ~n45513;
  assign n45515 = ~controllable_BtoR_REQ0 & ~n45514;
  assign n45516 = ~controllable_BtoR_REQ0 & ~n45515;
  assign n45517 = ~i_RtoB_ACK0 & ~n45516;
  assign n45518 = ~n45509 & ~n45517;
  assign n45519 = ~controllable_DEQ & ~n45518;
  assign n45520 = ~n11351 & ~n45519;
  assign n45521 = i_FULL & ~n45520;
  assign n45522 = ~n37124 & ~n37788;
  assign n45523 = i_RtoB_ACK1 & ~n45522;
  assign n45524 = ~n37826 & ~n45523;
  assign n45525 = controllable_BtoR_REQ1 & ~n45524;
  assign n45526 = ~n37826 & ~n45511;
  assign n45527 = ~controllable_BtoR_REQ1 & ~n45526;
  assign n45528 = ~n45525 & ~n45527;
  assign n45529 = ~controllable_BtoR_REQ0 & ~n45528;
  assign n45530 = ~controllable_BtoR_REQ0 & ~n45529;
  assign n45531 = ~i_RtoB_ACK0 & ~n45530;
  assign n45532 = ~n45509 & ~n45531;
  assign n45533 = ~controllable_DEQ & ~n45532;
  assign n45534 = ~n11364 & ~n45533;
  assign n45535 = ~i_FULL & ~n45534;
  assign n45536 = ~n45521 & ~n45535;
  assign n45537 = ~i_nEMPTY & ~n45536;
  assign n45538 = ~n45494 & ~n45537;
  assign n45539 = ~controllable_BtoS_ACK0 & ~n45538;
  assign n45540 = ~n45454 & ~n45539;
  assign n45541 = n4465 & ~n45540;
  assign n45542 = ~n11323 & ~n28073;
  assign n45543 = i_FULL & ~n45542;
  assign n45544 = ~n28082 & ~n45543;
  assign n45545 = i_nEMPTY & ~n45544;
  assign n45546 = ~n28101 & ~n45545;
  assign n45547 = ~controllable_BtoS_ACK0 & ~n45546;
  assign n45548 = ~n11296 & ~n45547;
  assign n45549 = ~n4465 & ~n45548;
  assign n45550 = ~n45541 & ~n45549;
  assign n45551 = ~i_StoB_REQ10 & ~n45550;
  assign n45552 = ~n45289 & ~n45551;
  assign n45553 = controllable_BtoS_ACK10 & ~n45552;
  assign n45554 = ~n14082 & ~n37915;
  assign n45555 = controllable_BtoR_REQ1 & ~n45554;
  assign n45556 = ~n11248 & ~n45555;
  assign n45557 = ~controllable_BtoR_REQ0 & ~n45556;
  assign n45558 = ~controllable_BtoR_REQ0 & ~n45557;
  assign n45559 = i_RtoB_ACK0 & ~n45558;
  assign n45560 = ~n20377 & ~n45385;
  assign n45561 = ~controllable_BtoR_REQ0 & ~n45560;
  assign n45562 = ~controllable_BtoR_REQ0 & ~n45561;
  assign n45563 = ~i_RtoB_ACK0 & ~n45562;
  assign n45564 = ~n45559 & ~n45563;
  assign n45565 = ~controllable_DEQ & ~n45564;
  assign n45566 = ~n28139 & ~n45565;
  assign n45567 = i_FULL & ~n45566;
  assign n45568 = ~n9517 & ~n37491;
  assign n45569 = ~controllable_BtoR_REQ1 & ~n45568;
  assign n45570 = ~n45397 & ~n45569;
  assign n45571 = ~controllable_BtoR_REQ0 & ~n45570;
  assign n45572 = ~controllable_BtoR_REQ0 & ~n45571;
  assign n45573 = ~i_RtoB_ACK0 & ~n45572;
  assign n45574 = ~n45559 & ~n45573;
  assign n45575 = ~controllable_DEQ & ~n45574;
  assign n45576 = ~n28139 & ~n45575;
  assign n45577 = ~i_FULL & ~n45576;
  assign n45578 = ~n45567 & ~n45577;
  assign n45579 = i_nEMPTY & ~n45578;
  assign n45580 = ~n14073 & ~n37948;
  assign n45581 = controllable_BtoR_REQ1 & ~n45580;
  assign n45582 = ~n11230 & ~n45581;
  assign n45583 = ~controllable_BtoR_REQ0 & ~n45582;
  assign n45584 = ~controllable_BtoR_REQ0 & ~n45583;
  assign n45585 = i_RtoB_ACK0 & ~n45584;
  assign n45586 = ~n20411 & ~n45425;
  assign n45587 = ~controllable_BtoR_REQ0 & ~n45586;
  assign n45588 = ~controllable_BtoR_REQ0 & ~n45587;
  assign n45589 = ~i_RtoB_ACK0 & ~n45588;
  assign n45590 = ~n45585 & ~n45589;
  assign n45591 = ~controllable_DEQ & ~n45590;
  assign n45592 = ~n28153 & ~n45591;
  assign n45593 = i_FULL & ~n45592;
  assign n45594 = ~n36897 & ~n37525;
  assign n45595 = i_RtoB_ACK1 & ~n45594;
  assign n45596 = ~n37491 & ~n45595;
  assign n45597 = controllable_BtoR_REQ1 & ~n45596;
  assign n45598 = ~n9571 & ~n37491;
  assign n45599 = ~controllable_BtoR_REQ1 & ~n45598;
  assign n45600 = ~n45597 & ~n45599;
  assign n45601 = ~controllable_BtoR_REQ0 & ~n45600;
  assign n45602 = ~controllable_BtoR_REQ0 & ~n45601;
  assign n45603 = ~i_RtoB_ACK0 & ~n45602;
  assign n45604 = ~n45585 & ~n45603;
  assign n45605 = ~controllable_DEQ & ~n45604;
  assign n45606 = ~n28163 & ~n45605;
  assign n45607 = ~i_FULL & ~n45606;
  assign n45608 = ~n45593 & ~n45607;
  assign n45609 = ~i_nEMPTY & ~n45608;
  assign n45610 = ~n45579 & ~n45609;
  assign n45611 = controllable_BtoS_ACK0 & ~n45610;
  assign n45612 = ~n14125 & ~n37999;
  assign n45613 = controllable_BtoR_REQ1 & ~n45612;
  assign n45614 = ~n11328 & ~n45613;
  assign n45615 = ~controllable_BtoR_REQ0 & ~n45614;
  assign n45616 = ~controllable_BtoR_REQ0 & ~n45615;
  assign n45617 = i_RtoB_ACK0 & ~n45616;
  assign n45618 = ~n19321 & ~n45470;
  assign n45619 = ~controllable_BtoR_REQ0 & ~n45618;
  assign n45620 = ~controllable_BtoR_REQ0 & ~n45619;
  assign n45621 = ~i_RtoB_ACK0 & ~n45620;
  assign n45622 = ~n45617 & ~n45621;
  assign n45623 = ~controllable_DEQ & ~n45622;
  assign n45624 = ~n28200 & ~n45623;
  assign n45625 = i_FULL & ~n45624;
  assign n45626 = ~n9664 & ~n37754;
  assign n45627 = ~controllable_BtoR_REQ1 & ~n45626;
  assign n45628 = ~n45482 & ~n45627;
  assign n45629 = ~controllable_BtoR_REQ0 & ~n45628;
  assign n45630 = ~controllable_BtoR_REQ0 & ~n45629;
  assign n45631 = ~i_RtoB_ACK0 & ~n45630;
  assign n45632 = ~n45617 & ~n45631;
  assign n45633 = ~controllable_DEQ & ~n45632;
  assign n45634 = ~n28200 & ~n45633;
  assign n45635 = ~i_FULL & ~n45634;
  assign n45636 = ~n45625 & ~n45635;
  assign n45637 = i_nEMPTY & ~n45636;
  assign n45638 = ~n14116 & ~n38032;
  assign n45639 = controllable_BtoR_REQ1 & ~n45638;
  assign n45640 = ~n11305 & ~n45639;
  assign n45641 = ~controllable_BtoR_REQ0 & ~n45640;
  assign n45642 = ~controllable_BtoR_REQ0 & ~n45641;
  assign n45643 = i_RtoB_ACK0 & ~n45642;
  assign n45644 = ~n19351 & ~n45510;
  assign n45645 = ~controllable_BtoR_REQ0 & ~n45644;
  assign n45646 = ~controllable_BtoR_REQ0 & ~n45645;
  assign n45647 = ~i_RtoB_ACK0 & ~n45646;
  assign n45648 = ~n45643 & ~n45647;
  assign n45649 = ~controllable_DEQ & ~n45648;
  assign n45650 = ~n28214 & ~n45649;
  assign n45651 = i_FULL & ~n45650;
  assign n45652 = ~n37078 & ~n37788;
  assign n45653 = i_RtoB_ACK1 & ~n45652;
  assign n45654 = ~n37754 & ~n45653;
  assign n45655 = controllable_BtoR_REQ1 & ~n45654;
  assign n45656 = ~n9718 & ~n37754;
  assign n45657 = ~controllable_BtoR_REQ1 & ~n45656;
  assign n45658 = ~n45655 & ~n45657;
  assign n45659 = ~controllable_BtoR_REQ0 & ~n45658;
  assign n45660 = ~controllable_BtoR_REQ0 & ~n45659;
  assign n45661 = ~i_RtoB_ACK0 & ~n45660;
  assign n45662 = ~n45643 & ~n45661;
  assign n45663 = ~controllable_DEQ & ~n45662;
  assign n45664 = ~n28224 & ~n45663;
  assign n45665 = ~i_FULL & ~n45664;
  assign n45666 = ~n45651 & ~n45665;
  assign n45667 = ~i_nEMPTY & ~n45666;
  assign n45668 = ~n45637 & ~n45667;
  assign n45669 = ~controllable_BtoS_ACK0 & ~n45668;
  assign n45670 = ~n45611 & ~n45669;
  assign n45671 = n4465 & ~n45670;
  assign n45672 = ~n28200 & ~n28258;
  assign n45673 = i_FULL & ~n45672;
  assign n45674 = ~n28264 & ~n45673;
  assign n45675 = i_nEMPTY & ~n45674;
  assign n45676 = ~n28275 & ~n45675;
  assign n45677 = ~controllable_BtoS_ACK0 & ~n45676;
  assign n45678 = ~n28248 & ~n45677;
  assign n45679 = ~n4465 & ~n45678;
  assign n45680 = ~n45671 & ~n45679;
  assign n45681 = i_StoB_REQ10 & ~n45680;
  assign n45682 = ~n45551 & ~n45681;
  assign n45683 = ~controllable_BtoS_ACK10 & ~n45682;
  assign n45684 = ~n45553 & ~n45683;
  assign n45685 = n4464 & ~n45684;
  assign n45686 = ~n5251 & ~n28296;
  assign n45687 = i_FULL & ~n45686;
  assign n45688 = ~n28305 & ~n45687;
  assign n45689 = i_nEMPTY & ~n45688;
  assign n45690 = ~n28322 & ~n45689;
  assign n45691 = controllable_BtoS_ACK0 & ~n45690;
  assign n45692 = ~n27884 & ~n28335;
  assign n45693 = i_FULL & ~n45692;
  assign n45694 = ~n28344 & ~n45693;
  assign n45695 = i_nEMPTY & ~n45694;
  assign n45696 = ~n28361 & ~n45695;
  assign n45697 = ~controllable_BtoS_ACK0 & ~n45696;
  assign n45698 = ~n45691 & ~n45697;
  assign n45699 = n4465 & ~n45698;
  assign n45700 = ~n5307 & ~n45697;
  assign n45701 = ~n4465 & ~n45700;
  assign n45702 = ~n45699 & ~n45701;
  assign n45703 = i_StoB_REQ10 & ~n45702;
  assign n45704 = ~n11244 & ~n28382;
  assign n45705 = i_FULL & ~n45704;
  assign n45706 = ~n28391 & ~n45705;
  assign n45707 = i_nEMPTY & ~n45706;
  assign n45708 = ~n28410 & ~n45707;
  assign n45709 = controllable_BtoS_ACK0 & ~n45708;
  assign n45710 = ~n11323 & ~n28425;
  assign n45711 = i_FULL & ~n45710;
  assign n45712 = ~n28434 & ~n45711;
  assign n45713 = i_nEMPTY & ~n45712;
  assign n45714 = ~n28453 & ~n45713;
  assign n45715 = ~controllable_BtoS_ACK0 & ~n45714;
  assign n45716 = ~n45709 & ~n45715;
  assign n45717 = n4465 & ~n45716;
  assign n45718 = ~n11296 & ~n45715;
  assign n45719 = ~n4465 & ~n45718;
  assign n45720 = ~n45717 & ~n45719;
  assign n45721 = ~i_StoB_REQ10 & ~n45720;
  assign n45722 = ~n45703 & ~n45721;
  assign n45723 = controllable_BtoS_ACK10 & ~n45722;
  assign n45724 = ~n28139 & ~n28473;
  assign n45725 = i_FULL & ~n45724;
  assign n45726 = ~n28479 & ~n45725;
  assign n45727 = i_nEMPTY & ~n45726;
  assign n45728 = ~n28490 & ~n45727;
  assign n45729 = controllable_BtoS_ACK0 & ~n45728;
  assign n45730 = ~n28200 & ~n28502;
  assign n45731 = i_FULL & ~n45730;
  assign n45732 = ~n28508 & ~n45731;
  assign n45733 = i_nEMPTY & ~n45732;
  assign n45734 = ~n28519 & ~n45733;
  assign n45735 = ~controllable_BtoS_ACK0 & ~n45734;
  assign n45736 = ~n45729 & ~n45735;
  assign n45737 = n4465 & ~n45736;
  assign n45738 = ~n28248 & ~n45735;
  assign n45739 = ~n4465 & ~n45738;
  assign n45740 = ~n45737 & ~n45739;
  assign n45741 = i_StoB_REQ10 & ~n45740;
  assign n45742 = ~n45721 & ~n45741;
  assign n45743 = ~controllable_BtoS_ACK10 & ~n45742;
  assign n45744 = ~n45723 & ~n45743;
  assign n45745 = ~n4464 & ~n45744;
  assign n45746 = ~n45685 & ~n45745;
  assign n45747 = n4463 & ~n45746;
  assign n45748 = ~n5254 & ~n45153;
  assign n45749 = ~controllable_BtoR_REQ0 & ~n45748;
  assign n45750 = ~controllable_BtoR_REQ0 & ~n45749;
  assign n45751 = i_RtoB_ACK0 & ~n45750;
  assign n45752 = ~n14082 & ~n36879;
  assign n45753 = ~controllable_BtoR_REQ0 & ~n45752;
  assign n45754 = ~controllable_BtoR_REQ0 & ~n45753;
  assign n45755 = ~i_RtoB_ACK0 & ~n45754;
  assign n45756 = ~n45751 & ~n45755;
  assign n45757 = ~controllable_DEQ & ~n45756;
  assign n45758 = ~n5251 & ~n45757;
  assign n45759 = i_nEMPTY & ~n45758;
  assign n45760 = ~n5224 & ~n45185;
  assign n45761 = ~controllable_BtoR_REQ0 & ~n45760;
  assign n45762 = ~controllable_BtoR_REQ0 & ~n45761;
  assign n45763 = i_RtoB_ACK0 & ~n45762;
  assign n45764 = ~n14073 & ~n36914;
  assign n45765 = ~controllable_BtoR_REQ0 & ~n45764;
  assign n45766 = ~controllable_BtoR_REQ0 & ~n45765;
  assign n45767 = ~i_RtoB_ACK0 & ~n45766;
  assign n45768 = ~n45763 & ~n45767;
  assign n45769 = ~controllable_DEQ & ~n45768;
  assign n45770 = ~n5281 & ~n45769;
  assign n45771 = i_FULL & ~n45770;
  assign n45772 = ~n36912 & ~n37038;
  assign n45773 = ~i_RtoB_ACK1 & ~n45772;
  assign n45774 = ~n14073 & ~n45773;
  assign n45775 = ~controllable_BtoR_REQ0 & ~n45774;
  assign n45776 = ~controllable_BtoR_REQ0 & ~n45775;
  assign n45777 = ~i_RtoB_ACK0 & ~n45776;
  assign n45778 = ~n45763 & ~n45777;
  assign n45779 = ~controllable_DEQ & ~n45778;
  assign n45780 = ~n5296 & ~n45779;
  assign n45781 = ~i_FULL & ~n45780;
  assign n45782 = ~n45771 & ~n45781;
  assign n45783 = ~i_nEMPTY & ~n45782;
  assign n45784 = ~n45759 & ~n45783;
  assign n45785 = controllable_BtoS_ACK0 & ~n45784;
  assign n45786 = ~n27867 & ~n45217;
  assign n45787 = ~controllable_BtoR_REQ0 & ~n45786;
  assign n45788 = ~controllable_BtoR_REQ0 & ~n45787;
  assign n45789 = i_RtoB_ACK0 & ~n45788;
  assign n45790 = ~n14125 & ~n37060;
  assign n45791 = ~controllable_BtoR_REQ0 & ~n45790;
  assign n45792 = ~controllable_BtoR_REQ0 & ~n45791;
  assign n45793 = ~i_RtoB_ACK0 & ~n45792;
  assign n45794 = ~n45789 & ~n45793;
  assign n45795 = ~controllable_DEQ & ~n45794;
  assign n45796 = ~n27884 & ~n45795;
  assign n45797 = i_nEMPTY & ~n45796;
  assign n45798 = ~n27855 & ~n45249;
  assign n45799 = ~controllable_BtoR_REQ0 & ~n45798;
  assign n45800 = ~controllable_BtoR_REQ0 & ~n45799;
  assign n45801 = i_RtoB_ACK0 & ~n45800;
  assign n45802 = ~n14116 & ~n37095;
  assign n45803 = ~controllable_BtoR_REQ0 & ~n45802;
  assign n45804 = ~controllable_BtoR_REQ0 & ~n45803;
  assign n45805 = ~i_RtoB_ACK0 & ~n45804;
  assign n45806 = ~n45801 & ~n45805;
  assign n45807 = ~controllable_DEQ & ~n45806;
  assign n45808 = ~n27900 & ~n45807;
  assign n45809 = i_FULL & ~n45808;
  assign n45810 = ~n37093 & ~n37124;
  assign n45811 = ~i_RtoB_ACK1 & ~n45810;
  assign n45812 = ~n14116 & ~n45811;
  assign n45813 = ~controllable_BtoR_REQ0 & ~n45812;
  assign n45814 = ~controllable_BtoR_REQ0 & ~n45813;
  assign n45815 = ~i_RtoB_ACK0 & ~n45814;
  assign n45816 = ~n45801 & ~n45815;
  assign n45817 = ~controllable_DEQ & ~n45816;
  assign n45818 = ~n27912 & ~n45817;
  assign n45819 = ~i_FULL & ~n45818;
  assign n45820 = ~n45809 & ~n45819;
  assign n45821 = ~i_nEMPTY & ~n45820;
  assign n45822 = ~n45797 & ~n45821;
  assign n45823 = ~controllable_BtoS_ACK0 & ~n45822;
  assign n45824 = ~n45785 & ~n45823;
  assign n45825 = n4465 & ~n45824;
  assign n45826 = ~n4465 & ~n28559;
  assign n45827 = ~n45825 & ~n45826;
  assign n45828 = i_StoB_REQ10 & ~n45827;
  assign n45829 = ~n11247 & ~n45380;
  assign n45830 = ~controllable_BtoR_REQ0 & ~n45829;
  assign n45831 = ~controllable_BtoR_REQ0 & ~n45830;
  assign n45832 = i_RtoB_ACK0 & ~n45831;
  assign n45833 = ~n37915 & ~n45386;
  assign n45834 = ~controllable_BtoR_REQ0 & ~n45833;
  assign n45835 = ~controllable_BtoR_REQ0 & ~n45834;
  assign n45836 = ~i_RtoB_ACK0 & ~n45835;
  assign n45837 = ~n45832 & ~n45836;
  assign n45838 = ~controllable_DEQ & ~n45837;
  assign n45839 = ~n11244 & ~n45838;
  assign n45840 = i_nEMPTY & ~n45839;
  assign n45841 = ~n11229 & ~n45420;
  assign n45842 = ~controllable_BtoR_REQ0 & ~n45841;
  assign n45843 = ~controllable_BtoR_REQ0 & ~n45842;
  assign n45844 = i_RtoB_ACK0 & ~n45843;
  assign n45845 = ~n37948 & ~n45426;
  assign n45846 = ~controllable_BtoR_REQ0 & ~n45845;
  assign n45847 = ~controllable_BtoR_REQ0 & ~n45846;
  assign n45848 = ~i_RtoB_ACK0 & ~n45847;
  assign n45849 = ~n45844 & ~n45848;
  assign n45850 = ~controllable_DEQ & ~n45849;
  assign n45851 = ~n11269 & ~n45850;
  assign n45852 = i_FULL & ~n45851;
  assign n45853 = ~n38877 & ~n45418;
  assign n45854 = i_RtoB_ACK1 & ~n45853;
  assign n45855 = ~n37525 & ~n37662;
  assign n45856 = ~i_RtoB_ACK1 & ~n45855;
  assign n45857 = ~n45854 & ~n45856;
  assign n45858 = controllable_BtoR_REQ1 & ~n45857;
  assign n45859 = ~n45426 & ~n45856;
  assign n45860 = ~controllable_BtoR_REQ1 & ~n45859;
  assign n45861 = ~n45858 & ~n45860;
  assign n45862 = ~controllable_BtoR_REQ0 & ~n45861;
  assign n45863 = ~controllable_BtoR_REQ0 & ~n45862;
  assign n45864 = ~i_RtoB_ACK0 & ~n45863;
  assign n45865 = ~n45844 & ~n45864;
  assign n45866 = ~controllable_DEQ & ~n45865;
  assign n45867 = ~n11282 & ~n45866;
  assign n45868 = ~i_FULL & ~n45867;
  assign n45869 = ~n45852 & ~n45868;
  assign n45870 = ~i_nEMPTY & ~n45869;
  assign n45871 = ~n45840 & ~n45870;
  assign n45872 = controllable_BtoS_ACK0 & ~n45871;
  assign n45873 = ~n11327 & ~n45465;
  assign n45874 = ~controllable_BtoR_REQ0 & ~n45873;
  assign n45875 = ~controllable_BtoR_REQ0 & ~n45874;
  assign n45876 = i_RtoB_ACK0 & ~n45875;
  assign n45877 = ~n37999 & ~n45471;
  assign n45878 = ~controllable_BtoR_REQ0 & ~n45877;
  assign n45879 = ~controllable_BtoR_REQ0 & ~n45878;
  assign n45880 = ~i_RtoB_ACK0 & ~n45879;
  assign n45881 = ~n45876 & ~n45880;
  assign n45882 = ~controllable_DEQ & ~n45881;
  assign n45883 = ~n11323 & ~n45882;
  assign n45884 = i_nEMPTY & ~n45883;
  assign n45885 = ~n11304 & ~n45505;
  assign n45886 = ~controllable_BtoR_REQ0 & ~n45885;
  assign n45887 = ~controllable_BtoR_REQ0 & ~n45886;
  assign n45888 = i_RtoB_ACK0 & ~n45887;
  assign n45889 = ~n38032 & ~n45511;
  assign n45890 = ~controllable_BtoR_REQ0 & ~n45889;
  assign n45891 = ~controllable_BtoR_REQ0 & ~n45890;
  assign n45892 = ~i_RtoB_ACK0 & ~n45891;
  assign n45893 = ~n45888 & ~n45892;
  assign n45894 = ~controllable_DEQ & ~n45893;
  assign n45895 = ~n11351 & ~n45894;
  assign n45896 = i_FULL & ~n45895;
  assign n45897 = ~n38972 & ~n45503;
  assign n45898 = i_RtoB_ACK1 & ~n45897;
  assign n45899 = ~n37788 & ~n37824;
  assign n45900 = ~i_RtoB_ACK1 & ~n45899;
  assign n45901 = ~n45898 & ~n45900;
  assign n45902 = controllable_BtoR_REQ1 & ~n45901;
  assign n45903 = ~n45511 & ~n45900;
  assign n45904 = ~controllable_BtoR_REQ1 & ~n45903;
  assign n45905 = ~n45902 & ~n45904;
  assign n45906 = ~controllable_BtoR_REQ0 & ~n45905;
  assign n45907 = ~controllable_BtoR_REQ0 & ~n45906;
  assign n45908 = ~i_RtoB_ACK0 & ~n45907;
  assign n45909 = ~n45888 & ~n45908;
  assign n45910 = ~controllable_DEQ & ~n45909;
  assign n45911 = ~n11364 & ~n45910;
  assign n45912 = ~i_FULL & ~n45911;
  assign n45913 = ~n45896 & ~n45912;
  assign n45914 = ~i_nEMPTY & ~n45913;
  assign n45915 = ~n45884 & ~n45914;
  assign n45916 = ~controllable_BtoS_ACK0 & ~n45915;
  assign n45917 = ~n45872 & ~n45916;
  assign n45918 = n4465 & ~n45917;
  assign n45919 = ~n4465 & ~n11379;
  assign n45920 = ~n45918 & ~n45919;
  assign n45921 = ~i_StoB_REQ10 & ~n45920;
  assign n45922 = ~n45828 & ~n45921;
  assign n45923 = controllable_BtoS_ACK10 & ~n45922;
  assign n45924 = ~n9517 & ~n37915;
  assign n45925 = ~controllable_BtoR_REQ0 & ~n45924;
  assign n45926 = ~controllable_BtoR_REQ0 & ~n45925;
  assign n45927 = ~i_RtoB_ACK0 & ~n45926;
  assign n45928 = ~n28127 & ~n45927;
  assign n45929 = ~controllable_DEQ & ~n45928;
  assign n45930 = ~n28139 & ~n45929;
  assign n45931 = i_nEMPTY & ~n45930;
  assign n45932 = ~n9571 & ~n37948;
  assign n45933 = ~controllable_BtoR_REQ0 & ~n45932;
  assign n45934 = ~controllable_BtoR_REQ0 & ~n45933;
  assign n45935 = ~i_RtoB_ACK0 & ~n45934;
  assign n45936 = ~n28114 & ~n45935;
  assign n45937 = ~controllable_DEQ & ~n45936;
  assign n45938 = ~n28153 & ~n45937;
  assign n45939 = i_FULL & ~n45938;
  assign n45940 = ~n37915 & ~n39107;
  assign n45941 = controllable_BtoR_REQ1 & ~n45940;
  assign n45942 = ~n9571 & ~n37915;
  assign n45943 = ~controllable_BtoR_REQ1 & ~n45942;
  assign n45944 = ~n45941 & ~n45943;
  assign n45945 = ~controllable_BtoR_REQ0 & ~n45944;
  assign n45946 = ~controllable_BtoR_REQ0 & ~n45945;
  assign n45947 = ~i_RtoB_ACK0 & ~n45946;
  assign n45948 = ~n28114 & ~n45947;
  assign n45949 = ~controllable_DEQ & ~n45948;
  assign n45950 = ~n28163 & ~n45949;
  assign n45951 = ~i_FULL & ~n45950;
  assign n45952 = ~n45939 & ~n45951;
  assign n45953 = ~i_nEMPTY & ~n45952;
  assign n45954 = ~n45931 & ~n45953;
  assign n45955 = controllable_BtoS_ACK0 & ~n45954;
  assign n45956 = ~n9664 & ~n37999;
  assign n45957 = ~controllable_BtoR_REQ0 & ~n45956;
  assign n45958 = ~controllable_BtoR_REQ0 & ~n45957;
  assign n45959 = ~i_RtoB_ACK0 & ~n45958;
  assign n45960 = ~n28188 & ~n45959;
  assign n45961 = ~controllable_DEQ & ~n45960;
  assign n45962 = ~n28200 & ~n45961;
  assign n45963 = i_nEMPTY & ~n45962;
  assign n45964 = ~n9718 & ~n38032;
  assign n45965 = ~controllable_BtoR_REQ0 & ~n45964;
  assign n45966 = ~controllable_BtoR_REQ0 & ~n45965;
  assign n45967 = ~i_RtoB_ACK0 & ~n45966;
  assign n45968 = ~n28175 & ~n45967;
  assign n45969 = ~controllable_DEQ & ~n45968;
  assign n45970 = ~n28214 & ~n45969;
  assign n45971 = i_FULL & ~n45970;
  assign n45972 = ~n37999 & ~n39180;
  assign n45973 = controllable_BtoR_REQ1 & ~n45972;
  assign n45974 = ~n9718 & ~n37999;
  assign n45975 = ~controllable_BtoR_REQ1 & ~n45974;
  assign n45976 = ~n45973 & ~n45975;
  assign n45977 = ~controllable_BtoR_REQ0 & ~n45976;
  assign n45978 = ~controllable_BtoR_REQ0 & ~n45977;
  assign n45979 = ~i_RtoB_ACK0 & ~n45978;
  assign n45980 = ~n28175 & ~n45979;
  assign n45981 = ~controllable_DEQ & ~n45980;
  assign n45982 = ~n28224 & ~n45981;
  assign n45983 = ~i_FULL & ~n45982;
  assign n45984 = ~n45971 & ~n45983;
  assign n45985 = ~i_nEMPTY & ~n45984;
  assign n45986 = ~n45963 & ~n45985;
  assign n45987 = ~controllable_BtoS_ACK0 & ~n45986;
  assign n45988 = ~n45955 & ~n45987;
  assign n45989 = n4465 & ~n45988;
  assign n45990 = ~n4465 & ~n28578;
  assign n45991 = ~n45989 & ~n45990;
  assign n45992 = i_StoB_REQ10 & ~n45991;
  assign n45993 = ~n45921 & ~n45992;
  assign n45994 = ~controllable_BtoS_ACK10 & ~n45993;
  assign n45995 = ~n45923 & ~n45994;
  assign n45996 = n4464 & ~n45995;
  assign n45997 = ~n4464 & ~n28582;
  assign n45998 = ~n45996 & ~n45997;
  assign n45999 = ~n4463 & ~n45998;
  assign n46000 = ~n45747 & ~n45999;
  assign n46001 = n4462 & ~n46000;
  assign n46002 = ~n28139 & ~n28598;
  assign n46003 = i_FULL & ~n46002;
  assign n46004 = ~n28607 & ~n46003;
  assign n46005 = i_nEMPTY & ~n46004;
  assign n46006 = ~n28621 & ~n46005;
  assign n46007 = controllable_BtoS_ACK0 & ~n46006;
  assign n46008 = ~n45677 & ~n46007;
  assign n46009 = n4465 & ~n46008;
  assign n46010 = ~n45679 & ~n46009;
  assign n46011 = i_StoB_REQ10 & ~n46010;
  assign n46012 = ~n11244 & ~n28637;
  assign n46013 = i_FULL & ~n46012;
  assign n46014 = ~n28643 & ~n46013;
  assign n46015 = i_nEMPTY & ~n46014;
  assign n46016 = ~n28659 & ~n46015;
  assign n46017 = controllable_BtoS_ACK0 & ~n46016;
  assign n46018 = ~n45547 & ~n46017;
  assign n46019 = n4465 & ~n46018;
  assign n46020 = ~n45549 & ~n46019;
  assign n46021 = ~i_StoB_REQ10 & ~n46020;
  assign n46022 = ~n46011 & ~n46021;
  assign n46023 = ~controllable_BtoS_ACK10 & ~n46022;
  assign n46024 = ~n28562 & ~n46023;
  assign n46025 = n4464 & ~n46024;
  assign n46026 = ~n28562 & ~n45743;
  assign n46027 = ~n4464 & ~n46026;
  assign n46028 = ~n46025 & ~n46027;
  assign n46029 = n4463 & ~n46028;
  assign n46030 = ~n28583 & ~n46029;
  assign n46031 = ~n4462 & ~n46030;
  assign n46032 = ~n46001 & ~n46031;
  assign n46033 = n4461 & ~n46032;
  assign n46034 = ~controllable_BtoR_REQ0 & ~n14083;
  assign n46035 = ~controllable_BtoR_REQ0 & ~n46034;
  assign n46036 = ~i_RtoB_ACK0 & ~n46035;
  assign n46037 = ~n45157 & ~n46036;
  assign n46038 = ~controllable_DEQ & ~n46037;
  assign n46039 = ~n5251 & ~n46038;
  assign n46040 = i_FULL & ~n46039;
  assign n46041 = ~controllable_BtoR_REQ0 & ~n45168;
  assign n46042 = ~controllable_BtoR_REQ0 & ~n46041;
  assign n46043 = ~i_RtoB_ACK0 & ~n46042;
  assign n46044 = ~n45157 & ~n46043;
  assign n46045 = ~controllable_DEQ & ~n46044;
  assign n46046 = ~n5251 & ~n46045;
  assign n46047 = ~i_FULL & ~n46046;
  assign n46048 = ~n46040 & ~n46047;
  assign n46049 = i_nEMPTY & ~n46048;
  assign n46050 = ~controllable_BtoR_REQ0 & ~n14093;
  assign n46051 = ~controllable_BtoR_REQ0 & ~n46050;
  assign n46052 = ~i_RtoB_ACK0 & ~n46051;
  assign n46053 = ~n45189 & ~n46052;
  assign n46054 = ~controllable_DEQ & ~n46053;
  assign n46055 = ~n5281 & ~n46054;
  assign n46056 = i_FULL & ~n46055;
  assign n46057 = ~controllable_BtoR_REQ0 & ~n45200;
  assign n46058 = ~controllable_BtoR_REQ0 & ~n46057;
  assign n46059 = ~i_RtoB_ACK0 & ~n46058;
  assign n46060 = ~n45189 & ~n46059;
  assign n46061 = ~controllable_DEQ & ~n46060;
  assign n46062 = ~n5296 & ~n46061;
  assign n46063 = ~i_FULL & ~n46062;
  assign n46064 = ~n46056 & ~n46063;
  assign n46065 = ~i_nEMPTY & ~n46064;
  assign n46066 = ~n46049 & ~n46065;
  assign n46067 = controllable_BtoS_ACK0 & ~n46066;
  assign n46068 = ~controllable_BtoR_REQ0 & ~n14126;
  assign n46069 = ~controllable_BtoR_REQ0 & ~n46068;
  assign n46070 = ~i_RtoB_ACK0 & ~n46069;
  assign n46071 = ~n45221 & ~n46070;
  assign n46072 = ~controllable_DEQ & ~n46071;
  assign n46073 = ~n27884 & ~n46072;
  assign n46074 = i_FULL & ~n46073;
  assign n46075 = ~controllable_BtoR_REQ0 & ~n45232;
  assign n46076 = ~controllable_BtoR_REQ0 & ~n46075;
  assign n46077 = ~i_RtoB_ACK0 & ~n46076;
  assign n46078 = ~n45221 & ~n46077;
  assign n46079 = ~controllable_DEQ & ~n46078;
  assign n46080 = ~n27884 & ~n46079;
  assign n46081 = ~i_FULL & ~n46080;
  assign n46082 = ~n46074 & ~n46081;
  assign n46083 = i_nEMPTY & ~n46082;
  assign n46084 = ~controllable_BtoR_REQ0 & ~n14136;
  assign n46085 = ~controllable_BtoR_REQ0 & ~n46084;
  assign n46086 = ~i_RtoB_ACK0 & ~n46085;
  assign n46087 = ~n45253 & ~n46086;
  assign n46088 = ~controllable_DEQ & ~n46087;
  assign n46089 = ~n27900 & ~n46088;
  assign n46090 = i_FULL & ~n46089;
  assign n46091 = ~controllable_BtoR_REQ0 & ~n45264;
  assign n46092 = ~controllable_BtoR_REQ0 & ~n46091;
  assign n46093 = ~i_RtoB_ACK0 & ~n46092;
  assign n46094 = ~n45253 & ~n46093;
  assign n46095 = ~controllable_DEQ & ~n46094;
  assign n46096 = ~n27912 & ~n46095;
  assign n46097 = ~i_FULL & ~n46096;
  assign n46098 = ~n46090 & ~n46097;
  assign n46099 = ~i_nEMPTY & ~n46098;
  assign n46100 = ~n46083 & ~n46099;
  assign n46101 = ~controllable_BtoS_ACK0 & ~n46100;
  assign n46102 = ~n46067 & ~n46101;
  assign n46103 = n4465 & ~n46102;
  assign n46104 = ~n45287 & ~n46103;
  assign n46105 = i_StoB_REQ10 & ~n46104;
  assign n46106 = ~controllable_BtoR_REQ0 & ~n45387;
  assign n46107 = ~controllable_BtoR_REQ0 & ~n46106;
  assign n46108 = ~i_RtoB_ACK0 & ~n46107;
  assign n46109 = ~n45384 & ~n46108;
  assign n46110 = ~controllable_DEQ & ~n46109;
  assign n46111 = ~n11244 & ~n46110;
  assign n46112 = i_FULL & ~n46111;
  assign n46113 = ~controllable_BtoR_REQ0 & ~n45398;
  assign n46114 = ~controllable_BtoR_REQ0 & ~n46113;
  assign n46115 = ~i_RtoB_ACK0 & ~n46114;
  assign n46116 = ~n45384 & ~n46115;
  assign n46117 = ~controllable_DEQ & ~n46116;
  assign n46118 = ~n11244 & ~n46117;
  assign n46119 = ~i_FULL & ~n46118;
  assign n46120 = ~n46112 & ~n46119;
  assign n46121 = i_nEMPTY & ~n46120;
  assign n46122 = ~controllable_BtoR_REQ0 & ~n45427;
  assign n46123 = ~controllable_BtoR_REQ0 & ~n46122;
  assign n46124 = ~i_RtoB_ACK0 & ~n46123;
  assign n46125 = ~n45424 & ~n46124;
  assign n46126 = ~controllable_DEQ & ~n46125;
  assign n46127 = ~n11269 & ~n46126;
  assign n46128 = i_FULL & ~n46127;
  assign n46129 = ~n37664 & ~n45854;
  assign n46130 = controllable_BtoR_REQ1 & ~n46129;
  assign n46131 = ~n45442 & ~n46130;
  assign n46132 = ~controllable_BtoR_REQ0 & ~n46131;
  assign n46133 = ~controllable_BtoR_REQ0 & ~n46132;
  assign n46134 = ~i_RtoB_ACK0 & ~n46133;
  assign n46135 = ~n45424 & ~n46134;
  assign n46136 = ~controllable_DEQ & ~n46135;
  assign n46137 = ~n11282 & ~n46136;
  assign n46138 = ~i_FULL & ~n46137;
  assign n46139 = ~n46128 & ~n46138;
  assign n46140 = ~i_nEMPTY & ~n46139;
  assign n46141 = ~n46121 & ~n46140;
  assign n46142 = controllable_BtoS_ACK0 & ~n46141;
  assign n46143 = ~controllable_BtoR_REQ0 & ~n45472;
  assign n46144 = ~controllable_BtoR_REQ0 & ~n46143;
  assign n46145 = ~i_RtoB_ACK0 & ~n46144;
  assign n46146 = ~n45469 & ~n46145;
  assign n46147 = ~controllable_DEQ & ~n46146;
  assign n46148 = ~n11323 & ~n46147;
  assign n46149 = i_FULL & ~n46148;
  assign n46150 = ~controllable_BtoR_REQ0 & ~n45483;
  assign n46151 = ~controllable_BtoR_REQ0 & ~n46150;
  assign n46152 = ~i_RtoB_ACK0 & ~n46151;
  assign n46153 = ~n45469 & ~n46152;
  assign n46154 = ~controllable_DEQ & ~n46153;
  assign n46155 = ~n11323 & ~n46154;
  assign n46156 = ~i_FULL & ~n46155;
  assign n46157 = ~n46149 & ~n46156;
  assign n46158 = i_nEMPTY & ~n46157;
  assign n46159 = ~controllable_BtoR_REQ0 & ~n45512;
  assign n46160 = ~controllable_BtoR_REQ0 & ~n46159;
  assign n46161 = ~i_RtoB_ACK0 & ~n46160;
  assign n46162 = ~n45509 & ~n46161;
  assign n46163 = ~controllable_DEQ & ~n46162;
  assign n46164 = ~n11351 & ~n46163;
  assign n46165 = i_FULL & ~n46164;
  assign n46166 = ~n37826 & ~n45898;
  assign n46167 = controllable_BtoR_REQ1 & ~n46166;
  assign n46168 = ~n45527 & ~n46167;
  assign n46169 = ~controllable_BtoR_REQ0 & ~n46168;
  assign n46170 = ~controllable_BtoR_REQ0 & ~n46169;
  assign n46171 = ~i_RtoB_ACK0 & ~n46170;
  assign n46172 = ~n45509 & ~n46171;
  assign n46173 = ~controllable_DEQ & ~n46172;
  assign n46174 = ~n11364 & ~n46173;
  assign n46175 = ~i_FULL & ~n46174;
  assign n46176 = ~n46165 & ~n46175;
  assign n46177 = ~i_nEMPTY & ~n46176;
  assign n46178 = ~n46158 & ~n46177;
  assign n46179 = ~controllable_BtoS_ACK0 & ~n46178;
  assign n46180 = ~n46142 & ~n46179;
  assign n46181 = n4465 & ~n46180;
  assign n46182 = ~n45549 & ~n46181;
  assign n46183 = ~i_StoB_REQ10 & ~n46182;
  assign n46184 = ~n46105 & ~n46183;
  assign n46185 = controllable_BtoS_ACK10 & ~n46184;
  assign n46186 = ~n28596 & ~n45559;
  assign n46187 = ~controllable_DEQ & ~n46186;
  assign n46188 = ~n28139 & ~n46187;
  assign n46189 = i_FULL & ~n46188;
  assign n46190 = ~controllable_BtoR_REQ0 & ~n45568;
  assign n46191 = ~controllable_BtoR_REQ0 & ~n46190;
  assign n46192 = ~i_RtoB_ACK0 & ~n46191;
  assign n46193 = ~n45559 & ~n46192;
  assign n46194 = ~controllable_DEQ & ~n46193;
  assign n46195 = ~n28139 & ~n46194;
  assign n46196 = ~i_FULL & ~n46195;
  assign n46197 = ~n46189 & ~n46196;
  assign n46198 = i_nEMPTY & ~n46197;
  assign n46199 = ~n28612 & ~n45585;
  assign n46200 = ~controllable_DEQ & ~n46199;
  assign n46201 = ~n28153 & ~n46200;
  assign n46202 = i_FULL & ~n46201;
  assign n46203 = ~n37491 & ~n39107;
  assign n46204 = controllable_BtoR_REQ1 & ~n46203;
  assign n46205 = ~n45599 & ~n46204;
  assign n46206 = ~controllable_BtoR_REQ0 & ~n46205;
  assign n46207 = ~controllable_BtoR_REQ0 & ~n46206;
  assign n46208 = ~i_RtoB_ACK0 & ~n46207;
  assign n46209 = ~n45585 & ~n46208;
  assign n46210 = ~controllable_DEQ & ~n46209;
  assign n46211 = ~n28163 & ~n46210;
  assign n46212 = ~i_FULL & ~n46211;
  assign n46213 = ~n46202 & ~n46212;
  assign n46214 = ~i_nEMPTY & ~n46213;
  assign n46215 = ~n46198 & ~n46214;
  assign n46216 = controllable_BtoS_ACK0 & ~n46215;
  assign n46217 = ~n28071 & ~n45617;
  assign n46218 = ~controllable_DEQ & ~n46217;
  assign n46219 = ~n28200 & ~n46218;
  assign n46220 = i_FULL & ~n46219;
  assign n46221 = ~controllable_BtoR_REQ0 & ~n45626;
  assign n46222 = ~controllable_BtoR_REQ0 & ~n46221;
  assign n46223 = ~i_RtoB_ACK0 & ~n46222;
  assign n46224 = ~n45617 & ~n46223;
  assign n46225 = ~controllable_DEQ & ~n46224;
  assign n46226 = ~n28200 & ~n46225;
  assign n46227 = ~i_FULL & ~n46226;
  assign n46228 = ~n46220 & ~n46227;
  assign n46229 = i_nEMPTY & ~n46228;
  assign n46230 = ~n28087 & ~n45643;
  assign n46231 = ~controllable_DEQ & ~n46230;
  assign n46232 = ~n28214 & ~n46231;
  assign n46233 = i_FULL & ~n46232;
  assign n46234 = ~n37754 & ~n39180;
  assign n46235 = controllable_BtoR_REQ1 & ~n46234;
  assign n46236 = ~n45657 & ~n46235;
  assign n46237 = ~controllable_BtoR_REQ0 & ~n46236;
  assign n46238 = ~controllable_BtoR_REQ0 & ~n46237;
  assign n46239 = ~i_RtoB_ACK0 & ~n46238;
  assign n46240 = ~n45643 & ~n46239;
  assign n46241 = ~controllable_DEQ & ~n46240;
  assign n46242 = ~n28224 & ~n46241;
  assign n46243 = ~i_FULL & ~n46242;
  assign n46244 = ~n46233 & ~n46243;
  assign n46245 = ~i_nEMPTY & ~n46244;
  assign n46246 = ~n46229 & ~n46245;
  assign n46247 = ~controllable_BtoS_ACK0 & ~n46246;
  assign n46248 = ~n46216 & ~n46247;
  assign n46249 = n4465 & ~n46248;
  assign n46250 = ~n45679 & ~n46249;
  assign n46251 = i_StoB_REQ10 & ~n46250;
  assign n46252 = ~n46183 & ~n46251;
  assign n46253 = ~controllable_BtoS_ACK10 & ~n46252;
  assign n46254 = ~n46185 & ~n46253;
  assign n46255 = n4464 & ~n46254;
  assign n46256 = ~n45745 & ~n46255;
  assign n46257 = n4463 & ~n46256;
  assign n46258 = ~n45999 & ~n46257;
  assign n46259 = n4462 & ~n46258;
  assign n46260 = ~n46031 & ~n46259;
  assign n46261 = ~n4461 & ~n46260;
  assign n46262 = ~n46033 & ~n46261;
  assign n46263 = ~n4459 & ~n46262;
  assign n46264 = ~controllable_BtoR_REQ1 & ~n45153;
  assign n46265 = ~controllable_BtoR_REQ0 & ~n46264;
  assign n46266 = ~n39895 & ~n46265;
  assign n46267 = i_RtoB_ACK0 & ~n46266;
  assign n46268 = i_RtoB_ACK1 & ~n37037;
  assign n46269 = ~n11156 & ~n46268;
  assign n46270 = ~controllable_BtoR_REQ1 & ~n46269;
  assign n46271 = ~controllable_BtoR_REQ1 & ~n46270;
  assign n46272 = controllable_BtoR_REQ0 & ~n46271;
  assign n46273 = ~controllable_BtoR_REQ1 & ~n45158;
  assign n46274 = ~controllable_BtoR_REQ0 & ~n46273;
  assign n46275 = ~n46272 & ~n46274;
  assign n46276 = ~i_RtoB_ACK0 & ~n46275;
  assign n46277 = ~n46267 & ~n46276;
  assign n46278 = ~controllable_DEQ & ~n46277;
  assign n46279 = ~n14755 & ~n46278;
  assign n46280 = i_FULL & ~n46279;
  assign n46281 = ~n36899 & ~n46268;
  assign n46282 = ~controllable_BtoR_REQ1 & ~n46281;
  assign n46283 = ~controllable_BtoR_REQ1 & ~n46282;
  assign n46284 = controllable_BtoR_REQ0 & ~n46283;
  assign n46285 = ~controllable_BtoR_REQ1 & ~n45169;
  assign n46286 = ~controllable_BtoR_REQ0 & ~n46285;
  assign n46287 = ~n46284 & ~n46286;
  assign n46288 = ~i_RtoB_ACK0 & ~n46287;
  assign n46289 = ~n46267 & ~n46288;
  assign n46290 = ~controllable_DEQ & ~n46289;
  assign n46291 = ~n14755 & ~n46290;
  assign n46292 = ~i_FULL & ~n46291;
  assign n46293 = ~n46280 & ~n46292;
  assign n46294 = i_nEMPTY & ~n46293;
  assign n46295 = ~controllable_BtoR_REQ1 & ~n45185;
  assign n46296 = ~controllable_BtoR_REQ0 & ~n46295;
  assign n46297 = ~n39905 & ~n46296;
  assign n46298 = i_RtoB_ACK0 & ~n46297;
  assign n46299 = i_RtoB_ACK1 & ~n45181;
  assign n46300 = ~n12214 & ~n46299;
  assign n46301 = ~controllable_BtoR_REQ1 & ~n46300;
  assign n46302 = ~controllable_BtoR_REQ1 & ~n46301;
  assign n46303 = controllable_BtoR_REQ0 & ~n46302;
  assign n46304 = ~controllable_BtoR_REQ1 & ~n45190;
  assign n46305 = ~controllable_BtoR_REQ0 & ~n46304;
  assign n46306 = ~n46303 & ~n46305;
  assign n46307 = ~i_RtoB_ACK0 & ~n46306;
  assign n46308 = ~n46298 & ~n46307;
  assign n46309 = ~controllable_DEQ & ~n46308;
  assign n46310 = ~n14780 & ~n46309;
  assign n46311 = i_FULL & ~n46310;
  assign n46312 = ~n37040 & ~n46299;
  assign n46313 = ~controllable_BtoR_REQ1 & ~n46312;
  assign n46314 = ~controllable_BtoR_REQ1 & ~n46313;
  assign n46315 = controllable_BtoR_REQ0 & ~n46314;
  assign n46316 = ~controllable_BtoR_REQ1 & ~n45201;
  assign n46317 = ~controllable_BtoR_REQ0 & ~n46316;
  assign n46318 = ~n46315 & ~n46317;
  assign n46319 = ~i_RtoB_ACK0 & ~n46318;
  assign n46320 = ~n46298 & ~n46319;
  assign n46321 = ~controllable_DEQ & ~n46320;
  assign n46322 = ~n14798 & ~n46321;
  assign n46323 = ~i_FULL & ~n46322;
  assign n46324 = ~n46311 & ~n46323;
  assign n46325 = ~i_nEMPTY & ~n46324;
  assign n46326 = ~n46294 & ~n46325;
  assign n46327 = controllable_BtoS_ACK0 & ~n46326;
  assign n46328 = ~controllable_BtoR_REQ1 & ~n45217;
  assign n46329 = ~controllable_BtoR_REQ0 & ~n46328;
  assign n46330 = ~n39923 & ~n46329;
  assign n46331 = i_RtoB_ACK0 & ~n46330;
  assign n46332 = i_RtoB_ACK1 & ~n37123;
  assign n46333 = ~n5349 & ~n46332;
  assign n46334 = ~controllable_BtoR_REQ1 & ~n46333;
  assign n46335 = ~controllable_BtoR_REQ1 & ~n46334;
  assign n46336 = controllable_BtoR_REQ0 & ~n46335;
  assign n46337 = ~controllable_BtoR_REQ1 & ~n45222;
  assign n46338 = ~controllable_BtoR_REQ0 & ~n46337;
  assign n46339 = ~n46336 & ~n46338;
  assign n46340 = ~i_RtoB_ACK0 & ~n46339;
  assign n46341 = ~n46331 & ~n46340;
  assign n46342 = ~controllable_DEQ & ~n46341;
  assign n46343 = ~n28757 & ~n46342;
  assign n46344 = i_FULL & ~n46343;
  assign n46345 = ~n37080 & ~n46332;
  assign n46346 = ~controllable_BtoR_REQ1 & ~n46345;
  assign n46347 = ~controllable_BtoR_REQ1 & ~n46346;
  assign n46348 = controllable_BtoR_REQ0 & ~n46347;
  assign n46349 = ~controllable_BtoR_REQ1 & ~n45233;
  assign n46350 = ~controllable_BtoR_REQ0 & ~n46349;
  assign n46351 = ~n46348 & ~n46350;
  assign n46352 = ~i_RtoB_ACK0 & ~n46351;
  assign n46353 = ~n46331 & ~n46352;
  assign n46354 = ~controllable_DEQ & ~n46353;
  assign n46355 = ~n28757 & ~n46354;
  assign n46356 = ~i_FULL & ~n46355;
  assign n46357 = ~n46344 & ~n46356;
  assign n46358 = i_nEMPTY & ~n46357;
  assign n46359 = ~controllable_BtoR_REQ1 & ~n45249;
  assign n46360 = ~controllable_BtoR_REQ0 & ~n46359;
  assign n46361 = ~n39933 & ~n46360;
  assign n46362 = i_RtoB_ACK0 & ~n46361;
  assign n46363 = i_RtoB_ACK1 & ~n45245;
  assign n46364 = ~n9026 & ~n46363;
  assign n46365 = ~controllable_BtoR_REQ1 & ~n46364;
  assign n46366 = ~controllable_BtoR_REQ1 & ~n46365;
  assign n46367 = controllable_BtoR_REQ0 & ~n46366;
  assign n46368 = ~controllable_BtoR_REQ1 & ~n45254;
  assign n46369 = ~controllable_BtoR_REQ0 & ~n46368;
  assign n46370 = ~n46367 & ~n46369;
  assign n46371 = ~i_RtoB_ACK0 & ~n46370;
  assign n46372 = ~n46362 & ~n46371;
  assign n46373 = ~controllable_DEQ & ~n46372;
  assign n46374 = ~n28773 & ~n46373;
  assign n46375 = i_FULL & ~n46374;
  assign n46376 = ~n37126 & ~n46363;
  assign n46377 = ~controllable_BtoR_REQ1 & ~n46376;
  assign n46378 = ~controllable_BtoR_REQ1 & ~n46377;
  assign n46379 = controllable_BtoR_REQ0 & ~n46378;
  assign n46380 = ~controllable_BtoR_REQ1 & ~n45265;
  assign n46381 = ~controllable_BtoR_REQ0 & ~n46380;
  assign n46382 = ~n46379 & ~n46381;
  assign n46383 = ~i_RtoB_ACK0 & ~n46382;
  assign n46384 = ~n46362 & ~n46383;
  assign n46385 = ~controllable_DEQ & ~n46384;
  assign n46386 = ~n28787 & ~n46385;
  assign n46387 = ~i_FULL & ~n46386;
  assign n46388 = ~n46375 & ~n46387;
  assign n46389 = ~i_nEMPTY & ~n46388;
  assign n46390 = ~n46358 & ~n46389;
  assign n46391 = ~controllable_BtoS_ACK0 & ~n46390;
  assign n46392 = ~n46327 & ~n46391;
  assign n46393 = n4465 & ~n46392;
  assign n46394 = ~n28757 & ~n28815;
  assign n46395 = i_FULL & ~n46394;
  assign n46396 = ~n28827 & ~n46395;
  assign n46397 = i_nEMPTY & ~n46396;
  assign n46398 = ~n28847 & ~n46397;
  assign n46399 = ~controllable_BtoS_ACK0 & ~n46398;
  assign n46400 = ~n14811 & ~n46399;
  assign n46401 = ~n4465 & ~n46400;
  assign n46402 = ~n46393 & ~n46401;
  assign n46403 = i_StoB_REQ10 & ~n46402;
  assign n46404 = ~n37915 & ~n38940;
  assign n46405 = ~controllable_BtoR_REQ1 & ~n46404;
  assign n46406 = ~controllable_BtoR_REQ1 & ~n46405;
  assign n46407 = controllable_BtoR_REQ0 & ~n46406;
  assign n46408 = ~controllable_BtoR_REQ1 & ~n45380;
  assign n46409 = ~controllable_BtoR_REQ0 & ~n46408;
  assign n46410 = ~n46407 & ~n46409;
  assign n46411 = i_RtoB_ACK0 & ~n46410;
  assign n46412 = i_RtoB_ACK1 & ~n37661;
  assign n46413 = ~n12387 & ~n46412;
  assign n46414 = ~controllable_BtoR_REQ1 & ~n46413;
  assign n46415 = ~controllable_BtoR_REQ1 & ~n46414;
  assign n46416 = controllable_BtoR_REQ0 & ~n46415;
  assign n46417 = ~controllable_BtoR_REQ1 & ~n45388;
  assign n46418 = ~controllable_BtoR_REQ0 & ~n46417;
  assign n46419 = ~n46416 & ~n46418;
  assign n46420 = ~i_RtoB_ACK0 & ~n46419;
  assign n46421 = ~n46411 & ~n46420;
  assign n46422 = ~controllable_DEQ & ~n46421;
  assign n46423 = ~n17626 & ~n46422;
  assign n46424 = i_FULL & ~n46423;
  assign n46425 = ~n37491 & ~n46412;
  assign n46426 = ~controllable_BtoR_REQ1 & ~n46425;
  assign n46427 = ~controllable_BtoR_REQ1 & ~n46426;
  assign n46428 = controllable_BtoR_REQ0 & ~n46427;
  assign n46429 = ~controllable_BtoR_REQ1 & ~n45399;
  assign n46430 = ~controllable_BtoR_REQ0 & ~n46429;
  assign n46431 = ~n46428 & ~n46430;
  assign n46432 = ~i_RtoB_ACK0 & ~n46431;
  assign n46433 = ~n46411 & ~n46432;
  assign n46434 = ~controllable_DEQ & ~n46433;
  assign n46435 = ~n17626 & ~n46434;
  assign n46436 = ~i_FULL & ~n46435;
  assign n46437 = ~n46424 & ~n46436;
  assign n46438 = i_nEMPTY & ~n46437;
  assign n46439 = ~n37948 & ~n45412;
  assign n46440 = ~controllable_BtoR_REQ1 & ~n46439;
  assign n46441 = ~controllable_BtoR_REQ1 & ~n46440;
  assign n46442 = controllable_BtoR_REQ0 & ~n46441;
  assign n46443 = ~controllable_BtoR_REQ1 & ~n45420;
  assign n46444 = ~controllable_BtoR_REQ0 & ~n46443;
  assign n46445 = ~n46442 & ~n46444;
  assign n46446 = i_RtoB_ACK0 & ~n46445;
  assign n46447 = i_RtoB_ACK1 & ~n45414;
  assign n46448 = ~n12431 & ~n46447;
  assign n46449 = ~controllable_BtoR_REQ1 & ~n46448;
  assign n46450 = ~controllable_BtoR_REQ1 & ~n46449;
  assign n46451 = controllable_BtoR_REQ0 & ~n46450;
  assign n46452 = ~controllable_BtoR_REQ1 & ~n45428;
  assign n46453 = ~controllable_BtoR_REQ0 & ~n46452;
  assign n46454 = ~n46451 & ~n46453;
  assign n46455 = ~i_RtoB_ACK0 & ~n46454;
  assign n46456 = ~n46446 & ~n46455;
  assign n46457 = ~controllable_DEQ & ~n46456;
  assign n46458 = ~n17651 & ~n46457;
  assign n46459 = i_FULL & ~n46458;
  assign n46460 = ~i_RtoB_ACK1 & ~n45437;
  assign n46461 = ~n45412 & ~n46460;
  assign n46462 = ~controllable_BtoR_REQ1 & ~n46461;
  assign n46463 = ~controllable_BtoR_REQ1 & ~n46462;
  assign n46464 = controllable_BtoR_REQ0 & ~n46463;
  assign n46465 = ~n46444 & ~n46464;
  assign n46466 = i_RtoB_ACK0 & ~n46465;
  assign n46467 = ~n37664 & ~n46447;
  assign n46468 = ~controllable_BtoR_REQ1 & ~n46467;
  assign n46469 = ~controllable_BtoR_REQ1 & ~n46468;
  assign n46470 = controllable_BtoR_REQ0 & ~n46469;
  assign n46471 = ~controllable_BtoR_REQ1 & ~n45442;
  assign n46472 = ~controllable_BtoR_REQ0 & ~n46471;
  assign n46473 = ~n46470 & ~n46472;
  assign n46474 = ~i_RtoB_ACK0 & ~n46473;
  assign n46475 = ~n46466 & ~n46474;
  assign n46476 = ~controllable_DEQ & ~n46475;
  assign n46477 = ~n17673 & ~n46476;
  assign n46478 = ~i_FULL & ~n46477;
  assign n46479 = ~n46459 & ~n46478;
  assign n46480 = ~i_nEMPTY & ~n46479;
  assign n46481 = ~n46438 & ~n46480;
  assign n46482 = controllable_BtoS_ACK0 & ~n46481;
  assign n46483 = ~n37999 & ~n39035;
  assign n46484 = ~controllable_BtoR_REQ1 & ~n46483;
  assign n46485 = ~controllable_BtoR_REQ1 & ~n46484;
  assign n46486 = controllable_BtoR_REQ0 & ~n46485;
  assign n46487 = ~controllable_BtoR_REQ1 & ~n45465;
  assign n46488 = ~controllable_BtoR_REQ0 & ~n46487;
  assign n46489 = ~n46486 & ~n46488;
  assign n46490 = i_RtoB_ACK0 & ~n46489;
  assign n46491 = i_RtoB_ACK1 & ~n37823;
  assign n46492 = ~n9913 & ~n46491;
  assign n46493 = ~controllable_BtoR_REQ1 & ~n46492;
  assign n46494 = ~controllable_BtoR_REQ1 & ~n46493;
  assign n46495 = controllable_BtoR_REQ0 & ~n46494;
  assign n46496 = ~controllable_BtoR_REQ1 & ~n45473;
  assign n46497 = ~controllable_BtoR_REQ0 & ~n46496;
  assign n46498 = ~n46495 & ~n46497;
  assign n46499 = ~i_RtoB_ACK0 & ~n46498;
  assign n46500 = ~n46490 & ~n46499;
  assign n46501 = ~controllable_DEQ & ~n46500;
  assign n46502 = ~n17705 & ~n46501;
  assign n46503 = i_FULL & ~n46502;
  assign n46504 = ~n37754 & ~n46491;
  assign n46505 = ~controllable_BtoR_REQ1 & ~n46504;
  assign n46506 = ~controllable_BtoR_REQ1 & ~n46505;
  assign n46507 = controllable_BtoR_REQ0 & ~n46506;
  assign n46508 = ~controllable_BtoR_REQ1 & ~n45484;
  assign n46509 = ~controllable_BtoR_REQ0 & ~n46508;
  assign n46510 = ~n46507 & ~n46509;
  assign n46511 = ~i_RtoB_ACK0 & ~n46510;
  assign n46512 = ~n46490 & ~n46511;
  assign n46513 = ~controllable_DEQ & ~n46512;
  assign n46514 = ~n17705 & ~n46513;
  assign n46515 = ~i_FULL & ~n46514;
  assign n46516 = ~n46503 & ~n46515;
  assign n46517 = i_nEMPTY & ~n46516;
  assign n46518 = ~n38032 & ~n45497;
  assign n46519 = ~controllable_BtoR_REQ1 & ~n46518;
  assign n46520 = ~controllable_BtoR_REQ1 & ~n46519;
  assign n46521 = controllable_BtoR_REQ0 & ~n46520;
  assign n46522 = ~controllable_BtoR_REQ1 & ~n45505;
  assign n46523 = ~controllable_BtoR_REQ0 & ~n46522;
  assign n46524 = ~n46521 & ~n46523;
  assign n46525 = i_RtoB_ACK0 & ~n46524;
  assign n46526 = i_RtoB_ACK1 & ~n45499;
  assign n46527 = ~n9961 & ~n46526;
  assign n46528 = ~controllable_BtoR_REQ1 & ~n46527;
  assign n46529 = ~controllable_BtoR_REQ1 & ~n46528;
  assign n46530 = controllable_BtoR_REQ0 & ~n46529;
  assign n46531 = ~controllable_BtoR_REQ1 & ~n45513;
  assign n46532 = ~controllable_BtoR_REQ0 & ~n46531;
  assign n46533 = ~n46530 & ~n46532;
  assign n46534 = ~i_RtoB_ACK0 & ~n46533;
  assign n46535 = ~n46525 & ~n46534;
  assign n46536 = ~controllable_DEQ & ~n46535;
  assign n46537 = ~n17741 & ~n46536;
  assign n46538 = i_FULL & ~n46537;
  assign n46539 = ~i_RtoB_ACK1 & ~n45522;
  assign n46540 = ~n45497 & ~n46539;
  assign n46541 = ~controllable_BtoR_REQ1 & ~n46540;
  assign n46542 = ~controllable_BtoR_REQ1 & ~n46541;
  assign n46543 = controllable_BtoR_REQ0 & ~n46542;
  assign n46544 = ~n46523 & ~n46543;
  assign n46545 = i_RtoB_ACK0 & ~n46544;
  assign n46546 = ~n37826 & ~n46526;
  assign n46547 = ~controllable_BtoR_REQ1 & ~n46546;
  assign n46548 = ~controllable_BtoR_REQ1 & ~n46547;
  assign n46549 = controllable_BtoR_REQ0 & ~n46548;
  assign n46550 = ~controllable_BtoR_REQ1 & ~n45527;
  assign n46551 = ~controllable_BtoR_REQ0 & ~n46550;
  assign n46552 = ~n46549 & ~n46551;
  assign n46553 = ~i_RtoB_ACK0 & ~n46552;
  assign n46554 = ~n46545 & ~n46553;
  assign n46555 = ~controllable_DEQ & ~n46554;
  assign n46556 = ~n17774 & ~n46555;
  assign n46557 = ~i_FULL & ~n46556;
  assign n46558 = ~n46538 & ~n46557;
  assign n46559 = ~i_nEMPTY & ~n46558;
  assign n46560 = ~n46517 & ~n46559;
  assign n46561 = ~controllable_BtoS_ACK0 & ~n46560;
  assign n46562 = ~n46482 & ~n46561;
  assign n46563 = n4465 & ~n46562;
  assign n46564 = ~n17705 & ~n28975;
  assign n46565 = i_FULL & ~n46564;
  assign n46566 = ~n28987 & ~n46565;
  assign n46567 = i_nEMPTY & ~n46566;
  assign n46568 = ~n29007 & ~n46567;
  assign n46569 = ~controllable_BtoS_ACK0 & ~n46568;
  assign n46570 = ~n17685 & ~n46569;
  assign n46571 = ~n4465 & ~n46570;
  assign n46572 = ~n46563 & ~n46571;
  assign n46573 = ~i_StoB_REQ10 & ~n46572;
  assign n46574 = ~n46403 & ~n46573;
  assign n46575 = controllable_BtoS_ACK10 & ~n46574;
  assign n46576 = ~controllable_BtoR_REQ1 & ~n45554;
  assign n46577 = ~controllable_BtoR_REQ1 & ~n46576;
  assign n46578 = controllable_BtoR_REQ0 & ~n46577;
  assign n46579 = ~n17628 & ~n46578;
  assign n46580 = i_RtoB_ACK0 & ~n46579;
  assign n46581 = controllable_BtoR_REQ0 & ~n40936;
  assign n46582 = ~n20379 & ~n46581;
  assign n46583 = ~i_RtoB_ACK0 & ~n46582;
  assign n46584 = ~n46580 & ~n46583;
  assign n46585 = ~controllable_DEQ & ~n46584;
  assign n46586 = ~n29030 & ~n46585;
  assign n46587 = i_FULL & ~n46586;
  assign n46588 = controllable_BtoR_REQ0 & ~n40952;
  assign n46589 = ~controllable_BtoR_REQ1 & ~n45569;
  assign n46590 = ~controllable_BtoR_REQ0 & ~n46589;
  assign n46591 = ~n46588 & ~n46590;
  assign n46592 = ~i_RtoB_ACK0 & ~n46591;
  assign n46593 = ~n46580 & ~n46592;
  assign n46594 = ~controllable_DEQ & ~n46593;
  assign n46595 = ~n29030 & ~n46594;
  assign n46596 = ~i_FULL & ~n46595;
  assign n46597 = ~n46587 & ~n46596;
  assign n46598 = i_nEMPTY & ~n46597;
  assign n46599 = ~controllable_BtoR_REQ1 & ~n45580;
  assign n46600 = ~controllable_BtoR_REQ1 & ~n46599;
  assign n46601 = controllable_BtoR_REQ0 & ~n46600;
  assign n46602 = ~n17613 & ~n46601;
  assign n46603 = i_RtoB_ACK0 & ~n46602;
  assign n46604 = controllable_BtoR_REQ0 & ~n40970;
  assign n46605 = ~n20413 & ~n46604;
  assign n46606 = ~i_RtoB_ACK0 & ~n46605;
  assign n46607 = ~n46603 & ~n46606;
  assign n46608 = ~controllable_DEQ & ~n46607;
  assign n46609 = ~n29040 & ~n46608;
  assign n46610 = i_FULL & ~n46609;
  assign n46611 = ~i_RtoB_ACK1 & ~n45594;
  assign n46612 = ~n14073 & ~n46611;
  assign n46613 = ~controllable_BtoR_REQ1 & ~n46612;
  assign n46614 = ~controllable_BtoR_REQ1 & ~n46613;
  assign n46615 = controllable_BtoR_REQ0 & ~n46614;
  assign n46616 = ~n17613 & ~n46615;
  assign n46617 = i_RtoB_ACK0 & ~n46616;
  assign n46618 = controllable_BtoR_REQ0 & ~n40985;
  assign n46619 = ~controllable_BtoR_REQ1 & ~n45599;
  assign n46620 = ~controllable_BtoR_REQ0 & ~n46619;
  assign n46621 = ~n46618 & ~n46620;
  assign n46622 = ~i_RtoB_ACK0 & ~n46621;
  assign n46623 = ~n46617 & ~n46622;
  assign n46624 = ~controllable_DEQ & ~n46623;
  assign n46625 = ~n29050 & ~n46624;
  assign n46626 = ~i_FULL & ~n46625;
  assign n46627 = ~n46610 & ~n46626;
  assign n46628 = ~i_nEMPTY & ~n46627;
  assign n46629 = ~n46598 & ~n46628;
  assign n46630 = controllable_BtoS_ACK0 & ~n46629;
  assign n46631 = ~controllable_BtoR_REQ1 & ~n45612;
  assign n46632 = ~controllable_BtoR_REQ1 & ~n46631;
  assign n46633 = controllable_BtoR_REQ0 & ~n46632;
  assign n46634 = ~n17711 & ~n46633;
  assign n46635 = i_RtoB_ACK0 & ~n46634;
  assign n46636 = controllable_BtoR_REQ0 & ~n41007;
  assign n46637 = ~n19323 & ~n46636;
  assign n46638 = ~i_RtoB_ACK0 & ~n46637;
  assign n46639 = ~n46635 & ~n46638;
  assign n46640 = ~controllable_DEQ & ~n46639;
  assign n46641 = ~n29072 & ~n46640;
  assign n46642 = i_FULL & ~n46641;
  assign n46643 = controllable_BtoR_REQ0 & ~n41023;
  assign n46644 = ~controllable_BtoR_REQ1 & ~n45627;
  assign n46645 = ~controllable_BtoR_REQ0 & ~n46644;
  assign n46646 = ~n46643 & ~n46645;
  assign n46647 = ~i_RtoB_ACK0 & ~n46646;
  assign n46648 = ~n46635 & ~n46647;
  assign n46649 = ~controllable_DEQ & ~n46648;
  assign n46650 = ~n29072 & ~n46649;
  assign n46651 = ~i_FULL & ~n46650;
  assign n46652 = ~n46642 & ~n46651;
  assign n46653 = i_nEMPTY & ~n46652;
  assign n46654 = ~controllable_BtoR_REQ1 & ~n45638;
  assign n46655 = ~controllable_BtoR_REQ1 & ~n46654;
  assign n46656 = controllable_BtoR_REQ0 & ~n46655;
  assign n46657 = ~n17692 & ~n46656;
  assign n46658 = i_RtoB_ACK0 & ~n46657;
  assign n46659 = controllable_BtoR_REQ0 & ~n41041;
  assign n46660 = ~n19353 & ~n46659;
  assign n46661 = ~i_RtoB_ACK0 & ~n46660;
  assign n46662 = ~n46658 & ~n46661;
  assign n46663 = ~controllable_DEQ & ~n46662;
  assign n46664 = ~n29082 & ~n46663;
  assign n46665 = i_FULL & ~n46664;
  assign n46666 = ~i_RtoB_ACK1 & ~n45652;
  assign n46667 = ~n14116 & ~n46666;
  assign n46668 = ~controllable_BtoR_REQ1 & ~n46667;
  assign n46669 = ~controllable_BtoR_REQ1 & ~n46668;
  assign n46670 = controllable_BtoR_REQ0 & ~n46669;
  assign n46671 = ~n17692 & ~n46670;
  assign n46672 = i_RtoB_ACK0 & ~n46671;
  assign n46673 = controllable_BtoR_REQ0 & ~n41056;
  assign n46674 = ~controllable_BtoR_REQ1 & ~n45657;
  assign n46675 = ~controllable_BtoR_REQ0 & ~n46674;
  assign n46676 = ~n46673 & ~n46675;
  assign n46677 = ~i_RtoB_ACK0 & ~n46676;
  assign n46678 = ~n46672 & ~n46677;
  assign n46679 = ~controllable_DEQ & ~n46678;
  assign n46680 = ~n29092 & ~n46679;
  assign n46681 = ~i_FULL & ~n46680;
  assign n46682 = ~n46665 & ~n46681;
  assign n46683 = ~i_nEMPTY & ~n46682;
  assign n46684 = ~n46653 & ~n46683;
  assign n46685 = ~controllable_BtoS_ACK0 & ~n46684;
  assign n46686 = ~n46630 & ~n46685;
  assign n46687 = n4465 & ~n46686;
  assign n46688 = ~n29072 & ~n29124;
  assign n46689 = i_FULL & ~n46688;
  assign n46690 = ~n29131 & ~n46689;
  assign n46691 = i_nEMPTY & ~n46690;
  assign n46692 = ~n29143 & ~n46691;
  assign n46693 = ~controllable_BtoS_ACK0 & ~n46692;
  assign n46694 = ~n29118 & ~n46693;
  assign n46695 = ~n4465 & ~n46694;
  assign n46696 = ~n46687 & ~n46695;
  assign n46697 = i_StoB_REQ10 & ~n46696;
  assign n46698 = ~n46573 & ~n46697;
  assign n46699 = ~controllable_BtoS_ACK10 & ~n46698;
  assign n46700 = ~n46575 & ~n46699;
  assign n46701 = n4464 & ~n46700;
  assign n46702 = ~n14755 & ~n29169;
  assign n46703 = i_FULL & ~n46702;
  assign n46704 = ~n29181 & ~n46703;
  assign n46705 = i_nEMPTY & ~n46704;
  assign n46706 = ~n29201 & ~n46705;
  assign n46707 = controllable_BtoS_ACK0 & ~n46706;
  assign n46708 = ~n28757 & ~n29219;
  assign n46709 = i_FULL & ~n46708;
  assign n46710 = ~n29231 & ~n46709;
  assign n46711 = i_nEMPTY & ~n46710;
  assign n46712 = ~n29251 & ~n46711;
  assign n46713 = ~controllable_BtoS_ACK0 & ~n46712;
  assign n46714 = ~n46707 & ~n46713;
  assign n46715 = n4465 & ~n46714;
  assign n46716 = ~n14811 & ~n46713;
  assign n46717 = ~n4465 & ~n46716;
  assign n46718 = ~n46715 & ~n46717;
  assign n46719 = i_StoB_REQ10 & ~n46718;
  assign n46720 = ~n17626 & ~n29275;
  assign n46721 = i_FULL & ~n46720;
  assign n46722 = ~n29287 & ~n46721;
  assign n46723 = i_nEMPTY & ~n46722;
  assign n46724 = ~n29307 & ~n46723;
  assign n46725 = controllable_BtoS_ACK0 & ~n46724;
  assign n46726 = ~n17705 & ~n29325;
  assign n46727 = i_FULL & ~n46726;
  assign n46728 = ~n29337 & ~n46727;
  assign n46729 = i_nEMPTY & ~n46728;
  assign n46730 = ~n29357 & ~n46729;
  assign n46731 = ~controllable_BtoS_ACK0 & ~n46730;
  assign n46732 = ~n46725 & ~n46731;
  assign n46733 = n4465 & ~n46732;
  assign n46734 = ~n17685 & ~n46731;
  assign n46735 = ~n4465 & ~n46734;
  assign n46736 = ~n46733 & ~n46735;
  assign n46737 = ~i_StoB_REQ10 & ~n46736;
  assign n46738 = ~n46719 & ~n46737;
  assign n46739 = controllable_BtoS_ACK10 & ~n46738;
  assign n46740 = ~n29030 & ~n29373;
  assign n46741 = i_FULL & ~n46740;
  assign n46742 = ~n29380 & ~n46741;
  assign n46743 = i_nEMPTY & ~n46742;
  assign n46744 = ~n29392 & ~n46743;
  assign n46745 = controllable_BtoS_ACK0 & ~n46744;
  assign n46746 = ~n29072 & ~n29400;
  assign n46747 = i_FULL & ~n46746;
  assign n46748 = ~n29407 & ~n46747;
  assign n46749 = i_nEMPTY & ~n46748;
  assign n46750 = ~n29419 & ~n46749;
  assign n46751 = ~controllable_BtoS_ACK0 & ~n46750;
  assign n46752 = ~n46745 & ~n46751;
  assign n46753 = n4465 & ~n46752;
  assign n46754 = ~n29118 & ~n46751;
  assign n46755 = ~n4465 & ~n46754;
  assign n46756 = ~n46753 & ~n46755;
  assign n46757 = i_StoB_REQ10 & ~n46756;
  assign n46758 = ~n46737 & ~n46757;
  assign n46759 = ~controllable_BtoS_ACK10 & ~n46758;
  assign n46760 = ~n46739 & ~n46759;
  assign n46761 = ~n4464 & ~n46760;
  assign n46762 = ~n46701 & ~n46761;
  assign n46763 = n4463 & ~n46762;
  assign n46764 = ~n18434 & ~n46265;
  assign n46765 = i_RtoB_ACK0 & ~n46764;
  assign n46766 = ~n46276 & ~n46765;
  assign n46767 = ~controllable_DEQ & ~n46766;
  assign n46768 = ~n14755 & ~n46767;
  assign n46769 = i_FULL & ~n46768;
  assign n46770 = ~n46288 & ~n46765;
  assign n46771 = ~controllable_DEQ & ~n46770;
  assign n46772 = ~n14755 & ~n46771;
  assign n46773 = ~i_FULL & ~n46772;
  assign n46774 = ~n46769 & ~n46773;
  assign n46775 = i_nEMPTY & ~n46774;
  assign n46776 = ~n18428 & ~n46296;
  assign n46777 = i_RtoB_ACK0 & ~n46776;
  assign n46778 = ~n46307 & ~n46777;
  assign n46779 = ~controllable_DEQ & ~n46778;
  assign n46780 = ~n14780 & ~n46779;
  assign n46781 = i_FULL & ~n46780;
  assign n46782 = ~n46319 & ~n46777;
  assign n46783 = ~controllable_DEQ & ~n46782;
  assign n46784 = ~n14798 & ~n46783;
  assign n46785 = ~i_FULL & ~n46784;
  assign n46786 = ~n46781 & ~n46785;
  assign n46787 = ~i_nEMPTY & ~n46786;
  assign n46788 = ~n46775 & ~n46787;
  assign n46789 = controllable_BtoS_ACK0 & ~n46788;
  assign n46790 = ~n18462 & ~n46329;
  assign n46791 = i_RtoB_ACK0 & ~n46790;
  assign n46792 = ~n46340 & ~n46791;
  assign n46793 = ~controllable_DEQ & ~n46792;
  assign n46794 = ~n28757 & ~n46793;
  assign n46795 = i_FULL & ~n46794;
  assign n46796 = ~n46352 & ~n46791;
  assign n46797 = ~controllable_DEQ & ~n46796;
  assign n46798 = ~n28757 & ~n46797;
  assign n46799 = ~i_FULL & ~n46798;
  assign n46800 = ~n46795 & ~n46799;
  assign n46801 = i_nEMPTY & ~n46800;
  assign n46802 = ~n18456 & ~n46360;
  assign n46803 = i_RtoB_ACK0 & ~n46802;
  assign n46804 = ~n46371 & ~n46803;
  assign n46805 = ~controllable_DEQ & ~n46804;
  assign n46806 = ~n28773 & ~n46805;
  assign n46807 = i_FULL & ~n46806;
  assign n46808 = ~n46383 & ~n46803;
  assign n46809 = ~controllable_DEQ & ~n46808;
  assign n46810 = ~n28787 & ~n46809;
  assign n46811 = ~i_FULL & ~n46810;
  assign n46812 = ~n46807 & ~n46811;
  assign n46813 = ~i_nEMPTY & ~n46812;
  assign n46814 = ~n46801 & ~n46813;
  assign n46815 = ~controllable_BtoS_ACK0 & ~n46814;
  assign n46816 = ~n46789 & ~n46815;
  assign n46817 = n4465 & ~n46816;
  assign n46818 = ~n46401 & ~n46817;
  assign n46819 = i_StoB_REQ10 & ~n46818;
  assign n46820 = ~i_RtoB_ACK1 & ~n45379;
  assign n46821 = ~n38940 & ~n46820;
  assign n46822 = ~controllable_BtoR_REQ1 & ~n46821;
  assign n46823 = ~controllable_BtoR_REQ1 & ~n46822;
  assign n46824 = controllable_BtoR_REQ0 & ~n46823;
  assign n46825 = ~n46409 & ~n46824;
  assign n46826 = i_RtoB_ACK0 & ~n46825;
  assign n46827 = ~n46420 & ~n46826;
  assign n46828 = ~controllable_DEQ & ~n46827;
  assign n46829 = ~n17626 & ~n46828;
  assign n46830 = i_FULL & ~n46829;
  assign n46831 = ~n46432 & ~n46826;
  assign n46832 = ~controllable_DEQ & ~n46831;
  assign n46833 = ~n17626 & ~n46832;
  assign n46834 = ~i_FULL & ~n46833;
  assign n46835 = ~n46830 & ~n46834;
  assign n46836 = i_nEMPTY & ~n46835;
  assign n46837 = ~i_RtoB_ACK1 & ~n45419;
  assign n46838 = ~n45412 & ~n46837;
  assign n46839 = ~controllable_BtoR_REQ1 & ~n46838;
  assign n46840 = ~controllable_BtoR_REQ1 & ~n46839;
  assign n46841 = controllable_BtoR_REQ0 & ~n46840;
  assign n46842 = ~n46444 & ~n46841;
  assign n46843 = i_RtoB_ACK0 & ~n46842;
  assign n46844 = ~n46455 & ~n46843;
  assign n46845 = ~controllable_DEQ & ~n46844;
  assign n46846 = ~n17651 & ~n46845;
  assign n46847 = i_FULL & ~n46846;
  assign n46848 = ~i_RtoB_ACK1 & ~n45853;
  assign n46849 = ~n45412 & ~n46848;
  assign n46850 = ~controllable_BtoR_REQ1 & ~n46849;
  assign n46851 = ~controllable_BtoR_REQ1 & ~n46850;
  assign n46852 = controllable_BtoR_REQ0 & ~n46851;
  assign n46853 = ~n46444 & ~n46852;
  assign n46854 = i_RtoB_ACK0 & ~n46853;
  assign n46855 = ~n46474 & ~n46854;
  assign n46856 = ~controllable_DEQ & ~n46855;
  assign n46857 = ~n17673 & ~n46856;
  assign n46858 = ~i_FULL & ~n46857;
  assign n46859 = ~n46847 & ~n46858;
  assign n46860 = ~i_nEMPTY & ~n46859;
  assign n46861 = ~n46836 & ~n46860;
  assign n46862 = controllable_BtoS_ACK0 & ~n46861;
  assign n46863 = ~i_RtoB_ACK1 & ~n45464;
  assign n46864 = ~n39035 & ~n46863;
  assign n46865 = ~controllable_BtoR_REQ1 & ~n46864;
  assign n46866 = ~controllable_BtoR_REQ1 & ~n46865;
  assign n46867 = controllable_BtoR_REQ0 & ~n46866;
  assign n46868 = ~n46488 & ~n46867;
  assign n46869 = i_RtoB_ACK0 & ~n46868;
  assign n46870 = ~n46499 & ~n46869;
  assign n46871 = ~controllable_DEQ & ~n46870;
  assign n46872 = ~n17705 & ~n46871;
  assign n46873 = i_FULL & ~n46872;
  assign n46874 = ~n46511 & ~n46869;
  assign n46875 = ~controllable_DEQ & ~n46874;
  assign n46876 = ~n17705 & ~n46875;
  assign n46877 = ~i_FULL & ~n46876;
  assign n46878 = ~n46873 & ~n46877;
  assign n46879 = i_nEMPTY & ~n46878;
  assign n46880 = ~i_RtoB_ACK1 & ~n45504;
  assign n46881 = ~n45497 & ~n46880;
  assign n46882 = ~controllable_BtoR_REQ1 & ~n46881;
  assign n46883 = ~controllable_BtoR_REQ1 & ~n46882;
  assign n46884 = controllable_BtoR_REQ0 & ~n46883;
  assign n46885 = ~n46523 & ~n46884;
  assign n46886 = i_RtoB_ACK0 & ~n46885;
  assign n46887 = ~n46534 & ~n46886;
  assign n46888 = ~controllable_DEQ & ~n46887;
  assign n46889 = ~n17741 & ~n46888;
  assign n46890 = i_FULL & ~n46889;
  assign n46891 = ~i_RtoB_ACK1 & ~n45897;
  assign n46892 = ~n45497 & ~n46891;
  assign n46893 = ~controllable_BtoR_REQ1 & ~n46892;
  assign n46894 = ~controllable_BtoR_REQ1 & ~n46893;
  assign n46895 = controllable_BtoR_REQ0 & ~n46894;
  assign n46896 = ~n46523 & ~n46895;
  assign n46897 = i_RtoB_ACK0 & ~n46896;
  assign n46898 = ~n46553 & ~n46897;
  assign n46899 = ~controllable_DEQ & ~n46898;
  assign n46900 = ~n17774 & ~n46899;
  assign n46901 = ~i_FULL & ~n46900;
  assign n46902 = ~n46890 & ~n46901;
  assign n46903 = ~i_nEMPTY & ~n46902;
  assign n46904 = ~n46879 & ~n46903;
  assign n46905 = ~controllable_BtoS_ACK0 & ~n46904;
  assign n46906 = ~n46862 & ~n46905;
  assign n46907 = n4465 & ~n46906;
  assign n46908 = ~n46571 & ~n46907;
  assign n46909 = ~i_StoB_REQ10 & ~n46908;
  assign n46910 = ~n46819 & ~n46909;
  assign n46911 = controllable_BtoS_ACK10 & ~n46910;
  assign n46912 = ~n9813 & ~n14082;
  assign n46913 = ~controllable_BtoR_REQ1 & ~n46912;
  assign n46914 = ~controllable_BtoR_REQ1 & ~n46913;
  assign n46915 = controllable_BtoR_REQ0 & ~n46914;
  assign n46916 = ~n17628 & ~n46915;
  assign n46917 = i_RtoB_ACK0 & ~n46916;
  assign n46918 = ~n46583 & ~n46917;
  assign n46919 = ~controllable_DEQ & ~n46918;
  assign n46920 = ~n29030 & ~n46919;
  assign n46921 = i_FULL & ~n46920;
  assign n46922 = ~n46592 & ~n46917;
  assign n46923 = ~controllable_DEQ & ~n46922;
  assign n46924 = ~n29030 & ~n46923;
  assign n46925 = ~i_FULL & ~n46924;
  assign n46926 = ~n46921 & ~n46925;
  assign n46927 = i_nEMPTY & ~n46926;
  assign n46928 = ~n9836 & ~n14073;
  assign n46929 = ~controllable_BtoR_REQ1 & ~n46928;
  assign n46930 = ~controllable_BtoR_REQ1 & ~n46929;
  assign n46931 = controllable_BtoR_REQ0 & ~n46930;
  assign n46932 = ~n17613 & ~n46931;
  assign n46933 = i_RtoB_ACK0 & ~n46932;
  assign n46934 = ~n46606 & ~n46933;
  assign n46935 = ~controllable_DEQ & ~n46934;
  assign n46936 = ~n29040 & ~n46935;
  assign n46937 = i_FULL & ~n46936;
  assign n46938 = ~n14073 & ~n40128;
  assign n46939 = ~controllable_BtoR_REQ1 & ~n46938;
  assign n46940 = ~controllable_BtoR_REQ1 & ~n46939;
  assign n46941 = controllable_BtoR_REQ0 & ~n46940;
  assign n46942 = ~n17613 & ~n46941;
  assign n46943 = i_RtoB_ACK0 & ~n46942;
  assign n46944 = ~n46622 & ~n46943;
  assign n46945 = ~controllable_DEQ & ~n46944;
  assign n46946 = ~n29050 & ~n46945;
  assign n46947 = ~i_FULL & ~n46946;
  assign n46948 = ~n46937 & ~n46947;
  assign n46949 = ~i_nEMPTY & ~n46948;
  assign n46950 = ~n46927 & ~n46949;
  assign n46951 = controllable_BtoS_ACK0 & ~n46950;
  assign n46952 = ~n9904 & ~n14125;
  assign n46953 = ~controllable_BtoR_REQ1 & ~n46952;
  assign n46954 = ~controllable_BtoR_REQ1 & ~n46953;
  assign n46955 = controllable_BtoR_REQ0 & ~n46954;
  assign n46956 = ~n17711 & ~n46955;
  assign n46957 = i_RtoB_ACK0 & ~n46956;
  assign n46958 = ~n46638 & ~n46957;
  assign n46959 = ~controllable_DEQ & ~n46958;
  assign n46960 = ~n29072 & ~n46959;
  assign n46961 = i_FULL & ~n46960;
  assign n46962 = ~n46647 & ~n46957;
  assign n46963 = ~controllable_DEQ & ~n46962;
  assign n46964 = ~n29072 & ~n46963;
  assign n46965 = ~i_FULL & ~n46964;
  assign n46966 = ~n46961 & ~n46965;
  assign n46967 = i_nEMPTY & ~n46966;
  assign n46968 = ~n9871 & ~n14116;
  assign n46969 = ~controllable_BtoR_REQ1 & ~n46968;
  assign n46970 = ~controllable_BtoR_REQ1 & ~n46969;
  assign n46971 = controllable_BtoR_REQ0 & ~n46970;
  assign n46972 = ~n17692 & ~n46971;
  assign n46973 = i_RtoB_ACK0 & ~n46972;
  assign n46974 = ~n46661 & ~n46973;
  assign n46975 = ~controllable_DEQ & ~n46974;
  assign n46976 = ~n29082 & ~n46975;
  assign n46977 = i_FULL & ~n46976;
  assign n46978 = ~n14116 & ~n40189;
  assign n46979 = ~controllable_BtoR_REQ1 & ~n46978;
  assign n46980 = ~controllable_BtoR_REQ1 & ~n46979;
  assign n46981 = controllable_BtoR_REQ0 & ~n46980;
  assign n46982 = ~n17692 & ~n46981;
  assign n46983 = i_RtoB_ACK0 & ~n46982;
  assign n46984 = ~n46677 & ~n46983;
  assign n46985 = ~controllable_DEQ & ~n46984;
  assign n46986 = ~n29092 & ~n46985;
  assign n46987 = ~i_FULL & ~n46986;
  assign n46988 = ~n46977 & ~n46987;
  assign n46989 = ~i_nEMPTY & ~n46988;
  assign n46990 = ~n46967 & ~n46989;
  assign n46991 = ~controllable_BtoS_ACK0 & ~n46990;
  assign n46992 = ~n46951 & ~n46991;
  assign n46993 = n4465 & ~n46992;
  assign n46994 = ~n46695 & ~n46993;
  assign n46995 = i_StoB_REQ10 & ~n46994;
  assign n46996 = ~n46909 & ~n46995;
  assign n46997 = ~controllable_BtoS_ACK10 & ~n46996;
  assign n46998 = ~n46911 & ~n46997;
  assign n46999 = n4464 & ~n46998;
  assign n47000 = ~n46761 & ~n46999;
  assign n47001 = ~n4463 & ~n47000;
  assign n47002 = ~n46763 & ~n47001;
  assign n47003 = n4462 & ~n47002;
  assign n47004 = ~n29030 & ~n29473;
  assign n47005 = i_FULL & ~n47004;
  assign n47006 = ~n29480 & ~n47005;
  assign n47007 = i_nEMPTY & ~n47006;
  assign n47008 = ~n29492 & ~n47007;
  assign n47009 = controllable_BtoS_ACK0 & ~n47008;
  assign n47010 = ~n46693 & ~n47009;
  assign n47011 = n4465 & ~n47010;
  assign n47012 = ~n46695 & ~n47011;
  assign n47013 = i_StoB_REQ10 & ~n47012;
  assign n47014 = ~n17626 & ~n29514;
  assign n47015 = i_FULL & ~n47014;
  assign n47016 = ~n29526 & ~n47015;
  assign n47017 = i_nEMPTY & ~n47016;
  assign n47018 = ~n29546 & ~n47017;
  assign n47019 = controllable_BtoS_ACK0 & ~n47018;
  assign n47020 = ~n46569 & ~n47019;
  assign n47021 = n4465 & ~n47020;
  assign n47022 = ~n46571 & ~n47021;
  assign n47023 = ~i_StoB_REQ10 & ~n47022;
  assign n47024 = ~n47013 & ~n47023;
  assign n47025 = ~controllable_BtoS_ACK10 & ~n47024;
  assign n47026 = ~n29467 & ~n47025;
  assign n47027 = n4464 & ~n47026;
  assign n47028 = ~n29467 & ~n46759;
  assign n47029 = ~n4464 & ~n47028;
  assign n47030 = ~n47027 & ~n47029;
  assign n47031 = ~n4462 & ~n47030;
  assign n47032 = ~n47003 & ~n47031;
  assign n47033 = n4461 & ~n47032;
  assign n47034 = ~n7111 & ~n36879;
  assign n47035 = ~controllable_BtoR_REQ1 & ~n47034;
  assign n47036 = ~controllable_BtoR_REQ1 & ~n47035;
  assign n47037 = controllable_BtoR_REQ0 & ~n47036;
  assign n47038 = ~controllable_BtoR_REQ1 & ~n45752;
  assign n47039 = ~controllable_BtoR_REQ1 & ~n47038;
  assign n47040 = ~controllable_BtoR_REQ0 & ~n47039;
  assign n47041 = ~n47037 & ~n47040;
  assign n47042 = ~i_RtoB_ACK0 & ~n47041;
  assign n47043 = ~n46765 & ~n47042;
  assign n47044 = ~controllable_DEQ & ~n47043;
  assign n47045 = ~n14755 & ~n47044;
  assign n47046 = i_nEMPTY & ~n47045;
  assign n47047 = ~n7054 & ~n36914;
  assign n47048 = ~controllable_BtoR_REQ1 & ~n47047;
  assign n47049 = ~controllable_BtoR_REQ1 & ~n47048;
  assign n47050 = controllable_BtoR_REQ0 & ~n47049;
  assign n47051 = ~controllable_BtoR_REQ1 & ~n45764;
  assign n47052 = ~controllable_BtoR_REQ1 & ~n47051;
  assign n47053 = ~controllable_BtoR_REQ0 & ~n47052;
  assign n47054 = ~n47050 & ~n47053;
  assign n47055 = ~i_RtoB_ACK0 & ~n47054;
  assign n47056 = ~n46777 & ~n47055;
  assign n47057 = ~controllable_DEQ & ~n47056;
  assign n47058 = ~n14780 & ~n47057;
  assign n47059 = i_FULL & ~n47058;
  assign n47060 = ~n7054 & ~n45773;
  assign n47061 = ~controllable_BtoR_REQ1 & ~n47060;
  assign n47062 = ~controllable_BtoR_REQ1 & ~n47061;
  assign n47063 = controllable_BtoR_REQ0 & ~n47062;
  assign n47064 = ~controllable_BtoR_REQ1 & ~n45774;
  assign n47065 = ~controllable_BtoR_REQ1 & ~n47064;
  assign n47066 = ~controllable_BtoR_REQ0 & ~n47065;
  assign n47067 = ~n47063 & ~n47066;
  assign n47068 = ~i_RtoB_ACK0 & ~n47067;
  assign n47069 = ~n46777 & ~n47068;
  assign n47070 = ~controllable_DEQ & ~n47069;
  assign n47071 = ~n14798 & ~n47070;
  assign n47072 = ~i_FULL & ~n47071;
  assign n47073 = ~n47059 & ~n47072;
  assign n47074 = ~i_nEMPTY & ~n47073;
  assign n47075 = ~n47046 & ~n47074;
  assign n47076 = controllable_BtoS_ACK0 & ~n47075;
  assign n47077 = ~n11324 & ~n37060;
  assign n47078 = ~controllable_BtoR_REQ1 & ~n47077;
  assign n47079 = ~controllable_BtoR_REQ1 & ~n47078;
  assign n47080 = controllable_BtoR_REQ0 & ~n47079;
  assign n47081 = ~controllable_BtoR_REQ1 & ~n45790;
  assign n47082 = ~controllable_BtoR_REQ1 & ~n47081;
  assign n47083 = ~controllable_BtoR_REQ0 & ~n47082;
  assign n47084 = ~n47080 & ~n47083;
  assign n47085 = ~i_RtoB_ACK0 & ~n47084;
  assign n47086 = ~n46791 & ~n47085;
  assign n47087 = ~controllable_DEQ & ~n47086;
  assign n47088 = ~n28757 & ~n47087;
  assign n47089 = i_nEMPTY & ~n47088;
  assign n47090 = ~n11299 & ~n37095;
  assign n47091 = ~controllable_BtoR_REQ1 & ~n47090;
  assign n47092 = ~controllable_BtoR_REQ1 & ~n47091;
  assign n47093 = controllable_BtoR_REQ0 & ~n47092;
  assign n47094 = ~controllable_BtoR_REQ1 & ~n45802;
  assign n47095 = ~controllable_BtoR_REQ1 & ~n47094;
  assign n47096 = ~controllable_BtoR_REQ0 & ~n47095;
  assign n47097 = ~n47093 & ~n47096;
  assign n47098 = ~i_RtoB_ACK0 & ~n47097;
  assign n47099 = ~n46803 & ~n47098;
  assign n47100 = ~controllable_DEQ & ~n47099;
  assign n47101 = ~n28773 & ~n47100;
  assign n47102 = i_FULL & ~n47101;
  assign n47103 = ~n11299 & ~n45811;
  assign n47104 = ~controllable_BtoR_REQ1 & ~n47103;
  assign n47105 = ~controllable_BtoR_REQ1 & ~n47104;
  assign n47106 = controllable_BtoR_REQ0 & ~n47105;
  assign n47107 = ~controllable_BtoR_REQ1 & ~n45812;
  assign n47108 = ~controllable_BtoR_REQ1 & ~n47107;
  assign n47109 = ~controllable_BtoR_REQ0 & ~n47108;
  assign n47110 = ~n47106 & ~n47109;
  assign n47111 = ~i_RtoB_ACK0 & ~n47110;
  assign n47112 = ~n46803 & ~n47111;
  assign n47113 = ~controllable_DEQ & ~n47112;
  assign n47114 = ~n28787 & ~n47113;
  assign n47115 = ~i_FULL & ~n47114;
  assign n47116 = ~n47102 & ~n47115;
  assign n47117 = ~i_nEMPTY & ~n47116;
  assign n47118 = ~n47089 & ~n47117;
  assign n47119 = ~controllable_BtoS_ACK0 & ~n47118;
  assign n47120 = ~n47076 & ~n47119;
  assign n47121 = n4465 & ~n47120;
  assign n47122 = ~n4465 & ~n29464;
  assign n47123 = ~n47121 & ~n47122;
  assign n47124 = i_StoB_REQ10 & ~n47123;
  assign n47125 = ~n7111 & ~n46820;
  assign n47126 = ~controllable_BtoR_REQ1 & ~n47125;
  assign n47127 = ~controllable_BtoR_REQ1 & ~n47126;
  assign n47128 = controllable_BtoR_REQ0 & ~n47127;
  assign n47129 = ~n46409 & ~n47128;
  assign n47130 = i_RtoB_ACK0 & ~n47129;
  assign n47131 = ~n17631 & ~n37915;
  assign n47132 = ~controllable_BtoR_REQ1 & ~n47131;
  assign n47133 = ~controllable_BtoR_REQ1 & ~n47132;
  assign n47134 = controllable_BtoR_REQ0 & ~n47133;
  assign n47135 = ~controllable_BtoR_REQ1 & ~n45833;
  assign n47136 = ~controllable_BtoR_REQ1 & ~n47135;
  assign n47137 = ~controllable_BtoR_REQ0 & ~n47136;
  assign n47138 = ~n47134 & ~n47137;
  assign n47139 = ~i_RtoB_ACK0 & ~n47138;
  assign n47140 = ~n47130 & ~n47139;
  assign n47141 = ~controllable_DEQ & ~n47140;
  assign n47142 = ~n17626 & ~n47141;
  assign n47143 = i_nEMPTY & ~n47142;
  assign n47144 = ~n7054 & ~n46837;
  assign n47145 = ~controllable_BtoR_REQ1 & ~n47144;
  assign n47146 = ~controllable_BtoR_REQ1 & ~n47145;
  assign n47147 = controllable_BtoR_REQ0 & ~n47146;
  assign n47148 = ~n46444 & ~n47147;
  assign n47149 = i_RtoB_ACK0 & ~n47148;
  assign n47150 = ~n17616 & ~n37948;
  assign n47151 = ~controllable_BtoR_REQ1 & ~n47150;
  assign n47152 = ~controllable_BtoR_REQ1 & ~n47151;
  assign n47153 = controllable_BtoR_REQ0 & ~n47152;
  assign n47154 = ~controllable_BtoR_REQ1 & ~n45845;
  assign n47155 = ~controllable_BtoR_REQ1 & ~n47154;
  assign n47156 = ~controllable_BtoR_REQ0 & ~n47155;
  assign n47157 = ~n47153 & ~n47156;
  assign n47158 = ~i_RtoB_ACK0 & ~n47157;
  assign n47159 = ~n47149 & ~n47158;
  assign n47160 = ~controllable_DEQ & ~n47159;
  assign n47161 = ~n17651 & ~n47160;
  assign n47162 = i_FULL & ~n47161;
  assign n47163 = ~n7054 & ~n46848;
  assign n47164 = ~controllable_BtoR_REQ1 & ~n47163;
  assign n47165 = ~controllable_BtoR_REQ1 & ~n47164;
  assign n47166 = controllable_BtoR_REQ0 & ~n47165;
  assign n47167 = ~n46444 & ~n47166;
  assign n47168 = i_RtoB_ACK0 & ~n47167;
  assign n47169 = ~n17616 & ~n45856;
  assign n47170 = ~controllable_BtoR_REQ1 & ~n47169;
  assign n47171 = ~controllable_BtoR_REQ1 & ~n47170;
  assign n47172 = controllable_BtoR_REQ0 & ~n47171;
  assign n47173 = ~controllable_BtoR_REQ1 & ~n45860;
  assign n47174 = ~controllable_BtoR_REQ0 & ~n47173;
  assign n47175 = ~n47172 & ~n47174;
  assign n47176 = ~i_RtoB_ACK0 & ~n47175;
  assign n47177 = ~n47168 & ~n47176;
  assign n47178 = ~controllable_DEQ & ~n47177;
  assign n47179 = ~n17673 & ~n47178;
  assign n47180 = ~i_FULL & ~n47179;
  assign n47181 = ~n47162 & ~n47180;
  assign n47182 = ~i_nEMPTY & ~n47181;
  assign n47183 = ~n47143 & ~n47182;
  assign n47184 = controllable_BtoS_ACK0 & ~n47183;
  assign n47185 = ~n11324 & ~n46863;
  assign n47186 = ~controllable_BtoR_REQ1 & ~n47185;
  assign n47187 = ~controllable_BtoR_REQ1 & ~n47186;
  assign n47188 = controllable_BtoR_REQ0 & ~n47187;
  assign n47189 = ~n46488 & ~n47188;
  assign n47190 = i_RtoB_ACK0 & ~n47189;
  assign n47191 = ~n17714 & ~n37999;
  assign n47192 = ~controllable_BtoR_REQ1 & ~n47191;
  assign n47193 = ~controllable_BtoR_REQ1 & ~n47192;
  assign n47194 = controllable_BtoR_REQ0 & ~n47193;
  assign n47195 = ~controllable_BtoR_REQ1 & ~n45877;
  assign n47196 = ~controllable_BtoR_REQ1 & ~n47195;
  assign n47197 = ~controllable_BtoR_REQ0 & ~n47196;
  assign n47198 = ~n47194 & ~n47197;
  assign n47199 = ~i_RtoB_ACK0 & ~n47198;
  assign n47200 = ~n47190 & ~n47199;
  assign n47201 = ~controllable_DEQ & ~n47200;
  assign n47202 = ~n17705 & ~n47201;
  assign n47203 = i_nEMPTY & ~n47202;
  assign n47204 = ~n11299 & ~n46880;
  assign n47205 = ~controllable_BtoR_REQ1 & ~n47204;
  assign n47206 = ~controllable_BtoR_REQ1 & ~n47205;
  assign n47207 = controllable_BtoR_REQ0 & ~n47206;
  assign n47208 = ~n46523 & ~n47207;
  assign n47209 = i_RtoB_ACK0 & ~n47208;
  assign n47210 = ~n17695 & ~n38032;
  assign n47211 = ~controllable_BtoR_REQ1 & ~n47210;
  assign n47212 = ~controllable_BtoR_REQ1 & ~n47211;
  assign n47213 = controllable_BtoR_REQ0 & ~n47212;
  assign n47214 = ~controllable_BtoR_REQ1 & ~n45889;
  assign n47215 = ~controllable_BtoR_REQ1 & ~n47214;
  assign n47216 = ~controllable_BtoR_REQ0 & ~n47215;
  assign n47217 = ~n47213 & ~n47216;
  assign n47218 = ~i_RtoB_ACK0 & ~n47217;
  assign n47219 = ~n47209 & ~n47218;
  assign n47220 = ~controllable_DEQ & ~n47219;
  assign n47221 = ~n17741 & ~n47220;
  assign n47222 = i_FULL & ~n47221;
  assign n47223 = ~n11299 & ~n46891;
  assign n47224 = ~controllable_BtoR_REQ1 & ~n47223;
  assign n47225 = ~controllable_BtoR_REQ1 & ~n47224;
  assign n47226 = controllable_BtoR_REQ0 & ~n47225;
  assign n47227 = ~n46523 & ~n47226;
  assign n47228 = i_RtoB_ACK0 & ~n47227;
  assign n47229 = ~n17695 & ~n45900;
  assign n47230 = ~controllable_BtoR_REQ1 & ~n47229;
  assign n47231 = ~controllable_BtoR_REQ1 & ~n47230;
  assign n47232 = controllable_BtoR_REQ0 & ~n47231;
  assign n47233 = ~controllable_BtoR_REQ1 & ~n45904;
  assign n47234 = ~controllable_BtoR_REQ0 & ~n47233;
  assign n47235 = ~n47232 & ~n47234;
  assign n47236 = ~i_RtoB_ACK0 & ~n47235;
  assign n47237 = ~n47228 & ~n47236;
  assign n47238 = ~controllable_DEQ & ~n47237;
  assign n47239 = ~n17774 & ~n47238;
  assign n47240 = ~i_FULL & ~n47239;
  assign n47241 = ~n47222 & ~n47240;
  assign n47242 = ~i_nEMPTY & ~n47241;
  assign n47243 = ~n47203 & ~n47242;
  assign n47244 = ~controllable_BtoS_ACK0 & ~n47243;
  assign n47245 = ~n47184 & ~n47244;
  assign n47246 = n4465 & ~n47245;
  assign n47247 = ~n4465 & ~n17787;
  assign n47248 = ~n47246 & ~n47247;
  assign n47249 = ~i_StoB_REQ10 & ~n47248;
  assign n47250 = ~n47124 & ~n47249;
  assign n47251 = controllable_BtoS_ACK10 & ~n47250;
  assign n47252 = ~controllable_BtoR_REQ1 & ~n45924;
  assign n47253 = ~controllable_BtoR_REQ1 & ~n47252;
  assign n47254 = ~i_RtoB_ACK0 & ~n47253;
  assign n47255 = ~n29022 & ~n47254;
  assign n47256 = ~controllable_DEQ & ~n47255;
  assign n47257 = ~n29030 & ~n47256;
  assign n47258 = i_nEMPTY & ~n47257;
  assign n47259 = ~controllable_BtoR_REQ1 & ~n45932;
  assign n47260 = ~controllable_BtoR_REQ1 & ~n47259;
  assign n47261 = ~i_RtoB_ACK0 & ~n47260;
  assign n47262 = ~n29042 & ~n47261;
  assign n47263 = ~controllable_DEQ & ~n47262;
  assign n47264 = ~n29040 & ~n47263;
  assign n47265 = i_FULL & ~n47264;
  assign n47266 = ~n5237 & ~n40128;
  assign n47267 = ~controllable_BtoR_REQ1 & ~n47266;
  assign n47268 = ~controllable_BtoR_REQ1 & ~n47267;
  assign n47269 = controllable_BtoR_REQ0 & ~n47268;
  assign n47270 = ~n17613 & ~n47269;
  assign n47271 = i_RtoB_ACK0 & ~n47270;
  assign n47272 = ~controllable_BtoR_REQ1 & ~n45943;
  assign n47273 = ~i_RtoB_ACK0 & ~n47272;
  assign n47274 = ~n47271 & ~n47273;
  assign n47275 = ~controllable_DEQ & ~n47274;
  assign n47276 = ~n29050 & ~n47275;
  assign n47277 = ~i_FULL & ~n47276;
  assign n47278 = ~n47265 & ~n47277;
  assign n47279 = ~i_nEMPTY & ~n47278;
  assign n47280 = ~n47258 & ~n47279;
  assign n47281 = controllable_BtoS_ACK0 & ~n47280;
  assign n47282 = ~controllable_BtoR_REQ1 & ~n45956;
  assign n47283 = ~controllable_BtoR_REQ1 & ~n47282;
  assign n47284 = ~i_RtoB_ACK0 & ~n47283;
  assign n47285 = ~n29064 & ~n47284;
  assign n47286 = ~controllable_DEQ & ~n47285;
  assign n47287 = ~n29072 & ~n47286;
  assign n47288 = i_nEMPTY & ~n47287;
  assign n47289 = ~controllable_BtoR_REQ1 & ~n45964;
  assign n47290 = ~controllable_BtoR_REQ1 & ~n47289;
  assign n47291 = ~i_RtoB_ACK0 & ~n47290;
  assign n47292 = ~n29084 & ~n47291;
  assign n47293 = ~controllable_DEQ & ~n47292;
  assign n47294 = ~n29082 & ~n47293;
  assign n47295 = i_FULL & ~n47294;
  assign n47296 = ~n8861 & ~n40189;
  assign n47297 = ~controllable_BtoR_REQ1 & ~n47296;
  assign n47298 = ~controllable_BtoR_REQ1 & ~n47297;
  assign n47299 = controllable_BtoR_REQ0 & ~n47298;
  assign n47300 = ~n17692 & ~n47299;
  assign n47301 = i_RtoB_ACK0 & ~n47300;
  assign n47302 = ~controllable_BtoR_REQ1 & ~n45975;
  assign n47303 = ~i_RtoB_ACK0 & ~n47302;
  assign n47304 = ~n47301 & ~n47303;
  assign n47305 = ~controllable_DEQ & ~n47304;
  assign n47306 = ~n29092 & ~n47305;
  assign n47307 = ~i_FULL & ~n47306;
  assign n47308 = ~n47295 & ~n47307;
  assign n47309 = ~i_nEMPTY & ~n47308;
  assign n47310 = ~n47288 & ~n47309;
  assign n47311 = ~controllable_BtoS_ACK0 & ~n47310;
  assign n47312 = ~n47281 & ~n47311;
  assign n47313 = n4465 & ~n47312;
  assign n47314 = ~n4465 & ~n29580;
  assign n47315 = ~n47313 & ~n47314;
  assign n47316 = i_StoB_REQ10 & ~n47315;
  assign n47317 = ~n47249 & ~n47316;
  assign n47318 = ~controllable_BtoS_ACK10 & ~n47317;
  assign n47319 = ~n47251 & ~n47318;
  assign n47320 = n4464 & ~n47319;
  assign n47321 = ~n4464 & ~n29584;
  assign n47322 = ~n47320 & ~n47321;
  assign n47323 = n4462 & ~n47322;
  assign n47324 = ~n4462 & ~n29584;
  assign n47325 = ~n47323 & ~n47324;
  assign n47326 = ~n4461 & ~n47325;
  assign n47327 = ~n47033 & ~n47326;
  assign n47328 = n4459 & ~n47327;
  assign n47329 = ~n46263 & ~n47328;
  assign n47330 = n4455 & ~n47329;
  assign n47331 = ~n39895 & ~n45155;
  assign n47332 = i_RtoB_ACK0 & ~n47331;
  assign n47333 = ~n45160 & ~n46272;
  assign n47334 = ~i_RtoB_ACK0 & ~n47333;
  assign n47335 = ~n47332 & ~n47334;
  assign n47336 = ~controllable_DEQ & ~n47335;
  assign n47337 = ~n20981 & ~n47336;
  assign n47338 = i_FULL & ~n47337;
  assign n47339 = ~n45171 & ~n46284;
  assign n47340 = ~i_RtoB_ACK0 & ~n47339;
  assign n47341 = ~n47332 & ~n47340;
  assign n47342 = ~controllable_DEQ & ~n47341;
  assign n47343 = ~n20981 & ~n47342;
  assign n47344 = ~i_FULL & ~n47343;
  assign n47345 = ~n47338 & ~n47344;
  assign n47346 = i_nEMPTY & ~n47345;
  assign n47347 = ~n39905 & ~n45187;
  assign n47348 = i_RtoB_ACK0 & ~n47347;
  assign n47349 = ~n45192 & ~n46303;
  assign n47350 = ~i_RtoB_ACK0 & ~n47349;
  assign n47351 = ~n47348 & ~n47350;
  assign n47352 = ~controllable_DEQ & ~n47351;
  assign n47353 = ~n20993 & ~n47352;
  assign n47354 = i_FULL & ~n47353;
  assign n47355 = ~n45203 & ~n46315;
  assign n47356 = ~i_RtoB_ACK0 & ~n47355;
  assign n47357 = ~n47348 & ~n47356;
  assign n47358 = ~controllable_DEQ & ~n47357;
  assign n47359 = ~n21003 & ~n47358;
  assign n47360 = ~i_FULL & ~n47359;
  assign n47361 = ~n47354 & ~n47360;
  assign n47362 = ~i_nEMPTY & ~n47361;
  assign n47363 = ~n47346 & ~n47362;
  assign n47364 = controllable_BtoS_ACK0 & ~n47363;
  assign n47365 = ~n39923 & ~n45219;
  assign n47366 = i_RtoB_ACK0 & ~n47365;
  assign n47367 = ~n45224 & ~n46336;
  assign n47368 = ~i_RtoB_ACK0 & ~n47367;
  assign n47369 = ~n47366 & ~n47368;
  assign n47370 = ~controllable_DEQ & ~n47369;
  assign n47371 = ~n29641 & ~n47370;
  assign n47372 = i_FULL & ~n47371;
  assign n47373 = ~n45235 & ~n46348;
  assign n47374 = ~i_RtoB_ACK0 & ~n47373;
  assign n47375 = ~n47366 & ~n47374;
  assign n47376 = ~controllable_DEQ & ~n47375;
  assign n47377 = ~n29641 & ~n47376;
  assign n47378 = ~i_FULL & ~n47377;
  assign n47379 = ~n47372 & ~n47378;
  assign n47380 = i_nEMPTY & ~n47379;
  assign n47381 = ~n39933 & ~n45251;
  assign n47382 = i_RtoB_ACK0 & ~n47381;
  assign n47383 = ~n45256 & ~n46367;
  assign n47384 = ~i_RtoB_ACK0 & ~n47383;
  assign n47385 = ~n47382 & ~n47384;
  assign n47386 = ~controllable_DEQ & ~n47385;
  assign n47387 = ~n29653 & ~n47386;
  assign n47388 = i_FULL & ~n47387;
  assign n47389 = ~n45267 & ~n46379;
  assign n47390 = ~i_RtoB_ACK0 & ~n47389;
  assign n47391 = ~n47382 & ~n47390;
  assign n47392 = ~controllable_DEQ & ~n47391;
  assign n47393 = ~n29663 & ~n47392;
  assign n47394 = ~i_FULL & ~n47393;
  assign n47395 = ~n47388 & ~n47394;
  assign n47396 = ~i_nEMPTY & ~n47395;
  assign n47397 = ~n47380 & ~n47396;
  assign n47398 = ~controllable_BtoS_ACK0 & ~n47397;
  assign n47399 = ~n47364 & ~n47398;
  assign n47400 = n4465 & ~n47399;
  assign n47401 = ~n29641 & ~n29683;
  assign n47402 = i_FULL & ~n47401;
  assign n47403 = ~n29691 & ~n47402;
  assign n47404 = i_nEMPTY & ~n47403;
  assign n47405 = ~n29707 & ~n47404;
  assign n47406 = ~controllable_BtoS_ACK0 & ~n47405;
  assign n47407 = ~n21013 & ~n47406;
  assign n47408 = ~n4465 & ~n47407;
  assign n47409 = ~n47400 & ~n47408;
  assign n47410 = i_StoB_REQ10 & ~n47409;
  assign n47411 = ~n45382 & ~n46407;
  assign n47412 = i_RtoB_ACK0 & ~n47411;
  assign n47413 = ~n45390 & ~n46416;
  assign n47414 = ~i_RtoB_ACK0 & ~n47413;
  assign n47415 = ~n47412 & ~n47414;
  assign n47416 = ~controllable_DEQ & ~n47415;
  assign n47417 = ~n23093 & ~n47416;
  assign n47418 = i_FULL & ~n47417;
  assign n47419 = ~n45401 & ~n46428;
  assign n47420 = ~i_RtoB_ACK0 & ~n47419;
  assign n47421 = ~n47412 & ~n47420;
  assign n47422 = ~controllable_DEQ & ~n47421;
  assign n47423 = ~n23093 & ~n47422;
  assign n47424 = ~i_FULL & ~n47423;
  assign n47425 = ~n47418 & ~n47424;
  assign n47426 = i_nEMPTY & ~n47425;
  assign n47427 = ~n45422 & ~n46442;
  assign n47428 = i_RtoB_ACK0 & ~n47427;
  assign n47429 = ~n45430 & ~n46451;
  assign n47430 = ~i_RtoB_ACK0 & ~n47429;
  assign n47431 = ~n47428 & ~n47430;
  assign n47432 = ~controllable_DEQ & ~n47431;
  assign n47433 = ~n23105 & ~n47432;
  assign n47434 = i_FULL & ~n47433;
  assign n47435 = ~n45422 & ~n46464;
  assign n47436 = i_RtoB_ACK0 & ~n47435;
  assign n47437 = ~n45444 & ~n46470;
  assign n47438 = ~i_RtoB_ACK0 & ~n47437;
  assign n47439 = ~n47436 & ~n47438;
  assign n47440 = ~controllable_DEQ & ~n47439;
  assign n47441 = ~n23117 & ~n47440;
  assign n47442 = ~i_FULL & ~n47441;
  assign n47443 = ~n47434 & ~n47442;
  assign n47444 = ~i_nEMPTY & ~n47443;
  assign n47445 = ~n47426 & ~n47444;
  assign n47446 = controllable_BtoS_ACK0 & ~n47445;
  assign n47447 = ~n45467 & ~n46486;
  assign n47448 = i_RtoB_ACK0 & ~n47447;
  assign n47449 = ~n45475 & ~n46495;
  assign n47450 = ~i_RtoB_ACK0 & ~n47449;
  assign n47451 = ~n47448 & ~n47450;
  assign n47452 = ~controllable_DEQ & ~n47451;
  assign n47453 = ~n23133 & ~n47452;
  assign n47454 = i_FULL & ~n47453;
  assign n47455 = ~n45486 & ~n46507;
  assign n47456 = ~i_RtoB_ACK0 & ~n47455;
  assign n47457 = ~n47448 & ~n47456;
  assign n47458 = ~controllable_DEQ & ~n47457;
  assign n47459 = ~n23133 & ~n47458;
  assign n47460 = ~i_FULL & ~n47459;
  assign n47461 = ~n47454 & ~n47460;
  assign n47462 = i_nEMPTY & ~n47461;
  assign n47463 = ~n45507 & ~n46521;
  assign n47464 = i_RtoB_ACK0 & ~n47463;
  assign n47465 = ~n45515 & ~n46530;
  assign n47466 = ~i_RtoB_ACK0 & ~n47465;
  assign n47467 = ~n47464 & ~n47466;
  assign n47468 = ~controllable_DEQ & ~n47467;
  assign n47469 = ~n23145 & ~n47468;
  assign n47470 = i_FULL & ~n47469;
  assign n47471 = ~n45507 & ~n46543;
  assign n47472 = i_RtoB_ACK0 & ~n47471;
  assign n47473 = ~n45529 & ~n46549;
  assign n47474 = ~i_RtoB_ACK0 & ~n47473;
  assign n47475 = ~n47472 & ~n47474;
  assign n47476 = ~controllable_DEQ & ~n47475;
  assign n47477 = ~n23157 & ~n47476;
  assign n47478 = ~i_FULL & ~n47477;
  assign n47479 = ~n47470 & ~n47478;
  assign n47480 = ~i_nEMPTY & ~n47479;
  assign n47481 = ~n47462 & ~n47480;
  assign n47482 = ~controllable_BtoS_ACK0 & ~n47481;
  assign n47483 = ~n47446 & ~n47482;
  assign n47484 = n4465 & ~n47483;
  assign n47485 = ~n23133 & ~n29791;
  assign n47486 = i_FULL & ~n47485;
  assign n47487 = ~n29799 & ~n47486;
  assign n47488 = i_nEMPTY & ~n47487;
  assign n47489 = ~n29815 & ~n47488;
  assign n47490 = ~controllable_BtoS_ACK0 & ~n47489;
  assign n47491 = ~n23127 & ~n47490;
  assign n47492 = ~n4465 & ~n47491;
  assign n47493 = ~n47484 & ~n47492;
  assign n47494 = ~i_StoB_REQ10 & ~n47493;
  assign n47495 = ~n47410 & ~n47494;
  assign n47496 = controllable_BtoS_ACK10 & ~n47495;
  assign n47497 = ~n45557 & ~n46578;
  assign n47498 = i_RtoB_ACK0 & ~n47497;
  assign n47499 = ~n45561 & ~n46581;
  assign n47500 = ~i_RtoB_ACK0 & ~n47499;
  assign n47501 = ~n47498 & ~n47500;
  assign n47502 = ~controllable_DEQ & ~n47501;
  assign n47503 = ~n29844 & ~n47502;
  assign n47504 = i_FULL & ~n47503;
  assign n47505 = ~n45571 & ~n46588;
  assign n47506 = ~i_RtoB_ACK0 & ~n47505;
  assign n47507 = ~n47498 & ~n47506;
  assign n47508 = ~controllable_DEQ & ~n47507;
  assign n47509 = ~n29844 & ~n47508;
  assign n47510 = ~i_FULL & ~n47509;
  assign n47511 = ~n47504 & ~n47510;
  assign n47512 = i_nEMPTY & ~n47511;
  assign n47513 = ~n45583 & ~n46601;
  assign n47514 = i_RtoB_ACK0 & ~n47513;
  assign n47515 = ~n45587 & ~n46604;
  assign n47516 = ~i_RtoB_ACK0 & ~n47515;
  assign n47517 = ~n47514 & ~n47516;
  assign n47518 = ~controllable_DEQ & ~n47517;
  assign n47519 = ~n29858 & ~n47518;
  assign n47520 = i_FULL & ~n47519;
  assign n47521 = ~n45583 & ~n46615;
  assign n47522 = i_RtoB_ACK0 & ~n47521;
  assign n47523 = ~n45601 & ~n46618;
  assign n47524 = ~i_RtoB_ACK0 & ~n47523;
  assign n47525 = ~n47522 & ~n47524;
  assign n47526 = ~controllable_DEQ & ~n47525;
  assign n47527 = ~n29872 & ~n47526;
  assign n47528 = ~i_FULL & ~n47527;
  assign n47529 = ~n47520 & ~n47528;
  assign n47530 = ~i_nEMPTY & ~n47529;
  assign n47531 = ~n47512 & ~n47530;
  assign n47532 = controllable_BtoS_ACK0 & ~n47531;
  assign n47533 = ~n45615 & ~n46633;
  assign n47534 = i_RtoB_ACK0 & ~n47533;
  assign n47535 = ~n45619 & ~n46636;
  assign n47536 = ~i_RtoB_ACK0 & ~n47535;
  assign n47537 = ~n47534 & ~n47536;
  assign n47538 = ~controllable_DEQ & ~n47537;
  assign n47539 = ~n29900 & ~n47538;
  assign n47540 = i_FULL & ~n47539;
  assign n47541 = ~n45629 & ~n46643;
  assign n47542 = ~i_RtoB_ACK0 & ~n47541;
  assign n47543 = ~n47534 & ~n47542;
  assign n47544 = ~controllable_DEQ & ~n47543;
  assign n47545 = ~n29900 & ~n47544;
  assign n47546 = ~i_FULL & ~n47545;
  assign n47547 = ~n47540 & ~n47546;
  assign n47548 = i_nEMPTY & ~n47547;
  assign n47549 = ~n45641 & ~n46656;
  assign n47550 = i_RtoB_ACK0 & ~n47549;
  assign n47551 = ~n45645 & ~n46659;
  assign n47552 = ~i_RtoB_ACK0 & ~n47551;
  assign n47553 = ~n47550 & ~n47552;
  assign n47554 = ~controllable_DEQ & ~n47553;
  assign n47555 = ~n29914 & ~n47554;
  assign n47556 = i_FULL & ~n47555;
  assign n47557 = ~n45641 & ~n46670;
  assign n47558 = i_RtoB_ACK0 & ~n47557;
  assign n47559 = ~n45659 & ~n46673;
  assign n47560 = ~i_RtoB_ACK0 & ~n47559;
  assign n47561 = ~n47558 & ~n47560;
  assign n47562 = ~controllable_DEQ & ~n47561;
  assign n47563 = ~n29928 & ~n47562;
  assign n47564 = ~i_FULL & ~n47563;
  assign n47565 = ~n47556 & ~n47564;
  assign n47566 = ~i_nEMPTY & ~n47565;
  assign n47567 = ~n47548 & ~n47566;
  assign n47568 = ~controllable_BtoS_ACK0 & ~n47567;
  assign n47569 = ~n47532 & ~n47568;
  assign n47570 = n4465 & ~n47569;
  assign n47571 = ~n29900 & ~n29968;
  assign n47572 = i_FULL & ~n47571;
  assign n47573 = ~n29977 & ~n47572;
  assign n47574 = i_nEMPTY & ~n47573;
  assign n47575 = ~n29991 & ~n47574;
  assign n47576 = ~controllable_BtoS_ACK0 & ~n47575;
  assign n47577 = ~n29958 & ~n47576;
  assign n47578 = ~n4465 & ~n47577;
  assign n47579 = ~n47570 & ~n47578;
  assign n47580 = i_StoB_REQ10 & ~n47579;
  assign n47581 = ~n47494 & ~n47580;
  assign n47582 = ~controllable_BtoS_ACK10 & ~n47581;
  assign n47583 = ~n47496 & ~n47582;
  assign n47584 = n4464 & ~n47583;
  assign n47585 = ~n20981 & ~n30009;
  assign n47586 = i_FULL & ~n47585;
  assign n47587 = ~n30017 & ~n47586;
  assign n47588 = i_nEMPTY & ~n47587;
  assign n47589 = ~n30033 & ~n47588;
  assign n47590 = controllable_BtoS_ACK0 & ~n47589;
  assign n47591 = ~n29641 & ~n30043;
  assign n47592 = i_FULL & ~n47591;
  assign n47593 = ~n30051 & ~n47592;
  assign n47594 = i_nEMPTY & ~n47593;
  assign n47595 = ~n30067 & ~n47594;
  assign n47596 = ~controllable_BtoS_ACK0 & ~n47595;
  assign n47597 = ~n47590 & ~n47596;
  assign n47598 = n4465 & ~n47597;
  assign n47599 = ~n21013 & ~n47596;
  assign n47600 = ~n4465 & ~n47599;
  assign n47601 = ~n47598 & ~n47600;
  assign n47602 = i_StoB_REQ10 & ~n47601;
  assign n47603 = ~n23093 & ~n30083;
  assign n47604 = i_FULL & ~n47603;
  assign n47605 = ~n30091 & ~n47604;
  assign n47606 = i_nEMPTY & ~n47605;
  assign n47607 = ~n30107 & ~n47606;
  assign n47608 = controllable_BtoS_ACK0 & ~n47607;
  assign n47609 = ~n23133 & ~n30117;
  assign n47610 = i_FULL & ~n47609;
  assign n47611 = ~n30125 & ~n47610;
  assign n47612 = i_nEMPTY & ~n47611;
  assign n47613 = ~n30141 & ~n47612;
  assign n47614 = ~controllable_BtoS_ACK0 & ~n47613;
  assign n47615 = ~n47608 & ~n47614;
  assign n47616 = n4465 & ~n47615;
  assign n47617 = ~n23127 & ~n47614;
  assign n47618 = ~n4465 & ~n47617;
  assign n47619 = ~n47616 & ~n47618;
  assign n47620 = ~i_StoB_REQ10 & ~n47619;
  assign n47621 = ~n47602 & ~n47620;
  assign n47622 = controllable_BtoS_ACK10 & ~n47621;
  assign n47623 = ~n29844 & ~n30161;
  assign n47624 = i_FULL & ~n47623;
  assign n47625 = ~n30170 & ~n47624;
  assign n47626 = i_nEMPTY & ~n47625;
  assign n47627 = ~n30184 & ~n47626;
  assign n47628 = controllable_BtoS_ACK0 & ~n47627;
  assign n47629 = ~n29900 & ~n30196;
  assign n47630 = i_FULL & ~n47629;
  assign n47631 = ~n30205 & ~n47630;
  assign n47632 = i_nEMPTY & ~n47631;
  assign n47633 = ~n30219 & ~n47632;
  assign n47634 = ~controllable_BtoS_ACK0 & ~n47633;
  assign n47635 = ~n47628 & ~n47634;
  assign n47636 = n4465 & ~n47635;
  assign n47637 = ~n29958 & ~n47634;
  assign n47638 = ~n4465 & ~n47637;
  assign n47639 = ~n47636 & ~n47638;
  assign n47640 = i_StoB_REQ10 & ~n47639;
  assign n47641 = ~n47620 & ~n47640;
  assign n47642 = ~controllable_BtoS_ACK10 & ~n47641;
  assign n47643 = ~n47622 & ~n47642;
  assign n47644 = ~n4464 & ~n47643;
  assign n47645 = ~n47584 & ~n47644;
  assign n47646 = n4463 & ~n47645;
  assign n47647 = ~n18434 & ~n45749;
  assign n47648 = i_RtoB_ACK0 & ~n47647;
  assign n47649 = ~n45753 & ~n46272;
  assign n47650 = ~i_RtoB_ACK0 & ~n47649;
  assign n47651 = ~n47648 & ~n47650;
  assign n47652 = ~controllable_DEQ & ~n47651;
  assign n47653 = ~n20981 & ~n47652;
  assign n47654 = i_FULL & ~n47653;
  assign n47655 = ~n45753 & ~n46284;
  assign n47656 = ~i_RtoB_ACK0 & ~n47655;
  assign n47657 = ~n47648 & ~n47656;
  assign n47658 = ~controllable_DEQ & ~n47657;
  assign n47659 = ~n20981 & ~n47658;
  assign n47660 = ~i_FULL & ~n47659;
  assign n47661 = ~n47654 & ~n47660;
  assign n47662 = i_nEMPTY & ~n47661;
  assign n47663 = ~n18428 & ~n45761;
  assign n47664 = i_RtoB_ACK0 & ~n47663;
  assign n47665 = ~n45765 & ~n46303;
  assign n47666 = ~i_RtoB_ACK0 & ~n47665;
  assign n47667 = ~n47664 & ~n47666;
  assign n47668 = ~controllable_DEQ & ~n47667;
  assign n47669 = ~n20993 & ~n47668;
  assign n47670 = i_FULL & ~n47669;
  assign n47671 = ~n45775 & ~n46315;
  assign n47672 = ~i_RtoB_ACK0 & ~n47671;
  assign n47673 = ~n47664 & ~n47672;
  assign n47674 = ~controllable_DEQ & ~n47673;
  assign n47675 = ~n21003 & ~n47674;
  assign n47676 = ~i_FULL & ~n47675;
  assign n47677 = ~n47670 & ~n47676;
  assign n47678 = ~i_nEMPTY & ~n47677;
  assign n47679 = ~n47662 & ~n47678;
  assign n47680 = controllable_BtoS_ACK0 & ~n47679;
  assign n47681 = ~n18462 & ~n45787;
  assign n47682 = i_RtoB_ACK0 & ~n47681;
  assign n47683 = ~n45791 & ~n46336;
  assign n47684 = ~i_RtoB_ACK0 & ~n47683;
  assign n47685 = ~n47682 & ~n47684;
  assign n47686 = ~controllable_DEQ & ~n47685;
  assign n47687 = ~n29641 & ~n47686;
  assign n47688 = i_FULL & ~n47687;
  assign n47689 = ~n45791 & ~n46348;
  assign n47690 = ~i_RtoB_ACK0 & ~n47689;
  assign n47691 = ~n47682 & ~n47690;
  assign n47692 = ~controllable_DEQ & ~n47691;
  assign n47693 = ~n29641 & ~n47692;
  assign n47694 = ~i_FULL & ~n47693;
  assign n47695 = ~n47688 & ~n47694;
  assign n47696 = i_nEMPTY & ~n47695;
  assign n47697 = ~n18456 & ~n45799;
  assign n47698 = i_RtoB_ACK0 & ~n47697;
  assign n47699 = ~n45803 & ~n46367;
  assign n47700 = ~i_RtoB_ACK0 & ~n47699;
  assign n47701 = ~n47698 & ~n47700;
  assign n47702 = ~controllable_DEQ & ~n47701;
  assign n47703 = ~n29653 & ~n47702;
  assign n47704 = i_FULL & ~n47703;
  assign n47705 = ~n45813 & ~n46379;
  assign n47706 = ~i_RtoB_ACK0 & ~n47705;
  assign n47707 = ~n47698 & ~n47706;
  assign n47708 = ~controllable_DEQ & ~n47707;
  assign n47709 = ~n29663 & ~n47708;
  assign n47710 = ~i_FULL & ~n47709;
  assign n47711 = ~n47704 & ~n47710;
  assign n47712 = ~i_nEMPTY & ~n47711;
  assign n47713 = ~n47696 & ~n47712;
  assign n47714 = ~controllable_BtoS_ACK0 & ~n47713;
  assign n47715 = ~n47680 & ~n47714;
  assign n47716 = n4465 & ~n47715;
  assign n47717 = ~n29641 & ~n30311;
  assign n47718 = i_FULL & ~n47717;
  assign n47719 = ~n30319 & ~n47718;
  assign n47720 = i_nEMPTY & ~n47719;
  assign n47721 = ~n30335 & ~n47720;
  assign n47722 = ~controllable_BtoS_ACK0 & ~n47721;
  assign n47723 = ~n21013 & ~n47722;
  assign n47724 = ~n4465 & ~n47723;
  assign n47725 = ~n47716 & ~n47724;
  assign n47726 = i_StoB_REQ10 & ~n47725;
  assign n47727 = ~n45830 & ~n46824;
  assign n47728 = i_RtoB_ACK0 & ~n47727;
  assign n47729 = ~n45834 & ~n46416;
  assign n47730 = ~i_RtoB_ACK0 & ~n47729;
  assign n47731 = ~n47728 & ~n47730;
  assign n47732 = ~controllable_DEQ & ~n47731;
  assign n47733 = ~n23093 & ~n47732;
  assign n47734 = i_FULL & ~n47733;
  assign n47735 = ~n45834 & ~n46428;
  assign n47736 = ~i_RtoB_ACK0 & ~n47735;
  assign n47737 = ~n47728 & ~n47736;
  assign n47738 = ~controllable_DEQ & ~n47737;
  assign n47739 = ~n23093 & ~n47738;
  assign n47740 = ~i_FULL & ~n47739;
  assign n47741 = ~n47734 & ~n47740;
  assign n47742 = i_nEMPTY & ~n47741;
  assign n47743 = ~n45842 & ~n46841;
  assign n47744 = i_RtoB_ACK0 & ~n47743;
  assign n47745 = ~n45846 & ~n46451;
  assign n47746 = ~i_RtoB_ACK0 & ~n47745;
  assign n47747 = ~n47744 & ~n47746;
  assign n47748 = ~controllable_DEQ & ~n47747;
  assign n47749 = ~n23105 & ~n47748;
  assign n47750 = i_FULL & ~n47749;
  assign n47751 = ~n45842 & ~n46852;
  assign n47752 = i_RtoB_ACK0 & ~n47751;
  assign n47753 = ~n45862 & ~n46470;
  assign n47754 = ~i_RtoB_ACK0 & ~n47753;
  assign n47755 = ~n47752 & ~n47754;
  assign n47756 = ~controllable_DEQ & ~n47755;
  assign n47757 = ~n23117 & ~n47756;
  assign n47758 = ~i_FULL & ~n47757;
  assign n47759 = ~n47750 & ~n47758;
  assign n47760 = ~i_nEMPTY & ~n47759;
  assign n47761 = ~n47742 & ~n47760;
  assign n47762 = controllable_BtoS_ACK0 & ~n47761;
  assign n47763 = ~n45874 & ~n46867;
  assign n47764 = i_RtoB_ACK0 & ~n47763;
  assign n47765 = ~n45878 & ~n46495;
  assign n47766 = ~i_RtoB_ACK0 & ~n47765;
  assign n47767 = ~n47764 & ~n47766;
  assign n47768 = ~controllable_DEQ & ~n47767;
  assign n47769 = ~n23133 & ~n47768;
  assign n47770 = i_FULL & ~n47769;
  assign n47771 = ~n45878 & ~n46507;
  assign n47772 = ~i_RtoB_ACK0 & ~n47771;
  assign n47773 = ~n47764 & ~n47772;
  assign n47774 = ~controllable_DEQ & ~n47773;
  assign n47775 = ~n23133 & ~n47774;
  assign n47776 = ~i_FULL & ~n47775;
  assign n47777 = ~n47770 & ~n47776;
  assign n47778 = i_nEMPTY & ~n47777;
  assign n47779 = ~n45886 & ~n46884;
  assign n47780 = i_RtoB_ACK0 & ~n47779;
  assign n47781 = ~n45890 & ~n46530;
  assign n47782 = ~i_RtoB_ACK0 & ~n47781;
  assign n47783 = ~n47780 & ~n47782;
  assign n47784 = ~controllable_DEQ & ~n47783;
  assign n47785 = ~n23145 & ~n47784;
  assign n47786 = i_FULL & ~n47785;
  assign n47787 = ~n45886 & ~n46895;
  assign n47788 = i_RtoB_ACK0 & ~n47787;
  assign n47789 = ~n45906 & ~n46549;
  assign n47790 = ~i_RtoB_ACK0 & ~n47789;
  assign n47791 = ~n47788 & ~n47790;
  assign n47792 = ~controllable_DEQ & ~n47791;
  assign n47793 = ~n23157 & ~n47792;
  assign n47794 = ~i_FULL & ~n47793;
  assign n47795 = ~n47786 & ~n47794;
  assign n47796 = ~i_nEMPTY & ~n47795;
  assign n47797 = ~n47778 & ~n47796;
  assign n47798 = ~controllable_BtoS_ACK0 & ~n47797;
  assign n47799 = ~n47762 & ~n47798;
  assign n47800 = n4465 & ~n47799;
  assign n47801 = ~n23133 & ~n30419;
  assign n47802 = i_FULL & ~n47801;
  assign n47803 = ~n30427 & ~n47802;
  assign n47804 = i_nEMPTY & ~n47803;
  assign n47805 = ~n30443 & ~n47804;
  assign n47806 = ~controllable_BtoS_ACK0 & ~n47805;
  assign n47807 = ~n23127 & ~n47806;
  assign n47808 = ~n4465 & ~n47807;
  assign n47809 = ~n47800 & ~n47808;
  assign n47810 = ~i_StoB_REQ10 & ~n47809;
  assign n47811 = ~n47726 & ~n47810;
  assign n47812 = controllable_BtoS_ACK10 & ~n47811;
  assign n47813 = ~n28125 & ~n46915;
  assign n47814 = i_RtoB_ACK0 & ~n47813;
  assign n47815 = ~n45925 & ~n46581;
  assign n47816 = ~i_RtoB_ACK0 & ~n47815;
  assign n47817 = ~n47814 & ~n47816;
  assign n47818 = ~controllable_DEQ & ~n47817;
  assign n47819 = ~n29844 & ~n47818;
  assign n47820 = i_FULL & ~n47819;
  assign n47821 = ~n45925 & ~n46588;
  assign n47822 = ~i_RtoB_ACK0 & ~n47821;
  assign n47823 = ~n47814 & ~n47822;
  assign n47824 = ~controllable_DEQ & ~n47823;
  assign n47825 = ~n29844 & ~n47824;
  assign n47826 = ~i_FULL & ~n47825;
  assign n47827 = ~n47820 & ~n47826;
  assign n47828 = i_nEMPTY & ~n47827;
  assign n47829 = ~n28112 & ~n46931;
  assign n47830 = i_RtoB_ACK0 & ~n47829;
  assign n47831 = ~n45933 & ~n46604;
  assign n47832 = ~i_RtoB_ACK0 & ~n47831;
  assign n47833 = ~n47830 & ~n47832;
  assign n47834 = ~controllable_DEQ & ~n47833;
  assign n47835 = ~n29858 & ~n47834;
  assign n47836 = i_FULL & ~n47835;
  assign n47837 = ~n28112 & ~n46941;
  assign n47838 = i_RtoB_ACK0 & ~n47837;
  assign n47839 = ~n45945 & ~n46618;
  assign n47840 = ~i_RtoB_ACK0 & ~n47839;
  assign n47841 = ~n47838 & ~n47840;
  assign n47842 = ~controllable_DEQ & ~n47841;
  assign n47843 = ~n29872 & ~n47842;
  assign n47844 = ~i_FULL & ~n47843;
  assign n47845 = ~n47836 & ~n47844;
  assign n47846 = ~i_nEMPTY & ~n47845;
  assign n47847 = ~n47828 & ~n47846;
  assign n47848 = controllable_BtoS_ACK0 & ~n47847;
  assign n47849 = ~n28186 & ~n46955;
  assign n47850 = i_RtoB_ACK0 & ~n47849;
  assign n47851 = ~n45957 & ~n46636;
  assign n47852 = ~i_RtoB_ACK0 & ~n47851;
  assign n47853 = ~n47850 & ~n47852;
  assign n47854 = ~controllable_DEQ & ~n47853;
  assign n47855 = ~n29900 & ~n47854;
  assign n47856 = i_FULL & ~n47855;
  assign n47857 = ~n45957 & ~n46643;
  assign n47858 = ~i_RtoB_ACK0 & ~n47857;
  assign n47859 = ~n47850 & ~n47858;
  assign n47860 = ~controllable_DEQ & ~n47859;
  assign n47861 = ~n29900 & ~n47860;
  assign n47862 = ~i_FULL & ~n47861;
  assign n47863 = ~n47856 & ~n47862;
  assign n47864 = i_nEMPTY & ~n47863;
  assign n47865 = ~n28173 & ~n46971;
  assign n47866 = i_RtoB_ACK0 & ~n47865;
  assign n47867 = ~n45965 & ~n46659;
  assign n47868 = ~i_RtoB_ACK0 & ~n47867;
  assign n47869 = ~n47866 & ~n47868;
  assign n47870 = ~controllable_DEQ & ~n47869;
  assign n47871 = ~n29914 & ~n47870;
  assign n47872 = i_FULL & ~n47871;
  assign n47873 = ~n28173 & ~n46981;
  assign n47874 = i_RtoB_ACK0 & ~n47873;
  assign n47875 = ~n45977 & ~n46673;
  assign n47876 = ~i_RtoB_ACK0 & ~n47875;
  assign n47877 = ~n47874 & ~n47876;
  assign n47878 = ~controllable_DEQ & ~n47877;
  assign n47879 = ~n29928 & ~n47878;
  assign n47880 = ~i_FULL & ~n47879;
  assign n47881 = ~n47872 & ~n47880;
  assign n47882 = ~i_nEMPTY & ~n47881;
  assign n47883 = ~n47864 & ~n47882;
  assign n47884 = ~controllable_BtoS_ACK0 & ~n47883;
  assign n47885 = ~n47848 & ~n47884;
  assign n47886 = n4465 & ~n47885;
  assign n47887 = ~n29900 & ~n30523;
  assign n47888 = i_FULL & ~n47887;
  assign n47889 = ~n30531 & ~n47888;
  assign n47890 = i_nEMPTY & ~n47889;
  assign n47891 = ~n30544 & ~n47890;
  assign n47892 = ~controllable_BtoS_ACK0 & ~n47891;
  assign n47893 = ~n29958 & ~n47892;
  assign n47894 = ~n4465 & ~n47893;
  assign n47895 = ~n47886 & ~n47894;
  assign n47896 = i_StoB_REQ10 & ~n47895;
  assign n47897 = ~n47810 & ~n47896;
  assign n47898 = ~controllable_BtoS_ACK10 & ~n47897;
  assign n47899 = ~n47812 & ~n47898;
  assign n47900 = n4464 & ~n47899;
  assign n47901 = ~n20981 & ~n30562;
  assign n47902 = i_FULL & ~n47901;
  assign n47903 = ~n30570 & ~n47902;
  assign n47904 = i_nEMPTY & ~n47903;
  assign n47905 = ~n30586 & ~n47904;
  assign n47906 = controllable_BtoS_ACK0 & ~n47905;
  assign n47907 = ~n29641 & ~n30596;
  assign n47908 = i_FULL & ~n47907;
  assign n47909 = ~n30604 & ~n47908;
  assign n47910 = i_nEMPTY & ~n47909;
  assign n47911 = ~n30620 & ~n47910;
  assign n47912 = ~controllable_BtoS_ACK0 & ~n47911;
  assign n47913 = ~n47906 & ~n47912;
  assign n47914 = n4465 & ~n47913;
  assign n47915 = ~n21013 & ~n47912;
  assign n47916 = ~n4465 & ~n47915;
  assign n47917 = ~n47914 & ~n47916;
  assign n47918 = i_StoB_REQ10 & ~n47917;
  assign n47919 = ~n23093 & ~n30636;
  assign n47920 = i_FULL & ~n47919;
  assign n47921 = ~n30644 & ~n47920;
  assign n47922 = i_nEMPTY & ~n47921;
  assign n47923 = ~n30660 & ~n47922;
  assign n47924 = controllable_BtoS_ACK0 & ~n47923;
  assign n47925 = ~n23133 & ~n30670;
  assign n47926 = i_FULL & ~n47925;
  assign n47927 = ~n30678 & ~n47926;
  assign n47928 = i_nEMPTY & ~n47927;
  assign n47929 = ~n30694 & ~n47928;
  assign n47930 = ~controllable_BtoS_ACK0 & ~n47929;
  assign n47931 = ~n47924 & ~n47930;
  assign n47932 = n4465 & ~n47931;
  assign n47933 = ~n23127 & ~n47930;
  assign n47934 = ~n4465 & ~n47933;
  assign n47935 = ~n47932 & ~n47934;
  assign n47936 = ~i_StoB_REQ10 & ~n47935;
  assign n47937 = ~n47918 & ~n47936;
  assign n47938 = controllable_BtoS_ACK10 & ~n47937;
  assign n47939 = ~n29844 & ~n30712;
  assign n47940 = i_FULL & ~n47939;
  assign n47941 = ~n30720 & ~n47940;
  assign n47942 = i_nEMPTY & ~n47941;
  assign n47943 = ~n30733 & ~n47942;
  assign n47944 = controllable_BtoS_ACK0 & ~n47943;
  assign n47945 = ~n29900 & ~n30743;
  assign n47946 = i_FULL & ~n47945;
  assign n47947 = ~n30751 & ~n47946;
  assign n47948 = i_nEMPTY & ~n47947;
  assign n47949 = ~n30764 & ~n47948;
  assign n47950 = ~controllable_BtoS_ACK0 & ~n47949;
  assign n47951 = ~n47944 & ~n47950;
  assign n47952 = n4465 & ~n47951;
  assign n47953 = ~n29958 & ~n47950;
  assign n47954 = ~n4465 & ~n47953;
  assign n47955 = ~n47952 & ~n47954;
  assign n47956 = i_StoB_REQ10 & ~n47955;
  assign n47957 = ~n47936 & ~n47956;
  assign n47958 = ~controllable_BtoS_ACK10 & ~n47957;
  assign n47959 = ~n47938 & ~n47958;
  assign n47960 = ~n4464 & ~n47959;
  assign n47961 = ~n47900 & ~n47960;
  assign n47962 = ~n4463 & ~n47961;
  assign n47963 = ~n47646 & ~n47962;
  assign n47964 = n4462 & ~n47963;
  assign n47965 = ~n29844 & ~n30816;
  assign n47966 = i_FULL & ~n47965;
  assign n47967 = ~n30825 & ~n47966;
  assign n47968 = i_nEMPTY & ~n47967;
  assign n47969 = ~n30839 & ~n47968;
  assign n47970 = controllable_BtoS_ACK0 & ~n47969;
  assign n47971 = ~n47576 & ~n47970;
  assign n47972 = n4465 & ~n47971;
  assign n47973 = ~n47578 & ~n47972;
  assign n47974 = i_StoB_REQ10 & ~n47973;
  assign n47975 = ~n23093 & ~n30853;
  assign n47976 = i_FULL & ~n47975;
  assign n47977 = ~n30861 & ~n47976;
  assign n47978 = i_nEMPTY & ~n47977;
  assign n47979 = ~n30877 & ~n47978;
  assign n47980 = controllable_BtoS_ACK0 & ~n47979;
  assign n47981 = ~n47490 & ~n47980;
  assign n47982 = n4465 & ~n47981;
  assign n47983 = ~n47492 & ~n47982;
  assign n47984 = ~i_StoB_REQ10 & ~n47983;
  assign n47985 = ~n47974 & ~n47984;
  assign n47986 = ~controllable_BtoS_ACK10 & ~n47985;
  assign n47987 = ~n30806 & ~n47986;
  assign n47988 = n4464 & ~n47987;
  assign n47989 = ~n30806 & ~n47642;
  assign n47990 = ~n4464 & ~n47989;
  assign n47991 = ~n47988 & ~n47990;
  assign n47992 = n4463 & ~n47991;
  assign n47993 = ~n29844 & ~n30899;
  assign n47994 = i_FULL & ~n47993;
  assign n47995 = ~n30907 & ~n47994;
  assign n47996 = i_nEMPTY & ~n47995;
  assign n47997 = ~n30920 & ~n47996;
  assign n47998 = controllable_BtoS_ACK0 & ~n47997;
  assign n47999 = ~n47892 & ~n47998;
  assign n48000 = n4465 & ~n47999;
  assign n48001 = ~n47894 & ~n48000;
  assign n48002 = i_StoB_REQ10 & ~n48001;
  assign n48003 = ~n23093 & ~n30934;
  assign n48004 = i_FULL & ~n48003;
  assign n48005 = ~n30942 & ~n48004;
  assign n48006 = i_nEMPTY & ~n48005;
  assign n48007 = ~n30958 & ~n48006;
  assign n48008 = controllable_BtoS_ACK0 & ~n48007;
  assign n48009 = ~n47806 & ~n48008;
  assign n48010 = n4465 & ~n48009;
  assign n48011 = ~n47808 & ~n48010;
  assign n48012 = ~i_StoB_REQ10 & ~n48011;
  assign n48013 = ~n48002 & ~n48012;
  assign n48014 = ~controllable_BtoS_ACK10 & ~n48013;
  assign n48015 = ~n30806 & ~n48014;
  assign n48016 = n4464 & ~n48015;
  assign n48017 = ~n30806 & ~n47958;
  assign n48018 = ~n4464 & ~n48017;
  assign n48019 = ~n48016 & ~n48018;
  assign n48020 = ~n4463 & ~n48019;
  assign n48021 = ~n47992 & ~n48020;
  assign n48022 = ~n4462 & ~n48021;
  assign n48023 = ~n47964 & ~n48022;
  assign n48024 = n4461 & ~n48023;
  assign n48025 = ~n18434 & ~n45155;
  assign n48026 = i_RtoB_ACK0 & ~n48025;
  assign n48027 = ~n46034 & ~n47037;
  assign n48028 = ~i_RtoB_ACK0 & ~n48027;
  assign n48029 = ~n48026 & ~n48028;
  assign n48030 = ~controllable_DEQ & ~n48029;
  assign n48031 = ~n20981 & ~n48030;
  assign n48032 = i_FULL & ~n48031;
  assign n48033 = ~n46041 & ~n47037;
  assign n48034 = ~i_RtoB_ACK0 & ~n48033;
  assign n48035 = ~n48026 & ~n48034;
  assign n48036 = ~controllable_DEQ & ~n48035;
  assign n48037 = ~n20981 & ~n48036;
  assign n48038 = ~i_FULL & ~n48037;
  assign n48039 = ~n48032 & ~n48038;
  assign n48040 = i_nEMPTY & ~n48039;
  assign n48041 = ~n18428 & ~n45187;
  assign n48042 = i_RtoB_ACK0 & ~n48041;
  assign n48043 = ~n46050 & ~n47050;
  assign n48044 = ~i_RtoB_ACK0 & ~n48043;
  assign n48045 = ~n48042 & ~n48044;
  assign n48046 = ~controllable_DEQ & ~n48045;
  assign n48047 = ~n20993 & ~n48046;
  assign n48048 = i_FULL & ~n48047;
  assign n48049 = ~n46057 & ~n47063;
  assign n48050 = ~i_RtoB_ACK0 & ~n48049;
  assign n48051 = ~n48042 & ~n48050;
  assign n48052 = ~controllable_DEQ & ~n48051;
  assign n48053 = ~n21003 & ~n48052;
  assign n48054 = ~i_FULL & ~n48053;
  assign n48055 = ~n48048 & ~n48054;
  assign n48056 = ~i_nEMPTY & ~n48055;
  assign n48057 = ~n48040 & ~n48056;
  assign n48058 = controllable_BtoS_ACK0 & ~n48057;
  assign n48059 = ~n18462 & ~n45219;
  assign n48060 = i_RtoB_ACK0 & ~n48059;
  assign n48061 = ~n46068 & ~n47080;
  assign n48062 = ~i_RtoB_ACK0 & ~n48061;
  assign n48063 = ~n48060 & ~n48062;
  assign n48064 = ~controllable_DEQ & ~n48063;
  assign n48065 = ~n29641 & ~n48064;
  assign n48066 = i_FULL & ~n48065;
  assign n48067 = ~n46075 & ~n47080;
  assign n48068 = ~i_RtoB_ACK0 & ~n48067;
  assign n48069 = ~n48060 & ~n48068;
  assign n48070 = ~controllable_DEQ & ~n48069;
  assign n48071 = ~n29641 & ~n48070;
  assign n48072 = ~i_FULL & ~n48071;
  assign n48073 = ~n48066 & ~n48072;
  assign n48074 = i_nEMPTY & ~n48073;
  assign n48075 = ~n18456 & ~n45251;
  assign n48076 = i_RtoB_ACK0 & ~n48075;
  assign n48077 = ~n46084 & ~n47093;
  assign n48078 = ~i_RtoB_ACK0 & ~n48077;
  assign n48079 = ~n48076 & ~n48078;
  assign n48080 = ~controllable_DEQ & ~n48079;
  assign n48081 = ~n29653 & ~n48080;
  assign n48082 = i_FULL & ~n48081;
  assign n48083 = ~n46091 & ~n47106;
  assign n48084 = ~i_RtoB_ACK0 & ~n48083;
  assign n48085 = ~n48076 & ~n48084;
  assign n48086 = ~controllable_DEQ & ~n48085;
  assign n48087 = ~n29663 & ~n48086;
  assign n48088 = ~i_FULL & ~n48087;
  assign n48089 = ~n48082 & ~n48088;
  assign n48090 = ~i_nEMPTY & ~n48089;
  assign n48091 = ~n48074 & ~n48090;
  assign n48092 = ~controllable_BtoS_ACK0 & ~n48091;
  assign n48093 = ~n48058 & ~n48092;
  assign n48094 = n4465 & ~n48093;
  assign n48095 = ~n29641 & ~n31054;
  assign n48096 = i_FULL & ~n48095;
  assign n48097 = ~n31062 & ~n48096;
  assign n48098 = i_nEMPTY & ~n48097;
  assign n48099 = ~n31078 & ~n48098;
  assign n48100 = ~controllable_BtoS_ACK0 & ~n48099;
  assign n48101 = ~n21013 & ~n48100;
  assign n48102 = ~n4465 & ~n48101;
  assign n48103 = ~n48094 & ~n48102;
  assign n48104 = i_StoB_REQ10 & ~n48103;
  assign n48105 = ~n45382 & ~n47128;
  assign n48106 = i_RtoB_ACK0 & ~n48105;
  assign n48107 = ~n46106 & ~n47134;
  assign n48108 = ~i_RtoB_ACK0 & ~n48107;
  assign n48109 = ~n48106 & ~n48108;
  assign n48110 = ~controllable_DEQ & ~n48109;
  assign n48111 = ~n23093 & ~n48110;
  assign n48112 = i_FULL & ~n48111;
  assign n48113 = ~n46113 & ~n47134;
  assign n48114 = ~i_RtoB_ACK0 & ~n48113;
  assign n48115 = ~n48106 & ~n48114;
  assign n48116 = ~controllable_DEQ & ~n48115;
  assign n48117 = ~n23093 & ~n48116;
  assign n48118 = ~i_FULL & ~n48117;
  assign n48119 = ~n48112 & ~n48118;
  assign n48120 = i_nEMPTY & ~n48119;
  assign n48121 = ~n45422 & ~n47147;
  assign n48122 = i_RtoB_ACK0 & ~n48121;
  assign n48123 = ~n46122 & ~n47153;
  assign n48124 = ~i_RtoB_ACK0 & ~n48123;
  assign n48125 = ~n48122 & ~n48124;
  assign n48126 = ~controllable_DEQ & ~n48125;
  assign n48127 = ~n23105 & ~n48126;
  assign n48128 = i_FULL & ~n48127;
  assign n48129 = ~n45422 & ~n47166;
  assign n48130 = i_RtoB_ACK0 & ~n48129;
  assign n48131 = ~n46132 & ~n47172;
  assign n48132 = ~i_RtoB_ACK0 & ~n48131;
  assign n48133 = ~n48130 & ~n48132;
  assign n48134 = ~controllable_DEQ & ~n48133;
  assign n48135 = ~n23117 & ~n48134;
  assign n48136 = ~i_FULL & ~n48135;
  assign n48137 = ~n48128 & ~n48136;
  assign n48138 = ~i_nEMPTY & ~n48137;
  assign n48139 = ~n48120 & ~n48138;
  assign n48140 = controllable_BtoS_ACK0 & ~n48139;
  assign n48141 = ~n45467 & ~n47188;
  assign n48142 = i_RtoB_ACK0 & ~n48141;
  assign n48143 = ~n46143 & ~n47194;
  assign n48144 = ~i_RtoB_ACK0 & ~n48143;
  assign n48145 = ~n48142 & ~n48144;
  assign n48146 = ~controllable_DEQ & ~n48145;
  assign n48147 = ~n23133 & ~n48146;
  assign n48148 = i_FULL & ~n48147;
  assign n48149 = ~n46150 & ~n47194;
  assign n48150 = ~i_RtoB_ACK0 & ~n48149;
  assign n48151 = ~n48142 & ~n48150;
  assign n48152 = ~controllable_DEQ & ~n48151;
  assign n48153 = ~n23133 & ~n48152;
  assign n48154 = ~i_FULL & ~n48153;
  assign n48155 = ~n48148 & ~n48154;
  assign n48156 = i_nEMPTY & ~n48155;
  assign n48157 = ~n45507 & ~n47207;
  assign n48158 = i_RtoB_ACK0 & ~n48157;
  assign n48159 = ~n46159 & ~n47213;
  assign n48160 = ~i_RtoB_ACK0 & ~n48159;
  assign n48161 = ~n48158 & ~n48160;
  assign n48162 = ~controllable_DEQ & ~n48161;
  assign n48163 = ~n23145 & ~n48162;
  assign n48164 = i_FULL & ~n48163;
  assign n48165 = ~n45507 & ~n47226;
  assign n48166 = i_RtoB_ACK0 & ~n48165;
  assign n48167 = ~n46169 & ~n47232;
  assign n48168 = ~i_RtoB_ACK0 & ~n48167;
  assign n48169 = ~n48166 & ~n48168;
  assign n48170 = ~controllable_DEQ & ~n48169;
  assign n48171 = ~n23157 & ~n48170;
  assign n48172 = ~i_FULL & ~n48171;
  assign n48173 = ~n48164 & ~n48172;
  assign n48174 = ~i_nEMPTY & ~n48173;
  assign n48175 = ~n48156 & ~n48174;
  assign n48176 = ~controllable_BtoS_ACK0 & ~n48175;
  assign n48177 = ~n48140 & ~n48176;
  assign n48178 = n4465 & ~n48177;
  assign n48179 = ~n23133 & ~n31162;
  assign n48180 = i_FULL & ~n48179;
  assign n48181 = ~n31170 & ~n48180;
  assign n48182 = i_nEMPTY & ~n48181;
  assign n48183 = ~n31186 & ~n48182;
  assign n48184 = ~controllable_BtoS_ACK0 & ~n48183;
  assign n48185 = ~n23127 & ~n48184;
  assign n48186 = ~n4465 & ~n48185;
  assign n48187 = ~n48178 & ~n48186;
  assign n48188 = ~i_StoB_REQ10 & ~n48187;
  assign n48189 = ~n48104 & ~n48188;
  assign n48190 = controllable_BtoS_ACK10 & ~n48189;
  assign n48191 = ~n17058 & ~n45557;
  assign n48192 = i_RtoB_ACK0 & ~n48191;
  assign n48193 = controllable_BtoR_REQ0 & ~n47253;
  assign n48194 = ~n28594 & ~n48193;
  assign n48195 = ~i_RtoB_ACK0 & ~n48194;
  assign n48196 = ~n48192 & ~n48195;
  assign n48197 = ~controllable_DEQ & ~n48196;
  assign n48198 = ~n29844 & ~n48197;
  assign n48199 = i_FULL & ~n48198;
  assign n48200 = ~n46190 & ~n48193;
  assign n48201 = ~i_RtoB_ACK0 & ~n48200;
  assign n48202 = ~n48192 & ~n48201;
  assign n48203 = ~controllable_DEQ & ~n48202;
  assign n48204 = ~n29844 & ~n48203;
  assign n48205 = ~i_FULL & ~n48204;
  assign n48206 = ~n48199 & ~n48205;
  assign n48207 = i_nEMPTY & ~n48206;
  assign n48208 = ~n17068 & ~n45583;
  assign n48209 = i_RtoB_ACK0 & ~n48208;
  assign n48210 = controllable_BtoR_REQ0 & ~n47260;
  assign n48211 = ~n28610 & ~n48210;
  assign n48212 = ~i_RtoB_ACK0 & ~n48211;
  assign n48213 = ~n48209 & ~n48212;
  assign n48214 = ~controllable_DEQ & ~n48213;
  assign n48215 = ~n29858 & ~n48214;
  assign n48216 = i_FULL & ~n48215;
  assign n48217 = ~n45583 & ~n47269;
  assign n48218 = i_RtoB_ACK0 & ~n48217;
  assign n48219 = controllable_BtoR_REQ0 & ~n47272;
  assign n48220 = ~n46206 & ~n48219;
  assign n48221 = ~i_RtoB_ACK0 & ~n48220;
  assign n48222 = ~n48218 & ~n48221;
  assign n48223 = ~controllable_DEQ & ~n48222;
  assign n48224 = ~n29872 & ~n48223;
  assign n48225 = ~i_FULL & ~n48224;
  assign n48226 = ~n48216 & ~n48225;
  assign n48227 = ~i_nEMPTY & ~n48226;
  assign n48228 = ~n48207 & ~n48227;
  assign n48229 = controllable_BtoS_ACK0 & ~n48228;
  assign n48230 = ~n18530 & ~n45615;
  assign n48231 = i_RtoB_ACK0 & ~n48230;
  assign n48232 = controllable_BtoR_REQ0 & ~n47283;
  assign n48233 = ~n28069 & ~n48232;
  assign n48234 = ~i_RtoB_ACK0 & ~n48233;
  assign n48235 = ~n48231 & ~n48234;
  assign n48236 = ~controllable_DEQ & ~n48235;
  assign n48237 = ~n29900 & ~n48236;
  assign n48238 = i_FULL & ~n48237;
  assign n48239 = ~n46221 & ~n48232;
  assign n48240 = ~i_RtoB_ACK0 & ~n48239;
  assign n48241 = ~n48231 & ~n48240;
  assign n48242 = ~controllable_DEQ & ~n48241;
  assign n48243 = ~n29900 & ~n48242;
  assign n48244 = ~i_FULL & ~n48243;
  assign n48245 = ~n48238 & ~n48244;
  assign n48246 = i_nEMPTY & ~n48245;
  assign n48247 = ~n18548 & ~n45641;
  assign n48248 = i_RtoB_ACK0 & ~n48247;
  assign n48249 = controllable_BtoR_REQ0 & ~n47290;
  assign n48250 = ~n28085 & ~n48249;
  assign n48251 = ~i_RtoB_ACK0 & ~n48250;
  assign n48252 = ~n48248 & ~n48251;
  assign n48253 = ~controllable_DEQ & ~n48252;
  assign n48254 = ~n29914 & ~n48253;
  assign n48255 = i_FULL & ~n48254;
  assign n48256 = ~n45641 & ~n47299;
  assign n48257 = i_RtoB_ACK0 & ~n48256;
  assign n48258 = controllable_BtoR_REQ0 & ~n47302;
  assign n48259 = ~n46237 & ~n48258;
  assign n48260 = ~i_RtoB_ACK0 & ~n48259;
  assign n48261 = ~n48257 & ~n48260;
  assign n48262 = ~controllable_DEQ & ~n48261;
  assign n48263 = ~n29928 & ~n48262;
  assign n48264 = ~i_FULL & ~n48263;
  assign n48265 = ~n48255 & ~n48264;
  assign n48266 = ~i_nEMPTY & ~n48265;
  assign n48267 = ~n48246 & ~n48266;
  assign n48268 = ~controllable_BtoS_ACK0 & ~n48267;
  assign n48269 = ~n48229 & ~n48268;
  assign n48270 = n4465 & ~n48269;
  assign n48271 = ~n29900 & ~n31268;
  assign n48272 = i_FULL & ~n48271;
  assign n48273 = ~n31276 & ~n48272;
  assign n48274 = i_nEMPTY & ~n48273;
  assign n48275 = ~n31289 & ~n48274;
  assign n48276 = ~controllable_BtoS_ACK0 & ~n48275;
  assign n48277 = ~n29958 & ~n48276;
  assign n48278 = ~n4465 & ~n48277;
  assign n48279 = ~n48270 & ~n48278;
  assign n48280 = i_StoB_REQ10 & ~n48279;
  assign n48281 = ~n48188 & ~n48280;
  assign n48282 = ~controllable_BtoS_ACK10 & ~n48281;
  assign n48283 = ~n48190 & ~n48282;
  assign n48284 = n4464 & ~n48283;
  assign n48285 = ~n20981 & ~n31307;
  assign n48286 = i_FULL & ~n48285;
  assign n48287 = ~n31315 & ~n48286;
  assign n48288 = i_nEMPTY & ~n48287;
  assign n48289 = ~n31331 & ~n48288;
  assign n48290 = controllable_BtoS_ACK0 & ~n48289;
  assign n48291 = ~n29641 & ~n31341;
  assign n48292 = i_FULL & ~n48291;
  assign n48293 = ~n31349 & ~n48292;
  assign n48294 = i_nEMPTY & ~n48293;
  assign n48295 = ~n31365 & ~n48294;
  assign n48296 = ~controllable_BtoS_ACK0 & ~n48295;
  assign n48297 = ~n48290 & ~n48296;
  assign n48298 = n4465 & ~n48297;
  assign n48299 = ~n21013 & ~n48296;
  assign n48300 = ~n4465 & ~n48299;
  assign n48301 = ~n48298 & ~n48300;
  assign n48302 = i_StoB_REQ10 & ~n48301;
  assign n48303 = ~n23093 & ~n31381;
  assign n48304 = i_FULL & ~n48303;
  assign n48305 = ~n31389 & ~n48304;
  assign n48306 = i_nEMPTY & ~n48305;
  assign n48307 = ~n31405 & ~n48306;
  assign n48308 = controllable_BtoS_ACK0 & ~n48307;
  assign n48309 = ~n23133 & ~n31415;
  assign n48310 = i_FULL & ~n48309;
  assign n48311 = ~n31423 & ~n48310;
  assign n48312 = i_nEMPTY & ~n48311;
  assign n48313 = ~n31439 & ~n48312;
  assign n48314 = ~controllable_BtoS_ACK0 & ~n48313;
  assign n48315 = ~n48308 & ~n48314;
  assign n48316 = n4465 & ~n48315;
  assign n48317 = ~n23127 & ~n48314;
  assign n48318 = ~n4465 & ~n48317;
  assign n48319 = ~n48316 & ~n48318;
  assign n48320 = ~i_StoB_REQ10 & ~n48319;
  assign n48321 = ~n48302 & ~n48320;
  assign n48322 = controllable_BtoS_ACK10 & ~n48321;
  assign n48323 = ~n29844 & ~n31457;
  assign n48324 = i_FULL & ~n48323;
  assign n48325 = ~n31465 & ~n48324;
  assign n48326 = i_nEMPTY & ~n48325;
  assign n48327 = ~n31478 & ~n48326;
  assign n48328 = controllable_BtoS_ACK0 & ~n48327;
  assign n48329 = ~n29900 & ~n31488;
  assign n48330 = i_FULL & ~n48329;
  assign n48331 = ~n31496 & ~n48330;
  assign n48332 = i_nEMPTY & ~n48331;
  assign n48333 = ~n31509 & ~n48332;
  assign n48334 = ~controllable_BtoS_ACK0 & ~n48333;
  assign n48335 = ~n48328 & ~n48334;
  assign n48336 = n4465 & ~n48335;
  assign n48337 = ~n29958 & ~n48334;
  assign n48338 = ~n4465 & ~n48337;
  assign n48339 = ~n48336 & ~n48338;
  assign n48340 = i_StoB_REQ10 & ~n48339;
  assign n48341 = ~n48320 & ~n48340;
  assign n48342 = ~controllable_BtoS_ACK10 & ~n48341;
  assign n48343 = ~n48322 & ~n48342;
  assign n48344 = ~n4464 & ~n48343;
  assign n48345 = ~n48284 & ~n48344;
  assign n48346 = n4463 & ~n48345;
  assign n48347 = ~n45753 & ~n47037;
  assign n48348 = ~i_RtoB_ACK0 & ~n48347;
  assign n48349 = ~n47648 & ~n48348;
  assign n48350 = ~controllable_DEQ & ~n48349;
  assign n48351 = ~n20981 & ~n48350;
  assign n48352 = i_nEMPTY & ~n48351;
  assign n48353 = ~n45765 & ~n47050;
  assign n48354 = ~i_RtoB_ACK0 & ~n48353;
  assign n48355 = ~n47664 & ~n48354;
  assign n48356 = ~controllable_DEQ & ~n48355;
  assign n48357 = ~n20993 & ~n48356;
  assign n48358 = i_FULL & ~n48357;
  assign n48359 = ~n45775 & ~n47063;
  assign n48360 = ~i_RtoB_ACK0 & ~n48359;
  assign n48361 = ~n47664 & ~n48360;
  assign n48362 = ~controllable_DEQ & ~n48361;
  assign n48363 = ~n21003 & ~n48362;
  assign n48364 = ~i_FULL & ~n48363;
  assign n48365 = ~n48358 & ~n48364;
  assign n48366 = ~i_nEMPTY & ~n48365;
  assign n48367 = ~n48352 & ~n48366;
  assign n48368 = controllable_BtoS_ACK0 & ~n48367;
  assign n48369 = ~n45791 & ~n47080;
  assign n48370 = ~i_RtoB_ACK0 & ~n48369;
  assign n48371 = ~n47682 & ~n48370;
  assign n48372 = ~controllable_DEQ & ~n48371;
  assign n48373 = ~n29641 & ~n48372;
  assign n48374 = i_nEMPTY & ~n48373;
  assign n48375 = ~n45803 & ~n47093;
  assign n48376 = ~i_RtoB_ACK0 & ~n48375;
  assign n48377 = ~n47698 & ~n48376;
  assign n48378 = ~controllable_DEQ & ~n48377;
  assign n48379 = ~n29653 & ~n48378;
  assign n48380 = i_FULL & ~n48379;
  assign n48381 = ~n45813 & ~n47106;
  assign n48382 = ~i_RtoB_ACK0 & ~n48381;
  assign n48383 = ~n47698 & ~n48382;
  assign n48384 = ~controllable_DEQ & ~n48383;
  assign n48385 = ~n29663 & ~n48384;
  assign n48386 = ~i_FULL & ~n48385;
  assign n48387 = ~n48380 & ~n48386;
  assign n48388 = ~i_nEMPTY & ~n48387;
  assign n48389 = ~n48374 & ~n48388;
  assign n48390 = ~controllable_BtoS_ACK0 & ~n48389;
  assign n48391 = ~n48368 & ~n48390;
  assign n48392 = n4465 & ~n48391;
  assign n48393 = ~n4465 & ~n30803;
  assign n48394 = ~n48392 & ~n48393;
  assign n48395 = i_StoB_REQ10 & ~n48394;
  assign n48396 = ~n45830 & ~n47128;
  assign n48397 = i_RtoB_ACK0 & ~n48396;
  assign n48398 = ~n45834 & ~n47134;
  assign n48399 = ~i_RtoB_ACK0 & ~n48398;
  assign n48400 = ~n48397 & ~n48399;
  assign n48401 = ~controllable_DEQ & ~n48400;
  assign n48402 = ~n23093 & ~n48401;
  assign n48403 = i_nEMPTY & ~n48402;
  assign n48404 = ~n45842 & ~n47147;
  assign n48405 = i_RtoB_ACK0 & ~n48404;
  assign n48406 = ~n45846 & ~n47153;
  assign n48407 = ~i_RtoB_ACK0 & ~n48406;
  assign n48408 = ~n48405 & ~n48407;
  assign n48409 = ~controllable_DEQ & ~n48408;
  assign n48410 = ~n23105 & ~n48409;
  assign n48411 = i_FULL & ~n48410;
  assign n48412 = ~n45842 & ~n47166;
  assign n48413 = i_RtoB_ACK0 & ~n48412;
  assign n48414 = ~n45862 & ~n47172;
  assign n48415 = ~i_RtoB_ACK0 & ~n48414;
  assign n48416 = ~n48413 & ~n48415;
  assign n48417 = ~controllable_DEQ & ~n48416;
  assign n48418 = ~n23117 & ~n48417;
  assign n48419 = ~i_FULL & ~n48418;
  assign n48420 = ~n48411 & ~n48419;
  assign n48421 = ~i_nEMPTY & ~n48420;
  assign n48422 = ~n48403 & ~n48421;
  assign n48423 = controllable_BtoS_ACK0 & ~n48422;
  assign n48424 = ~n45874 & ~n47188;
  assign n48425 = i_RtoB_ACK0 & ~n48424;
  assign n48426 = ~n45878 & ~n47194;
  assign n48427 = ~i_RtoB_ACK0 & ~n48426;
  assign n48428 = ~n48425 & ~n48427;
  assign n48429 = ~controllable_DEQ & ~n48428;
  assign n48430 = ~n23133 & ~n48429;
  assign n48431 = i_nEMPTY & ~n48430;
  assign n48432 = ~n45886 & ~n47207;
  assign n48433 = i_RtoB_ACK0 & ~n48432;
  assign n48434 = ~n45890 & ~n47213;
  assign n48435 = ~i_RtoB_ACK0 & ~n48434;
  assign n48436 = ~n48433 & ~n48435;
  assign n48437 = ~controllable_DEQ & ~n48436;
  assign n48438 = ~n23145 & ~n48437;
  assign n48439 = i_FULL & ~n48438;
  assign n48440 = ~n45886 & ~n47226;
  assign n48441 = i_RtoB_ACK0 & ~n48440;
  assign n48442 = ~n45906 & ~n47232;
  assign n48443 = ~i_RtoB_ACK0 & ~n48442;
  assign n48444 = ~n48441 & ~n48443;
  assign n48445 = ~controllable_DEQ & ~n48444;
  assign n48446 = ~n23157 & ~n48445;
  assign n48447 = ~i_FULL & ~n48446;
  assign n48448 = ~n48439 & ~n48447;
  assign n48449 = ~i_nEMPTY & ~n48448;
  assign n48450 = ~n48431 & ~n48449;
  assign n48451 = ~controllable_BtoS_ACK0 & ~n48450;
  assign n48452 = ~n48423 & ~n48451;
  assign n48453 = n4465 & ~n48452;
  assign n48454 = ~n4465 & ~n23168;
  assign n48455 = ~n48453 & ~n48454;
  assign n48456 = ~i_StoB_REQ10 & ~n48455;
  assign n48457 = ~n48395 & ~n48456;
  assign n48458 = controllable_BtoS_ACK10 & ~n48457;
  assign n48459 = ~n45925 & ~n48193;
  assign n48460 = ~i_RtoB_ACK0 & ~n48459;
  assign n48461 = ~n29832 & ~n48460;
  assign n48462 = ~controllable_DEQ & ~n48461;
  assign n48463 = ~n29844 & ~n48462;
  assign n48464 = i_nEMPTY & ~n48463;
  assign n48465 = ~n45933 & ~n48210;
  assign n48466 = ~i_RtoB_ACK0 & ~n48465;
  assign n48467 = ~n29860 & ~n48466;
  assign n48468 = ~controllable_DEQ & ~n48467;
  assign n48469 = ~n29858 & ~n48468;
  assign n48470 = i_FULL & ~n48469;
  assign n48471 = ~n28112 & ~n47269;
  assign n48472 = i_RtoB_ACK0 & ~n48471;
  assign n48473 = ~n45945 & ~n48219;
  assign n48474 = ~i_RtoB_ACK0 & ~n48473;
  assign n48475 = ~n48472 & ~n48474;
  assign n48476 = ~controllable_DEQ & ~n48475;
  assign n48477 = ~n29872 & ~n48476;
  assign n48478 = ~i_FULL & ~n48477;
  assign n48479 = ~n48470 & ~n48478;
  assign n48480 = ~i_nEMPTY & ~n48479;
  assign n48481 = ~n48464 & ~n48480;
  assign n48482 = controllable_BtoS_ACK0 & ~n48481;
  assign n48483 = ~n45957 & ~n48232;
  assign n48484 = ~i_RtoB_ACK0 & ~n48483;
  assign n48485 = ~n29888 & ~n48484;
  assign n48486 = ~controllable_DEQ & ~n48485;
  assign n48487 = ~n29900 & ~n48486;
  assign n48488 = i_nEMPTY & ~n48487;
  assign n48489 = ~n45965 & ~n48249;
  assign n48490 = ~i_RtoB_ACK0 & ~n48489;
  assign n48491 = ~n29916 & ~n48490;
  assign n48492 = ~controllable_DEQ & ~n48491;
  assign n48493 = ~n29914 & ~n48492;
  assign n48494 = i_FULL & ~n48493;
  assign n48495 = ~n28173 & ~n47299;
  assign n48496 = i_RtoB_ACK0 & ~n48495;
  assign n48497 = ~n45977 & ~n48258;
  assign n48498 = ~i_RtoB_ACK0 & ~n48497;
  assign n48499 = ~n48496 & ~n48498;
  assign n48500 = ~controllable_DEQ & ~n48499;
  assign n48501 = ~n29928 & ~n48500;
  assign n48502 = ~i_FULL & ~n48501;
  assign n48503 = ~n48494 & ~n48502;
  assign n48504 = ~i_nEMPTY & ~n48503;
  assign n48505 = ~n48488 & ~n48504;
  assign n48506 = ~controllable_BtoS_ACK0 & ~n48505;
  assign n48507 = ~n48482 & ~n48506;
  assign n48508 = n4465 & ~n48507;
  assign n48509 = ~n4465 & ~n31543;
  assign n48510 = ~n48508 & ~n48509;
  assign n48511 = i_StoB_REQ10 & ~n48510;
  assign n48512 = ~n48456 & ~n48511;
  assign n48513 = ~controllable_BtoS_ACK10 & ~n48512;
  assign n48514 = ~n48458 & ~n48513;
  assign n48515 = n4464 & ~n48514;
  assign n48516 = ~n4464 & ~n31547;
  assign n48517 = ~n48515 & ~n48516;
  assign n48518 = ~n4463 & ~n48517;
  assign n48519 = ~n48346 & ~n48518;
  assign n48520 = n4462 & ~n48519;
  assign n48521 = ~n29844 & ~n31558;
  assign n48522 = i_FULL & ~n48521;
  assign n48523 = ~n31566 & ~n48522;
  assign n48524 = i_nEMPTY & ~n48523;
  assign n48525 = ~n31579 & ~n48524;
  assign n48526 = controllable_BtoS_ACK0 & ~n48525;
  assign n48527 = ~n48276 & ~n48526;
  assign n48528 = n4465 & ~n48527;
  assign n48529 = ~n48278 & ~n48528;
  assign n48530 = i_StoB_REQ10 & ~n48529;
  assign n48531 = ~n23093 & ~n31593;
  assign n48532 = i_FULL & ~n48531;
  assign n48533 = ~n31601 & ~n48532;
  assign n48534 = i_nEMPTY & ~n48533;
  assign n48535 = ~n31617 & ~n48534;
  assign n48536 = controllable_BtoS_ACK0 & ~n48535;
  assign n48537 = ~n48184 & ~n48536;
  assign n48538 = n4465 & ~n48537;
  assign n48539 = ~n48186 & ~n48538;
  assign n48540 = ~i_StoB_REQ10 & ~n48539;
  assign n48541 = ~n48530 & ~n48540;
  assign n48542 = ~controllable_BtoS_ACK10 & ~n48541;
  assign n48543 = ~n30806 & ~n48542;
  assign n48544 = n4464 & ~n48543;
  assign n48545 = ~n30806 & ~n48342;
  assign n48546 = ~n4464 & ~n48545;
  assign n48547 = ~n48544 & ~n48546;
  assign n48548 = n4463 & ~n48547;
  assign n48549 = ~n31548 & ~n48548;
  assign n48550 = ~n4462 & ~n48549;
  assign n48551 = ~n48520 & ~n48550;
  assign n48552 = ~n4461 & ~n48551;
  assign n48553 = ~n48024 & ~n48552;
  assign n48554 = ~n4459 & ~n48553;
  assign n48555 = controllable_BtoR_REQ1 & ~n45752;
  assign n48556 = ~n45158 & ~n48555;
  assign n48557 = ~controllable_BtoR_REQ0 & ~n48556;
  assign n48558 = ~n46272 & ~n48557;
  assign n48559 = ~i_RtoB_ACK0 & ~n48558;
  assign n48560 = ~n47648 & ~n48559;
  assign n48561 = ~controllable_DEQ & ~n48560;
  assign n48562 = ~n20981 & ~n48561;
  assign n48563 = i_FULL & ~n48562;
  assign n48564 = ~n45169 & ~n48555;
  assign n48565 = ~controllable_BtoR_REQ0 & ~n48564;
  assign n48566 = ~n46284 & ~n48565;
  assign n48567 = ~i_RtoB_ACK0 & ~n48566;
  assign n48568 = ~n47648 & ~n48567;
  assign n48569 = ~controllable_DEQ & ~n48568;
  assign n48570 = ~n20981 & ~n48569;
  assign n48571 = ~i_FULL & ~n48570;
  assign n48572 = ~n48563 & ~n48571;
  assign n48573 = i_nEMPTY & ~n48572;
  assign n48574 = controllable_BtoR_REQ1 & ~n45764;
  assign n48575 = ~n45190 & ~n48574;
  assign n48576 = ~controllable_BtoR_REQ0 & ~n48575;
  assign n48577 = ~n46303 & ~n48576;
  assign n48578 = ~i_RtoB_ACK0 & ~n48577;
  assign n48579 = ~n47664 & ~n48578;
  assign n48580 = ~controllable_DEQ & ~n48579;
  assign n48581 = ~n20993 & ~n48580;
  assign n48582 = i_FULL & ~n48581;
  assign n48583 = controllable_BtoR_REQ1 & ~n45774;
  assign n48584 = ~n45201 & ~n48583;
  assign n48585 = ~controllable_BtoR_REQ0 & ~n48584;
  assign n48586 = ~n46315 & ~n48585;
  assign n48587 = ~i_RtoB_ACK0 & ~n48586;
  assign n48588 = ~n47664 & ~n48587;
  assign n48589 = ~controllable_DEQ & ~n48588;
  assign n48590 = ~n21003 & ~n48589;
  assign n48591 = ~i_FULL & ~n48590;
  assign n48592 = ~n48582 & ~n48591;
  assign n48593 = ~i_nEMPTY & ~n48592;
  assign n48594 = ~n48573 & ~n48593;
  assign n48595 = controllable_BtoS_ACK0 & ~n48594;
  assign n48596 = controllable_BtoR_REQ1 & ~n45790;
  assign n48597 = ~n45222 & ~n48596;
  assign n48598 = ~controllable_BtoR_REQ0 & ~n48597;
  assign n48599 = ~n46336 & ~n48598;
  assign n48600 = ~i_RtoB_ACK0 & ~n48599;
  assign n48601 = ~n47682 & ~n48600;
  assign n48602 = ~controllable_DEQ & ~n48601;
  assign n48603 = ~n29641 & ~n48602;
  assign n48604 = i_FULL & ~n48603;
  assign n48605 = ~n45233 & ~n48596;
  assign n48606 = ~controllable_BtoR_REQ0 & ~n48605;
  assign n48607 = ~n46348 & ~n48606;
  assign n48608 = ~i_RtoB_ACK0 & ~n48607;
  assign n48609 = ~n47682 & ~n48608;
  assign n48610 = ~controllable_DEQ & ~n48609;
  assign n48611 = ~n29641 & ~n48610;
  assign n48612 = ~i_FULL & ~n48611;
  assign n48613 = ~n48604 & ~n48612;
  assign n48614 = i_nEMPTY & ~n48613;
  assign n48615 = controllable_BtoR_REQ1 & ~n45802;
  assign n48616 = ~n45254 & ~n48615;
  assign n48617 = ~controllable_BtoR_REQ0 & ~n48616;
  assign n48618 = ~n46367 & ~n48617;
  assign n48619 = ~i_RtoB_ACK0 & ~n48618;
  assign n48620 = ~n47698 & ~n48619;
  assign n48621 = ~controllable_DEQ & ~n48620;
  assign n48622 = ~n29653 & ~n48621;
  assign n48623 = i_FULL & ~n48622;
  assign n48624 = controllable_BtoR_REQ1 & ~n45812;
  assign n48625 = ~n45265 & ~n48624;
  assign n48626 = ~controllable_BtoR_REQ0 & ~n48625;
  assign n48627 = ~n46379 & ~n48626;
  assign n48628 = ~i_RtoB_ACK0 & ~n48627;
  assign n48629 = ~n47698 & ~n48628;
  assign n48630 = ~controllable_DEQ & ~n48629;
  assign n48631 = ~n29663 & ~n48630;
  assign n48632 = ~i_FULL & ~n48631;
  assign n48633 = ~n48623 & ~n48632;
  assign n48634 = ~i_nEMPTY & ~n48633;
  assign n48635 = ~n48614 & ~n48634;
  assign n48636 = ~controllable_BtoS_ACK0 & ~n48635;
  assign n48637 = ~n48595 & ~n48636;
  assign n48638 = n4465 & ~n48637;
  assign n48639 = ~n29641 & ~n31743;
  assign n48640 = i_FULL & ~n48639;
  assign n48641 = ~n31753 & ~n48640;
  assign n48642 = i_nEMPTY & ~n48641;
  assign n48643 = ~n31773 & ~n48642;
  assign n48644 = ~controllable_BtoS_ACK0 & ~n48643;
  assign n48645 = ~n21013 & ~n48644;
  assign n48646 = ~n4465 & ~n48645;
  assign n48647 = ~n48638 & ~n48646;
  assign n48648 = i_StoB_REQ10 & ~n48647;
  assign n48649 = controllable_BtoR_REQ1 & ~n45833;
  assign n48650 = ~n45388 & ~n48649;
  assign n48651 = ~controllable_BtoR_REQ0 & ~n48650;
  assign n48652 = ~n46416 & ~n48651;
  assign n48653 = ~i_RtoB_ACK0 & ~n48652;
  assign n48654 = ~n47728 & ~n48653;
  assign n48655 = ~controllable_DEQ & ~n48654;
  assign n48656 = ~n23093 & ~n48655;
  assign n48657 = i_FULL & ~n48656;
  assign n48658 = ~n45399 & ~n48649;
  assign n48659 = ~controllable_BtoR_REQ0 & ~n48658;
  assign n48660 = ~n46428 & ~n48659;
  assign n48661 = ~i_RtoB_ACK0 & ~n48660;
  assign n48662 = ~n47728 & ~n48661;
  assign n48663 = ~controllable_DEQ & ~n48662;
  assign n48664 = ~n23093 & ~n48663;
  assign n48665 = ~i_FULL & ~n48664;
  assign n48666 = ~n48657 & ~n48665;
  assign n48667 = i_nEMPTY & ~n48666;
  assign n48668 = controllable_BtoR_REQ1 & ~n45845;
  assign n48669 = ~n45428 & ~n48668;
  assign n48670 = ~controllable_BtoR_REQ0 & ~n48669;
  assign n48671 = ~n46451 & ~n48670;
  assign n48672 = ~i_RtoB_ACK0 & ~n48671;
  assign n48673 = ~n47744 & ~n48672;
  assign n48674 = ~controllable_DEQ & ~n48673;
  assign n48675 = ~n23105 & ~n48674;
  assign n48676 = i_FULL & ~n48675;
  assign n48677 = ~n45442 & ~n45858;
  assign n48678 = ~controllable_BtoR_REQ0 & ~n48677;
  assign n48679 = ~n46470 & ~n48678;
  assign n48680 = ~i_RtoB_ACK0 & ~n48679;
  assign n48681 = ~n47752 & ~n48680;
  assign n48682 = ~controllable_DEQ & ~n48681;
  assign n48683 = ~n23117 & ~n48682;
  assign n48684 = ~i_FULL & ~n48683;
  assign n48685 = ~n48676 & ~n48684;
  assign n48686 = ~i_nEMPTY & ~n48685;
  assign n48687 = ~n48667 & ~n48686;
  assign n48688 = controllable_BtoS_ACK0 & ~n48687;
  assign n48689 = controllable_BtoR_REQ1 & ~n45877;
  assign n48690 = ~n45473 & ~n48689;
  assign n48691 = ~controllable_BtoR_REQ0 & ~n48690;
  assign n48692 = ~n46495 & ~n48691;
  assign n48693 = ~i_RtoB_ACK0 & ~n48692;
  assign n48694 = ~n47764 & ~n48693;
  assign n48695 = ~controllable_DEQ & ~n48694;
  assign n48696 = ~n23133 & ~n48695;
  assign n48697 = i_FULL & ~n48696;
  assign n48698 = ~n45484 & ~n48689;
  assign n48699 = ~controllable_BtoR_REQ0 & ~n48698;
  assign n48700 = ~n46507 & ~n48699;
  assign n48701 = ~i_RtoB_ACK0 & ~n48700;
  assign n48702 = ~n47764 & ~n48701;
  assign n48703 = ~controllable_DEQ & ~n48702;
  assign n48704 = ~n23133 & ~n48703;
  assign n48705 = ~i_FULL & ~n48704;
  assign n48706 = ~n48697 & ~n48705;
  assign n48707 = i_nEMPTY & ~n48706;
  assign n48708 = controllable_BtoR_REQ1 & ~n45889;
  assign n48709 = ~n45513 & ~n48708;
  assign n48710 = ~controllable_BtoR_REQ0 & ~n48709;
  assign n48711 = ~n46530 & ~n48710;
  assign n48712 = ~i_RtoB_ACK0 & ~n48711;
  assign n48713 = ~n47780 & ~n48712;
  assign n48714 = ~controllable_DEQ & ~n48713;
  assign n48715 = ~n23145 & ~n48714;
  assign n48716 = i_FULL & ~n48715;
  assign n48717 = ~n45527 & ~n45902;
  assign n48718 = ~controllable_BtoR_REQ0 & ~n48717;
  assign n48719 = ~n46549 & ~n48718;
  assign n48720 = ~i_RtoB_ACK0 & ~n48719;
  assign n48721 = ~n47788 & ~n48720;
  assign n48722 = ~controllable_DEQ & ~n48721;
  assign n48723 = ~n23157 & ~n48722;
  assign n48724 = ~i_FULL & ~n48723;
  assign n48725 = ~n48716 & ~n48724;
  assign n48726 = ~i_nEMPTY & ~n48725;
  assign n48727 = ~n48707 & ~n48726;
  assign n48728 = ~controllable_BtoS_ACK0 & ~n48727;
  assign n48729 = ~n48688 & ~n48728;
  assign n48730 = n4465 & ~n48729;
  assign n48731 = ~n23133 & ~n31885;
  assign n48732 = i_FULL & ~n48731;
  assign n48733 = ~n31895 & ~n48732;
  assign n48734 = i_nEMPTY & ~n48733;
  assign n48735 = ~n31915 & ~n48734;
  assign n48736 = ~controllable_BtoS_ACK0 & ~n48735;
  assign n48737 = ~n23127 & ~n48736;
  assign n48738 = ~n4465 & ~n48737;
  assign n48739 = ~n48730 & ~n48738;
  assign n48740 = ~i_StoB_REQ10 & ~n48739;
  assign n48741 = ~n48648 & ~n48740;
  assign n48742 = controllable_BtoS_ACK10 & ~n48741;
  assign n48743 = controllable_BtoR_REQ1 & ~n45924;
  assign n48744 = ~n20377 & ~n48743;
  assign n48745 = ~controllable_BtoR_REQ0 & ~n48744;
  assign n48746 = ~n46581 & ~n48745;
  assign n48747 = ~i_RtoB_ACK0 & ~n48746;
  assign n48748 = ~n47814 & ~n48747;
  assign n48749 = ~controllable_DEQ & ~n48748;
  assign n48750 = ~n29844 & ~n48749;
  assign n48751 = i_FULL & ~n48750;
  assign n48752 = ~n45569 & ~n48743;
  assign n48753 = ~controllable_BtoR_REQ0 & ~n48752;
  assign n48754 = ~n46588 & ~n48753;
  assign n48755 = ~i_RtoB_ACK0 & ~n48754;
  assign n48756 = ~n47814 & ~n48755;
  assign n48757 = ~controllable_DEQ & ~n48756;
  assign n48758 = ~n29844 & ~n48757;
  assign n48759 = ~i_FULL & ~n48758;
  assign n48760 = ~n48751 & ~n48759;
  assign n48761 = i_nEMPTY & ~n48760;
  assign n48762 = controllable_BtoR_REQ1 & ~n45932;
  assign n48763 = ~n20411 & ~n48762;
  assign n48764 = ~controllable_BtoR_REQ0 & ~n48763;
  assign n48765 = ~n46604 & ~n48764;
  assign n48766 = ~i_RtoB_ACK0 & ~n48765;
  assign n48767 = ~n47830 & ~n48766;
  assign n48768 = ~controllable_DEQ & ~n48767;
  assign n48769 = ~n29858 & ~n48768;
  assign n48770 = i_FULL & ~n48769;
  assign n48771 = ~n45599 & ~n45941;
  assign n48772 = ~controllable_BtoR_REQ0 & ~n48771;
  assign n48773 = ~n46618 & ~n48772;
  assign n48774 = ~i_RtoB_ACK0 & ~n48773;
  assign n48775 = ~n47838 & ~n48774;
  assign n48776 = ~controllable_DEQ & ~n48775;
  assign n48777 = ~n29872 & ~n48776;
  assign n48778 = ~i_FULL & ~n48777;
  assign n48779 = ~n48770 & ~n48778;
  assign n48780 = ~i_nEMPTY & ~n48779;
  assign n48781 = ~n48761 & ~n48780;
  assign n48782 = controllable_BtoS_ACK0 & ~n48781;
  assign n48783 = controllable_BtoR_REQ1 & ~n45956;
  assign n48784 = ~n19321 & ~n48783;
  assign n48785 = ~controllable_BtoR_REQ0 & ~n48784;
  assign n48786 = ~n46636 & ~n48785;
  assign n48787 = ~i_RtoB_ACK0 & ~n48786;
  assign n48788 = ~n47850 & ~n48787;
  assign n48789 = ~controllable_DEQ & ~n48788;
  assign n48790 = ~n29900 & ~n48789;
  assign n48791 = i_FULL & ~n48790;
  assign n48792 = ~n45627 & ~n48783;
  assign n48793 = ~controllable_BtoR_REQ0 & ~n48792;
  assign n48794 = ~n46643 & ~n48793;
  assign n48795 = ~i_RtoB_ACK0 & ~n48794;
  assign n48796 = ~n47850 & ~n48795;
  assign n48797 = ~controllable_DEQ & ~n48796;
  assign n48798 = ~n29900 & ~n48797;
  assign n48799 = ~i_FULL & ~n48798;
  assign n48800 = ~n48791 & ~n48799;
  assign n48801 = i_nEMPTY & ~n48800;
  assign n48802 = controllable_BtoR_REQ1 & ~n45964;
  assign n48803 = ~n19351 & ~n48802;
  assign n48804 = ~controllable_BtoR_REQ0 & ~n48803;
  assign n48805 = ~n46659 & ~n48804;
  assign n48806 = ~i_RtoB_ACK0 & ~n48805;
  assign n48807 = ~n47866 & ~n48806;
  assign n48808 = ~controllable_DEQ & ~n48807;
  assign n48809 = ~n29914 & ~n48808;
  assign n48810 = i_FULL & ~n48809;
  assign n48811 = ~n45657 & ~n45973;
  assign n48812 = ~controllable_BtoR_REQ0 & ~n48811;
  assign n48813 = ~n46673 & ~n48812;
  assign n48814 = ~i_RtoB_ACK0 & ~n48813;
  assign n48815 = ~n47874 & ~n48814;
  assign n48816 = ~controllable_DEQ & ~n48815;
  assign n48817 = ~n29928 & ~n48816;
  assign n48818 = ~i_FULL & ~n48817;
  assign n48819 = ~n48810 & ~n48818;
  assign n48820 = ~i_nEMPTY & ~n48819;
  assign n48821 = ~n48801 & ~n48820;
  assign n48822 = ~controllable_BtoS_ACK0 & ~n48821;
  assign n48823 = ~n48782 & ~n48822;
  assign n48824 = n4465 & ~n48823;
  assign n48825 = ~n29900 & ~n32001;
  assign n48826 = i_FULL & ~n48825;
  assign n48827 = ~n32009 & ~n48826;
  assign n48828 = i_nEMPTY & ~n48827;
  assign n48829 = ~n32022 & ~n48828;
  assign n48830 = ~controllable_BtoS_ACK0 & ~n48829;
  assign n48831 = ~n29958 & ~n48830;
  assign n48832 = ~n4465 & ~n48831;
  assign n48833 = ~n48824 & ~n48832;
  assign n48834 = i_StoB_REQ10 & ~n48833;
  assign n48835 = ~n48740 & ~n48834;
  assign n48836 = ~controllable_BtoS_ACK10 & ~n48835;
  assign n48837 = ~n48742 & ~n48836;
  assign n48838 = n4464 & ~n48837;
  assign n48839 = ~n20981 & ~n32044;
  assign n48840 = i_FULL & ~n48839;
  assign n48841 = ~n32054 & ~n48840;
  assign n48842 = i_nEMPTY & ~n48841;
  assign n48843 = ~n32074 & ~n48842;
  assign n48844 = controllable_BtoS_ACK0 & ~n48843;
  assign n48845 = ~n29641 & ~n32088;
  assign n48846 = i_FULL & ~n48845;
  assign n48847 = ~n32098 & ~n48846;
  assign n48848 = i_nEMPTY & ~n48847;
  assign n48849 = ~n32118 & ~n48848;
  assign n48850 = ~controllable_BtoS_ACK0 & ~n48849;
  assign n48851 = ~n48844 & ~n48850;
  assign n48852 = n4465 & ~n48851;
  assign n48853 = ~n21013 & ~n48850;
  assign n48854 = ~n4465 & ~n48853;
  assign n48855 = ~n48852 & ~n48854;
  assign n48856 = i_StoB_REQ10 & ~n48855;
  assign n48857 = ~n23093 & ~n32138;
  assign n48858 = i_FULL & ~n48857;
  assign n48859 = ~n32148 & ~n48858;
  assign n48860 = i_nEMPTY & ~n48859;
  assign n48861 = ~n32168 & ~n48860;
  assign n48862 = controllable_BtoS_ACK0 & ~n48861;
  assign n48863 = ~n23133 & ~n32182;
  assign n48864 = i_FULL & ~n48863;
  assign n48865 = ~n32192 & ~n48864;
  assign n48866 = i_nEMPTY & ~n48865;
  assign n48867 = ~n32212 & ~n48866;
  assign n48868 = ~controllable_BtoS_ACK0 & ~n48867;
  assign n48869 = ~n48862 & ~n48868;
  assign n48870 = n4465 & ~n48869;
  assign n48871 = ~n23127 & ~n48868;
  assign n48872 = ~n4465 & ~n48871;
  assign n48873 = ~n48870 & ~n48872;
  assign n48874 = ~i_StoB_REQ10 & ~n48873;
  assign n48875 = ~n48856 & ~n48874;
  assign n48876 = controllable_BtoS_ACK10 & ~n48875;
  assign n48877 = ~n29844 & ~n32232;
  assign n48878 = i_FULL & ~n48877;
  assign n48879 = ~n32240 & ~n48878;
  assign n48880 = i_nEMPTY & ~n48879;
  assign n48881 = ~n32253 & ~n48880;
  assign n48882 = controllable_BtoS_ACK0 & ~n48881;
  assign n48883 = ~n29900 & ~n32265;
  assign n48884 = i_FULL & ~n48883;
  assign n48885 = ~n32273 & ~n48884;
  assign n48886 = i_nEMPTY & ~n48885;
  assign n48887 = ~n32286 & ~n48886;
  assign n48888 = ~controllable_BtoS_ACK0 & ~n48887;
  assign n48889 = ~n48882 & ~n48888;
  assign n48890 = n4465 & ~n48889;
  assign n48891 = ~n29958 & ~n48888;
  assign n48892 = ~n4465 & ~n48891;
  assign n48893 = ~n48890 & ~n48892;
  assign n48894 = i_StoB_REQ10 & ~n48893;
  assign n48895 = ~n48874 & ~n48894;
  assign n48896 = ~controllable_BtoS_ACK10 & ~n48895;
  assign n48897 = ~n48876 & ~n48896;
  assign n48898 = ~n4464 & ~n48897;
  assign n48899 = ~n48838 & ~n48898;
  assign n48900 = ~n4463 & ~n48899;
  assign n48901 = ~n47646 & ~n48900;
  assign n48902 = n4462 & ~n48901;
  assign n48903 = ~n29844 & ~n32314;
  assign n48904 = i_FULL & ~n48903;
  assign n48905 = ~n32324 & ~n48904;
  assign n48906 = i_nEMPTY & ~n48905;
  assign n48907 = ~n32339 & ~n48906;
  assign n48908 = controllable_BtoS_ACK0 & ~n48907;
  assign n48909 = ~n48830 & ~n48908;
  assign n48910 = n4465 & ~n48909;
  assign n48911 = ~n48832 & ~n48910;
  assign n48912 = i_StoB_REQ10 & ~n48911;
  assign n48913 = ~n23093 & ~n32355;
  assign n48914 = i_FULL & ~n48913;
  assign n48915 = ~n32363 & ~n48914;
  assign n48916 = i_nEMPTY & ~n48915;
  assign n48917 = ~n32381 & ~n48916;
  assign n48918 = controllable_BtoS_ACK0 & ~n48917;
  assign n48919 = ~n48736 & ~n48918;
  assign n48920 = n4465 & ~n48919;
  assign n48921 = ~n48738 & ~n48920;
  assign n48922 = ~i_StoB_REQ10 & ~n48921;
  assign n48923 = ~n48912 & ~n48922;
  assign n48924 = ~controllable_BtoS_ACK10 & ~n48923;
  assign n48925 = ~n30806 & ~n48924;
  assign n48926 = n4464 & ~n48925;
  assign n48927 = ~n30806 & ~n48896;
  assign n48928 = ~n4464 & ~n48927;
  assign n48929 = ~n48926 & ~n48928;
  assign n48930 = ~n4463 & ~n48929;
  assign n48931 = ~n47992 & ~n48930;
  assign n48932 = ~n4462 & ~n48931;
  assign n48933 = ~n48902 & ~n48932;
  assign n48934 = n4461 & ~n48933;
  assign n48935 = ~n14084 & ~n47038;
  assign n48936 = ~controllable_BtoR_REQ0 & ~n48935;
  assign n48937 = ~n47037 & ~n48936;
  assign n48938 = ~i_RtoB_ACK0 & ~n48937;
  assign n48939 = ~n48026 & ~n48938;
  assign n48940 = ~controllable_DEQ & ~n48939;
  assign n48941 = ~n20981 & ~n48940;
  assign n48942 = i_FULL & ~n48941;
  assign n48943 = controllable_BtoR_REQ1 & ~n45168;
  assign n48944 = ~n47038 & ~n48943;
  assign n48945 = ~controllable_BtoR_REQ0 & ~n48944;
  assign n48946 = ~n47037 & ~n48945;
  assign n48947 = ~i_RtoB_ACK0 & ~n48946;
  assign n48948 = ~n48026 & ~n48947;
  assign n48949 = ~controllable_DEQ & ~n48948;
  assign n48950 = ~n20981 & ~n48949;
  assign n48951 = ~i_FULL & ~n48950;
  assign n48952 = ~n48942 & ~n48951;
  assign n48953 = i_nEMPTY & ~n48952;
  assign n48954 = ~n14094 & ~n47051;
  assign n48955 = ~controllable_BtoR_REQ0 & ~n48954;
  assign n48956 = ~n47050 & ~n48955;
  assign n48957 = ~i_RtoB_ACK0 & ~n48956;
  assign n48958 = ~n48042 & ~n48957;
  assign n48959 = ~controllable_DEQ & ~n48958;
  assign n48960 = ~n20993 & ~n48959;
  assign n48961 = i_FULL & ~n48960;
  assign n48962 = controllable_BtoR_REQ1 & ~n45200;
  assign n48963 = ~n47064 & ~n48962;
  assign n48964 = ~controllable_BtoR_REQ0 & ~n48963;
  assign n48965 = ~n47063 & ~n48964;
  assign n48966 = ~i_RtoB_ACK0 & ~n48965;
  assign n48967 = ~n48042 & ~n48966;
  assign n48968 = ~controllable_DEQ & ~n48967;
  assign n48969 = ~n21003 & ~n48968;
  assign n48970 = ~i_FULL & ~n48969;
  assign n48971 = ~n48961 & ~n48970;
  assign n48972 = ~i_nEMPTY & ~n48971;
  assign n48973 = ~n48953 & ~n48972;
  assign n48974 = controllable_BtoS_ACK0 & ~n48973;
  assign n48975 = ~n14127 & ~n47081;
  assign n48976 = ~controllable_BtoR_REQ0 & ~n48975;
  assign n48977 = ~n47080 & ~n48976;
  assign n48978 = ~i_RtoB_ACK0 & ~n48977;
  assign n48979 = ~n48060 & ~n48978;
  assign n48980 = ~controllable_DEQ & ~n48979;
  assign n48981 = ~n29641 & ~n48980;
  assign n48982 = i_FULL & ~n48981;
  assign n48983 = controllable_BtoR_REQ1 & ~n45232;
  assign n48984 = ~n47081 & ~n48983;
  assign n48985 = ~controllable_BtoR_REQ0 & ~n48984;
  assign n48986 = ~n47080 & ~n48985;
  assign n48987 = ~i_RtoB_ACK0 & ~n48986;
  assign n48988 = ~n48060 & ~n48987;
  assign n48989 = ~controllable_DEQ & ~n48988;
  assign n48990 = ~n29641 & ~n48989;
  assign n48991 = ~i_FULL & ~n48990;
  assign n48992 = ~n48982 & ~n48991;
  assign n48993 = i_nEMPTY & ~n48992;
  assign n48994 = ~n14137 & ~n47094;
  assign n48995 = ~controllable_BtoR_REQ0 & ~n48994;
  assign n48996 = ~n47093 & ~n48995;
  assign n48997 = ~i_RtoB_ACK0 & ~n48996;
  assign n48998 = ~n48076 & ~n48997;
  assign n48999 = ~controllable_DEQ & ~n48998;
  assign n49000 = ~n29653 & ~n48999;
  assign n49001 = i_FULL & ~n49000;
  assign n49002 = controllable_BtoR_REQ1 & ~n45264;
  assign n49003 = ~n47107 & ~n49002;
  assign n49004 = ~controllable_BtoR_REQ0 & ~n49003;
  assign n49005 = ~n47106 & ~n49004;
  assign n49006 = ~i_RtoB_ACK0 & ~n49005;
  assign n49007 = ~n48076 & ~n49006;
  assign n49008 = ~controllable_DEQ & ~n49007;
  assign n49009 = ~n29663 & ~n49008;
  assign n49010 = ~i_FULL & ~n49009;
  assign n49011 = ~n49001 & ~n49010;
  assign n49012 = ~i_nEMPTY & ~n49011;
  assign n49013 = ~n48993 & ~n49012;
  assign n49014 = ~controllable_BtoS_ACK0 & ~n49013;
  assign n49015 = ~n48974 & ~n49014;
  assign n49016 = n4465 & ~n49015;
  assign n49017 = ~n29641 & ~n32501;
  assign n49018 = i_FULL & ~n49017;
  assign n49019 = ~n32512 & ~n49018;
  assign n49020 = i_nEMPTY & ~n49019;
  assign n49021 = ~n32530 & ~n49020;
  assign n49022 = ~controllable_BtoS_ACK0 & ~n49021;
  assign n49023 = ~n21013 & ~n49022;
  assign n49024 = ~n4465 & ~n49023;
  assign n49025 = ~n49016 & ~n49024;
  assign n49026 = i_StoB_REQ10 & ~n49025;
  assign n49027 = controllable_BtoR_REQ1 & ~n45387;
  assign n49028 = ~n47135 & ~n49027;
  assign n49029 = ~controllable_BtoR_REQ0 & ~n49028;
  assign n49030 = ~n47134 & ~n49029;
  assign n49031 = ~i_RtoB_ACK0 & ~n49030;
  assign n49032 = ~n48106 & ~n49031;
  assign n49033 = ~controllable_DEQ & ~n49032;
  assign n49034 = ~n23093 & ~n49033;
  assign n49035 = i_FULL & ~n49034;
  assign n49036 = controllable_BtoR_REQ1 & ~n45398;
  assign n49037 = ~n47135 & ~n49036;
  assign n49038 = ~controllable_BtoR_REQ0 & ~n49037;
  assign n49039 = ~n47134 & ~n49038;
  assign n49040 = ~i_RtoB_ACK0 & ~n49039;
  assign n49041 = ~n48106 & ~n49040;
  assign n49042 = ~controllable_DEQ & ~n49041;
  assign n49043 = ~n23093 & ~n49042;
  assign n49044 = ~i_FULL & ~n49043;
  assign n49045 = ~n49035 & ~n49044;
  assign n49046 = i_nEMPTY & ~n49045;
  assign n49047 = controllable_BtoR_REQ1 & ~n45427;
  assign n49048 = ~n47154 & ~n49047;
  assign n49049 = ~controllable_BtoR_REQ0 & ~n49048;
  assign n49050 = ~n47153 & ~n49049;
  assign n49051 = ~i_RtoB_ACK0 & ~n49050;
  assign n49052 = ~n48122 & ~n49051;
  assign n49053 = ~controllable_DEQ & ~n49052;
  assign n49054 = ~n23105 & ~n49053;
  assign n49055 = i_FULL & ~n49054;
  assign n49056 = ~n45860 & ~n46130;
  assign n49057 = ~controllable_BtoR_REQ0 & ~n49056;
  assign n49058 = ~n47172 & ~n49057;
  assign n49059 = ~i_RtoB_ACK0 & ~n49058;
  assign n49060 = ~n48130 & ~n49059;
  assign n49061 = ~controllable_DEQ & ~n49060;
  assign n49062 = ~n23117 & ~n49061;
  assign n49063 = ~i_FULL & ~n49062;
  assign n49064 = ~n49055 & ~n49063;
  assign n49065 = ~i_nEMPTY & ~n49064;
  assign n49066 = ~n49046 & ~n49065;
  assign n49067 = controllable_BtoS_ACK0 & ~n49066;
  assign n49068 = controllable_BtoR_REQ1 & ~n45472;
  assign n49069 = ~n47195 & ~n49068;
  assign n49070 = ~controllable_BtoR_REQ0 & ~n49069;
  assign n49071 = ~n47194 & ~n49070;
  assign n49072 = ~i_RtoB_ACK0 & ~n49071;
  assign n49073 = ~n48142 & ~n49072;
  assign n49074 = ~controllable_DEQ & ~n49073;
  assign n49075 = ~n23133 & ~n49074;
  assign n49076 = i_FULL & ~n49075;
  assign n49077 = controllable_BtoR_REQ1 & ~n45483;
  assign n49078 = ~n47195 & ~n49077;
  assign n49079 = ~controllable_BtoR_REQ0 & ~n49078;
  assign n49080 = ~n47194 & ~n49079;
  assign n49081 = ~i_RtoB_ACK0 & ~n49080;
  assign n49082 = ~n48142 & ~n49081;
  assign n49083 = ~controllable_DEQ & ~n49082;
  assign n49084 = ~n23133 & ~n49083;
  assign n49085 = ~i_FULL & ~n49084;
  assign n49086 = ~n49076 & ~n49085;
  assign n49087 = i_nEMPTY & ~n49086;
  assign n49088 = controllable_BtoR_REQ1 & ~n45512;
  assign n49089 = ~n47214 & ~n49088;
  assign n49090 = ~controllable_BtoR_REQ0 & ~n49089;
  assign n49091 = ~n47213 & ~n49090;
  assign n49092 = ~i_RtoB_ACK0 & ~n49091;
  assign n49093 = ~n48158 & ~n49092;
  assign n49094 = ~controllable_DEQ & ~n49093;
  assign n49095 = ~n23145 & ~n49094;
  assign n49096 = i_FULL & ~n49095;
  assign n49097 = ~n45904 & ~n46167;
  assign n49098 = ~controllable_BtoR_REQ0 & ~n49097;
  assign n49099 = ~n47232 & ~n49098;
  assign n49100 = ~i_RtoB_ACK0 & ~n49099;
  assign n49101 = ~n48166 & ~n49100;
  assign n49102 = ~controllable_DEQ & ~n49101;
  assign n49103 = ~n23157 & ~n49102;
  assign n49104 = ~i_FULL & ~n49103;
  assign n49105 = ~n49096 & ~n49104;
  assign n49106 = ~i_nEMPTY & ~n49105;
  assign n49107 = ~n49087 & ~n49106;
  assign n49108 = ~controllable_BtoS_ACK0 & ~n49107;
  assign n49109 = ~n49067 & ~n49108;
  assign n49110 = n4465 & ~n49109;
  assign n49111 = ~n23133 & ~n32645;
  assign n49112 = i_FULL & ~n49111;
  assign n49113 = ~n32656 & ~n49112;
  assign n49114 = i_nEMPTY & ~n49113;
  assign n49115 = ~n32677 & ~n49114;
  assign n49116 = ~controllable_BtoS_ACK0 & ~n49115;
  assign n49117 = ~n23127 & ~n49116;
  assign n49118 = ~n4465 & ~n49117;
  assign n49119 = ~n49110 & ~n49118;
  assign n49120 = ~i_StoB_REQ10 & ~n49119;
  assign n49121 = ~n49026 & ~n49120;
  assign n49122 = controllable_BtoS_ACK10 & ~n49121;
  assign n49123 = ~n33071 & ~n47252;
  assign n49124 = ~controllable_BtoR_REQ0 & ~n49123;
  assign n49125 = ~n48193 & ~n49124;
  assign n49126 = ~i_RtoB_ACK0 & ~n49125;
  assign n49127 = ~n48192 & ~n49126;
  assign n49128 = ~controllable_DEQ & ~n49127;
  assign n49129 = ~n29844 & ~n49128;
  assign n49130 = i_FULL & ~n49129;
  assign n49131 = controllable_BtoR_REQ1 & ~n45568;
  assign n49132 = ~n47252 & ~n49131;
  assign n49133 = ~controllable_BtoR_REQ0 & ~n49132;
  assign n49134 = ~n48193 & ~n49133;
  assign n49135 = ~i_RtoB_ACK0 & ~n49134;
  assign n49136 = ~n48192 & ~n49135;
  assign n49137 = ~controllable_DEQ & ~n49136;
  assign n49138 = ~n29844 & ~n49137;
  assign n49139 = ~i_FULL & ~n49138;
  assign n49140 = ~n49130 & ~n49139;
  assign n49141 = i_nEMPTY & ~n49140;
  assign n49142 = ~n33091 & ~n47259;
  assign n49143 = ~controllable_BtoR_REQ0 & ~n49142;
  assign n49144 = ~n48210 & ~n49143;
  assign n49145 = ~i_RtoB_ACK0 & ~n49144;
  assign n49146 = ~n48209 & ~n49145;
  assign n49147 = ~controllable_DEQ & ~n49146;
  assign n49148 = ~n29858 & ~n49147;
  assign n49149 = i_FULL & ~n49148;
  assign n49150 = ~n45943 & ~n46204;
  assign n49151 = ~controllable_BtoR_REQ0 & ~n49150;
  assign n49152 = ~n48219 & ~n49151;
  assign n49153 = ~i_RtoB_ACK0 & ~n49152;
  assign n49154 = ~n48218 & ~n49153;
  assign n49155 = ~controllable_DEQ & ~n49154;
  assign n49156 = ~n29872 & ~n49155;
  assign n49157 = ~i_FULL & ~n49156;
  assign n49158 = ~n49149 & ~n49157;
  assign n49159 = ~i_nEMPTY & ~n49158;
  assign n49160 = ~n49141 & ~n49159;
  assign n49161 = controllable_BtoS_ACK0 & ~n49160;
  assign n49162 = ~n32639 & ~n47282;
  assign n49163 = ~controllable_BtoR_REQ0 & ~n49162;
  assign n49164 = ~n48232 & ~n49163;
  assign n49165 = ~i_RtoB_ACK0 & ~n49164;
  assign n49166 = ~n48231 & ~n49165;
  assign n49167 = ~controllable_DEQ & ~n49166;
  assign n49168 = ~n29900 & ~n49167;
  assign n49169 = i_FULL & ~n49168;
  assign n49170 = controllable_BtoR_REQ1 & ~n45626;
  assign n49171 = ~n47282 & ~n49170;
  assign n49172 = ~controllable_BtoR_REQ0 & ~n49171;
  assign n49173 = ~n48232 & ~n49172;
  assign n49174 = ~i_RtoB_ACK0 & ~n49173;
  assign n49175 = ~n48231 & ~n49174;
  assign n49176 = ~controllable_DEQ & ~n49175;
  assign n49177 = ~n29900 & ~n49176;
  assign n49178 = ~i_FULL & ~n49177;
  assign n49179 = ~n49169 & ~n49178;
  assign n49180 = i_nEMPTY & ~n49179;
  assign n49181 = ~n32659 & ~n47289;
  assign n49182 = ~controllable_BtoR_REQ0 & ~n49181;
  assign n49183 = ~n48249 & ~n49182;
  assign n49184 = ~i_RtoB_ACK0 & ~n49183;
  assign n49185 = ~n48248 & ~n49184;
  assign n49186 = ~controllable_DEQ & ~n49185;
  assign n49187 = ~n29914 & ~n49186;
  assign n49188 = i_FULL & ~n49187;
  assign n49189 = ~n45975 & ~n46235;
  assign n49190 = ~controllable_BtoR_REQ0 & ~n49189;
  assign n49191 = ~n48258 & ~n49190;
  assign n49192 = ~i_RtoB_ACK0 & ~n49191;
  assign n49193 = ~n48257 & ~n49192;
  assign n49194 = ~controllable_DEQ & ~n49193;
  assign n49195 = ~n29928 & ~n49194;
  assign n49196 = ~i_FULL & ~n49195;
  assign n49197 = ~n49188 & ~n49196;
  assign n49198 = ~i_nEMPTY & ~n49197;
  assign n49199 = ~n49180 & ~n49198;
  assign n49200 = ~controllable_BtoS_ACK0 & ~n49199;
  assign n49201 = ~n49161 & ~n49200;
  assign n49202 = n4465 & ~n49201;
  assign n49203 = ~n29900 & ~n32763;
  assign n49204 = i_FULL & ~n49203;
  assign n49205 = ~n32771 & ~n49204;
  assign n49206 = i_nEMPTY & ~n49205;
  assign n49207 = ~n32784 & ~n49206;
  assign n49208 = ~controllable_BtoS_ACK0 & ~n49207;
  assign n49209 = ~n29958 & ~n49208;
  assign n49210 = ~n4465 & ~n49209;
  assign n49211 = ~n49202 & ~n49210;
  assign n49212 = i_StoB_REQ10 & ~n49211;
  assign n49213 = ~n49120 & ~n49212;
  assign n49214 = ~controllable_BtoS_ACK10 & ~n49213;
  assign n49215 = ~n49122 & ~n49214;
  assign n49216 = n4464 & ~n49215;
  assign n49217 = ~n20981 & ~n32804;
  assign n49218 = i_FULL & ~n49217;
  assign n49219 = ~n32815 & ~n49218;
  assign n49220 = i_nEMPTY & ~n49219;
  assign n49221 = ~n32833 & ~n49220;
  assign n49222 = controllable_BtoS_ACK0 & ~n49221;
  assign n49223 = ~n29641 & ~n32845;
  assign n49224 = i_FULL & ~n49223;
  assign n49225 = ~n32856 & ~n49224;
  assign n49226 = i_nEMPTY & ~n49225;
  assign n49227 = ~n32874 & ~n49226;
  assign n49228 = ~controllable_BtoS_ACK0 & ~n49227;
  assign n49229 = ~n49222 & ~n49228;
  assign n49230 = n4465 & ~n49229;
  assign n49231 = ~n21013 & ~n49228;
  assign n49232 = ~n4465 & ~n49231;
  assign n49233 = ~n49230 & ~n49232;
  assign n49234 = i_StoB_REQ10 & ~n49233;
  assign n49235 = ~n23093 & ~n32895;
  assign n49236 = i_FULL & ~n49235;
  assign n49237 = ~n32906 & ~n49236;
  assign n49238 = i_nEMPTY & ~n49237;
  assign n49239 = ~n32927 & ~n49238;
  assign n49240 = controllable_BtoS_ACK0 & ~n49239;
  assign n49241 = ~n23133 & ~n32942;
  assign n49242 = i_FULL & ~n49241;
  assign n49243 = ~n32953 & ~n49242;
  assign n49244 = i_nEMPTY & ~n49243;
  assign n49245 = ~n32974 & ~n49244;
  assign n49246 = ~controllable_BtoS_ACK0 & ~n49245;
  assign n49247 = ~n49240 & ~n49246;
  assign n49248 = n4465 & ~n49247;
  assign n49249 = ~n23127 & ~n49246;
  assign n49250 = ~n4465 & ~n49249;
  assign n49251 = ~n49248 & ~n49250;
  assign n49252 = ~i_StoB_REQ10 & ~n49251;
  assign n49253 = ~n49234 & ~n49252;
  assign n49254 = controllable_BtoS_ACK10 & ~n49253;
  assign n49255 = ~n29844 & ~n32994;
  assign n49256 = i_FULL & ~n49255;
  assign n49257 = ~n33002 & ~n49256;
  assign n49258 = i_nEMPTY & ~n49257;
  assign n49259 = ~n33015 & ~n49258;
  assign n49260 = controllable_BtoS_ACK0 & ~n49259;
  assign n49261 = ~n29900 & ~n33027;
  assign n49262 = i_FULL & ~n49261;
  assign n49263 = ~n33035 & ~n49262;
  assign n49264 = i_nEMPTY & ~n49263;
  assign n49265 = ~n33048 & ~n49264;
  assign n49266 = ~controllable_BtoS_ACK0 & ~n49265;
  assign n49267 = ~n49260 & ~n49266;
  assign n49268 = n4465 & ~n49267;
  assign n49269 = ~n29958 & ~n49266;
  assign n49270 = ~n4465 & ~n49269;
  assign n49271 = ~n49268 & ~n49270;
  assign n49272 = i_StoB_REQ10 & ~n49271;
  assign n49273 = ~n49252 & ~n49272;
  assign n49274 = ~controllable_BtoS_ACK10 & ~n49273;
  assign n49275 = ~n49254 & ~n49274;
  assign n49276 = ~n4464 & ~n49275;
  assign n49277 = ~n49216 & ~n49276;
  assign n49278 = n4463 & ~n49277;
  assign n49279 = ~n48518 & ~n49278;
  assign n49280 = n4462 & ~n49279;
  assign n49281 = ~n29844 & ~n33077;
  assign n49282 = i_FULL & ~n49281;
  assign n49283 = ~n33088 & ~n49282;
  assign n49284 = i_nEMPTY & ~n49283;
  assign n49285 = ~n33104 & ~n49284;
  assign n49286 = controllable_BtoS_ACK0 & ~n49285;
  assign n49287 = ~n49208 & ~n49286;
  assign n49288 = n4465 & ~n49287;
  assign n49289 = ~n49210 & ~n49288;
  assign n49290 = i_StoB_REQ10 & ~n49289;
  assign n49291 = ~n23093 & ~n33120;
  assign n49292 = i_FULL & ~n49291;
  assign n49293 = ~n33128 & ~n49292;
  assign n49294 = i_nEMPTY & ~n49293;
  assign n49295 = ~n33146 & ~n49294;
  assign n49296 = controllable_BtoS_ACK0 & ~n49295;
  assign n49297 = ~n49116 & ~n49296;
  assign n49298 = n4465 & ~n49297;
  assign n49299 = ~n49118 & ~n49298;
  assign n49300 = ~i_StoB_REQ10 & ~n49299;
  assign n49301 = ~n49290 & ~n49300;
  assign n49302 = ~controllable_BtoS_ACK10 & ~n49301;
  assign n49303 = ~n30806 & ~n49302;
  assign n49304 = n4464 & ~n49303;
  assign n49305 = ~n30806 & ~n49274;
  assign n49306 = ~n4464 & ~n49305;
  assign n49307 = ~n49304 & ~n49306;
  assign n49308 = n4463 & ~n49307;
  assign n49309 = ~n31548 & ~n49308;
  assign n49310 = ~n4462 & ~n49309;
  assign n49311 = ~n49280 & ~n49310;
  assign n49312 = ~n4461 & ~n49311;
  assign n49313 = ~n48934 & ~n49312;
  assign n49314 = n4459 & ~n49313;
  assign n49315 = ~n48554 & ~n49314;
  assign n49316 = ~n4455 & ~n49315;
  assign n49317 = ~n47330 & ~n49316;
  assign n49318 = ~n4445 & ~n49317;
  assign n49319 = ~n45149 & ~n49318;
  assign n49320 = n4442 & ~n49319;
  assign n49321 = ~n7563 & ~n36879;
  assign n49322 = ~controllable_BtoR_REQ1 & ~n49321;
  assign n49323 = ~n48555 & ~n49322;
  assign n49324 = ~controllable_BtoR_REQ0 & ~n49323;
  assign n49325 = ~controllable_BtoR_REQ0 & ~n49324;
  assign n49326 = ~i_RtoB_ACK0 & ~n49325;
  assign n49327 = ~n5259 & ~n49326;
  assign n49328 = ~controllable_DEQ & ~n49327;
  assign n49329 = ~n5251 & ~n49328;
  assign n49330 = i_nEMPTY & ~n49329;
  assign n49331 = ~n5237 & ~n36914;
  assign n49332 = ~controllable_BtoR_REQ1 & ~n49331;
  assign n49333 = ~n48574 & ~n49332;
  assign n49334 = ~controllable_BtoR_REQ0 & ~n49333;
  assign n49335 = ~controllable_BtoR_REQ0 & ~n49334;
  assign n49336 = ~i_RtoB_ACK0 & ~n49335;
  assign n49337 = ~n5236 & ~n49336;
  assign n49338 = ~controllable_DEQ & ~n49337;
  assign n49339 = ~n5281 & ~n49338;
  assign n49340 = i_FULL & ~n49339;
  assign n49341 = ~n5237 & ~n45773;
  assign n49342 = ~controllable_BtoR_REQ1 & ~n49341;
  assign n49343 = ~n48583 & ~n49342;
  assign n49344 = ~controllable_BtoR_REQ0 & ~n49343;
  assign n49345 = ~controllable_BtoR_REQ0 & ~n49344;
  assign n49346 = ~i_RtoB_ACK0 & ~n49345;
  assign n49347 = ~n5236 & ~n49346;
  assign n49348 = ~controllable_DEQ & ~n49347;
  assign n49349 = ~n5296 & ~n49348;
  assign n49350 = ~i_FULL & ~n49349;
  assign n49351 = ~n49340 & ~n49350;
  assign n49352 = ~i_nEMPTY & ~n49351;
  assign n49353 = ~n49330 & ~n49352;
  assign n49354 = controllable_BtoS_ACK0 & ~n49353;
  assign n49355 = ~n8883 & ~n37060;
  assign n49356 = ~controllable_BtoR_REQ1 & ~n49355;
  assign n49357 = ~n48596 & ~n49356;
  assign n49358 = ~controllable_BtoR_REQ0 & ~n49357;
  assign n49359 = ~controllable_BtoR_REQ0 & ~n49358;
  assign n49360 = ~i_RtoB_ACK0 & ~n49359;
  assign n49361 = ~n27871 & ~n49360;
  assign n49362 = ~controllable_DEQ & ~n49361;
  assign n49363 = ~n27884 & ~n49362;
  assign n49364 = i_nEMPTY & ~n49363;
  assign n49365 = ~n8861 & ~n37095;
  assign n49366 = ~controllable_BtoR_REQ1 & ~n49365;
  assign n49367 = ~n48615 & ~n49366;
  assign n49368 = ~controllable_BtoR_REQ0 & ~n49367;
  assign n49369 = ~controllable_BtoR_REQ0 & ~n49368;
  assign n49370 = ~i_RtoB_ACK0 & ~n49369;
  assign n49371 = ~n27859 & ~n49370;
  assign n49372 = ~controllable_DEQ & ~n49371;
  assign n49373 = ~n27900 & ~n49372;
  assign n49374 = i_FULL & ~n49373;
  assign n49375 = ~n8861 & ~n45811;
  assign n49376 = ~controllable_BtoR_REQ1 & ~n49375;
  assign n49377 = ~n48624 & ~n49376;
  assign n49378 = ~controllable_BtoR_REQ0 & ~n49377;
  assign n49379 = ~controllable_BtoR_REQ0 & ~n49378;
  assign n49380 = ~i_RtoB_ACK0 & ~n49379;
  assign n49381 = ~n27859 & ~n49380;
  assign n49382 = ~controllable_DEQ & ~n49381;
  assign n49383 = ~n27912 & ~n49382;
  assign n49384 = ~i_FULL & ~n49383;
  assign n49385 = ~n49374 & ~n49384;
  assign n49386 = ~i_nEMPTY & ~n49385;
  assign n49387 = ~n49364 & ~n49386;
  assign n49388 = ~controllable_BtoS_ACK0 & ~n49387;
  assign n49389 = ~n49354 & ~n49388;
  assign n49390 = n4465 & ~n49389;
  assign n49391 = ~n45826 & ~n49390;
  assign n49392 = i_StoB_REQ10 & ~n49391;
  assign n49393 = ~n47252 & ~n48649;
  assign n49394 = ~controllable_BtoR_REQ0 & ~n49393;
  assign n49395 = ~controllable_BtoR_REQ0 & ~n49394;
  assign n49396 = ~i_RtoB_ACK0 & ~n49395;
  assign n49397 = ~n11252 & ~n49396;
  assign n49398 = ~controllable_DEQ & ~n49397;
  assign n49399 = ~n11244 & ~n49398;
  assign n49400 = i_nEMPTY & ~n49399;
  assign n49401 = ~n47259 & ~n48668;
  assign n49402 = ~controllable_BtoR_REQ0 & ~n49401;
  assign n49403 = ~controllable_BtoR_REQ0 & ~n49402;
  assign n49404 = ~i_RtoB_ACK0 & ~n49403;
  assign n49405 = ~n11234 & ~n49404;
  assign n49406 = ~controllable_DEQ & ~n49405;
  assign n49407 = ~n11269 & ~n49406;
  assign n49408 = i_FULL & ~n49407;
  assign n49409 = ~n9571 & ~n45856;
  assign n49410 = ~controllable_BtoR_REQ1 & ~n49409;
  assign n49411 = ~n45858 & ~n49410;
  assign n49412 = ~controllable_BtoR_REQ0 & ~n49411;
  assign n49413 = ~controllable_BtoR_REQ0 & ~n49412;
  assign n49414 = ~i_RtoB_ACK0 & ~n49413;
  assign n49415 = ~n11234 & ~n49414;
  assign n49416 = ~controllable_DEQ & ~n49415;
  assign n49417 = ~n11282 & ~n49416;
  assign n49418 = ~i_FULL & ~n49417;
  assign n49419 = ~n49408 & ~n49418;
  assign n49420 = ~i_nEMPTY & ~n49419;
  assign n49421 = ~n49400 & ~n49420;
  assign n49422 = controllable_BtoS_ACK0 & ~n49421;
  assign n49423 = ~n47282 & ~n48689;
  assign n49424 = ~controllable_BtoR_REQ0 & ~n49423;
  assign n49425 = ~controllable_BtoR_REQ0 & ~n49424;
  assign n49426 = ~i_RtoB_ACK0 & ~n49425;
  assign n49427 = ~n11332 & ~n49426;
  assign n49428 = ~controllable_DEQ & ~n49427;
  assign n49429 = ~n11323 & ~n49428;
  assign n49430 = i_nEMPTY & ~n49429;
  assign n49431 = ~n47289 & ~n48708;
  assign n49432 = ~controllable_BtoR_REQ0 & ~n49431;
  assign n49433 = ~controllable_BtoR_REQ0 & ~n49432;
  assign n49434 = ~i_RtoB_ACK0 & ~n49433;
  assign n49435 = ~n11309 & ~n49434;
  assign n49436 = ~controllable_DEQ & ~n49435;
  assign n49437 = ~n11351 & ~n49436;
  assign n49438 = i_FULL & ~n49437;
  assign n49439 = ~n9718 & ~n45900;
  assign n49440 = ~controllable_BtoR_REQ1 & ~n49439;
  assign n49441 = ~n45902 & ~n49440;
  assign n49442 = ~controllable_BtoR_REQ0 & ~n49441;
  assign n49443 = ~controllable_BtoR_REQ0 & ~n49442;
  assign n49444 = ~i_RtoB_ACK0 & ~n49443;
  assign n49445 = ~n11309 & ~n49444;
  assign n49446 = ~controllable_DEQ & ~n49445;
  assign n49447 = ~n11364 & ~n49446;
  assign n49448 = ~i_FULL & ~n49447;
  assign n49449 = ~n49438 & ~n49448;
  assign n49450 = ~i_nEMPTY & ~n49449;
  assign n49451 = ~n49430 & ~n49450;
  assign n49452 = ~controllable_BtoS_ACK0 & ~n49451;
  assign n49453 = ~n49422 & ~n49452;
  assign n49454 = n4465 & ~n49453;
  assign n49455 = ~n45919 & ~n49454;
  assign n49456 = ~i_StoB_REQ10 & ~n49455;
  assign n49457 = ~n49392 & ~n49456;
  assign n49458 = controllable_BtoS_ACK10 & ~n49457;
  assign n49459 = ~n45992 & ~n49456;
  assign n49460 = ~controllable_BtoS_ACK10 & ~n49459;
  assign n49461 = ~n49458 & ~n49460;
  assign n49462 = n4464 & ~n49461;
  assign n49463 = ~n45997 & ~n49462;
  assign n49464 = n4463 & ~n49463;
  assign n49465 = ~n7563 & ~n12185;
  assign n49466 = ~controllable_BtoR_REQ0 & ~n49465;
  assign n49467 = ~controllable_BtoR_REQ0 & ~n49466;
  assign n49468 = ~i_RtoB_ACK0 & ~n49467;
  assign n49469 = ~n5259 & ~n49468;
  assign n49470 = ~controllable_DEQ & ~n49469;
  assign n49471 = ~n5251 & ~n49470;
  assign n49472 = i_nEMPTY & ~n49471;
  assign n49473 = ~n5237 & ~n12164;
  assign n49474 = ~controllable_BtoR_REQ0 & ~n49473;
  assign n49475 = ~controllable_BtoR_REQ0 & ~n49474;
  assign n49476 = ~i_RtoB_ACK0 & ~n49475;
  assign n49477 = ~n5236 & ~n49476;
  assign n49478 = ~controllable_DEQ & ~n49477;
  assign n49479 = ~n5281 & ~n49478;
  assign n49480 = i_FULL & ~n49479;
  assign n49481 = ~n12162 & ~n38877;
  assign n49482 = ~i_RtoB_ACK1 & ~n49481;
  assign n49483 = ~n5237 & ~n49482;
  assign n49484 = ~controllable_BtoR_REQ0 & ~n49483;
  assign n49485 = ~controllable_BtoR_REQ0 & ~n49484;
  assign n49486 = ~i_RtoB_ACK0 & ~n49485;
  assign n49487 = ~n5236 & ~n49486;
  assign n49488 = ~controllable_DEQ & ~n49487;
  assign n49489 = ~n5296 & ~n49488;
  assign n49490 = ~i_FULL & ~n49489;
  assign n49491 = ~n49480 & ~n49490;
  assign n49492 = ~i_nEMPTY & ~n49491;
  assign n49493 = ~n49472 & ~n49492;
  assign n49494 = controllable_BtoS_ACK0 & ~n49493;
  assign n49495 = ~n8883 & ~n12275;
  assign n49496 = ~controllable_BtoR_REQ0 & ~n49495;
  assign n49497 = ~controllable_BtoR_REQ0 & ~n49496;
  assign n49498 = ~i_RtoB_ACK0 & ~n49497;
  assign n49499 = ~n27871 & ~n49498;
  assign n49500 = ~controllable_DEQ & ~n49499;
  assign n49501 = ~n27884 & ~n49500;
  assign n49502 = i_nEMPTY & ~n49501;
  assign n49503 = ~n8861 & ~n12257;
  assign n49504 = ~controllable_BtoR_REQ0 & ~n49503;
  assign n49505 = ~controllable_BtoR_REQ0 & ~n49504;
  assign n49506 = ~i_RtoB_ACK0 & ~n49505;
  assign n49507 = ~n27859 & ~n49506;
  assign n49508 = ~controllable_DEQ & ~n49507;
  assign n49509 = ~n27900 & ~n49508;
  assign n49510 = i_FULL & ~n49509;
  assign n49511 = ~n12255 & ~n38972;
  assign n49512 = ~i_RtoB_ACK1 & ~n49511;
  assign n49513 = ~n8861 & ~n49512;
  assign n49514 = ~controllable_BtoR_REQ0 & ~n49513;
  assign n49515 = ~controllable_BtoR_REQ0 & ~n49514;
  assign n49516 = ~i_RtoB_ACK0 & ~n49515;
  assign n49517 = ~n27859 & ~n49516;
  assign n49518 = ~controllable_DEQ & ~n49517;
  assign n49519 = ~n27912 & ~n49518;
  assign n49520 = ~i_FULL & ~n49519;
  assign n49521 = ~n49510 & ~n49520;
  assign n49522 = ~i_nEMPTY & ~n49521;
  assign n49523 = ~n49502 & ~n49522;
  assign n49524 = ~controllable_BtoS_ACK0 & ~n49523;
  assign n49525 = ~n49494 & ~n49524;
  assign n49526 = n4465 & ~n49525;
  assign n49527 = ~n45826 & ~n49526;
  assign n49528 = i_StoB_REQ10 & ~n49527;
  assign n49529 = ~n9517 & ~n46820;
  assign n49530 = ~controllable_BtoR_REQ0 & ~n49529;
  assign n49531 = ~controllable_BtoR_REQ0 & ~n49530;
  assign n49532 = ~i_RtoB_ACK0 & ~n49531;
  assign n49533 = ~n11252 & ~n49532;
  assign n49534 = ~controllable_DEQ & ~n49533;
  assign n49535 = ~n11244 & ~n49534;
  assign n49536 = i_nEMPTY & ~n49535;
  assign n49537 = ~n9571 & ~n46837;
  assign n49538 = ~controllable_BtoR_REQ0 & ~n49537;
  assign n49539 = ~controllable_BtoR_REQ0 & ~n49538;
  assign n49540 = ~i_RtoB_ACK0 & ~n49539;
  assign n49541 = ~n11234 & ~n49540;
  assign n49542 = ~controllable_DEQ & ~n49541;
  assign n49543 = ~n11269 & ~n49542;
  assign n49544 = i_FULL & ~n49543;
  assign n49545 = i_StoB_REQ14 & ~n38870;
  assign n49546 = i_StoB_REQ0 & ~n38868;
  assign n49547 = controllable_BtoS_ACK13 & ~n38864;
  assign n49548 = ~controllable_BtoS_ACK13 & ~n45367;
  assign n49549 = ~n49547 & ~n49548;
  assign n49550 = i_StoB_REQ13 & ~n49549;
  assign n49551 = i_StoB_REQ12 & ~n38857;
  assign n49552 = i_StoB_REQ11 & ~n38848;
  assign n49553 = i_StoB_REQ9 & ~n38839;
  assign n49554 = i_StoB_REQ7 & ~n38829;
  assign n49555 = i_StoB_REQ6 & ~n38822;
  assign n49556 = i_StoB_REQ8 & ~n38812;
  assign n49557 = i_StoB_REQ5 & ~n38804;
  assign n49558 = i_StoB_REQ4 & ~n38796;
  assign n49559 = i_StoB_REQ3 & ~n38788;
  assign n49560 = ~n37567 & ~n38785;
  assign n49561 = n4476 & ~n49560;
  assign n49562 = ~n37570 & ~n49561;
  assign n49563 = ~i_StoB_REQ3 & ~n49562;
  assign n49564 = ~n49559 & ~n49563;
  assign n49565 = controllable_BtoS_ACK3 & ~n49564;
  assign n49566 = i_StoB_REQ3 & ~n45295;
  assign n49567 = ~n49563 & ~n49566;
  assign n49568 = ~controllable_BtoS_ACK3 & ~n49567;
  assign n49569 = ~n49565 & ~n49568;
  assign n49570 = n4475 & ~n49569;
  assign n49571 = ~n37579 & ~n49570;
  assign n49572 = ~i_StoB_REQ4 & ~n49571;
  assign n49573 = ~n49558 & ~n49572;
  assign n49574 = controllable_BtoS_ACK4 & ~n49573;
  assign n49575 = i_StoB_REQ4 & ~n45303;
  assign n49576 = ~n49572 & ~n49575;
  assign n49577 = ~controllable_BtoS_ACK4 & ~n49576;
  assign n49578 = ~n49574 & ~n49577;
  assign n49579 = n4474 & ~n49578;
  assign n49580 = ~n37588 & ~n49579;
  assign n49581 = ~i_StoB_REQ5 & ~n49580;
  assign n49582 = ~n49557 & ~n49581;
  assign n49583 = controllable_BtoS_ACK5 & ~n49582;
  assign n49584 = i_StoB_REQ5 & ~n45311;
  assign n49585 = ~n49581 & ~n49584;
  assign n49586 = ~controllable_BtoS_ACK5 & ~n49585;
  assign n49587 = ~n49583 & ~n49586;
  assign n49588 = n4473 & ~n49587;
  assign n49589 = ~n37597 & ~n49588;
  assign n49590 = ~i_StoB_REQ8 & ~n49589;
  assign n49591 = ~n49556 & ~n49590;
  assign n49592 = controllable_BtoS_ACK8 & ~n49591;
  assign n49593 = i_StoB_REQ8 & ~n45319;
  assign n49594 = ~n49590 & ~n49593;
  assign n49595 = ~controllable_BtoS_ACK8 & ~n49594;
  assign n49596 = ~n49592 & ~n49595;
  assign n49597 = n4472 & ~n49596;
  assign n49598 = ~n37606 & ~n49597;
  assign n49599 = n4471 & ~n49598;
  assign n49600 = ~n6345 & ~n49599;
  assign n49601 = ~i_StoB_REQ6 & ~n49600;
  assign n49602 = ~n49555 & ~n49601;
  assign n49603 = controllable_BtoS_ACK6 & ~n49602;
  assign n49604 = i_StoB_REQ6 & ~n45329;
  assign n49605 = ~n49601 & ~n49604;
  assign n49606 = ~controllable_BtoS_ACK6 & ~n49605;
  assign n49607 = ~n49603 & ~n49606;
  assign n49608 = ~i_StoB_REQ7 & ~n49607;
  assign n49609 = ~n49554 & ~n49608;
  assign n49610 = controllable_BtoS_ACK7 & ~n49609;
  assign n49611 = i_StoB_REQ7 & ~n45335;
  assign n49612 = ~n49608 & ~n49611;
  assign n49613 = ~controllable_BtoS_ACK7 & ~n49612;
  assign n49614 = ~n49610 & ~n49613;
  assign n49615 = n4470 & ~n49614;
  assign n49616 = ~n37623 & ~n49615;
  assign n49617 = n4469 & ~n49616;
  assign n49618 = ~n6408 & ~n49617;
  assign n49619 = ~i_StoB_REQ9 & ~n49618;
  assign n49620 = ~n49553 & ~n49619;
  assign n49621 = controllable_BtoS_ACK9 & ~n49620;
  assign n49622 = i_StoB_REQ9 & ~n45345;
  assign n49623 = ~n49619 & ~n49622;
  assign n49624 = ~controllable_BtoS_ACK9 & ~n49623;
  assign n49625 = ~n49621 & ~n49624;
  assign n49626 = n4468 & ~n49625;
  assign n49627 = ~n6436 & ~n49626;
  assign n49628 = ~i_StoB_REQ11 & ~n49627;
  assign n49629 = ~n49552 & ~n49628;
  assign n49630 = controllable_BtoS_ACK11 & ~n49629;
  assign n49631 = i_StoB_REQ11 & ~n45353;
  assign n49632 = ~n49628 & ~n49631;
  assign n49633 = ~controllable_BtoS_ACK11 & ~n49632;
  assign n49634 = ~n49630 & ~n49633;
  assign n49635 = n4467 & ~n49634;
  assign n49636 = ~n6466 & ~n49635;
  assign n49637 = ~i_StoB_REQ12 & ~n49636;
  assign n49638 = ~n49551 & ~n49637;
  assign n49639 = controllable_BtoS_ACK12 & ~n49638;
  assign n49640 = i_StoB_REQ12 & ~n45361;
  assign n49641 = ~n49637 & ~n49640;
  assign n49642 = ~controllable_BtoS_ACK12 & ~n49641;
  assign n49643 = ~n49639 & ~n49642;
  assign n49644 = ~i_StoB_REQ13 & ~n49643;
  assign n49645 = ~n49550 & ~n49644;
  assign n49646 = n4466 & ~n49645;
  assign n49647 = ~n37652 & ~n49646;
  assign n49648 = ~i_StoB_REQ0 & ~n49647;
  assign n49649 = ~n49546 & ~n49648;
  assign n49650 = ~i_StoB_REQ14 & ~n49649;
  assign n49651 = ~n49545 & ~n49650;
  assign n49652 = controllable_BtoS_ACK14 & ~n49651;
  assign n49653 = i_StoB_REQ14 & ~n45373;
  assign n49654 = ~n49650 & ~n49653;
  assign n49655 = ~controllable_BtoS_ACK14 & ~n49654;
  assign n49656 = ~n49652 & ~n49655;
  assign n49657 = ~controllable_ENQ & ~n49656;
  assign n49658 = ~n45418 & ~n49657;
  assign n49659 = ~i_RtoB_ACK1 & ~n49658;
  assign n49660 = ~n9789 & ~n49659;
  assign n49661 = controllable_BtoR_REQ1 & ~n49660;
  assign n49662 = ~n9571 & ~n49659;
  assign n49663 = ~controllable_BtoR_REQ1 & ~n49662;
  assign n49664 = ~n49661 & ~n49663;
  assign n49665 = ~controllable_BtoR_REQ0 & ~n49664;
  assign n49666 = ~controllable_BtoR_REQ0 & ~n49665;
  assign n49667 = ~i_RtoB_ACK0 & ~n49666;
  assign n49668 = ~n11234 & ~n49667;
  assign n49669 = ~controllable_DEQ & ~n49668;
  assign n49670 = ~n11282 & ~n49669;
  assign n49671 = ~i_FULL & ~n49670;
  assign n49672 = ~n49544 & ~n49671;
  assign n49673 = ~i_nEMPTY & ~n49672;
  assign n49674 = ~n49536 & ~n49673;
  assign n49675 = controllable_BtoS_ACK0 & ~n49674;
  assign n49676 = ~n9664 & ~n46863;
  assign n49677 = ~controllable_BtoR_REQ0 & ~n49676;
  assign n49678 = ~controllable_BtoR_REQ0 & ~n49677;
  assign n49679 = ~i_RtoB_ACK0 & ~n49678;
  assign n49680 = ~n11332 & ~n49679;
  assign n49681 = ~controllable_DEQ & ~n49680;
  assign n49682 = ~n11323 & ~n49681;
  assign n49683 = i_nEMPTY & ~n49682;
  assign n49684 = ~n9718 & ~n46880;
  assign n49685 = ~controllable_BtoR_REQ0 & ~n49684;
  assign n49686 = ~controllable_BtoR_REQ0 & ~n49685;
  assign n49687 = ~i_RtoB_ACK0 & ~n49686;
  assign n49688 = ~n11309 & ~n49687;
  assign n49689 = ~controllable_DEQ & ~n49688;
  assign n49690 = ~n11351 & ~n49689;
  assign n49691 = i_FULL & ~n49690;
  assign n49692 = i_StoB_REQ14 & ~n38965;
  assign n49693 = i_StoB_REQ0 & ~n45371;
  assign n49694 = ~n49648 & ~n49693;
  assign n49695 = ~i_StoB_REQ14 & ~n49694;
  assign n49696 = ~n49692 & ~n49695;
  assign n49697 = controllable_BtoS_ACK14 & ~n49696;
  assign n49698 = i_StoB_REQ14 & ~n45458;
  assign n49699 = ~n49695 & ~n49698;
  assign n49700 = ~controllable_BtoS_ACK14 & ~n49699;
  assign n49701 = ~n49697 & ~n49700;
  assign n49702 = ~controllable_ENQ & ~n49701;
  assign n49703 = ~n45503 & ~n49702;
  assign n49704 = ~i_RtoB_ACK1 & ~n49703;
  assign n49705 = ~n11311 & ~n49704;
  assign n49706 = controllable_BtoR_REQ1 & ~n49705;
  assign n49707 = ~n9718 & ~n49704;
  assign n49708 = ~controllable_BtoR_REQ1 & ~n49707;
  assign n49709 = ~n49706 & ~n49708;
  assign n49710 = ~controllable_BtoR_REQ0 & ~n49709;
  assign n49711 = ~controllable_BtoR_REQ0 & ~n49710;
  assign n49712 = ~i_RtoB_ACK0 & ~n49711;
  assign n49713 = ~n11309 & ~n49712;
  assign n49714 = ~controllable_DEQ & ~n49713;
  assign n49715 = ~n11364 & ~n49714;
  assign n49716 = ~i_FULL & ~n49715;
  assign n49717 = ~n49691 & ~n49716;
  assign n49718 = ~i_nEMPTY & ~n49717;
  assign n49719 = ~n49683 & ~n49718;
  assign n49720 = ~controllable_BtoS_ACK0 & ~n49719;
  assign n49721 = ~n49675 & ~n49720;
  assign n49722 = n4465 & ~n49721;
  assign n49723 = ~n45919 & ~n49722;
  assign n49724 = ~i_StoB_REQ10 & ~n49723;
  assign n49725 = ~n49528 & ~n49724;
  assign n49726 = controllable_BtoS_ACK10 & ~n49725;
  assign n49727 = ~controllable_ENQ & ~n45379;
  assign n49728 = ~n9302 & ~n49727;
  assign n49729 = ~i_RtoB_ACK1 & ~n49728;
  assign n49730 = ~n10149 & ~n49729;
  assign n49731 = controllable_BtoR_REQ1 & ~n49730;
  assign n49732 = ~n9571 & ~n49729;
  assign n49733 = ~controllable_BtoR_REQ1 & ~n49732;
  assign n49734 = ~n49731 & ~n49733;
  assign n49735 = ~controllable_BtoR_REQ0 & ~n49734;
  assign n49736 = ~controllable_BtoR_REQ0 & ~n49735;
  assign n49737 = ~i_RtoB_ACK0 & ~n49736;
  assign n49738 = ~n28114 & ~n49737;
  assign n49739 = ~controllable_DEQ & ~n49738;
  assign n49740 = ~n28163 & ~n49739;
  assign n49741 = ~i_FULL & ~n49740;
  assign n49742 = ~n28241 & ~n49741;
  assign n49743 = ~i_nEMPTY & ~n49742;
  assign n49744 = ~n28237 & ~n49743;
  assign n49745 = controllable_BtoS_ACK0 & ~n49744;
  assign n49746 = ~controllable_ENQ & ~n45464;
  assign n49747 = ~n9635 & ~n49746;
  assign n49748 = ~i_RtoB_ACK1 & ~n49747;
  assign n49749 = ~n12462 & ~n49748;
  assign n49750 = controllable_BtoR_REQ1 & ~n49749;
  assign n49751 = ~n9718 & ~n49748;
  assign n49752 = ~controllable_BtoR_REQ1 & ~n49751;
  assign n49753 = ~n49750 & ~n49752;
  assign n49754 = ~controllable_BtoR_REQ0 & ~n49753;
  assign n49755 = ~controllable_BtoR_REQ0 & ~n49754;
  assign n49756 = ~i_RtoB_ACK0 & ~n49755;
  assign n49757 = ~n28175 & ~n49756;
  assign n49758 = ~controllable_DEQ & ~n49757;
  assign n49759 = ~n28224 & ~n49758;
  assign n49760 = ~i_FULL & ~n49759;
  assign n49761 = ~n28570 & ~n49760;
  assign n49762 = ~i_nEMPTY & ~n49761;
  assign n49763 = ~n28566 & ~n49762;
  assign n49764 = ~controllable_BtoS_ACK0 & ~n49763;
  assign n49765 = ~n49745 & ~n49764;
  assign n49766 = n4465 & ~n49765;
  assign n49767 = ~n45990 & ~n49766;
  assign n49768 = i_StoB_REQ10 & ~n49767;
  assign n49769 = ~n49724 & ~n49768;
  assign n49770 = ~controllable_BtoS_ACK10 & ~n49769;
  assign n49771 = ~n49726 & ~n49770;
  assign n49772 = n4464 & ~n49771;
  assign n49773 = ~n45997 & ~n49772;
  assign n49774 = ~n4463 & ~n49773;
  assign n49775 = ~n49464 & ~n49774;
  assign n49776 = n4462 & ~n49775;
  assign n49777 = ~n4462 & ~n28582;
  assign n49778 = ~n49776 & ~n49777;
  assign n49779 = ~n4459 & ~n49778;
  assign n49780 = ~n14759 & ~n18434;
  assign n49781 = i_RtoB_ACK0 & ~n49780;
  assign n49782 = ~controllable_BtoR_REQ1 & ~n49322;
  assign n49783 = ~controllable_BtoR_REQ0 & ~n49782;
  assign n49784 = ~n47037 & ~n49783;
  assign n49785 = ~i_RtoB_ACK0 & ~n49784;
  assign n49786 = ~n49781 & ~n49785;
  assign n49787 = ~controllable_DEQ & ~n49786;
  assign n49788 = ~n14755 & ~n49787;
  assign n49789 = i_nEMPTY & ~n49788;
  assign n49790 = ~n14743 & ~n18428;
  assign n49791 = i_RtoB_ACK0 & ~n49790;
  assign n49792 = ~controllable_BtoR_REQ1 & ~n49332;
  assign n49793 = ~controllable_BtoR_REQ0 & ~n49792;
  assign n49794 = ~n47050 & ~n49793;
  assign n49795 = ~i_RtoB_ACK0 & ~n49794;
  assign n49796 = ~n49791 & ~n49795;
  assign n49797 = ~controllable_DEQ & ~n49796;
  assign n49798 = ~n14780 & ~n49797;
  assign n49799 = i_FULL & ~n49798;
  assign n49800 = ~controllable_BtoR_REQ1 & ~n49342;
  assign n49801 = ~controllable_BtoR_REQ0 & ~n49800;
  assign n49802 = ~n47063 & ~n49801;
  assign n49803 = ~i_RtoB_ACK0 & ~n49802;
  assign n49804 = ~n49791 & ~n49803;
  assign n49805 = ~controllable_DEQ & ~n49804;
  assign n49806 = ~n14798 & ~n49805;
  assign n49807 = ~i_FULL & ~n49806;
  assign n49808 = ~n49799 & ~n49807;
  assign n49809 = ~i_nEMPTY & ~n49808;
  assign n49810 = ~n49789 & ~n49809;
  assign n49811 = controllable_BtoS_ACK0 & ~n49810;
  assign n49812 = ~n18462 & ~n20330;
  assign n49813 = i_RtoB_ACK0 & ~n49812;
  assign n49814 = ~controllable_BtoR_REQ1 & ~n49356;
  assign n49815 = ~controllable_BtoR_REQ0 & ~n49814;
  assign n49816 = ~n47080 & ~n49815;
  assign n49817 = ~i_RtoB_ACK0 & ~n49816;
  assign n49818 = ~n49813 & ~n49817;
  assign n49819 = ~controllable_DEQ & ~n49818;
  assign n49820 = ~n28757 & ~n49819;
  assign n49821 = i_nEMPTY & ~n49820;
  assign n49822 = ~n18456 & ~n20339;
  assign n49823 = i_RtoB_ACK0 & ~n49822;
  assign n49824 = ~controllable_BtoR_REQ1 & ~n49366;
  assign n49825 = ~controllable_BtoR_REQ0 & ~n49824;
  assign n49826 = ~n47093 & ~n49825;
  assign n49827 = ~i_RtoB_ACK0 & ~n49826;
  assign n49828 = ~n49823 & ~n49827;
  assign n49829 = ~controllable_DEQ & ~n49828;
  assign n49830 = ~n28773 & ~n49829;
  assign n49831 = i_FULL & ~n49830;
  assign n49832 = ~controllable_BtoR_REQ1 & ~n49376;
  assign n49833 = ~controllable_BtoR_REQ0 & ~n49832;
  assign n49834 = ~n47106 & ~n49833;
  assign n49835 = ~i_RtoB_ACK0 & ~n49834;
  assign n49836 = ~n49823 & ~n49835;
  assign n49837 = ~controllable_DEQ & ~n49836;
  assign n49838 = ~n28787 & ~n49837;
  assign n49839 = ~i_FULL & ~n49838;
  assign n49840 = ~n49831 & ~n49839;
  assign n49841 = ~i_nEMPTY & ~n49840;
  assign n49842 = ~n49821 & ~n49841;
  assign n49843 = ~controllable_BtoS_ACK0 & ~n49842;
  assign n49844 = ~n49811 & ~n49843;
  assign n49845 = n4465 & ~n49844;
  assign n49846 = ~n47122 & ~n49845;
  assign n49847 = i_StoB_REQ10 & ~n49846;
  assign n49848 = ~n17628 & ~n47128;
  assign n49849 = i_RtoB_ACK0 & ~n49848;
  assign n49850 = ~controllable_BtoR_REQ0 & ~n47253;
  assign n49851 = ~n47134 & ~n49850;
  assign n49852 = ~i_RtoB_ACK0 & ~n49851;
  assign n49853 = ~n49849 & ~n49852;
  assign n49854 = ~controllable_DEQ & ~n49853;
  assign n49855 = ~n17626 & ~n49854;
  assign n49856 = i_nEMPTY & ~n49855;
  assign n49857 = ~n17613 & ~n47147;
  assign n49858 = i_RtoB_ACK0 & ~n49857;
  assign n49859 = ~controllable_BtoR_REQ0 & ~n47260;
  assign n49860 = ~n47153 & ~n49859;
  assign n49861 = ~i_RtoB_ACK0 & ~n49860;
  assign n49862 = ~n49858 & ~n49861;
  assign n49863 = ~controllable_DEQ & ~n49862;
  assign n49864 = ~n17651 & ~n49863;
  assign n49865 = i_FULL & ~n49864;
  assign n49866 = ~n17613 & ~n47166;
  assign n49867 = i_RtoB_ACK0 & ~n49866;
  assign n49868 = ~controllable_BtoR_REQ1 & ~n49410;
  assign n49869 = ~controllable_BtoR_REQ0 & ~n49868;
  assign n49870 = ~n47172 & ~n49869;
  assign n49871 = ~i_RtoB_ACK0 & ~n49870;
  assign n49872 = ~n49867 & ~n49871;
  assign n49873 = ~controllable_DEQ & ~n49872;
  assign n49874 = ~n17673 & ~n49873;
  assign n49875 = ~i_FULL & ~n49874;
  assign n49876 = ~n49865 & ~n49875;
  assign n49877 = ~i_nEMPTY & ~n49876;
  assign n49878 = ~n49856 & ~n49877;
  assign n49879 = controllable_BtoS_ACK0 & ~n49878;
  assign n49880 = ~n17711 & ~n47188;
  assign n49881 = i_RtoB_ACK0 & ~n49880;
  assign n49882 = ~controllable_BtoR_REQ0 & ~n47283;
  assign n49883 = ~n47194 & ~n49882;
  assign n49884 = ~i_RtoB_ACK0 & ~n49883;
  assign n49885 = ~n49881 & ~n49884;
  assign n49886 = ~controllable_DEQ & ~n49885;
  assign n49887 = ~n17705 & ~n49886;
  assign n49888 = i_nEMPTY & ~n49887;
  assign n49889 = ~n17692 & ~n47207;
  assign n49890 = i_RtoB_ACK0 & ~n49889;
  assign n49891 = ~controllable_BtoR_REQ0 & ~n47290;
  assign n49892 = ~n47213 & ~n49891;
  assign n49893 = ~i_RtoB_ACK0 & ~n49892;
  assign n49894 = ~n49890 & ~n49893;
  assign n49895 = ~controllable_DEQ & ~n49894;
  assign n49896 = ~n17741 & ~n49895;
  assign n49897 = i_FULL & ~n49896;
  assign n49898 = ~n17692 & ~n47226;
  assign n49899 = i_RtoB_ACK0 & ~n49898;
  assign n49900 = ~controllable_BtoR_REQ1 & ~n49440;
  assign n49901 = ~controllable_BtoR_REQ0 & ~n49900;
  assign n49902 = ~n47232 & ~n49901;
  assign n49903 = ~i_RtoB_ACK0 & ~n49902;
  assign n49904 = ~n49899 & ~n49903;
  assign n49905 = ~controllable_DEQ & ~n49904;
  assign n49906 = ~n17774 & ~n49905;
  assign n49907 = ~i_FULL & ~n49906;
  assign n49908 = ~n49897 & ~n49907;
  assign n49909 = ~i_nEMPTY & ~n49908;
  assign n49910 = ~n49888 & ~n49909;
  assign n49911 = ~controllable_BtoS_ACK0 & ~n49910;
  assign n49912 = ~n49879 & ~n49911;
  assign n49913 = n4465 & ~n49912;
  assign n49914 = ~n47247 & ~n49913;
  assign n49915 = ~i_StoB_REQ10 & ~n49914;
  assign n49916 = ~n49847 & ~n49915;
  assign n49917 = controllable_BtoS_ACK10 & ~n49916;
  assign n49918 = ~n47316 & ~n49915;
  assign n49919 = ~controllable_BtoS_ACK10 & ~n49918;
  assign n49920 = ~n49917 & ~n49919;
  assign n49921 = n4464 & ~n49920;
  assign n49922 = ~n47321 & ~n49921;
  assign n49923 = n4462 & ~n49922;
  assign n49924 = ~n47324 & ~n49923;
  assign n49925 = n4461 & ~n49924;
  assign n49926 = ~n7111 & ~n12185;
  assign n49927 = ~controllable_BtoR_REQ1 & ~n49926;
  assign n49928 = ~controllable_BtoR_REQ1 & ~n49927;
  assign n49929 = controllable_BtoR_REQ0 & ~n49928;
  assign n49930 = ~controllable_BtoR_REQ1 & ~n49465;
  assign n49931 = ~controllable_BtoR_REQ1 & ~n49930;
  assign n49932 = ~controllable_BtoR_REQ0 & ~n49931;
  assign n49933 = ~n49929 & ~n49932;
  assign n49934 = ~i_RtoB_ACK0 & ~n49933;
  assign n49935 = ~n14761 & ~n49934;
  assign n49936 = ~controllable_DEQ & ~n49935;
  assign n49937 = ~n14755 & ~n49936;
  assign n49938 = i_nEMPTY & ~n49937;
  assign n49939 = ~n7054 & ~n12164;
  assign n49940 = ~controllable_BtoR_REQ1 & ~n49939;
  assign n49941 = ~controllable_BtoR_REQ1 & ~n49940;
  assign n49942 = controllable_BtoR_REQ0 & ~n49941;
  assign n49943 = ~controllable_BtoR_REQ1 & ~n49473;
  assign n49944 = ~controllable_BtoR_REQ1 & ~n49943;
  assign n49945 = ~controllable_BtoR_REQ0 & ~n49944;
  assign n49946 = ~n49942 & ~n49945;
  assign n49947 = ~i_RtoB_ACK0 & ~n49946;
  assign n49948 = ~n14745 & ~n49947;
  assign n49949 = ~controllable_DEQ & ~n49948;
  assign n49950 = ~n14780 & ~n49949;
  assign n49951 = i_FULL & ~n49950;
  assign n49952 = ~n7054 & ~n49482;
  assign n49953 = ~controllable_BtoR_REQ1 & ~n49952;
  assign n49954 = ~controllable_BtoR_REQ1 & ~n49953;
  assign n49955 = controllable_BtoR_REQ0 & ~n49954;
  assign n49956 = ~controllable_BtoR_REQ1 & ~n49483;
  assign n49957 = ~controllable_BtoR_REQ1 & ~n49956;
  assign n49958 = ~controllable_BtoR_REQ0 & ~n49957;
  assign n49959 = ~n49955 & ~n49958;
  assign n49960 = ~i_RtoB_ACK0 & ~n49959;
  assign n49961 = ~n14745 & ~n49960;
  assign n49962 = ~controllable_DEQ & ~n49961;
  assign n49963 = ~n14798 & ~n49962;
  assign n49964 = ~i_FULL & ~n49963;
  assign n49965 = ~n49951 & ~n49964;
  assign n49966 = ~i_nEMPTY & ~n49965;
  assign n49967 = ~n49938 & ~n49966;
  assign n49968 = controllable_BtoS_ACK0 & ~n49967;
  assign n49969 = ~n11324 & ~n12275;
  assign n49970 = ~controllable_BtoR_REQ1 & ~n49969;
  assign n49971 = ~controllable_BtoR_REQ1 & ~n49970;
  assign n49972 = controllable_BtoR_REQ0 & ~n49971;
  assign n49973 = ~controllable_BtoR_REQ1 & ~n49495;
  assign n49974 = ~controllable_BtoR_REQ1 & ~n49973;
  assign n49975 = ~controllable_BtoR_REQ0 & ~n49974;
  assign n49976 = ~n49972 & ~n49975;
  assign n49977 = ~i_RtoB_ACK0 & ~n49976;
  assign n49978 = ~n28739 & ~n49977;
  assign n49979 = ~controllable_DEQ & ~n49978;
  assign n49980 = ~n28757 & ~n49979;
  assign n49981 = i_nEMPTY & ~n49980;
  assign n49982 = ~n11299 & ~n12257;
  assign n49983 = ~controllable_BtoR_REQ1 & ~n49982;
  assign n49984 = ~controllable_BtoR_REQ1 & ~n49983;
  assign n49985 = controllable_BtoR_REQ0 & ~n49984;
  assign n49986 = ~controllable_BtoR_REQ1 & ~n49503;
  assign n49987 = ~controllable_BtoR_REQ1 & ~n49986;
  assign n49988 = ~controllable_BtoR_REQ0 & ~n49987;
  assign n49989 = ~n49985 & ~n49988;
  assign n49990 = ~i_RtoB_ACK0 & ~n49989;
  assign n49991 = ~n28729 & ~n49990;
  assign n49992 = ~controllable_DEQ & ~n49991;
  assign n49993 = ~n28773 & ~n49992;
  assign n49994 = i_FULL & ~n49993;
  assign n49995 = ~n11299 & ~n49512;
  assign n49996 = ~controllable_BtoR_REQ1 & ~n49995;
  assign n49997 = ~controllable_BtoR_REQ1 & ~n49996;
  assign n49998 = controllable_BtoR_REQ0 & ~n49997;
  assign n49999 = ~controllable_BtoR_REQ1 & ~n49513;
  assign n50000 = ~controllable_BtoR_REQ1 & ~n49999;
  assign n50001 = ~controllable_BtoR_REQ0 & ~n50000;
  assign n50002 = ~n49998 & ~n50001;
  assign n50003 = ~i_RtoB_ACK0 & ~n50002;
  assign n50004 = ~n28729 & ~n50003;
  assign n50005 = ~controllable_DEQ & ~n50004;
  assign n50006 = ~n28787 & ~n50005;
  assign n50007 = ~i_FULL & ~n50006;
  assign n50008 = ~n49994 & ~n50007;
  assign n50009 = ~i_nEMPTY & ~n50008;
  assign n50010 = ~n49981 & ~n50009;
  assign n50011 = ~controllable_BtoS_ACK0 & ~n50010;
  assign n50012 = ~n49968 & ~n50011;
  assign n50013 = n4465 & ~n50012;
  assign n50014 = ~n47122 & ~n50013;
  assign n50015 = i_StoB_REQ10 & ~n50014;
  assign n50016 = ~n17631 & ~n46820;
  assign n50017 = ~controllable_BtoR_REQ1 & ~n50016;
  assign n50018 = ~controllable_BtoR_REQ1 & ~n50017;
  assign n50019 = controllable_BtoR_REQ0 & ~n50018;
  assign n50020 = ~controllable_BtoR_REQ1 & ~n49529;
  assign n50021 = ~controllable_BtoR_REQ1 & ~n50020;
  assign n50022 = ~controllable_BtoR_REQ0 & ~n50021;
  assign n50023 = ~n50019 & ~n50022;
  assign n50024 = ~i_RtoB_ACK0 & ~n50023;
  assign n50025 = ~n17630 & ~n50024;
  assign n50026 = ~controllable_DEQ & ~n50025;
  assign n50027 = ~n17626 & ~n50026;
  assign n50028 = i_nEMPTY & ~n50027;
  assign n50029 = ~n17616 & ~n46837;
  assign n50030 = ~controllable_BtoR_REQ1 & ~n50029;
  assign n50031 = ~controllable_BtoR_REQ1 & ~n50030;
  assign n50032 = controllable_BtoR_REQ0 & ~n50031;
  assign n50033 = ~controllable_BtoR_REQ1 & ~n49537;
  assign n50034 = ~controllable_BtoR_REQ1 & ~n50033;
  assign n50035 = ~controllable_BtoR_REQ0 & ~n50034;
  assign n50036 = ~n50032 & ~n50035;
  assign n50037 = ~i_RtoB_ACK0 & ~n50036;
  assign n50038 = ~n17653 & ~n50037;
  assign n50039 = ~controllable_DEQ & ~n50038;
  assign n50040 = ~n17651 & ~n50039;
  assign n50041 = i_FULL & ~n50040;
  assign n50042 = ~n17616 & ~n49659;
  assign n50043 = ~controllable_BtoR_REQ1 & ~n50042;
  assign n50044 = ~controllable_BtoR_REQ1 & ~n50043;
  assign n50045 = controllable_BtoR_REQ0 & ~n50044;
  assign n50046 = ~controllable_BtoR_REQ1 & ~n49663;
  assign n50047 = ~controllable_BtoR_REQ0 & ~n50046;
  assign n50048 = ~n50045 & ~n50047;
  assign n50049 = ~i_RtoB_ACK0 & ~n50048;
  assign n50050 = ~n17615 & ~n50049;
  assign n50051 = ~controllable_DEQ & ~n50050;
  assign n50052 = ~n17673 & ~n50051;
  assign n50053 = ~i_FULL & ~n50052;
  assign n50054 = ~n50041 & ~n50053;
  assign n50055 = ~i_nEMPTY & ~n50054;
  assign n50056 = ~n50028 & ~n50055;
  assign n50057 = controllable_BtoS_ACK0 & ~n50056;
  assign n50058 = ~n17714 & ~n46863;
  assign n50059 = ~controllable_BtoR_REQ1 & ~n50058;
  assign n50060 = ~controllable_BtoR_REQ1 & ~n50059;
  assign n50061 = controllable_BtoR_REQ0 & ~n50060;
  assign n50062 = ~controllable_BtoR_REQ1 & ~n49676;
  assign n50063 = ~controllable_BtoR_REQ1 & ~n50062;
  assign n50064 = ~controllable_BtoR_REQ0 & ~n50063;
  assign n50065 = ~n50061 & ~n50064;
  assign n50066 = ~i_RtoB_ACK0 & ~n50065;
  assign n50067 = ~n17713 & ~n50066;
  assign n50068 = ~controllable_DEQ & ~n50067;
  assign n50069 = ~n17705 & ~n50068;
  assign n50070 = i_nEMPTY & ~n50069;
  assign n50071 = ~n17695 & ~n46880;
  assign n50072 = ~controllable_BtoR_REQ1 & ~n50071;
  assign n50073 = ~controllable_BtoR_REQ1 & ~n50072;
  assign n50074 = controllable_BtoR_REQ0 & ~n50073;
  assign n50075 = ~controllable_BtoR_REQ1 & ~n49684;
  assign n50076 = ~controllable_BtoR_REQ1 & ~n50075;
  assign n50077 = ~controllable_BtoR_REQ0 & ~n50076;
  assign n50078 = ~n50074 & ~n50077;
  assign n50079 = ~i_RtoB_ACK0 & ~n50078;
  assign n50080 = ~n17747 & ~n50079;
  assign n50081 = ~controllable_DEQ & ~n50080;
  assign n50082 = ~n17741 & ~n50081;
  assign n50083 = i_FULL & ~n50082;
  assign n50084 = ~n17695 & ~n49704;
  assign n50085 = ~controllable_BtoR_REQ1 & ~n50084;
  assign n50086 = ~controllable_BtoR_REQ1 & ~n50085;
  assign n50087 = controllable_BtoR_REQ0 & ~n50086;
  assign n50088 = ~controllable_BtoR_REQ1 & ~n49708;
  assign n50089 = ~controllable_BtoR_REQ0 & ~n50088;
  assign n50090 = ~n50087 & ~n50089;
  assign n50091 = ~i_RtoB_ACK0 & ~n50090;
  assign n50092 = ~n17694 & ~n50091;
  assign n50093 = ~controllable_DEQ & ~n50092;
  assign n50094 = ~n17774 & ~n50093;
  assign n50095 = ~i_FULL & ~n50094;
  assign n50096 = ~n50083 & ~n50095;
  assign n50097 = ~i_nEMPTY & ~n50096;
  assign n50098 = ~n50070 & ~n50097;
  assign n50099 = ~controllable_BtoS_ACK0 & ~n50098;
  assign n50100 = ~n50057 & ~n50099;
  assign n50101 = n4465 & ~n50100;
  assign n50102 = ~n47247 & ~n50101;
  assign n50103 = ~i_StoB_REQ10 & ~n50102;
  assign n50104 = ~n50015 & ~n50103;
  assign n50105 = controllable_BtoS_ACK10 & ~n50104;
  assign n50106 = ~controllable_BtoR_REQ1 & ~n49733;
  assign n50107 = ~i_RtoB_ACK0 & ~n50106;
  assign n50108 = ~n29017 & ~n50107;
  assign n50109 = ~controllable_DEQ & ~n50108;
  assign n50110 = ~n29050 & ~n50109;
  assign n50111 = ~i_FULL & ~n50110;
  assign n50112 = ~n29111 & ~n50111;
  assign n50113 = ~i_nEMPTY & ~n50112;
  assign n50114 = ~n29106 & ~n50113;
  assign n50115 = controllable_BtoS_ACK0 & ~n50114;
  assign n50116 = ~controllable_BtoR_REQ1 & ~n49752;
  assign n50117 = ~i_RtoB_ACK0 & ~n50116;
  assign n50118 = ~n29059 & ~n50117;
  assign n50119 = ~controllable_DEQ & ~n50118;
  assign n50120 = ~n29092 & ~n50119;
  assign n50121 = ~i_FULL & ~n50120;
  assign n50122 = ~n29572 & ~n50121;
  assign n50123 = ~i_nEMPTY & ~n50122;
  assign n50124 = ~n29567 & ~n50123;
  assign n50125 = ~controllable_BtoS_ACK0 & ~n50124;
  assign n50126 = ~n50115 & ~n50125;
  assign n50127 = n4465 & ~n50126;
  assign n50128 = ~n47314 & ~n50127;
  assign n50129 = i_StoB_REQ10 & ~n50128;
  assign n50130 = ~n50103 & ~n50129;
  assign n50131 = ~controllable_BtoS_ACK10 & ~n50130;
  assign n50132 = ~n50105 & ~n50131;
  assign n50133 = n4464 & ~n50132;
  assign n50134 = ~n47321 & ~n50133;
  assign n50135 = n4462 & ~n50134;
  assign n50136 = ~n47324 & ~n50135;
  assign n50137 = ~n4461 & ~n50136;
  assign n50138 = ~n49925 & ~n50137;
  assign n50139 = n4459 & ~n50138;
  assign n50140 = ~n49779 & ~n50139;
  assign n50141 = n4455 & ~n50140;
  assign n50142 = ~n5257 & ~n18434;
  assign n50143 = i_RtoB_ACK0 & ~n50142;
  assign n50144 = ~n47037 & ~n49324;
  assign n50145 = ~i_RtoB_ACK0 & ~n50144;
  assign n50146 = ~n50143 & ~n50145;
  assign n50147 = ~controllable_DEQ & ~n50146;
  assign n50148 = ~n20981 & ~n50147;
  assign n50149 = i_nEMPTY & ~n50148;
  assign n50150 = ~n5234 & ~n18428;
  assign n50151 = i_RtoB_ACK0 & ~n50150;
  assign n50152 = ~n47050 & ~n49334;
  assign n50153 = ~i_RtoB_ACK0 & ~n50152;
  assign n50154 = ~n50151 & ~n50153;
  assign n50155 = ~controllable_DEQ & ~n50154;
  assign n50156 = ~n20993 & ~n50155;
  assign n50157 = i_FULL & ~n50156;
  assign n50158 = ~n47063 & ~n49344;
  assign n50159 = ~i_RtoB_ACK0 & ~n50158;
  assign n50160 = ~n50151 & ~n50159;
  assign n50161 = ~controllable_DEQ & ~n50160;
  assign n50162 = ~n21003 & ~n50161;
  assign n50163 = ~i_FULL & ~n50162;
  assign n50164 = ~n50157 & ~n50163;
  assign n50165 = ~i_nEMPTY & ~n50164;
  assign n50166 = ~n50149 & ~n50165;
  assign n50167 = controllable_BtoS_ACK0 & ~n50166;
  assign n50168 = ~n18462 & ~n27869;
  assign n50169 = i_RtoB_ACK0 & ~n50168;
  assign n50170 = ~n47080 & ~n49358;
  assign n50171 = ~i_RtoB_ACK0 & ~n50170;
  assign n50172 = ~n50169 & ~n50171;
  assign n50173 = ~controllable_DEQ & ~n50172;
  assign n50174 = ~n29641 & ~n50173;
  assign n50175 = i_nEMPTY & ~n50174;
  assign n50176 = ~n18456 & ~n27857;
  assign n50177 = i_RtoB_ACK0 & ~n50176;
  assign n50178 = ~n47093 & ~n49368;
  assign n50179 = ~i_RtoB_ACK0 & ~n50178;
  assign n50180 = ~n50177 & ~n50179;
  assign n50181 = ~controllable_DEQ & ~n50180;
  assign n50182 = ~n29653 & ~n50181;
  assign n50183 = i_FULL & ~n50182;
  assign n50184 = ~n47106 & ~n49378;
  assign n50185 = ~i_RtoB_ACK0 & ~n50184;
  assign n50186 = ~n50177 & ~n50185;
  assign n50187 = ~controllable_DEQ & ~n50186;
  assign n50188 = ~n29663 & ~n50187;
  assign n50189 = ~i_FULL & ~n50188;
  assign n50190 = ~n50183 & ~n50189;
  assign n50191 = ~i_nEMPTY & ~n50190;
  assign n50192 = ~n50175 & ~n50191;
  assign n50193 = ~controllable_BtoS_ACK0 & ~n50192;
  assign n50194 = ~n50167 & ~n50193;
  assign n50195 = n4465 & ~n50194;
  assign n50196 = ~n48393 & ~n50195;
  assign n50197 = i_StoB_REQ10 & ~n50196;
  assign n50198 = ~n11250 & ~n47128;
  assign n50199 = i_RtoB_ACK0 & ~n50198;
  assign n50200 = ~n47134 & ~n49394;
  assign n50201 = ~i_RtoB_ACK0 & ~n50200;
  assign n50202 = ~n50199 & ~n50201;
  assign n50203 = ~controllable_DEQ & ~n50202;
  assign n50204 = ~n23093 & ~n50203;
  assign n50205 = i_nEMPTY & ~n50204;
  assign n50206 = ~n11232 & ~n47147;
  assign n50207 = i_RtoB_ACK0 & ~n50206;
  assign n50208 = ~n47153 & ~n49402;
  assign n50209 = ~i_RtoB_ACK0 & ~n50208;
  assign n50210 = ~n50207 & ~n50209;
  assign n50211 = ~controllable_DEQ & ~n50210;
  assign n50212 = ~n23105 & ~n50211;
  assign n50213 = i_FULL & ~n50212;
  assign n50214 = ~n11232 & ~n47166;
  assign n50215 = i_RtoB_ACK0 & ~n50214;
  assign n50216 = ~n47172 & ~n49412;
  assign n50217 = ~i_RtoB_ACK0 & ~n50216;
  assign n50218 = ~n50215 & ~n50217;
  assign n50219 = ~controllable_DEQ & ~n50218;
  assign n50220 = ~n23117 & ~n50219;
  assign n50221 = ~i_FULL & ~n50220;
  assign n50222 = ~n50213 & ~n50221;
  assign n50223 = ~i_nEMPTY & ~n50222;
  assign n50224 = ~n50205 & ~n50223;
  assign n50225 = controllable_BtoS_ACK0 & ~n50224;
  assign n50226 = ~n11330 & ~n47188;
  assign n50227 = i_RtoB_ACK0 & ~n50226;
  assign n50228 = ~n47194 & ~n49424;
  assign n50229 = ~i_RtoB_ACK0 & ~n50228;
  assign n50230 = ~n50227 & ~n50229;
  assign n50231 = ~controllable_DEQ & ~n50230;
  assign n50232 = ~n23133 & ~n50231;
  assign n50233 = i_nEMPTY & ~n50232;
  assign n50234 = ~n11307 & ~n47207;
  assign n50235 = i_RtoB_ACK0 & ~n50234;
  assign n50236 = ~n47213 & ~n49432;
  assign n50237 = ~i_RtoB_ACK0 & ~n50236;
  assign n50238 = ~n50235 & ~n50237;
  assign n50239 = ~controllable_DEQ & ~n50238;
  assign n50240 = ~n23145 & ~n50239;
  assign n50241 = i_FULL & ~n50240;
  assign n50242 = ~n11307 & ~n47226;
  assign n50243 = i_RtoB_ACK0 & ~n50242;
  assign n50244 = ~n47232 & ~n49442;
  assign n50245 = ~i_RtoB_ACK0 & ~n50244;
  assign n50246 = ~n50243 & ~n50245;
  assign n50247 = ~controllable_DEQ & ~n50246;
  assign n50248 = ~n23157 & ~n50247;
  assign n50249 = ~i_FULL & ~n50248;
  assign n50250 = ~n50241 & ~n50249;
  assign n50251 = ~i_nEMPTY & ~n50250;
  assign n50252 = ~n50233 & ~n50251;
  assign n50253 = ~controllable_BtoS_ACK0 & ~n50252;
  assign n50254 = ~n50225 & ~n50253;
  assign n50255 = n4465 & ~n50254;
  assign n50256 = ~n48454 & ~n50255;
  assign n50257 = ~i_StoB_REQ10 & ~n50256;
  assign n50258 = ~n50197 & ~n50257;
  assign n50259 = controllable_BtoS_ACK10 & ~n50258;
  assign n50260 = ~n48511 & ~n50257;
  assign n50261 = ~controllable_BtoS_ACK10 & ~n50260;
  assign n50262 = ~n50259 & ~n50261;
  assign n50263 = n4464 & ~n50262;
  assign n50264 = ~n48516 & ~n50263;
  assign n50265 = n4463 & ~n50264;
  assign n50266 = ~n47037 & ~n49466;
  assign n50267 = ~i_RtoB_ACK0 & ~n50266;
  assign n50268 = ~n50143 & ~n50267;
  assign n50269 = ~controllable_DEQ & ~n50268;
  assign n50270 = ~n20981 & ~n50269;
  assign n50271 = i_nEMPTY & ~n50270;
  assign n50272 = ~n47050 & ~n49474;
  assign n50273 = ~i_RtoB_ACK0 & ~n50272;
  assign n50274 = ~n50151 & ~n50273;
  assign n50275 = ~controllable_DEQ & ~n50274;
  assign n50276 = ~n20993 & ~n50275;
  assign n50277 = i_FULL & ~n50276;
  assign n50278 = ~n47063 & ~n49484;
  assign n50279 = ~i_RtoB_ACK0 & ~n50278;
  assign n50280 = ~n50151 & ~n50279;
  assign n50281 = ~controllable_DEQ & ~n50280;
  assign n50282 = ~n21003 & ~n50281;
  assign n50283 = ~i_FULL & ~n50282;
  assign n50284 = ~n50277 & ~n50283;
  assign n50285 = ~i_nEMPTY & ~n50284;
  assign n50286 = ~n50271 & ~n50285;
  assign n50287 = controllable_BtoS_ACK0 & ~n50286;
  assign n50288 = ~n47080 & ~n49496;
  assign n50289 = ~i_RtoB_ACK0 & ~n50288;
  assign n50290 = ~n50169 & ~n50289;
  assign n50291 = ~controllable_DEQ & ~n50290;
  assign n50292 = ~n29641 & ~n50291;
  assign n50293 = i_nEMPTY & ~n50292;
  assign n50294 = ~n47093 & ~n49504;
  assign n50295 = ~i_RtoB_ACK0 & ~n50294;
  assign n50296 = ~n50177 & ~n50295;
  assign n50297 = ~controllable_DEQ & ~n50296;
  assign n50298 = ~n29653 & ~n50297;
  assign n50299 = i_FULL & ~n50298;
  assign n50300 = ~n47106 & ~n49514;
  assign n50301 = ~i_RtoB_ACK0 & ~n50300;
  assign n50302 = ~n50177 & ~n50301;
  assign n50303 = ~controllable_DEQ & ~n50302;
  assign n50304 = ~n29663 & ~n50303;
  assign n50305 = ~i_FULL & ~n50304;
  assign n50306 = ~n50299 & ~n50305;
  assign n50307 = ~i_nEMPTY & ~n50306;
  assign n50308 = ~n50293 & ~n50307;
  assign n50309 = ~controllable_BtoS_ACK0 & ~n50308;
  assign n50310 = ~n50287 & ~n50309;
  assign n50311 = n4465 & ~n50310;
  assign n50312 = ~n48393 & ~n50311;
  assign n50313 = i_StoB_REQ10 & ~n50312;
  assign n50314 = ~n47134 & ~n49530;
  assign n50315 = ~i_RtoB_ACK0 & ~n50314;
  assign n50316 = ~n50199 & ~n50315;
  assign n50317 = ~controllable_DEQ & ~n50316;
  assign n50318 = ~n23093 & ~n50317;
  assign n50319 = i_nEMPTY & ~n50318;
  assign n50320 = ~n47153 & ~n49538;
  assign n50321 = ~i_RtoB_ACK0 & ~n50320;
  assign n50322 = ~n50207 & ~n50321;
  assign n50323 = ~controllable_DEQ & ~n50322;
  assign n50324 = ~n23105 & ~n50323;
  assign n50325 = i_FULL & ~n50324;
  assign n50326 = ~n47172 & ~n49665;
  assign n50327 = ~i_RtoB_ACK0 & ~n50326;
  assign n50328 = ~n50215 & ~n50327;
  assign n50329 = ~controllable_DEQ & ~n50328;
  assign n50330 = ~n23117 & ~n50329;
  assign n50331 = ~i_FULL & ~n50330;
  assign n50332 = ~n50325 & ~n50331;
  assign n50333 = ~i_nEMPTY & ~n50332;
  assign n50334 = ~n50319 & ~n50333;
  assign n50335 = controllable_BtoS_ACK0 & ~n50334;
  assign n50336 = ~n47194 & ~n49677;
  assign n50337 = ~i_RtoB_ACK0 & ~n50336;
  assign n50338 = ~n50227 & ~n50337;
  assign n50339 = ~controllable_DEQ & ~n50338;
  assign n50340 = ~n23133 & ~n50339;
  assign n50341 = i_nEMPTY & ~n50340;
  assign n50342 = ~n47213 & ~n49685;
  assign n50343 = ~i_RtoB_ACK0 & ~n50342;
  assign n50344 = ~n50235 & ~n50343;
  assign n50345 = ~controllable_DEQ & ~n50344;
  assign n50346 = ~n23145 & ~n50345;
  assign n50347 = i_FULL & ~n50346;
  assign n50348 = ~n47232 & ~n49710;
  assign n50349 = ~i_RtoB_ACK0 & ~n50348;
  assign n50350 = ~n50243 & ~n50349;
  assign n50351 = ~controllable_DEQ & ~n50350;
  assign n50352 = ~n23157 & ~n50351;
  assign n50353 = ~i_FULL & ~n50352;
  assign n50354 = ~n50347 & ~n50353;
  assign n50355 = ~i_nEMPTY & ~n50354;
  assign n50356 = ~n50341 & ~n50355;
  assign n50357 = ~controllable_BtoS_ACK0 & ~n50356;
  assign n50358 = ~n50335 & ~n50357;
  assign n50359 = n4465 & ~n50358;
  assign n50360 = ~n48454 & ~n50359;
  assign n50361 = ~i_StoB_REQ10 & ~n50360;
  assign n50362 = ~n50313 & ~n50361;
  assign n50363 = controllable_BtoS_ACK10 & ~n50362;
  assign n50364 = ~n11253 & ~n48193;
  assign n50365 = ~i_RtoB_ACK0 & ~n50364;
  assign n50366 = ~n29832 & ~n50365;
  assign n50367 = ~controllable_DEQ & ~n50366;
  assign n50368 = ~n29844 & ~n50367;
  assign n50369 = i_nEMPTY & ~n50368;
  assign n50370 = ~n11270 & ~n48210;
  assign n50371 = ~i_RtoB_ACK0 & ~n50370;
  assign n50372 = ~n29860 & ~n50371;
  assign n50373 = ~controllable_DEQ & ~n50372;
  assign n50374 = ~n29858 & ~n50373;
  assign n50375 = i_FULL & ~n50374;
  assign n50376 = ~n48219 & ~n49735;
  assign n50377 = ~i_RtoB_ACK0 & ~n50376;
  assign n50378 = ~n48472 & ~n50377;
  assign n50379 = ~controllable_DEQ & ~n50378;
  assign n50380 = ~n29872 & ~n50379;
  assign n50381 = ~i_FULL & ~n50380;
  assign n50382 = ~n50375 & ~n50381;
  assign n50383 = ~i_nEMPTY & ~n50382;
  assign n50384 = ~n50369 & ~n50383;
  assign n50385 = controllable_BtoS_ACK0 & ~n50384;
  assign n50386 = ~n11333 & ~n48232;
  assign n50387 = ~i_RtoB_ACK0 & ~n50386;
  assign n50388 = ~n29888 & ~n50387;
  assign n50389 = ~controllable_DEQ & ~n50388;
  assign n50390 = ~n29900 & ~n50389;
  assign n50391 = i_nEMPTY & ~n50390;
  assign n50392 = ~n11352 & ~n48249;
  assign n50393 = ~i_RtoB_ACK0 & ~n50392;
  assign n50394 = ~n29916 & ~n50393;
  assign n50395 = ~controllable_DEQ & ~n50394;
  assign n50396 = ~n29914 & ~n50395;
  assign n50397 = i_FULL & ~n50396;
  assign n50398 = ~n48258 & ~n49754;
  assign n50399 = ~i_RtoB_ACK0 & ~n50398;
  assign n50400 = ~n48496 & ~n50399;
  assign n50401 = ~controllable_DEQ & ~n50400;
  assign n50402 = ~n29928 & ~n50401;
  assign n50403 = ~i_FULL & ~n50402;
  assign n50404 = ~n50397 & ~n50403;
  assign n50405 = ~i_nEMPTY & ~n50404;
  assign n50406 = ~n50391 & ~n50405;
  assign n50407 = ~controllable_BtoS_ACK0 & ~n50406;
  assign n50408 = ~n50385 & ~n50407;
  assign n50409 = n4465 & ~n50408;
  assign n50410 = ~n48509 & ~n50409;
  assign n50411 = i_StoB_REQ10 & ~n50410;
  assign n50412 = ~n50361 & ~n50411;
  assign n50413 = ~controllable_BtoS_ACK10 & ~n50412;
  assign n50414 = ~n50363 & ~n50413;
  assign n50415 = n4464 & ~n50414;
  assign n50416 = ~n48516 & ~n50415;
  assign n50417 = ~n4463 & ~n50416;
  assign n50418 = ~n50265 & ~n50417;
  assign n50419 = n4462 & ~n50418;
  assign n50420 = ~n4462 & ~n31547;
  assign n50421 = ~n50419 & ~n50420;
  assign n50422 = n4461 & ~n50421;
  assign n50423 = ~n49324 & ~n49929;
  assign n50424 = ~i_RtoB_ACK0 & ~n50423;
  assign n50425 = ~n20983 & ~n50424;
  assign n50426 = ~controllable_DEQ & ~n50425;
  assign n50427 = ~n20981 & ~n50426;
  assign n50428 = i_nEMPTY & ~n50427;
  assign n50429 = ~n49334 & ~n49942;
  assign n50430 = ~i_RtoB_ACK0 & ~n50429;
  assign n50431 = ~n20977 & ~n50430;
  assign n50432 = ~controllable_DEQ & ~n50431;
  assign n50433 = ~n20993 & ~n50432;
  assign n50434 = i_FULL & ~n50433;
  assign n50435 = ~n49344 & ~n49955;
  assign n50436 = ~i_RtoB_ACK0 & ~n50435;
  assign n50437 = ~n20977 & ~n50436;
  assign n50438 = ~controllable_DEQ & ~n50437;
  assign n50439 = ~n21003 & ~n50438;
  assign n50440 = ~i_FULL & ~n50439;
  assign n50441 = ~n50434 & ~n50440;
  assign n50442 = ~i_nEMPTY & ~n50441;
  assign n50443 = ~n50428 & ~n50442;
  assign n50444 = controllable_BtoS_ACK0 & ~n50443;
  assign n50445 = ~n49358 & ~n49972;
  assign n50446 = ~i_RtoB_ACK0 & ~n50445;
  assign n50447 = ~n29631 & ~n50446;
  assign n50448 = ~controllable_DEQ & ~n50447;
  assign n50449 = ~n29641 & ~n50448;
  assign n50450 = i_nEMPTY & ~n50449;
  assign n50451 = ~n49368 & ~n49985;
  assign n50452 = ~i_RtoB_ACK0 & ~n50451;
  assign n50453 = ~n29625 & ~n50452;
  assign n50454 = ~controllable_DEQ & ~n50453;
  assign n50455 = ~n29653 & ~n50454;
  assign n50456 = i_FULL & ~n50455;
  assign n50457 = ~n49378 & ~n49998;
  assign n50458 = ~i_RtoB_ACK0 & ~n50457;
  assign n50459 = ~n29625 & ~n50458;
  assign n50460 = ~controllable_DEQ & ~n50459;
  assign n50461 = ~n29663 & ~n50460;
  assign n50462 = ~i_FULL & ~n50461;
  assign n50463 = ~n50456 & ~n50462;
  assign n50464 = ~i_nEMPTY & ~n50463;
  assign n50465 = ~n50450 & ~n50464;
  assign n50466 = ~controllable_BtoS_ACK0 & ~n50465;
  assign n50467 = ~n50444 & ~n50466;
  assign n50468 = n4465 & ~n50467;
  assign n50469 = ~n48393 & ~n50468;
  assign n50470 = i_StoB_REQ10 & ~n50469;
  assign n50471 = ~n49394 & ~n50019;
  assign n50472 = ~i_RtoB_ACK0 & ~n50471;
  assign n50473 = ~n23095 & ~n50472;
  assign n50474 = ~controllable_DEQ & ~n50473;
  assign n50475 = ~n23093 & ~n50474;
  assign n50476 = i_nEMPTY & ~n50475;
  assign n50477 = ~n49402 & ~n50032;
  assign n50478 = ~i_RtoB_ACK0 & ~n50477;
  assign n50479 = ~n23107 & ~n50478;
  assign n50480 = ~controllable_DEQ & ~n50479;
  assign n50481 = ~n23105 & ~n50480;
  assign n50482 = i_FULL & ~n50481;
  assign n50483 = ~n49412 & ~n50045;
  assign n50484 = ~i_RtoB_ACK0 & ~n50483;
  assign n50485 = ~n23089 & ~n50484;
  assign n50486 = ~controllable_DEQ & ~n50485;
  assign n50487 = ~n23117 & ~n50486;
  assign n50488 = ~i_FULL & ~n50487;
  assign n50489 = ~n50482 & ~n50488;
  assign n50490 = ~i_nEMPTY & ~n50489;
  assign n50491 = ~n50476 & ~n50490;
  assign n50492 = controllable_BtoS_ACK0 & ~n50491;
  assign n50493 = ~n49424 & ~n50061;
  assign n50494 = ~i_RtoB_ACK0 & ~n50493;
  assign n50495 = ~n23135 & ~n50494;
  assign n50496 = ~controllable_DEQ & ~n50495;
  assign n50497 = ~n23133 & ~n50496;
  assign n50498 = i_nEMPTY & ~n50497;
  assign n50499 = ~n49432 & ~n50074;
  assign n50500 = ~i_RtoB_ACK0 & ~n50499;
  assign n50501 = ~n23147 & ~n50500;
  assign n50502 = ~controllable_DEQ & ~n50501;
  assign n50503 = ~n23145 & ~n50502;
  assign n50504 = i_FULL & ~n50503;
  assign n50505 = ~n49442 & ~n50087;
  assign n50506 = ~i_RtoB_ACK0 & ~n50505;
  assign n50507 = ~n23129 & ~n50506;
  assign n50508 = ~controllable_DEQ & ~n50507;
  assign n50509 = ~n23157 & ~n50508;
  assign n50510 = ~i_FULL & ~n50509;
  assign n50511 = ~n50504 & ~n50510;
  assign n50512 = ~i_nEMPTY & ~n50511;
  assign n50513 = ~n50498 & ~n50512;
  assign n50514 = ~controllable_BtoS_ACK0 & ~n50513;
  assign n50515 = ~n50492 & ~n50514;
  assign n50516 = n4465 & ~n50515;
  assign n50517 = ~n48454 & ~n50516;
  assign n50518 = ~i_StoB_REQ10 & ~n50517;
  assign n50519 = ~n50470 & ~n50518;
  assign n50520 = controllable_BtoS_ACK10 & ~n50519;
  assign n50521 = ~n29938 & ~n45925;
  assign n50522 = ~i_RtoB_ACK0 & ~n50521;
  assign n50523 = ~n29832 & ~n50522;
  assign n50524 = ~controllable_DEQ & ~n50523;
  assign n50525 = ~n29844 & ~n50524;
  assign n50526 = i_nEMPTY & ~n50525;
  assign n50527 = ~n29945 & ~n45933;
  assign n50528 = ~i_RtoB_ACK0 & ~n50527;
  assign n50529 = ~n29860 & ~n50528;
  assign n50530 = ~controllable_DEQ & ~n50529;
  assign n50531 = ~n29858 & ~n50530;
  assign n50532 = i_FULL & ~n50531;
  assign n50533 = controllable_BtoR_REQ0 & ~n50106;
  assign n50534 = ~n45945 & ~n50533;
  assign n50535 = ~i_RtoB_ACK0 & ~n50534;
  assign n50536 = ~n29825 & ~n50535;
  assign n50537 = ~controllable_DEQ & ~n50536;
  assign n50538 = ~n29872 & ~n50537;
  assign n50539 = ~i_FULL & ~n50538;
  assign n50540 = ~n50532 & ~n50539;
  assign n50541 = ~i_nEMPTY & ~n50540;
  assign n50542 = ~n50526 & ~n50541;
  assign n50543 = controllable_BtoS_ACK0 & ~n50542;
  assign n50544 = ~n31230 & ~n45957;
  assign n50545 = ~i_RtoB_ACK0 & ~n50544;
  assign n50546 = ~n29888 & ~n50545;
  assign n50547 = ~controllable_DEQ & ~n50546;
  assign n50548 = ~n29900 & ~n50547;
  assign n50549 = i_nEMPTY & ~n50548;
  assign n50550 = ~n31245 & ~n45965;
  assign n50551 = ~i_RtoB_ACK0 & ~n50550;
  assign n50552 = ~n29916 & ~n50551;
  assign n50553 = ~controllable_DEQ & ~n50552;
  assign n50554 = ~n29914 & ~n50553;
  assign n50555 = i_FULL & ~n50554;
  assign n50556 = controllable_BtoR_REQ0 & ~n50116;
  assign n50557 = ~n45977 & ~n50556;
  assign n50558 = ~i_RtoB_ACK0 & ~n50557;
  assign n50559 = ~n29881 & ~n50558;
  assign n50560 = ~controllable_DEQ & ~n50559;
  assign n50561 = ~n29928 & ~n50560;
  assign n50562 = ~i_FULL & ~n50561;
  assign n50563 = ~n50555 & ~n50562;
  assign n50564 = ~i_nEMPTY & ~n50563;
  assign n50565 = ~n50549 & ~n50564;
  assign n50566 = ~controllable_BtoS_ACK0 & ~n50565;
  assign n50567 = ~n50543 & ~n50566;
  assign n50568 = n4465 & ~n50567;
  assign n50569 = ~n48509 & ~n50568;
  assign n50570 = i_StoB_REQ10 & ~n50569;
  assign n50571 = ~n50518 & ~n50570;
  assign n50572 = ~controllable_BtoS_ACK10 & ~n50571;
  assign n50573 = ~n50520 & ~n50572;
  assign n50574 = n4464 & ~n50573;
  assign n50575 = ~n48516 & ~n50574;
  assign n50576 = n4463 & ~n50575;
  assign n50577 = ~n49466 & ~n49929;
  assign n50578 = ~i_RtoB_ACK0 & ~n50577;
  assign n50579 = ~n20983 & ~n50578;
  assign n50580 = ~controllable_DEQ & ~n50579;
  assign n50581 = ~n20981 & ~n50580;
  assign n50582 = i_nEMPTY & ~n50581;
  assign n50583 = ~n49474 & ~n49942;
  assign n50584 = ~i_RtoB_ACK0 & ~n50583;
  assign n50585 = ~n20977 & ~n50584;
  assign n50586 = ~controllable_DEQ & ~n50585;
  assign n50587 = ~n20993 & ~n50586;
  assign n50588 = i_FULL & ~n50587;
  assign n50589 = ~n49484 & ~n49955;
  assign n50590 = ~i_RtoB_ACK0 & ~n50589;
  assign n50591 = ~n20977 & ~n50590;
  assign n50592 = ~controllable_DEQ & ~n50591;
  assign n50593 = ~n21003 & ~n50592;
  assign n50594 = ~i_FULL & ~n50593;
  assign n50595 = ~n50588 & ~n50594;
  assign n50596 = ~i_nEMPTY & ~n50595;
  assign n50597 = ~n50582 & ~n50596;
  assign n50598 = controllable_BtoS_ACK0 & ~n50597;
  assign n50599 = ~n49496 & ~n49972;
  assign n50600 = ~i_RtoB_ACK0 & ~n50599;
  assign n50601 = ~n29631 & ~n50600;
  assign n50602 = ~controllable_DEQ & ~n50601;
  assign n50603 = ~n29641 & ~n50602;
  assign n50604 = i_nEMPTY & ~n50603;
  assign n50605 = ~n49504 & ~n49985;
  assign n50606 = ~i_RtoB_ACK0 & ~n50605;
  assign n50607 = ~n29625 & ~n50606;
  assign n50608 = ~controllable_DEQ & ~n50607;
  assign n50609 = ~n29653 & ~n50608;
  assign n50610 = i_FULL & ~n50609;
  assign n50611 = ~n49514 & ~n49998;
  assign n50612 = ~i_RtoB_ACK0 & ~n50611;
  assign n50613 = ~n29625 & ~n50612;
  assign n50614 = ~controllable_DEQ & ~n50613;
  assign n50615 = ~n29663 & ~n50614;
  assign n50616 = ~i_FULL & ~n50615;
  assign n50617 = ~n50610 & ~n50616;
  assign n50618 = ~i_nEMPTY & ~n50617;
  assign n50619 = ~n50604 & ~n50618;
  assign n50620 = ~controllable_BtoS_ACK0 & ~n50619;
  assign n50621 = ~n50598 & ~n50620;
  assign n50622 = n4465 & ~n50621;
  assign n50623 = ~n48393 & ~n50622;
  assign n50624 = i_StoB_REQ10 & ~n50623;
  assign n50625 = ~n49530 & ~n50019;
  assign n50626 = ~i_RtoB_ACK0 & ~n50625;
  assign n50627 = ~n23095 & ~n50626;
  assign n50628 = ~controllable_DEQ & ~n50627;
  assign n50629 = ~n23093 & ~n50628;
  assign n50630 = i_nEMPTY & ~n50629;
  assign n50631 = ~n49538 & ~n50032;
  assign n50632 = ~i_RtoB_ACK0 & ~n50631;
  assign n50633 = ~n23107 & ~n50632;
  assign n50634 = ~controllable_DEQ & ~n50633;
  assign n50635 = ~n23105 & ~n50634;
  assign n50636 = i_FULL & ~n50635;
  assign n50637 = ~n49665 & ~n50045;
  assign n50638 = ~i_RtoB_ACK0 & ~n50637;
  assign n50639 = ~n23089 & ~n50638;
  assign n50640 = ~controllable_DEQ & ~n50639;
  assign n50641 = ~n23117 & ~n50640;
  assign n50642 = ~i_FULL & ~n50641;
  assign n50643 = ~n50636 & ~n50642;
  assign n50644 = ~i_nEMPTY & ~n50643;
  assign n50645 = ~n50630 & ~n50644;
  assign n50646 = controllable_BtoS_ACK0 & ~n50645;
  assign n50647 = ~n49677 & ~n50061;
  assign n50648 = ~i_RtoB_ACK0 & ~n50647;
  assign n50649 = ~n23135 & ~n50648;
  assign n50650 = ~controllable_DEQ & ~n50649;
  assign n50651 = ~n23133 & ~n50650;
  assign n50652 = i_nEMPTY & ~n50651;
  assign n50653 = ~n49685 & ~n50074;
  assign n50654 = ~i_RtoB_ACK0 & ~n50653;
  assign n50655 = ~n23147 & ~n50654;
  assign n50656 = ~controllable_DEQ & ~n50655;
  assign n50657 = ~n23145 & ~n50656;
  assign n50658 = i_FULL & ~n50657;
  assign n50659 = ~n49710 & ~n50087;
  assign n50660 = ~i_RtoB_ACK0 & ~n50659;
  assign n50661 = ~n23129 & ~n50660;
  assign n50662 = ~controllable_DEQ & ~n50661;
  assign n50663 = ~n23157 & ~n50662;
  assign n50664 = ~i_FULL & ~n50663;
  assign n50665 = ~n50658 & ~n50664;
  assign n50666 = ~i_nEMPTY & ~n50665;
  assign n50667 = ~n50652 & ~n50666;
  assign n50668 = ~controllable_BtoS_ACK0 & ~n50667;
  assign n50669 = ~n50646 & ~n50668;
  assign n50670 = n4465 & ~n50669;
  assign n50671 = ~n48454 & ~n50670;
  assign n50672 = ~i_StoB_REQ10 & ~n50671;
  assign n50673 = ~n50624 & ~n50672;
  assign n50674 = controllable_BtoS_ACK10 & ~n50673;
  assign n50675 = ~n49735 & ~n50533;
  assign n50676 = ~i_RtoB_ACK0 & ~n50675;
  assign n50677 = ~n29825 & ~n50676;
  assign n50678 = ~controllable_DEQ & ~n50677;
  assign n50679 = ~n29872 & ~n50678;
  assign n50680 = ~i_FULL & ~n50679;
  assign n50681 = ~n29951 & ~n50680;
  assign n50682 = ~i_nEMPTY & ~n50681;
  assign n50683 = ~n29944 & ~n50682;
  assign n50684 = controllable_BtoS_ACK0 & ~n50683;
  assign n50685 = ~n49754 & ~n50556;
  assign n50686 = ~i_RtoB_ACK0 & ~n50685;
  assign n50687 = ~n29881 & ~n50686;
  assign n50688 = ~controllable_DEQ & ~n50687;
  assign n50689 = ~n29928 & ~n50688;
  assign n50690 = ~i_FULL & ~n50689;
  assign n50691 = ~n31535 & ~n50690;
  assign n50692 = ~i_nEMPTY & ~n50691;
  assign n50693 = ~n31529 & ~n50692;
  assign n50694 = ~controllable_BtoS_ACK0 & ~n50693;
  assign n50695 = ~n50684 & ~n50694;
  assign n50696 = n4465 & ~n50695;
  assign n50697 = ~n48509 & ~n50696;
  assign n50698 = i_StoB_REQ10 & ~n50697;
  assign n50699 = ~n50672 & ~n50698;
  assign n50700 = ~controllable_BtoS_ACK10 & ~n50699;
  assign n50701 = ~n50674 & ~n50700;
  assign n50702 = n4464 & ~n50701;
  assign n50703 = ~n48516 & ~n50702;
  assign n50704 = ~n4463 & ~n50703;
  assign n50705 = ~n50576 & ~n50704;
  assign n50706 = n4462 & ~n50705;
  assign n50707 = ~n50420 & ~n50706;
  assign n50708 = ~n4461 & ~n50707;
  assign n50709 = ~n50422 & ~n50708;
  assign n50710 = ~n4459 & ~n50709;
  assign n50711 = controllable_BtoR_REQ1 & ~n49465;
  assign n50712 = ~n49322 & ~n50711;
  assign n50713 = ~controllable_BtoR_REQ0 & ~n50712;
  assign n50714 = ~n47037 & ~n50713;
  assign n50715 = ~i_RtoB_ACK0 & ~n50714;
  assign n50716 = ~n50143 & ~n50715;
  assign n50717 = ~controllable_DEQ & ~n50716;
  assign n50718 = ~n20981 & ~n50717;
  assign n50719 = i_nEMPTY & ~n50718;
  assign n50720 = controllable_BtoR_REQ1 & ~n49473;
  assign n50721 = ~n49332 & ~n50720;
  assign n50722 = ~controllable_BtoR_REQ0 & ~n50721;
  assign n50723 = ~n47050 & ~n50722;
  assign n50724 = ~i_RtoB_ACK0 & ~n50723;
  assign n50725 = ~n50151 & ~n50724;
  assign n50726 = ~controllable_DEQ & ~n50725;
  assign n50727 = ~n20993 & ~n50726;
  assign n50728 = i_FULL & ~n50727;
  assign n50729 = controllable_BtoR_REQ1 & ~n49483;
  assign n50730 = ~n49342 & ~n50729;
  assign n50731 = ~controllable_BtoR_REQ0 & ~n50730;
  assign n50732 = ~n47063 & ~n50731;
  assign n50733 = ~i_RtoB_ACK0 & ~n50732;
  assign n50734 = ~n50151 & ~n50733;
  assign n50735 = ~controllable_DEQ & ~n50734;
  assign n50736 = ~n21003 & ~n50735;
  assign n50737 = ~i_FULL & ~n50736;
  assign n50738 = ~n50728 & ~n50737;
  assign n50739 = ~i_nEMPTY & ~n50738;
  assign n50740 = ~n50719 & ~n50739;
  assign n50741 = controllable_BtoS_ACK0 & ~n50740;
  assign n50742 = controllable_BtoR_REQ1 & ~n49495;
  assign n50743 = ~n49356 & ~n50742;
  assign n50744 = ~controllable_BtoR_REQ0 & ~n50743;
  assign n50745 = ~n47080 & ~n50744;
  assign n50746 = ~i_RtoB_ACK0 & ~n50745;
  assign n50747 = ~n50169 & ~n50746;
  assign n50748 = ~controllable_DEQ & ~n50747;
  assign n50749 = ~n29641 & ~n50748;
  assign n50750 = i_nEMPTY & ~n50749;
  assign n50751 = controllable_BtoR_REQ1 & ~n49503;
  assign n50752 = ~n49366 & ~n50751;
  assign n50753 = ~controllable_BtoR_REQ0 & ~n50752;
  assign n50754 = ~n47093 & ~n50753;
  assign n50755 = ~i_RtoB_ACK0 & ~n50754;
  assign n50756 = ~n50177 & ~n50755;
  assign n50757 = ~controllable_DEQ & ~n50756;
  assign n50758 = ~n29653 & ~n50757;
  assign n50759 = i_FULL & ~n50758;
  assign n50760 = controllable_BtoR_REQ1 & ~n49513;
  assign n50761 = ~n49376 & ~n50760;
  assign n50762 = ~controllable_BtoR_REQ0 & ~n50761;
  assign n50763 = ~n47106 & ~n50762;
  assign n50764 = ~i_RtoB_ACK0 & ~n50763;
  assign n50765 = ~n50177 & ~n50764;
  assign n50766 = ~controllable_DEQ & ~n50765;
  assign n50767 = ~n29663 & ~n50766;
  assign n50768 = ~i_FULL & ~n50767;
  assign n50769 = ~n50759 & ~n50768;
  assign n50770 = ~i_nEMPTY & ~n50769;
  assign n50771 = ~n50750 & ~n50770;
  assign n50772 = ~controllable_BtoS_ACK0 & ~n50771;
  assign n50773 = ~n50741 & ~n50772;
  assign n50774 = n4465 & ~n50773;
  assign n50775 = ~n48393 & ~n50774;
  assign n50776 = i_StoB_REQ10 & ~n50775;
  assign n50777 = controllable_BtoR_REQ1 & ~n49529;
  assign n50778 = ~n47252 & ~n50777;
  assign n50779 = ~controllable_BtoR_REQ0 & ~n50778;
  assign n50780 = ~n47134 & ~n50779;
  assign n50781 = ~i_RtoB_ACK0 & ~n50780;
  assign n50782 = ~n50199 & ~n50781;
  assign n50783 = ~controllable_DEQ & ~n50782;
  assign n50784 = ~n23093 & ~n50783;
  assign n50785 = i_nEMPTY & ~n50784;
  assign n50786 = controllable_BtoR_REQ1 & ~n49537;
  assign n50787 = ~n47259 & ~n50786;
  assign n50788 = ~controllable_BtoR_REQ0 & ~n50787;
  assign n50789 = ~n47153 & ~n50788;
  assign n50790 = ~i_RtoB_ACK0 & ~n50789;
  assign n50791 = ~n50207 & ~n50790;
  assign n50792 = ~controllable_DEQ & ~n50791;
  assign n50793 = ~n23105 & ~n50792;
  assign n50794 = i_FULL & ~n50793;
  assign n50795 = ~n49410 & ~n49661;
  assign n50796 = ~controllable_BtoR_REQ0 & ~n50795;
  assign n50797 = ~n47172 & ~n50796;
  assign n50798 = ~i_RtoB_ACK0 & ~n50797;
  assign n50799 = ~n50215 & ~n50798;
  assign n50800 = ~controllable_DEQ & ~n50799;
  assign n50801 = ~n23117 & ~n50800;
  assign n50802 = ~i_FULL & ~n50801;
  assign n50803 = ~n50794 & ~n50802;
  assign n50804 = ~i_nEMPTY & ~n50803;
  assign n50805 = ~n50785 & ~n50804;
  assign n50806 = controllable_BtoS_ACK0 & ~n50805;
  assign n50807 = controllable_BtoR_REQ1 & ~n49676;
  assign n50808 = ~n47282 & ~n50807;
  assign n50809 = ~controllable_BtoR_REQ0 & ~n50808;
  assign n50810 = ~n47194 & ~n50809;
  assign n50811 = ~i_RtoB_ACK0 & ~n50810;
  assign n50812 = ~n50227 & ~n50811;
  assign n50813 = ~controllable_DEQ & ~n50812;
  assign n50814 = ~n23133 & ~n50813;
  assign n50815 = i_nEMPTY & ~n50814;
  assign n50816 = controllable_BtoR_REQ1 & ~n49684;
  assign n50817 = ~n47289 & ~n50816;
  assign n50818 = ~controllable_BtoR_REQ0 & ~n50817;
  assign n50819 = ~n47213 & ~n50818;
  assign n50820 = ~i_RtoB_ACK0 & ~n50819;
  assign n50821 = ~n50235 & ~n50820;
  assign n50822 = ~controllable_DEQ & ~n50821;
  assign n50823 = ~n23145 & ~n50822;
  assign n50824 = i_FULL & ~n50823;
  assign n50825 = ~n49440 & ~n49706;
  assign n50826 = ~controllable_BtoR_REQ0 & ~n50825;
  assign n50827 = ~n47232 & ~n50826;
  assign n50828 = ~i_RtoB_ACK0 & ~n50827;
  assign n50829 = ~n50243 & ~n50828;
  assign n50830 = ~controllable_DEQ & ~n50829;
  assign n50831 = ~n23157 & ~n50830;
  assign n50832 = ~i_FULL & ~n50831;
  assign n50833 = ~n50824 & ~n50832;
  assign n50834 = ~i_nEMPTY & ~n50833;
  assign n50835 = ~n50815 & ~n50834;
  assign n50836 = ~controllable_BtoS_ACK0 & ~n50835;
  assign n50837 = ~n50806 & ~n50836;
  assign n50838 = n4465 & ~n50837;
  assign n50839 = ~n48454 & ~n50838;
  assign n50840 = ~i_StoB_REQ10 & ~n50839;
  assign n50841 = ~n50776 & ~n50840;
  assign n50842 = controllable_BtoS_ACK10 & ~n50841;
  assign n50843 = ~n31786 & ~n47252;
  assign n50844 = ~controllable_BtoR_REQ0 & ~n50843;
  assign n50845 = ~n48193 & ~n50844;
  assign n50846 = ~i_RtoB_ACK0 & ~n50845;
  assign n50847 = ~n29832 & ~n50846;
  assign n50848 = ~controllable_DEQ & ~n50847;
  assign n50849 = ~n29844 & ~n50848;
  assign n50850 = i_nEMPTY & ~n50849;
  assign n50851 = ~n31805 & ~n47259;
  assign n50852 = ~controllable_BtoR_REQ0 & ~n50851;
  assign n50853 = ~n48210 & ~n50852;
  assign n50854 = ~i_RtoB_ACK0 & ~n50853;
  assign n50855 = ~n29860 & ~n50854;
  assign n50856 = ~controllable_DEQ & ~n50855;
  assign n50857 = ~n29858 & ~n50856;
  assign n50858 = i_FULL & ~n50857;
  assign n50859 = ~n45943 & ~n49731;
  assign n50860 = ~controllable_BtoR_REQ0 & ~n50859;
  assign n50861 = ~n48219 & ~n50860;
  assign n50862 = ~i_RtoB_ACK0 & ~n50861;
  assign n50863 = ~n48472 & ~n50862;
  assign n50864 = ~controllable_DEQ & ~n50863;
  assign n50865 = ~n29872 & ~n50864;
  assign n50866 = ~i_FULL & ~n50865;
  assign n50867 = ~n50858 & ~n50866;
  assign n50868 = ~i_nEMPTY & ~n50867;
  assign n50869 = ~n50850 & ~n50868;
  assign n50870 = controllable_BtoS_ACK0 & ~n50869;
  assign n50871 = ~n31832 & ~n47282;
  assign n50872 = ~controllable_BtoR_REQ0 & ~n50871;
  assign n50873 = ~n48232 & ~n50872;
  assign n50874 = ~i_RtoB_ACK0 & ~n50873;
  assign n50875 = ~n29888 & ~n50874;
  assign n50876 = ~controllable_DEQ & ~n50875;
  assign n50877 = ~n29900 & ~n50876;
  assign n50878 = i_nEMPTY & ~n50877;
  assign n50879 = ~n31851 & ~n47289;
  assign n50880 = ~controllable_BtoR_REQ0 & ~n50879;
  assign n50881 = ~n48249 & ~n50880;
  assign n50882 = ~i_RtoB_ACK0 & ~n50881;
  assign n50883 = ~n29916 & ~n50882;
  assign n50884 = ~controllable_DEQ & ~n50883;
  assign n50885 = ~n29914 & ~n50884;
  assign n50886 = i_FULL & ~n50885;
  assign n50887 = ~n45975 & ~n49750;
  assign n50888 = ~controllable_BtoR_REQ0 & ~n50887;
  assign n50889 = ~n48258 & ~n50888;
  assign n50890 = ~i_RtoB_ACK0 & ~n50889;
  assign n50891 = ~n48496 & ~n50890;
  assign n50892 = ~controllable_DEQ & ~n50891;
  assign n50893 = ~n29928 & ~n50892;
  assign n50894 = ~i_FULL & ~n50893;
  assign n50895 = ~n50886 & ~n50894;
  assign n50896 = ~i_nEMPTY & ~n50895;
  assign n50897 = ~n50878 & ~n50896;
  assign n50898 = ~controllable_BtoS_ACK0 & ~n50897;
  assign n50899 = ~n50870 & ~n50898;
  assign n50900 = n4465 & ~n50899;
  assign n50901 = ~n48509 & ~n50900;
  assign n50902 = i_StoB_REQ10 & ~n50901;
  assign n50903 = ~n50840 & ~n50902;
  assign n50904 = ~controllable_BtoS_ACK10 & ~n50903;
  assign n50905 = ~n50842 & ~n50904;
  assign n50906 = n4464 & ~n50905;
  assign n50907 = ~n48516 & ~n50906;
  assign n50908 = ~n4463 & ~n50907;
  assign n50909 = ~n50265 & ~n50908;
  assign n50910 = n4462 & ~n50909;
  assign n50911 = ~n50420 & ~n50910;
  assign n50912 = n4461 & ~n50911;
  assign n50913 = ~n48555 & ~n49930;
  assign n50914 = ~controllable_BtoR_REQ0 & ~n50913;
  assign n50915 = ~n49929 & ~n50914;
  assign n50916 = ~i_RtoB_ACK0 & ~n50915;
  assign n50917 = ~n20983 & ~n50916;
  assign n50918 = ~controllable_DEQ & ~n50917;
  assign n50919 = ~n20981 & ~n50918;
  assign n50920 = i_nEMPTY & ~n50919;
  assign n50921 = ~n48574 & ~n49943;
  assign n50922 = ~controllable_BtoR_REQ0 & ~n50921;
  assign n50923 = ~n49942 & ~n50922;
  assign n50924 = ~i_RtoB_ACK0 & ~n50923;
  assign n50925 = ~n20977 & ~n50924;
  assign n50926 = ~controllable_DEQ & ~n50925;
  assign n50927 = ~n20993 & ~n50926;
  assign n50928 = i_FULL & ~n50927;
  assign n50929 = ~n48583 & ~n49956;
  assign n50930 = ~controllable_BtoR_REQ0 & ~n50929;
  assign n50931 = ~n49955 & ~n50930;
  assign n50932 = ~i_RtoB_ACK0 & ~n50931;
  assign n50933 = ~n20977 & ~n50932;
  assign n50934 = ~controllable_DEQ & ~n50933;
  assign n50935 = ~n21003 & ~n50934;
  assign n50936 = ~i_FULL & ~n50935;
  assign n50937 = ~n50928 & ~n50936;
  assign n50938 = ~i_nEMPTY & ~n50937;
  assign n50939 = ~n50920 & ~n50938;
  assign n50940 = controllable_BtoS_ACK0 & ~n50939;
  assign n50941 = ~n48596 & ~n49973;
  assign n50942 = ~controllable_BtoR_REQ0 & ~n50941;
  assign n50943 = ~n49972 & ~n50942;
  assign n50944 = ~i_RtoB_ACK0 & ~n50943;
  assign n50945 = ~n29631 & ~n50944;
  assign n50946 = ~controllable_DEQ & ~n50945;
  assign n50947 = ~n29641 & ~n50946;
  assign n50948 = i_nEMPTY & ~n50947;
  assign n50949 = ~n48615 & ~n49986;
  assign n50950 = ~controllable_BtoR_REQ0 & ~n50949;
  assign n50951 = ~n49985 & ~n50950;
  assign n50952 = ~i_RtoB_ACK0 & ~n50951;
  assign n50953 = ~n29625 & ~n50952;
  assign n50954 = ~controllable_DEQ & ~n50953;
  assign n50955 = ~n29653 & ~n50954;
  assign n50956 = i_FULL & ~n50955;
  assign n50957 = ~n48624 & ~n49999;
  assign n50958 = ~controllable_BtoR_REQ0 & ~n50957;
  assign n50959 = ~n49998 & ~n50958;
  assign n50960 = ~i_RtoB_ACK0 & ~n50959;
  assign n50961 = ~n29625 & ~n50960;
  assign n50962 = ~controllable_DEQ & ~n50961;
  assign n50963 = ~n29663 & ~n50962;
  assign n50964 = ~i_FULL & ~n50963;
  assign n50965 = ~n50956 & ~n50964;
  assign n50966 = ~i_nEMPTY & ~n50965;
  assign n50967 = ~n50948 & ~n50966;
  assign n50968 = ~controllable_BtoS_ACK0 & ~n50967;
  assign n50969 = ~n50940 & ~n50968;
  assign n50970 = n4465 & ~n50969;
  assign n50971 = ~n48393 & ~n50970;
  assign n50972 = i_StoB_REQ10 & ~n50971;
  assign n50973 = ~n48649 & ~n50020;
  assign n50974 = ~controllable_BtoR_REQ0 & ~n50973;
  assign n50975 = ~n50019 & ~n50974;
  assign n50976 = ~i_RtoB_ACK0 & ~n50975;
  assign n50977 = ~n23095 & ~n50976;
  assign n50978 = ~controllable_DEQ & ~n50977;
  assign n50979 = ~n23093 & ~n50978;
  assign n50980 = i_nEMPTY & ~n50979;
  assign n50981 = ~n48668 & ~n50033;
  assign n50982 = ~controllable_BtoR_REQ0 & ~n50981;
  assign n50983 = ~n50032 & ~n50982;
  assign n50984 = ~i_RtoB_ACK0 & ~n50983;
  assign n50985 = ~n23107 & ~n50984;
  assign n50986 = ~controllable_DEQ & ~n50985;
  assign n50987 = ~n23105 & ~n50986;
  assign n50988 = i_FULL & ~n50987;
  assign n50989 = ~n45858 & ~n49663;
  assign n50990 = ~controllable_BtoR_REQ0 & ~n50989;
  assign n50991 = ~n50045 & ~n50990;
  assign n50992 = ~i_RtoB_ACK0 & ~n50991;
  assign n50993 = ~n23089 & ~n50992;
  assign n50994 = ~controllable_DEQ & ~n50993;
  assign n50995 = ~n23117 & ~n50994;
  assign n50996 = ~i_FULL & ~n50995;
  assign n50997 = ~n50988 & ~n50996;
  assign n50998 = ~i_nEMPTY & ~n50997;
  assign n50999 = ~n50980 & ~n50998;
  assign n51000 = controllable_BtoS_ACK0 & ~n50999;
  assign n51001 = ~n48689 & ~n50062;
  assign n51002 = ~controllable_BtoR_REQ0 & ~n51001;
  assign n51003 = ~n50061 & ~n51002;
  assign n51004 = ~i_RtoB_ACK0 & ~n51003;
  assign n51005 = ~n23135 & ~n51004;
  assign n51006 = ~controllable_DEQ & ~n51005;
  assign n51007 = ~n23133 & ~n51006;
  assign n51008 = i_nEMPTY & ~n51007;
  assign n51009 = ~n48708 & ~n50075;
  assign n51010 = ~controllable_BtoR_REQ0 & ~n51009;
  assign n51011 = ~n50074 & ~n51010;
  assign n51012 = ~i_RtoB_ACK0 & ~n51011;
  assign n51013 = ~n23147 & ~n51012;
  assign n51014 = ~controllable_DEQ & ~n51013;
  assign n51015 = ~n23145 & ~n51014;
  assign n51016 = i_FULL & ~n51015;
  assign n51017 = ~n45902 & ~n49708;
  assign n51018 = ~controllable_BtoR_REQ0 & ~n51017;
  assign n51019 = ~n50087 & ~n51018;
  assign n51020 = ~i_RtoB_ACK0 & ~n51019;
  assign n51021 = ~n23129 & ~n51020;
  assign n51022 = ~controllable_DEQ & ~n51021;
  assign n51023 = ~n23157 & ~n51022;
  assign n51024 = ~i_FULL & ~n51023;
  assign n51025 = ~n51016 & ~n51024;
  assign n51026 = ~i_nEMPTY & ~n51025;
  assign n51027 = ~n51008 & ~n51026;
  assign n51028 = ~controllable_BtoS_ACK0 & ~n51027;
  assign n51029 = ~n51000 & ~n51028;
  assign n51030 = n4465 & ~n51029;
  assign n51031 = ~n48454 & ~n51030;
  assign n51032 = ~i_StoB_REQ10 & ~n51031;
  assign n51033 = ~n50972 & ~n51032;
  assign n51034 = controllable_BtoS_ACK10 & ~n51033;
  assign n51035 = ~n11248 & ~n48743;
  assign n51036 = ~controllable_BtoR_REQ0 & ~n51035;
  assign n51037 = ~n29938 & ~n51036;
  assign n51038 = ~i_RtoB_ACK0 & ~n51037;
  assign n51039 = ~n29832 & ~n51038;
  assign n51040 = ~controllable_DEQ & ~n51039;
  assign n51041 = ~n29844 & ~n51040;
  assign n51042 = i_nEMPTY & ~n51041;
  assign n51043 = ~n11230 & ~n48762;
  assign n51044 = ~controllable_BtoR_REQ0 & ~n51043;
  assign n51045 = ~n29945 & ~n51044;
  assign n51046 = ~i_RtoB_ACK0 & ~n51045;
  assign n51047 = ~n29860 & ~n51046;
  assign n51048 = ~controllable_DEQ & ~n51047;
  assign n51049 = ~n29858 & ~n51048;
  assign n51050 = i_FULL & ~n51049;
  assign n51051 = ~n45941 & ~n49733;
  assign n51052 = ~controllable_BtoR_REQ0 & ~n51051;
  assign n51053 = ~n50533 & ~n51052;
  assign n51054 = ~i_RtoB_ACK0 & ~n51053;
  assign n51055 = ~n29825 & ~n51054;
  assign n51056 = ~controllable_DEQ & ~n51055;
  assign n51057 = ~n29872 & ~n51056;
  assign n51058 = ~i_FULL & ~n51057;
  assign n51059 = ~n51050 & ~n51058;
  assign n51060 = ~i_nEMPTY & ~n51059;
  assign n51061 = ~n51042 & ~n51060;
  assign n51062 = controllable_BtoS_ACK0 & ~n51061;
  assign n51063 = ~n11328 & ~n48783;
  assign n51064 = ~controllable_BtoR_REQ0 & ~n51063;
  assign n51065 = ~n31230 & ~n51064;
  assign n51066 = ~i_RtoB_ACK0 & ~n51065;
  assign n51067 = ~n29888 & ~n51066;
  assign n51068 = ~controllable_DEQ & ~n51067;
  assign n51069 = ~n29900 & ~n51068;
  assign n51070 = i_nEMPTY & ~n51069;
  assign n51071 = ~n11305 & ~n48802;
  assign n51072 = ~controllable_BtoR_REQ0 & ~n51071;
  assign n51073 = ~n31245 & ~n51072;
  assign n51074 = ~i_RtoB_ACK0 & ~n51073;
  assign n51075 = ~n29916 & ~n51074;
  assign n51076 = ~controllable_DEQ & ~n51075;
  assign n51077 = ~n29914 & ~n51076;
  assign n51078 = i_FULL & ~n51077;
  assign n51079 = ~n45973 & ~n49752;
  assign n51080 = ~controllable_BtoR_REQ0 & ~n51079;
  assign n51081 = ~n50556 & ~n51080;
  assign n51082 = ~i_RtoB_ACK0 & ~n51081;
  assign n51083 = ~n29881 & ~n51082;
  assign n51084 = ~controllable_DEQ & ~n51083;
  assign n51085 = ~n29928 & ~n51084;
  assign n51086 = ~i_FULL & ~n51085;
  assign n51087 = ~n51078 & ~n51086;
  assign n51088 = ~i_nEMPTY & ~n51087;
  assign n51089 = ~n51070 & ~n51088;
  assign n51090 = ~controllable_BtoS_ACK0 & ~n51089;
  assign n51091 = ~n51062 & ~n51090;
  assign n51092 = n4465 & ~n51091;
  assign n51093 = ~n48509 & ~n51092;
  assign n51094 = i_StoB_REQ10 & ~n51093;
  assign n51095 = ~n51032 & ~n51094;
  assign n51096 = ~controllable_BtoS_ACK10 & ~n51095;
  assign n51097 = ~n51034 & ~n51096;
  assign n51098 = n4464 & ~n51097;
  assign n51099 = ~n48516 & ~n51098;
  assign n51100 = n4463 & ~n51099;
  assign n51101 = ~n50704 & ~n51100;
  assign n51102 = n4462 & ~n51101;
  assign n51103 = ~n50420 & ~n51102;
  assign n51104 = ~n4461 & ~n51103;
  assign n51105 = ~n50912 & ~n51104;
  assign n51106 = n4459 & ~n51105;
  assign n51107 = ~n50710 & ~n51106;
  assign n51108 = ~n4455 & ~n51107;
  assign n51109 = ~n50141 & ~n51108;
  assign n51110 = n4445 & ~n51109;
  assign n51111 = n4463 & ~n49773;
  assign n51112 = ~n28583 & ~n51111;
  assign n51113 = n4462 & ~n51112;
  assign n51114 = ~n49777 & ~n51113;
  assign n51115 = ~n4459 & ~n51114;
  assign n51116 = n4461 & ~n50136;
  assign n51117 = ~n29585 & ~n51116;
  assign n51118 = n4459 & ~n51117;
  assign n51119 = ~n51115 & ~n51118;
  assign n51120 = n4455 & ~n51119;
  assign n51121 = n4463 & ~n50703;
  assign n51122 = ~n5260 & ~n49929;
  assign n51123 = ~i_RtoB_ACK0 & ~n51122;
  assign n51124 = ~n20983 & ~n51123;
  assign n51125 = ~controllable_DEQ & ~n51124;
  assign n51126 = ~n20981 & ~n51125;
  assign n51127 = i_nEMPTY & ~n51126;
  assign n51128 = ~n5282 & ~n49942;
  assign n51129 = ~i_RtoB_ACK0 & ~n51128;
  assign n51130 = ~n20977 & ~n51129;
  assign n51131 = ~controllable_DEQ & ~n51130;
  assign n51132 = ~n20993 & ~n51131;
  assign n51133 = i_FULL & ~n51132;
  assign n51134 = ~n5297 & ~n49955;
  assign n51135 = ~i_RtoB_ACK0 & ~n51134;
  assign n51136 = ~n20977 & ~n51135;
  assign n51137 = ~controllable_DEQ & ~n51136;
  assign n51138 = ~n21003 & ~n51137;
  assign n51139 = ~i_FULL & ~n51138;
  assign n51140 = ~n51133 & ~n51139;
  assign n51141 = ~i_nEMPTY & ~n51140;
  assign n51142 = ~n51127 & ~n51141;
  assign n51143 = controllable_BtoS_ACK0 & ~n51142;
  assign n51144 = ~n28534 & ~n49972;
  assign n51145 = ~i_RtoB_ACK0 & ~n51144;
  assign n51146 = ~n29631 & ~n51145;
  assign n51147 = ~controllable_DEQ & ~n51146;
  assign n51148 = ~n29641 & ~n51147;
  assign n51149 = i_nEMPTY & ~n51148;
  assign n51150 = ~n28541 & ~n49985;
  assign n51151 = ~i_RtoB_ACK0 & ~n51150;
  assign n51152 = ~n29625 & ~n51151;
  assign n51153 = ~controllable_DEQ & ~n51152;
  assign n51154 = ~n29653 & ~n51153;
  assign n51155 = i_FULL & ~n51154;
  assign n51156 = ~n28548 & ~n49998;
  assign n51157 = ~i_RtoB_ACK0 & ~n51156;
  assign n51158 = ~n29625 & ~n51157;
  assign n51159 = ~controllable_DEQ & ~n51158;
  assign n51160 = ~n29663 & ~n51159;
  assign n51161 = ~i_FULL & ~n51160;
  assign n51162 = ~n51155 & ~n51161;
  assign n51163 = ~i_nEMPTY & ~n51162;
  assign n51164 = ~n51149 & ~n51163;
  assign n51165 = ~controllable_BtoS_ACK0 & ~n51164;
  assign n51166 = ~n51143 & ~n51165;
  assign n51167 = n4465 & ~n51166;
  assign n51168 = ~n48393 & ~n51167;
  assign n51169 = i_StoB_REQ10 & ~n51168;
  assign n51170 = ~n11253 & ~n50019;
  assign n51171 = ~i_RtoB_ACK0 & ~n51170;
  assign n51172 = ~n23095 & ~n51171;
  assign n51173 = ~controllable_DEQ & ~n51172;
  assign n51174 = ~n23093 & ~n51173;
  assign n51175 = i_nEMPTY & ~n51174;
  assign n51176 = ~n11270 & ~n50032;
  assign n51177 = ~i_RtoB_ACK0 & ~n51176;
  assign n51178 = ~n23107 & ~n51177;
  assign n51179 = ~controllable_DEQ & ~n51178;
  assign n51180 = ~n23105 & ~n51179;
  assign n51181 = i_FULL & ~n51180;
  assign n51182 = ~n11286 & ~n50045;
  assign n51183 = ~i_RtoB_ACK0 & ~n51182;
  assign n51184 = ~n23089 & ~n51183;
  assign n51185 = ~controllable_DEQ & ~n51184;
  assign n51186 = ~n23117 & ~n51185;
  assign n51187 = ~i_FULL & ~n51186;
  assign n51188 = ~n51181 & ~n51187;
  assign n51189 = ~i_nEMPTY & ~n51188;
  assign n51190 = ~n51175 & ~n51189;
  assign n51191 = controllable_BtoS_ACK0 & ~n51190;
  assign n51192 = ~n11333 & ~n50061;
  assign n51193 = ~i_RtoB_ACK0 & ~n51192;
  assign n51194 = ~n23135 & ~n51193;
  assign n51195 = ~controllable_DEQ & ~n51194;
  assign n51196 = ~n23133 & ~n51195;
  assign n51197 = i_nEMPTY & ~n51196;
  assign n51198 = ~n11352 & ~n50074;
  assign n51199 = ~i_RtoB_ACK0 & ~n51198;
  assign n51200 = ~n23147 & ~n51199;
  assign n51201 = ~controllable_DEQ & ~n51200;
  assign n51202 = ~n23145 & ~n51201;
  assign n51203 = i_FULL & ~n51202;
  assign n51204 = ~n11368 & ~n50087;
  assign n51205 = ~i_RtoB_ACK0 & ~n51204;
  assign n51206 = ~n23129 & ~n51205;
  assign n51207 = ~controllable_DEQ & ~n51206;
  assign n51208 = ~n23157 & ~n51207;
  assign n51209 = ~i_FULL & ~n51208;
  assign n51210 = ~n51203 & ~n51209;
  assign n51211 = ~i_nEMPTY & ~n51210;
  assign n51212 = ~n51197 & ~n51211;
  assign n51213 = ~controllable_BtoS_ACK0 & ~n51212;
  assign n51214 = ~n51191 & ~n51213;
  assign n51215 = n4465 & ~n51214;
  assign n51216 = ~n48454 & ~n51215;
  assign n51217 = ~i_StoB_REQ10 & ~n51216;
  assign n51218 = ~n51169 & ~n51217;
  assign n51219 = controllable_BtoS_ACK10 & ~n51218;
  assign n51220 = ~n28135 & ~n50533;
  assign n51221 = ~i_RtoB_ACK0 & ~n51220;
  assign n51222 = ~n29825 & ~n51221;
  assign n51223 = ~controllable_DEQ & ~n51222;
  assign n51224 = ~n29872 & ~n51223;
  assign n51225 = ~i_FULL & ~n51224;
  assign n51226 = ~n29951 & ~n51225;
  assign n51227 = ~i_nEMPTY & ~n51226;
  assign n51228 = ~n29944 & ~n51227;
  assign n51229 = controllable_BtoS_ACK0 & ~n51228;
  assign n51230 = ~n28196 & ~n50556;
  assign n51231 = ~i_RtoB_ACK0 & ~n51230;
  assign n51232 = ~n29881 & ~n51231;
  assign n51233 = ~controllable_DEQ & ~n51232;
  assign n51234 = ~n29928 & ~n51233;
  assign n51235 = ~i_FULL & ~n51234;
  assign n51236 = ~n31535 & ~n51235;
  assign n51237 = ~i_nEMPTY & ~n51236;
  assign n51238 = ~n31529 & ~n51237;
  assign n51239 = ~controllable_BtoS_ACK0 & ~n51238;
  assign n51240 = ~n51229 & ~n51239;
  assign n51241 = n4465 & ~n51240;
  assign n51242 = ~n48509 & ~n51241;
  assign n51243 = i_StoB_REQ10 & ~n51242;
  assign n51244 = ~n51217 & ~n51243;
  assign n51245 = ~controllable_BtoS_ACK10 & ~n51244;
  assign n51246 = ~n51219 & ~n51245;
  assign n51247 = n4464 & ~n51246;
  assign n51248 = ~n48516 & ~n51247;
  assign n51249 = ~n4463 & ~n51248;
  assign n51250 = ~n51121 & ~n51249;
  assign n51251 = n4462 & ~n51250;
  assign n51252 = ~n50420 & ~n51251;
  assign n51253 = n4461 & ~n51252;
  assign n51254 = ~n14765 & ~n49466;
  assign n51255 = ~i_RtoB_ACK0 & ~n51254;
  assign n51256 = ~n20983 & ~n51255;
  assign n51257 = ~controllable_DEQ & ~n51256;
  assign n51258 = ~n20981 & ~n51257;
  assign n51259 = i_nEMPTY & ~n51258;
  assign n51260 = ~n14784 & ~n49474;
  assign n51261 = ~i_RtoB_ACK0 & ~n51260;
  assign n51262 = ~n20977 & ~n51261;
  assign n51263 = ~controllable_DEQ & ~n51262;
  assign n51264 = ~n20993 & ~n51263;
  assign n51265 = i_FULL & ~n51264;
  assign n51266 = ~n14749 & ~n49484;
  assign n51267 = ~i_RtoB_ACK0 & ~n51266;
  assign n51268 = ~n20977 & ~n51267;
  assign n51269 = ~controllable_DEQ & ~n51268;
  assign n51270 = ~n21003 & ~n51269;
  assign n51271 = ~i_FULL & ~n51270;
  assign n51272 = ~n51265 & ~n51271;
  assign n51273 = ~i_nEMPTY & ~n51272;
  assign n51274 = ~n51259 & ~n51273;
  assign n51275 = controllable_BtoS_ACK0 & ~n51274;
  assign n51276 = ~n29437 & ~n49496;
  assign n51277 = ~i_RtoB_ACK0 & ~n51276;
  assign n51278 = ~n29631 & ~n51277;
  assign n51279 = ~controllable_DEQ & ~n51278;
  assign n51280 = ~n29641 & ~n51279;
  assign n51281 = i_nEMPTY & ~n51280;
  assign n51282 = ~n29447 & ~n49504;
  assign n51283 = ~i_RtoB_ACK0 & ~n51282;
  assign n51284 = ~n29625 & ~n51283;
  assign n51285 = ~controllable_DEQ & ~n51284;
  assign n51286 = ~n29653 & ~n51285;
  assign n51287 = i_FULL & ~n51286;
  assign n51288 = ~n28753 & ~n49514;
  assign n51289 = ~i_RtoB_ACK0 & ~n51288;
  assign n51290 = ~n29625 & ~n51289;
  assign n51291 = ~controllable_DEQ & ~n51290;
  assign n51292 = ~n29663 & ~n51291;
  assign n51293 = ~i_FULL & ~n51292;
  assign n51294 = ~n51287 & ~n51293;
  assign n51295 = ~i_nEMPTY & ~n51294;
  assign n51296 = ~n51281 & ~n51295;
  assign n51297 = ~controllable_BtoS_ACK0 & ~n51296;
  assign n51298 = ~n51275 & ~n51297;
  assign n51299 = n4465 & ~n51298;
  assign n51300 = ~n48393 & ~n51299;
  assign n51301 = i_StoB_REQ10 & ~n51300;
  assign n51302 = ~n17635 & ~n49530;
  assign n51303 = ~i_RtoB_ACK0 & ~n51302;
  assign n51304 = ~n23095 & ~n51303;
  assign n51305 = ~controllable_DEQ & ~n51304;
  assign n51306 = ~n23093 & ~n51305;
  assign n51307 = i_nEMPTY & ~n51306;
  assign n51308 = ~n17657 & ~n49538;
  assign n51309 = ~i_RtoB_ACK0 & ~n51308;
  assign n51310 = ~n23107 & ~n51309;
  assign n51311 = ~controllable_DEQ & ~n51310;
  assign n51312 = ~n23105 & ~n51311;
  assign n51313 = i_FULL & ~n51312;
  assign n51314 = ~n17620 & ~n49665;
  assign n51315 = ~i_RtoB_ACK0 & ~n51314;
  assign n51316 = ~n23089 & ~n51315;
  assign n51317 = ~controllable_DEQ & ~n51316;
  assign n51318 = ~n23117 & ~n51317;
  assign n51319 = ~i_FULL & ~n51318;
  assign n51320 = ~n51313 & ~n51319;
  assign n51321 = ~i_nEMPTY & ~n51320;
  assign n51322 = ~n51307 & ~n51321;
  assign n51323 = controllable_BtoS_ACK0 & ~n51322;
  assign n51324 = ~n17718 & ~n49677;
  assign n51325 = ~i_RtoB_ACK0 & ~n51324;
  assign n51326 = ~n23135 & ~n51325;
  assign n51327 = ~controllable_DEQ & ~n51326;
  assign n51328 = ~n23133 & ~n51327;
  assign n51329 = i_nEMPTY & ~n51328;
  assign n51330 = ~n17751 & ~n49685;
  assign n51331 = ~i_RtoB_ACK0 & ~n51330;
  assign n51332 = ~n23147 & ~n51331;
  assign n51333 = ~controllable_DEQ & ~n51332;
  assign n51334 = ~n23145 & ~n51333;
  assign n51335 = i_FULL & ~n51334;
  assign n51336 = ~n17699 & ~n49710;
  assign n51337 = ~i_RtoB_ACK0 & ~n51336;
  assign n51338 = ~n23129 & ~n51337;
  assign n51339 = ~controllable_DEQ & ~n51338;
  assign n51340 = ~n23157 & ~n51339;
  assign n51341 = ~i_FULL & ~n51340;
  assign n51342 = ~n51335 & ~n51341;
  assign n51343 = ~i_nEMPTY & ~n51342;
  assign n51344 = ~n51329 & ~n51343;
  assign n51345 = ~controllable_BtoS_ACK0 & ~n51344;
  assign n51346 = ~n51323 & ~n51345;
  assign n51347 = n4465 & ~n51346;
  assign n51348 = ~n48454 & ~n51347;
  assign n51349 = ~i_StoB_REQ10 & ~n51348;
  assign n51350 = ~n51301 & ~n51349;
  assign n51351 = controllable_BtoS_ACK10 & ~n51350;
  assign n51352 = ~n29840 & ~n49735;
  assign n51353 = ~i_RtoB_ACK0 & ~n51352;
  assign n51354 = ~n29825 & ~n51353;
  assign n51355 = ~controllable_DEQ & ~n51354;
  assign n51356 = ~n29872 & ~n51355;
  assign n51357 = ~i_FULL & ~n51356;
  assign n51358 = ~n29951 & ~n51357;
  assign n51359 = ~i_nEMPTY & ~n51358;
  assign n51360 = ~n29944 & ~n51359;
  assign n51361 = controllable_BtoS_ACK0 & ~n51360;
  assign n51362 = ~n29896 & ~n49754;
  assign n51363 = ~i_RtoB_ACK0 & ~n51362;
  assign n51364 = ~n29881 & ~n51363;
  assign n51365 = ~controllable_DEQ & ~n51364;
  assign n51366 = ~n29928 & ~n51365;
  assign n51367 = ~i_FULL & ~n51366;
  assign n51368 = ~n31535 & ~n51367;
  assign n51369 = ~i_nEMPTY & ~n51368;
  assign n51370 = ~n31529 & ~n51369;
  assign n51371 = ~controllable_BtoS_ACK0 & ~n51370;
  assign n51372 = ~n51361 & ~n51371;
  assign n51373 = n4465 & ~n51372;
  assign n51374 = ~n48509 & ~n51373;
  assign n51375 = i_StoB_REQ10 & ~n51374;
  assign n51376 = ~n51349 & ~n51375;
  assign n51377 = ~controllable_BtoS_ACK10 & ~n51376;
  assign n51378 = ~n51351 & ~n51377;
  assign n51379 = n4464 & ~n51378;
  assign n51380 = ~n48516 & ~n51379;
  assign n51381 = n4463 & ~n51380;
  assign n51382 = ~n31548 & ~n51381;
  assign n51383 = n4462 & ~n51382;
  assign n51384 = ~n50420 & ~n51383;
  assign n51385 = ~n4461 & ~n51384;
  assign n51386 = ~n51253 & ~n51385;
  assign n51387 = ~n4459 & ~n51386;
  assign n51388 = ~n31644 & ~n49930;
  assign n51389 = ~controllable_BtoR_REQ0 & ~n51388;
  assign n51390 = ~n49929 & ~n51389;
  assign n51391 = ~i_RtoB_ACK0 & ~n51390;
  assign n51392 = ~n20983 & ~n51391;
  assign n51393 = ~controllable_DEQ & ~n51392;
  assign n51394 = ~n20981 & ~n51393;
  assign n51395 = i_nEMPTY & ~n51394;
  assign n51396 = ~n31663 & ~n49943;
  assign n51397 = ~controllable_BtoR_REQ0 & ~n51396;
  assign n51398 = ~n49942 & ~n51397;
  assign n51399 = ~i_RtoB_ACK0 & ~n51398;
  assign n51400 = ~n20977 & ~n51399;
  assign n51401 = ~controllable_DEQ & ~n51400;
  assign n51402 = ~n20993 & ~n51401;
  assign n51403 = i_FULL & ~n51402;
  assign n51404 = ~n5242 & ~n49956;
  assign n51405 = ~controllable_BtoR_REQ0 & ~n51404;
  assign n51406 = ~n49955 & ~n51405;
  assign n51407 = ~i_RtoB_ACK0 & ~n51406;
  assign n51408 = ~n20977 & ~n51407;
  assign n51409 = ~controllable_DEQ & ~n51408;
  assign n51410 = ~n21003 & ~n51409;
  assign n51411 = ~i_FULL & ~n51410;
  assign n51412 = ~n51403 & ~n51411;
  assign n51413 = ~i_nEMPTY & ~n51412;
  assign n51414 = ~n51395 & ~n51413;
  assign n51415 = controllable_BtoS_ACK0 & ~n51414;
  assign n51416 = ~n31690 & ~n49973;
  assign n51417 = ~controllable_BtoR_REQ0 & ~n51416;
  assign n51418 = ~n49972 & ~n51417;
  assign n51419 = ~i_RtoB_ACK0 & ~n51418;
  assign n51420 = ~n29631 & ~n51419;
  assign n51421 = ~controllable_DEQ & ~n51420;
  assign n51422 = ~n29641 & ~n51421;
  assign n51423 = i_nEMPTY & ~n51422;
  assign n51424 = ~n31709 & ~n49986;
  assign n51425 = ~controllable_BtoR_REQ0 & ~n51424;
  assign n51426 = ~n49985 & ~n51425;
  assign n51427 = ~i_RtoB_ACK0 & ~n51426;
  assign n51428 = ~n29625 & ~n51427;
  assign n51429 = ~controllable_DEQ & ~n51428;
  assign n51430 = ~n29653 & ~n51429;
  assign n51431 = i_FULL & ~n51430;
  assign n51432 = ~n27878 & ~n49999;
  assign n51433 = ~controllable_BtoR_REQ0 & ~n51432;
  assign n51434 = ~n49998 & ~n51433;
  assign n51435 = ~i_RtoB_ACK0 & ~n51434;
  assign n51436 = ~n29625 & ~n51435;
  assign n51437 = ~controllable_DEQ & ~n51436;
  assign n51438 = ~n29663 & ~n51437;
  assign n51439 = ~i_FULL & ~n51438;
  assign n51440 = ~n51431 & ~n51439;
  assign n51441 = ~i_nEMPTY & ~n51440;
  assign n51442 = ~n51423 & ~n51441;
  assign n51443 = ~controllable_BtoS_ACK0 & ~n51442;
  assign n51444 = ~n51415 & ~n51443;
  assign n51445 = n4465 & ~n51444;
  assign n51446 = ~n48393 & ~n51445;
  assign n51447 = i_StoB_REQ10 & ~n51446;
  assign n51448 = ~n31786 & ~n50020;
  assign n51449 = ~controllable_BtoR_REQ0 & ~n51448;
  assign n51450 = ~n50019 & ~n51449;
  assign n51451 = ~i_RtoB_ACK0 & ~n51450;
  assign n51452 = ~n23095 & ~n51451;
  assign n51453 = ~controllable_DEQ & ~n51452;
  assign n51454 = ~n23093 & ~n51453;
  assign n51455 = i_nEMPTY & ~n51454;
  assign n51456 = ~n31805 & ~n50033;
  assign n51457 = ~controllable_BtoR_REQ0 & ~n51456;
  assign n51458 = ~n50032 & ~n51457;
  assign n51459 = ~i_RtoB_ACK0 & ~n51458;
  assign n51460 = ~n23107 & ~n51459;
  assign n51461 = ~controllable_DEQ & ~n51460;
  assign n51462 = ~n23105 & ~n51461;
  assign n51463 = i_FULL & ~n51462;
  assign n51464 = ~n11236 & ~n49663;
  assign n51465 = ~controllable_BtoR_REQ0 & ~n51464;
  assign n51466 = ~n50045 & ~n51465;
  assign n51467 = ~i_RtoB_ACK0 & ~n51466;
  assign n51468 = ~n23089 & ~n51467;
  assign n51469 = ~controllable_DEQ & ~n51468;
  assign n51470 = ~n23117 & ~n51469;
  assign n51471 = ~i_FULL & ~n51470;
  assign n51472 = ~n51463 & ~n51471;
  assign n51473 = ~i_nEMPTY & ~n51472;
  assign n51474 = ~n51455 & ~n51473;
  assign n51475 = controllable_BtoS_ACK0 & ~n51474;
  assign n51476 = ~n31832 & ~n50062;
  assign n51477 = ~controllable_BtoR_REQ0 & ~n51476;
  assign n51478 = ~n50061 & ~n51477;
  assign n51479 = ~i_RtoB_ACK0 & ~n51478;
  assign n51480 = ~n23135 & ~n51479;
  assign n51481 = ~controllable_DEQ & ~n51480;
  assign n51482 = ~n23133 & ~n51481;
  assign n51483 = i_nEMPTY & ~n51482;
  assign n51484 = ~n31851 & ~n50075;
  assign n51485 = ~controllable_BtoR_REQ0 & ~n51484;
  assign n51486 = ~n50074 & ~n51485;
  assign n51487 = ~i_RtoB_ACK0 & ~n51486;
  assign n51488 = ~n23147 & ~n51487;
  assign n51489 = ~controllable_DEQ & ~n51488;
  assign n51490 = ~n23145 & ~n51489;
  assign n51491 = i_FULL & ~n51490;
  assign n51492 = ~n11315 & ~n49708;
  assign n51493 = ~controllable_BtoR_REQ0 & ~n51492;
  assign n51494 = ~n50087 & ~n51493;
  assign n51495 = ~i_RtoB_ACK0 & ~n51494;
  assign n51496 = ~n23129 & ~n51495;
  assign n51497 = ~controllable_DEQ & ~n51496;
  assign n51498 = ~n23157 & ~n51497;
  assign n51499 = ~i_FULL & ~n51498;
  assign n51500 = ~n51491 & ~n51499;
  assign n51501 = ~i_nEMPTY & ~n51500;
  assign n51502 = ~n51483 & ~n51501;
  assign n51503 = ~controllable_BtoS_ACK0 & ~n51502;
  assign n51504 = ~n51475 & ~n51503;
  assign n51505 = n4465 & ~n51504;
  assign n51506 = ~n48454 & ~n51505;
  assign n51507 = ~i_StoB_REQ10 & ~n51506;
  assign n51508 = ~n51447 & ~n51507;
  assign n51509 = controllable_BtoS_ACK10 & ~n51508;
  assign n51510 = ~n28133 & ~n49733;
  assign n51511 = ~controllable_BtoR_REQ0 & ~n51510;
  assign n51512 = ~n50533 & ~n51511;
  assign n51513 = ~i_RtoB_ACK0 & ~n51512;
  assign n51514 = ~n29825 & ~n51513;
  assign n51515 = ~controllable_DEQ & ~n51514;
  assign n51516 = ~n29872 & ~n51515;
  assign n51517 = ~i_FULL & ~n51516;
  assign n51518 = ~n29951 & ~n51517;
  assign n51519 = ~i_nEMPTY & ~n51518;
  assign n51520 = ~n29944 & ~n51519;
  assign n51521 = controllable_BtoS_ACK0 & ~n51520;
  assign n51522 = ~n28194 & ~n49752;
  assign n51523 = ~controllable_BtoR_REQ0 & ~n51522;
  assign n51524 = ~n50556 & ~n51523;
  assign n51525 = ~i_RtoB_ACK0 & ~n51524;
  assign n51526 = ~n29881 & ~n51525;
  assign n51527 = ~controllable_DEQ & ~n51526;
  assign n51528 = ~n29928 & ~n51527;
  assign n51529 = ~i_FULL & ~n51528;
  assign n51530 = ~n31535 & ~n51529;
  assign n51531 = ~i_nEMPTY & ~n51530;
  assign n51532 = ~n31529 & ~n51531;
  assign n51533 = ~controllable_BtoS_ACK0 & ~n51532;
  assign n51534 = ~n51521 & ~n51533;
  assign n51535 = n4465 & ~n51534;
  assign n51536 = ~n48509 & ~n51535;
  assign n51537 = i_StoB_REQ10 & ~n51536;
  assign n51538 = ~n51507 & ~n51537;
  assign n51539 = ~controllable_BtoS_ACK10 & ~n51538;
  assign n51540 = ~n51509 & ~n51539;
  assign n51541 = n4464 & ~n51540;
  assign n51542 = ~n48516 & ~n51541;
  assign n51543 = ~n4463 & ~n51542;
  assign n51544 = ~n51121 & ~n51543;
  assign n51545 = n4462 & ~n51544;
  assign n51546 = ~n50420 & ~n51545;
  assign n51547 = n4461 & ~n51546;
  assign n51548 = ~n5255 & ~n50711;
  assign n51549 = ~controllable_BtoR_REQ0 & ~n51548;
  assign n51550 = ~n14765 & ~n51549;
  assign n51551 = ~i_RtoB_ACK0 & ~n51550;
  assign n51552 = ~n20983 & ~n51551;
  assign n51553 = ~controllable_DEQ & ~n51552;
  assign n51554 = ~n20981 & ~n51553;
  assign n51555 = i_nEMPTY & ~n51554;
  assign n51556 = ~n5232 & ~n50720;
  assign n51557 = ~controllable_BtoR_REQ0 & ~n51556;
  assign n51558 = ~n14784 & ~n51557;
  assign n51559 = ~i_RtoB_ACK0 & ~n51558;
  assign n51560 = ~n20977 & ~n51559;
  assign n51561 = ~controllable_DEQ & ~n51560;
  assign n51562 = ~n20993 & ~n51561;
  assign n51563 = i_FULL & ~n51562;
  assign n51564 = ~n14799 & ~n50729;
  assign n51565 = ~controllable_BtoR_REQ0 & ~n51564;
  assign n51566 = ~n14749 & ~n51565;
  assign n51567 = ~i_RtoB_ACK0 & ~n51566;
  assign n51568 = ~n20977 & ~n51567;
  assign n51569 = ~controllable_DEQ & ~n51568;
  assign n51570 = ~n21003 & ~n51569;
  assign n51571 = ~i_FULL & ~n51570;
  assign n51572 = ~n51563 & ~n51571;
  assign n51573 = ~i_nEMPTY & ~n51572;
  assign n51574 = ~n51555 & ~n51573;
  assign n51575 = controllable_BtoS_ACK0 & ~n51574;
  assign n51576 = ~n20328 & ~n50742;
  assign n51577 = ~controllable_BtoR_REQ0 & ~n51576;
  assign n51578 = ~n29437 & ~n51577;
  assign n51579 = ~i_RtoB_ACK0 & ~n51578;
  assign n51580 = ~n29631 & ~n51579;
  assign n51581 = ~controllable_DEQ & ~n51580;
  assign n51582 = ~n29641 & ~n51581;
  assign n51583 = i_nEMPTY & ~n51582;
  assign n51584 = ~n20337 & ~n50751;
  assign n51585 = ~controllable_BtoR_REQ0 & ~n51584;
  assign n51586 = ~n29447 & ~n51585;
  assign n51587 = ~i_RtoB_ACK0 & ~n51586;
  assign n51588 = ~n29625 & ~n51587;
  assign n51589 = ~controllable_DEQ & ~n51588;
  assign n51590 = ~n29653 & ~n51589;
  assign n51591 = i_FULL & ~n51590;
  assign n51592 = ~n20347 & ~n50760;
  assign n51593 = ~controllable_BtoR_REQ0 & ~n51592;
  assign n51594 = ~n28753 & ~n51593;
  assign n51595 = ~i_RtoB_ACK0 & ~n51594;
  assign n51596 = ~n29625 & ~n51595;
  assign n51597 = ~controllable_DEQ & ~n51596;
  assign n51598 = ~n29663 & ~n51597;
  assign n51599 = ~i_FULL & ~n51598;
  assign n51600 = ~n51591 & ~n51599;
  assign n51601 = ~i_nEMPTY & ~n51600;
  assign n51602 = ~n51583 & ~n51601;
  assign n51603 = ~controllable_BtoS_ACK0 & ~n51602;
  assign n51604 = ~n51575 & ~n51603;
  assign n51605 = n4465 & ~n51604;
  assign n51606 = ~n48393 & ~n51605;
  assign n51607 = i_StoB_REQ10 & ~n51606;
  assign n51608 = ~n11248 & ~n50777;
  assign n51609 = ~controllable_BtoR_REQ0 & ~n51608;
  assign n51610 = ~n17635 & ~n51609;
  assign n51611 = ~i_RtoB_ACK0 & ~n51610;
  assign n51612 = ~n23095 & ~n51611;
  assign n51613 = ~controllable_DEQ & ~n51612;
  assign n51614 = ~n23093 & ~n51613;
  assign n51615 = i_nEMPTY & ~n51614;
  assign n51616 = ~n11230 & ~n50786;
  assign n51617 = ~controllable_BtoR_REQ0 & ~n51616;
  assign n51618 = ~n17657 & ~n51617;
  assign n51619 = ~i_RtoB_ACK0 & ~n51618;
  assign n51620 = ~n23107 & ~n51619;
  assign n51621 = ~controllable_DEQ & ~n51620;
  assign n51622 = ~n23105 & ~n51621;
  assign n51623 = i_FULL & ~n51622;
  assign n51624 = ~n11284 & ~n49661;
  assign n51625 = ~controllable_BtoR_REQ0 & ~n51624;
  assign n51626 = ~n17620 & ~n51625;
  assign n51627 = ~i_RtoB_ACK0 & ~n51626;
  assign n51628 = ~n23089 & ~n51627;
  assign n51629 = ~controllable_DEQ & ~n51628;
  assign n51630 = ~n23117 & ~n51629;
  assign n51631 = ~i_FULL & ~n51630;
  assign n51632 = ~n51623 & ~n51631;
  assign n51633 = ~i_nEMPTY & ~n51632;
  assign n51634 = ~n51615 & ~n51633;
  assign n51635 = controllable_BtoS_ACK0 & ~n51634;
  assign n51636 = ~n11328 & ~n50807;
  assign n51637 = ~controllable_BtoR_REQ0 & ~n51636;
  assign n51638 = ~n17718 & ~n51637;
  assign n51639 = ~i_RtoB_ACK0 & ~n51638;
  assign n51640 = ~n23135 & ~n51639;
  assign n51641 = ~controllable_DEQ & ~n51640;
  assign n51642 = ~n23133 & ~n51641;
  assign n51643 = i_nEMPTY & ~n51642;
  assign n51644 = ~n11305 & ~n50816;
  assign n51645 = ~controllable_BtoR_REQ0 & ~n51644;
  assign n51646 = ~n17751 & ~n51645;
  assign n51647 = ~i_RtoB_ACK0 & ~n51646;
  assign n51648 = ~n23147 & ~n51647;
  assign n51649 = ~controllable_DEQ & ~n51648;
  assign n51650 = ~n23145 & ~n51649;
  assign n51651 = i_FULL & ~n51650;
  assign n51652 = ~n11366 & ~n49706;
  assign n51653 = ~controllable_BtoR_REQ0 & ~n51652;
  assign n51654 = ~n17699 & ~n51653;
  assign n51655 = ~i_RtoB_ACK0 & ~n51654;
  assign n51656 = ~n23129 & ~n51655;
  assign n51657 = ~controllable_DEQ & ~n51656;
  assign n51658 = ~n23157 & ~n51657;
  assign n51659 = ~i_FULL & ~n51658;
  assign n51660 = ~n51651 & ~n51659;
  assign n51661 = ~i_nEMPTY & ~n51660;
  assign n51662 = ~n51643 & ~n51661;
  assign n51663 = ~controllable_BtoS_ACK0 & ~n51662;
  assign n51664 = ~n51635 & ~n51663;
  assign n51665 = n4465 & ~n51664;
  assign n51666 = ~n48454 & ~n51665;
  assign n51667 = ~i_StoB_REQ10 & ~n51666;
  assign n51668 = ~n51607 & ~n51667;
  assign n51669 = controllable_BtoS_ACK10 & ~n51668;
  assign n51670 = ~n11238 & ~n49731;
  assign n51671 = ~controllable_BtoR_REQ0 & ~n51670;
  assign n51672 = ~n29840 & ~n51671;
  assign n51673 = ~i_RtoB_ACK0 & ~n51672;
  assign n51674 = ~n29825 & ~n51673;
  assign n51675 = ~controllable_DEQ & ~n51674;
  assign n51676 = ~n29872 & ~n51675;
  assign n51677 = ~i_FULL & ~n51676;
  assign n51678 = ~n29951 & ~n51677;
  assign n51679 = ~i_nEMPTY & ~n51678;
  assign n51680 = ~n29944 & ~n51679;
  assign n51681 = controllable_BtoS_ACK0 & ~n51680;
  assign n51682 = ~n11317 & ~n49750;
  assign n51683 = ~controllable_BtoR_REQ0 & ~n51682;
  assign n51684 = ~n29896 & ~n51683;
  assign n51685 = ~i_RtoB_ACK0 & ~n51684;
  assign n51686 = ~n29881 & ~n51685;
  assign n51687 = ~controllable_DEQ & ~n51686;
  assign n51688 = ~n29928 & ~n51687;
  assign n51689 = ~i_FULL & ~n51688;
  assign n51690 = ~n31535 & ~n51689;
  assign n51691 = ~i_nEMPTY & ~n51690;
  assign n51692 = ~n31529 & ~n51691;
  assign n51693 = ~controllable_BtoS_ACK0 & ~n51692;
  assign n51694 = ~n51681 & ~n51693;
  assign n51695 = n4465 & ~n51694;
  assign n51696 = ~n48509 & ~n51695;
  assign n51697 = i_StoB_REQ10 & ~n51696;
  assign n51698 = ~n51667 & ~n51697;
  assign n51699 = ~controllable_BtoS_ACK10 & ~n51698;
  assign n51700 = ~n51669 & ~n51699;
  assign n51701 = n4464 & ~n51700;
  assign n51702 = ~n48516 & ~n51701;
  assign n51703 = n4463 & ~n51702;
  assign n51704 = ~n31548 & ~n51703;
  assign n51705 = n4462 & ~n51704;
  assign n51706 = ~n50420 & ~n51705;
  assign n51707 = ~n4461 & ~n51706;
  assign n51708 = ~n51547 & ~n51707;
  assign n51709 = n4459 & ~n51708;
  assign n51710 = ~n51387 & ~n51709;
  assign n51711 = ~n4455 & ~n51710;
  assign n51712 = ~n51120 & ~n51711;
  assign n51713 = ~n4445 & ~n51712;
  assign n51714 = ~n51110 & ~n51713;
  assign n51715 = ~n4442 & ~n51714;
  assign n51716 = ~n49320 & ~n51715;
  assign n51717 = ~n4438 & ~n51716;
  assign n51718 = ~n4438 & ~n51717;
  assign n51719 = n4386 & ~n51718;
  assign n51720 = ~n4438 & ~n36619;
  assign n51721 = ~n4438 & ~n51720;
  assign n51722 = ~n4386 & ~n51721;
  assign n51723 = ~n51719 & ~n51722;
  assign n51724 = n4384 & n51723;
  assign n51725 = n4384 & ~n51724;
  assign n51726 = ~n4244 & ~n51725;
  assign n51727 = ~n36628 & ~n51726;
  assign inductivity_check  = ~n4150 & n51727;
endmodule


