// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module factorization16_simplified ( i2[15], i2[14], i2[13], i2[12], i2[11], i2[10], i2[9], i2[8], i1[15], i1[14], i1[13], i1[12], i1[11], i1[10], i1[9], i1[8], a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], o_1 );
input i2[15];
input i2[14];
input i2[13];
input i2[12];
input i2[11];
input i2[10];
input i2[9];
input i2[8];
input i1[15];
input i1[14];
input i1[13];
input i1[12];
input i1[11];
input i1[10];
input i1[9];
input i1[8];
input a[0];
input a[1];
input a[2];
input a[3];
input a[4];
input a[5];
input a[6];
input a[7];
input a[8];
input a[9];
input a[10];
input a[11];
input a[12];
input a[13];
input a[14];
input a[15];
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
assign n_1 =  i2[8] &  i1[8];
assign n_2 =  i2[8] &  i1[9];
assign n_3 =  i2[8] &  i1[10];
assign n_4 =  i2[8] &  i1[11];
assign n_5 =  i2[8] &  i1[12];
assign n_6 =  i2[8] &  i1[13];
assign n_7 =  i2[9] &  i1[14];
assign n_8 =  i2[8] &  i1[15];
assign n_9 =  n_7 &  n_8;
assign n_10 =  i2[10] &  i1[14];
assign n_11 =  i2[9] &  i1[15];
assign n_12 =  n_10 &  n_11;
assign n_13 =  i2[11] &  i1[14];
assign n_14 =  i2[10] &  i1[15];
assign n_15 =  n_13 &  n_14;
assign n_16 =  i2[12] &  i1[14];
assign n_17 =  i2[11] &  i1[15];
assign n_18 =  n_16 &  n_17;
assign n_19 =  i2[13] &  i1[14];
assign n_20 =  i2[12] &  i1[15];
assign n_21 =  n_19 &  n_20;
assign n_22 =  i2[14] &  i1[15];
assign n_23 =  i2[15] &  i1[14];
assign n_24 =  n_22 &  n_23;
assign n_25 =  i2[14] &  i1[14];
assign n_26 =  i2[13] &  i1[15];
assign n_27 =  n_25 &  n_26;
assign n_28 = ~n_24 & ~n_27;
assign n_29 = ~n_19 & ~n_20;
assign n_30 = ~n_29 & ~n_21;
assign n_31 = ~n_28 &  n_30;
assign n_32 = ~n_21 & ~n_31;
assign n_33 = ~n_16 & ~n_17;
assign n_34 = ~n_33 & ~n_18;
assign n_35 = ~n_32 &  n_34;
assign n_36 = ~n_18 & ~n_35;
assign n_37 = ~n_13 & ~n_14;
assign n_38 = ~n_37 & ~n_15;
assign n_39 = ~n_36 &  n_38;
assign n_40 = ~n_15 & ~n_39;
assign n_41 = ~n_10 & ~n_11;
assign n_42 = ~n_41 & ~n_12;
assign n_43 = ~n_40 &  n_42;
assign n_44 = ~n_12 & ~n_43;
assign n_45 = ~n_7 & ~n_8;
assign n_46 = ~n_45 & ~n_9;
assign n_47 = ~n_44 &  n_46;
assign n_48 = ~n_9 & ~n_47;
assign n_49 =  i2[8] &  i1[14];
assign n_50 = ~n_48 &  n_49;
assign n_51 =  n_6 &  n_50;
assign n_52 =  i2[9] &  i1[13];
assign n_53 =  n_48 & ~n_49;
assign n_54 = ~n_50 & ~n_53;
assign n_55 =  n_52 &  n_54;
assign n_56 =  n_44 & ~n_46;
assign n_57 = ~n_47 & ~n_56;
assign n_58 =  i2[10] &  i1[13];
assign n_59 =  n_57 &  n_58;
assign n_60 =  n_40 & ~n_42;
assign n_61 = ~n_43 & ~n_60;
assign n_62 =  i2[11] &  i1[13];
assign n_63 =  n_61 &  n_62;
assign n_64 =  n_36 & ~n_38;
assign n_65 = ~n_39 & ~n_64;
assign n_66 =  i2[12] &  i1[13];
assign n_67 =  n_65 &  n_66;
assign n_68 =  n_32 & ~n_34;
assign n_69 = ~n_35 & ~n_68;
assign n_70 =  i2[13] &  i1[13];
assign n_71 =  n_69 &  n_70;
assign n_72 =  n_28 & ~n_30;
assign n_73 = ~n_31 & ~n_72;
assign n_74 =  i2[14] &  i1[13];
assign n_75 =  n_73 &  n_74;
assign n_76 =  i2[15] &  i1[13];
assign n_77 =  n_24 &  n_27;
assign n_78 = ~n_28 & ~n_77;
assign n_79 = ~n_25 & ~n_26;
assign n_80 = ~n_78 & ~n_79;
assign n_81 =  n_76 &  n_80;
assign n_82 = ~n_73 & ~n_74;
assign n_83 = ~n_75 & ~n_82;
assign n_84 =  n_81 &  n_83;
assign n_85 = ~n_75 & ~n_84;
assign n_86 = ~n_69 & ~n_70;
assign n_87 = ~n_71 & ~n_86;
assign n_88 = ~n_85 &  n_87;
assign n_89 = ~n_71 & ~n_88;
assign n_90 = ~n_65 & ~n_66;
assign n_91 = ~n_67 & ~n_90;
assign n_92 = ~n_89 &  n_91;
assign n_93 = ~n_67 & ~n_92;
assign n_94 = ~n_61 & ~n_62;
assign n_95 = ~n_63 & ~n_94;
assign n_96 = ~n_93 &  n_95;
assign n_97 = ~n_63 & ~n_96;
assign n_98 = ~n_57 & ~n_58;
assign n_99 = ~n_59 & ~n_98;
assign n_100 = ~n_97 &  n_99;
assign n_101 = ~n_59 & ~n_100;
assign n_102 = ~n_52 & ~n_54;
assign n_103 = ~n_55 & ~n_102;
assign n_104 = ~n_101 &  n_103;
assign n_105 = ~n_55 & ~n_104;
assign n_106 = ~n_6 & ~n_50;
assign n_107 = ~n_51 & ~n_106;
assign n_108 = ~n_105 &  n_107;
assign n_109 = ~n_51 & ~n_108;
assign n_110 =  n_5 & ~n_109;
assign n_111 =  i2[9] &  i1[12];
assign n_112 =  n_105 & ~n_107;
assign n_113 = ~n_108 & ~n_112;
assign n_114 =  n_111 &  n_113;
assign n_115 =  i2[10] &  i1[12];
assign n_116 =  n_101 & ~n_103;
assign n_117 = ~n_104 & ~n_116;
assign n_118 =  n_115 &  n_117;
assign n_119 =  n_97 & ~n_99;
assign n_120 = ~n_100 & ~n_119;
assign n_121 =  i2[11] &  i1[12];
assign n_122 =  n_120 &  n_121;
assign n_123 =  n_93 & ~n_95;
assign n_124 = ~n_96 & ~n_123;
assign n_125 =  i2[12] &  i1[12];
assign n_126 =  n_124 &  n_125;
assign n_127 =  n_89 & ~n_91;
assign n_128 = ~n_92 & ~n_127;
assign n_129 =  i2[13] &  i1[12];
assign n_130 =  n_128 &  n_129;
assign n_131 =  n_85 & ~n_87;
assign n_132 = ~n_88 & ~n_131;
assign n_133 =  i2[14] &  i1[12];
assign n_134 =  n_132 &  n_133;
assign n_135 = ~n_81 & ~n_83;
assign n_136 = ~n_84 & ~n_135;
assign n_137 =  i2[15] &  i1[12];
assign n_138 =  n_136 &  n_137;
assign n_139 = ~n_132 & ~n_133;
assign n_140 = ~n_134 & ~n_139;
assign n_141 =  n_138 &  n_140;
assign n_142 = ~n_134 & ~n_141;
assign n_143 = ~n_128 & ~n_129;
assign n_144 = ~n_130 & ~n_143;
assign n_145 = ~n_142 &  n_144;
assign n_146 = ~n_130 & ~n_145;
assign n_147 = ~n_124 & ~n_125;
assign n_148 = ~n_126 & ~n_147;
assign n_149 = ~n_146 &  n_148;
assign n_150 = ~n_126 & ~n_149;
assign n_151 = ~n_120 & ~n_121;
assign n_152 = ~n_122 & ~n_151;
assign n_153 = ~n_150 &  n_152;
assign n_154 = ~n_122 & ~n_153;
assign n_155 = ~n_115 & ~n_117;
assign n_156 = ~n_118 & ~n_155;
assign n_157 = ~n_154 &  n_156;
assign n_158 = ~n_118 & ~n_157;
assign n_159 = ~n_111 & ~n_113;
assign n_160 = ~n_114 & ~n_159;
assign n_161 = ~n_158 &  n_160;
assign n_162 = ~n_114 & ~n_161;
assign n_163 = ~n_5 &  n_109;
assign n_164 = ~n_110 & ~n_163;
assign n_165 = ~n_162 &  n_164;
assign n_166 = ~n_110 & ~n_165;
assign n_167 =  n_4 & ~n_166;
assign n_168 =  i2[9] &  i1[11];
assign n_169 =  n_162 & ~n_164;
assign n_170 = ~n_165 & ~n_169;
assign n_171 =  n_168 &  n_170;
assign n_172 =  i2[10] &  i1[11];
assign n_173 =  n_158 & ~n_160;
assign n_174 = ~n_161 & ~n_173;
assign n_175 =  n_172 &  n_174;
assign n_176 =  i2[11] &  i1[11];
assign n_177 =  n_154 & ~n_156;
assign n_178 = ~n_157 & ~n_177;
assign n_179 =  n_176 &  n_178;
assign n_180 =  n_150 & ~n_152;
assign n_181 = ~n_153 & ~n_180;
assign n_182 =  i2[12] &  i1[11];
assign n_183 =  n_181 &  n_182;
assign n_184 =  n_146 & ~n_148;
assign n_185 = ~n_149 & ~n_184;
assign n_186 =  i2[13] &  i1[11];
assign n_187 =  n_185 &  n_186;
assign n_188 =  n_142 & ~n_144;
assign n_189 = ~n_145 & ~n_188;
assign n_190 =  i2[14] &  i1[11];
assign n_191 =  n_189 &  n_190;
assign n_192 = ~n_138 & ~n_140;
assign n_193 = ~n_141 & ~n_192;
assign n_194 =  i2[15] &  i1[11];
assign n_195 =  n_193 &  n_194;
assign n_196 = ~n_189 & ~n_190;
assign n_197 = ~n_191 & ~n_196;
assign n_198 =  n_195 &  n_197;
assign n_199 = ~n_191 & ~n_198;
assign n_200 = ~n_185 & ~n_186;
assign n_201 = ~n_187 & ~n_200;
assign n_202 = ~n_199 &  n_201;
assign n_203 = ~n_187 & ~n_202;
assign n_204 = ~n_181 & ~n_182;
assign n_205 = ~n_183 & ~n_204;
assign n_206 = ~n_203 &  n_205;
assign n_207 = ~n_183 & ~n_206;
assign n_208 = ~n_176 & ~n_178;
assign n_209 = ~n_179 & ~n_208;
assign n_210 = ~n_207 &  n_209;
assign n_211 = ~n_179 & ~n_210;
assign n_212 = ~n_172 & ~n_174;
assign n_213 = ~n_175 & ~n_212;
assign n_214 = ~n_211 &  n_213;
assign n_215 = ~n_175 & ~n_214;
assign n_216 = ~n_168 & ~n_170;
assign n_217 = ~n_171 & ~n_216;
assign n_218 = ~n_215 &  n_217;
assign n_219 = ~n_171 & ~n_218;
assign n_220 = ~n_4 &  n_166;
assign n_221 = ~n_167 & ~n_220;
assign n_222 = ~n_219 &  n_221;
assign n_223 = ~n_167 & ~n_222;
assign n_224 =  n_3 & ~n_223;
assign n_225 =  i2[9] &  i1[10];
assign n_226 =  n_219 & ~n_221;
assign n_227 = ~n_222 & ~n_226;
assign n_228 =  n_225 &  n_227;
assign n_229 =  i2[10] &  i1[10];
assign n_230 =  n_215 & ~n_217;
assign n_231 = ~n_218 & ~n_230;
assign n_232 =  n_229 &  n_231;
assign n_233 =  i2[11] &  i1[10];
assign n_234 =  n_211 & ~n_213;
assign n_235 = ~n_214 & ~n_234;
assign n_236 =  n_233 &  n_235;
assign n_237 =  i2[12] &  i1[10];
assign n_238 =  n_207 & ~n_209;
assign n_239 = ~n_210 & ~n_238;
assign n_240 =  n_237 &  n_239;
assign n_241 =  n_203 & ~n_205;
assign n_242 = ~n_206 & ~n_241;
assign n_243 =  i2[13] &  i1[10];
assign n_244 =  n_242 &  n_243;
assign n_245 =  n_199 & ~n_201;
assign n_246 = ~n_202 & ~n_245;
assign n_247 =  i2[14] &  i1[10];
assign n_248 =  n_246 &  n_247;
assign n_249 = ~n_195 & ~n_197;
assign n_250 = ~n_198 & ~n_249;
assign n_251 =  i2[15] &  i1[10];
assign n_252 =  n_250 &  n_251;
assign n_253 = ~n_246 & ~n_247;
assign n_254 = ~n_248 & ~n_253;
assign n_255 =  n_252 &  n_254;
assign n_256 = ~n_248 & ~n_255;
assign n_257 = ~n_242 & ~n_243;
assign n_258 = ~n_244 & ~n_257;
assign n_259 = ~n_256 &  n_258;
assign n_260 = ~n_244 & ~n_259;
assign n_261 = ~n_237 & ~n_239;
assign n_262 = ~n_240 & ~n_261;
assign n_263 = ~n_260 &  n_262;
assign n_264 = ~n_240 & ~n_263;
assign n_265 = ~n_233 & ~n_235;
assign n_266 = ~n_236 & ~n_265;
assign n_267 = ~n_264 &  n_266;
assign n_268 = ~n_236 & ~n_267;
assign n_269 = ~n_229 & ~n_231;
assign n_270 = ~n_232 & ~n_269;
assign n_271 = ~n_268 &  n_270;
assign n_272 = ~n_232 & ~n_271;
assign n_273 = ~n_225 & ~n_227;
assign n_274 = ~n_228 & ~n_273;
assign n_275 = ~n_272 &  n_274;
assign n_276 = ~n_228 & ~n_275;
assign n_277 = ~n_3 &  n_223;
assign n_278 = ~n_224 & ~n_277;
assign n_279 = ~n_276 &  n_278;
assign n_280 = ~n_224 & ~n_279;
assign n_281 =  n_2 & ~n_280;
assign n_282 =  i2[9] &  i1[9];
assign n_283 =  n_276 & ~n_278;
assign n_284 = ~n_279 & ~n_283;
assign n_285 =  n_282 &  n_284;
assign n_286 =  i2[10] &  i1[9];
assign n_287 =  n_272 & ~n_274;
assign n_288 = ~n_275 & ~n_287;
assign n_289 =  n_286 &  n_288;
assign n_290 =  i2[11] &  i1[9];
assign n_291 =  n_268 & ~n_270;
assign n_292 = ~n_271 & ~n_291;
assign n_293 =  n_290 &  n_292;
assign n_294 =  i2[12] &  i1[9];
assign n_295 =  n_264 & ~n_266;
assign n_296 = ~n_267 & ~n_295;
assign n_297 =  n_294 &  n_296;
assign n_298 =  i2[13] &  i1[9];
assign n_299 =  n_260 & ~n_262;
assign n_300 = ~n_263 & ~n_299;
assign n_301 =  n_298 &  n_300;
assign n_302 =  n_256 & ~n_258;
assign n_303 = ~n_259 & ~n_302;
assign n_304 =  i2[14] &  i1[9];
assign n_305 =  n_303 &  n_304;
assign n_306 = ~n_252 & ~n_254;
assign n_307 = ~n_255 & ~n_306;
assign n_308 =  i2[15] &  i1[9];
assign n_309 =  n_307 &  n_308;
assign n_310 = ~n_303 & ~n_304;
assign n_311 = ~n_305 & ~n_310;
assign n_312 =  n_309 &  n_311;
assign n_313 = ~n_305 & ~n_312;
assign n_314 = ~n_298 & ~n_300;
assign n_315 = ~n_301 & ~n_314;
assign n_316 = ~n_313 &  n_315;
assign n_317 = ~n_301 & ~n_316;
assign n_318 = ~n_294 & ~n_296;
assign n_319 = ~n_297 & ~n_318;
assign n_320 = ~n_317 &  n_319;
assign n_321 = ~n_297 & ~n_320;
assign n_322 = ~n_290 & ~n_292;
assign n_323 = ~n_293 & ~n_322;
assign n_324 = ~n_321 &  n_323;
assign n_325 = ~n_293 & ~n_324;
assign n_326 = ~n_286 & ~n_288;
assign n_327 = ~n_289 & ~n_326;
assign n_328 = ~n_325 &  n_327;
assign n_329 = ~n_289 & ~n_328;
assign n_330 = ~n_282 & ~n_284;
assign n_331 = ~n_285 & ~n_330;
assign n_332 = ~n_329 &  n_331;
assign n_333 = ~n_285 & ~n_332;
assign n_334 = ~n_2 &  n_280;
assign n_335 = ~n_281 & ~n_334;
assign n_336 = ~n_333 &  n_335;
assign n_337 = ~n_281 & ~n_336;
assign n_338 =  n_1 & ~n_337;
assign n_339 =  i2[9] &  i1[8];
assign n_340 =  n_333 & ~n_335;
assign n_341 = ~n_336 & ~n_340;
assign n_342 =  n_339 &  n_341;
assign n_343 =  i2[10] &  i1[8];
assign n_344 =  n_329 & ~n_331;
assign n_345 = ~n_332 & ~n_344;
assign n_346 =  n_343 &  n_345;
assign n_347 =  i2[11] &  i1[8];
assign n_348 =  n_325 & ~n_327;
assign n_349 = ~n_328 & ~n_348;
assign n_350 =  n_347 &  n_349;
assign n_351 =  i2[12] &  i1[8];
assign n_352 =  n_321 & ~n_323;
assign n_353 = ~n_324 & ~n_352;
assign n_354 =  n_351 &  n_353;
assign n_355 =  i2[13] &  i1[8];
assign n_356 =  n_317 & ~n_319;
assign n_357 = ~n_320 & ~n_356;
assign n_358 =  n_355 &  n_357;
assign n_359 =  i2[14] &  i1[8];
assign n_360 =  n_313 & ~n_315;
assign n_361 = ~n_316 & ~n_360;
assign n_362 =  n_359 &  n_361;
assign n_363 = ~n_309 & ~n_311;
assign n_364 = ~n_312 & ~n_363;
assign n_365 =  i2[15] &  i1[8];
assign n_366 =  n_364 &  n_365;
assign n_367 = ~n_359 & ~n_361;
assign n_368 = ~n_362 & ~n_367;
assign n_369 =  n_366 &  n_368;
assign n_370 = ~n_362 & ~n_369;
assign n_371 = ~n_355 & ~n_357;
assign n_372 = ~n_358 & ~n_371;
assign n_373 = ~n_370 &  n_372;
assign n_374 = ~n_358 & ~n_373;
assign n_375 = ~n_351 & ~n_353;
assign n_376 = ~n_354 & ~n_375;
assign n_377 = ~n_374 &  n_376;
assign n_378 = ~n_354 & ~n_377;
assign n_379 = ~n_347 & ~n_349;
assign n_380 = ~n_350 & ~n_379;
assign n_381 = ~n_378 &  n_380;
assign n_382 = ~n_350 & ~n_381;
assign n_383 = ~n_343 & ~n_345;
assign n_384 = ~n_346 & ~n_383;
assign n_385 = ~n_382 &  n_384;
assign n_386 = ~n_346 & ~n_385;
assign n_387 = ~n_339 & ~n_341;
assign n_388 = ~n_342 & ~n_387;
assign n_389 = ~n_386 &  n_388;
assign n_390 = ~n_342 & ~n_389;
assign n_391 = ~n_1 &  n_337;
assign n_392 = ~n_338 & ~n_391;
assign n_393 = ~n_390 &  n_392;
assign n_394 = ~n_338 & ~n_393;
assign n_395 =  a[0] &  n_394;
assign n_396 = ~a[0] & ~n_394;
assign n_397 =  n_390 & ~n_392;
assign n_398 = ~n_393 & ~n_397;
assign n_399 = ~a[1] &  n_398;
assign n_400 =  a[1] & ~n_398;
assign n_401 =  n_386 & ~n_388;
assign n_402 = ~n_389 & ~n_401;
assign n_403 = ~a[2] &  n_402;
assign n_404 =  a[2] & ~n_402;
assign n_405 =  n_382 & ~n_384;
assign n_406 = ~n_385 & ~n_405;
assign n_407 = ~a[3] &  n_406;
assign n_408 =  a[3] & ~n_406;
assign n_409 =  n_378 & ~n_380;
assign n_410 = ~n_381 & ~n_409;
assign n_411 = ~a[4] &  n_410;
assign n_412 =  a[4] & ~n_410;
assign n_413 =  n_374 & ~n_376;
assign n_414 = ~n_377 & ~n_413;
assign n_415 = ~a[5] &  n_414;
assign n_416 =  a[5] & ~n_414;
assign n_417 =  n_370 & ~n_372;
assign n_418 = ~n_373 & ~n_417;
assign n_419 = ~a[6] &  n_418;
assign n_420 =  a[6] & ~n_418;
assign n_421 = ~n_366 & ~n_368;
assign n_422 = ~n_369 & ~n_421;
assign n_423 = ~a[7] &  n_422;
assign n_424 =  a[7] & ~n_422;
assign n_425 = ~n_364 & ~n_365;
assign n_426 = ~n_366 & ~n_425;
assign n_427 = ~a[8] &  n_426;
assign n_428 =  a[8] & ~n_426;
assign n_429 = ~n_307 & ~n_308;
assign n_430 = ~n_309 & ~n_429;
assign n_431 = ~a[9] &  n_430;
assign n_432 =  a[9] & ~n_430;
assign n_433 = ~n_250 & ~n_251;
assign n_434 = ~n_252 & ~n_433;
assign n_435 = ~a[10] &  n_434;
assign n_436 =  a[10] & ~n_434;
assign n_437 = ~n_193 & ~n_194;
assign n_438 = ~n_195 & ~n_437;
assign n_439 = ~a[11] &  n_438;
assign n_440 =  a[11] & ~n_438;
assign n_441 = ~n_136 & ~n_137;
assign n_442 = ~n_138 & ~n_441;
assign n_443 = ~a[12] &  n_442;
assign n_444 =  a[12] & ~n_442;
assign n_445 = ~n_76 & ~n_80;
assign n_446 = ~n_81 & ~n_445;
assign n_447 = ~a[13] &  n_446;
assign n_448 =  a[13] & ~n_446;
assign n_449 =  i2[15] &  i1[15];
assign n_450 = ~a[15] & ~n_449;
assign n_451 =  a[15] &  n_449;
assign n_452 = ~n_450 & ~n_451;
assign n_453 = ~n_22 & ~n_23;
assign n_454 = ~n_24 & ~n_453;
assign n_455 =  a[14] & ~n_454;
assign n_456 = ~n_452 & ~n_455;
assign n_457 = ~i2[11] & ~i2[10];
assign n_458 = ~i2[9] & ~i2[8];
assign n_459 =  n_457 &  n_458;
assign n_460 =  i2[15] & ~i2[14];
assign n_461 = ~i2[13] & ~i2[12];
assign n_462 =  n_460 &  n_461;
assign n_463 =  n_459 &  n_462;
assign n_464 = ~i1[11] & ~i1[10];
assign n_465 = ~i1[9] & ~i1[8];
assign n_466 =  n_464 &  n_465;
assign n_467 =  i1[15] & ~i1[14];
assign n_468 = ~i1[13] & ~i1[12];
assign n_469 =  n_467 &  n_468;
assign n_470 =  n_466 &  n_469;
assign n_471 = ~a[14] &  n_454;
assign n_472 = ~n_470 & ~n_471;
assign n_473 = ~n_463 &  n_472;
assign n_474 =  n_456 &  n_473;
assign n_475 = ~n_448 &  n_474;
assign n_476 = ~n_447 &  n_475;
assign n_477 = ~n_444 &  n_476;
assign n_478 = ~n_443 &  n_477;
assign n_479 = ~n_440 &  n_478;
assign n_480 = ~n_439 &  n_479;
assign n_481 = ~n_436 &  n_480;
assign n_482 = ~n_435 &  n_481;
assign n_483 = ~n_432 &  n_482;
assign n_484 = ~n_431 &  n_483;
assign n_485 = ~n_428 &  n_484;
assign n_486 = ~n_427 &  n_485;
assign n_487 = ~n_424 &  n_486;
assign n_488 = ~n_423 &  n_487;
assign n_489 = ~n_420 &  n_488;
assign n_490 = ~n_419 &  n_489;
assign n_491 = ~n_416 &  n_490;
assign n_492 = ~n_415 &  n_491;
assign n_493 = ~n_412 &  n_492;
assign n_494 = ~n_411 &  n_493;
assign n_495 = ~n_408 &  n_494;
assign n_496 = ~n_407 &  n_495;
assign n_497 = ~n_404 &  n_496;
assign n_498 = ~n_403 &  n_497;
assign n_499 = ~n_400 &  n_498;
assign n_500 = ~n_399 &  n_499;
assign n_501 = ~n_396 &  n_500;
assign n_502 = ~n_395 &  n_501;
assign o_1 =  n_502;
endmodule

