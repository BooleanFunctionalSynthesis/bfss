// Generated using findDep.cpp 
module mult_bool_matrix_17_17_17.sat (v_20, v_15, v_63, v_68, v_73, v_78, v_83, v_88, v_25, v_58, v_53, v_48, v_43, v_38, v_33, v_28, v_9, v_18, v_13, v_65, v_70, v_75, v_80, v_85, v_90, v_23, v_60, v_55, v_50, v_45, v_40, v_35, v_30, v_6, v_291, v_287, v_328, v_332, v_336, v_340, v_344, v_348, v_295, v_324, v_320, v_316, v_312, v_308, v_304, v_300, v_283, v_551, v_547, v_588, v_592, v_596, v_600, v_604, v_608, v_555, v_584, v_580, v_576, v_572, v_568, v_564, v_560, v_543, v_811, v_807, v_848, v_852, v_856, v_860, v_864, v_868, v_815, v_844, v_840, v_836, v_832, v_828, v_824, v_820, v_803, v_1071, v_1067, v_1108, v_1112, v_1116, v_1120, v_1124, v_1128, v_1075, v_1104, v_1100, v_1096, v_1092, v_1088, v_1084, v_1080, v_1063, v_1331, v_1327, v_1368, v_1372, v_1376, v_1380, v_1384, v_1388, v_1335, v_1364, v_1360, v_1356, v_1352, v_1348, v_1344, v_1340, v_1323, v_1591, v_1587, v_1628, v_1632, v_1636, v_1640, v_1644, v_1648, v_1595, v_1624, v_1620, v_1616, v_1612, v_1608, v_1604, v_1600, v_1583, v_1851, v_1847, v_1888, v_1892, v_1896, v_1900, v_1904, v_1908, v_1855, v_1884, v_1880, v_1876, v_1872, v_1868, v_1864, v_1860, v_1843, v_2111, v_2107, v_2148, v_2152, v_2156, v_2160, v_2164, v_2168, v_2115, v_2144, v_2140, v_2136, v_2132, v_2128, v_2124, v_2120, v_2103, v_2371, v_2367, v_2408, v_2412, v_2416, v_2420, v_2424, v_2428, v_2375, v_2404, v_2400, v_2396, v_2392, v_2388, v_2384, v_2380, v_2363, v_2631, v_2627, v_2668, v_2672, v_2676, v_2680, v_2684, v_2688, v_2635, v_2664, v_2660, v_2656, v_2652, v_2648, v_2644, v_2640, v_2623, v_2891, v_2887, v_2928, v_2932, v_2936, v_2940, v_2944, v_2948, v_2895, v_2924, v_2920, v_2916, v_2912, v_2908, v_2904, v_2900, v_2883, v_3151, v_3147, v_3188, v_3192, v_3196, v_3200, v_3204, v_3208, v_3155, v_3184, v_3180, v_3176, v_3172, v_3168, v_3164, v_3160, v_3143, v_3411, v_3407, v_3448, v_3452, v_3456, v_3460, v_3464, v_3468, v_3415, v_3444, v_3440, v_3436, v_3432, v_3428, v_3424, v_3420, v_3403, v_3671, v_3667, v_3708, v_3712, v_3716, v_3720, v_3724, v_3728, v_3675, v_3704, v_3700, v_3696, v_3692, v_3688, v_3684, v_3680, v_3663, v_3931, v_3927, v_3968, v_3972, v_3976, v_3980, v_3984, v_3988, v_3935, v_3964, v_3960, v_3956, v_3952, v_3948, v_3944, v_3940, v_3923, v_4190, v_4186, v_4227, v_4231, v_4235, v_4239, v_4243, v_4247, v_4194, v_4223, v_4219, v_4215, v_4211, v_4207, v_4203, v_4199, v_4182, v_4452, v_4448, v_4487, v_4491, v_4495, v_4499, v_4503, v_4507, v_4456, v_4483, v_4479, v_4475, v_4471, v_4467, v_4463, v_4459, v_4444, v_8600, v_8596, v_8635, v_8639, v_8643, v_8647, v_8651, v_8655, v_8604, v_8631, v_8627, v_8623, v_8619, v_8615, v_8611, v_8607, v_8592, v_12748, v_12744, v_12783, v_12787, v_12791, v_12795, v_12799, v_12803, v_12752, v_12779, v_12775, v_12771, v_12767, v_12763, v_12759, v_12755, v_12740, v_16896, v_16892, v_16931, v_16935, v_16939, v_16943, v_16947, v_16951, v_16900, v_16927, v_16923, v_16919, v_16915, v_16911, v_16907, v_16903, v_16888, v_21044, v_21040, v_21079, v_21083, v_21087, v_21091, v_21095, v_21099, v_21048, v_21075, v_21071, v_21067, v_21063, v_21059, v_21055, v_21051, v_21036, v_25192, v_25188, v_25227, v_25231, v_25235, v_25239, v_25243, v_25247, v_25196, v_25223, v_25219, v_25215, v_25211, v_25207, v_25203, v_25199, v_25184, v_29340, v_29336, v_29375, v_29379, v_29383, v_29387, v_29391, v_29395, v_29344, v_29371, v_29367, v_29363, v_29359, v_29355, v_29351, v_29347, v_29332, v_33488, v_33484, v_33523, v_33527, v_33531, v_33535, v_33539, v_33543, v_33492, v_33519, v_33515, v_33511, v_33507, v_33503, v_33499, v_33495, v_33480, v_37636, v_37632, v_37671, v_37675, v_37679, v_37683, v_37687, v_37691, v_37640, v_37667, v_37663, v_37659, v_37655, v_37651, v_37647, v_37643, v_37628, v_41784, v_41780, v_41819, v_41823, v_41827, v_41831, v_41835, v_41839, v_41788, v_41815, v_41811, v_41807, v_41803, v_41799, v_41795, v_41791, v_41776, v_45932, v_45928, v_45967, v_45971, v_45975, v_45979, v_45983, v_45987, v_45936, v_45963, v_45959, v_45955, v_45951, v_45947, v_45943, v_45939, v_45924, v_50080, v_50076, v_50115, v_50119, v_50123, v_50127, v_50131, v_50135, v_50084, v_50111, v_50107, v_50103, v_50099, v_50095, v_50091, v_50087, v_50072, v_54228, v_54224, v_54263, v_54267, v_54271, v_54275, v_54279, v_54283, v_54232, v_54259, v_54255, v_54251, v_54247, v_54243, v_54239, v_54235, v_54220, v_58376, v_58372, v_58411, v_58415, v_58419, v_58423, v_58427, v_58431, v_58380, v_58407, v_58403, v_58399, v_58395, v_58391, v_58387, v_58383, v_58368, v_62524, v_62520, v_62559, v_62563, v_62567, v_62571, v_62575, v_62579, v_62528, v_62555, v_62551, v_62547, v_62543, v_62539, v_62535, v_62531, v_62516, v_66671, v_66667, v_66706, v_66710, v_66714, v_66718, v_66722, v_66726, v_66675, v_66702, v_66698, v_66694, v_66690, v_66686, v_66682, v_66678, v_66663, v_1, v_5, v_282, v_542, v_802, v_1062, v_1322, v_1582, v_1842, v_2102, v_2362, v_2622, v_2882, v_3142, v_3402, v_3662, v_3922, v_4348, v_4442, v_4702, v_4945, v_5188, v_5431, v_5674, v_5917, v_6160, v_6403, v_6646, v_6889, v_7132, v_7375, v_7618, v_7861, v_8104, v_8496, v_8590, v_8850, v_9093, v_9336, v_9579, v_9822, v_10065, v_10308, v_10551, v_10794, v_11037, v_11280, v_11523, v_11766, v_12009, v_12252, v_12644, v_12738, v_12998, v_13241, v_13484, v_13727, v_13970, v_14213, v_14456, v_14699, v_14942, v_15185, v_15428, v_15671, v_15914, v_16157, v_16400, v_16792, v_16886, v_17146, v_17389, v_17632, v_17875, v_18118, v_18361, v_18604, v_18847, v_19090, v_19333, v_19576, v_19819, v_20062, v_20305, v_20548, v_20940, v_21034, v_21294, v_21537, v_21780, v_22023, v_22266, v_22509, v_22752, v_22995, v_23238, v_23481, v_23724, v_23967, v_24210, v_24453, v_24696, v_25088, v_25182, v_25442, v_25685, v_25928, v_26171, v_26414, v_26657, v_26900, v_27143, v_27386, v_27629, v_27872, v_28115, v_28358, v_28601, v_28844, v_29236, v_29330, v_29590, v_29833, v_30076, v_30319, v_30562, v_30805, v_31048, v_31291, v_31534, v_31777, v_32020, v_32263, v_32506, v_32749, v_32992, v_33384, v_33478, v_33738, v_33981, v_34224, v_34467, v_34710, v_34953, v_35196, v_35439, v_35682, v_35925, v_36168, v_36411, v_36654, v_36897, v_37140, v_37532, v_37626, v_37886, v_38129, v_38372, v_38615, v_38858, v_39101, v_39344, v_39587, v_39830, v_40073, v_40316, v_40559, v_40802, v_41045, v_41288, v_41680, v_41774, v_42034, v_42277, v_42520, v_42763, v_43006, v_43249, v_43492, v_43735, v_43978, v_44221, v_44464, v_44707, v_44950, v_45193, v_45436, v_45828, v_45922, v_46182, v_46425, v_46668, v_46911, v_47154, v_47397, v_47640, v_47883, v_48126, v_48369, v_48612, v_48855, v_49098, v_49341, v_49584, v_49976, v_50070, v_50330, v_50573, v_50816, v_51059, v_51302, v_51545, v_51788, v_52031, v_52274, v_52517, v_52760, v_53003, v_53246, v_53489, v_53732, v_54124, v_54218, v_54478, v_54721, v_54964, v_55207, v_55450, v_55693, v_55936, v_56179, v_56422, v_56665, v_56908, v_57151, v_57394, v_57637, v_57880, v_58272, v_58366, v_58626, v_58869, v_59112, v_59355, v_59598, v_59841, v_60084, v_60327, v_60570, v_60813, v_61056, v_61299, v_61542, v_61785, v_62028, v_62420, v_62514, v_62774, v_63017, v_63260, v_63503, v_63746, v_63989, v_64232, v_64475, v_64718, v_64961, v_65204, v_65447, v_65690, v_65933, v_66176, v_66568, v_66828, v_67071, v_67314, v_67557, v_67800, v_68043, v_68286, v_68529, v_68772, v_69015, v_69258, v_69501, v_69744, v_69987, v_70230, v_70473, v_70716, v_4, o_1);
input v_20;
input v_15;
input v_63;
input v_68;
input v_73;
input v_78;
input v_83;
input v_88;
input v_25;
input v_58;
input v_53;
input v_48;
input v_43;
input v_38;
input v_33;
input v_28;
input v_9;
input v_18;
input v_13;
input v_65;
input v_70;
input v_75;
input v_80;
input v_85;
input v_90;
input v_23;
input v_60;
input v_55;
input v_50;
input v_45;
input v_40;
input v_35;
input v_30;
input v_6;
input v_291;
input v_287;
input v_328;
input v_332;
input v_336;
input v_340;
input v_344;
input v_348;
input v_295;
input v_324;
input v_320;
input v_316;
input v_312;
input v_308;
input v_304;
input v_300;
input v_283;
input v_551;
input v_547;
input v_588;
input v_592;
input v_596;
input v_600;
input v_604;
input v_608;
input v_555;
input v_584;
input v_580;
input v_576;
input v_572;
input v_568;
input v_564;
input v_560;
input v_543;
input v_811;
input v_807;
input v_848;
input v_852;
input v_856;
input v_860;
input v_864;
input v_868;
input v_815;
input v_844;
input v_840;
input v_836;
input v_832;
input v_828;
input v_824;
input v_820;
input v_803;
input v_1071;
input v_1067;
input v_1108;
input v_1112;
input v_1116;
input v_1120;
input v_1124;
input v_1128;
input v_1075;
input v_1104;
input v_1100;
input v_1096;
input v_1092;
input v_1088;
input v_1084;
input v_1080;
input v_1063;
input v_1331;
input v_1327;
input v_1368;
input v_1372;
input v_1376;
input v_1380;
input v_1384;
input v_1388;
input v_1335;
input v_1364;
input v_1360;
input v_1356;
input v_1352;
input v_1348;
input v_1344;
input v_1340;
input v_1323;
input v_1591;
input v_1587;
input v_1628;
input v_1632;
input v_1636;
input v_1640;
input v_1644;
input v_1648;
input v_1595;
input v_1624;
input v_1620;
input v_1616;
input v_1612;
input v_1608;
input v_1604;
input v_1600;
input v_1583;
input v_1851;
input v_1847;
input v_1888;
input v_1892;
input v_1896;
input v_1900;
input v_1904;
input v_1908;
input v_1855;
input v_1884;
input v_1880;
input v_1876;
input v_1872;
input v_1868;
input v_1864;
input v_1860;
input v_1843;
input v_2111;
input v_2107;
input v_2148;
input v_2152;
input v_2156;
input v_2160;
input v_2164;
input v_2168;
input v_2115;
input v_2144;
input v_2140;
input v_2136;
input v_2132;
input v_2128;
input v_2124;
input v_2120;
input v_2103;
input v_2371;
input v_2367;
input v_2408;
input v_2412;
input v_2416;
input v_2420;
input v_2424;
input v_2428;
input v_2375;
input v_2404;
input v_2400;
input v_2396;
input v_2392;
input v_2388;
input v_2384;
input v_2380;
input v_2363;
input v_2631;
input v_2627;
input v_2668;
input v_2672;
input v_2676;
input v_2680;
input v_2684;
input v_2688;
input v_2635;
input v_2664;
input v_2660;
input v_2656;
input v_2652;
input v_2648;
input v_2644;
input v_2640;
input v_2623;
input v_2891;
input v_2887;
input v_2928;
input v_2932;
input v_2936;
input v_2940;
input v_2944;
input v_2948;
input v_2895;
input v_2924;
input v_2920;
input v_2916;
input v_2912;
input v_2908;
input v_2904;
input v_2900;
input v_2883;
input v_3151;
input v_3147;
input v_3188;
input v_3192;
input v_3196;
input v_3200;
input v_3204;
input v_3208;
input v_3155;
input v_3184;
input v_3180;
input v_3176;
input v_3172;
input v_3168;
input v_3164;
input v_3160;
input v_3143;
input v_3411;
input v_3407;
input v_3448;
input v_3452;
input v_3456;
input v_3460;
input v_3464;
input v_3468;
input v_3415;
input v_3444;
input v_3440;
input v_3436;
input v_3432;
input v_3428;
input v_3424;
input v_3420;
input v_3403;
input v_3671;
input v_3667;
input v_3708;
input v_3712;
input v_3716;
input v_3720;
input v_3724;
input v_3728;
input v_3675;
input v_3704;
input v_3700;
input v_3696;
input v_3692;
input v_3688;
input v_3684;
input v_3680;
input v_3663;
input v_3931;
input v_3927;
input v_3968;
input v_3972;
input v_3976;
input v_3980;
input v_3984;
input v_3988;
input v_3935;
input v_3964;
input v_3960;
input v_3956;
input v_3952;
input v_3948;
input v_3944;
input v_3940;
input v_3923;
input v_4190;
input v_4186;
input v_4227;
input v_4231;
input v_4235;
input v_4239;
input v_4243;
input v_4247;
input v_4194;
input v_4223;
input v_4219;
input v_4215;
input v_4211;
input v_4207;
input v_4203;
input v_4199;
input v_4182;
input v_4452;
input v_4448;
input v_4487;
input v_4491;
input v_4495;
input v_4499;
input v_4503;
input v_4507;
input v_4456;
input v_4483;
input v_4479;
input v_4475;
input v_4471;
input v_4467;
input v_4463;
input v_4459;
input v_4444;
input v_8600;
input v_8596;
input v_8635;
input v_8639;
input v_8643;
input v_8647;
input v_8651;
input v_8655;
input v_8604;
input v_8631;
input v_8627;
input v_8623;
input v_8619;
input v_8615;
input v_8611;
input v_8607;
input v_8592;
input v_12748;
input v_12744;
input v_12783;
input v_12787;
input v_12791;
input v_12795;
input v_12799;
input v_12803;
input v_12752;
input v_12779;
input v_12775;
input v_12771;
input v_12767;
input v_12763;
input v_12759;
input v_12755;
input v_12740;
input v_16896;
input v_16892;
input v_16931;
input v_16935;
input v_16939;
input v_16943;
input v_16947;
input v_16951;
input v_16900;
input v_16927;
input v_16923;
input v_16919;
input v_16915;
input v_16911;
input v_16907;
input v_16903;
input v_16888;
input v_21044;
input v_21040;
input v_21079;
input v_21083;
input v_21087;
input v_21091;
input v_21095;
input v_21099;
input v_21048;
input v_21075;
input v_21071;
input v_21067;
input v_21063;
input v_21059;
input v_21055;
input v_21051;
input v_21036;
input v_25192;
input v_25188;
input v_25227;
input v_25231;
input v_25235;
input v_25239;
input v_25243;
input v_25247;
input v_25196;
input v_25223;
input v_25219;
input v_25215;
input v_25211;
input v_25207;
input v_25203;
input v_25199;
input v_25184;
input v_29340;
input v_29336;
input v_29375;
input v_29379;
input v_29383;
input v_29387;
input v_29391;
input v_29395;
input v_29344;
input v_29371;
input v_29367;
input v_29363;
input v_29359;
input v_29355;
input v_29351;
input v_29347;
input v_29332;
input v_33488;
input v_33484;
input v_33523;
input v_33527;
input v_33531;
input v_33535;
input v_33539;
input v_33543;
input v_33492;
input v_33519;
input v_33515;
input v_33511;
input v_33507;
input v_33503;
input v_33499;
input v_33495;
input v_33480;
input v_37636;
input v_37632;
input v_37671;
input v_37675;
input v_37679;
input v_37683;
input v_37687;
input v_37691;
input v_37640;
input v_37667;
input v_37663;
input v_37659;
input v_37655;
input v_37651;
input v_37647;
input v_37643;
input v_37628;
input v_41784;
input v_41780;
input v_41819;
input v_41823;
input v_41827;
input v_41831;
input v_41835;
input v_41839;
input v_41788;
input v_41815;
input v_41811;
input v_41807;
input v_41803;
input v_41799;
input v_41795;
input v_41791;
input v_41776;
input v_45932;
input v_45928;
input v_45967;
input v_45971;
input v_45975;
input v_45979;
input v_45983;
input v_45987;
input v_45936;
input v_45963;
input v_45959;
input v_45955;
input v_45951;
input v_45947;
input v_45943;
input v_45939;
input v_45924;
input v_50080;
input v_50076;
input v_50115;
input v_50119;
input v_50123;
input v_50127;
input v_50131;
input v_50135;
input v_50084;
input v_50111;
input v_50107;
input v_50103;
input v_50099;
input v_50095;
input v_50091;
input v_50087;
input v_50072;
input v_54228;
input v_54224;
input v_54263;
input v_54267;
input v_54271;
input v_54275;
input v_54279;
input v_54283;
input v_54232;
input v_54259;
input v_54255;
input v_54251;
input v_54247;
input v_54243;
input v_54239;
input v_54235;
input v_54220;
input v_58376;
input v_58372;
input v_58411;
input v_58415;
input v_58419;
input v_58423;
input v_58427;
input v_58431;
input v_58380;
input v_58407;
input v_58403;
input v_58399;
input v_58395;
input v_58391;
input v_58387;
input v_58383;
input v_58368;
input v_62524;
input v_62520;
input v_62559;
input v_62563;
input v_62567;
input v_62571;
input v_62575;
input v_62579;
input v_62528;
input v_62555;
input v_62551;
input v_62547;
input v_62543;
input v_62539;
input v_62535;
input v_62531;
input v_62516;
input v_66671;
input v_66667;
input v_66706;
input v_66710;
input v_66714;
input v_66718;
input v_66722;
input v_66726;
input v_66675;
input v_66702;
input v_66698;
input v_66694;
input v_66690;
input v_66686;
input v_66682;
input v_66678;
input v_66663;
input v_1;
input v_5;
input v_282;
input v_542;
input v_802;
input v_1062;
input v_1322;
input v_1582;
input v_1842;
input v_2102;
input v_2362;
input v_2622;
input v_2882;
input v_3142;
input v_3402;
input v_3662;
input v_3922;
input v_4348;
input v_4442;
input v_4702;
input v_4945;
input v_5188;
input v_5431;
input v_5674;
input v_5917;
input v_6160;
input v_6403;
input v_6646;
input v_6889;
input v_7132;
input v_7375;
input v_7618;
input v_7861;
input v_8104;
input v_8496;
input v_8590;
input v_8850;
input v_9093;
input v_9336;
input v_9579;
input v_9822;
input v_10065;
input v_10308;
input v_10551;
input v_10794;
input v_11037;
input v_11280;
input v_11523;
input v_11766;
input v_12009;
input v_12252;
input v_12644;
input v_12738;
input v_12998;
input v_13241;
input v_13484;
input v_13727;
input v_13970;
input v_14213;
input v_14456;
input v_14699;
input v_14942;
input v_15185;
input v_15428;
input v_15671;
input v_15914;
input v_16157;
input v_16400;
input v_16792;
input v_16886;
input v_17146;
input v_17389;
input v_17632;
input v_17875;
input v_18118;
input v_18361;
input v_18604;
input v_18847;
input v_19090;
input v_19333;
input v_19576;
input v_19819;
input v_20062;
input v_20305;
input v_20548;
input v_20940;
input v_21034;
input v_21294;
input v_21537;
input v_21780;
input v_22023;
input v_22266;
input v_22509;
input v_22752;
input v_22995;
input v_23238;
input v_23481;
input v_23724;
input v_23967;
input v_24210;
input v_24453;
input v_24696;
input v_25088;
input v_25182;
input v_25442;
input v_25685;
input v_25928;
input v_26171;
input v_26414;
input v_26657;
input v_26900;
input v_27143;
input v_27386;
input v_27629;
input v_27872;
input v_28115;
input v_28358;
input v_28601;
input v_28844;
input v_29236;
input v_29330;
input v_29590;
input v_29833;
input v_30076;
input v_30319;
input v_30562;
input v_30805;
input v_31048;
input v_31291;
input v_31534;
input v_31777;
input v_32020;
input v_32263;
input v_32506;
input v_32749;
input v_32992;
input v_33384;
input v_33478;
input v_33738;
input v_33981;
input v_34224;
input v_34467;
input v_34710;
input v_34953;
input v_35196;
input v_35439;
input v_35682;
input v_35925;
input v_36168;
input v_36411;
input v_36654;
input v_36897;
input v_37140;
input v_37532;
input v_37626;
input v_37886;
input v_38129;
input v_38372;
input v_38615;
input v_38858;
input v_39101;
input v_39344;
input v_39587;
input v_39830;
input v_40073;
input v_40316;
input v_40559;
input v_40802;
input v_41045;
input v_41288;
input v_41680;
input v_41774;
input v_42034;
input v_42277;
input v_42520;
input v_42763;
input v_43006;
input v_43249;
input v_43492;
input v_43735;
input v_43978;
input v_44221;
input v_44464;
input v_44707;
input v_44950;
input v_45193;
input v_45436;
input v_45828;
input v_45922;
input v_46182;
input v_46425;
input v_46668;
input v_46911;
input v_47154;
input v_47397;
input v_47640;
input v_47883;
input v_48126;
input v_48369;
input v_48612;
input v_48855;
input v_49098;
input v_49341;
input v_49584;
input v_49976;
input v_50070;
input v_50330;
input v_50573;
input v_50816;
input v_51059;
input v_51302;
input v_51545;
input v_51788;
input v_52031;
input v_52274;
input v_52517;
input v_52760;
input v_53003;
input v_53246;
input v_53489;
input v_53732;
input v_54124;
input v_54218;
input v_54478;
input v_54721;
input v_54964;
input v_55207;
input v_55450;
input v_55693;
input v_55936;
input v_56179;
input v_56422;
input v_56665;
input v_56908;
input v_57151;
input v_57394;
input v_57637;
input v_57880;
input v_58272;
input v_58366;
input v_58626;
input v_58869;
input v_59112;
input v_59355;
input v_59598;
input v_59841;
input v_60084;
input v_60327;
input v_60570;
input v_60813;
input v_61056;
input v_61299;
input v_61542;
input v_61785;
input v_62028;
input v_62420;
input v_62514;
input v_62774;
input v_63017;
input v_63260;
input v_63503;
input v_63746;
input v_63989;
input v_64232;
input v_64475;
input v_64718;
input v_64961;
input v_65204;
input v_65447;
input v_65690;
input v_65933;
input v_66176;
input v_66568;
input v_66828;
input v_67071;
input v_67314;
input v_67557;
input v_67800;
input v_68043;
input v_68286;
input v_68529;
input v_68772;
input v_69015;
input v_69258;
input v_69501;
input v_69744;
input v_69987;
input v_70230;
input v_70473;
input v_70716;
input v_4;
output o_1;
wire v_2;
wire v_3;
wire v_7;
wire v_8;
wire v_10;
wire v_11;
wire v_12;
wire v_14;
wire v_16;
wire v_17;
wire v_19;
wire v_21;
wire v_22;
wire v_24;
wire v_26;
wire v_27;
wire v_29;
wire v_31;
wire v_32;
wire v_34;
wire v_36;
wire v_37;
wire v_39;
wire v_41;
wire v_42;
wire v_44;
wire v_46;
wire v_47;
wire v_49;
wire v_51;
wire v_52;
wire v_54;
wire v_56;
wire v_57;
wire v_59;
wire v_61;
wire v_62;
wire v_64;
wire v_66;
wire v_67;
wire v_69;
wire v_71;
wire v_72;
wire v_74;
wire v_76;
wire v_77;
wire v_79;
wire v_81;
wire v_82;
wire v_84;
wire v_86;
wire v_87;
wire v_89;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_284;
wire v_285;
wire v_286;
wire v_288;
wire v_289;
wire v_290;
wire v_292;
wire v_293;
wire v_294;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_301;
wire v_302;
wire v_303;
wire v_305;
wire v_306;
wire v_307;
wire v_309;
wire v_310;
wire v_311;
wire v_313;
wire v_314;
wire v_315;
wire v_317;
wire v_318;
wire v_319;
wire v_321;
wire v_322;
wire v_323;
wire v_325;
wire v_326;
wire v_327;
wire v_329;
wire v_330;
wire v_331;
wire v_333;
wire v_334;
wire v_335;
wire v_337;
wire v_338;
wire v_339;
wire v_341;
wire v_342;
wire v_343;
wire v_345;
wire v_346;
wire v_347;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_452;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_459;
wire v_460;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_471;
wire v_472;
wire v_473;
wire v_474;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_481;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_496;
wire v_497;
wire v_498;
wire v_499;
wire v_500;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_511;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_544;
wire v_545;
wire v_546;
wire v_548;
wire v_549;
wire v_550;
wire v_552;
wire v_553;
wire v_554;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_561;
wire v_562;
wire v_563;
wire v_565;
wire v_566;
wire v_567;
wire v_569;
wire v_570;
wire v_571;
wire v_573;
wire v_574;
wire v_575;
wire v_577;
wire v_578;
wire v_579;
wire v_581;
wire v_582;
wire v_583;
wire v_585;
wire v_586;
wire v_587;
wire v_589;
wire v_590;
wire v_591;
wire v_593;
wire v_594;
wire v_595;
wire v_597;
wire v_598;
wire v_599;
wire v_601;
wire v_602;
wire v_603;
wire v_605;
wire v_606;
wire v_607;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_804;
wire v_805;
wire v_806;
wire v_808;
wire v_809;
wire v_810;
wire v_812;
wire v_813;
wire v_814;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_821;
wire v_822;
wire v_823;
wire v_825;
wire v_826;
wire v_827;
wire v_829;
wire v_830;
wire v_831;
wire v_833;
wire v_834;
wire v_835;
wire v_837;
wire v_838;
wire v_839;
wire v_841;
wire v_842;
wire v_843;
wire v_845;
wire v_846;
wire v_847;
wire v_849;
wire v_850;
wire v_851;
wire v_853;
wire v_854;
wire v_855;
wire v_857;
wire v_858;
wire v_859;
wire v_861;
wire v_862;
wire v_863;
wire v_865;
wire v_866;
wire v_867;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1008;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2116;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2121;
wire v_2122;
wire v_2123;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2157;
wire v_2158;
wire v_2159;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2169;
wire v_2170;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2181;
wire v_2182;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2218;
wire v_2219;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2226;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2265;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2364;
wire v_2365;
wire v_2366;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2744;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2755;
wire v_2756;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2764;
wire v_2765;
wire v_2766;
wire v_2767;
wire v_2768;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2786;
wire v_2787;
wire v_2788;
wire v_2789;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2795;
wire v_2796;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2804;
wire v_2805;
wire v_2806;
wire v_2807;
wire v_2808;
wire v_2809;
wire v_2810;
wire v_2811;
wire v_2812;
wire v_2813;
wire v_2814;
wire v_2815;
wire v_2816;
wire v_2817;
wire v_2818;
wire v_2819;
wire v_2820;
wire v_2821;
wire v_2822;
wire v_2823;
wire v_2824;
wire v_2825;
wire v_2826;
wire v_2827;
wire v_2828;
wire v_2829;
wire v_2830;
wire v_2831;
wire v_2832;
wire v_2833;
wire v_2834;
wire v_2835;
wire v_2836;
wire v_2837;
wire v_2838;
wire v_2839;
wire v_2840;
wire v_2841;
wire v_2842;
wire v_2843;
wire v_2844;
wire v_2845;
wire v_2846;
wire v_2847;
wire v_2848;
wire v_2849;
wire v_2850;
wire v_2851;
wire v_2852;
wire v_2853;
wire v_2854;
wire v_2855;
wire v_2856;
wire v_2857;
wire v_2858;
wire v_2859;
wire v_2860;
wire v_2861;
wire v_2862;
wire v_2863;
wire v_2864;
wire v_2865;
wire v_2866;
wire v_2867;
wire v_2868;
wire v_2869;
wire v_2870;
wire v_2871;
wire v_2872;
wire v_2873;
wire v_2874;
wire v_2875;
wire v_2876;
wire v_2877;
wire v_2878;
wire v_2879;
wire v_2880;
wire v_2881;
wire v_2884;
wire v_2885;
wire v_2886;
wire v_2888;
wire v_2889;
wire v_2890;
wire v_2892;
wire v_2893;
wire v_2894;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2899;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2921;
wire v_2922;
wire v_2923;
wire v_2925;
wire v_2926;
wire v_2927;
wire v_2929;
wire v_2930;
wire v_2931;
wire v_2933;
wire v_2934;
wire v_2935;
wire v_2937;
wire v_2938;
wire v_2939;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2945;
wire v_2946;
wire v_2947;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2952;
wire v_2953;
wire v_2954;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2967;
wire v_2968;
wire v_2969;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2988;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3011;
wire v_3012;
wire v_3013;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3023;
wire v_3024;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3028;
wire v_3029;
wire v_3030;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3035;
wire v_3036;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3044;
wire v_3045;
wire v_3046;
wire v_3047;
wire v_3048;
wire v_3049;
wire v_3050;
wire v_3051;
wire v_3052;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3059;
wire v_3060;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3071;
wire v_3072;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3080;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3088;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3099;
wire v_3100;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3109;
wire v_3110;
wire v_3111;
wire v_3112;
wire v_3113;
wire v_3114;
wire v_3115;
wire v_3116;
wire v_3117;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3134;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3139;
wire v_3140;
wire v_3141;
wire v_3144;
wire v_3145;
wire v_3146;
wire v_3148;
wire v_3149;
wire v_3150;
wire v_3152;
wire v_3153;
wire v_3154;
wire v_3156;
wire v_3157;
wire v_3158;
wire v_3159;
wire v_3161;
wire v_3162;
wire v_3163;
wire v_3165;
wire v_3166;
wire v_3167;
wire v_3169;
wire v_3170;
wire v_3171;
wire v_3173;
wire v_3174;
wire v_3175;
wire v_3177;
wire v_3178;
wire v_3179;
wire v_3181;
wire v_3182;
wire v_3183;
wire v_3185;
wire v_3186;
wire v_3187;
wire v_3189;
wire v_3190;
wire v_3191;
wire v_3193;
wire v_3194;
wire v_3195;
wire v_3197;
wire v_3198;
wire v_3199;
wire v_3201;
wire v_3202;
wire v_3203;
wire v_3205;
wire v_3206;
wire v_3207;
wire v_3209;
wire v_3210;
wire v_3211;
wire v_3212;
wire v_3213;
wire v_3214;
wire v_3215;
wire v_3216;
wire v_3217;
wire v_3218;
wire v_3219;
wire v_3220;
wire v_3221;
wire v_3222;
wire v_3223;
wire v_3224;
wire v_3225;
wire v_3226;
wire v_3227;
wire v_3228;
wire v_3229;
wire v_3230;
wire v_3231;
wire v_3232;
wire v_3233;
wire v_3234;
wire v_3235;
wire v_3236;
wire v_3237;
wire v_3238;
wire v_3239;
wire v_3240;
wire v_3241;
wire v_3242;
wire v_3243;
wire v_3244;
wire v_3245;
wire v_3246;
wire v_3247;
wire v_3248;
wire v_3249;
wire v_3250;
wire v_3251;
wire v_3252;
wire v_3253;
wire v_3254;
wire v_3255;
wire v_3256;
wire v_3257;
wire v_3258;
wire v_3259;
wire v_3260;
wire v_3261;
wire v_3262;
wire v_3263;
wire v_3264;
wire v_3265;
wire v_3266;
wire v_3267;
wire v_3268;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3277;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3293;
wire v_3294;
wire v_3295;
wire v_3296;
wire v_3297;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3305;
wire v_3306;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3315;
wire v_3316;
wire v_3317;
wire v_3318;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3329;
wire v_3330;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3341;
wire v_3342;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3348;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3353;
wire v_3354;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire v_3364;
wire v_3365;
wire v_3366;
wire v_3367;
wire v_3368;
wire v_3369;
wire v_3370;
wire v_3371;
wire v_3372;
wire v_3373;
wire v_3374;
wire v_3375;
wire v_3376;
wire v_3377;
wire v_3378;
wire v_3379;
wire v_3380;
wire v_3381;
wire v_3382;
wire v_3383;
wire v_3384;
wire v_3385;
wire v_3386;
wire v_3387;
wire v_3388;
wire v_3389;
wire v_3390;
wire v_3391;
wire v_3392;
wire v_3393;
wire v_3394;
wire v_3395;
wire v_3396;
wire v_3397;
wire v_3398;
wire v_3399;
wire v_3400;
wire v_3401;
wire v_3404;
wire v_3405;
wire v_3406;
wire v_3408;
wire v_3409;
wire v_3410;
wire v_3412;
wire v_3413;
wire v_3414;
wire v_3416;
wire v_3417;
wire v_3418;
wire v_3419;
wire v_3421;
wire v_3422;
wire v_3423;
wire v_3425;
wire v_3426;
wire v_3427;
wire v_3429;
wire v_3430;
wire v_3431;
wire v_3433;
wire v_3434;
wire v_3435;
wire v_3437;
wire v_3438;
wire v_3439;
wire v_3441;
wire v_3442;
wire v_3443;
wire v_3445;
wire v_3446;
wire v_3447;
wire v_3449;
wire v_3450;
wire v_3451;
wire v_3453;
wire v_3454;
wire v_3455;
wire v_3457;
wire v_3458;
wire v_3459;
wire v_3461;
wire v_3462;
wire v_3463;
wire v_3465;
wire v_3466;
wire v_3467;
wire v_3469;
wire v_3470;
wire v_3471;
wire v_3472;
wire v_3473;
wire v_3474;
wire v_3475;
wire v_3476;
wire v_3477;
wire v_3478;
wire v_3479;
wire v_3480;
wire v_3481;
wire v_3482;
wire v_3483;
wire v_3484;
wire v_3485;
wire v_3486;
wire v_3487;
wire v_3488;
wire v_3489;
wire v_3490;
wire v_3491;
wire v_3492;
wire v_3493;
wire v_3494;
wire v_3495;
wire v_3496;
wire v_3497;
wire v_3498;
wire v_3499;
wire v_3500;
wire v_3501;
wire v_3502;
wire v_3503;
wire v_3504;
wire v_3505;
wire v_3506;
wire v_3507;
wire v_3508;
wire v_3509;
wire v_3510;
wire v_3511;
wire v_3512;
wire v_3513;
wire v_3514;
wire v_3515;
wire v_3516;
wire v_3517;
wire v_3518;
wire v_3519;
wire v_3520;
wire v_3521;
wire v_3522;
wire v_3523;
wire v_3524;
wire v_3525;
wire v_3526;
wire v_3527;
wire v_3528;
wire v_3529;
wire v_3530;
wire v_3531;
wire v_3532;
wire v_3533;
wire v_3534;
wire v_3535;
wire v_3536;
wire v_3537;
wire v_3538;
wire v_3539;
wire v_3540;
wire v_3541;
wire v_3542;
wire v_3543;
wire v_3544;
wire v_3545;
wire v_3546;
wire v_3547;
wire v_3548;
wire v_3549;
wire v_3550;
wire v_3551;
wire v_3552;
wire v_3553;
wire v_3554;
wire v_3555;
wire v_3556;
wire v_3557;
wire v_3558;
wire v_3559;
wire v_3560;
wire v_3561;
wire v_3562;
wire v_3563;
wire v_3564;
wire v_3565;
wire v_3566;
wire v_3567;
wire v_3568;
wire v_3569;
wire v_3570;
wire v_3571;
wire v_3572;
wire v_3573;
wire v_3574;
wire v_3575;
wire v_3576;
wire v_3577;
wire v_3578;
wire v_3579;
wire v_3580;
wire v_3581;
wire v_3582;
wire v_3583;
wire v_3584;
wire v_3585;
wire v_3586;
wire v_3587;
wire v_3588;
wire v_3589;
wire v_3590;
wire v_3591;
wire v_3592;
wire v_3593;
wire v_3594;
wire v_3595;
wire v_3596;
wire v_3597;
wire v_3598;
wire v_3599;
wire v_3600;
wire v_3601;
wire v_3602;
wire v_3603;
wire v_3604;
wire v_3605;
wire v_3606;
wire v_3607;
wire v_3608;
wire v_3609;
wire v_3610;
wire v_3611;
wire v_3612;
wire v_3613;
wire v_3614;
wire v_3615;
wire v_3616;
wire v_3617;
wire v_3618;
wire v_3619;
wire v_3620;
wire v_3621;
wire v_3622;
wire v_3623;
wire v_3624;
wire v_3625;
wire v_3626;
wire v_3627;
wire v_3628;
wire v_3629;
wire v_3630;
wire v_3631;
wire v_3632;
wire v_3633;
wire v_3634;
wire v_3635;
wire v_3636;
wire v_3637;
wire v_3638;
wire v_3639;
wire v_3640;
wire v_3641;
wire v_3642;
wire v_3643;
wire v_3644;
wire v_3645;
wire v_3646;
wire v_3647;
wire v_3648;
wire v_3649;
wire v_3650;
wire v_3651;
wire v_3652;
wire v_3653;
wire v_3654;
wire v_3655;
wire v_3656;
wire v_3657;
wire v_3658;
wire v_3659;
wire v_3660;
wire v_3661;
wire v_3664;
wire v_3665;
wire v_3666;
wire v_3668;
wire v_3669;
wire v_3670;
wire v_3672;
wire v_3673;
wire v_3674;
wire v_3676;
wire v_3677;
wire v_3678;
wire v_3679;
wire v_3681;
wire v_3682;
wire v_3683;
wire v_3685;
wire v_3686;
wire v_3687;
wire v_3689;
wire v_3690;
wire v_3691;
wire v_3693;
wire v_3694;
wire v_3695;
wire v_3697;
wire v_3698;
wire v_3699;
wire v_3701;
wire v_3702;
wire v_3703;
wire v_3705;
wire v_3706;
wire v_3707;
wire v_3709;
wire v_3710;
wire v_3711;
wire v_3713;
wire v_3714;
wire v_3715;
wire v_3717;
wire v_3718;
wire v_3719;
wire v_3721;
wire v_3722;
wire v_3723;
wire v_3725;
wire v_3726;
wire v_3727;
wire v_3729;
wire v_3730;
wire v_3731;
wire v_3732;
wire v_3733;
wire v_3734;
wire v_3735;
wire v_3736;
wire v_3737;
wire v_3738;
wire v_3739;
wire v_3740;
wire v_3741;
wire v_3742;
wire v_3743;
wire v_3744;
wire v_3745;
wire v_3746;
wire v_3747;
wire v_3748;
wire v_3749;
wire v_3750;
wire v_3751;
wire v_3752;
wire v_3753;
wire v_3754;
wire v_3755;
wire v_3756;
wire v_3757;
wire v_3758;
wire v_3759;
wire v_3760;
wire v_3761;
wire v_3762;
wire v_3763;
wire v_3764;
wire v_3765;
wire v_3766;
wire v_3767;
wire v_3768;
wire v_3769;
wire v_3770;
wire v_3771;
wire v_3772;
wire v_3773;
wire v_3774;
wire v_3775;
wire v_3776;
wire v_3777;
wire v_3778;
wire v_3779;
wire v_3780;
wire v_3781;
wire v_3782;
wire v_3783;
wire v_3784;
wire v_3785;
wire v_3786;
wire v_3787;
wire v_3788;
wire v_3789;
wire v_3790;
wire v_3791;
wire v_3792;
wire v_3793;
wire v_3794;
wire v_3795;
wire v_3796;
wire v_3797;
wire v_3798;
wire v_3799;
wire v_3800;
wire v_3801;
wire v_3802;
wire v_3803;
wire v_3804;
wire v_3805;
wire v_3806;
wire v_3807;
wire v_3808;
wire v_3809;
wire v_3810;
wire v_3811;
wire v_3812;
wire v_3813;
wire v_3814;
wire v_3815;
wire v_3816;
wire v_3817;
wire v_3818;
wire v_3819;
wire v_3820;
wire v_3821;
wire v_3822;
wire v_3823;
wire v_3824;
wire v_3825;
wire v_3826;
wire v_3827;
wire v_3828;
wire v_3829;
wire v_3830;
wire v_3831;
wire v_3832;
wire v_3833;
wire v_3834;
wire v_3835;
wire v_3836;
wire v_3837;
wire v_3838;
wire v_3839;
wire v_3840;
wire v_3841;
wire v_3842;
wire v_3843;
wire v_3844;
wire v_3845;
wire v_3846;
wire v_3847;
wire v_3848;
wire v_3849;
wire v_3850;
wire v_3851;
wire v_3852;
wire v_3853;
wire v_3854;
wire v_3855;
wire v_3856;
wire v_3857;
wire v_3858;
wire v_3859;
wire v_3860;
wire v_3861;
wire v_3862;
wire v_3863;
wire v_3864;
wire v_3865;
wire v_3866;
wire v_3867;
wire v_3868;
wire v_3869;
wire v_3870;
wire v_3871;
wire v_3872;
wire v_3873;
wire v_3874;
wire v_3875;
wire v_3876;
wire v_3877;
wire v_3878;
wire v_3879;
wire v_3880;
wire v_3881;
wire v_3882;
wire v_3883;
wire v_3884;
wire v_3885;
wire v_3886;
wire v_3887;
wire v_3888;
wire v_3889;
wire v_3890;
wire v_3891;
wire v_3892;
wire v_3893;
wire v_3894;
wire v_3895;
wire v_3896;
wire v_3897;
wire v_3898;
wire v_3899;
wire v_3900;
wire v_3901;
wire v_3902;
wire v_3903;
wire v_3904;
wire v_3905;
wire v_3906;
wire v_3907;
wire v_3908;
wire v_3909;
wire v_3910;
wire v_3911;
wire v_3912;
wire v_3913;
wire v_3914;
wire v_3915;
wire v_3916;
wire v_3917;
wire v_3918;
wire v_3919;
wire v_3920;
wire v_3921;
wire v_3924;
wire v_3925;
wire v_3926;
wire v_3928;
wire v_3929;
wire v_3930;
wire v_3932;
wire v_3933;
wire v_3934;
wire v_3936;
wire v_3937;
wire v_3938;
wire v_3939;
wire v_3941;
wire v_3942;
wire v_3943;
wire v_3945;
wire v_3946;
wire v_3947;
wire v_3949;
wire v_3950;
wire v_3951;
wire v_3953;
wire v_3954;
wire v_3955;
wire v_3957;
wire v_3958;
wire v_3959;
wire v_3961;
wire v_3962;
wire v_3963;
wire v_3965;
wire v_3966;
wire v_3967;
wire v_3969;
wire v_3970;
wire v_3971;
wire v_3973;
wire v_3974;
wire v_3975;
wire v_3977;
wire v_3978;
wire v_3979;
wire v_3981;
wire v_3982;
wire v_3983;
wire v_3985;
wire v_3986;
wire v_3987;
wire v_3989;
wire v_3990;
wire v_3991;
wire v_3992;
wire v_3993;
wire v_3994;
wire v_3995;
wire v_3996;
wire v_3997;
wire v_3998;
wire v_3999;
wire v_4000;
wire v_4001;
wire v_4002;
wire v_4003;
wire v_4004;
wire v_4005;
wire v_4006;
wire v_4007;
wire v_4008;
wire v_4009;
wire v_4010;
wire v_4011;
wire v_4012;
wire v_4013;
wire v_4014;
wire v_4015;
wire v_4016;
wire v_4017;
wire v_4018;
wire v_4019;
wire v_4020;
wire v_4021;
wire v_4022;
wire v_4023;
wire v_4024;
wire v_4025;
wire v_4026;
wire v_4027;
wire v_4028;
wire v_4029;
wire v_4030;
wire v_4031;
wire v_4032;
wire v_4033;
wire v_4034;
wire v_4035;
wire v_4036;
wire v_4037;
wire v_4038;
wire v_4039;
wire v_4040;
wire v_4041;
wire v_4042;
wire v_4043;
wire v_4044;
wire v_4045;
wire v_4046;
wire v_4047;
wire v_4048;
wire v_4049;
wire v_4050;
wire v_4051;
wire v_4052;
wire v_4053;
wire v_4054;
wire v_4055;
wire v_4056;
wire v_4057;
wire v_4058;
wire v_4059;
wire v_4060;
wire v_4061;
wire v_4062;
wire v_4063;
wire v_4064;
wire v_4065;
wire v_4066;
wire v_4067;
wire v_4068;
wire v_4069;
wire v_4070;
wire v_4071;
wire v_4072;
wire v_4073;
wire v_4074;
wire v_4075;
wire v_4076;
wire v_4077;
wire v_4078;
wire v_4079;
wire v_4080;
wire v_4081;
wire v_4082;
wire v_4083;
wire v_4084;
wire v_4085;
wire v_4086;
wire v_4087;
wire v_4088;
wire v_4089;
wire v_4090;
wire v_4091;
wire v_4092;
wire v_4093;
wire v_4094;
wire v_4095;
wire v_4096;
wire v_4097;
wire v_4098;
wire v_4099;
wire v_4100;
wire v_4101;
wire v_4102;
wire v_4103;
wire v_4104;
wire v_4105;
wire v_4106;
wire v_4107;
wire v_4108;
wire v_4109;
wire v_4110;
wire v_4111;
wire v_4112;
wire v_4113;
wire v_4114;
wire v_4115;
wire v_4116;
wire v_4117;
wire v_4118;
wire v_4119;
wire v_4120;
wire v_4121;
wire v_4122;
wire v_4123;
wire v_4124;
wire v_4125;
wire v_4126;
wire v_4127;
wire v_4128;
wire v_4129;
wire v_4130;
wire v_4131;
wire v_4132;
wire v_4133;
wire v_4134;
wire v_4135;
wire v_4136;
wire v_4137;
wire v_4138;
wire v_4139;
wire v_4140;
wire v_4141;
wire v_4142;
wire v_4143;
wire v_4144;
wire v_4145;
wire v_4146;
wire v_4147;
wire v_4148;
wire v_4149;
wire v_4150;
wire v_4151;
wire v_4152;
wire v_4153;
wire v_4154;
wire v_4155;
wire v_4156;
wire v_4157;
wire v_4158;
wire v_4159;
wire v_4160;
wire v_4161;
wire v_4162;
wire v_4163;
wire v_4164;
wire v_4165;
wire v_4166;
wire v_4167;
wire v_4168;
wire v_4169;
wire v_4170;
wire v_4171;
wire v_4172;
wire v_4173;
wire v_4174;
wire v_4175;
wire v_4176;
wire v_4177;
wire v_4178;
wire v_4179;
wire v_4180;
wire v_4181;
wire v_4183;
wire v_4184;
wire v_4185;
wire v_4187;
wire v_4188;
wire v_4189;
wire v_4191;
wire v_4192;
wire v_4193;
wire v_4195;
wire v_4196;
wire v_4197;
wire v_4198;
wire v_4200;
wire v_4201;
wire v_4202;
wire v_4204;
wire v_4205;
wire v_4206;
wire v_4208;
wire v_4209;
wire v_4210;
wire v_4212;
wire v_4213;
wire v_4214;
wire v_4216;
wire v_4217;
wire v_4218;
wire v_4220;
wire v_4221;
wire v_4222;
wire v_4224;
wire v_4225;
wire v_4226;
wire v_4228;
wire v_4229;
wire v_4230;
wire v_4232;
wire v_4233;
wire v_4234;
wire v_4236;
wire v_4237;
wire v_4238;
wire v_4240;
wire v_4241;
wire v_4242;
wire v_4244;
wire v_4245;
wire v_4246;
wire v_4248;
wire v_4249;
wire v_4250;
wire v_4251;
wire v_4252;
wire v_4253;
wire v_4254;
wire v_4255;
wire v_4256;
wire v_4257;
wire v_4258;
wire v_4259;
wire v_4260;
wire v_4261;
wire v_4262;
wire v_4263;
wire v_4264;
wire v_4265;
wire v_4266;
wire v_4267;
wire v_4268;
wire v_4269;
wire v_4270;
wire v_4271;
wire v_4272;
wire v_4273;
wire v_4274;
wire v_4275;
wire v_4276;
wire v_4277;
wire v_4278;
wire v_4279;
wire v_4280;
wire v_4281;
wire v_4282;
wire v_4283;
wire v_4284;
wire v_4285;
wire v_4286;
wire v_4287;
wire v_4288;
wire v_4289;
wire v_4290;
wire v_4291;
wire v_4292;
wire v_4293;
wire v_4294;
wire v_4295;
wire v_4296;
wire v_4297;
wire v_4298;
wire v_4299;
wire v_4300;
wire v_4301;
wire v_4302;
wire v_4303;
wire v_4304;
wire v_4305;
wire v_4306;
wire v_4307;
wire v_4308;
wire v_4309;
wire v_4310;
wire v_4311;
wire v_4312;
wire v_4313;
wire v_4314;
wire v_4315;
wire v_4316;
wire v_4317;
wire v_4318;
wire v_4319;
wire v_4320;
wire v_4321;
wire v_4322;
wire v_4323;
wire v_4324;
wire v_4325;
wire v_4326;
wire v_4327;
wire v_4328;
wire v_4329;
wire v_4330;
wire v_4331;
wire v_4332;
wire v_4333;
wire v_4334;
wire v_4335;
wire v_4336;
wire v_4337;
wire v_4338;
wire v_4339;
wire v_4340;
wire v_4341;
wire v_4342;
wire v_4343;
wire v_4344;
wire v_4345;
wire v_4346;
wire v_4347;
wire v_4349;
wire v_4350;
wire v_4351;
wire v_4352;
wire v_4353;
wire v_4354;
wire v_4355;
wire v_4356;
wire v_4357;
wire v_4358;
wire v_4359;
wire v_4360;
wire v_4361;
wire v_4362;
wire v_4363;
wire v_4364;
wire v_4365;
wire v_4366;
wire v_4367;
wire v_4368;
wire v_4369;
wire v_4370;
wire v_4371;
wire v_4372;
wire v_4373;
wire v_4374;
wire v_4375;
wire v_4376;
wire v_4377;
wire v_4378;
wire v_4379;
wire v_4380;
wire v_4381;
wire v_4382;
wire v_4383;
wire v_4384;
wire v_4385;
wire v_4386;
wire v_4387;
wire v_4388;
wire v_4389;
wire v_4390;
wire v_4391;
wire v_4392;
wire v_4393;
wire v_4394;
wire v_4395;
wire v_4396;
wire v_4397;
wire v_4398;
wire v_4399;
wire v_4400;
wire v_4401;
wire v_4402;
wire v_4403;
wire v_4404;
wire v_4405;
wire v_4406;
wire v_4407;
wire v_4408;
wire v_4409;
wire v_4410;
wire v_4411;
wire v_4412;
wire v_4413;
wire v_4414;
wire v_4415;
wire v_4416;
wire v_4417;
wire v_4418;
wire v_4419;
wire v_4420;
wire v_4421;
wire v_4422;
wire v_4423;
wire v_4424;
wire v_4425;
wire v_4426;
wire v_4427;
wire v_4428;
wire v_4429;
wire v_4430;
wire v_4431;
wire v_4432;
wire v_4433;
wire v_4434;
wire v_4435;
wire v_4436;
wire v_4437;
wire v_4438;
wire v_4439;
wire v_4440;
wire v_4441;
wire v_4443;
wire v_4445;
wire v_4446;
wire v_4447;
wire v_4449;
wire v_4450;
wire v_4451;
wire v_4453;
wire v_4454;
wire v_4455;
wire v_4457;
wire v_4458;
wire v_4460;
wire v_4461;
wire v_4462;
wire v_4464;
wire v_4465;
wire v_4466;
wire v_4468;
wire v_4469;
wire v_4470;
wire v_4472;
wire v_4473;
wire v_4474;
wire v_4476;
wire v_4477;
wire v_4478;
wire v_4480;
wire v_4481;
wire v_4482;
wire v_4484;
wire v_4485;
wire v_4486;
wire v_4488;
wire v_4489;
wire v_4490;
wire v_4492;
wire v_4493;
wire v_4494;
wire v_4496;
wire v_4497;
wire v_4498;
wire v_4500;
wire v_4501;
wire v_4502;
wire v_4504;
wire v_4505;
wire v_4506;
wire v_4508;
wire v_4509;
wire v_4510;
wire v_4511;
wire v_4512;
wire v_4513;
wire v_4514;
wire v_4515;
wire v_4516;
wire v_4517;
wire v_4518;
wire v_4519;
wire v_4520;
wire v_4521;
wire v_4522;
wire v_4523;
wire v_4524;
wire v_4525;
wire v_4526;
wire v_4527;
wire v_4528;
wire v_4529;
wire v_4530;
wire v_4531;
wire v_4532;
wire v_4533;
wire v_4534;
wire v_4535;
wire v_4536;
wire v_4537;
wire v_4538;
wire v_4539;
wire v_4540;
wire v_4541;
wire v_4542;
wire v_4543;
wire v_4544;
wire v_4545;
wire v_4546;
wire v_4547;
wire v_4548;
wire v_4549;
wire v_4550;
wire v_4551;
wire v_4552;
wire v_4553;
wire v_4554;
wire v_4555;
wire v_4556;
wire v_4557;
wire v_4558;
wire v_4559;
wire v_4560;
wire v_4561;
wire v_4562;
wire v_4563;
wire v_4564;
wire v_4565;
wire v_4566;
wire v_4567;
wire v_4568;
wire v_4569;
wire v_4570;
wire v_4571;
wire v_4572;
wire v_4573;
wire v_4574;
wire v_4575;
wire v_4576;
wire v_4577;
wire v_4578;
wire v_4579;
wire v_4580;
wire v_4581;
wire v_4582;
wire v_4583;
wire v_4584;
wire v_4585;
wire v_4586;
wire v_4587;
wire v_4588;
wire v_4589;
wire v_4590;
wire v_4591;
wire v_4592;
wire v_4593;
wire v_4594;
wire v_4595;
wire v_4596;
wire v_4597;
wire v_4598;
wire v_4599;
wire v_4600;
wire v_4601;
wire v_4602;
wire v_4603;
wire v_4604;
wire v_4605;
wire v_4606;
wire v_4607;
wire v_4608;
wire v_4609;
wire v_4610;
wire v_4611;
wire v_4612;
wire v_4613;
wire v_4614;
wire v_4615;
wire v_4616;
wire v_4617;
wire v_4618;
wire v_4619;
wire v_4620;
wire v_4621;
wire v_4622;
wire v_4623;
wire v_4624;
wire v_4625;
wire v_4626;
wire v_4627;
wire v_4628;
wire v_4629;
wire v_4630;
wire v_4631;
wire v_4632;
wire v_4633;
wire v_4634;
wire v_4635;
wire v_4636;
wire v_4637;
wire v_4638;
wire v_4639;
wire v_4640;
wire v_4641;
wire v_4642;
wire v_4643;
wire v_4644;
wire v_4645;
wire v_4646;
wire v_4647;
wire v_4648;
wire v_4649;
wire v_4650;
wire v_4651;
wire v_4652;
wire v_4653;
wire v_4654;
wire v_4655;
wire v_4656;
wire v_4657;
wire v_4658;
wire v_4659;
wire v_4660;
wire v_4661;
wire v_4662;
wire v_4663;
wire v_4664;
wire v_4665;
wire v_4666;
wire v_4667;
wire v_4668;
wire v_4669;
wire v_4670;
wire v_4671;
wire v_4672;
wire v_4673;
wire v_4674;
wire v_4675;
wire v_4676;
wire v_4677;
wire v_4678;
wire v_4679;
wire v_4680;
wire v_4681;
wire v_4682;
wire v_4683;
wire v_4684;
wire v_4685;
wire v_4686;
wire v_4687;
wire v_4688;
wire v_4689;
wire v_4690;
wire v_4691;
wire v_4692;
wire v_4693;
wire v_4694;
wire v_4695;
wire v_4696;
wire v_4697;
wire v_4698;
wire v_4699;
wire v_4700;
wire v_4701;
wire v_4703;
wire v_4704;
wire v_4705;
wire v_4706;
wire v_4707;
wire v_4708;
wire v_4709;
wire v_4710;
wire v_4711;
wire v_4712;
wire v_4713;
wire v_4714;
wire v_4715;
wire v_4716;
wire v_4717;
wire v_4718;
wire v_4719;
wire v_4720;
wire v_4721;
wire v_4722;
wire v_4723;
wire v_4724;
wire v_4725;
wire v_4726;
wire v_4727;
wire v_4728;
wire v_4729;
wire v_4730;
wire v_4731;
wire v_4732;
wire v_4733;
wire v_4734;
wire v_4735;
wire v_4736;
wire v_4737;
wire v_4738;
wire v_4739;
wire v_4740;
wire v_4741;
wire v_4742;
wire v_4743;
wire v_4744;
wire v_4745;
wire v_4746;
wire v_4747;
wire v_4748;
wire v_4749;
wire v_4750;
wire v_4751;
wire v_4752;
wire v_4753;
wire v_4754;
wire v_4755;
wire v_4756;
wire v_4757;
wire v_4758;
wire v_4759;
wire v_4760;
wire v_4761;
wire v_4762;
wire v_4763;
wire v_4764;
wire v_4765;
wire v_4766;
wire v_4767;
wire v_4768;
wire v_4769;
wire v_4770;
wire v_4771;
wire v_4772;
wire v_4773;
wire v_4774;
wire v_4775;
wire v_4776;
wire v_4777;
wire v_4778;
wire v_4779;
wire v_4780;
wire v_4781;
wire v_4782;
wire v_4783;
wire v_4784;
wire v_4785;
wire v_4786;
wire v_4787;
wire v_4788;
wire v_4789;
wire v_4790;
wire v_4791;
wire v_4792;
wire v_4793;
wire v_4794;
wire v_4795;
wire v_4796;
wire v_4797;
wire v_4798;
wire v_4799;
wire v_4800;
wire v_4801;
wire v_4802;
wire v_4803;
wire v_4804;
wire v_4805;
wire v_4806;
wire v_4807;
wire v_4808;
wire v_4809;
wire v_4810;
wire v_4811;
wire v_4812;
wire v_4813;
wire v_4814;
wire v_4815;
wire v_4816;
wire v_4817;
wire v_4818;
wire v_4819;
wire v_4820;
wire v_4821;
wire v_4822;
wire v_4823;
wire v_4824;
wire v_4825;
wire v_4826;
wire v_4827;
wire v_4828;
wire v_4829;
wire v_4830;
wire v_4831;
wire v_4832;
wire v_4833;
wire v_4834;
wire v_4835;
wire v_4836;
wire v_4837;
wire v_4838;
wire v_4839;
wire v_4840;
wire v_4841;
wire v_4842;
wire v_4843;
wire v_4844;
wire v_4845;
wire v_4846;
wire v_4847;
wire v_4848;
wire v_4849;
wire v_4850;
wire v_4851;
wire v_4852;
wire v_4853;
wire v_4854;
wire v_4855;
wire v_4856;
wire v_4857;
wire v_4858;
wire v_4859;
wire v_4860;
wire v_4861;
wire v_4862;
wire v_4863;
wire v_4864;
wire v_4865;
wire v_4866;
wire v_4867;
wire v_4868;
wire v_4869;
wire v_4870;
wire v_4871;
wire v_4872;
wire v_4873;
wire v_4874;
wire v_4875;
wire v_4876;
wire v_4877;
wire v_4878;
wire v_4879;
wire v_4880;
wire v_4881;
wire v_4882;
wire v_4883;
wire v_4884;
wire v_4885;
wire v_4886;
wire v_4887;
wire v_4888;
wire v_4889;
wire v_4890;
wire v_4891;
wire v_4892;
wire v_4893;
wire v_4894;
wire v_4895;
wire v_4896;
wire v_4897;
wire v_4898;
wire v_4899;
wire v_4900;
wire v_4901;
wire v_4902;
wire v_4903;
wire v_4904;
wire v_4905;
wire v_4906;
wire v_4907;
wire v_4908;
wire v_4909;
wire v_4910;
wire v_4911;
wire v_4912;
wire v_4913;
wire v_4914;
wire v_4915;
wire v_4916;
wire v_4917;
wire v_4918;
wire v_4919;
wire v_4920;
wire v_4921;
wire v_4922;
wire v_4923;
wire v_4924;
wire v_4925;
wire v_4926;
wire v_4927;
wire v_4928;
wire v_4929;
wire v_4930;
wire v_4931;
wire v_4932;
wire v_4933;
wire v_4934;
wire v_4935;
wire v_4936;
wire v_4937;
wire v_4938;
wire v_4939;
wire v_4940;
wire v_4941;
wire v_4942;
wire v_4943;
wire v_4944;
wire v_4946;
wire v_4947;
wire v_4948;
wire v_4949;
wire v_4950;
wire v_4951;
wire v_4952;
wire v_4953;
wire v_4954;
wire v_4955;
wire v_4956;
wire v_4957;
wire v_4958;
wire v_4959;
wire v_4960;
wire v_4961;
wire v_4962;
wire v_4963;
wire v_4964;
wire v_4965;
wire v_4966;
wire v_4967;
wire v_4968;
wire v_4969;
wire v_4970;
wire v_4971;
wire v_4972;
wire v_4973;
wire v_4974;
wire v_4975;
wire v_4976;
wire v_4977;
wire v_4978;
wire v_4979;
wire v_4980;
wire v_4981;
wire v_4982;
wire v_4983;
wire v_4984;
wire v_4985;
wire v_4986;
wire v_4987;
wire v_4988;
wire v_4989;
wire v_4990;
wire v_4991;
wire v_4992;
wire v_4993;
wire v_4994;
wire v_4995;
wire v_4996;
wire v_4997;
wire v_4998;
wire v_4999;
wire v_5000;
wire v_5001;
wire v_5002;
wire v_5003;
wire v_5004;
wire v_5005;
wire v_5006;
wire v_5007;
wire v_5008;
wire v_5009;
wire v_5010;
wire v_5011;
wire v_5012;
wire v_5013;
wire v_5014;
wire v_5015;
wire v_5016;
wire v_5017;
wire v_5018;
wire v_5019;
wire v_5020;
wire v_5021;
wire v_5022;
wire v_5023;
wire v_5024;
wire v_5025;
wire v_5026;
wire v_5027;
wire v_5028;
wire v_5029;
wire v_5030;
wire v_5031;
wire v_5032;
wire v_5033;
wire v_5034;
wire v_5035;
wire v_5036;
wire v_5037;
wire v_5038;
wire v_5039;
wire v_5040;
wire v_5041;
wire v_5042;
wire v_5043;
wire v_5044;
wire v_5045;
wire v_5046;
wire v_5047;
wire v_5048;
wire v_5049;
wire v_5050;
wire v_5051;
wire v_5052;
wire v_5053;
wire v_5054;
wire v_5055;
wire v_5056;
wire v_5057;
wire v_5058;
wire v_5059;
wire v_5060;
wire v_5061;
wire v_5062;
wire v_5063;
wire v_5064;
wire v_5065;
wire v_5066;
wire v_5067;
wire v_5068;
wire v_5069;
wire v_5070;
wire v_5071;
wire v_5072;
wire v_5073;
wire v_5074;
wire v_5075;
wire v_5076;
wire v_5077;
wire v_5078;
wire v_5079;
wire v_5080;
wire v_5081;
wire v_5082;
wire v_5083;
wire v_5084;
wire v_5085;
wire v_5086;
wire v_5087;
wire v_5088;
wire v_5089;
wire v_5090;
wire v_5091;
wire v_5092;
wire v_5093;
wire v_5094;
wire v_5095;
wire v_5096;
wire v_5097;
wire v_5098;
wire v_5099;
wire v_5100;
wire v_5101;
wire v_5102;
wire v_5103;
wire v_5104;
wire v_5105;
wire v_5106;
wire v_5107;
wire v_5108;
wire v_5109;
wire v_5110;
wire v_5111;
wire v_5112;
wire v_5113;
wire v_5114;
wire v_5115;
wire v_5116;
wire v_5117;
wire v_5118;
wire v_5119;
wire v_5120;
wire v_5121;
wire v_5122;
wire v_5123;
wire v_5124;
wire v_5125;
wire v_5126;
wire v_5127;
wire v_5128;
wire v_5129;
wire v_5130;
wire v_5131;
wire v_5132;
wire v_5133;
wire v_5134;
wire v_5135;
wire v_5136;
wire v_5137;
wire v_5138;
wire v_5139;
wire v_5140;
wire v_5141;
wire v_5142;
wire v_5143;
wire v_5144;
wire v_5145;
wire v_5146;
wire v_5147;
wire v_5148;
wire v_5149;
wire v_5150;
wire v_5151;
wire v_5152;
wire v_5153;
wire v_5154;
wire v_5155;
wire v_5156;
wire v_5157;
wire v_5158;
wire v_5159;
wire v_5160;
wire v_5161;
wire v_5162;
wire v_5163;
wire v_5164;
wire v_5165;
wire v_5166;
wire v_5167;
wire v_5168;
wire v_5169;
wire v_5170;
wire v_5171;
wire v_5172;
wire v_5173;
wire v_5174;
wire v_5175;
wire v_5176;
wire v_5177;
wire v_5178;
wire v_5179;
wire v_5180;
wire v_5181;
wire v_5182;
wire v_5183;
wire v_5184;
wire v_5185;
wire v_5186;
wire v_5187;
wire v_5189;
wire v_5190;
wire v_5191;
wire v_5192;
wire v_5193;
wire v_5194;
wire v_5195;
wire v_5196;
wire v_5197;
wire v_5198;
wire v_5199;
wire v_5200;
wire v_5201;
wire v_5202;
wire v_5203;
wire v_5204;
wire v_5205;
wire v_5206;
wire v_5207;
wire v_5208;
wire v_5209;
wire v_5210;
wire v_5211;
wire v_5212;
wire v_5213;
wire v_5214;
wire v_5215;
wire v_5216;
wire v_5217;
wire v_5218;
wire v_5219;
wire v_5220;
wire v_5221;
wire v_5222;
wire v_5223;
wire v_5224;
wire v_5225;
wire v_5226;
wire v_5227;
wire v_5228;
wire v_5229;
wire v_5230;
wire v_5231;
wire v_5232;
wire v_5233;
wire v_5234;
wire v_5235;
wire v_5236;
wire v_5237;
wire v_5238;
wire v_5239;
wire v_5240;
wire v_5241;
wire v_5242;
wire v_5243;
wire v_5244;
wire v_5245;
wire v_5246;
wire v_5247;
wire v_5248;
wire v_5249;
wire v_5250;
wire v_5251;
wire v_5252;
wire v_5253;
wire v_5254;
wire v_5255;
wire v_5256;
wire v_5257;
wire v_5258;
wire v_5259;
wire v_5260;
wire v_5261;
wire v_5262;
wire v_5263;
wire v_5264;
wire v_5265;
wire v_5266;
wire v_5267;
wire v_5268;
wire v_5269;
wire v_5270;
wire v_5271;
wire v_5272;
wire v_5273;
wire v_5274;
wire v_5275;
wire v_5276;
wire v_5277;
wire v_5278;
wire v_5279;
wire v_5280;
wire v_5281;
wire v_5282;
wire v_5283;
wire v_5284;
wire v_5285;
wire v_5286;
wire v_5287;
wire v_5288;
wire v_5289;
wire v_5290;
wire v_5291;
wire v_5292;
wire v_5293;
wire v_5294;
wire v_5295;
wire v_5296;
wire v_5297;
wire v_5298;
wire v_5299;
wire v_5300;
wire v_5301;
wire v_5302;
wire v_5303;
wire v_5304;
wire v_5305;
wire v_5306;
wire v_5307;
wire v_5308;
wire v_5309;
wire v_5310;
wire v_5311;
wire v_5312;
wire v_5313;
wire v_5314;
wire v_5315;
wire v_5316;
wire v_5317;
wire v_5318;
wire v_5319;
wire v_5320;
wire v_5321;
wire v_5322;
wire v_5323;
wire v_5324;
wire v_5325;
wire v_5326;
wire v_5327;
wire v_5328;
wire v_5329;
wire v_5330;
wire v_5331;
wire v_5332;
wire v_5333;
wire v_5334;
wire v_5335;
wire v_5336;
wire v_5337;
wire v_5338;
wire v_5339;
wire v_5340;
wire v_5341;
wire v_5342;
wire v_5343;
wire v_5344;
wire v_5345;
wire v_5346;
wire v_5347;
wire v_5348;
wire v_5349;
wire v_5350;
wire v_5351;
wire v_5352;
wire v_5353;
wire v_5354;
wire v_5355;
wire v_5356;
wire v_5357;
wire v_5358;
wire v_5359;
wire v_5360;
wire v_5361;
wire v_5362;
wire v_5363;
wire v_5364;
wire v_5365;
wire v_5366;
wire v_5367;
wire v_5368;
wire v_5369;
wire v_5370;
wire v_5371;
wire v_5372;
wire v_5373;
wire v_5374;
wire v_5375;
wire v_5376;
wire v_5377;
wire v_5378;
wire v_5379;
wire v_5380;
wire v_5381;
wire v_5382;
wire v_5383;
wire v_5384;
wire v_5385;
wire v_5386;
wire v_5387;
wire v_5388;
wire v_5389;
wire v_5390;
wire v_5391;
wire v_5392;
wire v_5393;
wire v_5394;
wire v_5395;
wire v_5396;
wire v_5397;
wire v_5398;
wire v_5399;
wire v_5400;
wire v_5401;
wire v_5402;
wire v_5403;
wire v_5404;
wire v_5405;
wire v_5406;
wire v_5407;
wire v_5408;
wire v_5409;
wire v_5410;
wire v_5411;
wire v_5412;
wire v_5413;
wire v_5414;
wire v_5415;
wire v_5416;
wire v_5417;
wire v_5418;
wire v_5419;
wire v_5420;
wire v_5421;
wire v_5422;
wire v_5423;
wire v_5424;
wire v_5425;
wire v_5426;
wire v_5427;
wire v_5428;
wire v_5429;
wire v_5430;
wire v_5432;
wire v_5433;
wire v_5434;
wire v_5435;
wire v_5436;
wire v_5437;
wire v_5438;
wire v_5439;
wire v_5440;
wire v_5441;
wire v_5442;
wire v_5443;
wire v_5444;
wire v_5445;
wire v_5446;
wire v_5447;
wire v_5448;
wire v_5449;
wire v_5450;
wire v_5451;
wire v_5452;
wire v_5453;
wire v_5454;
wire v_5455;
wire v_5456;
wire v_5457;
wire v_5458;
wire v_5459;
wire v_5460;
wire v_5461;
wire v_5462;
wire v_5463;
wire v_5464;
wire v_5465;
wire v_5466;
wire v_5467;
wire v_5468;
wire v_5469;
wire v_5470;
wire v_5471;
wire v_5472;
wire v_5473;
wire v_5474;
wire v_5475;
wire v_5476;
wire v_5477;
wire v_5478;
wire v_5479;
wire v_5480;
wire v_5481;
wire v_5482;
wire v_5483;
wire v_5484;
wire v_5485;
wire v_5486;
wire v_5487;
wire v_5488;
wire v_5489;
wire v_5490;
wire v_5491;
wire v_5492;
wire v_5493;
wire v_5494;
wire v_5495;
wire v_5496;
wire v_5497;
wire v_5498;
wire v_5499;
wire v_5500;
wire v_5501;
wire v_5502;
wire v_5503;
wire v_5504;
wire v_5505;
wire v_5506;
wire v_5507;
wire v_5508;
wire v_5509;
wire v_5510;
wire v_5511;
wire v_5512;
wire v_5513;
wire v_5514;
wire v_5515;
wire v_5516;
wire v_5517;
wire v_5518;
wire v_5519;
wire v_5520;
wire v_5521;
wire v_5522;
wire v_5523;
wire v_5524;
wire v_5525;
wire v_5526;
wire v_5527;
wire v_5528;
wire v_5529;
wire v_5530;
wire v_5531;
wire v_5532;
wire v_5533;
wire v_5534;
wire v_5535;
wire v_5536;
wire v_5537;
wire v_5538;
wire v_5539;
wire v_5540;
wire v_5541;
wire v_5542;
wire v_5543;
wire v_5544;
wire v_5545;
wire v_5546;
wire v_5547;
wire v_5548;
wire v_5549;
wire v_5550;
wire v_5551;
wire v_5552;
wire v_5553;
wire v_5554;
wire v_5555;
wire v_5556;
wire v_5557;
wire v_5558;
wire v_5559;
wire v_5560;
wire v_5561;
wire v_5562;
wire v_5563;
wire v_5564;
wire v_5565;
wire v_5566;
wire v_5567;
wire v_5568;
wire v_5569;
wire v_5570;
wire v_5571;
wire v_5572;
wire v_5573;
wire v_5574;
wire v_5575;
wire v_5576;
wire v_5577;
wire v_5578;
wire v_5579;
wire v_5580;
wire v_5581;
wire v_5582;
wire v_5583;
wire v_5584;
wire v_5585;
wire v_5586;
wire v_5587;
wire v_5588;
wire v_5589;
wire v_5590;
wire v_5591;
wire v_5592;
wire v_5593;
wire v_5594;
wire v_5595;
wire v_5596;
wire v_5597;
wire v_5598;
wire v_5599;
wire v_5600;
wire v_5601;
wire v_5602;
wire v_5603;
wire v_5604;
wire v_5605;
wire v_5606;
wire v_5607;
wire v_5608;
wire v_5609;
wire v_5610;
wire v_5611;
wire v_5612;
wire v_5613;
wire v_5614;
wire v_5615;
wire v_5616;
wire v_5617;
wire v_5618;
wire v_5619;
wire v_5620;
wire v_5621;
wire v_5622;
wire v_5623;
wire v_5624;
wire v_5625;
wire v_5626;
wire v_5627;
wire v_5628;
wire v_5629;
wire v_5630;
wire v_5631;
wire v_5632;
wire v_5633;
wire v_5634;
wire v_5635;
wire v_5636;
wire v_5637;
wire v_5638;
wire v_5639;
wire v_5640;
wire v_5641;
wire v_5642;
wire v_5643;
wire v_5644;
wire v_5645;
wire v_5646;
wire v_5647;
wire v_5648;
wire v_5649;
wire v_5650;
wire v_5651;
wire v_5652;
wire v_5653;
wire v_5654;
wire v_5655;
wire v_5656;
wire v_5657;
wire v_5658;
wire v_5659;
wire v_5660;
wire v_5661;
wire v_5662;
wire v_5663;
wire v_5664;
wire v_5665;
wire v_5666;
wire v_5667;
wire v_5668;
wire v_5669;
wire v_5670;
wire v_5671;
wire v_5672;
wire v_5673;
wire v_5675;
wire v_5676;
wire v_5677;
wire v_5678;
wire v_5679;
wire v_5680;
wire v_5681;
wire v_5682;
wire v_5683;
wire v_5684;
wire v_5685;
wire v_5686;
wire v_5687;
wire v_5688;
wire v_5689;
wire v_5690;
wire v_5691;
wire v_5692;
wire v_5693;
wire v_5694;
wire v_5695;
wire v_5696;
wire v_5697;
wire v_5698;
wire v_5699;
wire v_5700;
wire v_5701;
wire v_5702;
wire v_5703;
wire v_5704;
wire v_5705;
wire v_5706;
wire v_5707;
wire v_5708;
wire v_5709;
wire v_5710;
wire v_5711;
wire v_5712;
wire v_5713;
wire v_5714;
wire v_5715;
wire v_5716;
wire v_5717;
wire v_5718;
wire v_5719;
wire v_5720;
wire v_5721;
wire v_5722;
wire v_5723;
wire v_5724;
wire v_5725;
wire v_5726;
wire v_5727;
wire v_5728;
wire v_5729;
wire v_5730;
wire v_5731;
wire v_5732;
wire v_5733;
wire v_5734;
wire v_5735;
wire v_5736;
wire v_5737;
wire v_5738;
wire v_5739;
wire v_5740;
wire v_5741;
wire v_5742;
wire v_5743;
wire v_5744;
wire v_5745;
wire v_5746;
wire v_5747;
wire v_5748;
wire v_5749;
wire v_5750;
wire v_5751;
wire v_5752;
wire v_5753;
wire v_5754;
wire v_5755;
wire v_5756;
wire v_5757;
wire v_5758;
wire v_5759;
wire v_5760;
wire v_5761;
wire v_5762;
wire v_5763;
wire v_5764;
wire v_5765;
wire v_5766;
wire v_5767;
wire v_5768;
wire v_5769;
wire v_5770;
wire v_5771;
wire v_5772;
wire v_5773;
wire v_5774;
wire v_5775;
wire v_5776;
wire v_5777;
wire v_5778;
wire v_5779;
wire v_5780;
wire v_5781;
wire v_5782;
wire v_5783;
wire v_5784;
wire v_5785;
wire v_5786;
wire v_5787;
wire v_5788;
wire v_5789;
wire v_5790;
wire v_5791;
wire v_5792;
wire v_5793;
wire v_5794;
wire v_5795;
wire v_5796;
wire v_5797;
wire v_5798;
wire v_5799;
wire v_5800;
wire v_5801;
wire v_5802;
wire v_5803;
wire v_5804;
wire v_5805;
wire v_5806;
wire v_5807;
wire v_5808;
wire v_5809;
wire v_5810;
wire v_5811;
wire v_5812;
wire v_5813;
wire v_5814;
wire v_5815;
wire v_5816;
wire v_5817;
wire v_5818;
wire v_5819;
wire v_5820;
wire v_5821;
wire v_5822;
wire v_5823;
wire v_5824;
wire v_5825;
wire v_5826;
wire v_5827;
wire v_5828;
wire v_5829;
wire v_5830;
wire v_5831;
wire v_5832;
wire v_5833;
wire v_5834;
wire v_5835;
wire v_5836;
wire v_5837;
wire v_5838;
wire v_5839;
wire v_5840;
wire v_5841;
wire v_5842;
wire v_5843;
wire v_5844;
wire v_5845;
wire v_5846;
wire v_5847;
wire v_5848;
wire v_5849;
wire v_5850;
wire v_5851;
wire v_5852;
wire v_5853;
wire v_5854;
wire v_5855;
wire v_5856;
wire v_5857;
wire v_5858;
wire v_5859;
wire v_5860;
wire v_5861;
wire v_5862;
wire v_5863;
wire v_5864;
wire v_5865;
wire v_5866;
wire v_5867;
wire v_5868;
wire v_5869;
wire v_5870;
wire v_5871;
wire v_5872;
wire v_5873;
wire v_5874;
wire v_5875;
wire v_5876;
wire v_5877;
wire v_5878;
wire v_5879;
wire v_5880;
wire v_5881;
wire v_5882;
wire v_5883;
wire v_5884;
wire v_5885;
wire v_5886;
wire v_5887;
wire v_5888;
wire v_5889;
wire v_5890;
wire v_5891;
wire v_5892;
wire v_5893;
wire v_5894;
wire v_5895;
wire v_5896;
wire v_5897;
wire v_5898;
wire v_5899;
wire v_5900;
wire v_5901;
wire v_5902;
wire v_5903;
wire v_5904;
wire v_5905;
wire v_5906;
wire v_5907;
wire v_5908;
wire v_5909;
wire v_5910;
wire v_5911;
wire v_5912;
wire v_5913;
wire v_5914;
wire v_5915;
wire v_5916;
wire v_5918;
wire v_5919;
wire v_5920;
wire v_5921;
wire v_5922;
wire v_5923;
wire v_5924;
wire v_5925;
wire v_5926;
wire v_5927;
wire v_5928;
wire v_5929;
wire v_5930;
wire v_5931;
wire v_5932;
wire v_5933;
wire v_5934;
wire v_5935;
wire v_5936;
wire v_5937;
wire v_5938;
wire v_5939;
wire v_5940;
wire v_5941;
wire v_5942;
wire v_5943;
wire v_5944;
wire v_5945;
wire v_5946;
wire v_5947;
wire v_5948;
wire v_5949;
wire v_5950;
wire v_5951;
wire v_5952;
wire v_5953;
wire v_5954;
wire v_5955;
wire v_5956;
wire v_5957;
wire v_5958;
wire v_5959;
wire v_5960;
wire v_5961;
wire v_5962;
wire v_5963;
wire v_5964;
wire v_5965;
wire v_5966;
wire v_5967;
wire v_5968;
wire v_5969;
wire v_5970;
wire v_5971;
wire v_5972;
wire v_5973;
wire v_5974;
wire v_5975;
wire v_5976;
wire v_5977;
wire v_5978;
wire v_5979;
wire v_5980;
wire v_5981;
wire v_5982;
wire v_5983;
wire v_5984;
wire v_5985;
wire v_5986;
wire v_5987;
wire v_5988;
wire v_5989;
wire v_5990;
wire v_5991;
wire v_5992;
wire v_5993;
wire v_5994;
wire v_5995;
wire v_5996;
wire v_5997;
wire v_5998;
wire v_5999;
wire v_6000;
wire v_6001;
wire v_6002;
wire v_6003;
wire v_6004;
wire v_6005;
wire v_6006;
wire v_6007;
wire v_6008;
wire v_6009;
wire v_6010;
wire v_6011;
wire v_6012;
wire v_6013;
wire v_6014;
wire v_6015;
wire v_6016;
wire v_6017;
wire v_6018;
wire v_6019;
wire v_6020;
wire v_6021;
wire v_6022;
wire v_6023;
wire v_6024;
wire v_6025;
wire v_6026;
wire v_6027;
wire v_6028;
wire v_6029;
wire v_6030;
wire v_6031;
wire v_6032;
wire v_6033;
wire v_6034;
wire v_6035;
wire v_6036;
wire v_6037;
wire v_6038;
wire v_6039;
wire v_6040;
wire v_6041;
wire v_6042;
wire v_6043;
wire v_6044;
wire v_6045;
wire v_6046;
wire v_6047;
wire v_6048;
wire v_6049;
wire v_6050;
wire v_6051;
wire v_6052;
wire v_6053;
wire v_6054;
wire v_6055;
wire v_6056;
wire v_6057;
wire v_6058;
wire v_6059;
wire v_6060;
wire v_6061;
wire v_6062;
wire v_6063;
wire v_6064;
wire v_6065;
wire v_6066;
wire v_6067;
wire v_6068;
wire v_6069;
wire v_6070;
wire v_6071;
wire v_6072;
wire v_6073;
wire v_6074;
wire v_6075;
wire v_6076;
wire v_6077;
wire v_6078;
wire v_6079;
wire v_6080;
wire v_6081;
wire v_6082;
wire v_6083;
wire v_6084;
wire v_6085;
wire v_6086;
wire v_6087;
wire v_6088;
wire v_6089;
wire v_6090;
wire v_6091;
wire v_6092;
wire v_6093;
wire v_6094;
wire v_6095;
wire v_6096;
wire v_6097;
wire v_6098;
wire v_6099;
wire v_6100;
wire v_6101;
wire v_6102;
wire v_6103;
wire v_6104;
wire v_6105;
wire v_6106;
wire v_6107;
wire v_6108;
wire v_6109;
wire v_6110;
wire v_6111;
wire v_6112;
wire v_6113;
wire v_6114;
wire v_6115;
wire v_6116;
wire v_6117;
wire v_6118;
wire v_6119;
wire v_6120;
wire v_6121;
wire v_6122;
wire v_6123;
wire v_6124;
wire v_6125;
wire v_6126;
wire v_6127;
wire v_6128;
wire v_6129;
wire v_6130;
wire v_6131;
wire v_6132;
wire v_6133;
wire v_6134;
wire v_6135;
wire v_6136;
wire v_6137;
wire v_6138;
wire v_6139;
wire v_6140;
wire v_6141;
wire v_6142;
wire v_6143;
wire v_6144;
wire v_6145;
wire v_6146;
wire v_6147;
wire v_6148;
wire v_6149;
wire v_6150;
wire v_6151;
wire v_6152;
wire v_6153;
wire v_6154;
wire v_6155;
wire v_6156;
wire v_6157;
wire v_6158;
wire v_6159;
wire v_6161;
wire v_6162;
wire v_6163;
wire v_6164;
wire v_6165;
wire v_6166;
wire v_6167;
wire v_6168;
wire v_6169;
wire v_6170;
wire v_6171;
wire v_6172;
wire v_6173;
wire v_6174;
wire v_6175;
wire v_6176;
wire v_6177;
wire v_6178;
wire v_6179;
wire v_6180;
wire v_6181;
wire v_6182;
wire v_6183;
wire v_6184;
wire v_6185;
wire v_6186;
wire v_6187;
wire v_6188;
wire v_6189;
wire v_6190;
wire v_6191;
wire v_6192;
wire v_6193;
wire v_6194;
wire v_6195;
wire v_6196;
wire v_6197;
wire v_6198;
wire v_6199;
wire v_6200;
wire v_6201;
wire v_6202;
wire v_6203;
wire v_6204;
wire v_6205;
wire v_6206;
wire v_6207;
wire v_6208;
wire v_6209;
wire v_6210;
wire v_6211;
wire v_6212;
wire v_6213;
wire v_6214;
wire v_6215;
wire v_6216;
wire v_6217;
wire v_6218;
wire v_6219;
wire v_6220;
wire v_6221;
wire v_6222;
wire v_6223;
wire v_6224;
wire v_6225;
wire v_6226;
wire v_6227;
wire v_6228;
wire v_6229;
wire v_6230;
wire v_6231;
wire v_6232;
wire v_6233;
wire v_6234;
wire v_6235;
wire v_6236;
wire v_6237;
wire v_6238;
wire v_6239;
wire v_6240;
wire v_6241;
wire v_6242;
wire v_6243;
wire v_6244;
wire v_6245;
wire v_6246;
wire v_6247;
wire v_6248;
wire v_6249;
wire v_6250;
wire v_6251;
wire v_6252;
wire v_6253;
wire v_6254;
wire v_6255;
wire v_6256;
wire v_6257;
wire v_6258;
wire v_6259;
wire v_6260;
wire v_6261;
wire v_6262;
wire v_6263;
wire v_6264;
wire v_6265;
wire v_6266;
wire v_6267;
wire v_6268;
wire v_6269;
wire v_6270;
wire v_6271;
wire v_6272;
wire v_6273;
wire v_6274;
wire v_6275;
wire v_6276;
wire v_6277;
wire v_6278;
wire v_6279;
wire v_6280;
wire v_6281;
wire v_6282;
wire v_6283;
wire v_6284;
wire v_6285;
wire v_6286;
wire v_6287;
wire v_6288;
wire v_6289;
wire v_6290;
wire v_6291;
wire v_6292;
wire v_6293;
wire v_6294;
wire v_6295;
wire v_6296;
wire v_6297;
wire v_6298;
wire v_6299;
wire v_6300;
wire v_6301;
wire v_6302;
wire v_6303;
wire v_6304;
wire v_6305;
wire v_6306;
wire v_6307;
wire v_6308;
wire v_6309;
wire v_6310;
wire v_6311;
wire v_6312;
wire v_6313;
wire v_6314;
wire v_6315;
wire v_6316;
wire v_6317;
wire v_6318;
wire v_6319;
wire v_6320;
wire v_6321;
wire v_6322;
wire v_6323;
wire v_6324;
wire v_6325;
wire v_6326;
wire v_6327;
wire v_6328;
wire v_6329;
wire v_6330;
wire v_6331;
wire v_6332;
wire v_6333;
wire v_6334;
wire v_6335;
wire v_6336;
wire v_6337;
wire v_6338;
wire v_6339;
wire v_6340;
wire v_6341;
wire v_6342;
wire v_6343;
wire v_6344;
wire v_6345;
wire v_6346;
wire v_6347;
wire v_6348;
wire v_6349;
wire v_6350;
wire v_6351;
wire v_6352;
wire v_6353;
wire v_6354;
wire v_6355;
wire v_6356;
wire v_6357;
wire v_6358;
wire v_6359;
wire v_6360;
wire v_6361;
wire v_6362;
wire v_6363;
wire v_6364;
wire v_6365;
wire v_6366;
wire v_6367;
wire v_6368;
wire v_6369;
wire v_6370;
wire v_6371;
wire v_6372;
wire v_6373;
wire v_6374;
wire v_6375;
wire v_6376;
wire v_6377;
wire v_6378;
wire v_6379;
wire v_6380;
wire v_6381;
wire v_6382;
wire v_6383;
wire v_6384;
wire v_6385;
wire v_6386;
wire v_6387;
wire v_6388;
wire v_6389;
wire v_6390;
wire v_6391;
wire v_6392;
wire v_6393;
wire v_6394;
wire v_6395;
wire v_6396;
wire v_6397;
wire v_6398;
wire v_6399;
wire v_6400;
wire v_6401;
wire v_6402;
wire v_6404;
wire v_6405;
wire v_6406;
wire v_6407;
wire v_6408;
wire v_6409;
wire v_6410;
wire v_6411;
wire v_6412;
wire v_6413;
wire v_6414;
wire v_6415;
wire v_6416;
wire v_6417;
wire v_6418;
wire v_6419;
wire v_6420;
wire v_6421;
wire v_6422;
wire v_6423;
wire v_6424;
wire v_6425;
wire v_6426;
wire v_6427;
wire v_6428;
wire v_6429;
wire v_6430;
wire v_6431;
wire v_6432;
wire v_6433;
wire v_6434;
wire v_6435;
wire v_6436;
wire v_6437;
wire v_6438;
wire v_6439;
wire v_6440;
wire v_6441;
wire v_6442;
wire v_6443;
wire v_6444;
wire v_6445;
wire v_6446;
wire v_6447;
wire v_6448;
wire v_6449;
wire v_6450;
wire v_6451;
wire v_6452;
wire v_6453;
wire v_6454;
wire v_6455;
wire v_6456;
wire v_6457;
wire v_6458;
wire v_6459;
wire v_6460;
wire v_6461;
wire v_6462;
wire v_6463;
wire v_6464;
wire v_6465;
wire v_6466;
wire v_6467;
wire v_6468;
wire v_6469;
wire v_6470;
wire v_6471;
wire v_6472;
wire v_6473;
wire v_6474;
wire v_6475;
wire v_6476;
wire v_6477;
wire v_6478;
wire v_6479;
wire v_6480;
wire v_6481;
wire v_6482;
wire v_6483;
wire v_6484;
wire v_6485;
wire v_6486;
wire v_6487;
wire v_6488;
wire v_6489;
wire v_6490;
wire v_6491;
wire v_6492;
wire v_6493;
wire v_6494;
wire v_6495;
wire v_6496;
wire v_6497;
wire v_6498;
wire v_6499;
wire v_6500;
wire v_6501;
wire v_6502;
wire v_6503;
wire v_6504;
wire v_6505;
wire v_6506;
wire v_6507;
wire v_6508;
wire v_6509;
wire v_6510;
wire v_6511;
wire v_6512;
wire v_6513;
wire v_6514;
wire v_6515;
wire v_6516;
wire v_6517;
wire v_6518;
wire v_6519;
wire v_6520;
wire v_6521;
wire v_6522;
wire v_6523;
wire v_6524;
wire v_6525;
wire v_6526;
wire v_6527;
wire v_6528;
wire v_6529;
wire v_6530;
wire v_6531;
wire v_6532;
wire v_6533;
wire v_6534;
wire v_6535;
wire v_6536;
wire v_6537;
wire v_6538;
wire v_6539;
wire v_6540;
wire v_6541;
wire v_6542;
wire v_6543;
wire v_6544;
wire v_6545;
wire v_6546;
wire v_6547;
wire v_6548;
wire v_6549;
wire v_6550;
wire v_6551;
wire v_6552;
wire v_6553;
wire v_6554;
wire v_6555;
wire v_6556;
wire v_6557;
wire v_6558;
wire v_6559;
wire v_6560;
wire v_6561;
wire v_6562;
wire v_6563;
wire v_6564;
wire v_6565;
wire v_6566;
wire v_6567;
wire v_6568;
wire v_6569;
wire v_6570;
wire v_6571;
wire v_6572;
wire v_6573;
wire v_6574;
wire v_6575;
wire v_6576;
wire v_6577;
wire v_6578;
wire v_6579;
wire v_6580;
wire v_6581;
wire v_6582;
wire v_6583;
wire v_6584;
wire v_6585;
wire v_6586;
wire v_6587;
wire v_6588;
wire v_6589;
wire v_6590;
wire v_6591;
wire v_6592;
wire v_6593;
wire v_6594;
wire v_6595;
wire v_6596;
wire v_6597;
wire v_6598;
wire v_6599;
wire v_6600;
wire v_6601;
wire v_6602;
wire v_6603;
wire v_6604;
wire v_6605;
wire v_6606;
wire v_6607;
wire v_6608;
wire v_6609;
wire v_6610;
wire v_6611;
wire v_6612;
wire v_6613;
wire v_6614;
wire v_6615;
wire v_6616;
wire v_6617;
wire v_6618;
wire v_6619;
wire v_6620;
wire v_6621;
wire v_6622;
wire v_6623;
wire v_6624;
wire v_6625;
wire v_6626;
wire v_6627;
wire v_6628;
wire v_6629;
wire v_6630;
wire v_6631;
wire v_6632;
wire v_6633;
wire v_6634;
wire v_6635;
wire v_6636;
wire v_6637;
wire v_6638;
wire v_6639;
wire v_6640;
wire v_6641;
wire v_6642;
wire v_6643;
wire v_6644;
wire v_6645;
wire v_6647;
wire v_6648;
wire v_6649;
wire v_6650;
wire v_6651;
wire v_6652;
wire v_6653;
wire v_6654;
wire v_6655;
wire v_6656;
wire v_6657;
wire v_6658;
wire v_6659;
wire v_6660;
wire v_6661;
wire v_6662;
wire v_6663;
wire v_6664;
wire v_6665;
wire v_6666;
wire v_6667;
wire v_6668;
wire v_6669;
wire v_6670;
wire v_6671;
wire v_6672;
wire v_6673;
wire v_6674;
wire v_6675;
wire v_6676;
wire v_6677;
wire v_6678;
wire v_6679;
wire v_6680;
wire v_6681;
wire v_6682;
wire v_6683;
wire v_6684;
wire v_6685;
wire v_6686;
wire v_6687;
wire v_6688;
wire v_6689;
wire v_6690;
wire v_6691;
wire v_6692;
wire v_6693;
wire v_6694;
wire v_6695;
wire v_6696;
wire v_6697;
wire v_6698;
wire v_6699;
wire v_6700;
wire v_6701;
wire v_6702;
wire v_6703;
wire v_6704;
wire v_6705;
wire v_6706;
wire v_6707;
wire v_6708;
wire v_6709;
wire v_6710;
wire v_6711;
wire v_6712;
wire v_6713;
wire v_6714;
wire v_6715;
wire v_6716;
wire v_6717;
wire v_6718;
wire v_6719;
wire v_6720;
wire v_6721;
wire v_6722;
wire v_6723;
wire v_6724;
wire v_6725;
wire v_6726;
wire v_6727;
wire v_6728;
wire v_6729;
wire v_6730;
wire v_6731;
wire v_6732;
wire v_6733;
wire v_6734;
wire v_6735;
wire v_6736;
wire v_6737;
wire v_6738;
wire v_6739;
wire v_6740;
wire v_6741;
wire v_6742;
wire v_6743;
wire v_6744;
wire v_6745;
wire v_6746;
wire v_6747;
wire v_6748;
wire v_6749;
wire v_6750;
wire v_6751;
wire v_6752;
wire v_6753;
wire v_6754;
wire v_6755;
wire v_6756;
wire v_6757;
wire v_6758;
wire v_6759;
wire v_6760;
wire v_6761;
wire v_6762;
wire v_6763;
wire v_6764;
wire v_6765;
wire v_6766;
wire v_6767;
wire v_6768;
wire v_6769;
wire v_6770;
wire v_6771;
wire v_6772;
wire v_6773;
wire v_6774;
wire v_6775;
wire v_6776;
wire v_6777;
wire v_6778;
wire v_6779;
wire v_6780;
wire v_6781;
wire v_6782;
wire v_6783;
wire v_6784;
wire v_6785;
wire v_6786;
wire v_6787;
wire v_6788;
wire v_6789;
wire v_6790;
wire v_6791;
wire v_6792;
wire v_6793;
wire v_6794;
wire v_6795;
wire v_6796;
wire v_6797;
wire v_6798;
wire v_6799;
wire v_6800;
wire v_6801;
wire v_6802;
wire v_6803;
wire v_6804;
wire v_6805;
wire v_6806;
wire v_6807;
wire v_6808;
wire v_6809;
wire v_6810;
wire v_6811;
wire v_6812;
wire v_6813;
wire v_6814;
wire v_6815;
wire v_6816;
wire v_6817;
wire v_6818;
wire v_6819;
wire v_6820;
wire v_6821;
wire v_6822;
wire v_6823;
wire v_6824;
wire v_6825;
wire v_6826;
wire v_6827;
wire v_6828;
wire v_6829;
wire v_6830;
wire v_6831;
wire v_6832;
wire v_6833;
wire v_6834;
wire v_6835;
wire v_6836;
wire v_6837;
wire v_6838;
wire v_6839;
wire v_6840;
wire v_6841;
wire v_6842;
wire v_6843;
wire v_6844;
wire v_6845;
wire v_6846;
wire v_6847;
wire v_6848;
wire v_6849;
wire v_6850;
wire v_6851;
wire v_6852;
wire v_6853;
wire v_6854;
wire v_6855;
wire v_6856;
wire v_6857;
wire v_6858;
wire v_6859;
wire v_6860;
wire v_6861;
wire v_6862;
wire v_6863;
wire v_6864;
wire v_6865;
wire v_6866;
wire v_6867;
wire v_6868;
wire v_6869;
wire v_6870;
wire v_6871;
wire v_6872;
wire v_6873;
wire v_6874;
wire v_6875;
wire v_6876;
wire v_6877;
wire v_6878;
wire v_6879;
wire v_6880;
wire v_6881;
wire v_6882;
wire v_6883;
wire v_6884;
wire v_6885;
wire v_6886;
wire v_6887;
wire v_6888;
wire v_6890;
wire v_6891;
wire v_6892;
wire v_6893;
wire v_6894;
wire v_6895;
wire v_6896;
wire v_6897;
wire v_6898;
wire v_6899;
wire v_6900;
wire v_6901;
wire v_6902;
wire v_6903;
wire v_6904;
wire v_6905;
wire v_6906;
wire v_6907;
wire v_6908;
wire v_6909;
wire v_6910;
wire v_6911;
wire v_6912;
wire v_6913;
wire v_6914;
wire v_6915;
wire v_6916;
wire v_6917;
wire v_6918;
wire v_6919;
wire v_6920;
wire v_6921;
wire v_6922;
wire v_6923;
wire v_6924;
wire v_6925;
wire v_6926;
wire v_6927;
wire v_6928;
wire v_6929;
wire v_6930;
wire v_6931;
wire v_6932;
wire v_6933;
wire v_6934;
wire v_6935;
wire v_6936;
wire v_6937;
wire v_6938;
wire v_6939;
wire v_6940;
wire v_6941;
wire v_6942;
wire v_6943;
wire v_6944;
wire v_6945;
wire v_6946;
wire v_6947;
wire v_6948;
wire v_6949;
wire v_6950;
wire v_6951;
wire v_6952;
wire v_6953;
wire v_6954;
wire v_6955;
wire v_6956;
wire v_6957;
wire v_6958;
wire v_6959;
wire v_6960;
wire v_6961;
wire v_6962;
wire v_6963;
wire v_6964;
wire v_6965;
wire v_6966;
wire v_6967;
wire v_6968;
wire v_6969;
wire v_6970;
wire v_6971;
wire v_6972;
wire v_6973;
wire v_6974;
wire v_6975;
wire v_6976;
wire v_6977;
wire v_6978;
wire v_6979;
wire v_6980;
wire v_6981;
wire v_6982;
wire v_6983;
wire v_6984;
wire v_6985;
wire v_6986;
wire v_6987;
wire v_6988;
wire v_6989;
wire v_6990;
wire v_6991;
wire v_6992;
wire v_6993;
wire v_6994;
wire v_6995;
wire v_6996;
wire v_6997;
wire v_6998;
wire v_6999;
wire v_7000;
wire v_7001;
wire v_7002;
wire v_7003;
wire v_7004;
wire v_7005;
wire v_7006;
wire v_7007;
wire v_7008;
wire v_7009;
wire v_7010;
wire v_7011;
wire v_7012;
wire v_7013;
wire v_7014;
wire v_7015;
wire v_7016;
wire v_7017;
wire v_7018;
wire v_7019;
wire v_7020;
wire v_7021;
wire v_7022;
wire v_7023;
wire v_7024;
wire v_7025;
wire v_7026;
wire v_7027;
wire v_7028;
wire v_7029;
wire v_7030;
wire v_7031;
wire v_7032;
wire v_7033;
wire v_7034;
wire v_7035;
wire v_7036;
wire v_7037;
wire v_7038;
wire v_7039;
wire v_7040;
wire v_7041;
wire v_7042;
wire v_7043;
wire v_7044;
wire v_7045;
wire v_7046;
wire v_7047;
wire v_7048;
wire v_7049;
wire v_7050;
wire v_7051;
wire v_7052;
wire v_7053;
wire v_7054;
wire v_7055;
wire v_7056;
wire v_7057;
wire v_7058;
wire v_7059;
wire v_7060;
wire v_7061;
wire v_7062;
wire v_7063;
wire v_7064;
wire v_7065;
wire v_7066;
wire v_7067;
wire v_7068;
wire v_7069;
wire v_7070;
wire v_7071;
wire v_7072;
wire v_7073;
wire v_7074;
wire v_7075;
wire v_7076;
wire v_7077;
wire v_7078;
wire v_7079;
wire v_7080;
wire v_7081;
wire v_7082;
wire v_7083;
wire v_7084;
wire v_7085;
wire v_7086;
wire v_7087;
wire v_7088;
wire v_7089;
wire v_7090;
wire v_7091;
wire v_7092;
wire v_7093;
wire v_7094;
wire v_7095;
wire v_7096;
wire v_7097;
wire v_7098;
wire v_7099;
wire v_7100;
wire v_7101;
wire v_7102;
wire v_7103;
wire v_7104;
wire v_7105;
wire v_7106;
wire v_7107;
wire v_7108;
wire v_7109;
wire v_7110;
wire v_7111;
wire v_7112;
wire v_7113;
wire v_7114;
wire v_7115;
wire v_7116;
wire v_7117;
wire v_7118;
wire v_7119;
wire v_7120;
wire v_7121;
wire v_7122;
wire v_7123;
wire v_7124;
wire v_7125;
wire v_7126;
wire v_7127;
wire v_7128;
wire v_7129;
wire v_7130;
wire v_7131;
wire v_7133;
wire v_7134;
wire v_7135;
wire v_7136;
wire v_7137;
wire v_7138;
wire v_7139;
wire v_7140;
wire v_7141;
wire v_7142;
wire v_7143;
wire v_7144;
wire v_7145;
wire v_7146;
wire v_7147;
wire v_7148;
wire v_7149;
wire v_7150;
wire v_7151;
wire v_7152;
wire v_7153;
wire v_7154;
wire v_7155;
wire v_7156;
wire v_7157;
wire v_7158;
wire v_7159;
wire v_7160;
wire v_7161;
wire v_7162;
wire v_7163;
wire v_7164;
wire v_7165;
wire v_7166;
wire v_7167;
wire v_7168;
wire v_7169;
wire v_7170;
wire v_7171;
wire v_7172;
wire v_7173;
wire v_7174;
wire v_7175;
wire v_7176;
wire v_7177;
wire v_7178;
wire v_7179;
wire v_7180;
wire v_7181;
wire v_7182;
wire v_7183;
wire v_7184;
wire v_7185;
wire v_7186;
wire v_7187;
wire v_7188;
wire v_7189;
wire v_7190;
wire v_7191;
wire v_7192;
wire v_7193;
wire v_7194;
wire v_7195;
wire v_7196;
wire v_7197;
wire v_7198;
wire v_7199;
wire v_7200;
wire v_7201;
wire v_7202;
wire v_7203;
wire v_7204;
wire v_7205;
wire v_7206;
wire v_7207;
wire v_7208;
wire v_7209;
wire v_7210;
wire v_7211;
wire v_7212;
wire v_7213;
wire v_7214;
wire v_7215;
wire v_7216;
wire v_7217;
wire v_7218;
wire v_7219;
wire v_7220;
wire v_7221;
wire v_7222;
wire v_7223;
wire v_7224;
wire v_7225;
wire v_7226;
wire v_7227;
wire v_7228;
wire v_7229;
wire v_7230;
wire v_7231;
wire v_7232;
wire v_7233;
wire v_7234;
wire v_7235;
wire v_7236;
wire v_7237;
wire v_7238;
wire v_7239;
wire v_7240;
wire v_7241;
wire v_7242;
wire v_7243;
wire v_7244;
wire v_7245;
wire v_7246;
wire v_7247;
wire v_7248;
wire v_7249;
wire v_7250;
wire v_7251;
wire v_7252;
wire v_7253;
wire v_7254;
wire v_7255;
wire v_7256;
wire v_7257;
wire v_7258;
wire v_7259;
wire v_7260;
wire v_7261;
wire v_7262;
wire v_7263;
wire v_7264;
wire v_7265;
wire v_7266;
wire v_7267;
wire v_7268;
wire v_7269;
wire v_7270;
wire v_7271;
wire v_7272;
wire v_7273;
wire v_7274;
wire v_7275;
wire v_7276;
wire v_7277;
wire v_7278;
wire v_7279;
wire v_7280;
wire v_7281;
wire v_7282;
wire v_7283;
wire v_7284;
wire v_7285;
wire v_7286;
wire v_7287;
wire v_7288;
wire v_7289;
wire v_7290;
wire v_7291;
wire v_7292;
wire v_7293;
wire v_7294;
wire v_7295;
wire v_7296;
wire v_7297;
wire v_7298;
wire v_7299;
wire v_7300;
wire v_7301;
wire v_7302;
wire v_7303;
wire v_7304;
wire v_7305;
wire v_7306;
wire v_7307;
wire v_7308;
wire v_7309;
wire v_7310;
wire v_7311;
wire v_7312;
wire v_7313;
wire v_7314;
wire v_7315;
wire v_7316;
wire v_7317;
wire v_7318;
wire v_7319;
wire v_7320;
wire v_7321;
wire v_7322;
wire v_7323;
wire v_7324;
wire v_7325;
wire v_7326;
wire v_7327;
wire v_7328;
wire v_7329;
wire v_7330;
wire v_7331;
wire v_7332;
wire v_7333;
wire v_7334;
wire v_7335;
wire v_7336;
wire v_7337;
wire v_7338;
wire v_7339;
wire v_7340;
wire v_7341;
wire v_7342;
wire v_7343;
wire v_7344;
wire v_7345;
wire v_7346;
wire v_7347;
wire v_7348;
wire v_7349;
wire v_7350;
wire v_7351;
wire v_7352;
wire v_7353;
wire v_7354;
wire v_7355;
wire v_7356;
wire v_7357;
wire v_7358;
wire v_7359;
wire v_7360;
wire v_7361;
wire v_7362;
wire v_7363;
wire v_7364;
wire v_7365;
wire v_7366;
wire v_7367;
wire v_7368;
wire v_7369;
wire v_7370;
wire v_7371;
wire v_7372;
wire v_7373;
wire v_7374;
wire v_7376;
wire v_7377;
wire v_7378;
wire v_7379;
wire v_7380;
wire v_7381;
wire v_7382;
wire v_7383;
wire v_7384;
wire v_7385;
wire v_7386;
wire v_7387;
wire v_7388;
wire v_7389;
wire v_7390;
wire v_7391;
wire v_7392;
wire v_7393;
wire v_7394;
wire v_7395;
wire v_7396;
wire v_7397;
wire v_7398;
wire v_7399;
wire v_7400;
wire v_7401;
wire v_7402;
wire v_7403;
wire v_7404;
wire v_7405;
wire v_7406;
wire v_7407;
wire v_7408;
wire v_7409;
wire v_7410;
wire v_7411;
wire v_7412;
wire v_7413;
wire v_7414;
wire v_7415;
wire v_7416;
wire v_7417;
wire v_7418;
wire v_7419;
wire v_7420;
wire v_7421;
wire v_7422;
wire v_7423;
wire v_7424;
wire v_7425;
wire v_7426;
wire v_7427;
wire v_7428;
wire v_7429;
wire v_7430;
wire v_7431;
wire v_7432;
wire v_7433;
wire v_7434;
wire v_7435;
wire v_7436;
wire v_7437;
wire v_7438;
wire v_7439;
wire v_7440;
wire v_7441;
wire v_7442;
wire v_7443;
wire v_7444;
wire v_7445;
wire v_7446;
wire v_7447;
wire v_7448;
wire v_7449;
wire v_7450;
wire v_7451;
wire v_7452;
wire v_7453;
wire v_7454;
wire v_7455;
wire v_7456;
wire v_7457;
wire v_7458;
wire v_7459;
wire v_7460;
wire v_7461;
wire v_7462;
wire v_7463;
wire v_7464;
wire v_7465;
wire v_7466;
wire v_7467;
wire v_7468;
wire v_7469;
wire v_7470;
wire v_7471;
wire v_7472;
wire v_7473;
wire v_7474;
wire v_7475;
wire v_7476;
wire v_7477;
wire v_7478;
wire v_7479;
wire v_7480;
wire v_7481;
wire v_7482;
wire v_7483;
wire v_7484;
wire v_7485;
wire v_7486;
wire v_7487;
wire v_7488;
wire v_7489;
wire v_7490;
wire v_7491;
wire v_7492;
wire v_7493;
wire v_7494;
wire v_7495;
wire v_7496;
wire v_7497;
wire v_7498;
wire v_7499;
wire v_7500;
wire v_7501;
wire v_7502;
wire v_7503;
wire v_7504;
wire v_7505;
wire v_7506;
wire v_7507;
wire v_7508;
wire v_7509;
wire v_7510;
wire v_7511;
wire v_7512;
wire v_7513;
wire v_7514;
wire v_7515;
wire v_7516;
wire v_7517;
wire v_7518;
wire v_7519;
wire v_7520;
wire v_7521;
wire v_7522;
wire v_7523;
wire v_7524;
wire v_7525;
wire v_7526;
wire v_7527;
wire v_7528;
wire v_7529;
wire v_7530;
wire v_7531;
wire v_7532;
wire v_7533;
wire v_7534;
wire v_7535;
wire v_7536;
wire v_7537;
wire v_7538;
wire v_7539;
wire v_7540;
wire v_7541;
wire v_7542;
wire v_7543;
wire v_7544;
wire v_7545;
wire v_7546;
wire v_7547;
wire v_7548;
wire v_7549;
wire v_7550;
wire v_7551;
wire v_7552;
wire v_7553;
wire v_7554;
wire v_7555;
wire v_7556;
wire v_7557;
wire v_7558;
wire v_7559;
wire v_7560;
wire v_7561;
wire v_7562;
wire v_7563;
wire v_7564;
wire v_7565;
wire v_7566;
wire v_7567;
wire v_7568;
wire v_7569;
wire v_7570;
wire v_7571;
wire v_7572;
wire v_7573;
wire v_7574;
wire v_7575;
wire v_7576;
wire v_7577;
wire v_7578;
wire v_7579;
wire v_7580;
wire v_7581;
wire v_7582;
wire v_7583;
wire v_7584;
wire v_7585;
wire v_7586;
wire v_7587;
wire v_7588;
wire v_7589;
wire v_7590;
wire v_7591;
wire v_7592;
wire v_7593;
wire v_7594;
wire v_7595;
wire v_7596;
wire v_7597;
wire v_7598;
wire v_7599;
wire v_7600;
wire v_7601;
wire v_7602;
wire v_7603;
wire v_7604;
wire v_7605;
wire v_7606;
wire v_7607;
wire v_7608;
wire v_7609;
wire v_7610;
wire v_7611;
wire v_7612;
wire v_7613;
wire v_7614;
wire v_7615;
wire v_7616;
wire v_7617;
wire v_7619;
wire v_7620;
wire v_7621;
wire v_7622;
wire v_7623;
wire v_7624;
wire v_7625;
wire v_7626;
wire v_7627;
wire v_7628;
wire v_7629;
wire v_7630;
wire v_7631;
wire v_7632;
wire v_7633;
wire v_7634;
wire v_7635;
wire v_7636;
wire v_7637;
wire v_7638;
wire v_7639;
wire v_7640;
wire v_7641;
wire v_7642;
wire v_7643;
wire v_7644;
wire v_7645;
wire v_7646;
wire v_7647;
wire v_7648;
wire v_7649;
wire v_7650;
wire v_7651;
wire v_7652;
wire v_7653;
wire v_7654;
wire v_7655;
wire v_7656;
wire v_7657;
wire v_7658;
wire v_7659;
wire v_7660;
wire v_7661;
wire v_7662;
wire v_7663;
wire v_7664;
wire v_7665;
wire v_7666;
wire v_7667;
wire v_7668;
wire v_7669;
wire v_7670;
wire v_7671;
wire v_7672;
wire v_7673;
wire v_7674;
wire v_7675;
wire v_7676;
wire v_7677;
wire v_7678;
wire v_7679;
wire v_7680;
wire v_7681;
wire v_7682;
wire v_7683;
wire v_7684;
wire v_7685;
wire v_7686;
wire v_7687;
wire v_7688;
wire v_7689;
wire v_7690;
wire v_7691;
wire v_7692;
wire v_7693;
wire v_7694;
wire v_7695;
wire v_7696;
wire v_7697;
wire v_7698;
wire v_7699;
wire v_7700;
wire v_7701;
wire v_7702;
wire v_7703;
wire v_7704;
wire v_7705;
wire v_7706;
wire v_7707;
wire v_7708;
wire v_7709;
wire v_7710;
wire v_7711;
wire v_7712;
wire v_7713;
wire v_7714;
wire v_7715;
wire v_7716;
wire v_7717;
wire v_7718;
wire v_7719;
wire v_7720;
wire v_7721;
wire v_7722;
wire v_7723;
wire v_7724;
wire v_7725;
wire v_7726;
wire v_7727;
wire v_7728;
wire v_7729;
wire v_7730;
wire v_7731;
wire v_7732;
wire v_7733;
wire v_7734;
wire v_7735;
wire v_7736;
wire v_7737;
wire v_7738;
wire v_7739;
wire v_7740;
wire v_7741;
wire v_7742;
wire v_7743;
wire v_7744;
wire v_7745;
wire v_7746;
wire v_7747;
wire v_7748;
wire v_7749;
wire v_7750;
wire v_7751;
wire v_7752;
wire v_7753;
wire v_7754;
wire v_7755;
wire v_7756;
wire v_7757;
wire v_7758;
wire v_7759;
wire v_7760;
wire v_7761;
wire v_7762;
wire v_7763;
wire v_7764;
wire v_7765;
wire v_7766;
wire v_7767;
wire v_7768;
wire v_7769;
wire v_7770;
wire v_7771;
wire v_7772;
wire v_7773;
wire v_7774;
wire v_7775;
wire v_7776;
wire v_7777;
wire v_7778;
wire v_7779;
wire v_7780;
wire v_7781;
wire v_7782;
wire v_7783;
wire v_7784;
wire v_7785;
wire v_7786;
wire v_7787;
wire v_7788;
wire v_7789;
wire v_7790;
wire v_7791;
wire v_7792;
wire v_7793;
wire v_7794;
wire v_7795;
wire v_7796;
wire v_7797;
wire v_7798;
wire v_7799;
wire v_7800;
wire v_7801;
wire v_7802;
wire v_7803;
wire v_7804;
wire v_7805;
wire v_7806;
wire v_7807;
wire v_7808;
wire v_7809;
wire v_7810;
wire v_7811;
wire v_7812;
wire v_7813;
wire v_7814;
wire v_7815;
wire v_7816;
wire v_7817;
wire v_7818;
wire v_7819;
wire v_7820;
wire v_7821;
wire v_7822;
wire v_7823;
wire v_7824;
wire v_7825;
wire v_7826;
wire v_7827;
wire v_7828;
wire v_7829;
wire v_7830;
wire v_7831;
wire v_7832;
wire v_7833;
wire v_7834;
wire v_7835;
wire v_7836;
wire v_7837;
wire v_7838;
wire v_7839;
wire v_7840;
wire v_7841;
wire v_7842;
wire v_7843;
wire v_7844;
wire v_7845;
wire v_7846;
wire v_7847;
wire v_7848;
wire v_7849;
wire v_7850;
wire v_7851;
wire v_7852;
wire v_7853;
wire v_7854;
wire v_7855;
wire v_7856;
wire v_7857;
wire v_7858;
wire v_7859;
wire v_7860;
wire v_7862;
wire v_7863;
wire v_7864;
wire v_7865;
wire v_7866;
wire v_7867;
wire v_7868;
wire v_7869;
wire v_7870;
wire v_7871;
wire v_7872;
wire v_7873;
wire v_7874;
wire v_7875;
wire v_7876;
wire v_7877;
wire v_7878;
wire v_7879;
wire v_7880;
wire v_7881;
wire v_7882;
wire v_7883;
wire v_7884;
wire v_7885;
wire v_7886;
wire v_7887;
wire v_7888;
wire v_7889;
wire v_7890;
wire v_7891;
wire v_7892;
wire v_7893;
wire v_7894;
wire v_7895;
wire v_7896;
wire v_7897;
wire v_7898;
wire v_7899;
wire v_7900;
wire v_7901;
wire v_7902;
wire v_7903;
wire v_7904;
wire v_7905;
wire v_7906;
wire v_7907;
wire v_7908;
wire v_7909;
wire v_7910;
wire v_7911;
wire v_7912;
wire v_7913;
wire v_7914;
wire v_7915;
wire v_7916;
wire v_7917;
wire v_7918;
wire v_7919;
wire v_7920;
wire v_7921;
wire v_7922;
wire v_7923;
wire v_7924;
wire v_7925;
wire v_7926;
wire v_7927;
wire v_7928;
wire v_7929;
wire v_7930;
wire v_7931;
wire v_7932;
wire v_7933;
wire v_7934;
wire v_7935;
wire v_7936;
wire v_7937;
wire v_7938;
wire v_7939;
wire v_7940;
wire v_7941;
wire v_7942;
wire v_7943;
wire v_7944;
wire v_7945;
wire v_7946;
wire v_7947;
wire v_7948;
wire v_7949;
wire v_7950;
wire v_7951;
wire v_7952;
wire v_7953;
wire v_7954;
wire v_7955;
wire v_7956;
wire v_7957;
wire v_7958;
wire v_7959;
wire v_7960;
wire v_7961;
wire v_7962;
wire v_7963;
wire v_7964;
wire v_7965;
wire v_7966;
wire v_7967;
wire v_7968;
wire v_7969;
wire v_7970;
wire v_7971;
wire v_7972;
wire v_7973;
wire v_7974;
wire v_7975;
wire v_7976;
wire v_7977;
wire v_7978;
wire v_7979;
wire v_7980;
wire v_7981;
wire v_7982;
wire v_7983;
wire v_7984;
wire v_7985;
wire v_7986;
wire v_7987;
wire v_7988;
wire v_7989;
wire v_7990;
wire v_7991;
wire v_7992;
wire v_7993;
wire v_7994;
wire v_7995;
wire v_7996;
wire v_7997;
wire v_7998;
wire v_7999;
wire v_8000;
wire v_8001;
wire v_8002;
wire v_8003;
wire v_8004;
wire v_8005;
wire v_8006;
wire v_8007;
wire v_8008;
wire v_8009;
wire v_8010;
wire v_8011;
wire v_8012;
wire v_8013;
wire v_8014;
wire v_8015;
wire v_8016;
wire v_8017;
wire v_8018;
wire v_8019;
wire v_8020;
wire v_8021;
wire v_8022;
wire v_8023;
wire v_8024;
wire v_8025;
wire v_8026;
wire v_8027;
wire v_8028;
wire v_8029;
wire v_8030;
wire v_8031;
wire v_8032;
wire v_8033;
wire v_8034;
wire v_8035;
wire v_8036;
wire v_8037;
wire v_8038;
wire v_8039;
wire v_8040;
wire v_8041;
wire v_8042;
wire v_8043;
wire v_8044;
wire v_8045;
wire v_8046;
wire v_8047;
wire v_8048;
wire v_8049;
wire v_8050;
wire v_8051;
wire v_8052;
wire v_8053;
wire v_8054;
wire v_8055;
wire v_8056;
wire v_8057;
wire v_8058;
wire v_8059;
wire v_8060;
wire v_8061;
wire v_8062;
wire v_8063;
wire v_8064;
wire v_8065;
wire v_8066;
wire v_8067;
wire v_8068;
wire v_8069;
wire v_8070;
wire v_8071;
wire v_8072;
wire v_8073;
wire v_8074;
wire v_8075;
wire v_8076;
wire v_8077;
wire v_8078;
wire v_8079;
wire v_8080;
wire v_8081;
wire v_8082;
wire v_8083;
wire v_8084;
wire v_8085;
wire v_8086;
wire v_8087;
wire v_8088;
wire v_8089;
wire v_8090;
wire v_8091;
wire v_8092;
wire v_8093;
wire v_8094;
wire v_8095;
wire v_8096;
wire v_8097;
wire v_8098;
wire v_8099;
wire v_8100;
wire v_8101;
wire v_8102;
wire v_8103;
wire v_8105;
wire v_8106;
wire v_8107;
wire v_8108;
wire v_8109;
wire v_8110;
wire v_8111;
wire v_8112;
wire v_8113;
wire v_8114;
wire v_8115;
wire v_8116;
wire v_8117;
wire v_8118;
wire v_8119;
wire v_8120;
wire v_8121;
wire v_8122;
wire v_8123;
wire v_8124;
wire v_8125;
wire v_8126;
wire v_8127;
wire v_8128;
wire v_8129;
wire v_8130;
wire v_8131;
wire v_8132;
wire v_8133;
wire v_8134;
wire v_8135;
wire v_8136;
wire v_8137;
wire v_8138;
wire v_8139;
wire v_8140;
wire v_8141;
wire v_8142;
wire v_8143;
wire v_8144;
wire v_8145;
wire v_8146;
wire v_8147;
wire v_8148;
wire v_8149;
wire v_8150;
wire v_8151;
wire v_8152;
wire v_8153;
wire v_8154;
wire v_8155;
wire v_8156;
wire v_8157;
wire v_8158;
wire v_8159;
wire v_8160;
wire v_8161;
wire v_8162;
wire v_8163;
wire v_8164;
wire v_8165;
wire v_8166;
wire v_8167;
wire v_8168;
wire v_8169;
wire v_8170;
wire v_8171;
wire v_8172;
wire v_8173;
wire v_8174;
wire v_8175;
wire v_8176;
wire v_8177;
wire v_8178;
wire v_8179;
wire v_8180;
wire v_8181;
wire v_8182;
wire v_8183;
wire v_8184;
wire v_8185;
wire v_8186;
wire v_8187;
wire v_8188;
wire v_8189;
wire v_8190;
wire v_8191;
wire v_8192;
wire v_8193;
wire v_8194;
wire v_8195;
wire v_8196;
wire v_8197;
wire v_8198;
wire v_8199;
wire v_8200;
wire v_8201;
wire v_8202;
wire v_8203;
wire v_8204;
wire v_8205;
wire v_8206;
wire v_8207;
wire v_8208;
wire v_8209;
wire v_8210;
wire v_8211;
wire v_8212;
wire v_8213;
wire v_8214;
wire v_8215;
wire v_8216;
wire v_8217;
wire v_8218;
wire v_8219;
wire v_8220;
wire v_8221;
wire v_8222;
wire v_8223;
wire v_8224;
wire v_8225;
wire v_8226;
wire v_8227;
wire v_8228;
wire v_8229;
wire v_8230;
wire v_8231;
wire v_8232;
wire v_8233;
wire v_8234;
wire v_8235;
wire v_8236;
wire v_8237;
wire v_8238;
wire v_8239;
wire v_8240;
wire v_8241;
wire v_8242;
wire v_8243;
wire v_8244;
wire v_8245;
wire v_8246;
wire v_8247;
wire v_8248;
wire v_8249;
wire v_8250;
wire v_8251;
wire v_8252;
wire v_8253;
wire v_8254;
wire v_8255;
wire v_8256;
wire v_8257;
wire v_8258;
wire v_8259;
wire v_8260;
wire v_8261;
wire v_8262;
wire v_8263;
wire v_8264;
wire v_8265;
wire v_8266;
wire v_8267;
wire v_8268;
wire v_8269;
wire v_8270;
wire v_8271;
wire v_8272;
wire v_8273;
wire v_8274;
wire v_8275;
wire v_8276;
wire v_8277;
wire v_8278;
wire v_8279;
wire v_8280;
wire v_8281;
wire v_8282;
wire v_8283;
wire v_8284;
wire v_8285;
wire v_8286;
wire v_8287;
wire v_8288;
wire v_8289;
wire v_8290;
wire v_8291;
wire v_8292;
wire v_8293;
wire v_8294;
wire v_8295;
wire v_8296;
wire v_8297;
wire v_8298;
wire v_8299;
wire v_8300;
wire v_8301;
wire v_8302;
wire v_8303;
wire v_8304;
wire v_8305;
wire v_8306;
wire v_8307;
wire v_8308;
wire v_8309;
wire v_8310;
wire v_8311;
wire v_8312;
wire v_8313;
wire v_8314;
wire v_8315;
wire v_8316;
wire v_8317;
wire v_8318;
wire v_8319;
wire v_8320;
wire v_8321;
wire v_8322;
wire v_8323;
wire v_8324;
wire v_8325;
wire v_8326;
wire v_8327;
wire v_8328;
wire v_8329;
wire v_8330;
wire v_8331;
wire v_8332;
wire v_8333;
wire v_8334;
wire v_8335;
wire v_8336;
wire v_8337;
wire v_8338;
wire v_8339;
wire v_8340;
wire v_8341;
wire v_8342;
wire v_8343;
wire v_8344;
wire v_8345;
wire v_8346;
wire v_8347;
wire v_8348;
wire v_8349;
wire v_8350;
wire v_8351;
wire v_8352;
wire v_8353;
wire v_8354;
wire v_8355;
wire v_8356;
wire v_8357;
wire v_8358;
wire v_8359;
wire v_8360;
wire v_8361;
wire v_8362;
wire v_8363;
wire v_8364;
wire v_8365;
wire v_8366;
wire v_8367;
wire v_8368;
wire v_8369;
wire v_8370;
wire v_8371;
wire v_8372;
wire v_8373;
wire v_8374;
wire v_8375;
wire v_8376;
wire v_8377;
wire v_8378;
wire v_8379;
wire v_8380;
wire v_8381;
wire v_8382;
wire v_8383;
wire v_8384;
wire v_8385;
wire v_8386;
wire v_8387;
wire v_8388;
wire v_8389;
wire v_8390;
wire v_8391;
wire v_8392;
wire v_8393;
wire v_8394;
wire v_8395;
wire v_8396;
wire v_8397;
wire v_8398;
wire v_8399;
wire v_8400;
wire v_8401;
wire v_8402;
wire v_8403;
wire v_8404;
wire v_8405;
wire v_8406;
wire v_8407;
wire v_8408;
wire v_8409;
wire v_8410;
wire v_8411;
wire v_8412;
wire v_8413;
wire v_8414;
wire v_8415;
wire v_8416;
wire v_8417;
wire v_8418;
wire v_8419;
wire v_8420;
wire v_8421;
wire v_8422;
wire v_8423;
wire v_8424;
wire v_8425;
wire v_8426;
wire v_8427;
wire v_8428;
wire v_8429;
wire v_8430;
wire v_8431;
wire v_8432;
wire v_8433;
wire v_8434;
wire v_8435;
wire v_8436;
wire v_8437;
wire v_8438;
wire v_8439;
wire v_8440;
wire v_8441;
wire v_8442;
wire v_8443;
wire v_8444;
wire v_8445;
wire v_8446;
wire v_8447;
wire v_8448;
wire v_8449;
wire v_8450;
wire v_8451;
wire v_8452;
wire v_8453;
wire v_8454;
wire v_8455;
wire v_8456;
wire v_8457;
wire v_8458;
wire v_8459;
wire v_8460;
wire v_8461;
wire v_8462;
wire v_8463;
wire v_8464;
wire v_8465;
wire v_8466;
wire v_8467;
wire v_8468;
wire v_8469;
wire v_8470;
wire v_8471;
wire v_8472;
wire v_8473;
wire v_8474;
wire v_8475;
wire v_8476;
wire v_8477;
wire v_8478;
wire v_8479;
wire v_8480;
wire v_8481;
wire v_8482;
wire v_8483;
wire v_8484;
wire v_8485;
wire v_8486;
wire v_8487;
wire v_8488;
wire v_8489;
wire v_8490;
wire v_8491;
wire v_8492;
wire v_8493;
wire v_8494;
wire v_8495;
wire v_8497;
wire v_8498;
wire v_8499;
wire v_8500;
wire v_8501;
wire v_8502;
wire v_8503;
wire v_8504;
wire v_8505;
wire v_8506;
wire v_8507;
wire v_8508;
wire v_8509;
wire v_8510;
wire v_8511;
wire v_8512;
wire v_8513;
wire v_8514;
wire v_8515;
wire v_8516;
wire v_8517;
wire v_8518;
wire v_8519;
wire v_8520;
wire v_8521;
wire v_8522;
wire v_8523;
wire v_8524;
wire v_8525;
wire v_8526;
wire v_8527;
wire v_8528;
wire v_8529;
wire v_8530;
wire v_8531;
wire v_8532;
wire v_8533;
wire v_8534;
wire v_8535;
wire v_8536;
wire v_8537;
wire v_8538;
wire v_8539;
wire v_8540;
wire v_8541;
wire v_8542;
wire v_8543;
wire v_8544;
wire v_8545;
wire v_8546;
wire v_8547;
wire v_8548;
wire v_8549;
wire v_8550;
wire v_8551;
wire v_8552;
wire v_8553;
wire v_8554;
wire v_8555;
wire v_8556;
wire v_8557;
wire v_8558;
wire v_8559;
wire v_8560;
wire v_8561;
wire v_8562;
wire v_8563;
wire v_8564;
wire v_8565;
wire v_8566;
wire v_8567;
wire v_8568;
wire v_8569;
wire v_8570;
wire v_8571;
wire v_8572;
wire v_8573;
wire v_8574;
wire v_8575;
wire v_8576;
wire v_8577;
wire v_8578;
wire v_8579;
wire v_8580;
wire v_8581;
wire v_8582;
wire v_8583;
wire v_8584;
wire v_8585;
wire v_8586;
wire v_8587;
wire v_8588;
wire v_8589;
wire v_8591;
wire v_8593;
wire v_8594;
wire v_8595;
wire v_8597;
wire v_8598;
wire v_8599;
wire v_8601;
wire v_8602;
wire v_8603;
wire v_8605;
wire v_8606;
wire v_8608;
wire v_8609;
wire v_8610;
wire v_8612;
wire v_8613;
wire v_8614;
wire v_8616;
wire v_8617;
wire v_8618;
wire v_8620;
wire v_8621;
wire v_8622;
wire v_8624;
wire v_8625;
wire v_8626;
wire v_8628;
wire v_8629;
wire v_8630;
wire v_8632;
wire v_8633;
wire v_8634;
wire v_8636;
wire v_8637;
wire v_8638;
wire v_8640;
wire v_8641;
wire v_8642;
wire v_8644;
wire v_8645;
wire v_8646;
wire v_8648;
wire v_8649;
wire v_8650;
wire v_8652;
wire v_8653;
wire v_8654;
wire v_8656;
wire v_8657;
wire v_8658;
wire v_8659;
wire v_8660;
wire v_8661;
wire v_8662;
wire v_8663;
wire v_8664;
wire v_8665;
wire v_8666;
wire v_8667;
wire v_8668;
wire v_8669;
wire v_8670;
wire v_8671;
wire v_8672;
wire v_8673;
wire v_8674;
wire v_8675;
wire v_8676;
wire v_8677;
wire v_8678;
wire v_8679;
wire v_8680;
wire v_8681;
wire v_8682;
wire v_8683;
wire v_8684;
wire v_8685;
wire v_8686;
wire v_8687;
wire v_8688;
wire v_8689;
wire v_8690;
wire v_8691;
wire v_8692;
wire v_8693;
wire v_8694;
wire v_8695;
wire v_8696;
wire v_8697;
wire v_8698;
wire v_8699;
wire v_8700;
wire v_8701;
wire v_8702;
wire v_8703;
wire v_8704;
wire v_8705;
wire v_8706;
wire v_8707;
wire v_8708;
wire v_8709;
wire v_8710;
wire v_8711;
wire v_8712;
wire v_8713;
wire v_8714;
wire v_8715;
wire v_8716;
wire v_8717;
wire v_8718;
wire v_8719;
wire v_8720;
wire v_8721;
wire v_8722;
wire v_8723;
wire v_8724;
wire v_8725;
wire v_8726;
wire v_8727;
wire v_8728;
wire v_8729;
wire v_8730;
wire v_8731;
wire v_8732;
wire v_8733;
wire v_8734;
wire v_8735;
wire v_8736;
wire v_8737;
wire v_8738;
wire v_8739;
wire v_8740;
wire v_8741;
wire v_8742;
wire v_8743;
wire v_8744;
wire v_8745;
wire v_8746;
wire v_8747;
wire v_8748;
wire v_8749;
wire v_8750;
wire v_8751;
wire v_8752;
wire v_8753;
wire v_8754;
wire v_8755;
wire v_8756;
wire v_8757;
wire v_8758;
wire v_8759;
wire v_8760;
wire v_8761;
wire v_8762;
wire v_8763;
wire v_8764;
wire v_8765;
wire v_8766;
wire v_8767;
wire v_8768;
wire v_8769;
wire v_8770;
wire v_8771;
wire v_8772;
wire v_8773;
wire v_8774;
wire v_8775;
wire v_8776;
wire v_8777;
wire v_8778;
wire v_8779;
wire v_8780;
wire v_8781;
wire v_8782;
wire v_8783;
wire v_8784;
wire v_8785;
wire v_8786;
wire v_8787;
wire v_8788;
wire v_8789;
wire v_8790;
wire v_8791;
wire v_8792;
wire v_8793;
wire v_8794;
wire v_8795;
wire v_8796;
wire v_8797;
wire v_8798;
wire v_8799;
wire v_8800;
wire v_8801;
wire v_8802;
wire v_8803;
wire v_8804;
wire v_8805;
wire v_8806;
wire v_8807;
wire v_8808;
wire v_8809;
wire v_8810;
wire v_8811;
wire v_8812;
wire v_8813;
wire v_8814;
wire v_8815;
wire v_8816;
wire v_8817;
wire v_8818;
wire v_8819;
wire v_8820;
wire v_8821;
wire v_8822;
wire v_8823;
wire v_8824;
wire v_8825;
wire v_8826;
wire v_8827;
wire v_8828;
wire v_8829;
wire v_8830;
wire v_8831;
wire v_8832;
wire v_8833;
wire v_8834;
wire v_8835;
wire v_8836;
wire v_8837;
wire v_8838;
wire v_8839;
wire v_8840;
wire v_8841;
wire v_8842;
wire v_8843;
wire v_8844;
wire v_8845;
wire v_8846;
wire v_8847;
wire v_8848;
wire v_8849;
wire v_8851;
wire v_8852;
wire v_8853;
wire v_8854;
wire v_8855;
wire v_8856;
wire v_8857;
wire v_8858;
wire v_8859;
wire v_8860;
wire v_8861;
wire v_8862;
wire v_8863;
wire v_8864;
wire v_8865;
wire v_8866;
wire v_8867;
wire v_8868;
wire v_8869;
wire v_8870;
wire v_8871;
wire v_8872;
wire v_8873;
wire v_8874;
wire v_8875;
wire v_8876;
wire v_8877;
wire v_8878;
wire v_8879;
wire v_8880;
wire v_8881;
wire v_8882;
wire v_8883;
wire v_8884;
wire v_8885;
wire v_8886;
wire v_8887;
wire v_8888;
wire v_8889;
wire v_8890;
wire v_8891;
wire v_8892;
wire v_8893;
wire v_8894;
wire v_8895;
wire v_8896;
wire v_8897;
wire v_8898;
wire v_8899;
wire v_8900;
wire v_8901;
wire v_8902;
wire v_8903;
wire v_8904;
wire v_8905;
wire v_8906;
wire v_8907;
wire v_8908;
wire v_8909;
wire v_8910;
wire v_8911;
wire v_8912;
wire v_8913;
wire v_8914;
wire v_8915;
wire v_8916;
wire v_8917;
wire v_8918;
wire v_8919;
wire v_8920;
wire v_8921;
wire v_8922;
wire v_8923;
wire v_8924;
wire v_8925;
wire v_8926;
wire v_8927;
wire v_8928;
wire v_8929;
wire v_8930;
wire v_8931;
wire v_8932;
wire v_8933;
wire v_8934;
wire v_8935;
wire v_8936;
wire v_8937;
wire v_8938;
wire v_8939;
wire v_8940;
wire v_8941;
wire v_8942;
wire v_8943;
wire v_8944;
wire v_8945;
wire v_8946;
wire v_8947;
wire v_8948;
wire v_8949;
wire v_8950;
wire v_8951;
wire v_8952;
wire v_8953;
wire v_8954;
wire v_8955;
wire v_8956;
wire v_8957;
wire v_8958;
wire v_8959;
wire v_8960;
wire v_8961;
wire v_8962;
wire v_8963;
wire v_8964;
wire v_8965;
wire v_8966;
wire v_8967;
wire v_8968;
wire v_8969;
wire v_8970;
wire v_8971;
wire v_8972;
wire v_8973;
wire v_8974;
wire v_8975;
wire v_8976;
wire v_8977;
wire v_8978;
wire v_8979;
wire v_8980;
wire v_8981;
wire v_8982;
wire v_8983;
wire v_8984;
wire v_8985;
wire v_8986;
wire v_8987;
wire v_8988;
wire v_8989;
wire v_8990;
wire v_8991;
wire v_8992;
wire v_8993;
wire v_8994;
wire v_8995;
wire v_8996;
wire v_8997;
wire v_8998;
wire v_8999;
wire v_9000;
wire v_9001;
wire v_9002;
wire v_9003;
wire v_9004;
wire v_9005;
wire v_9006;
wire v_9007;
wire v_9008;
wire v_9009;
wire v_9010;
wire v_9011;
wire v_9012;
wire v_9013;
wire v_9014;
wire v_9015;
wire v_9016;
wire v_9017;
wire v_9018;
wire v_9019;
wire v_9020;
wire v_9021;
wire v_9022;
wire v_9023;
wire v_9024;
wire v_9025;
wire v_9026;
wire v_9027;
wire v_9028;
wire v_9029;
wire v_9030;
wire v_9031;
wire v_9032;
wire v_9033;
wire v_9034;
wire v_9035;
wire v_9036;
wire v_9037;
wire v_9038;
wire v_9039;
wire v_9040;
wire v_9041;
wire v_9042;
wire v_9043;
wire v_9044;
wire v_9045;
wire v_9046;
wire v_9047;
wire v_9048;
wire v_9049;
wire v_9050;
wire v_9051;
wire v_9052;
wire v_9053;
wire v_9054;
wire v_9055;
wire v_9056;
wire v_9057;
wire v_9058;
wire v_9059;
wire v_9060;
wire v_9061;
wire v_9062;
wire v_9063;
wire v_9064;
wire v_9065;
wire v_9066;
wire v_9067;
wire v_9068;
wire v_9069;
wire v_9070;
wire v_9071;
wire v_9072;
wire v_9073;
wire v_9074;
wire v_9075;
wire v_9076;
wire v_9077;
wire v_9078;
wire v_9079;
wire v_9080;
wire v_9081;
wire v_9082;
wire v_9083;
wire v_9084;
wire v_9085;
wire v_9086;
wire v_9087;
wire v_9088;
wire v_9089;
wire v_9090;
wire v_9091;
wire v_9092;
wire v_9094;
wire v_9095;
wire v_9096;
wire v_9097;
wire v_9098;
wire v_9099;
wire v_9100;
wire v_9101;
wire v_9102;
wire v_9103;
wire v_9104;
wire v_9105;
wire v_9106;
wire v_9107;
wire v_9108;
wire v_9109;
wire v_9110;
wire v_9111;
wire v_9112;
wire v_9113;
wire v_9114;
wire v_9115;
wire v_9116;
wire v_9117;
wire v_9118;
wire v_9119;
wire v_9120;
wire v_9121;
wire v_9122;
wire v_9123;
wire v_9124;
wire v_9125;
wire v_9126;
wire v_9127;
wire v_9128;
wire v_9129;
wire v_9130;
wire v_9131;
wire v_9132;
wire v_9133;
wire v_9134;
wire v_9135;
wire v_9136;
wire v_9137;
wire v_9138;
wire v_9139;
wire v_9140;
wire v_9141;
wire v_9142;
wire v_9143;
wire v_9144;
wire v_9145;
wire v_9146;
wire v_9147;
wire v_9148;
wire v_9149;
wire v_9150;
wire v_9151;
wire v_9152;
wire v_9153;
wire v_9154;
wire v_9155;
wire v_9156;
wire v_9157;
wire v_9158;
wire v_9159;
wire v_9160;
wire v_9161;
wire v_9162;
wire v_9163;
wire v_9164;
wire v_9165;
wire v_9166;
wire v_9167;
wire v_9168;
wire v_9169;
wire v_9170;
wire v_9171;
wire v_9172;
wire v_9173;
wire v_9174;
wire v_9175;
wire v_9176;
wire v_9177;
wire v_9178;
wire v_9179;
wire v_9180;
wire v_9181;
wire v_9182;
wire v_9183;
wire v_9184;
wire v_9185;
wire v_9186;
wire v_9187;
wire v_9188;
wire v_9189;
wire v_9190;
wire v_9191;
wire v_9192;
wire v_9193;
wire v_9194;
wire v_9195;
wire v_9196;
wire v_9197;
wire v_9198;
wire v_9199;
wire v_9200;
wire v_9201;
wire v_9202;
wire v_9203;
wire v_9204;
wire v_9205;
wire v_9206;
wire v_9207;
wire v_9208;
wire v_9209;
wire v_9210;
wire v_9211;
wire v_9212;
wire v_9213;
wire v_9214;
wire v_9215;
wire v_9216;
wire v_9217;
wire v_9218;
wire v_9219;
wire v_9220;
wire v_9221;
wire v_9222;
wire v_9223;
wire v_9224;
wire v_9225;
wire v_9226;
wire v_9227;
wire v_9228;
wire v_9229;
wire v_9230;
wire v_9231;
wire v_9232;
wire v_9233;
wire v_9234;
wire v_9235;
wire v_9236;
wire v_9237;
wire v_9238;
wire v_9239;
wire v_9240;
wire v_9241;
wire v_9242;
wire v_9243;
wire v_9244;
wire v_9245;
wire v_9246;
wire v_9247;
wire v_9248;
wire v_9249;
wire v_9250;
wire v_9251;
wire v_9252;
wire v_9253;
wire v_9254;
wire v_9255;
wire v_9256;
wire v_9257;
wire v_9258;
wire v_9259;
wire v_9260;
wire v_9261;
wire v_9262;
wire v_9263;
wire v_9264;
wire v_9265;
wire v_9266;
wire v_9267;
wire v_9268;
wire v_9269;
wire v_9270;
wire v_9271;
wire v_9272;
wire v_9273;
wire v_9274;
wire v_9275;
wire v_9276;
wire v_9277;
wire v_9278;
wire v_9279;
wire v_9280;
wire v_9281;
wire v_9282;
wire v_9283;
wire v_9284;
wire v_9285;
wire v_9286;
wire v_9287;
wire v_9288;
wire v_9289;
wire v_9290;
wire v_9291;
wire v_9292;
wire v_9293;
wire v_9294;
wire v_9295;
wire v_9296;
wire v_9297;
wire v_9298;
wire v_9299;
wire v_9300;
wire v_9301;
wire v_9302;
wire v_9303;
wire v_9304;
wire v_9305;
wire v_9306;
wire v_9307;
wire v_9308;
wire v_9309;
wire v_9310;
wire v_9311;
wire v_9312;
wire v_9313;
wire v_9314;
wire v_9315;
wire v_9316;
wire v_9317;
wire v_9318;
wire v_9319;
wire v_9320;
wire v_9321;
wire v_9322;
wire v_9323;
wire v_9324;
wire v_9325;
wire v_9326;
wire v_9327;
wire v_9328;
wire v_9329;
wire v_9330;
wire v_9331;
wire v_9332;
wire v_9333;
wire v_9334;
wire v_9335;
wire v_9337;
wire v_9338;
wire v_9339;
wire v_9340;
wire v_9341;
wire v_9342;
wire v_9343;
wire v_9344;
wire v_9345;
wire v_9346;
wire v_9347;
wire v_9348;
wire v_9349;
wire v_9350;
wire v_9351;
wire v_9352;
wire v_9353;
wire v_9354;
wire v_9355;
wire v_9356;
wire v_9357;
wire v_9358;
wire v_9359;
wire v_9360;
wire v_9361;
wire v_9362;
wire v_9363;
wire v_9364;
wire v_9365;
wire v_9366;
wire v_9367;
wire v_9368;
wire v_9369;
wire v_9370;
wire v_9371;
wire v_9372;
wire v_9373;
wire v_9374;
wire v_9375;
wire v_9376;
wire v_9377;
wire v_9378;
wire v_9379;
wire v_9380;
wire v_9381;
wire v_9382;
wire v_9383;
wire v_9384;
wire v_9385;
wire v_9386;
wire v_9387;
wire v_9388;
wire v_9389;
wire v_9390;
wire v_9391;
wire v_9392;
wire v_9393;
wire v_9394;
wire v_9395;
wire v_9396;
wire v_9397;
wire v_9398;
wire v_9399;
wire v_9400;
wire v_9401;
wire v_9402;
wire v_9403;
wire v_9404;
wire v_9405;
wire v_9406;
wire v_9407;
wire v_9408;
wire v_9409;
wire v_9410;
wire v_9411;
wire v_9412;
wire v_9413;
wire v_9414;
wire v_9415;
wire v_9416;
wire v_9417;
wire v_9418;
wire v_9419;
wire v_9420;
wire v_9421;
wire v_9422;
wire v_9423;
wire v_9424;
wire v_9425;
wire v_9426;
wire v_9427;
wire v_9428;
wire v_9429;
wire v_9430;
wire v_9431;
wire v_9432;
wire v_9433;
wire v_9434;
wire v_9435;
wire v_9436;
wire v_9437;
wire v_9438;
wire v_9439;
wire v_9440;
wire v_9441;
wire v_9442;
wire v_9443;
wire v_9444;
wire v_9445;
wire v_9446;
wire v_9447;
wire v_9448;
wire v_9449;
wire v_9450;
wire v_9451;
wire v_9452;
wire v_9453;
wire v_9454;
wire v_9455;
wire v_9456;
wire v_9457;
wire v_9458;
wire v_9459;
wire v_9460;
wire v_9461;
wire v_9462;
wire v_9463;
wire v_9464;
wire v_9465;
wire v_9466;
wire v_9467;
wire v_9468;
wire v_9469;
wire v_9470;
wire v_9471;
wire v_9472;
wire v_9473;
wire v_9474;
wire v_9475;
wire v_9476;
wire v_9477;
wire v_9478;
wire v_9479;
wire v_9480;
wire v_9481;
wire v_9482;
wire v_9483;
wire v_9484;
wire v_9485;
wire v_9486;
wire v_9487;
wire v_9488;
wire v_9489;
wire v_9490;
wire v_9491;
wire v_9492;
wire v_9493;
wire v_9494;
wire v_9495;
wire v_9496;
wire v_9497;
wire v_9498;
wire v_9499;
wire v_9500;
wire v_9501;
wire v_9502;
wire v_9503;
wire v_9504;
wire v_9505;
wire v_9506;
wire v_9507;
wire v_9508;
wire v_9509;
wire v_9510;
wire v_9511;
wire v_9512;
wire v_9513;
wire v_9514;
wire v_9515;
wire v_9516;
wire v_9517;
wire v_9518;
wire v_9519;
wire v_9520;
wire v_9521;
wire v_9522;
wire v_9523;
wire v_9524;
wire v_9525;
wire v_9526;
wire v_9527;
wire v_9528;
wire v_9529;
wire v_9530;
wire v_9531;
wire v_9532;
wire v_9533;
wire v_9534;
wire v_9535;
wire v_9536;
wire v_9537;
wire v_9538;
wire v_9539;
wire v_9540;
wire v_9541;
wire v_9542;
wire v_9543;
wire v_9544;
wire v_9545;
wire v_9546;
wire v_9547;
wire v_9548;
wire v_9549;
wire v_9550;
wire v_9551;
wire v_9552;
wire v_9553;
wire v_9554;
wire v_9555;
wire v_9556;
wire v_9557;
wire v_9558;
wire v_9559;
wire v_9560;
wire v_9561;
wire v_9562;
wire v_9563;
wire v_9564;
wire v_9565;
wire v_9566;
wire v_9567;
wire v_9568;
wire v_9569;
wire v_9570;
wire v_9571;
wire v_9572;
wire v_9573;
wire v_9574;
wire v_9575;
wire v_9576;
wire v_9577;
wire v_9578;
wire v_9580;
wire v_9581;
wire v_9582;
wire v_9583;
wire v_9584;
wire v_9585;
wire v_9586;
wire v_9587;
wire v_9588;
wire v_9589;
wire v_9590;
wire v_9591;
wire v_9592;
wire v_9593;
wire v_9594;
wire v_9595;
wire v_9596;
wire v_9597;
wire v_9598;
wire v_9599;
wire v_9600;
wire v_9601;
wire v_9602;
wire v_9603;
wire v_9604;
wire v_9605;
wire v_9606;
wire v_9607;
wire v_9608;
wire v_9609;
wire v_9610;
wire v_9611;
wire v_9612;
wire v_9613;
wire v_9614;
wire v_9615;
wire v_9616;
wire v_9617;
wire v_9618;
wire v_9619;
wire v_9620;
wire v_9621;
wire v_9622;
wire v_9623;
wire v_9624;
wire v_9625;
wire v_9626;
wire v_9627;
wire v_9628;
wire v_9629;
wire v_9630;
wire v_9631;
wire v_9632;
wire v_9633;
wire v_9634;
wire v_9635;
wire v_9636;
wire v_9637;
wire v_9638;
wire v_9639;
wire v_9640;
wire v_9641;
wire v_9642;
wire v_9643;
wire v_9644;
wire v_9645;
wire v_9646;
wire v_9647;
wire v_9648;
wire v_9649;
wire v_9650;
wire v_9651;
wire v_9652;
wire v_9653;
wire v_9654;
wire v_9655;
wire v_9656;
wire v_9657;
wire v_9658;
wire v_9659;
wire v_9660;
wire v_9661;
wire v_9662;
wire v_9663;
wire v_9664;
wire v_9665;
wire v_9666;
wire v_9667;
wire v_9668;
wire v_9669;
wire v_9670;
wire v_9671;
wire v_9672;
wire v_9673;
wire v_9674;
wire v_9675;
wire v_9676;
wire v_9677;
wire v_9678;
wire v_9679;
wire v_9680;
wire v_9681;
wire v_9682;
wire v_9683;
wire v_9684;
wire v_9685;
wire v_9686;
wire v_9687;
wire v_9688;
wire v_9689;
wire v_9690;
wire v_9691;
wire v_9692;
wire v_9693;
wire v_9694;
wire v_9695;
wire v_9696;
wire v_9697;
wire v_9698;
wire v_9699;
wire v_9700;
wire v_9701;
wire v_9702;
wire v_9703;
wire v_9704;
wire v_9705;
wire v_9706;
wire v_9707;
wire v_9708;
wire v_9709;
wire v_9710;
wire v_9711;
wire v_9712;
wire v_9713;
wire v_9714;
wire v_9715;
wire v_9716;
wire v_9717;
wire v_9718;
wire v_9719;
wire v_9720;
wire v_9721;
wire v_9722;
wire v_9723;
wire v_9724;
wire v_9725;
wire v_9726;
wire v_9727;
wire v_9728;
wire v_9729;
wire v_9730;
wire v_9731;
wire v_9732;
wire v_9733;
wire v_9734;
wire v_9735;
wire v_9736;
wire v_9737;
wire v_9738;
wire v_9739;
wire v_9740;
wire v_9741;
wire v_9742;
wire v_9743;
wire v_9744;
wire v_9745;
wire v_9746;
wire v_9747;
wire v_9748;
wire v_9749;
wire v_9750;
wire v_9751;
wire v_9752;
wire v_9753;
wire v_9754;
wire v_9755;
wire v_9756;
wire v_9757;
wire v_9758;
wire v_9759;
wire v_9760;
wire v_9761;
wire v_9762;
wire v_9763;
wire v_9764;
wire v_9765;
wire v_9766;
wire v_9767;
wire v_9768;
wire v_9769;
wire v_9770;
wire v_9771;
wire v_9772;
wire v_9773;
wire v_9774;
wire v_9775;
wire v_9776;
wire v_9777;
wire v_9778;
wire v_9779;
wire v_9780;
wire v_9781;
wire v_9782;
wire v_9783;
wire v_9784;
wire v_9785;
wire v_9786;
wire v_9787;
wire v_9788;
wire v_9789;
wire v_9790;
wire v_9791;
wire v_9792;
wire v_9793;
wire v_9794;
wire v_9795;
wire v_9796;
wire v_9797;
wire v_9798;
wire v_9799;
wire v_9800;
wire v_9801;
wire v_9802;
wire v_9803;
wire v_9804;
wire v_9805;
wire v_9806;
wire v_9807;
wire v_9808;
wire v_9809;
wire v_9810;
wire v_9811;
wire v_9812;
wire v_9813;
wire v_9814;
wire v_9815;
wire v_9816;
wire v_9817;
wire v_9818;
wire v_9819;
wire v_9820;
wire v_9821;
wire v_9823;
wire v_9824;
wire v_9825;
wire v_9826;
wire v_9827;
wire v_9828;
wire v_9829;
wire v_9830;
wire v_9831;
wire v_9832;
wire v_9833;
wire v_9834;
wire v_9835;
wire v_9836;
wire v_9837;
wire v_9838;
wire v_9839;
wire v_9840;
wire v_9841;
wire v_9842;
wire v_9843;
wire v_9844;
wire v_9845;
wire v_9846;
wire v_9847;
wire v_9848;
wire v_9849;
wire v_9850;
wire v_9851;
wire v_9852;
wire v_9853;
wire v_9854;
wire v_9855;
wire v_9856;
wire v_9857;
wire v_9858;
wire v_9859;
wire v_9860;
wire v_9861;
wire v_9862;
wire v_9863;
wire v_9864;
wire v_9865;
wire v_9866;
wire v_9867;
wire v_9868;
wire v_9869;
wire v_9870;
wire v_9871;
wire v_9872;
wire v_9873;
wire v_9874;
wire v_9875;
wire v_9876;
wire v_9877;
wire v_9878;
wire v_9879;
wire v_9880;
wire v_9881;
wire v_9882;
wire v_9883;
wire v_9884;
wire v_9885;
wire v_9886;
wire v_9887;
wire v_9888;
wire v_9889;
wire v_9890;
wire v_9891;
wire v_9892;
wire v_9893;
wire v_9894;
wire v_9895;
wire v_9896;
wire v_9897;
wire v_9898;
wire v_9899;
wire v_9900;
wire v_9901;
wire v_9902;
wire v_9903;
wire v_9904;
wire v_9905;
wire v_9906;
wire v_9907;
wire v_9908;
wire v_9909;
wire v_9910;
wire v_9911;
wire v_9912;
wire v_9913;
wire v_9914;
wire v_9915;
wire v_9916;
wire v_9917;
wire v_9918;
wire v_9919;
wire v_9920;
wire v_9921;
wire v_9922;
wire v_9923;
wire v_9924;
wire v_9925;
wire v_9926;
wire v_9927;
wire v_9928;
wire v_9929;
wire v_9930;
wire v_9931;
wire v_9932;
wire v_9933;
wire v_9934;
wire v_9935;
wire v_9936;
wire v_9937;
wire v_9938;
wire v_9939;
wire v_9940;
wire v_9941;
wire v_9942;
wire v_9943;
wire v_9944;
wire v_9945;
wire v_9946;
wire v_9947;
wire v_9948;
wire v_9949;
wire v_9950;
wire v_9951;
wire v_9952;
wire v_9953;
wire v_9954;
wire v_9955;
wire v_9956;
wire v_9957;
wire v_9958;
wire v_9959;
wire v_9960;
wire v_9961;
wire v_9962;
wire v_9963;
wire v_9964;
wire v_9965;
wire v_9966;
wire v_9967;
wire v_9968;
wire v_9969;
wire v_9970;
wire v_9971;
wire v_9972;
wire v_9973;
wire v_9974;
wire v_9975;
wire v_9976;
wire v_9977;
wire v_9978;
wire v_9979;
wire v_9980;
wire v_9981;
wire v_9982;
wire v_9983;
wire v_9984;
wire v_9985;
wire v_9986;
wire v_9987;
wire v_9988;
wire v_9989;
wire v_9990;
wire v_9991;
wire v_9992;
wire v_9993;
wire v_9994;
wire v_9995;
wire v_9996;
wire v_9997;
wire v_9998;
wire v_9999;
wire v_10000;
wire v_10001;
wire v_10002;
wire v_10003;
wire v_10004;
wire v_10005;
wire v_10006;
wire v_10007;
wire v_10008;
wire v_10009;
wire v_10010;
wire v_10011;
wire v_10012;
wire v_10013;
wire v_10014;
wire v_10015;
wire v_10016;
wire v_10017;
wire v_10018;
wire v_10019;
wire v_10020;
wire v_10021;
wire v_10022;
wire v_10023;
wire v_10024;
wire v_10025;
wire v_10026;
wire v_10027;
wire v_10028;
wire v_10029;
wire v_10030;
wire v_10031;
wire v_10032;
wire v_10033;
wire v_10034;
wire v_10035;
wire v_10036;
wire v_10037;
wire v_10038;
wire v_10039;
wire v_10040;
wire v_10041;
wire v_10042;
wire v_10043;
wire v_10044;
wire v_10045;
wire v_10046;
wire v_10047;
wire v_10048;
wire v_10049;
wire v_10050;
wire v_10051;
wire v_10052;
wire v_10053;
wire v_10054;
wire v_10055;
wire v_10056;
wire v_10057;
wire v_10058;
wire v_10059;
wire v_10060;
wire v_10061;
wire v_10062;
wire v_10063;
wire v_10064;
wire v_10066;
wire v_10067;
wire v_10068;
wire v_10069;
wire v_10070;
wire v_10071;
wire v_10072;
wire v_10073;
wire v_10074;
wire v_10075;
wire v_10076;
wire v_10077;
wire v_10078;
wire v_10079;
wire v_10080;
wire v_10081;
wire v_10082;
wire v_10083;
wire v_10084;
wire v_10085;
wire v_10086;
wire v_10087;
wire v_10088;
wire v_10089;
wire v_10090;
wire v_10091;
wire v_10092;
wire v_10093;
wire v_10094;
wire v_10095;
wire v_10096;
wire v_10097;
wire v_10098;
wire v_10099;
wire v_10100;
wire v_10101;
wire v_10102;
wire v_10103;
wire v_10104;
wire v_10105;
wire v_10106;
wire v_10107;
wire v_10108;
wire v_10109;
wire v_10110;
wire v_10111;
wire v_10112;
wire v_10113;
wire v_10114;
wire v_10115;
wire v_10116;
wire v_10117;
wire v_10118;
wire v_10119;
wire v_10120;
wire v_10121;
wire v_10122;
wire v_10123;
wire v_10124;
wire v_10125;
wire v_10126;
wire v_10127;
wire v_10128;
wire v_10129;
wire v_10130;
wire v_10131;
wire v_10132;
wire v_10133;
wire v_10134;
wire v_10135;
wire v_10136;
wire v_10137;
wire v_10138;
wire v_10139;
wire v_10140;
wire v_10141;
wire v_10142;
wire v_10143;
wire v_10144;
wire v_10145;
wire v_10146;
wire v_10147;
wire v_10148;
wire v_10149;
wire v_10150;
wire v_10151;
wire v_10152;
wire v_10153;
wire v_10154;
wire v_10155;
wire v_10156;
wire v_10157;
wire v_10158;
wire v_10159;
wire v_10160;
wire v_10161;
wire v_10162;
wire v_10163;
wire v_10164;
wire v_10165;
wire v_10166;
wire v_10167;
wire v_10168;
wire v_10169;
wire v_10170;
wire v_10171;
wire v_10172;
wire v_10173;
wire v_10174;
wire v_10175;
wire v_10176;
wire v_10177;
wire v_10178;
wire v_10179;
wire v_10180;
wire v_10181;
wire v_10182;
wire v_10183;
wire v_10184;
wire v_10185;
wire v_10186;
wire v_10187;
wire v_10188;
wire v_10189;
wire v_10190;
wire v_10191;
wire v_10192;
wire v_10193;
wire v_10194;
wire v_10195;
wire v_10196;
wire v_10197;
wire v_10198;
wire v_10199;
wire v_10200;
wire v_10201;
wire v_10202;
wire v_10203;
wire v_10204;
wire v_10205;
wire v_10206;
wire v_10207;
wire v_10208;
wire v_10209;
wire v_10210;
wire v_10211;
wire v_10212;
wire v_10213;
wire v_10214;
wire v_10215;
wire v_10216;
wire v_10217;
wire v_10218;
wire v_10219;
wire v_10220;
wire v_10221;
wire v_10222;
wire v_10223;
wire v_10224;
wire v_10225;
wire v_10226;
wire v_10227;
wire v_10228;
wire v_10229;
wire v_10230;
wire v_10231;
wire v_10232;
wire v_10233;
wire v_10234;
wire v_10235;
wire v_10236;
wire v_10237;
wire v_10238;
wire v_10239;
wire v_10240;
wire v_10241;
wire v_10242;
wire v_10243;
wire v_10244;
wire v_10245;
wire v_10246;
wire v_10247;
wire v_10248;
wire v_10249;
wire v_10250;
wire v_10251;
wire v_10252;
wire v_10253;
wire v_10254;
wire v_10255;
wire v_10256;
wire v_10257;
wire v_10258;
wire v_10259;
wire v_10260;
wire v_10261;
wire v_10262;
wire v_10263;
wire v_10264;
wire v_10265;
wire v_10266;
wire v_10267;
wire v_10268;
wire v_10269;
wire v_10270;
wire v_10271;
wire v_10272;
wire v_10273;
wire v_10274;
wire v_10275;
wire v_10276;
wire v_10277;
wire v_10278;
wire v_10279;
wire v_10280;
wire v_10281;
wire v_10282;
wire v_10283;
wire v_10284;
wire v_10285;
wire v_10286;
wire v_10287;
wire v_10288;
wire v_10289;
wire v_10290;
wire v_10291;
wire v_10292;
wire v_10293;
wire v_10294;
wire v_10295;
wire v_10296;
wire v_10297;
wire v_10298;
wire v_10299;
wire v_10300;
wire v_10301;
wire v_10302;
wire v_10303;
wire v_10304;
wire v_10305;
wire v_10306;
wire v_10307;
wire v_10309;
wire v_10310;
wire v_10311;
wire v_10312;
wire v_10313;
wire v_10314;
wire v_10315;
wire v_10316;
wire v_10317;
wire v_10318;
wire v_10319;
wire v_10320;
wire v_10321;
wire v_10322;
wire v_10323;
wire v_10324;
wire v_10325;
wire v_10326;
wire v_10327;
wire v_10328;
wire v_10329;
wire v_10330;
wire v_10331;
wire v_10332;
wire v_10333;
wire v_10334;
wire v_10335;
wire v_10336;
wire v_10337;
wire v_10338;
wire v_10339;
wire v_10340;
wire v_10341;
wire v_10342;
wire v_10343;
wire v_10344;
wire v_10345;
wire v_10346;
wire v_10347;
wire v_10348;
wire v_10349;
wire v_10350;
wire v_10351;
wire v_10352;
wire v_10353;
wire v_10354;
wire v_10355;
wire v_10356;
wire v_10357;
wire v_10358;
wire v_10359;
wire v_10360;
wire v_10361;
wire v_10362;
wire v_10363;
wire v_10364;
wire v_10365;
wire v_10366;
wire v_10367;
wire v_10368;
wire v_10369;
wire v_10370;
wire v_10371;
wire v_10372;
wire v_10373;
wire v_10374;
wire v_10375;
wire v_10376;
wire v_10377;
wire v_10378;
wire v_10379;
wire v_10380;
wire v_10381;
wire v_10382;
wire v_10383;
wire v_10384;
wire v_10385;
wire v_10386;
wire v_10387;
wire v_10388;
wire v_10389;
wire v_10390;
wire v_10391;
wire v_10392;
wire v_10393;
wire v_10394;
wire v_10395;
wire v_10396;
wire v_10397;
wire v_10398;
wire v_10399;
wire v_10400;
wire v_10401;
wire v_10402;
wire v_10403;
wire v_10404;
wire v_10405;
wire v_10406;
wire v_10407;
wire v_10408;
wire v_10409;
wire v_10410;
wire v_10411;
wire v_10412;
wire v_10413;
wire v_10414;
wire v_10415;
wire v_10416;
wire v_10417;
wire v_10418;
wire v_10419;
wire v_10420;
wire v_10421;
wire v_10422;
wire v_10423;
wire v_10424;
wire v_10425;
wire v_10426;
wire v_10427;
wire v_10428;
wire v_10429;
wire v_10430;
wire v_10431;
wire v_10432;
wire v_10433;
wire v_10434;
wire v_10435;
wire v_10436;
wire v_10437;
wire v_10438;
wire v_10439;
wire v_10440;
wire v_10441;
wire v_10442;
wire v_10443;
wire v_10444;
wire v_10445;
wire v_10446;
wire v_10447;
wire v_10448;
wire v_10449;
wire v_10450;
wire v_10451;
wire v_10452;
wire v_10453;
wire v_10454;
wire v_10455;
wire v_10456;
wire v_10457;
wire v_10458;
wire v_10459;
wire v_10460;
wire v_10461;
wire v_10462;
wire v_10463;
wire v_10464;
wire v_10465;
wire v_10466;
wire v_10467;
wire v_10468;
wire v_10469;
wire v_10470;
wire v_10471;
wire v_10472;
wire v_10473;
wire v_10474;
wire v_10475;
wire v_10476;
wire v_10477;
wire v_10478;
wire v_10479;
wire v_10480;
wire v_10481;
wire v_10482;
wire v_10483;
wire v_10484;
wire v_10485;
wire v_10486;
wire v_10487;
wire v_10488;
wire v_10489;
wire v_10490;
wire v_10491;
wire v_10492;
wire v_10493;
wire v_10494;
wire v_10495;
wire v_10496;
wire v_10497;
wire v_10498;
wire v_10499;
wire v_10500;
wire v_10501;
wire v_10502;
wire v_10503;
wire v_10504;
wire v_10505;
wire v_10506;
wire v_10507;
wire v_10508;
wire v_10509;
wire v_10510;
wire v_10511;
wire v_10512;
wire v_10513;
wire v_10514;
wire v_10515;
wire v_10516;
wire v_10517;
wire v_10518;
wire v_10519;
wire v_10520;
wire v_10521;
wire v_10522;
wire v_10523;
wire v_10524;
wire v_10525;
wire v_10526;
wire v_10527;
wire v_10528;
wire v_10529;
wire v_10530;
wire v_10531;
wire v_10532;
wire v_10533;
wire v_10534;
wire v_10535;
wire v_10536;
wire v_10537;
wire v_10538;
wire v_10539;
wire v_10540;
wire v_10541;
wire v_10542;
wire v_10543;
wire v_10544;
wire v_10545;
wire v_10546;
wire v_10547;
wire v_10548;
wire v_10549;
wire v_10550;
wire v_10552;
wire v_10553;
wire v_10554;
wire v_10555;
wire v_10556;
wire v_10557;
wire v_10558;
wire v_10559;
wire v_10560;
wire v_10561;
wire v_10562;
wire v_10563;
wire v_10564;
wire v_10565;
wire v_10566;
wire v_10567;
wire v_10568;
wire v_10569;
wire v_10570;
wire v_10571;
wire v_10572;
wire v_10573;
wire v_10574;
wire v_10575;
wire v_10576;
wire v_10577;
wire v_10578;
wire v_10579;
wire v_10580;
wire v_10581;
wire v_10582;
wire v_10583;
wire v_10584;
wire v_10585;
wire v_10586;
wire v_10587;
wire v_10588;
wire v_10589;
wire v_10590;
wire v_10591;
wire v_10592;
wire v_10593;
wire v_10594;
wire v_10595;
wire v_10596;
wire v_10597;
wire v_10598;
wire v_10599;
wire v_10600;
wire v_10601;
wire v_10602;
wire v_10603;
wire v_10604;
wire v_10605;
wire v_10606;
wire v_10607;
wire v_10608;
wire v_10609;
wire v_10610;
wire v_10611;
wire v_10612;
wire v_10613;
wire v_10614;
wire v_10615;
wire v_10616;
wire v_10617;
wire v_10618;
wire v_10619;
wire v_10620;
wire v_10621;
wire v_10622;
wire v_10623;
wire v_10624;
wire v_10625;
wire v_10626;
wire v_10627;
wire v_10628;
wire v_10629;
wire v_10630;
wire v_10631;
wire v_10632;
wire v_10633;
wire v_10634;
wire v_10635;
wire v_10636;
wire v_10637;
wire v_10638;
wire v_10639;
wire v_10640;
wire v_10641;
wire v_10642;
wire v_10643;
wire v_10644;
wire v_10645;
wire v_10646;
wire v_10647;
wire v_10648;
wire v_10649;
wire v_10650;
wire v_10651;
wire v_10652;
wire v_10653;
wire v_10654;
wire v_10655;
wire v_10656;
wire v_10657;
wire v_10658;
wire v_10659;
wire v_10660;
wire v_10661;
wire v_10662;
wire v_10663;
wire v_10664;
wire v_10665;
wire v_10666;
wire v_10667;
wire v_10668;
wire v_10669;
wire v_10670;
wire v_10671;
wire v_10672;
wire v_10673;
wire v_10674;
wire v_10675;
wire v_10676;
wire v_10677;
wire v_10678;
wire v_10679;
wire v_10680;
wire v_10681;
wire v_10682;
wire v_10683;
wire v_10684;
wire v_10685;
wire v_10686;
wire v_10687;
wire v_10688;
wire v_10689;
wire v_10690;
wire v_10691;
wire v_10692;
wire v_10693;
wire v_10694;
wire v_10695;
wire v_10696;
wire v_10697;
wire v_10698;
wire v_10699;
wire v_10700;
wire v_10701;
wire v_10702;
wire v_10703;
wire v_10704;
wire v_10705;
wire v_10706;
wire v_10707;
wire v_10708;
wire v_10709;
wire v_10710;
wire v_10711;
wire v_10712;
wire v_10713;
wire v_10714;
wire v_10715;
wire v_10716;
wire v_10717;
wire v_10718;
wire v_10719;
wire v_10720;
wire v_10721;
wire v_10722;
wire v_10723;
wire v_10724;
wire v_10725;
wire v_10726;
wire v_10727;
wire v_10728;
wire v_10729;
wire v_10730;
wire v_10731;
wire v_10732;
wire v_10733;
wire v_10734;
wire v_10735;
wire v_10736;
wire v_10737;
wire v_10738;
wire v_10739;
wire v_10740;
wire v_10741;
wire v_10742;
wire v_10743;
wire v_10744;
wire v_10745;
wire v_10746;
wire v_10747;
wire v_10748;
wire v_10749;
wire v_10750;
wire v_10751;
wire v_10752;
wire v_10753;
wire v_10754;
wire v_10755;
wire v_10756;
wire v_10757;
wire v_10758;
wire v_10759;
wire v_10760;
wire v_10761;
wire v_10762;
wire v_10763;
wire v_10764;
wire v_10765;
wire v_10766;
wire v_10767;
wire v_10768;
wire v_10769;
wire v_10770;
wire v_10771;
wire v_10772;
wire v_10773;
wire v_10774;
wire v_10775;
wire v_10776;
wire v_10777;
wire v_10778;
wire v_10779;
wire v_10780;
wire v_10781;
wire v_10782;
wire v_10783;
wire v_10784;
wire v_10785;
wire v_10786;
wire v_10787;
wire v_10788;
wire v_10789;
wire v_10790;
wire v_10791;
wire v_10792;
wire v_10793;
wire v_10795;
wire v_10796;
wire v_10797;
wire v_10798;
wire v_10799;
wire v_10800;
wire v_10801;
wire v_10802;
wire v_10803;
wire v_10804;
wire v_10805;
wire v_10806;
wire v_10807;
wire v_10808;
wire v_10809;
wire v_10810;
wire v_10811;
wire v_10812;
wire v_10813;
wire v_10814;
wire v_10815;
wire v_10816;
wire v_10817;
wire v_10818;
wire v_10819;
wire v_10820;
wire v_10821;
wire v_10822;
wire v_10823;
wire v_10824;
wire v_10825;
wire v_10826;
wire v_10827;
wire v_10828;
wire v_10829;
wire v_10830;
wire v_10831;
wire v_10832;
wire v_10833;
wire v_10834;
wire v_10835;
wire v_10836;
wire v_10837;
wire v_10838;
wire v_10839;
wire v_10840;
wire v_10841;
wire v_10842;
wire v_10843;
wire v_10844;
wire v_10845;
wire v_10846;
wire v_10847;
wire v_10848;
wire v_10849;
wire v_10850;
wire v_10851;
wire v_10852;
wire v_10853;
wire v_10854;
wire v_10855;
wire v_10856;
wire v_10857;
wire v_10858;
wire v_10859;
wire v_10860;
wire v_10861;
wire v_10862;
wire v_10863;
wire v_10864;
wire v_10865;
wire v_10866;
wire v_10867;
wire v_10868;
wire v_10869;
wire v_10870;
wire v_10871;
wire v_10872;
wire v_10873;
wire v_10874;
wire v_10875;
wire v_10876;
wire v_10877;
wire v_10878;
wire v_10879;
wire v_10880;
wire v_10881;
wire v_10882;
wire v_10883;
wire v_10884;
wire v_10885;
wire v_10886;
wire v_10887;
wire v_10888;
wire v_10889;
wire v_10890;
wire v_10891;
wire v_10892;
wire v_10893;
wire v_10894;
wire v_10895;
wire v_10896;
wire v_10897;
wire v_10898;
wire v_10899;
wire v_10900;
wire v_10901;
wire v_10902;
wire v_10903;
wire v_10904;
wire v_10905;
wire v_10906;
wire v_10907;
wire v_10908;
wire v_10909;
wire v_10910;
wire v_10911;
wire v_10912;
wire v_10913;
wire v_10914;
wire v_10915;
wire v_10916;
wire v_10917;
wire v_10918;
wire v_10919;
wire v_10920;
wire v_10921;
wire v_10922;
wire v_10923;
wire v_10924;
wire v_10925;
wire v_10926;
wire v_10927;
wire v_10928;
wire v_10929;
wire v_10930;
wire v_10931;
wire v_10932;
wire v_10933;
wire v_10934;
wire v_10935;
wire v_10936;
wire v_10937;
wire v_10938;
wire v_10939;
wire v_10940;
wire v_10941;
wire v_10942;
wire v_10943;
wire v_10944;
wire v_10945;
wire v_10946;
wire v_10947;
wire v_10948;
wire v_10949;
wire v_10950;
wire v_10951;
wire v_10952;
wire v_10953;
wire v_10954;
wire v_10955;
wire v_10956;
wire v_10957;
wire v_10958;
wire v_10959;
wire v_10960;
wire v_10961;
wire v_10962;
wire v_10963;
wire v_10964;
wire v_10965;
wire v_10966;
wire v_10967;
wire v_10968;
wire v_10969;
wire v_10970;
wire v_10971;
wire v_10972;
wire v_10973;
wire v_10974;
wire v_10975;
wire v_10976;
wire v_10977;
wire v_10978;
wire v_10979;
wire v_10980;
wire v_10981;
wire v_10982;
wire v_10983;
wire v_10984;
wire v_10985;
wire v_10986;
wire v_10987;
wire v_10988;
wire v_10989;
wire v_10990;
wire v_10991;
wire v_10992;
wire v_10993;
wire v_10994;
wire v_10995;
wire v_10996;
wire v_10997;
wire v_10998;
wire v_10999;
wire v_11000;
wire v_11001;
wire v_11002;
wire v_11003;
wire v_11004;
wire v_11005;
wire v_11006;
wire v_11007;
wire v_11008;
wire v_11009;
wire v_11010;
wire v_11011;
wire v_11012;
wire v_11013;
wire v_11014;
wire v_11015;
wire v_11016;
wire v_11017;
wire v_11018;
wire v_11019;
wire v_11020;
wire v_11021;
wire v_11022;
wire v_11023;
wire v_11024;
wire v_11025;
wire v_11026;
wire v_11027;
wire v_11028;
wire v_11029;
wire v_11030;
wire v_11031;
wire v_11032;
wire v_11033;
wire v_11034;
wire v_11035;
wire v_11036;
wire v_11038;
wire v_11039;
wire v_11040;
wire v_11041;
wire v_11042;
wire v_11043;
wire v_11044;
wire v_11045;
wire v_11046;
wire v_11047;
wire v_11048;
wire v_11049;
wire v_11050;
wire v_11051;
wire v_11052;
wire v_11053;
wire v_11054;
wire v_11055;
wire v_11056;
wire v_11057;
wire v_11058;
wire v_11059;
wire v_11060;
wire v_11061;
wire v_11062;
wire v_11063;
wire v_11064;
wire v_11065;
wire v_11066;
wire v_11067;
wire v_11068;
wire v_11069;
wire v_11070;
wire v_11071;
wire v_11072;
wire v_11073;
wire v_11074;
wire v_11075;
wire v_11076;
wire v_11077;
wire v_11078;
wire v_11079;
wire v_11080;
wire v_11081;
wire v_11082;
wire v_11083;
wire v_11084;
wire v_11085;
wire v_11086;
wire v_11087;
wire v_11088;
wire v_11089;
wire v_11090;
wire v_11091;
wire v_11092;
wire v_11093;
wire v_11094;
wire v_11095;
wire v_11096;
wire v_11097;
wire v_11098;
wire v_11099;
wire v_11100;
wire v_11101;
wire v_11102;
wire v_11103;
wire v_11104;
wire v_11105;
wire v_11106;
wire v_11107;
wire v_11108;
wire v_11109;
wire v_11110;
wire v_11111;
wire v_11112;
wire v_11113;
wire v_11114;
wire v_11115;
wire v_11116;
wire v_11117;
wire v_11118;
wire v_11119;
wire v_11120;
wire v_11121;
wire v_11122;
wire v_11123;
wire v_11124;
wire v_11125;
wire v_11126;
wire v_11127;
wire v_11128;
wire v_11129;
wire v_11130;
wire v_11131;
wire v_11132;
wire v_11133;
wire v_11134;
wire v_11135;
wire v_11136;
wire v_11137;
wire v_11138;
wire v_11139;
wire v_11140;
wire v_11141;
wire v_11142;
wire v_11143;
wire v_11144;
wire v_11145;
wire v_11146;
wire v_11147;
wire v_11148;
wire v_11149;
wire v_11150;
wire v_11151;
wire v_11152;
wire v_11153;
wire v_11154;
wire v_11155;
wire v_11156;
wire v_11157;
wire v_11158;
wire v_11159;
wire v_11160;
wire v_11161;
wire v_11162;
wire v_11163;
wire v_11164;
wire v_11165;
wire v_11166;
wire v_11167;
wire v_11168;
wire v_11169;
wire v_11170;
wire v_11171;
wire v_11172;
wire v_11173;
wire v_11174;
wire v_11175;
wire v_11176;
wire v_11177;
wire v_11178;
wire v_11179;
wire v_11180;
wire v_11181;
wire v_11182;
wire v_11183;
wire v_11184;
wire v_11185;
wire v_11186;
wire v_11187;
wire v_11188;
wire v_11189;
wire v_11190;
wire v_11191;
wire v_11192;
wire v_11193;
wire v_11194;
wire v_11195;
wire v_11196;
wire v_11197;
wire v_11198;
wire v_11199;
wire v_11200;
wire v_11201;
wire v_11202;
wire v_11203;
wire v_11204;
wire v_11205;
wire v_11206;
wire v_11207;
wire v_11208;
wire v_11209;
wire v_11210;
wire v_11211;
wire v_11212;
wire v_11213;
wire v_11214;
wire v_11215;
wire v_11216;
wire v_11217;
wire v_11218;
wire v_11219;
wire v_11220;
wire v_11221;
wire v_11222;
wire v_11223;
wire v_11224;
wire v_11225;
wire v_11226;
wire v_11227;
wire v_11228;
wire v_11229;
wire v_11230;
wire v_11231;
wire v_11232;
wire v_11233;
wire v_11234;
wire v_11235;
wire v_11236;
wire v_11237;
wire v_11238;
wire v_11239;
wire v_11240;
wire v_11241;
wire v_11242;
wire v_11243;
wire v_11244;
wire v_11245;
wire v_11246;
wire v_11247;
wire v_11248;
wire v_11249;
wire v_11250;
wire v_11251;
wire v_11252;
wire v_11253;
wire v_11254;
wire v_11255;
wire v_11256;
wire v_11257;
wire v_11258;
wire v_11259;
wire v_11260;
wire v_11261;
wire v_11262;
wire v_11263;
wire v_11264;
wire v_11265;
wire v_11266;
wire v_11267;
wire v_11268;
wire v_11269;
wire v_11270;
wire v_11271;
wire v_11272;
wire v_11273;
wire v_11274;
wire v_11275;
wire v_11276;
wire v_11277;
wire v_11278;
wire v_11279;
wire v_11281;
wire v_11282;
wire v_11283;
wire v_11284;
wire v_11285;
wire v_11286;
wire v_11287;
wire v_11288;
wire v_11289;
wire v_11290;
wire v_11291;
wire v_11292;
wire v_11293;
wire v_11294;
wire v_11295;
wire v_11296;
wire v_11297;
wire v_11298;
wire v_11299;
wire v_11300;
wire v_11301;
wire v_11302;
wire v_11303;
wire v_11304;
wire v_11305;
wire v_11306;
wire v_11307;
wire v_11308;
wire v_11309;
wire v_11310;
wire v_11311;
wire v_11312;
wire v_11313;
wire v_11314;
wire v_11315;
wire v_11316;
wire v_11317;
wire v_11318;
wire v_11319;
wire v_11320;
wire v_11321;
wire v_11322;
wire v_11323;
wire v_11324;
wire v_11325;
wire v_11326;
wire v_11327;
wire v_11328;
wire v_11329;
wire v_11330;
wire v_11331;
wire v_11332;
wire v_11333;
wire v_11334;
wire v_11335;
wire v_11336;
wire v_11337;
wire v_11338;
wire v_11339;
wire v_11340;
wire v_11341;
wire v_11342;
wire v_11343;
wire v_11344;
wire v_11345;
wire v_11346;
wire v_11347;
wire v_11348;
wire v_11349;
wire v_11350;
wire v_11351;
wire v_11352;
wire v_11353;
wire v_11354;
wire v_11355;
wire v_11356;
wire v_11357;
wire v_11358;
wire v_11359;
wire v_11360;
wire v_11361;
wire v_11362;
wire v_11363;
wire v_11364;
wire v_11365;
wire v_11366;
wire v_11367;
wire v_11368;
wire v_11369;
wire v_11370;
wire v_11371;
wire v_11372;
wire v_11373;
wire v_11374;
wire v_11375;
wire v_11376;
wire v_11377;
wire v_11378;
wire v_11379;
wire v_11380;
wire v_11381;
wire v_11382;
wire v_11383;
wire v_11384;
wire v_11385;
wire v_11386;
wire v_11387;
wire v_11388;
wire v_11389;
wire v_11390;
wire v_11391;
wire v_11392;
wire v_11393;
wire v_11394;
wire v_11395;
wire v_11396;
wire v_11397;
wire v_11398;
wire v_11399;
wire v_11400;
wire v_11401;
wire v_11402;
wire v_11403;
wire v_11404;
wire v_11405;
wire v_11406;
wire v_11407;
wire v_11408;
wire v_11409;
wire v_11410;
wire v_11411;
wire v_11412;
wire v_11413;
wire v_11414;
wire v_11415;
wire v_11416;
wire v_11417;
wire v_11418;
wire v_11419;
wire v_11420;
wire v_11421;
wire v_11422;
wire v_11423;
wire v_11424;
wire v_11425;
wire v_11426;
wire v_11427;
wire v_11428;
wire v_11429;
wire v_11430;
wire v_11431;
wire v_11432;
wire v_11433;
wire v_11434;
wire v_11435;
wire v_11436;
wire v_11437;
wire v_11438;
wire v_11439;
wire v_11440;
wire v_11441;
wire v_11442;
wire v_11443;
wire v_11444;
wire v_11445;
wire v_11446;
wire v_11447;
wire v_11448;
wire v_11449;
wire v_11450;
wire v_11451;
wire v_11452;
wire v_11453;
wire v_11454;
wire v_11455;
wire v_11456;
wire v_11457;
wire v_11458;
wire v_11459;
wire v_11460;
wire v_11461;
wire v_11462;
wire v_11463;
wire v_11464;
wire v_11465;
wire v_11466;
wire v_11467;
wire v_11468;
wire v_11469;
wire v_11470;
wire v_11471;
wire v_11472;
wire v_11473;
wire v_11474;
wire v_11475;
wire v_11476;
wire v_11477;
wire v_11478;
wire v_11479;
wire v_11480;
wire v_11481;
wire v_11482;
wire v_11483;
wire v_11484;
wire v_11485;
wire v_11486;
wire v_11487;
wire v_11488;
wire v_11489;
wire v_11490;
wire v_11491;
wire v_11492;
wire v_11493;
wire v_11494;
wire v_11495;
wire v_11496;
wire v_11497;
wire v_11498;
wire v_11499;
wire v_11500;
wire v_11501;
wire v_11502;
wire v_11503;
wire v_11504;
wire v_11505;
wire v_11506;
wire v_11507;
wire v_11508;
wire v_11509;
wire v_11510;
wire v_11511;
wire v_11512;
wire v_11513;
wire v_11514;
wire v_11515;
wire v_11516;
wire v_11517;
wire v_11518;
wire v_11519;
wire v_11520;
wire v_11521;
wire v_11522;
wire v_11524;
wire v_11525;
wire v_11526;
wire v_11527;
wire v_11528;
wire v_11529;
wire v_11530;
wire v_11531;
wire v_11532;
wire v_11533;
wire v_11534;
wire v_11535;
wire v_11536;
wire v_11537;
wire v_11538;
wire v_11539;
wire v_11540;
wire v_11541;
wire v_11542;
wire v_11543;
wire v_11544;
wire v_11545;
wire v_11546;
wire v_11547;
wire v_11548;
wire v_11549;
wire v_11550;
wire v_11551;
wire v_11552;
wire v_11553;
wire v_11554;
wire v_11555;
wire v_11556;
wire v_11557;
wire v_11558;
wire v_11559;
wire v_11560;
wire v_11561;
wire v_11562;
wire v_11563;
wire v_11564;
wire v_11565;
wire v_11566;
wire v_11567;
wire v_11568;
wire v_11569;
wire v_11570;
wire v_11571;
wire v_11572;
wire v_11573;
wire v_11574;
wire v_11575;
wire v_11576;
wire v_11577;
wire v_11578;
wire v_11579;
wire v_11580;
wire v_11581;
wire v_11582;
wire v_11583;
wire v_11584;
wire v_11585;
wire v_11586;
wire v_11587;
wire v_11588;
wire v_11589;
wire v_11590;
wire v_11591;
wire v_11592;
wire v_11593;
wire v_11594;
wire v_11595;
wire v_11596;
wire v_11597;
wire v_11598;
wire v_11599;
wire v_11600;
wire v_11601;
wire v_11602;
wire v_11603;
wire v_11604;
wire v_11605;
wire v_11606;
wire v_11607;
wire v_11608;
wire v_11609;
wire v_11610;
wire v_11611;
wire v_11612;
wire v_11613;
wire v_11614;
wire v_11615;
wire v_11616;
wire v_11617;
wire v_11618;
wire v_11619;
wire v_11620;
wire v_11621;
wire v_11622;
wire v_11623;
wire v_11624;
wire v_11625;
wire v_11626;
wire v_11627;
wire v_11628;
wire v_11629;
wire v_11630;
wire v_11631;
wire v_11632;
wire v_11633;
wire v_11634;
wire v_11635;
wire v_11636;
wire v_11637;
wire v_11638;
wire v_11639;
wire v_11640;
wire v_11641;
wire v_11642;
wire v_11643;
wire v_11644;
wire v_11645;
wire v_11646;
wire v_11647;
wire v_11648;
wire v_11649;
wire v_11650;
wire v_11651;
wire v_11652;
wire v_11653;
wire v_11654;
wire v_11655;
wire v_11656;
wire v_11657;
wire v_11658;
wire v_11659;
wire v_11660;
wire v_11661;
wire v_11662;
wire v_11663;
wire v_11664;
wire v_11665;
wire v_11666;
wire v_11667;
wire v_11668;
wire v_11669;
wire v_11670;
wire v_11671;
wire v_11672;
wire v_11673;
wire v_11674;
wire v_11675;
wire v_11676;
wire v_11677;
wire v_11678;
wire v_11679;
wire v_11680;
wire v_11681;
wire v_11682;
wire v_11683;
wire v_11684;
wire v_11685;
wire v_11686;
wire v_11687;
wire v_11688;
wire v_11689;
wire v_11690;
wire v_11691;
wire v_11692;
wire v_11693;
wire v_11694;
wire v_11695;
wire v_11696;
wire v_11697;
wire v_11698;
wire v_11699;
wire v_11700;
wire v_11701;
wire v_11702;
wire v_11703;
wire v_11704;
wire v_11705;
wire v_11706;
wire v_11707;
wire v_11708;
wire v_11709;
wire v_11710;
wire v_11711;
wire v_11712;
wire v_11713;
wire v_11714;
wire v_11715;
wire v_11716;
wire v_11717;
wire v_11718;
wire v_11719;
wire v_11720;
wire v_11721;
wire v_11722;
wire v_11723;
wire v_11724;
wire v_11725;
wire v_11726;
wire v_11727;
wire v_11728;
wire v_11729;
wire v_11730;
wire v_11731;
wire v_11732;
wire v_11733;
wire v_11734;
wire v_11735;
wire v_11736;
wire v_11737;
wire v_11738;
wire v_11739;
wire v_11740;
wire v_11741;
wire v_11742;
wire v_11743;
wire v_11744;
wire v_11745;
wire v_11746;
wire v_11747;
wire v_11748;
wire v_11749;
wire v_11750;
wire v_11751;
wire v_11752;
wire v_11753;
wire v_11754;
wire v_11755;
wire v_11756;
wire v_11757;
wire v_11758;
wire v_11759;
wire v_11760;
wire v_11761;
wire v_11762;
wire v_11763;
wire v_11764;
wire v_11765;
wire v_11767;
wire v_11768;
wire v_11769;
wire v_11770;
wire v_11771;
wire v_11772;
wire v_11773;
wire v_11774;
wire v_11775;
wire v_11776;
wire v_11777;
wire v_11778;
wire v_11779;
wire v_11780;
wire v_11781;
wire v_11782;
wire v_11783;
wire v_11784;
wire v_11785;
wire v_11786;
wire v_11787;
wire v_11788;
wire v_11789;
wire v_11790;
wire v_11791;
wire v_11792;
wire v_11793;
wire v_11794;
wire v_11795;
wire v_11796;
wire v_11797;
wire v_11798;
wire v_11799;
wire v_11800;
wire v_11801;
wire v_11802;
wire v_11803;
wire v_11804;
wire v_11805;
wire v_11806;
wire v_11807;
wire v_11808;
wire v_11809;
wire v_11810;
wire v_11811;
wire v_11812;
wire v_11813;
wire v_11814;
wire v_11815;
wire v_11816;
wire v_11817;
wire v_11818;
wire v_11819;
wire v_11820;
wire v_11821;
wire v_11822;
wire v_11823;
wire v_11824;
wire v_11825;
wire v_11826;
wire v_11827;
wire v_11828;
wire v_11829;
wire v_11830;
wire v_11831;
wire v_11832;
wire v_11833;
wire v_11834;
wire v_11835;
wire v_11836;
wire v_11837;
wire v_11838;
wire v_11839;
wire v_11840;
wire v_11841;
wire v_11842;
wire v_11843;
wire v_11844;
wire v_11845;
wire v_11846;
wire v_11847;
wire v_11848;
wire v_11849;
wire v_11850;
wire v_11851;
wire v_11852;
wire v_11853;
wire v_11854;
wire v_11855;
wire v_11856;
wire v_11857;
wire v_11858;
wire v_11859;
wire v_11860;
wire v_11861;
wire v_11862;
wire v_11863;
wire v_11864;
wire v_11865;
wire v_11866;
wire v_11867;
wire v_11868;
wire v_11869;
wire v_11870;
wire v_11871;
wire v_11872;
wire v_11873;
wire v_11874;
wire v_11875;
wire v_11876;
wire v_11877;
wire v_11878;
wire v_11879;
wire v_11880;
wire v_11881;
wire v_11882;
wire v_11883;
wire v_11884;
wire v_11885;
wire v_11886;
wire v_11887;
wire v_11888;
wire v_11889;
wire v_11890;
wire v_11891;
wire v_11892;
wire v_11893;
wire v_11894;
wire v_11895;
wire v_11896;
wire v_11897;
wire v_11898;
wire v_11899;
wire v_11900;
wire v_11901;
wire v_11902;
wire v_11903;
wire v_11904;
wire v_11905;
wire v_11906;
wire v_11907;
wire v_11908;
wire v_11909;
wire v_11910;
wire v_11911;
wire v_11912;
wire v_11913;
wire v_11914;
wire v_11915;
wire v_11916;
wire v_11917;
wire v_11918;
wire v_11919;
wire v_11920;
wire v_11921;
wire v_11922;
wire v_11923;
wire v_11924;
wire v_11925;
wire v_11926;
wire v_11927;
wire v_11928;
wire v_11929;
wire v_11930;
wire v_11931;
wire v_11932;
wire v_11933;
wire v_11934;
wire v_11935;
wire v_11936;
wire v_11937;
wire v_11938;
wire v_11939;
wire v_11940;
wire v_11941;
wire v_11942;
wire v_11943;
wire v_11944;
wire v_11945;
wire v_11946;
wire v_11947;
wire v_11948;
wire v_11949;
wire v_11950;
wire v_11951;
wire v_11952;
wire v_11953;
wire v_11954;
wire v_11955;
wire v_11956;
wire v_11957;
wire v_11958;
wire v_11959;
wire v_11960;
wire v_11961;
wire v_11962;
wire v_11963;
wire v_11964;
wire v_11965;
wire v_11966;
wire v_11967;
wire v_11968;
wire v_11969;
wire v_11970;
wire v_11971;
wire v_11972;
wire v_11973;
wire v_11974;
wire v_11975;
wire v_11976;
wire v_11977;
wire v_11978;
wire v_11979;
wire v_11980;
wire v_11981;
wire v_11982;
wire v_11983;
wire v_11984;
wire v_11985;
wire v_11986;
wire v_11987;
wire v_11988;
wire v_11989;
wire v_11990;
wire v_11991;
wire v_11992;
wire v_11993;
wire v_11994;
wire v_11995;
wire v_11996;
wire v_11997;
wire v_11998;
wire v_11999;
wire v_12000;
wire v_12001;
wire v_12002;
wire v_12003;
wire v_12004;
wire v_12005;
wire v_12006;
wire v_12007;
wire v_12008;
wire v_12010;
wire v_12011;
wire v_12012;
wire v_12013;
wire v_12014;
wire v_12015;
wire v_12016;
wire v_12017;
wire v_12018;
wire v_12019;
wire v_12020;
wire v_12021;
wire v_12022;
wire v_12023;
wire v_12024;
wire v_12025;
wire v_12026;
wire v_12027;
wire v_12028;
wire v_12029;
wire v_12030;
wire v_12031;
wire v_12032;
wire v_12033;
wire v_12034;
wire v_12035;
wire v_12036;
wire v_12037;
wire v_12038;
wire v_12039;
wire v_12040;
wire v_12041;
wire v_12042;
wire v_12043;
wire v_12044;
wire v_12045;
wire v_12046;
wire v_12047;
wire v_12048;
wire v_12049;
wire v_12050;
wire v_12051;
wire v_12052;
wire v_12053;
wire v_12054;
wire v_12055;
wire v_12056;
wire v_12057;
wire v_12058;
wire v_12059;
wire v_12060;
wire v_12061;
wire v_12062;
wire v_12063;
wire v_12064;
wire v_12065;
wire v_12066;
wire v_12067;
wire v_12068;
wire v_12069;
wire v_12070;
wire v_12071;
wire v_12072;
wire v_12073;
wire v_12074;
wire v_12075;
wire v_12076;
wire v_12077;
wire v_12078;
wire v_12079;
wire v_12080;
wire v_12081;
wire v_12082;
wire v_12083;
wire v_12084;
wire v_12085;
wire v_12086;
wire v_12087;
wire v_12088;
wire v_12089;
wire v_12090;
wire v_12091;
wire v_12092;
wire v_12093;
wire v_12094;
wire v_12095;
wire v_12096;
wire v_12097;
wire v_12098;
wire v_12099;
wire v_12100;
wire v_12101;
wire v_12102;
wire v_12103;
wire v_12104;
wire v_12105;
wire v_12106;
wire v_12107;
wire v_12108;
wire v_12109;
wire v_12110;
wire v_12111;
wire v_12112;
wire v_12113;
wire v_12114;
wire v_12115;
wire v_12116;
wire v_12117;
wire v_12118;
wire v_12119;
wire v_12120;
wire v_12121;
wire v_12122;
wire v_12123;
wire v_12124;
wire v_12125;
wire v_12126;
wire v_12127;
wire v_12128;
wire v_12129;
wire v_12130;
wire v_12131;
wire v_12132;
wire v_12133;
wire v_12134;
wire v_12135;
wire v_12136;
wire v_12137;
wire v_12138;
wire v_12139;
wire v_12140;
wire v_12141;
wire v_12142;
wire v_12143;
wire v_12144;
wire v_12145;
wire v_12146;
wire v_12147;
wire v_12148;
wire v_12149;
wire v_12150;
wire v_12151;
wire v_12152;
wire v_12153;
wire v_12154;
wire v_12155;
wire v_12156;
wire v_12157;
wire v_12158;
wire v_12159;
wire v_12160;
wire v_12161;
wire v_12162;
wire v_12163;
wire v_12164;
wire v_12165;
wire v_12166;
wire v_12167;
wire v_12168;
wire v_12169;
wire v_12170;
wire v_12171;
wire v_12172;
wire v_12173;
wire v_12174;
wire v_12175;
wire v_12176;
wire v_12177;
wire v_12178;
wire v_12179;
wire v_12180;
wire v_12181;
wire v_12182;
wire v_12183;
wire v_12184;
wire v_12185;
wire v_12186;
wire v_12187;
wire v_12188;
wire v_12189;
wire v_12190;
wire v_12191;
wire v_12192;
wire v_12193;
wire v_12194;
wire v_12195;
wire v_12196;
wire v_12197;
wire v_12198;
wire v_12199;
wire v_12200;
wire v_12201;
wire v_12202;
wire v_12203;
wire v_12204;
wire v_12205;
wire v_12206;
wire v_12207;
wire v_12208;
wire v_12209;
wire v_12210;
wire v_12211;
wire v_12212;
wire v_12213;
wire v_12214;
wire v_12215;
wire v_12216;
wire v_12217;
wire v_12218;
wire v_12219;
wire v_12220;
wire v_12221;
wire v_12222;
wire v_12223;
wire v_12224;
wire v_12225;
wire v_12226;
wire v_12227;
wire v_12228;
wire v_12229;
wire v_12230;
wire v_12231;
wire v_12232;
wire v_12233;
wire v_12234;
wire v_12235;
wire v_12236;
wire v_12237;
wire v_12238;
wire v_12239;
wire v_12240;
wire v_12241;
wire v_12242;
wire v_12243;
wire v_12244;
wire v_12245;
wire v_12246;
wire v_12247;
wire v_12248;
wire v_12249;
wire v_12250;
wire v_12251;
wire v_12253;
wire v_12254;
wire v_12255;
wire v_12256;
wire v_12257;
wire v_12258;
wire v_12259;
wire v_12260;
wire v_12261;
wire v_12262;
wire v_12263;
wire v_12264;
wire v_12265;
wire v_12266;
wire v_12267;
wire v_12268;
wire v_12269;
wire v_12270;
wire v_12271;
wire v_12272;
wire v_12273;
wire v_12274;
wire v_12275;
wire v_12276;
wire v_12277;
wire v_12278;
wire v_12279;
wire v_12280;
wire v_12281;
wire v_12282;
wire v_12283;
wire v_12284;
wire v_12285;
wire v_12286;
wire v_12287;
wire v_12288;
wire v_12289;
wire v_12290;
wire v_12291;
wire v_12292;
wire v_12293;
wire v_12294;
wire v_12295;
wire v_12296;
wire v_12297;
wire v_12298;
wire v_12299;
wire v_12300;
wire v_12301;
wire v_12302;
wire v_12303;
wire v_12304;
wire v_12305;
wire v_12306;
wire v_12307;
wire v_12308;
wire v_12309;
wire v_12310;
wire v_12311;
wire v_12312;
wire v_12313;
wire v_12314;
wire v_12315;
wire v_12316;
wire v_12317;
wire v_12318;
wire v_12319;
wire v_12320;
wire v_12321;
wire v_12322;
wire v_12323;
wire v_12324;
wire v_12325;
wire v_12326;
wire v_12327;
wire v_12328;
wire v_12329;
wire v_12330;
wire v_12331;
wire v_12332;
wire v_12333;
wire v_12334;
wire v_12335;
wire v_12336;
wire v_12337;
wire v_12338;
wire v_12339;
wire v_12340;
wire v_12341;
wire v_12342;
wire v_12343;
wire v_12344;
wire v_12345;
wire v_12346;
wire v_12347;
wire v_12348;
wire v_12349;
wire v_12350;
wire v_12351;
wire v_12352;
wire v_12353;
wire v_12354;
wire v_12355;
wire v_12356;
wire v_12357;
wire v_12358;
wire v_12359;
wire v_12360;
wire v_12361;
wire v_12362;
wire v_12363;
wire v_12364;
wire v_12365;
wire v_12366;
wire v_12367;
wire v_12368;
wire v_12369;
wire v_12370;
wire v_12371;
wire v_12372;
wire v_12373;
wire v_12374;
wire v_12375;
wire v_12376;
wire v_12377;
wire v_12378;
wire v_12379;
wire v_12380;
wire v_12381;
wire v_12382;
wire v_12383;
wire v_12384;
wire v_12385;
wire v_12386;
wire v_12387;
wire v_12388;
wire v_12389;
wire v_12390;
wire v_12391;
wire v_12392;
wire v_12393;
wire v_12394;
wire v_12395;
wire v_12396;
wire v_12397;
wire v_12398;
wire v_12399;
wire v_12400;
wire v_12401;
wire v_12402;
wire v_12403;
wire v_12404;
wire v_12405;
wire v_12406;
wire v_12407;
wire v_12408;
wire v_12409;
wire v_12410;
wire v_12411;
wire v_12412;
wire v_12413;
wire v_12414;
wire v_12415;
wire v_12416;
wire v_12417;
wire v_12418;
wire v_12419;
wire v_12420;
wire v_12421;
wire v_12422;
wire v_12423;
wire v_12424;
wire v_12425;
wire v_12426;
wire v_12427;
wire v_12428;
wire v_12429;
wire v_12430;
wire v_12431;
wire v_12432;
wire v_12433;
wire v_12434;
wire v_12435;
wire v_12436;
wire v_12437;
wire v_12438;
wire v_12439;
wire v_12440;
wire v_12441;
wire v_12442;
wire v_12443;
wire v_12444;
wire v_12445;
wire v_12446;
wire v_12447;
wire v_12448;
wire v_12449;
wire v_12450;
wire v_12451;
wire v_12452;
wire v_12453;
wire v_12454;
wire v_12455;
wire v_12456;
wire v_12457;
wire v_12458;
wire v_12459;
wire v_12460;
wire v_12461;
wire v_12462;
wire v_12463;
wire v_12464;
wire v_12465;
wire v_12466;
wire v_12467;
wire v_12468;
wire v_12469;
wire v_12470;
wire v_12471;
wire v_12472;
wire v_12473;
wire v_12474;
wire v_12475;
wire v_12476;
wire v_12477;
wire v_12478;
wire v_12479;
wire v_12480;
wire v_12481;
wire v_12482;
wire v_12483;
wire v_12484;
wire v_12485;
wire v_12486;
wire v_12487;
wire v_12488;
wire v_12489;
wire v_12490;
wire v_12491;
wire v_12492;
wire v_12493;
wire v_12494;
wire v_12495;
wire v_12496;
wire v_12497;
wire v_12498;
wire v_12499;
wire v_12500;
wire v_12501;
wire v_12502;
wire v_12503;
wire v_12504;
wire v_12505;
wire v_12506;
wire v_12507;
wire v_12508;
wire v_12509;
wire v_12510;
wire v_12511;
wire v_12512;
wire v_12513;
wire v_12514;
wire v_12515;
wire v_12516;
wire v_12517;
wire v_12518;
wire v_12519;
wire v_12520;
wire v_12521;
wire v_12522;
wire v_12523;
wire v_12524;
wire v_12525;
wire v_12526;
wire v_12527;
wire v_12528;
wire v_12529;
wire v_12530;
wire v_12531;
wire v_12532;
wire v_12533;
wire v_12534;
wire v_12535;
wire v_12536;
wire v_12537;
wire v_12538;
wire v_12539;
wire v_12540;
wire v_12541;
wire v_12542;
wire v_12543;
wire v_12544;
wire v_12545;
wire v_12546;
wire v_12547;
wire v_12548;
wire v_12549;
wire v_12550;
wire v_12551;
wire v_12552;
wire v_12553;
wire v_12554;
wire v_12555;
wire v_12556;
wire v_12557;
wire v_12558;
wire v_12559;
wire v_12560;
wire v_12561;
wire v_12562;
wire v_12563;
wire v_12564;
wire v_12565;
wire v_12566;
wire v_12567;
wire v_12568;
wire v_12569;
wire v_12570;
wire v_12571;
wire v_12572;
wire v_12573;
wire v_12574;
wire v_12575;
wire v_12576;
wire v_12577;
wire v_12578;
wire v_12579;
wire v_12580;
wire v_12581;
wire v_12582;
wire v_12583;
wire v_12584;
wire v_12585;
wire v_12586;
wire v_12587;
wire v_12588;
wire v_12589;
wire v_12590;
wire v_12591;
wire v_12592;
wire v_12593;
wire v_12594;
wire v_12595;
wire v_12596;
wire v_12597;
wire v_12598;
wire v_12599;
wire v_12600;
wire v_12601;
wire v_12602;
wire v_12603;
wire v_12604;
wire v_12605;
wire v_12606;
wire v_12607;
wire v_12608;
wire v_12609;
wire v_12610;
wire v_12611;
wire v_12612;
wire v_12613;
wire v_12614;
wire v_12615;
wire v_12616;
wire v_12617;
wire v_12618;
wire v_12619;
wire v_12620;
wire v_12621;
wire v_12622;
wire v_12623;
wire v_12624;
wire v_12625;
wire v_12626;
wire v_12627;
wire v_12628;
wire v_12629;
wire v_12630;
wire v_12631;
wire v_12632;
wire v_12633;
wire v_12634;
wire v_12635;
wire v_12636;
wire v_12637;
wire v_12638;
wire v_12639;
wire v_12640;
wire v_12641;
wire v_12642;
wire v_12643;
wire v_12645;
wire v_12646;
wire v_12647;
wire v_12648;
wire v_12649;
wire v_12650;
wire v_12651;
wire v_12652;
wire v_12653;
wire v_12654;
wire v_12655;
wire v_12656;
wire v_12657;
wire v_12658;
wire v_12659;
wire v_12660;
wire v_12661;
wire v_12662;
wire v_12663;
wire v_12664;
wire v_12665;
wire v_12666;
wire v_12667;
wire v_12668;
wire v_12669;
wire v_12670;
wire v_12671;
wire v_12672;
wire v_12673;
wire v_12674;
wire v_12675;
wire v_12676;
wire v_12677;
wire v_12678;
wire v_12679;
wire v_12680;
wire v_12681;
wire v_12682;
wire v_12683;
wire v_12684;
wire v_12685;
wire v_12686;
wire v_12687;
wire v_12688;
wire v_12689;
wire v_12690;
wire v_12691;
wire v_12692;
wire v_12693;
wire v_12694;
wire v_12695;
wire v_12696;
wire v_12697;
wire v_12698;
wire v_12699;
wire v_12700;
wire v_12701;
wire v_12702;
wire v_12703;
wire v_12704;
wire v_12705;
wire v_12706;
wire v_12707;
wire v_12708;
wire v_12709;
wire v_12710;
wire v_12711;
wire v_12712;
wire v_12713;
wire v_12714;
wire v_12715;
wire v_12716;
wire v_12717;
wire v_12718;
wire v_12719;
wire v_12720;
wire v_12721;
wire v_12722;
wire v_12723;
wire v_12724;
wire v_12725;
wire v_12726;
wire v_12727;
wire v_12728;
wire v_12729;
wire v_12730;
wire v_12731;
wire v_12732;
wire v_12733;
wire v_12734;
wire v_12735;
wire v_12736;
wire v_12737;
wire v_12739;
wire v_12741;
wire v_12742;
wire v_12743;
wire v_12745;
wire v_12746;
wire v_12747;
wire v_12749;
wire v_12750;
wire v_12751;
wire v_12753;
wire v_12754;
wire v_12756;
wire v_12757;
wire v_12758;
wire v_12760;
wire v_12761;
wire v_12762;
wire v_12764;
wire v_12765;
wire v_12766;
wire v_12768;
wire v_12769;
wire v_12770;
wire v_12772;
wire v_12773;
wire v_12774;
wire v_12776;
wire v_12777;
wire v_12778;
wire v_12780;
wire v_12781;
wire v_12782;
wire v_12784;
wire v_12785;
wire v_12786;
wire v_12788;
wire v_12789;
wire v_12790;
wire v_12792;
wire v_12793;
wire v_12794;
wire v_12796;
wire v_12797;
wire v_12798;
wire v_12800;
wire v_12801;
wire v_12802;
wire v_12804;
wire v_12805;
wire v_12806;
wire v_12807;
wire v_12808;
wire v_12809;
wire v_12810;
wire v_12811;
wire v_12812;
wire v_12813;
wire v_12814;
wire v_12815;
wire v_12816;
wire v_12817;
wire v_12818;
wire v_12819;
wire v_12820;
wire v_12821;
wire v_12822;
wire v_12823;
wire v_12824;
wire v_12825;
wire v_12826;
wire v_12827;
wire v_12828;
wire v_12829;
wire v_12830;
wire v_12831;
wire v_12832;
wire v_12833;
wire v_12834;
wire v_12835;
wire v_12836;
wire v_12837;
wire v_12838;
wire v_12839;
wire v_12840;
wire v_12841;
wire v_12842;
wire v_12843;
wire v_12844;
wire v_12845;
wire v_12846;
wire v_12847;
wire v_12848;
wire v_12849;
wire v_12850;
wire v_12851;
wire v_12852;
wire v_12853;
wire v_12854;
wire v_12855;
wire v_12856;
wire v_12857;
wire v_12858;
wire v_12859;
wire v_12860;
wire v_12861;
wire v_12862;
wire v_12863;
wire v_12864;
wire v_12865;
wire v_12866;
wire v_12867;
wire v_12868;
wire v_12869;
wire v_12870;
wire v_12871;
wire v_12872;
wire v_12873;
wire v_12874;
wire v_12875;
wire v_12876;
wire v_12877;
wire v_12878;
wire v_12879;
wire v_12880;
wire v_12881;
wire v_12882;
wire v_12883;
wire v_12884;
wire v_12885;
wire v_12886;
wire v_12887;
wire v_12888;
wire v_12889;
wire v_12890;
wire v_12891;
wire v_12892;
wire v_12893;
wire v_12894;
wire v_12895;
wire v_12896;
wire v_12897;
wire v_12898;
wire v_12899;
wire v_12900;
wire v_12901;
wire v_12902;
wire v_12903;
wire v_12904;
wire v_12905;
wire v_12906;
wire v_12907;
wire v_12908;
wire v_12909;
wire v_12910;
wire v_12911;
wire v_12912;
wire v_12913;
wire v_12914;
wire v_12915;
wire v_12916;
wire v_12917;
wire v_12918;
wire v_12919;
wire v_12920;
wire v_12921;
wire v_12922;
wire v_12923;
wire v_12924;
wire v_12925;
wire v_12926;
wire v_12927;
wire v_12928;
wire v_12929;
wire v_12930;
wire v_12931;
wire v_12932;
wire v_12933;
wire v_12934;
wire v_12935;
wire v_12936;
wire v_12937;
wire v_12938;
wire v_12939;
wire v_12940;
wire v_12941;
wire v_12942;
wire v_12943;
wire v_12944;
wire v_12945;
wire v_12946;
wire v_12947;
wire v_12948;
wire v_12949;
wire v_12950;
wire v_12951;
wire v_12952;
wire v_12953;
wire v_12954;
wire v_12955;
wire v_12956;
wire v_12957;
wire v_12958;
wire v_12959;
wire v_12960;
wire v_12961;
wire v_12962;
wire v_12963;
wire v_12964;
wire v_12965;
wire v_12966;
wire v_12967;
wire v_12968;
wire v_12969;
wire v_12970;
wire v_12971;
wire v_12972;
wire v_12973;
wire v_12974;
wire v_12975;
wire v_12976;
wire v_12977;
wire v_12978;
wire v_12979;
wire v_12980;
wire v_12981;
wire v_12982;
wire v_12983;
wire v_12984;
wire v_12985;
wire v_12986;
wire v_12987;
wire v_12988;
wire v_12989;
wire v_12990;
wire v_12991;
wire v_12992;
wire v_12993;
wire v_12994;
wire v_12995;
wire v_12996;
wire v_12997;
wire v_12999;
wire v_13000;
wire v_13001;
wire v_13002;
wire v_13003;
wire v_13004;
wire v_13005;
wire v_13006;
wire v_13007;
wire v_13008;
wire v_13009;
wire v_13010;
wire v_13011;
wire v_13012;
wire v_13013;
wire v_13014;
wire v_13015;
wire v_13016;
wire v_13017;
wire v_13018;
wire v_13019;
wire v_13020;
wire v_13021;
wire v_13022;
wire v_13023;
wire v_13024;
wire v_13025;
wire v_13026;
wire v_13027;
wire v_13028;
wire v_13029;
wire v_13030;
wire v_13031;
wire v_13032;
wire v_13033;
wire v_13034;
wire v_13035;
wire v_13036;
wire v_13037;
wire v_13038;
wire v_13039;
wire v_13040;
wire v_13041;
wire v_13042;
wire v_13043;
wire v_13044;
wire v_13045;
wire v_13046;
wire v_13047;
wire v_13048;
wire v_13049;
wire v_13050;
wire v_13051;
wire v_13052;
wire v_13053;
wire v_13054;
wire v_13055;
wire v_13056;
wire v_13057;
wire v_13058;
wire v_13059;
wire v_13060;
wire v_13061;
wire v_13062;
wire v_13063;
wire v_13064;
wire v_13065;
wire v_13066;
wire v_13067;
wire v_13068;
wire v_13069;
wire v_13070;
wire v_13071;
wire v_13072;
wire v_13073;
wire v_13074;
wire v_13075;
wire v_13076;
wire v_13077;
wire v_13078;
wire v_13079;
wire v_13080;
wire v_13081;
wire v_13082;
wire v_13083;
wire v_13084;
wire v_13085;
wire v_13086;
wire v_13087;
wire v_13088;
wire v_13089;
wire v_13090;
wire v_13091;
wire v_13092;
wire v_13093;
wire v_13094;
wire v_13095;
wire v_13096;
wire v_13097;
wire v_13098;
wire v_13099;
wire v_13100;
wire v_13101;
wire v_13102;
wire v_13103;
wire v_13104;
wire v_13105;
wire v_13106;
wire v_13107;
wire v_13108;
wire v_13109;
wire v_13110;
wire v_13111;
wire v_13112;
wire v_13113;
wire v_13114;
wire v_13115;
wire v_13116;
wire v_13117;
wire v_13118;
wire v_13119;
wire v_13120;
wire v_13121;
wire v_13122;
wire v_13123;
wire v_13124;
wire v_13125;
wire v_13126;
wire v_13127;
wire v_13128;
wire v_13129;
wire v_13130;
wire v_13131;
wire v_13132;
wire v_13133;
wire v_13134;
wire v_13135;
wire v_13136;
wire v_13137;
wire v_13138;
wire v_13139;
wire v_13140;
wire v_13141;
wire v_13142;
wire v_13143;
wire v_13144;
wire v_13145;
wire v_13146;
wire v_13147;
wire v_13148;
wire v_13149;
wire v_13150;
wire v_13151;
wire v_13152;
wire v_13153;
wire v_13154;
wire v_13155;
wire v_13156;
wire v_13157;
wire v_13158;
wire v_13159;
wire v_13160;
wire v_13161;
wire v_13162;
wire v_13163;
wire v_13164;
wire v_13165;
wire v_13166;
wire v_13167;
wire v_13168;
wire v_13169;
wire v_13170;
wire v_13171;
wire v_13172;
wire v_13173;
wire v_13174;
wire v_13175;
wire v_13176;
wire v_13177;
wire v_13178;
wire v_13179;
wire v_13180;
wire v_13181;
wire v_13182;
wire v_13183;
wire v_13184;
wire v_13185;
wire v_13186;
wire v_13187;
wire v_13188;
wire v_13189;
wire v_13190;
wire v_13191;
wire v_13192;
wire v_13193;
wire v_13194;
wire v_13195;
wire v_13196;
wire v_13197;
wire v_13198;
wire v_13199;
wire v_13200;
wire v_13201;
wire v_13202;
wire v_13203;
wire v_13204;
wire v_13205;
wire v_13206;
wire v_13207;
wire v_13208;
wire v_13209;
wire v_13210;
wire v_13211;
wire v_13212;
wire v_13213;
wire v_13214;
wire v_13215;
wire v_13216;
wire v_13217;
wire v_13218;
wire v_13219;
wire v_13220;
wire v_13221;
wire v_13222;
wire v_13223;
wire v_13224;
wire v_13225;
wire v_13226;
wire v_13227;
wire v_13228;
wire v_13229;
wire v_13230;
wire v_13231;
wire v_13232;
wire v_13233;
wire v_13234;
wire v_13235;
wire v_13236;
wire v_13237;
wire v_13238;
wire v_13239;
wire v_13240;
wire v_13242;
wire v_13243;
wire v_13244;
wire v_13245;
wire v_13246;
wire v_13247;
wire v_13248;
wire v_13249;
wire v_13250;
wire v_13251;
wire v_13252;
wire v_13253;
wire v_13254;
wire v_13255;
wire v_13256;
wire v_13257;
wire v_13258;
wire v_13259;
wire v_13260;
wire v_13261;
wire v_13262;
wire v_13263;
wire v_13264;
wire v_13265;
wire v_13266;
wire v_13267;
wire v_13268;
wire v_13269;
wire v_13270;
wire v_13271;
wire v_13272;
wire v_13273;
wire v_13274;
wire v_13275;
wire v_13276;
wire v_13277;
wire v_13278;
wire v_13279;
wire v_13280;
wire v_13281;
wire v_13282;
wire v_13283;
wire v_13284;
wire v_13285;
wire v_13286;
wire v_13287;
wire v_13288;
wire v_13289;
wire v_13290;
wire v_13291;
wire v_13292;
wire v_13293;
wire v_13294;
wire v_13295;
wire v_13296;
wire v_13297;
wire v_13298;
wire v_13299;
wire v_13300;
wire v_13301;
wire v_13302;
wire v_13303;
wire v_13304;
wire v_13305;
wire v_13306;
wire v_13307;
wire v_13308;
wire v_13309;
wire v_13310;
wire v_13311;
wire v_13312;
wire v_13313;
wire v_13314;
wire v_13315;
wire v_13316;
wire v_13317;
wire v_13318;
wire v_13319;
wire v_13320;
wire v_13321;
wire v_13322;
wire v_13323;
wire v_13324;
wire v_13325;
wire v_13326;
wire v_13327;
wire v_13328;
wire v_13329;
wire v_13330;
wire v_13331;
wire v_13332;
wire v_13333;
wire v_13334;
wire v_13335;
wire v_13336;
wire v_13337;
wire v_13338;
wire v_13339;
wire v_13340;
wire v_13341;
wire v_13342;
wire v_13343;
wire v_13344;
wire v_13345;
wire v_13346;
wire v_13347;
wire v_13348;
wire v_13349;
wire v_13350;
wire v_13351;
wire v_13352;
wire v_13353;
wire v_13354;
wire v_13355;
wire v_13356;
wire v_13357;
wire v_13358;
wire v_13359;
wire v_13360;
wire v_13361;
wire v_13362;
wire v_13363;
wire v_13364;
wire v_13365;
wire v_13366;
wire v_13367;
wire v_13368;
wire v_13369;
wire v_13370;
wire v_13371;
wire v_13372;
wire v_13373;
wire v_13374;
wire v_13375;
wire v_13376;
wire v_13377;
wire v_13378;
wire v_13379;
wire v_13380;
wire v_13381;
wire v_13382;
wire v_13383;
wire v_13384;
wire v_13385;
wire v_13386;
wire v_13387;
wire v_13388;
wire v_13389;
wire v_13390;
wire v_13391;
wire v_13392;
wire v_13393;
wire v_13394;
wire v_13395;
wire v_13396;
wire v_13397;
wire v_13398;
wire v_13399;
wire v_13400;
wire v_13401;
wire v_13402;
wire v_13403;
wire v_13404;
wire v_13405;
wire v_13406;
wire v_13407;
wire v_13408;
wire v_13409;
wire v_13410;
wire v_13411;
wire v_13412;
wire v_13413;
wire v_13414;
wire v_13415;
wire v_13416;
wire v_13417;
wire v_13418;
wire v_13419;
wire v_13420;
wire v_13421;
wire v_13422;
wire v_13423;
wire v_13424;
wire v_13425;
wire v_13426;
wire v_13427;
wire v_13428;
wire v_13429;
wire v_13430;
wire v_13431;
wire v_13432;
wire v_13433;
wire v_13434;
wire v_13435;
wire v_13436;
wire v_13437;
wire v_13438;
wire v_13439;
wire v_13440;
wire v_13441;
wire v_13442;
wire v_13443;
wire v_13444;
wire v_13445;
wire v_13446;
wire v_13447;
wire v_13448;
wire v_13449;
wire v_13450;
wire v_13451;
wire v_13452;
wire v_13453;
wire v_13454;
wire v_13455;
wire v_13456;
wire v_13457;
wire v_13458;
wire v_13459;
wire v_13460;
wire v_13461;
wire v_13462;
wire v_13463;
wire v_13464;
wire v_13465;
wire v_13466;
wire v_13467;
wire v_13468;
wire v_13469;
wire v_13470;
wire v_13471;
wire v_13472;
wire v_13473;
wire v_13474;
wire v_13475;
wire v_13476;
wire v_13477;
wire v_13478;
wire v_13479;
wire v_13480;
wire v_13481;
wire v_13482;
wire v_13483;
wire v_13485;
wire v_13486;
wire v_13487;
wire v_13488;
wire v_13489;
wire v_13490;
wire v_13491;
wire v_13492;
wire v_13493;
wire v_13494;
wire v_13495;
wire v_13496;
wire v_13497;
wire v_13498;
wire v_13499;
wire v_13500;
wire v_13501;
wire v_13502;
wire v_13503;
wire v_13504;
wire v_13505;
wire v_13506;
wire v_13507;
wire v_13508;
wire v_13509;
wire v_13510;
wire v_13511;
wire v_13512;
wire v_13513;
wire v_13514;
wire v_13515;
wire v_13516;
wire v_13517;
wire v_13518;
wire v_13519;
wire v_13520;
wire v_13521;
wire v_13522;
wire v_13523;
wire v_13524;
wire v_13525;
wire v_13526;
wire v_13527;
wire v_13528;
wire v_13529;
wire v_13530;
wire v_13531;
wire v_13532;
wire v_13533;
wire v_13534;
wire v_13535;
wire v_13536;
wire v_13537;
wire v_13538;
wire v_13539;
wire v_13540;
wire v_13541;
wire v_13542;
wire v_13543;
wire v_13544;
wire v_13545;
wire v_13546;
wire v_13547;
wire v_13548;
wire v_13549;
wire v_13550;
wire v_13551;
wire v_13552;
wire v_13553;
wire v_13554;
wire v_13555;
wire v_13556;
wire v_13557;
wire v_13558;
wire v_13559;
wire v_13560;
wire v_13561;
wire v_13562;
wire v_13563;
wire v_13564;
wire v_13565;
wire v_13566;
wire v_13567;
wire v_13568;
wire v_13569;
wire v_13570;
wire v_13571;
wire v_13572;
wire v_13573;
wire v_13574;
wire v_13575;
wire v_13576;
wire v_13577;
wire v_13578;
wire v_13579;
wire v_13580;
wire v_13581;
wire v_13582;
wire v_13583;
wire v_13584;
wire v_13585;
wire v_13586;
wire v_13587;
wire v_13588;
wire v_13589;
wire v_13590;
wire v_13591;
wire v_13592;
wire v_13593;
wire v_13594;
wire v_13595;
wire v_13596;
wire v_13597;
wire v_13598;
wire v_13599;
wire v_13600;
wire v_13601;
wire v_13602;
wire v_13603;
wire v_13604;
wire v_13605;
wire v_13606;
wire v_13607;
wire v_13608;
wire v_13609;
wire v_13610;
wire v_13611;
wire v_13612;
wire v_13613;
wire v_13614;
wire v_13615;
wire v_13616;
wire v_13617;
wire v_13618;
wire v_13619;
wire v_13620;
wire v_13621;
wire v_13622;
wire v_13623;
wire v_13624;
wire v_13625;
wire v_13626;
wire v_13627;
wire v_13628;
wire v_13629;
wire v_13630;
wire v_13631;
wire v_13632;
wire v_13633;
wire v_13634;
wire v_13635;
wire v_13636;
wire v_13637;
wire v_13638;
wire v_13639;
wire v_13640;
wire v_13641;
wire v_13642;
wire v_13643;
wire v_13644;
wire v_13645;
wire v_13646;
wire v_13647;
wire v_13648;
wire v_13649;
wire v_13650;
wire v_13651;
wire v_13652;
wire v_13653;
wire v_13654;
wire v_13655;
wire v_13656;
wire v_13657;
wire v_13658;
wire v_13659;
wire v_13660;
wire v_13661;
wire v_13662;
wire v_13663;
wire v_13664;
wire v_13665;
wire v_13666;
wire v_13667;
wire v_13668;
wire v_13669;
wire v_13670;
wire v_13671;
wire v_13672;
wire v_13673;
wire v_13674;
wire v_13675;
wire v_13676;
wire v_13677;
wire v_13678;
wire v_13679;
wire v_13680;
wire v_13681;
wire v_13682;
wire v_13683;
wire v_13684;
wire v_13685;
wire v_13686;
wire v_13687;
wire v_13688;
wire v_13689;
wire v_13690;
wire v_13691;
wire v_13692;
wire v_13693;
wire v_13694;
wire v_13695;
wire v_13696;
wire v_13697;
wire v_13698;
wire v_13699;
wire v_13700;
wire v_13701;
wire v_13702;
wire v_13703;
wire v_13704;
wire v_13705;
wire v_13706;
wire v_13707;
wire v_13708;
wire v_13709;
wire v_13710;
wire v_13711;
wire v_13712;
wire v_13713;
wire v_13714;
wire v_13715;
wire v_13716;
wire v_13717;
wire v_13718;
wire v_13719;
wire v_13720;
wire v_13721;
wire v_13722;
wire v_13723;
wire v_13724;
wire v_13725;
wire v_13726;
wire v_13728;
wire v_13729;
wire v_13730;
wire v_13731;
wire v_13732;
wire v_13733;
wire v_13734;
wire v_13735;
wire v_13736;
wire v_13737;
wire v_13738;
wire v_13739;
wire v_13740;
wire v_13741;
wire v_13742;
wire v_13743;
wire v_13744;
wire v_13745;
wire v_13746;
wire v_13747;
wire v_13748;
wire v_13749;
wire v_13750;
wire v_13751;
wire v_13752;
wire v_13753;
wire v_13754;
wire v_13755;
wire v_13756;
wire v_13757;
wire v_13758;
wire v_13759;
wire v_13760;
wire v_13761;
wire v_13762;
wire v_13763;
wire v_13764;
wire v_13765;
wire v_13766;
wire v_13767;
wire v_13768;
wire v_13769;
wire v_13770;
wire v_13771;
wire v_13772;
wire v_13773;
wire v_13774;
wire v_13775;
wire v_13776;
wire v_13777;
wire v_13778;
wire v_13779;
wire v_13780;
wire v_13781;
wire v_13782;
wire v_13783;
wire v_13784;
wire v_13785;
wire v_13786;
wire v_13787;
wire v_13788;
wire v_13789;
wire v_13790;
wire v_13791;
wire v_13792;
wire v_13793;
wire v_13794;
wire v_13795;
wire v_13796;
wire v_13797;
wire v_13798;
wire v_13799;
wire v_13800;
wire v_13801;
wire v_13802;
wire v_13803;
wire v_13804;
wire v_13805;
wire v_13806;
wire v_13807;
wire v_13808;
wire v_13809;
wire v_13810;
wire v_13811;
wire v_13812;
wire v_13813;
wire v_13814;
wire v_13815;
wire v_13816;
wire v_13817;
wire v_13818;
wire v_13819;
wire v_13820;
wire v_13821;
wire v_13822;
wire v_13823;
wire v_13824;
wire v_13825;
wire v_13826;
wire v_13827;
wire v_13828;
wire v_13829;
wire v_13830;
wire v_13831;
wire v_13832;
wire v_13833;
wire v_13834;
wire v_13835;
wire v_13836;
wire v_13837;
wire v_13838;
wire v_13839;
wire v_13840;
wire v_13841;
wire v_13842;
wire v_13843;
wire v_13844;
wire v_13845;
wire v_13846;
wire v_13847;
wire v_13848;
wire v_13849;
wire v_13850;
wire v_13851;
wire v_13852;
wire v_13853;
wire v_13854;
wire v_13855;
wire v_13856;
wire v_13857;
wire v_13858;
wire v_13859;
wire v_13860;
wire v_13861;
wire v_13862;
wire v_13863;
wire v_13864;
wire v_13865;
wire v_13866;
wire v_13867;
wire v_13868;
wire v_13869;
wire v_13870;
wire v_13871;
wire v_13872;
wire v_13873;
wire v_13874;
wire v_13875;
wire v_13876;
wire v_13877;
wire v_13878;
wire v_13879;
wire v_13880;
wire v_13881;
wire v_13882;
wire v_13883;
wire v_13884;
wire v_13885;
wire v_13886;
wire v_13887;
wire v_13888;
wire v_13889;
wire v_13890;
wire v_13891;
wire v_13892;
wire v_13893;
wire v_13894;
wire v_13895;
wire v_13896;
wire v_13897;
wire v_13898;
wire v_13899;
wire v_13900;
wire v_13901;
wire v_13902;
wire v_13903;
wire v_13904;
wire v_13905;
wire v_13906;
wire v_13907;
wire v_13908;
wire v_13909;
wire v_13910;
wire v_13911;
wire v_13912;
wire v_13913;
wire v_13914;
wire v_13915;
wire v_13916;
wire v_13917;
wire v_13918;
wire v_13919;
wire v_13920;
wire v_13921;
wire v_13922;
wire v_13923;
wire v_13924;
wire v_13925;
wire v_13926;
wire v_13927;
wire v_13928;
wire v_13929;
wire v_13930;
wire v_13931;
wire v_13932;
wire v_13933;
wire v_13934;
wire v_13935;
wire v_13936;
wire v_13937;
wire v_13938;
wire v_13939;
wire v_13940;
wire v_13941;
wire v_13942;
wire v_13943;
wire v_13944;
wire v_13945;
wire v_13946;
wire v_13947;
wire v_13948;
wire v_13949;
wire v_13950;
wire v_13951;
wire v_13952;
wire v_13953;
wire v_13954;
wire v_13955;
wire v_13956;
wire v_13957;
wire v_13958;
wire v_13959;
wire v_13960;
wire v_13961;
wire v_13962;
wire v_13963;
wire v_13964;
wire v_13965;
wire v_13966;
wire v_13967;
wire v_13968;
wire v_13969;
wire v_13971;
wire v_13972;
wire v_13973;
wire v_13974;
wire v_13975;
wire v_13976;
wire v_13977;
wire v_13978;
wire v_13979;
wire v_13980;
wire v_13981;
wire v_13982;
wire v_13983;
wire v_13984;
wire v_13985;
wire v_13986;
wire v_13987;
wire v_13988;
wire v_13989;
wire v_13990;
wire v_13991;
wire v_13992;
wire v_13993;
wire v_13994;
wire v_13995;
wire v_13996;
wire v_13997;
wire v_13998;
wire v_13999;
wire v_14000;
wire v_14001;
wire v_14002;
wire v_14003;
wire v_14004;
wire v_14005;
wire v_14006;
wire v_14007;
wire v_14008;
wire v_14009;
wire v_14010;
wire v_14011;
wire v_14012;
wire v_14013;
wire v_14014;
wire v_14015;
wire v_14016;
wire v_14017;
wire v_14018;
wire v_14019;
wire v_14020;
wire v_14021;
wire v_14022;
wire v_14023;
wire v_14024;
wire v_14025;
wire v_14026;
wire v_14027;
wire v_14028;
wire v_14029;
wire v_14030;
wire v_14031;
wire v_14032;
wire v_14033;
wire v_14034;
wire v_14035;
wire v_14036;
wire v_14037;
wire v_14038;
wire v_14039;
wire v_14040;
wire v_14041;
wire v_14042;
wire v_14043;
wire v_14044;
wire v_14045;
wire v_14046;
wire v_14047;
wire v_14048;
wire v_14049;
wire v_14050;
wire v_14051;
wire v_14052;
wire v_14053;
wire v_14054;
wire v_14055;
wire v_14056;
wire v_14057;
wire v_14058;
wire v_14059;
wire v_14060;
wire v_14061;
wire v_14062;
wire v_14063;
wire v_14064;
wire v_14065;
wire v_14066;
wire v_14067;
wire v_14068;
wire v_14069;
wire v_14070;
wire v_14071;
wire v_14072;
wire v_14073;
wire v_14074;
wire v_14075;
wire v_14076;
wire v_14077;
wire v_14078;
wire v_14079;
wire v_14080;
wire v_14081;
wire v_14082;
wire v_14083;
wire v_14084;
wire v_14085;
wire v_14086;
wire v_14087;
wire v_14088;
wire v_14089;
wire v_14090;
wire v_14091;
wire v_14092;
wire v_14093;
wire v_14094;
wire v_14095;
wire v_14096;
wire v_14097;
wire v_14098;
wire v_14099;
wire v_14100;
wire v_14101;
wire v_14102;
wire v_14103;
wire v_14104;
wire v_14105;
wire v_14106;
wire v_14107;
wire v_14108;
wire v_14109;
wire v_14110;
wire v_14111;
wire v_14112;
wire v_14113;
wire v_14114;
wire v_14115;
wire v_14116;
wire v_14117;
wire v_14118;
wire v_14119;
wire v_14120;
wire v_14121;
wire v_14122;
wire v_14123;
wire v_14124;
wire v_14125;
wire v_14126;
wire v_14127;
wire v_14128;
wire v_14129;
wire v_14130;
wire v_14131;
wire v_14132;
wire v_14133;
wire v_14134;
wire v_14135;
wire v_14136;
wire v_14137;
wire v_14138;
wire v_14139;
wire v_14140;
wire v_14141;
wire v_14142;
wire v_14143;
wire v_14144;
wire v_14145;
wire v_14146;
wire v_14147;
wire v_14148;
wire v_14149;
wire v_14150;
wire v_14151;
wire v_14152;
wire v_14153;
wire v_14154;
wire v_14155;
wire v_14156;
wire v_14157;
wire v_14158;
wire v_14159;
wire v_14160;
wire v_14161;
wire v_14162;
wire v_14163;
wire v_14164;
wire v_14165;
wire v_14166;
wire v_14167;
wire v_14168;
wire v_14169;
wire v_14170;
wire v_14171;
wire v_14172;
wire v_14173;
wire v_14174;
wire v_14175;
wire v_14176;
wire v_14177;
wire v_14178;
wire v_14179;
wire v_14180;
wire v_14181;
wire v_14182;
wire v_14183;
wire v_14184;
wire v_14185;
wire v_14186;
wire v_14187;
wire v_14188;
wire v_14189;
wire v_14190;
wire v_14191;
wire v_14192;
wire v_14193;
wire v_14194;
wire v_14195;
wire v_14196;
wire v_14197;
wire v_14198;
wire v_14199;
wire v_14200;
wire v_14201;
wire v_14202;
wire v_14203;
wire v_14204;
wire v_14205;
wire v_14206;
wire v_14207;
wire v_14208;
wire v_14209;
wire v_14210;
wire v_14211;
wire v_14212;
wire v_14214;
wire v_14215;
wire v_14216;
wire v_14217;
wire v_14218;
wire v_14219;
wire v_14220;
wire v_14221;
wire v_14222;
wire v_14223;
wire v_14224;
wire v_14225;
wire v_14226;
wire v_14227;
wire v_14228;
wire v_14229;
wire v_14230;
wire v_14231;
wire v_14232;
wire v_14233;
wire v_14234;
wire v_14235;
wire v_14236;
wire v_14237;
wire v_14238;
wire v_14239;
wire v_14240;
wire v_14241;
wire v_14242;
wire v_14243;
wire v_14244;
wire v_14245;
wire v_14246;
wire v_14247;
wire v_14248;
wire v_14249;
wire v_14250;
wire v_14251;
wire v_14252;
wire v_14253;
wire v_14254;
wire v_14255;
wire v_14256;
wire v_14257;
wire v_14258;
wire v_14259;
wire v_14260;
wire v_14261;
wire v_14262;
wire v_14263;
wire v_14264;
wire v_14265;
wire v_14266;
wire v_14267;
wire v_14268;
wire v_14269;
wire v_14270;
wire v_14271;
wire v_14272;
wire v_14273;
wire v_14274;
wire v_14275;
wire v_14276;
wire v_14277;
wire v_14278;
wire v_14279;
wire v_14280;
wire v_14281;
wire v_14282;
wire v_14283;
wire v_14284;
wire v_14285;
wire v_14286;
wire v_14287;
wire v_14288;
wire v_14289;
wire v_14290;
wire v_14291;
wire v_14292;
wire v_14293;
wire v_14294;
wire v_14295;
wire v_14296;
wire v_14297;
wire v_14298;
wire v_14299;
wire v_14300;
wire v_14301;
wire v_14302;
wire v_14303;
wire v_14304;
wire v_14305;
wire v_14306;
wire v_14307;
wire v_14308;
wire v_14309;
wire v_14310;
wire v_14311;
wire v_14312;
wire v_14313;
wire v_14314;
wire v_14315;
wire v_14316;
wire v_14317;
wire v_14318;
wire v_14319;
wire v_14320;
wire v_14321;
wire v_14322;
wire v_14323;
wire v_14324;
wire v_14325;
wire v_14326;
wire v_14327;
wire v_14328;
wire v_14329;
wire v_14330;
wire v_14331;
wire v_14332;
wire v_14333;
wire v_14334;
wire v_14335;
wire v_14336;
wire v_14337;
wire v_14338;
wire v_14339;
wire v_14340;
wire v_14341;
wire v_14342;
wire v_14343;
wire v_14344;
wire v_14345;
wire v_14346;
wire v_14347;
wire v_14348;
wire v_14349;
wire v_14350;
wire v_14351;
wire v_14352;
wire v_14353;
wire v_14354;
wire v_14355;
wire v_14356;
wire v_14357;
wire v_14358;
wire v_14359;
wire v_14360;
wire v_14361;
wire v_14362;
wire v_14363;
wire v_14364;
wire v_14365;
wire v_14366;
wire v_14367;
wire v_14368;
wire v_14369;
wire v_14370;
wire v_14371;
wire v_14372;
wire v_14373;
wire v_14374;
wire v_14375;
wire v_14376;
wire v_14377;
wire v_14378;
wire v_14379;
wire v_14380;
wire v_14381;
wire v_14382;
wire v_14383;
wire v_14384;
wire v_14385;
wire v_14386;
wire v_14387;
wire v_14388;
wire v_14389;
wire v_14390;
wire v_14391;
wire v_14392;
wire v_14393;
wire v_14394;
wire v_14395;
wire v_14396;
wire v_14397;
wire v_14398;
wire v_14399;
wire v_14400;
wire v_14401;
wire v_14402;
wire v_14403;
wire v_14404;
wire v_14405;
wire v_14406;
wire v_14407;
wire v_14408;
wire v_14409;
wire v_14410;
wire v_14411;
wire v_14412;
wire v_14413;
wire v_14414;
wire v_14415;
wire v_14416;
wire v_14417;
wire v_14418;
wire v_14419;
wire v_14420;
wire v_14421;
wire v_14422;
wire v_14423;
wire v_14424;
wire v_14425;
wire v_14426;
wire v_14427;
wire v_14428;
wire v_14429;
wire v_14430;
wire v_14431;
wire v_14432;
wire v_14433;
wire v_14434;
wire v_14435;
wire v_14436;
wire v_14437;
wire v_14438;
wire v_14439;
wire v_14440;
wire v_14441;
wire v_14442;
wire v_14443;
wire v_14444;
wire v_14445;
wire v_14446;
wire v_14447;
wire v_14448;
wire v_14449;
wire v_14450;
wire v_14451;
wire v_14452;
wire v_14453;
wire v_14454;
wire v_14455;
wire v_14457;
wire v_14458;
wire v_14459;
wire v_14460;
wire v_14461;
wire v_14462;
wire v_14463;
wire v_14464;
wire v_14465;
wire v_14466;
wire v_14467;
wire v_14468;
wire v_14469;
wire v_14470;
wire v_14471;
wire v_14472;
wire v_14473;
wire v_14474;
wire v_14475;
wire v_14476;
wire v_14477;
wire v_14478;
wire v_14479;
wire v_14480;
wire v_14481;
wire v_14482;
wire v_14483;
wire v_14484;
wire v_14485;
wire v_14486;
wire v_14487;
wire v_14488;
wire v_14489;
wire v_14490;
wire v_14491;
wire v_14492;
wire v_14493;
wire v_14494;
wire v_14495;
wire v_14496;
wire v_14497;
wire v_14498;
wire v_14499;
wire v_14500;
wire v_14501;
wire v_14502;
wire v_14503;
wire v_14504;
wire v_14505;
wire v_14506;
wire v_14507;
wire v_14508;
wire v_14509;
wire v_14510;
wire v_14511;
wire v_14512;
wire v_14513;
wire v_14514;
wire v_14515;
wire v_14516;
wire v_14517;
wire v_14518;
wire v_14519;
wire v_14520;
wire v_14521;
wire v_14522;
wire v_14523;
wire v_14524;
wire v_14525;
wire v_14526;
wire v_14527;
wire v_14528;
wire v_14529;
wire v_14530;
wire v_14531;
wire v_14532;
wire v_14533;
wire v_14534;
wire v_14535;
wire v_14536;
wire v_14537;
wire v_14538;
wire v_14539;
wire v_14540;
wire v_14541;
wire v_14542;
wire v_14543;
wire v_14544;
wire v_14545;
wire v_14546;
wire v_14547;
wire v_14548;
wire v_14549;
wire v_14550;
wire v_14551;
wire v_14552;
wire v_14553;
wire v_14554;
wire v_14555;
wire v_14556;
wire v_14557;
wire v_14558;
wire v_14559;
wire v_14560;
wire v_14561;
wire v_14562;
wire v_14563;
wire v_14564;
wire v_14565;
wire v_14566;
wire v_14567;
wire v_14568;
wire v_14569;
wire v_14570;
wire v_14571;
wire v_14572;
wire v_14573;
wire v_14574;
wire v_14575;
wire v_14576;
wire v_14577;
wire v_14578;
wire v_14579;
wire v_14580;
wire v_14581;
wire v_14582;
wire v_14583;
wire v_14584;
wire v_14585;
wire v_14586;
wire v_14587;
wire v_14588;
wire v_14589;
wire v_14590;
wire v_14591;
wire v_14592;
wire v_14593;
wire v_14594;
wire v_14595;
wire v_14596;
wire v_14597;
wire v_14598;
wire v_14599;
wire v_14600;
wire v_14601;
wire v_14602;
wire v_14603;
wire v_14604;
wire v_14605;
wire v_14606;
wire v_14607;
wire v_14608;
wire v_14609;
wire v_14610;
wire v_14611;
wire v_14612;
wire v_14613;
wire v_14614;
wire v_14615;
wire v_14616;
wire v_14617;
wire v_14618;
wire v_14619;
wire v_14620;
wire v_14621;
wire v_14622;
wire v_14623;
wire v_14624;
wire v_14625;
wire v_14626;
wire v_14627;
wire v_14628;
wire v_14629;
wire v_14630;
wire v_14631;
wire v_14632;
wire v_14633;
wire v_14634;
wire v_14635;
wire v_14636;
wire v_14637;
wire v_14638;
wire v_14639;
wire v_14640;
wire v_14641;
wire v_14642;
wire v_14643;
wire v_14644;
wire v_14645;
wire v_14646;
wire v_14647;
wire v_14648;
wire v_14649;
wire v_14650;
wire v_14651;
wire v_14652;
wire v_14653;
wire v_14654;
wire v_14655;
wire v_14656;
wire v_14657;
wire v_14658;
wire v_14659;
wire v_14660;
wire v_14661;
wire v_14662;
wire v_14663;
wire v_14664;
wire v_14665;
wire v_14666;
wire v_14667;
wire v_14668;
wire v_14669;
wire v_14670;
wire v_14671;
wire v_14672;
wire v_14673;
wire v_14674;
wire v_14675;
wire v_14676;
wire v_14677;
wire v_14678;
wire v_14679;
wire v_14680;
wire v_14681;
wire v_14682;
wire v_14683;
wire v_14684;
wire v_14685;
wire v_14686;
wire v_14687;
wire v_14688;
wire v_14689;
wire v_14690;
wire v_14691;
wire v_14692;
wire v_14693;
wire v_14694;
wire v_14695;
wire v_14696;
wire v_14697;
wire v_14698;
wire v_14700;
wire v_14701;
wire v_14702;
wire v_14703;
wire v_14704;
wire v_14705;
wire v_14706;
wire v_14707;
wire v_14708;
wire v_14709;
wire v_14710;
wire v_14711;
wire v_14712;
wire v_14713;
wire v_14714;
wire v_14715;
wire v_14716;
wire v_14717;
wire v_14718;
wire v_14719;
wire v_14720;
wire v_14721;
wire v_14722;
wire v_14723;
wire v_14724;
wire v_14725;
wire v_14726;
wire v_14727;
wire v_14728;
wire v_14729;
wire v_14730;
wire v_14731;
wire v_14732;
wire v_14733;
wire v_14734;
wire v_14735;
wire v_14736;
wire v_14737;
wire v_14738;
wire v_14739;
wire v_14740;
wire v_14741;
wire v_14742;
wire v_14743;
wire v_14744;
wire v_14745;
wire v_14746;
wire v_14747;
wire v_14748;
wire v_14749;
wire v_14750;
wire v_14751;
wire v_14752;
wire v_14753;
wire v_14754;
wire v_14755;
wire v_14756;
wire v_14757;
wire v_14758;
wire v_14759;
wire v_14760;
wire v_14761;
wire v_14762;
wire v_14763;
wire v_14764;
wire v_14765;
wire v_14766;
wire v_14767;
wire v_14768;
wire v_14769;
wire v_14770;
wire v_14771;
wire v_14772;
wire v_14773;
wire v_14774;
wire v_14775;
wire v_14776;
wire v_14777;
wire v_14778;
wire v_14779;
wire v_14780;
wire v_14781;
wire v_14782;
wire v_14783;
wire v_14784;
wire v_14785;
wire v_14786;
wire v_14787;
wire v_14788;
wire v_14789;
wire v_14790;
wire v_14791;
wire v_14792;
wire v_14793;
wire v_14794;
wire v_14795;
wire v_14796;
wire v_14797;
wire v_14798;
wire v_14799;
wire v_14800;
wire v_14801;
wire v_14802;
wire v_14803;
wire v_14804;
wire v_14805;
wire v_14806;
wire v_14807;
wire v_14808;
wire v_14809;
wire v_14810;
wire v_14811;
wire v_14812;
wire v_14813;
wire v_14814;
wire v_14815;
wire v_14816;
wire v_14817;
wire v_14818;
wire v_14819;
wire v_14820;
wire v_14821;
wire v_14822;
wire v_14823;
wire v_14824;
wire v_14825;
wire v_14826;
wire v_14827;
wire v_14828;
wire v_14829;
wire v_14830;
wire v_14831;
wire v_14832;
wire v_14833;
wire v_14834;
wire v_14835;
wire v_14836;
wire v_14837;
wire v_14838;
wire v_14839;
wire v_14840;
wire v_14841;
wire v_14842;
wire v_14843;
wire v_14844;
wire v_14845;
wire v_14846;
wire v_14847;
wire v_14848;
wire v_14849;
wire v_14850;
wire v_14851;
wire v_14852;
wire v_14853;
wire v_14854;
wire v_14855;
wire v_14856;
wire v_14857;
wire v_14858;
wire v_14859;
wire v_14860;
wire v_14861;
wire v_14862;
wire v_14863;
wire v_14864;
wire v_14865;
wire v_14866;
wire v_14867;
wire v_14868;
wire v_14869;
wire v_14870;
wire v_14871;
wire v_14872;
wire v_14873;
wire v_14874;
wire v_14875;
wire v_14876;
wire v_14877;
wire v_14878;
wire v_14879;
wire v_14880;
wire v_14881;
wire v_14882;
wire v_14883;
wire v_14884;
wire v_14885;
wire v_14886;
wire v_14887;
wire v_14888;
wire v_14889;
wire v_14890;
wire v_14891;
wire v_14892;
wire v_14893;
wire v_14894;
wire v_14895;
wire v_14896;
wire v_14897;
wire v_14898;
wire v_14899;
wire v_14900;
wire v_14901;
wire v_14902;
wire v_14903;
wire v_14904;
wire v_14905;
wire v_14906;
wire v_14907;
wire v_14908;
wire v_14909;
wire v_14910;
wire v_14911;
wire v_14912;
wire v_14913;
wire v_14914;
wire v_14915;
wire v_14916;
wire v_14917;
wire v_14918;
wire v_14919;
wire v_14920;
wire v_14921;
wire v_14922;
wire v_14923;
wire v_14924;
wire v_14925;
wire v_14926;
wire v_14927;
wire v_14928;
wire v_14929;
wire v_14930;
wire v_14931;
wire v_14932;
wire v_14933;
wire v_14934;
wire v_14935;
wire v_14936;
wire v_14937;
wire v_14938;
wire v_14939;
wire v_14940;
wire v_14941;
wire v_14943;
wire v_14944;
wire v_14945;
wire v_14946;
wire v_14947;
wire v_14948;
wire v_14949;
wire v_14950;
wire v_14951;
wire v_14952;
wire v_14953;
wire v_14954;
wire v_14955;
wire v_14956;
wire v_14957;
wire v_14958;
wire v_14959;
wire v_14960;
wire v_14961;
wire v_14962;
wire v_14963;
wire v_14964;
wire v_14965;
wire v_14966;
wire v_14967;
wire v_14968;
wire v_14969;
wire v_14970;
wire v_14971;
wire v_14972;
wire v_14973;
wire v_14974;
wire v_14975;
wire v_14976;
wire v_14977;
wire v_14978;
wire v_14979;
wire v_14980;
wire v_14981;
wire v_14982;
wire v_14983;
wire v_14984;
wire v_14985;
wire v_14986;
wire v_14987;
wire v_14988;
wire v_14989;
wire v_14990;
wire v_14991;
wire v_14992;
wire v_14993;
wire v_14994;
wire v_14995;
wire v_14996;
wire v_14997;
wire v_14998;
wire v_14999;
wire v_15000;
wire v_15001;
wire v_15002;
wire v_15003;
wire v_15004;
wire v_15005;
wire v_15006;
wire v_15007;
wire v_15008;
wire v_15009;
wire v_15010;
wire v_15011;
wire v_15012;
wire v_15013;
wire v_15014;
wire v_15015;
wire v_15016;
wire v_15017;
wire v_15018;
wire v_15019;
wire v_15020;
wire v_15021;
wire v_15022;
wire v_15023;
wire v_15024;
wire v_15025;
wire v_15026;
wire v_15027;
wire v_15028;
wire v_15029;
wire v_15030;
wire v_15031;
wire v_15032;
wire v_15033;
wire v_15034;
wire v_15035;
wire v_15036;
wire v_15037;
wire v_15038;
wire v_15039;
wire v_15040;
wire v_15041;
wire v_15042;
wire v_15043;
wire v_15044;
wire v_15045;
wire v_15046;
wire v_15047;
wire v_15048;
wire v_15049;
wire v_15050;
wire v_15051;
wire v_15052;
wire v_15053;
wire v_15054;
wire v_15055;
wire v_15056;
wire v_15057;
wire v_15058;
wire v_15059;
wire v_15060;
wire v_15061;
wire v_15062;
wire v_15063;
wire v_15064;
wire v_15065;
wire v_15066;
wire v_15067;
wire v_15068;
wire v_15069;
wire v_15070;
wire v_15071;
wire v_15072;
wire v_15073;
wire v_15074;
wire v_15075;
wire v_15076;
wire v_15077;
wire v_15078;
wire v_15079;
wire v_15080;
wire v_15081;
wire v_15082;
wire v_15083;
wire v_15084;
wire v_15085;
wire v_15086;
wire v_15087;
wire v_15088;
wire v_15089;
wire v_15090;
wire v_15091;
wire v_15092;
wire v_15093;
wire v_15094;
wire v_15095;
wire v_15096;
wire v_15097;
wire v_15098;
wire v_15099;
wire v_15100;
wire v_15101;
wire v_15102;
wire v_15103;
wire v_15104;
wire v_15105;
wire v_15106;
wire v_15107;
wire v_15108;
wire v_15109;
wire v_15110;
wire v_15111;
wire v_15112;
wire v_15113;
wire v_15114;
wire v_15115;
wire v_15116;
wire v_15117;
wire v_15118;
wire v_15119;
wire v_15120;
wire v_15121;
wire v_15122;
wire v_15123;
wire v_15124;
wire v_15125;
wire v_15126;
wire v_15127;
wire v_15128;
wire v_15129;
wire v_15130;
wire v_15131;
wire v_15132;
wire v_15133;
wire v_15134;
wire v_15135;
wire v_15136;
wire v_15137;
wire v_15138;
wire v_15139;
wire v_15140;
wire v_15141;
wire v_15142;
wire v_15143;
wire v_15144;
wire v_15145;
wire v_15146;
wire v_15147;
wire v_15148;
wire v_15149;
wire v_15150;
wire v_15151;
wire v_15152;
wire v_15153;
wire v_15154;
wire v_15155;
wire v_15156;
wire v_15157;
wire v_15158;
wire v_15159;
wire v_15160;
wire v_15161;
wire v_15162;
wire v_15163;
wire v_15164;
wire v_15165;
wire v_15166;
wire v_15167;
wire v_15168;
wire v_15169;
wire v_15170;
wire v_15171;
wire v_15172;
wire v_15173;
wire v_15174;
wire v_15175;
wire v_15176;
wire v_15177;
wire v_15178;
wire v_15179;
wire v_15180;
wire v_15181;
wire v_15182;
wire v_15183;
wire v_15184;
wire v_15186;
wire v_15187;
wire v_15188;
wire v_15189;
wire v_15190;
wire v_15191;
wire v_15192;
wire v_15193;
wire v_15194;
wire v_15195;
wire v_15196;
wire v_15197;
wire v_15198;
wire v_15199;
wire v_15200;
wire v_15201;
wire v_15202;
wire v_15203;
wire v_15204;
wire v_15205;
wire v_15206;
wire v_15207;
wire v_15208;
wire v_15209;
wire v_15210;
wire v_15211;
wire v_15212;
wire v_15213;
wire v_15214;
wire v_15215;
wire v_15216;
wire v_15217;
wire v_15218;
wire v_15219;
wire v_15220;
wire v_15221;
wire v_15222;
wire v_15223;
wire v_15224;
wire v_15225;
wire v_15226;
wire v_15227;
wire v_15228;
wire v_15229;
wire v_15230;
wire v_15231;
wire v_15232;
wire v_15233;
wire v_15234;
wire v_15235;
wire v_15236;
wire v_15237;
wire v_15238;
wire v_15239;
wire v_15240;
wire v_15241;
wire v_15242;
wire v_15243;
wire v_15244;
wire v_15245;
wire v_15246;
wire v_15247;
wire v_15248;
wire v_15249;
wire v_15250;
wire v_15251;
wire v_15252;
wire v_15253;
wire v_15254;
wire v_15255;
wire v_15256;
wire v_15257;
wire v_15258;
wire v_15259;
wire v_15260;
wire v_15261;
wire v_15262;
wire v_15263;
wire v_15264;
wire v_15265;
wire v_15266;
wire v_15267;
wire v_15268;
wire v_15269;
wire v_15270;
wire v_15271;
wire v_15272;
wire v_15273;
wire v_15274;
wire v_15275;
wire v_15276;
wire v_15277;
wire v_15278;
wire v_15279;
wire v_15280;
wire v_15281;
wire v_15282;
wire v_15283;
wire v_15284;
wire v_15285;
wire v_15286;
wire v_15287;
wire v_15288;
wire v_15289;
wire v_15290;
wire v_15291;
wire v_15292;
wire v_15293;
wire v_15294;
wire v_15295;
wire v_15296;
wire v_15297;
wire v_15298;
wire v_15299;
wire v_15300;
wire v_15301;
wire v_15302;
wire v_15303;
wire v_15304;
wire v_15305;
wire v_15306;
wire v_15307;
wire v_15308;
wire v_15309;
wire v_15310;
wire v_15311;
wire v_15312;
wire v_15313;
wire v_15314;
wire v_15315;
wire v_15316;
wire v_15317;
wire v_15318;
wire v_15319;
wire v_15320;
wire v_15321;
wire v_15322;
wire v_15323;
wire v_15324;
wire v_15325;
wire v_15326;
wire v_15327;
wire v_15328;
wire v_15329;
wire v_15330;
wire v_15331;
wire v_15332;
wire v_15333;
wire v_15334;
wire v_15335;
wire v_15336;
wire v_15337;
wire v_15338;
wire v_15339;
wire v_15340;
wire v_15341;
wire v_15342;
wire v_15343;
wire v_15344;
wire v_15345;
wire v_15346;
wire v_15347;
wire v_15348;
wire v_15349;
wire v_15350;
wire v_15351;
wire v_15352;
wire v_15353;
wire v_15354;
wire v_15355;
wire v_15356;
wire v_15357;
wire v_15358;
wire v_15359;
wire v_15360;
wire v_15361;
wire v_15362;
wire v_15363;
wire v_15364;
wire v_15365;
wire v_15366;
wire v_15367;
wire v_15368;
wire v_15369;
wire v_15370;
wire v_15371;
wire v_15372;
wire v_15373;
wire v_15374;
wire v_15375;
wire v_15376;
wire v_15377;
wire v_15378;
wire v_15379;
wire v_15380;
wire v_15381;
wire v_15382;
wire v_15383;
wire v_15384;
wire v_15385;
wire v_15386;
wire v_15387;
wire v_15388;
wire v_15389;
wire v_15390;
wire v_15391;
wire v_15392;
wire v_15393;
wire v_15394;
wire v_15395;
wire v_15396;
wire v_15397;
wire v_15398;
wire v_15399;
wire v_15400;
wire v_15401;
wire v_15402;
wire v_15403;
wire v_15404;
wire v_15405;
wire v_15406;
wire v_15407;
wire v_15408;
wire v_15409;
wire v_15410;
wire v_15411;
wire v_15412;
wire v_15413;
wire v_15414;
wire v_15415;
wire v_15416;
wire v_15417;
wire v_15418;
wire v_15419;
wire v_15420;
wire v_15421;
wire v_15422;
wire v_15423;
wire v_15424;
wire v_15425;
wire v_15426;
wire v_15427;
wire v_15429;
wire v_15430;
wire v_15431;
wire v_15432;
wire v_15433;
wire v_15434;
wire v_15435;
wire v_15436;
wire v_15437;
wire v_15438;
wire v_15439;
wire v_15440;
wire v_15441;
wire v_15442;
wire v_15443;
wire v_15444;
wire v_15445;
wire v_15446;
wire v_15447;
wire v_15448;
wire v_15449;
wire v_15450;
wire v_15451;
wire v_15452;
wire v_15453;
wire v_15454;
wire v_15455;
wire v_15456;
wire v_15457;
wire v_15458;
wire v_15459;
wire v_15460;
wire v_15461;
wire v_15462;
wire v_15463;
wire v_15464;
wire v_15465;
wire v_15466;
wire v_15467;
wire v_15468;
wire v_15469;
wire v_15470;
wire v_15471;
wire v_15472;
wire v_15473;
wire v_15474;
wire v_15475;
wire v_15476;
wire v_15477;
wire v_15478;
wire v_15479;
wire v_15480;
wire v_15481;
wire v_15482;
wire v_15483;
wire v_15484;
wire v_15485;
wire v_15486;
wire v_15487;
wire v_15488;
wire v_15489;
wire v_15490;
wire v_15491;
wire v_15492;
wire v_15493;
wire v_15494;
wire v_15495;
wire v_15496;
wire v_15497;
wire v_15498;
wire v_15499;
wire v_15500;
wire v_15501;
wire v_15502;
wire v_15503;
wire v_15504;
wire v_15505;
wire v_15506;
wire v_15507;
wire v_15508;
wire v_15509;
wire v_15510;
wire v_15511;
wire v_15512;
wire v_15513;
wire v_15514;
wire v_15515;
wire v_15516;
wire v_15517;
wire v_15518;
wire v_15519;
wire v_15520;
wire v_15521;
wire v_15522;
wire v_15523;
wire v_15524;
wire v_15525;
wire v_15526;
wire v_15527;
wire v_15528;
wire v_15529;
wire v_15530;
wire v_15531;
wire v_15532;
wire v_15533;
wire v_15534;
wire v_15535;
wire v_15536;
wire v_15537;
wire v_15538;
wire v_15539;
wire v_15540;
wire v_15541;
wire v_15542;
wire v_15543;
wire v_15544;
wire v_15545;
wire v_15546;
wire v_15547;
wire v_15548;
wire v_15549;
wire v_15550;
wire v_15551;
wire v_15552;
wire v_15553;
wire v_15554;
wire v_15555;
wire v_15556;
wire v_15557;
wire v_15558;
wire v_15559;
wire v_15560;
wire v_15561;
wire v_15562;
wire v_15563;
wire v_15564;
wire v_15565;
wire v_15566;
wire v_15567;
wire v_15568;
wire v_15569;
wire v_15570;
wire v_15571;
wire v_15572;
wire v_15573;
wire v_15574;
wire v_15575;
wire v_15576;
wire v_15577;
wire v_15578;
wire v_15579;
wire v_15580;
wire v_15581;
wire v_15582;
wire v_15583;
wire v_15584;
wire v_15585;
wire v_15586;
wire v_15587;
wire v_15588;
wire v_15589;
wire v_15590;
wire v_15591;
wire v_15592;
wire v_15593;
wire v_15594;
wire v_15595;
wire v_15596;
wire v_15597;
wire v_15598;
wire v_15599;
wire v_15600;
wire v_15601;
wire v_15602;
wire v_15603;
wire v_15604;
wire v_15605;
wire v_15606;
wire v_15607;
wire v_15608;
wire v_15609;
wire v_15610;
wire v_15611;
wire v_15612;
wire v_15613;
wire v_15614;
wire v_15615;
wire v_15616;
wire v_15617;
wire v_15618;
wire v_15619;
wire v_15620;
wire v_15621;
wire v_15622;
wire v_15623;
wire v_15624;
wire v_15625;
wire v_15626;
wire v_15627;
wire v_15628;
wire v_15629;
wire v_15630;
wire v_15631;
wire v_15632;
wire v_15633;
wire v_15634;
wire v_15635;
wire v_15636;
wire v_15637;
wire v_15638;
wire v_15639;
wire v_15640;
wire v_15641;
wire v_15642;
wire v_15643;
wire v_15644;
wire v_15645;
wire v_15646;
wire v_15647;
wire v_15648;
wire v_15649;
wire v_15650;
wire v_15651;
wire v_15652;
wire v_15653;
wire v_15654;
wire v_15655;
wire v_15656;
wire v_15657;
wire v_15658;
wire v_15659;
wire v_15660;
wire v_15661;
wire v_15662;
wire v_15663;
wire v_15664;
wire v_15665;
wire v_15666;
wire v_15667;
wire v_15668;
wire v_15669;
wire v_15670;
wire v_15672;
wire v_15673;
wire v_15674;
wire v_15675;
wire v_15676;
wire v_15677;
wire v_15678;
wire v_15679;
wire v_15680;
wire v_15681;
wire v_15682;
wire v_15683;
wire v_15684;
wire v_15685;
wire v_15686;
wire v_15687;
wire v_15688;
wire v_15689;
wire v_15690;
wire v_15691;
wire v_15692;
wire v_15693;
wire v_15694;
wire v_15695;
wire v_15696;
wire v_15697;
wire v_15698;
wire v_15699;
wire v_15700;
wire v_15701;
wire v_15702;
wire v_15703;
wire v_15704;
wire v_15705;
wire v_15706;
wire v_15707;
wire v_15708;
wire v_15709;
wire v_15710;
wire v_15711;
wire v_15712;
wire v_15713;
wire v_15714;
wire v_15715;
wire v_15716;
wire v_15717;
wire v_15718;
wire v_15719;
wire v_15720;
wire v_15721;
wire v_15722;
wire v_15723;
wire v_15724;
wire v_15725;
wire v_15726;
wire v_15727;
wire v_15728;
wire v_15729;
wire v_15730;
wire v_15731;
wire v_15732;
wire v_15733;
wire v_15734;
wire v_15735;
wire v_15736;
wire v_15737;
wire v_15738;
wire v_15739;
wire v_15740;
wire v_15741;
wire v_15742;
wire v_15743;
wire v_15744;
wire v_15745;
wire v_15746;
wire v_15747;
wire v_15748;
wire v_15749;
wire v_15750;
wire v_15751;
wire v_15752;
wire v_15753;
wire v_15754;
wire v_15755;
wire v_15756;
wire v_15757;
wire v_15758;
wire v_15759;
wire v_15760;
wire v_15761;
wire v_15762;
wire v_15763;
wire v_15764;
wire v_15765;
wire v_15766;
wire v_15767;
wire v_15768;
wire v_15769;
wire v_15770;
wire v_15771;
wire v_15772;
wire v_15773;
wire v_15774;
wire v_15775;
wire v_15776;
wire v_15777;
wire v_15778;
wire v_15779;
wire v_15780;
wire v_15781;
wire v_15782;
wire v_15783;
wire v_15784;
wire v_15785;
wire v_15786;
wire v_15787;
wire v_15788;
wire v_15789;
wire v_15790;
wire v_15791;
wire v_15792;
wire v_15793;
wire v_15794;
wire v_15795;
wire v_15796;
wire v_15797;
wire v_15798;
wire v_15799;
wire v_15800;
wire v_15801;
wire v_15802;
wire v_15803;
wire v_15804;
wire v_15805;
wire v_15806;
wire v_15807;
wire v_15808;
wire v_15809;
wire v_15810;
wire v_15811;
wire v_15812;
wire v_15813;
wire v_15814;
wire v_15815;
wire v_15816;
wire v_15817;
wire v_15818;
wire v_15819;
wire v_15820;
wire v_15821;
wire v_15822;
wire v_15823;
wire v_15824;
wire v_15825;
wire v_15826;
wire v_15827;
wire v_15828;
wire v_15829;
wire v_15830;
wire v_15831;
wire v_15832;
wire v_15833;
wire v_15834;
wire v_15835;
wire v_15836;
wire v_15837;
wire v_15838;
wire v_15839;
wire v_15840;
wire v_15841;
wire v_15842;
wire v_15843;
wire v_15844;
wire v_15845;
wire v_15846;
wire v_15847;
wire v_15848;
wire v_15849;
wire v_15850;
wire v_15851;
wire v_15852;
wire v_15853;
wire v_15854;
wire v_15855;
wire v_15856;
wire v_15857;
wire v_15858;
wire v_15859;
wire v_15860;
wire v_15861;
wire v_15862;
wire v_15863;
wire v_15864;
wire v_15865;
wire v_15866;
wire v_15867;
wire v_15868;
wire v_15869;
wire v_15870;
wire v_15871;
wire v_15872;
wire v_15873;
wire v_15874;
wire v_15875;
wire v_15876;
wire v_15877;
wire v_15878;
wire v_15879;
wire v_15880;
wire v_15881;
wire v_15882;
wire v_15883;
wire v_15884;
wire v_15885;
wire v_15886;
wire v_15887;
wire v_15888;
wire v_15889;
wire v_15890;
wire v_15891;
wire v_15892;
wire v_15893;
wire v_15894;
wire v_15895;
wire v_15896;
wire v_15897;
wire v_15898;
wire v_15899;
wire v_15900;
wire v_15901;
wire v_15902;
wire v_15903;
wire v_15904;
wire v_15905;
wire v_15906;
wire v_15907;
wire v_15908;
wire v_15909;
wire v_15910;
wire v_15911;
wire v_15912;
wire v_15913;
wire v_15915;
wire v_15916;
wire v_15917;
wire v_15918;
wire v_15919;
wire v_15920;
wire v_15921;
wire v_15922;
wire v_15923;
wire v_15924;
wire v_15925;
wire v_15926;
wire v_15927;
wire v_15928;
wire v_15929;
wire v_15930;
wire v_15931;
wire v_15932;
wire v_15933;
wire v_15934;
wire v_15935;
wire v_15936;
wire v_15937;
wire v_15938;
wire v_15939;
wire v_15940;
wire v_15941;
wire v_15942;
wire v_15943;
wire v_15944;
wire v_15945;
wire v_15946;
wire v_15947;
wire v_15948;
wire v_15949;
wire v_15950;
wire v_15951;
wire v_15952;
wire v_15953;
wire v_15954;
wire v_15955;
wire v_15956;
wire v_15957;
wire v_15958;
wire v_15959;
wire v_15960;
wire v_15961;
wire v_15962;
wire v_15963;
wire v_15964;
wire v_15965;
wire v_15966;
wire v_15967;
wire v_15968;
wire v_15969;
wire v_15970;
wire v_15971;
wire v_15972;
wire v_15973;
wire v_15974;
wire v_15975;
wire v_15976;
wire v_15977;
wire v_15978;
wire v_15979;
wire v_15980;
wire v_15981;
wire v_15982;
wire v_15983;
wire v_15984;
wire v_15985;
wire v_15986;
wire v_15987;
wire v_15988;
wire v_15989;
wire v_15990;
wire v_15991;
wire v_15992;
wire v_15993;
wire v_15994;
wire v_15995;
wire v_15996;
wire v_15997;
wire v_15998;
wire v_15999;
wire v_16000;
wire v_16001;
wire v_16002;
wire v_16003;
wire v_16004;
wire v_16005;
wire v_16006;
wire v_16007;
wire v_16008;
wire v_16009;
wire v_16010;
wire v_16011;
wire v_16012;
wire v_16013;
wire v_16014;
wire v_16015;
wire v_16016;
wire v_16017;
wire v_16018;
wire v_16019;
wire v_16020;
wire v_16021;
wire v_16022;
wire v_16023;
wire v_16024;
wire v_16025;
wire v_16026;
wire v_16027;
wire v_16028;
wire v_16029;
wire v_16030;
wire v_16031;
wire v_16032;
wire v_16033;
wire v_16034;
wire v_16035;
wire v_16036;
wire v_16037;
wire v_16038;
wire v_16039;
wire v_16040;
wire v_16041;
wire v_16042;
wire v_16043;
wire v_16044;
wire v_16045;
wire v_16046;
wire v_16047;
wire v_16048;
wire v_16049;
wire v_16050;
wire v_16051;
wire v_16052;
wire v_16053;
wire v_16054;
wire v_16055;
wire v_16056;
wire v_16057;
wire v_16058;
wire v_16059;
wire v_16060;
wire v_16061;
wire v_16062;
wire v_16063;
wire v_16064;
wire v_16065;
wire v_16066;
wire v_16067;
wire v_16068;
wire v_16069;
wire v_16070;
wire v_16071;
wire v_16072;
wire v_16073;
wire v_16074;
wire v_16075;
wire v_16076;
wire v_16077;
wire v_16078;
wire v_16079;
wire v_16080;
wire v_16081;
wire v_16082;
wire v_16083;
wire v_16084;
wire v_16085;
wire v_16086;
wire v_16087;
wire v_16088;
wire v_16089;
wire v_16090;
wire v_16091;
wire v_16092;
wire v_16093;
wire v_16094;
wire v_16095;
wire v_16096;
wire v_16097;
wire v_16098;
wire v_16099;
wire v_16100;
wire v_16101;
wire v_16102;
wire v_16103;
wire v_16104;
wire v_16105;
wire v_16106;
wire v_16107;
wire v_16108;
wire v_16109;
wire v_16110;
wire v_16111;
wire v_16112;
wire v_16113;
wire v_16114;
wire v_16115;
wire v_16116;
wire v_16117;
wire v_16118;
wire v_16119;
wire v_16120;
wire v_16121;
wire v_16122;
wire v_16123;
wire v_16124;
wire v_16125;
wire v_16126;
wire v_16127;
wire v_16128;
wire v_16129;
wire v_16130;
wire v_16131;
wire v_16132;
wire v_16133;
wire v_16134;
wire v_16135;
wire v_16136;
wire v_16137;
wire v_16138;
wire v_16139;
wire v_16140;
wire v_16141;
wire v_16142;
wire v_16143;
wire v_16144;
wire v_16145;
wire v_16146;
wire v_16147;
wire v_16148;
wire v_16149;
wire v_16150;
wire v_16151;
wire v_16152;
wire v_16153;
wire v_16154;
wire v_16155;
wire v_16156;
wire v_16158;
wire v_16159;
wire v_16160;
wire v_16161;
wire v_16162;
wire v_16163;
wire v_16164;
wire v_16165;
wire v_16166;
wire v_16167;
wire v_16168;
wire v_16169;
wire v_16170;
wire v_16171;
wire v_16172;
wire v_16173;
wire v_16174;
wire v_16175;
wire v_16176;
wire v_16177;
wire v_16178;
wire v_16179;
wire v_16180;
wire v_16181;
wire v_16182;
wire v_16183;
wire v_16184;
wire v_16185;
wire v_16186;
wire v_16187;
wire v_16188;
wire v_16189;
wire v_16190;
wire v_16191;
wire v_16192;
wire v_16193;
wire v_16194;
wire v_16195;
wire v_16196;
wire v_16197;
wire v_16198;
wire v_16199;
wire v_16200;
wire v_16201;
wire v_16202;
wire v_16203;
wire v_16204;
wire v_16205;
wire v_16206;
wire v_16207;
wire v_16208;
wire v_16209;
wire v_16210;
wire v_16211;
wire v_16212;
wire v_16213;
wire v_16214;
wire v_16215;
wire v_16216;
wire v_16217;
wire v_16218;
wire v_16219;
wire v_16220;
wire v_16221;
wire v_16222;
wire v_16223;
wire v_16224;
wire v_16225;
wire v_16226;
wire v_16227;
wire v_16228;
wire v_16229;
wire v_16230;
wire v_16231;
wire v_16232;
wire v_16233;
wire v_16234;
wire v_16235;
wire v_16236;
wire v_16237;
wire v_16238;
wire v_16239;
wire v_16240;
wire v_16241;
wire v_16242;
wire v_16243;
wire v_16244;
wire v_16245;
wire v_16246;
wire v_16247;
wire v_16248;
wire v_16249;
wire v_16250;
wire v_16251;
wire v_16252;
wire v_16253;
wire v_16254;
wire v_16255;
wire v_16256;
wire v_16257;
wire v_16258;
wire v_16259;
wire v_16260;
wire v_16261;
wire v_16262;
wire v_16263;
wire v_16264;
wire v_16265;
wire v_16266;
wire v_16267;
wire v_16268;
wire v_16269;
wire v_16270;
wire v_16271;
wire v_16272;
wire v_16273;
wire v_16274;
wire v_16275;
wire v_16276;
wire v_16277;
wire v_16278;
wire v_16279;
wire v_16280;
wire v_16281;
wire v_16282;
wire v_16283;
wire v_16284;
wire v_16285;
wire v_16286;
wire v_16287;
wire v_16288;
wire v_16289;
wire v_16290;
wire v_16291;
wire v_16292;
wire v_16293;
wire v_16294;
wire v_16295;
wire v_16296;
wire v_16297;
wire v_16298;
wire v_16299;
wire v_16300;
wire v_16301;
wire v_16302;
wire v_16303;
wire v_16304;
wire v_16305;
wire v_16306;
wire v_16307;
wire v_16308;
wire v_16309;
wire v_16310;
wire v_16311;
wire v_16312;
wire v_16313;
wire v_16314;
wire v_16315;
wire v_16316;
wire v_16317;
wire v_16318;
wire v_16319;
wire v_16320;
wire v_16321;
wire v_16322;
wire v_16323;
wire v_16324;
wire v_16325;
wire v_16326;
wire v_16327;
wire v_16328;
wire v_16329;
wire v_16330;
wire v_16331;
wire v_16332;
wire v_16333;
wire v_16334;
wire v_16335;
wire v_16336;
wire v_16337;
wire v_16338;
wire v_16339;
wire v_16340;
wire v_16341;
wire v_16342;
wire v_16343;
wire v_16344;
wire v_16345;
wire v_16346;
wire v_16347;
wire v_16348;
wire v_16349;
wire v_16350;
wire v_16351;
wire v_16352;
wire v_16353;
wire v_16354;
wire v_16355;
wire v_16356;
wire v_16357;
wire v_16358;
wire v_16359;
wire v_16360;
wire v_16361;
wire v_16362;
wire v_16363;
wire v_16364;
wire v_16365;
wire v_16366;
wire v_16367;
wire v_16368;
wire v_16369;
wire v_16370;
wire v_16371;
wire v_16372;
wire v_16373;
wire v_16374;
wire v_16375;
wire v_16376;
wire v_16377;
wire v_16378;
wire v_16379;
wire v_16380;
wire v_16381;
wire v_16382;
wire v_16383;
wire v_16384;
wire v_16385;
wire v_16386;
wire v_16387;
wire v_16388;
wire v_16389;
wire v_16390;
wire v_16391;
wire v_16392;
wire v_16393;
wire v_16394;
wire v_16395;
wire v_16396;
wire v_16397;
wire v_16398;
wire v_16399;
wire v_16401;
wire v_16402;
wire v_16403;
wire v_16404;
wire v_16405;
wire v_16406;
wire v_16407;
wire v_16408;
wire v_16409;
wire v_16410;
wire v_16411;
wire v_16412;
wire v_16413;
wire v_16414;
wire v_16415;
wire v_16416;
wire v_16417;
wire v_16418;
wire v_16419;
wire v_16420;
wire v_16421;
wire v_16422;
wire v_16423;
wire v_16424;
wire v_16425;
wire v_16426;
wire v_16427;
wire v_16428;
wire v_16429;
wire v_16430;
wire v_16431;
wire v_16432;
wire v_16433;
wire v_16434;
wire v_16435;
wire v_16436;
wire v_16437;
wire v_16438;
wire v_16439;
wire v_16440;
wire v_16441;
wire v_16442;
wire v_16443;
wire v_16444;
wire v_16445;
wire v_16446;
wire v_16447;
wire v_16448;
wire v_16449;
wire v_16450;
wire v_16451;
wire v_16452;
wire v_16453;
wire v_16454;
wire v_16455;
wire v_16456;
wire v_16457;
wire v_16458;
wire v_16459;
wire v_16460;
wire v_16461;
wire v_16462;
wire v_16463;
wire v_16464;
wire v_16465;
wire v_16466;
wire v_16467;
wire v_16468;
wire v_16469;
wire v_16470;
wire v_16471;
wire v_16472;
wire v_16473;
wire v_16474;
wire v_16475;
wire v_16476;
wire v_16477;
wire v_16478;
wire v_16479;
wire v_16480;
wire v_16481;
wire v_16482;
wire v_16483;
wire v_16484;
wire v_16485;
wire v_16486;
wire v_16487;
wire v_16488;
wire v_16489;
wire v_16490;
wire v_16491;
wire v_16492;
wire v_16493;
wire v_16494;
wire v_16495;
wire v_16496;
wire v_16497;
wire v_16498;
wire v_16499;
wire v_16500;
wire v_16501;
wire v_16502;
wire v_16503;
wire v_16504;
wire v_16505;
wire v_16506;
wire v_16507;
wire v_16508;
wire v_16509;
wire v_16510;
wire v_16511;
wire v_16512;
wire v_16513;
wire v_16514;
wire v_16515;
wire v_16516;
wire v_16517;
wire v_16518;
wire v_16519;
wire v_16520;
wire v_16521;
wire v_16522;
wire v_16523;
wire v_16524;
wire v_16525;
wire v_16526;
wire v_16527;
wire v_16528;
wire v_16529;
wire v_16530;
wire v_16531;
wire v_16532;
wire v_16533;
wire v_16534;
wire v_16535;
wire v_16536;
wire v_16537;
wire v_16538;
wire v_16539;
wire v_16540;
wire v_16541;
wire v_16542;
wire v_16543;
wire v_16544;
wire v_16545;
wire v_16546;
wire v_16547;
wire v_16548;
wire v_16549;
wire v_16550;
wire v_16551;
wire v_16552;
wire v_16553;
wire v_16554;
wire v_16555;
wire v_16556;
wire v_16557;
wire v_16558;
wire v_16559;
wire v_16560;
wire v_16561;
wire v_16562;
wire v_16563;
wire v_16564;
wire v_16565;
wire v_16566;
wire v_16567;
wire v_16568;
wire v_16569;
wire v_16570;
wire v_16571;
wire v_16572;
wire v_16573;
wire v_16574;
wire v_16575;
wire v_16576;
wire v_16577;
wire v_16578;
wire v_16579;
wire v_16580;
wire v_16581;
wire v_16582;
wire v_16583;
wire v_16584;
wire v_16585;
wire v_16586;
wire v_16587;
wire v_16588;
wire v_16589;
wire v_16590;
wire v_16591;
wire v_16592;
wire v_16593;
wire v_16594;
wire v_16595;
wire v_16596;
wire v_16597;
wire v_16598;
wire v_16599;
wire v_16600;
wire v_16601;
wire v_16602;
wire v_16603;
wire v_16604;
wire v_16605;
wire v_16606;
wire v_16607;
wire v_16608;
wire v_16609;
wire v_16610;
wire v_16611;
wire v_16612;
wire v_16613;
wire v_16614;
wire v_16615;
wire v_16616;
wire v_16617;
wire v_16618;
wire v_16619;
wire v_16620;
wire v_16621;
wire v_16622;
wire v_16623;
wire v_16624;
wire v_16625;
wire v_16626;
wire v_16627;
wire v_16628;
wire v_16629;
wire v_16630;
wire v_16631;
wire v_16632;
wire v_16633;
wire v_16634;
wire v_16635;
wire v_16636;
wire v_16637;
wire v_16638;
wire v_16639;
wire v_16640;
wire v_16641;
wire v_16642;
wire v_16643;
wire v_16644;
wire v_16645;
wire v_16646;
wire v_16647;
wire v_16648;
wire v_16649;
wire v_16650;
wire v_16651;
wire v_16652;
wire v_16653;
wire v_16654;
wire v_16655;
wire v_16656;
wire v_16657;
wire v_16658;
wire v_16659;
wire v_16660;
wire v_16661;
wire v_16662;
wire v_16663;
wire v_16664;
wire v_16665;
wire v_16666;
wire v_16667;
wire v_16668;
wire v_16669;
wire v_16670;
wire v_16671;
wire v_16672;
wire v_16673;
wire v_16674;
wire v_16675;
wire v_16676;
wire v_16677;
wire v_16678;
wire v_16679;
wire v_16680;
wire v_16681;
wire v_16682;
wire v_16683;
wire v_16684;
wire v_16685;
wire v_16686;
wire v_16687;
wire v_16688;
wire v_16689;
wire v_16690;
wire v_16691;
wire v_16692;
wire v_16693;
wire v_16694;
wire v_16695;
wire v_16696;
wire v_16697;
wire v_16698;
wire v_16699;
wire v_16700;
wire v_16701;
wire v_16702;
wire v_16703;
wire v_16704;
wire v_16705;
wire v_16706;
wire v_16707;
wire v_16708;
wire v_16709;
wire v_16710;
wire v_16711;
wire v_16712;
wire v_16713;
wire v_16714;
wire v_16715;
wire v_16716;
wire v_16717;
wire v_16718;
wire v_16719;
wire v_16720;
wire v_16721;
wire v_16722;
wire v_16723;
wire v_16724;
wire v_16725;
wire v_16726;
wire v_16727;
wire v_16728;
wire v_16729;
wire v_16730;
wire v_16731;
wire v_16732;
wire v_16733;
wire v_16734;
wire v_16735;
wire v_16736;
wire v_16737;
wire v_16738;
wire v_16739;
wire v_16740;
wire v_16741;
wire v_16742;
wire v_16743;
wire v_16744;
wire v_16745;
wire v_16746;
wire v_16747;
wire v_16748;
wire v_16749;
wire v_16750;
wire v_16751;
wire v_16752;
wire v_16753;
wire v_16754;
wire v_16755;
wire v_16756;
wire v_16757;
wire v_16758;
wire v_16759;
wire v_16760;
wire v_16761;
wire v_16762;
wire v_16763;
wire v_16764;
wire v_16765;
wire v_16766;
wire v_16767;
wire v_16768;
wire v_16769;
wire v_16770;
wire v_16771;
wire v_16772;
wire v_16773;
wire v_16774;
wire v_16775;
wire v_16776;
wire v_16777;
wire v_16778;
wire v_16779;
wire v_16780;
wire v_16781;
wire v_16782;
wire v_16783;
wire v_16784;
wire v_16785;
wire v_16786;
wire v_16787;
wire v_16788;
wire v_16789;
wire v_16790;
wire v_16791;
wire v_16793;
wire v_16794;
wire v_16795;
wire v_16796;
wire v_16797;
wire v_16798;
wire v_16799;
wire v_16800;
wire v_16801;
wire v_16802;
wire v_16803;
wire v_16804;
wire v_16805;
wire v_16806;
wire v_16807;
wire v_16808;
wire v_16809;
wire v_16810;
wire v_16811;
wire v_16812;
wire v_16813;
wire v_16814;
wire v_16815;
wire v_16816;
wire v_16817;
wire v_16818;
wire v_16819;
wire v_16820;
wire v_16821;
wire v_16822;
wire v_16823;
wire v_16824;
wire v_16825;
wire v_16826;
wire v_16827;
wire v_16828;
wire v_16829;
wire v_16830;
wire v_16831;
wire v_16832;
wire v_16833;
wire v_16834;
wire v_16835;
wire v_16836;
wire v_16837;
wire v_16838;
wire v_16839;
wire v_16840;
wire v_16841;
wire v_16842;
wire v_16843;
wire v_16844;
wire v_16845;
wire v_16846;
wire v_16847;
wire v_16848;
wire v_16849;
wire v_16850;
wire v_16851;
wire v_16852;
wire v_16853;
wire v_16854;
wire v_16855;
wire v_16856;
wire v_16857;
wire v_16858;
wire v_16859;
wire v_16860;
wire v_16861;
wire v_16862;
wire v_16863;
wire v_16864;
wire v_16865;
wire v_16866;
wire v_16867;
wire v_16868;
wire v_16869;
wire v_16870;
wire v_16871;
wire v_16872;
wire v_16873;
wire v_16874;
wire v_16875;
wire v_16876;
wire v_16877;
wire v_16878;
wire v_16879;
wire v_16880;
wire v_16881;
wire v_16882;
wire v_16883;
wire v_16884;
wire v_16885;
wire v_16887;
wire v_16889;
wire v_16890;
wire v_16891;
wire v_16893;
wire v_16894;
wire v_16895;
wire v_16897;
wire v_16898;
wire v_16899;
wire v_16901;
wire v_16902;
wire v_16904;
wire v_16905;
wire v_16906;
wire v_16908;
wire v_16909;
wire v_16910;
wire v_16912;
wire v_16913;
wire v_16914;
wire v_16916;
wire v_16917;
wire v_16918;
wire v_16920;
wire v_16921;
wire v_16922;
wire v_16924;
wire v_16925;
wire v_16926;
wire v_16928;
wire v_16929;
wire v_16930;
wire v_16932;
wire v_16933;
wire v_16934;
wire v_16936;
wire v_16937;
wire v_16938;
wire v_16940;
wire v_16941;
wire v_16942;
wire v_16944;
wire v_16945;
wire v_16946;
wire v_16948;
wire v_16949;
wire v_16950;
wire v_16952;
wire v_16953;
wire v_16954;
wire v_16955;
wire v_16956;
wire v_16957;
wire v_16958;
wire v_16959;
wire v_16960;
wire v_16961;
wire v_16962;
wire v_16963;
wire v_16964;
wire v_16965;
wire v_16966;
wire v_16967;
wire v_16968;
wire v_16969;
wire v_16970;
wire v_16971;
wire v_16972;
wire v_16973;
wire v_16974;
wire v_16975;
wire v_16976;
wire v_16977;
wire v_16978;
wire v_16979;
wire v_16980;
wire v_16981;
wire v_16982;
wire v_16983;
wire v_16984;
wire v_16985;
wire v_16986;
wire v_16987;
wire v_16988;
wire v_16989;
wire v_16990;
wire v_16991;
wire v_16992;
wire v_16993;
wire v_16994;
wire v_16995;
wire v_16996;
wire v_16997;
wire v_16998;
wire v_16999;
wire v_17000;
wire v_17001;
wire v_17002;
wire v_17003;
wire v_17004;
wire v_17005;
wire v_17006;
wire v_17007;
wire v_17008;
wire v_17009;
wire v_17010;
wire v_17011;
wire v_17012;
wire v_17013;
wire v_17014;
wire v_17015;
wire v_17016;
wire v_17017;
wire v_17018;
wire v_17019;
wire v_17020;
wire v_17021;
wire v_17022;
wire v_17023;
wire v_17024;
wire v_17025;
wire v_17026;
wire v_17027;
wire v_17028;
wire v_17029;
wire v_17030;
wire v_17031;
wire v_17032;
wire v_17033;
wire v_17034;
wire v_17035;
wire v_17036;
wire v_17037;
wire v_17038;
wire v_17039;
wire v_17040;
wire v_17041;
wire v_17042;
wire v_17043;
wire v_17044;
wire v_17045;
wire v_17046;
wire v_17047;
wire v_17048;
wire v_17049;
wire v_17050;
wire v_17051;
wire v_17052;
wire v_17053;
wire v_17054;
wire v_17055;
wire v_17056;
wire v_17057;
wire v_17058;
wire v_17059;
wire v_17060;
wire v_17061;
wire v_17062;
wire v_17063;
wire v_17064;
wire v_17065;
wire v_17066;
wire v_17067;
wire v_17068;
wire v_17069;
wire v_17070;
wire v_17071;
wire v_17072;
wire v_17073;
wire v_17074;
wire v_17075;
wire v_17076;
wire v_17077;
wire v_17078;
wire v_17079;
wire v_17080;
wire v_17081;
wire v_17082;
wire v_17083;
wire v_17084;
wire v_17085;
wire v_17086;
wire v_17087;
wire v_17088;
wire v_17089;
wire v_17090;
wire v_17091;
wire v_17092;
wire v_17093;
wire v_17094;
wire v_17095;
wire v_17096;
wire v_17097;
wire v_17098;
wire v_17099;
wire v_17100;
wire v_17101;
wire v_17102;
wire v_17103;
wire v_17104;
wire v_17105;
wire v_17106;
wire v_17107;
wire v_17108;
wire v_17109;
wire v_17110;
wire v_17111;
wire v_17112;
wire v_17113;
wire v_17114;
wire v_17115;
wire v_17116;
wire v_17117;
wire v_17118;
wire v_17119;
wire v_17120;
wire v_17121;
wire v_17122;
wire v_17123;
wire v_17124;
wire v_17125;
wire v_17126;
wire v_17127;
wire v_17128;
wire v_17129;
wire v_17130;
wire v_17131;
wire v_17132;
wire v_17133;
wire v_17134;
wire v_17135;
wire v_17136;
wire v_17137;
wire v_17138;
wire v_17139;
wire v_17140;
wire v_17141;
wire v_17142;
wire v_17143;
wire v_17144;
wire v_17145;
wire v_17147;
wire v_17148;
wire v_17149;
wire v_17150;
wire v_17151;
wire v_17152;
wire v_17153;
wire v_17154;
wire v_17155;
wire v_17156;
wire v_17157;
wire v_17158;
wire v_17159;
wire v_17160;
wire v_17161;
wire v_17162;
wire v_17163;
wire v_17164;
wire v_17165;
wire v_17166;
wire v_17167;
wire v_17168;
wire v_17169;
wire v_17170;
wire v_17171;
wire v_17172;
wire v_17173;
wire v_17174;
wire v_17175;
wire v_17176;
wire v_17177;
wire v_17178;
wire v_17179;
wire v_17180;
wire v_17181;
wire v_17182;
wire v_17183;
wire v_17184;
wire v_17185;
wire v_17186;
wire v_17187;
wire v_17188;
wire v_17189;
wire v_17190;
wire v_17191;
wire v_17192;
wire v_17193;
wire v_17194;
wire v_17195;
wire v_17196;
wire v_17197;
wire v_17198;
wire v_17199;
wire v_17200;
wire v_17201;
wire v_17202;
wire v_17203;
wire v_17204;
wire v_17205;
wire v_17206;
wire v_17207;
wire v_17208;
wire v_17209;
wire v_17210;
wire v_17211;
wire v_17212;
wire v_17213;
wire v_17214;
wire v_17215;
wire v_17216;
wire v_17217;
wire v_17218;
wire v_17219;
wire v_17220;
wire v_17221;
wire v_17222;
wire v_17223;
wire v_17224;
wire v_17225;
wire v_17226;
wire v_17227;
wire v_17228;
wire v_17229;
wire v_17230;
wire v_17231;
wire v_17232;
wire v_17233;
wire v_17234;
wire v_17235;
wire v_17236;
wire v_17237;
wire v_17238;
wire v_17239;
wire v_17240;
wire v_17241;
wire v_17242;
wire v_17243;
wire v_17244;
wire v_17245;
wire v_17246;
wire v_17247;
wire v_17248;
wire v_17249;
wire v_17250;
wire v_17251;
wire v_17252;
wire v_17253;
wire v_17254;
wire v_17255;
wire v_17256;
wire v_17257;
wire v_17258;
wire v_17259;
wire v_17260;
wire v_17261;
wire v_17262;
wire v_17263;
wire v_17264;
wire v_17265;
wire v_17266;
wire v_17267;
wire v_17268;
wire v_17269;
wire v_17270;
wire v_17271;
wire v_17272;
wire v_17273;
wire v_17274;
wire v_17275;
wire v_17276;
wire v_17277;
wire v_17278;
wire v_17279;
wire v_17280;
wire v_17281;
wire v_17282;
wire v_17283;
wire v_17284;
wire v_17285;
wire v_17286;
wire v_17287;
wire v_17288;
wire v_17289;
wire v_17290;
wire v_17291;
wire v_17292;
wire v_17293;
wire v_17294;
wire v_17295;
wire v_17296;
wire v_17297;
wire v_17298;
wire v_17299;
wire v_17300;
wire v_17301;
wire v_17302;
wire v_17303;
wire v_17304;
wire v_17305;
wire v_17306;
wire v_17307;
wire v_17308;
wire v_17309;
wire v_17310;
wire v_17311;
wire v_17312;
wire v_17313;
wire v_17314;
wire v_17315;
wire v_17316;
wire v_17317;
wire v_17318;
wire v_17319;
wire v_17320;
wire v_17321;
wire v_17322;
wire v_17323;
wire v_17324;
wire v_17325;
wire v_17326;
wire v_17327;
wire v_17328;
wire v_17329;
wire v_17330;
wire v_17331;
wire v_17332;
wire v_17333;
wire v_17334;
wire v_17335;
wire v_17336;
wire v_17337;
wire v_17338;
wire v_17339;
wire v_17340;
wire v_17341;
wire v_17342;
wire v_17343;
wire v_17344;
wire v_17345;
wire v_17346;
wire v_17347;
wire v_17348;
wire v_17349;
wire v_17350;
wire v_17351;
wire v_17352;
wire v_17353;
wire v_17354;
wire v_17355;
wire v_17356;
wire v_17357;
wire v_17358;
wire v_17359;
wire v_17360;
wire v_17361;
wire v_17362;
wire v_17363;
wire v_17364;
wire v_17365;
wire v_17366;
wire v_17367;
wire v_17368;
wire v_17369;
wire v_17370;
wire v_17371;
wire v_17372;
wire v_17373;
wire v_17374;
wire v_17375;
wire v_17376;
wire v_17377;
wire v_17378;
wire v_17379;
wire v_17380;
wire v_17381;
wire v_17382;
wire v_17383;
wire v_17384;
wire v_17385;
wire v_17386;
wire v_17387;
wire v_17388;
wire v_17390;
wire v_17391;
wire v_17392;
wire v_17393;
wire v_17394;
wire v_17395;
wire v_17396;
wire v_17397;
wire v_17398;
wire v_17399;
wire v_17400;
wire v_17401;
wire v_17402;
wire v_17403;
wire v_17404;
wire v_17405;
wire v_17406;
wire v_17407;
wire v_17408;
wire v_17409;
wire v_17410;
wire v_17411;
wire v_17412;
wire v_17413;
wire v_17414;
wire v_17415;
wire v_17416;
wire v_17417;
wire v_17418;
wire v_17419;
wire v_17420;
wire v_17421;
wire v_17422;
wire v_17423;
wire v_17424;
wire v_17425;
wire v_17426;
wire v_17427;
wire v_17428;
wire v_17429;
wire v_17430;
wire v_17431;
wire v_17432;
wire v_17433;
wire v_17434;
wire v_17435;
wire v_17436;
wire v_17437;
wire v_17438;
wire v_17439;
wire v_17440;
wire v_17441;
wire v_17442;
wire v_17443;
wire v_17444;
wire v_17445;
wire v_17446;
wire v_17447;
wire v_17448;
wire v_17449;
wire v_17450;
wire v_17451;
wire v_17452;
wire v_17453;
wire v_17454;
wire v_17455;
wire v_17456;
wire v_17457;
wire v_17458;
wire v_17459;
wire v_17460;
wire v_17461;
wire v_17462;
wire v_17463;
wire v_17464;
wire v_17465;
wire v_17466;
wire v_17467;
wire v_17468;
wire v_17469;
wire v_17470;
wire v_17471;
wire v_17472;
wire v_17473;
wire v_17474;
wire v_17475;
wire v_17476;
wire v_17477;
wire v_17478;
wire v_17479;
wire v_17480;
wire v_17481;
wire v_17482;
wire v_17483;
wire v_17484;
wire v_17485;
wire v_17486;
wire v_17487;
wire v_17488;
wire v_17489;
wire v_17490;
wire v_17491;
wire v_17492;
wire v_17493;
wire v_17494;
wire v_17495;
wire v_17496;
wire v_17497;
wire v_17498;
wire v_17499;
wire v_17500;
wire v_17501;
wire v_17502;
wire v_17503;
wire v_17504;
wire v_17505;
wire v_17506;
wire v_17507;
wire v_17508;
wire v_17509;
wire v_17510;
wire v_17511;
wire v_17512;
wire v_17513;
wire v_17514;
wire v_17515;
wire v_17516;
wire v_17517;
wire v_17518;
wire v_17519;
wire v_17520;
wire v_17521;
wire v_17522;
wire v_17523;
wire v_17524;
wire v_17525;
wire v_17526;
wire v_17527;
wire v_17528;
wire v_17529;
wire v_17530;
wire v_17531;
wire v_17532;
wire v_17533;
wire v_17534;
wire v_17535;
wire v_17536;
wire v_17537;
wire v_17538;
wire v_17539;
wire v_17540;
wire v_17541;
wire v_17542;
wire v_17543;
wire v_17544;
wire v_17545;
wire v_17546;
wire v_17547;
wire v_17548;
wire v_17549;
wire v_17550;
wire v_17551;
wire v_17552;
wire v_17553;
wire v_17554;
wire v_17555;
wire v_17556;
wire v_17557;
wire v_17558;
wire v_17559;
wire v_17560;
wire v_17561;
wire v_17562;
wire v_17563;
wire v_17564;
wire v_17565;
wire v_17566;
wire v_17567;
wire v_17568;
wire v_17569;
wire v_17570;
wire v_17571;
wire v_17572;
wire v_17573;
wire v_17574;
wire v_17575;
wire v_17576;
wire v_17577;
wire v_17578;
wire v_17579;
wire v_17580;
wire v_17581;
wire v_17582;
wire v_17583;
wire v_17584;
wire v_17585;
wire v_17586;
wire v_17587;
wire v_17588;
wire v_17589;
wire v_17590;
wire v_17591;
wire v_17592;
wire v_17593;
wire v_17594;
wire v_17595;
wire v_17596;
wire v_17597;
wire v_17598;
wire v_17599;
wire v_17600;
wire v_17601;
wire v_17602;
wire v_17603;
wire v_17604;
wire v_17605;
wire v_17606;
wire v_17607;
wire v_17608;
wire v_17609;
wire v_17610;
wire v_17611;
wire v_17612;
wire v_17613;
wire v_17614;
wire v_17615;
wire v_17616;
wire v_17617;
wire v_17618;
wire v_17619;
wire v_17620;
wire v_17621;
wire v_17622;
wire v_17623;
wire v_17624;
wire v_17625;
wire v_17626;
wire v_17627;
wire v_17628;
wire v_17629;
wire v_17630;
wire v_17631;
wire v_17633;
wire v_17634;
wire v_17635;
wire v_17636;
wire v_17637;
wire v_17638;
wire v_17639;
wire v_17640;
wire v_17641;
wire v_17642;
wire v_17643;
wire v_17644;
wire v_17645;
wire v_17646;
wire v_17647;
wire v_17648;
wire v_17649;
wire v_17650;
wire v_17651;
wire v_17652;
wire v_17653;
wire v_17654;
wire v_17655;
wire v_17656;
wire v_17657;
wire v_17658;
wire v_17659;
wire v_17660;
wire v_17661;
wire v_17662;
wire v_17663;
wire v_17664;
wire v_17665;
wire v_17666;
wire v_17667;
wire v_17668;
wire v_17669;
wire v_17670;
wire v_17671;
wire v_17672;
wire v_17673;
wire v_17674;
wire v_17675;
wire v_17676;
wire v_17677;
wire v_17678;
wire v_17679;
wire v_17680;
wire v_17681;
wire v_17682;
wire v_17683;
wire v_17684;
wire v_17685;
wire v_17686;
wire v_17687;
wire v_17688;
wire v_17689;
wire v_17690;
wire v_17691;
wire v_17692;
wire v_17693;
wire v_17694;
wire v_17695;
wire v_17696;
wire v_17697;
wire v_17698;
wire v_17699;
wire v_17700;
wire v_17701;
wire v_17702;
wire v_17703;
wire v_17704;
wire v_17705;
wire v_17706;
wire v_17707;
wire v_17708;
wire v_17709;
wire v_17710;
wire v_17711;
wire v_17712;
wire v_17713;
wire v_17714;
wire v_17715;
wire v_17716;
wire v_17717;
wire v_17718;
wire v_17719;
wire v_17720;
wire v_17721;
wire v_17722;
wire v_17723;
wire v_17724;
wire v_17725;
wire v_17726;
wire v_17727;
wire v_17728;
wire v_17729;
wire v_17730;
wire v_17731;
wire v_17732;
wire v_17733;
wire v_17734;
wire v_17735;
wire v_17736;
wire v_17737;
wire v_17738;
wire v_17739;
wire v_17740;
wire v_17741;
wire v_17742;
wire v_17743;
wire v_17744;
wire v_17745;
wire v_17746;
wire v_17747;
wire v_17748;
wire v_17749;
wire v_17750;
wire v_17751;
wire v_17752;
wire v_17753;
wire v_17754;
wire v_17755;
wire v_17756;
wire v_17757;
wire v_17758;
wire v_17759;
wire v_17760;
wire v_17761;
wire v_17762;
wire v_17763;
wire v_17764;
wire v_17765;
wire v_17766;
wire v_17767;
wire v_17768;
wire v_17769;
wire v_17770;
wire v_17771;
wire v_17772;
wire v_17773;
wire v_17774;
wire v_17775;
wire v_17776;
wire v_17777;
wire v_17778;
wire v_17779;
wire v_17780;
wire v_17781;
wire v_17782;
wire v_17783;
wire v_17784;
wire v_17785;
wire v_17786;
wire v_17787;
wire v_17788;
wire v_17789;
wire v_17790;
wire v_17791;
wire v_17792;
wire v_17793;
wire v_17794;
wire v_17795;
wire v_17796;
wire v_17797;
wire v_17798;
wire v_17799;
wire v_17800;
wire v_17801;
wire v_17802;
wire v_17803;
wire v_17804;
wire v_17805;
wire v_17806;
wire v_17807;
wire v_17808;
wire v_17809;
wire v_17810;
wire v_17811;
wire v_17812;
wire v_17813;
wire v_17814;
wire v_17815;
wire v_17816;
wire v_17817;
wire v_17818;
wire v_17819;
wire v_17820;
wire v_17821;
wire v_17822;
wire v_17823;
wire v_17824;
wire v_17825;
wire v_17826;
wire v_17827;
wire v_17828;
wire v_17829;
wire v_17830;
wire v_17831;
wire v_17832;
wire v_17833;
wire v_17834;
wire v_17835;
wire v_17836;
wire v_17837;
wire v_17838;
wire v_17839;
wire v_17840;
wire v_17841;
wire v_17842;
wire v_17843;
wire v_17844;
wire v_17845;
wire v_17846;
wire v_17847;
wire v_17848;
wire v_17849;
wire v_17850;
wire v_17851;
wire v_17852;
wire v_17853;
wire v_17854;
wire v_17855;
wire v_17856;
wire v_17857;
wire v_17858;
wire v_17859;
wire v_17860;
wire v_17861;
wire v_17862;
wire v_17863;
wire v_17864;
wire v_17865;
wire v_17866;
wire v_17867;
wire v_17868;
wire v_17869;
wire v_17870;
wire v_17871;
wire v_17872;
wire v_17873;
wire v_17874;
wire v_17876;
wire v_17877;
wire v_17878;
wire v_17879;
wire v_17880;
wire v_17881;
wire v_17882;
wire v_17883;
wire v_17884;
wire v_17885;
wire v_17886;
wire v_17887;
wire v_17888;
wire v_17889;
wire v_17890;
wire v_17891;
wire v_17892;
wire v_17893;
wire v_17894;
wire v_17895;
wire v_17896;
wire v_17897;
wire v_17898;
wire v_17899;
wire v_17900;
wire v_17901;
wire v_17902;
wire v_17903;
wire v_17904;
wire v_17905;
wire v_17906;
wire v_17907;
wire v_17908;
wire v_17909;
wire v_17910;
wire v_17911;
wire v_17912;
wire v_17913;
wire v_17914;
wire v_17915;
wire v_17916;
wire v_17917;
wire v_17918;
wire v_17919;
wire v_17920;
wire v_17921;
wire v_17922;
wire v_17923;
wire v_17924;
wire v_17925;
wire v_17926;
wire v_17927;
wire v_17928;
wire v_17929;
wire v_17930;
wire v_17931;
wire v_17932;
wire v_17933;
wire v_17934;
wire v_17935;
wire v_17936;
wire v_17937;
wire v_17938;
wire v_17939;
wire v_17940;
wire v_17941;
wire v_17942;
wire v_17943;
wire v_17944;
wire v_17945;
wire v_17946;
wire v_17947;
wire v_17948;
wire v_17949;
wire v_17950;
wire v_17951;
wire v_17952;
wire v_17953;
wire v_17954;
wire v_17955;
wire v_17956;
wire v_17957;
wire v_17958;
wire v_17959;
wire v_17960;
wire v_17961;
wire v_17962;
wire v_17963;
wire v_17964;
wire v_17965;
wire v_17966;
wire v_17967;
wire v_17968;
wire v_17969;
wire v_17970;
wire v_17971;
wire v_17972;
wire v_17973;
wire v_17974;
wire v_17975;
wire v_17976;
wire v_17977;
wire v_17978;
wire v_17979;
wire v_17980;
wire v_17981;
wire v_17982;
wire v_17983;
wire v_17984;
wire v_17985;
wire v_17986;
wire v_17987;
wire v_17988;
wire v_17989;
wire v_17990;
wire v_17991;
wire v_17992;
wire v_17993;
wire v_17994;
wire v_17995;
wire v_17996;
wire v_17997;
wire v_17998;
wire v_17999;
wire v_18000;
wire v_18001;
wire v_18002;
wire v_18003;
wire v_18004;
wire v_18005;
wire v_18006;
wire v_18007;
wire v_18008;
wire v_18009;
wire v_18010;
wire v_18011;
wire v_18012;
wire v_18013;
wire v_18014;
wire v_18015;
wire v_18016;
wire v_18017;
wire v_18018;
wire v_18019;
wire v_18020;
wire v_18021;
wire v_18022;
wire v_18023;
wire v_18024;
wire v_18025;
wire v_18026;
wire v_18027;
wire v_18028;
wire v_18029;
wire v_18030;
wire v_18031;
wire v_18032;
wire v_18033;
wire v_18034;
wire v_18035;
wire v_18036;
wire v_18037;
wire v_18038;
wire v_18039;
wire v_18040;
wire v_18041;
wire v_18042;
wire v_18043;
wire v_18044;
wire v_18045;
wire v_18046;
wire v_18047;
wire v_18048;
wire v_18049;
wire v_18050;
wire v_18051;
wire v_18052;
wire v_18053;
wire v_18054;
wire v_18055;
wire v_18056;
wire v_18057;
wire v_18058;
wire v_18059;
wire v_18060;
wire v_18061;
wire v_18062;
wire v_18063;
wire v_18064;
wire v_18065;
wire v_18066;
wire v_18067;
wire v_18068;
wire v_18069;
wire v_18070;
wire v_18071;
wire v_18072;
wire v_18073;
wire v_18074;
wire v_18075;
wire v_18076;
wire v_18077;
wire v_18078;
wire v_18079;
wire v_18080;
wire v_18081;
wire v_18082;
wire v_18083;
wire v_18084;
wire v_18085;
wire v_18086;
wire v_18087;
wire v_18088;
wire v_18089;
wire v_18090;
wire v_18091;
wire v_18092;
wire v_18093;
wire v_18094;
wire v_18095;
wire v_18096;
wire v_18097;
wire v_18098;
wire v_18099;
wire v_18100;
wire v_18101;
wire v_18102;
wire v_18103;
wire v_18104;
wire v_18105;
wire v_18106;
wire v_18107;
wire v_18108;
wire v_18109;
wire v_18110;
wire v_18111;
wire v_18112;
wire v_18113;
wire v_18114;
wire v_18115;
wire v_18116;
wire v_18117;
wire v_18119;
wire v_18120;
wire v_18121;
wire v_18122;
wire v_18123;
wire v_18124;
wire v_18125;
wire v_18126;
wire v_18127;
wire v_18128;
wire v_18129;
wire v_18130;
wire v_18131;
wire v_18132;
wire v_18133;
wire v_18134;
wire v_18135;
wire v_18136;
wire v_18137;
wire v_18138;
wire v_18139;
wire v_18140;
wire v_18141;
wire v_18142;
wire v_18143;
wire v_18144;
wire v_18145;
wire v_18146;
wire v_18147;
wire v_18148;
wire v_18149;
wire v_18150;
wire v_18151;
wire v_18152;
wire v_18153;
wire v_18154;
wire v_18155;
wire v_18156;
wire v_18157;
wire v_18158;
wire v_18159;
wire v_18160;
wire v_18161;
wire v_18162;
wire v_18163;
wire v_18164;
wire v_18165;
wire v_18166;
wire v_18167;
wire v_18168;
wire v_18169;
wire v_18170;
wire v_18171;
wire v_18172;
wire v_18173;
wire v_18174;
wire v_18175;
wire v_18176;
wire v_18177;
wire v_18178;
wire v_18179;
wire v_18180;
wire v_18181;
wire v_18182;
wire v_18183;
wire v_18184;
wire v_18185;
wire v_18186;
wire v_18187;
wire v_18188;
wire v_18189;
wire v_18190;
wire v_18191;
wire v_18192;
wire v_18193;
wire v_18194;
wire v_18195;
wire v_18196;
wire v_18197;
wire v_18198;
wire v_18199;
wire v_18200;
wire v_18201;
wire v_18202;
wire v_18203;
wire v_18204;
wire v_18205;
wire v_18206;
wire v_18207;
wire v_18208;
wire v_18209;
wire v_18210;
wire v_18211;
wire v_18212;
wire v_18213;
wire v_18214;
wire v_18215;
wire v_18216;
wire v_18217;
wire v_18218;
wire v_18219;
wire v_18220;
wire v_18221;
wire v_18222;
wire v_18223;
wire v_18224;
wire v_18225;
wire v_18226;
wire v_18227;
wire v_18228;
wire v_18229;
wire v_18230;
wire v_18231;
wire v_18232;
wire v_18233;
wire v_18234;
wire v_18235;
wire v_18236;
wire v_18237;
wire v_18238;
wire v_18239;
wire v_18240;
wire v_18241;
wire v_18242;
wire v_18243;
wire v_18244;
wire v_18245;
wire v_18246;
wire v_18247;
wire v_18248;
wire v_18249;
wire v_18250;
wire v_18251;
wire v_18252;
wire v_18253;
wire v_18254;
wire v_18255;
wire v_18256;
wire v_18257;
wire v_18258;
wire v_18259;
wire v_18260;
wire v_18261;
wire v_18262;
wire v_18263;
wire v_18264;
wire v_18265;
wire v_18266;
wire v_18267;
wire v_18268;
wire v_18269;
wire v_18270;
wire v_18271;
wire v_18272;
wire v_18273;
wire v_18274;
wire v_18275;
wire v_18276;
wire v_18277;
wire v_18278;
wire v_18279;
wire v_18280;
wire v_18281;
wire v_18282;
wire v_18283;
wire v_18284;
wire v_18285;
wire v_18286;
wire v_18287;
wire v_18288;
wire v_18289;
wire v_18290;
wire v_18291;
wire v_18292;
wire v_18293;
wire v_18294;
wire v_18295;
wire v_18296;
wire v_18297;
wire v_18298;
wire v_18299;
wire v_18300;
wire v_18301;
wire v_18302;
wire v_18303;
wire v_18304;
wire v_18305;
wire v_18306;
wire v_18307;
wire v_18308;
wire v_18309;
wire v_18310;
wire v_18311;
wire v_18312;
wire v_18313;
wire v_18314;
wire v_18315;
wire v_18316;
wire v_18317;
wire v_18318;
wire v_18319;
wire v_18320;
wire v_18321;
wire v_18322;
wire v_18323;
wire v_18324;
wire v_18325;
wire v_18326;
wire v_18327;
wire v_18328;
wire v_18329;
wire v_18330;
wire v_18331;
wire v_18332;
wire v_18333;
wire v_18334;
wire v_18335;
wire v_18336;
wire v_18337;
wire v_18338;
wire v_18339;
wire v_18340;
wire v_18341;
wire v_18342;
wire v_18343;
wire v_18344;
wire v_18345;
wire v_18346;
wire v_18347;
wire v_18348;
wire v_18349;
wire v_18350;
wire v_18351;
wire v_18352;
wire v_18353;
wire v_18354;
wire v_18355;
wire v_18356;
wire v_18357;
wire v_18358;
wire v_18359;
wire v_18360;
wire v_18362;
wire v_18363;
wire v_18364;
wire v_18365;
wire v_18366;
wire v_18367;
wire v_18368;
wire v_18369;
wire v_18370;
wire v_18371;
wire v_18372;
wire v_18373;
wire v_18374;
wire v_18375;
wire v_18376;
wire v_18377;
wire v_18378;
wire v_18379;
wire v_18380;
wire v_18381;
wire v_18382;
wire v_18383;
wire v_18384;
wire v_18385;
wire v_18386;
wire v_18387;
wire v_18388;
wire v_18389;
wire v_18390;
wire v_18391;
wire v_18392;
wire v_18393;
wire v_18394;
wire v_18395;
wire v_18396;
wire v_18397;
wire v_18398;
wire v_18399;
wire v_18400;
wire v_18401;
wire v_18402;
wire v_18403;
wire v_18404;
wire v_18405;
wire v_18406;
wire v_18407;
wire v_18408;
wire v_18409;
wire v_18410;
wire v_18411;
wire v_18412;
wire v_18413;
wire v_18414;
wire v_18415;
wire v_18416;
wire v_18417;
wire v_18418;
wire v_18419;
wire v_18420;
wire v_18421;
wire v_18422;
wire v_18423;
wire v_18424;
wire v_18425;
wire v_18426;
wire v_18427;
wire v_18428;
wire v_18429;
wire v_18430;
wire v_18431;
wire v_18432;
wire v_18433;
wire v_18434;
wire v_18435;
wire v_18436;
wire v_18437;
wire v_18438;
wire v_18439;
wire v_18440;
wire v_18441;
wire v_18442;
wire v_18443;
wire v_18444;
wire v_18445;
wire v_18446;
wire v_18447;
wire v_18448;
wire v_18449;
wire v_18450;
wire v_18451;
wire v_18452;
wire v_18453;
wire v_18454;
wire v_18455;
wire v_18456;
wire v_18457;
wire v_18458;
wire v_18459;
wire v_18460;
wire v_18461;
wire v_18462;
wire v_18463;
wire v_18464;
wire v_18465;
wire v_18466;
wire v_18467;
wire v_18468;
wire v_18469;
wire v_18470;
wire v_18471;
wire v_18472;
wire v_18473;
wire v_18474;
wire v_18475;
wire v_18476;
wire v_18477;
wire v_18478;
wire v_18479;
wire v_18480;
wire v_18481;
wire v_18482;
wire v_18483;
wire v_18484;
wire v_18485;
wire v_18486;
wire v_18487;
wire v_18488;
wire v_18489;
wire v_18490;
wire v_18491;
wire v_18492;
wire v_18493;
wire v_18494;
wire v_18495;
wire v_18496;
wire v_18497;
wire v_18498;
wire v_18499;
wire v_18500;
wire v_18501;
wire v_18502;
wire v_18503;
wire v_18504;
wire v_18505;
wire v_18506;
wire v_18507;
wire v_18508;
wire v_18509;
wire v_18510;
wire v_18511;
wire v_18512;
wire v_18513;
wire v_18514;
wire v_18515;
wire v_18516;
wire v_18517;
wire v_18518;
wire v_18519;
wire v_18520;
wire v_18521;
wire v_18522;
wire v_18523;
wire v_18524;
wire v_18525;
wire v_18526;
wire v_18527;
wire v_18528;
wire v_18529;
wire v_18530;
wire v_18531;
wire v_18532;
wire v_18533;
wire v_18534;
wire v_18535;
wire v_18536;
wire v_18537;
wire v_18538;
wire v_18539;
wire v_18540;
wire v_18541;
wire v_18542;
wire v_18543;
wire v_18544;
wire v_18545;
wire v_18546;
wire v_18547;
wire v_18548;
wire v_18549;
wire v_18550;
wire v_18551;
wire v_18552;
wire v_18553;
wire v_18554;
wire v_18555;
wire v_18556;
wire v_18557;
wire v_18558;
wire v_18559;
wire v_18560;
wire v_18561;
wire v_18562;
wire v_18563;
wire v_18564;
wire v_18565;
wire v_18566;
wire v_18567;
wire v_18568;
wire v_18569;
wire v_18570;
wire v_18571;
wire v_18572;
wire v_18573;
wire v_18574;
wire v_18575;
wire v_18576;
wire v_18577;
wire v_18578;
wire v_18579;
wire v_18580;
wire v_18581;
wire v_18582;
wire v_18583;
wire v_18584;
wire v_18585;
wire v_18586;
wire v_18587;
wire v_18588;
wire v_18589;
wire v_18590;
wire v_18591;
wire v_18592;
wire v_18593;
wire v_18594;
wire v_18595;
wire v_18596;
wire v_18597;
wire v_18598;
wire v_18599;
wire v_18600;
wire v_18601;
wire v_18602;
wire v_18603;
wire v_18605;
wire v_18606;
wire v_18607;
wire v_18608;
wire v_18609;
wire v_18610;
wire v_18611;
wire v_18612;
wire v_18613;
wire v_18614;
wire v_18615;
wire v_18616;
wire v_18617;
wire v_18618;
wire v_18619;
wire v_18620;
wire v_18621;
wire v_18622;
wire v_18623;
wire v_18624;
wire v_18625;
wire v_18626;
wire v_18627;
wire v_18628;
wire v_18629;
wire v_18630;
wire v_18631;
wire v_18632;
wire v_18633;
wire v_18634;
wire v_18635;
wire v_18636;
wire v_18637;
wire v_18638;
wire v_18639;
wire v_18640;
wire v_18641;
wire v_18642;
wire v_18643;
wire v_18644;
wire v_18645;
wire v_18646;
wire v_18647;
wire v_18648;
wire v_18649;
wire v_18650;
wire v_18651;
wire v_18652;
wire v_18653;
wire v_18654;
wire v_18655;
wire v_18656;
wire v_18657;
wire v_18658;
wire v_18659;
wire v_18660;
wire v_18661;
wire v_18662;
wire v_18663;
wire v_18664;
wire v_18665;
wire v_18666;
wire v_18667;
wire v_18668;
wire v_18669;
wire v_18670;
wire v_18671;
wire v_18672;
wire v_18673;
wire v_18674;
wire v_18675;
wire v_18676;
wire v_18677;
wire v_18678;
wire v_18679;
wire v_18680;
wire v_18681;
wire v_18682;
wire v_18683;
wire v_18684;
wire v_18685;
wire v_18686;
wire v_18687;
wire v_18688;
wire v_18689;
wire v_18690;
wire v_18691;
wire v_18692;
wire v_18693;
wire v_18694;
wire v_18695;
wire v_18696;
wire v_18697;
wire v_18698;
wire v_18699;
wire v_18700;
wire v_18701;
wire v_18702;
wire v_18703;
wire v_18704;
wire v_18705;
wire v_18706;
wire v_18707;
wire v_18708;
wire v_18709;
wire v_18710;
wire v_18711;
wire v_18712;
wire v_18713;
wire v_18714;
wire v_18715;
wire v_18716;
wire v_18717;
wire v_18718;
wire v_18719;
wire v_18720;
wire v_18721;
wire v_18722;
wire v_18723;
wire v_18724;
wire v_18725;
wire v_18726;
wire v_18727;
wire v_18728;
wire v_18729;
wire v_18730;
wire v_18731;
wire v_18732;
wire v_18733;
wire v_18734;
wire v_18735;
wire v_18736;
wire v_18737;
wire v_18738;
wire v_18739;
wire v_18740;
wire v_18741;
wire v_18742;
wire v_18743;
wire v_18744;
wire v_18745;
wire v_18746;
wire v_18747;
wire v_18748;
wire v_18749;
wire v_18750;
wire v_18751;
wire v_18752;
wire v_18753;
wire v_18754;
wire v_18755;
wire v_18756;
wire v_18757;
wire v_18758;
wire v_18759;
wire v_18760;
wire v_18761;
wire v_18762;
wire v_18763;
wire v_18764;
wire v_18765;
wire v_18766;
wire v_18767;
wire v_18768;
wire v_18769;
wire v_18770;
wire v_18771;
wire v_18772;
wire v_18773;
wire v_18774;
wire v_18775;
wire v_18776;
wire v_18777;
wire v_18778;
wire v_18779;
wire v_18780;
wire v_18781;
wire v_18782;
wire v_18783;
wire v_18784;
wire v_18785;
wire v_18786;
wire v_18787;
wire v_18788;
wire v_18789;
wire v_18790;
wire v_18791;
wire v_18792;
wire v_18793;
wire v_18794;
wire v_18795;
wire v_18796;
wire v_18797;
wire v_18798;
wire v_18799;
wire v_18800;
wire v_18801;
wire v_18802;
wire v_18803;
wire v_18804;
wire v_18805;
wire v_18806;
wire v_18807;
wire v_18808;
wire v_18809;
wire v_18810;
wire v_18811;
wire v_18812;
wire v_18813;
wire v_18814;
wire v_18815;
wire v_18816;
wire v_18817;
wire v_18818;
wire v_18819;
wire v_18820;
wire v_18821;
wire v_18822;
wire v_18823;
wire v_18824;
wire v_18825;
wire v_18826;
wire v_18827;
wire v_18828;
wire v_18829;
wire v_18830;
wire v_18831;
wire v_18832;
wire v_18833;
wire v_18834;
wire v_18835;
wire v_18836;
wire v_18837;
wire v_18838;
wire v_18839;
wire v_18840;
wire v_18841;
wire v_18842;
wire v_18843;
wire v_18844;
wire v_18845;
wire v_18846;
wire v_18848;
wire v_18849;
wire v_18850;
wire v_18851;
wire v_18852;
wire v_18853;
wire v_18854;
wire v_18855;
wire v_18856;
wire v_18857;
wire v_18858;
wire v_18859;
wire v_18860;
wire v_18861;
wire v_18862;
wire v_18863;
wire v_18864;
wire v_18865;
wire v_18866;
wire v_18867;
wire v_18868;
wire v_18869;
wire v_18870;
wire v_18871;
wire v_18872;
wire v_18873;
wire v_18874;
wire v_18875;
wire v_18876;
wire v_18877;
wire v_18878;
wire v_18879;
wire v_18880;
wire v_18881;
wire v_18882;
wire v_18883;
wire v_18884;
wire v_18885;
wire v_18886;
wire v_18887;
wire v_18888;
wire v_18889;
wire v_18890;
wire v_18891;
wire v_18892;
wire v_18893;
wire v_18894;
wire v_18895;
wire v_18896;
wire v_18897;
wire v_18898;
wire v_18899;
wire v_18900;
wire v_18901;
wire v_18902;
wire v_18903;
wire v_18904;
wire v_18905;
wire v_18906;
wire v_18907;
wire v_18908;
wire v_18909;
wire v_18910;
wire v_18911;
wire v_18912;
wire v_18913;
wire v_18914;
wire v_18915;
wire v_18916;
wire v_18917;
wire v_18918;
wire v_18919;
wire v_18920;
wire v_18921;
wire v_18922;
wire v_18923;
wire v_18924;
wire v_18925;
wire v_18926;
wire v_18927;
wire v_18928;
wire v_18929;
wire v_18930;
wire v_18931;
wire v_18932;
wire v_18933;
wire v_18934;
wire v_18935;
wire v_18936;
wire v_18937;
wire v_18938;
wire v_18939;
wire v_18940;
wire v_18941;
wire v_18942;
wire v_18943;
wire v_18944;
wire v_18945;
wire v_18946;
wire v_18947;
wire v_18948;
wire v_18949;
wire v_18950;
wire v_18951;
wire v_18952;
wire v_18953;
wire v_18954;
wire v_18955;
wire v_18956;
wire v_18957;
wire v_18958;
wire v_18959;
wire v_18960;
wire v_18961;
wire v_18962;
wire v_18963;
wire v_18964;
wire v_18965;
wire v_18966;
wire v_18967;
wire v_18968;
wire v_18969;
wire v_18970;
wire v_18971;
wire v_18972;
wire v_18973;
wire v_18974;
wire v_18975;
wire v_18976;
wire v_18977;
wire v_18978;
wire v_18979;
wire v_18980;
wire v_18981;
wire v_18982;
wire v_18983;
wire v_18984;
wire v_18985;
wire v_18986;
wire v_18987;
wire v_18988;
wire v_18989;
wire v_18990;
wire v_18991;
wire v_18992;
wire v_18993;
wire v_18994;
wire v_18995;
wire v_18996;
wire v_18997;
wire v_18998;
wire v_18999;
wire v_19000;
wire v_19001;
wire v_19002;
wire v_19003;
wire v_19004;
wire v_19005;
wire v_19006;
wire v_19007;
wire v_19008;
wire v_19009;
wire v_19010;
wire v_19011;
wire v_19012;
wire v_19013;
wire v_19014;
wire v_19015;
wire v_19016;
wire v_19017;
wire v_19018;
wire v_19019;
wire v_19020;
wire v_19021;
wire v_19022;
wire v_19023;
wire v_19024;
wire v_19025;
wire v_19026;
wire v_19027;
wire v_19028;
wire v_19029;
wire v_19030;
wire v_19031;
wire v_19032;
wire v_19033;
wire v_19034;
wire v_19035;
wire v_19036;
wire v_19037;
wire v_19038;
wire v_19039;
wire v_19040;
wire v_19041;
wire v_19042;
wire v_19043;
wire v_19044;
wire v_19045;
wire v_19046;
wire v_19047;
wire v_19048;
wire v_19049;
wire v_19050;
wire v_19051;
wire v_19052;
wire v_19053;
wire v_19054;
wire v_19055;
wire v_19056;
wire v_19057;
wire v_19058;
wire v_19059;
wire v_19060;
wire v_19061;
wire v_19062;
wire v_19063;
wire v_19064;
wire v_19065;
wire v_19066;
wire v_19067;
wire v_19068;
wire v_19069;
wire v_19070;
wire v_19071;
wire v_19072;
wire v_19073;
wire v_19074;
wire v_19075;
wire v_19076;
wire v_19077;
wire v_19078;
wire v_19079;
wire v_19080;
wire v_19081;
wire v_19082;
wire v_19083;
wire v_19084;
wire v_19085;
wire v_19086;
wire v_19087;
wire v_19088;
wire v_19089;
wire v_19091;
wire v_19092;
wire v_19093;
wire v_19094;
wire v_19095;
wire v_19096;
wire v_19097;
wire v_19098;
wire v_19099;
wire v_19100;
wire v_19101;
wire v_19102;
wire v_19103;
wire v_19104;
wire v_19105;
wire v_19106;
wire v_19107;
wire v_19108;
wire v_19109;
wire v_19110;
wire v_19111;
wire v_19112;
wire v_19113;
wire v_19114;
wire v_19115;
wire v_19116;
wire v_19117;
wire v_19118;
wire v_19119;
wire v_19120;
wire v_19121;
wire v_19122;
wire v_19123;
wire v_19124;
wire v_19125;
wire v_19126;
wire v_19127;
wire v_19128;
wire v_19129;
wire v_19130;
wire v_19131;
wire v_19132;
wire v_19133;
wire v_19134;
wire v_19135;
wire v_19136;
wire v_19137;
wire v_19138;
wire v_19139;
wire v_19140;
wire v_19141;
wire v_19142;
wire v_19143;
wire v_19144;
wire v_19145;
wire v_19146;
wire v_19147;
wire v_19148;
wire v_19149;
wire v_19150;
wire v_19151;
wire v_19152;
wire v_19153;
wire v_19154;
wire v_19155;
wire v_19156;
wire v_19157;
wire v_19158;
wire v_19159;
wire v_19160;
wire v_19161;
wire v_19162;
wire v_19163;
wire v_19164;
wire v_19165;
wire v_19166;
wire v_19167;
wire v_19168;
wire v_19169;
wire v_19170;
wire v_19171;
wire v_19172;
wire v_19173;
wire v_19174;
wire v_19175;
wire v_19176;
wire v_19177;
wire v_19178;
wire v_19179;
wire v_19180;
wire v_19181;
wire v_19182;
wire v_19183;
wire v_19184;
wire v_19185;
wire v_19186;
wire v_19187;
wire v_19188;
wire v_19189;
wire v_19190;
wire v_19191;
wire v_19192;
wire v_19193;
wire v_19194;
wire v_19195;
wire v_19196;
wire v_19197;
wire v_19198;
wire v_19199;
wire v_19200;
wire v_19201;
wire v_19202;
wire v_19203;
wire v_19204;
wire v_19205;
wire v_19206;
wire v_19207;
wire v_19208;
wire v_19209;
wire v_19210;
wire v_19211;
wire v_19212;
wire v_19213;
wire v_19214;
wire v_19215;
wire v_19216;
wire v_19217;
wire v_19218;
wire v_19219;
wire v_19220;
wire v_19221;
wire v_19222;
wire v_19223;
wire v_19224;
wire v_19225;
wire v_19226;
wire v_19227;
wire v_19228;
wire v_19229;
wire v_19230;
wire v_19231;
wire v_19232;
wire v_19233;
wire v_19234;
wire v_19235;
wire v_19236;
wire v_19237;
wire v_19238;
wire v_19239;
wire v_19240;
wire v_19241;
wire v_19242;
wire v_19243;
wire v_19244;
wire v_19245;
wire v_19246;
wire v_19247;
wire v_19248;
wire v_19249;
wire v_19250;
wire v_19251;
wire v_19252;
wire v_19253;
wire v_19254;
wire v_19255;
wire v_19256;
wire v_19257;
wire v_19258;
wire v_19259;
wire v_19260;
wire v_19261;
wire v_19262;
wire v_19263;
wire v_19264;
wire v_19265;
wire v_19266;
wire v_19267;
wire v_19268;
wire v_19269;
wire v_19270;
wire v_19271;
wire v_19272;
wire v_19273;
wire v_19274;
wire v_19275;
wire v_19276;
wire v_19277;
wire v_19278;
wire v_19279;
wire v_19280;
wire v_19281;
wire v_19282;
wire v_19283;
wire v_19284;
wire v_19285;
wire v_19286;
wire v_19287;
wire v_19288;
wire v_19289;
wire v_19290;
wire v_19291;
wire v_19292;
wire v_19293;
wire v_19294;
wire v_19295;
wire v_19296;
wire v_19297;
wire v_19298;
wire v_19299;
wire v_19300;
wire v_19301;
wire v_19302;
wire v_19303;
wire v_19304;
wire v_19305;
wire v_19306;
wire v_19307;
wire v_19308;
wire v_19309;
wire v_19310;
wire v_19311;
wire v_19312;
wire v_19313;
wire v_19314;
wire v_19315;
wire v_19316;
wire v_19317;
wire v_19318;
wire v_19319;
wire v_19320;
wire v_19321;
wire v_19322;
wire v_19323;
wire v_19324;
wire v_19325;
wire v_19326;
wire v_19327;
wire v_19328;
wire v_19329;
wire v_19330;
wire v_19331;
wire v_19332;
wire v_19334;
wire v_19335;
wire v_19336;
wire v_19337;
wire v_19338;
wire v_19339;
wire v_19340;
wire v_19341;
wire v_19342;
wire v_19343;
wire v_19344;
wire v_19345;
wire v_19346;
wire v_19347;
wire v_19348;
wire v_19349;
wire v_19350;
wire v_19351;
wire v_19352;
wire v_19353;
wire v_19354;
wire v_19355;
wire v_19356;
wire v_19357;
wire v_19358;
wire v_19359;
wire v_19360;
wire v_19361;
wire v_19362;
wire v_19363;
wire v_19364;
wire v_19365;
wire v_19366;
wire v_19367;
wire v_19368;
wire v_19369;
wire v_19370;
wire v_19371;
wire v_19372;
wire v_19373;
wire v_19374;
wire v_19375;
wire v_19376;
wire v_19377;
wire v_19378;
wire v_19379;
wire v_19380;
wire v_19381;
wire v_19382;
wire v_19383;
wire v_19384;
wire v_19385;
wire v_19386;
wire v_19387;
wire v_19388;
wire v_19389;
wire v_19390;
wire v_19391;
wire v_19392;
wire v_19393;
wire v_19394;
wire v_19395;
wire v_19396;
wire v_19397;
wire v_19398;
wire v_19399;
wire v_19400;
wire v_19401;
wire v_19402;
wire v_19403;
wire v_19404;
wire v_19405;
wire v_19406;
wire v_19407;
wire v_19408;
wire v_19409;
wire v_19410;
wire v_19411;
wire v_19412;
wire v_19413;
wire v_19414;
wire v_19415;
wire v_19416;
wire v_19417;
wire v_19418;
wire v_19419;
wire v_19420;
wire v_19421;
wire v_19422;
wire v_19423;
wire v_19424;
wire v_19425;
wire v_19426;
wire v_19427;
wire v_19428;
wire v_19429;
wire v_19430;
wire v_19431;
wire v_19432;
wire v_19433;
wire v_19434;
wire v_19435;
wire v_19436;
wire v_19437;
wire v_19438;
wire v_19439;
wire v_19440;
wire v_19441;
wire v_19442;
wire v_19443;
wire v_19444;
wire v_19445;
wire v_19446;
wire v_19447;
wire v_19448;
wire v_19449;
wire v_19450;
wire v_19451;
wire v_19452;
wire v_19453;
wire v_19454;
wire v_19455;
wire v_19456;
wire v_19457;
wire v_19458;
wire v_19459;
wire v_19460;
wire v_19461;
wire v_19462;
wire v_19463;
wire v_19464;
wire v_19465;
wire v_19466;
wire v_19467;
wire v_19468;
wire v_19469;
wire v_19470;
wire v_19471;
wire v_19472;
wire v_19473;
wire v_19474;
wire v_19475;
wire v_19476;
wire v_19477;
wire v_19478;
wire v_19479;
wire v_19480;
wire v_19481;
wire v_19482;
wire v_19483;
wire v_19484;
wire v_19485;
wire v_19486;
wire v_19487;
wire v_19488;
wire v_19489;
wire v_19490;
wire v_19491;
wire v_19492;
wire v_19493;
wire v_19494;
wire v_19495;
wire v_19496;
wire v_19497;
wire v_19498;
wire v_19499;
wire v_19500;
wire v_19501;
wire v_19502;
wire v_19503;
wire v_19504;
wire v_19505;
wire v_19506;
wire v_19507;
wire v_19508;
wire v_19509;
wire v_19510;
wire v_19511;
wire v_19512;
wire v_19513;
wire v_19514;
wire v_19515;
wire v_19516;
wire v_19517;
wire v_19518;
wire v_19519;
wire v_19520;
wire v_19521;
wire v_19522;
wire v_19523;
wire v_19524;
wire v_19525;
wire v_19526;
wire v_19527;
wire v_19528;
wire v_19529;
wire v_19530;
wire v_19531;
wire v_19532;
wire v_19533;
wire v_19534;
wire v_19535;
wire v_19536;
wire v_19537;
wire v_19538;
wire v_19539;
wire v_19540;
wire v_19541;
wire v_19542;
wire v_19543;
wire v_19544;
wire v_19545;
wire v_19546;
wire v_19547;
wire v_19548;
wire v_19549;
wire v_19550;
wire v_19551;
wire v_19552;
wire v_19553;
wire v_19554;
wire v_19555;
wire v_19556;
wire v_19557;
wire v_19558;
wire v_19559;
wire v_19560;
wire v_19561;
wire v_19562;
wire v_19563;
wire v_19564;
wire v_19565;
wire v_19566;
wire v_19567;
wire v_19568;
wire v_19569;
wire v_19570;
wire v_19571;
wire v_19572;
wire v_19573;
wire v_19574;
wire v_19575;
wire v_19577;
wire v_19578;
wire v_19579;
wire v_19580;
wire v_19581;
wire v_19582;
wire v_19583;
wire v_19584;
wire v_19585;
wire v_19586;
wire v_19587;
wire v_19588;
wire v_19589;
wire v_19590;
wire v_19591;
wire v_19592;
wire v_19593;
wire v_19594;
wire v_19595;
wire v_19596;
wire v_19597;
wire v_19598;
wire v_19599;
wire v_19600;
wire v_19601;
wire v_19602;
wire v_19603;
wire v_19604;
wire v_19605;
wire v_19606;
wire v_19607;
wire v_19608;
wire v_19609;
wire v_19610;
wire v_19611;
wire v_19612;
wire v_19613;
wire v_19614;
wire v_19615;
wire v_19616;
wire v_19617;
wire v_19618;
wire v_19619;
wire v_19620;
wire v_19621;
wire v_19622;
wire v_19623;
wire v_19624;
wire v_19625;
wire v_19626;
wire v_19627;
wire v_19628;
wire v_19629;
wire v_19630;
wire v_19631;
wire v_19632;
wire v_19633;
wire v_19634;
wire v_19635;
wire v_19636;
wire v_19637;
wire v_19638;
wire v_19639;
wire v_19640;
wire v_19641;
wire v_19642;
wire v_19643;
wire v_19644;
wire v_19645;
wire v_19646;
wire v_19647;
wire v_19648;
wire v_19649;
wire v_19650;
wire v_19651;
wire v_19652;
wire v_19653;
wire v_19654;
wire v_19655;
wire v_19656;
wire v_19657;
wire v_19658;
wire v_19659;
wire v_19660;
wire v_19661;
wire v_19662;
wire v_19663;
wire v_19664;
wire v_19665;
wire v_19666;
wire v_19667;
wire v_19668;
wire v_19669;
wire v_19670;
wire v_19671;
wire v_19672;
wire v_19673;
wire v_19674;
wire v_19675;
wire v_19676;
wire v_19677;
wire v_19678;
wire v_19679;
wire v_19680;
wire v_19681;
wire v_19682;
wire v_19683;
wire v_19684;
wire v_19685;
wire v_19686;
wire v_19687;
wire v_19688;
wire v_19689;
wire v_19690;
wire v_19691;
wire v_19692;
wire v_19693;
wire v_19694;
wire v_19695;
wire v_19696;
wire v_19697;
wire v_19698;
wire v_19699;
wire v_19700;
wire v_19701;
wire v_19702;
wire v_19703;
wire v_19704;
wire v_19705;
wire v_19706;
wire v_19707;
wire v_19708;
wire v_19709;
wire v_19710;
wire v_19711;
wire v_19712;
wire v_19713;
wire v_19714;
wire v_19715;
wire v_19716;
wire v_19717;
wire v_19718;
wire v_19719;
wire v_19720;
wire v_19721;
wire v_19722;
wire v_19723;
wire v_19724;
wire v_19725;
wire v_19726;
wire v_19727;
wire v_19728;
wire v_19729;
wire v_19730;
wire v_19731;
wire v_19732;
wire v_19733;
wire v_19734;
wire v_19735;
wire v_19736;
wire v_19737;
wire v_19738;
wire v_19739;
wire v_19740;
wire v_19741;
wire v_19742;
wire v_19743;
wire v_19744;
wire v_19745;
wire v_19746;
wire v_19747;
wire v_19748;
wire v_19749;
wire v_19750;
wire v_19751;
wire v_19752;
wire v_19753;
wire v_19754;
wire v_19755;
wire v_19756;
wire v_19757;
wire v_19758;
wire v_19759;
wire v_19760;
wire v_19761;
wire v_19762;
wire v_19763;
wire v_19764;
wire v_19765;
wire v_19766;
wire v_19767;
wire v_19768;
wire v_19769;
wire v_19770;
wire v_19771;
wire v_19772;
wire v_19773;
wire v_19774;
wire v_19775;
wire v_19776;
wire v_19777;
wire v_19778;
wire v_19779;
wire v_19780;
wire v_19781;
wire v_19782;
wire v_19783;
wire v_19784;
wire v_19785;
wire v_19786;
wire v_19787;
wire v_19788;
wire v_19789;
wire v_19790;
wire v_19791;
wire v_19792;
wire v_19793;
wire v_19794;
wire v_19795;
wire v_19796;
wire v_19797;
wire v_19798;
wire v_19799;
wire v_19800;
wire v_19801;
wire v_19802;
wire v_19803;
wire v_19804;
wire v_19805;
wire v_19806;
wire v_19807;
wire v_19808;
wire v_19809;
wire v_19810;
wire v_19811;
wire v_19812;
wire v_19813;
wire v_19814;
wire v_19815;
wire v_19816;
wire v_19817;
wire v_19818;
wire v_19820;
wire v_19821;
wire v_19822;
wire v_19823;
wire v_19824;
wire v_19825;
wire v_19826;
wire v_19827;
wire v_19828;
wire v_19829;
wire v_19830;
wire v_19831;
wire v_19832;
wire v_19833;
wire v_19834;
wire v_19835;
wire v_19836;
wire v_19837;
wire v_19838;
wire v_19839;
wire v_19840;
wire v_19841;
wire v_19842;
wire v_19843;
wire v_19844;
wire v_19845;
wire v_19846;
wire v_19847;
wire v_19848;
wire v_19849;
wire v_19850;
wire v_19851;
wire v_19852;
wire v_19853;
wire v_19854;
wire v_19855;
wire v_19856;
wire v_19857;
wire v_19858;
wire v_19859;
wire v_19860;
wire v_19861;
wire v_19862;
wire v_19863;
wire v_19864;
wire v_19865;
wire v_19866;
wire v_19867;
wire v_19868;
wire v_19869;
wire v_19870;
wire v_19871;
wire v_19872;
wire v_19873;
wire v_19874;
wire v_19875;
wire v_19876;
wire v_19877;
wire v_19878;
wire v_19879;
wire v_19880;
wire v_19881;
wire v_19882;
wire v_19883;
wire v_19884;
wire v_19885;
wire v_19886;
wire v_19887;
wire v_19888;
wire v_19889;
wire v_19890;
wire v_19891;
wire v_19892;
wire v_19893;
wire v_19894;
wire v_19895;
wire v_19896;
wire v_19897;
wire v_19898;
wire v_19899;
wire v_19900;
wire v_19901;
wire v_19902;
wire v_19903;
wire v_19904;
wire v_19905;
wire v_19906;
wire v_19907;
wire v_19908;
wire v_19909;
wire v_19910;
wire v_19911;
wire v_19912;
wire v_19913;
wire v_19914;
wire v_19915;
wire v_19916;
wire v_19917;
wire v_19918;
wire v_19919;
wire v_19920;
wire v_19921;
wire v_19922;
wire v_19923;
wire v_19924;
wire v_19925;
wire v_19926;
wire v_19927;
wire v_19928;
wire v_19929;
wire v_19930;
wire v_19931;
wire v_19932;
wire v_19933;
wire v_19934;
wire v_19935;
wire v_19936;
wire v_19937;
wire v_19938;
wire v_19939;
wire v_19940;
wire v_19941;
wire v_19942;
wire v_19943;
wire v_19944;
wire v_19945;
wire v_19946;
wire v_19947;
wire v_19948;
wire v_19949;
wire v_19950;
wire v_19951;
wire v_19952;
wire v_19953;
wire v_19954;
wire v_19955;
wire v_19956;
wire v_19957;
wire v_19958;
wire v_19959;
wire v_19960;
wire v_19961;
wire v_19962;
wire v_19963;
wire v_19964;
wire v_19965;
wire v_19966;
wire v_19967;
wire v_19968;
wire v_19969;
wire v_19970;
wire v_19971;
wire v_19972;
wire v_19973;
wire v_19974;
wire v_19975;
wire v_19976;
wire v_19977;
wire v_19978;
wire v_19979;
wire v_19980;
wire v_19981;
wire v_19982;
wire v_19983;
wire v_19984;
wire v_19985;
wire v_19986;
wire v_19987;
wire v_19988;
wire v_19989;
wire v_19990;
wire v_19991;
wire v_19992;
wire v_19993;
wire v_19994;
wire v_19995;
wire v_19996;
wire v_19997;
wire v_19998;
wire v_19999;
wire v_20000;
wire v_20001;
wire v_20002;
wire v_20003;
wire v_20004;
wire v_20005;
wire v_20006;
wire v_20007;
wire v_20008;
wire v_20009;
wire v_20010;
wire v_20011;
wire v_20012;
wire v_20013;
wire v_20014;
wire v_20015;
wire v_20016;
wire v_20017;
wire v_20018;
wire v_20019;
wire v_20020;
wire v_20021;
wire v_20022;
wire v_20023;
wire v_20024;
wire v_20025;
wire v_20026;
wire v_20027;
wire v_20028;
wire v_20029;
wire v_20030;
wire v_20031;
wire v_20032;
wire v_20033;
wire v_20034;
wire v_20035;
wire v_20036;
wire v_20037;
wire v_20038;
wire v_20039;
wire v_20040;
wire v_20041;
wire v_20042;
wire v_20043;
wire v_20044;
wire v_20045;
wire v_20046;
wire v_20047;
wire v_20048;
wire v_20049;
wire v_20050;
wire v_20051;
wire v_20052;
wire v_20053;
wire v_20054;
wire v_20055;
wire v_20056;
wire v_20057;
wire v_20058;
wire v_20059;
wire v_20060;
wire v_20061;
wire v_20063;
wire v_20064;
wire v_20065;
wire v_20066;
wire v_20067;
wire v_20068;
wire v_20069;
wire v_20070;
wire v_20071;
wire v_20072;
wire v_20073;
wire v_20074;
wire v_20075;
wire v_20076;
wire v_20077;
wire v_20078;
wire v_20079;
wire v_20080;
wire v_20081;
wire v_20082;
wire v_20083;
wire v_20084;
wire v_20085;
wire v_20086;
wire v_20087;
wire v_20088;
wire v_20089;
wire v_20090;
wire v_20091;
wire v_20092;
wire v_20093;
wire v_20094;
wire v_20095;
wire v_20096;
wire v_20097;
wire v_20098;
wire v_20099;
wire v_20100;
wire v_20101;
wire v_20102;
wire v_20103;
wire v_20104;
wire v_20105;
wire v_20106;
wire v_20107;
wire v_20108;
wire v_20109;
wire v_20110;
wire v_20111;
wire v_20112;
wire v_20113;
wire v_20114;
wire v_20115;
wire v_20116;
wire v_20117;
wire v_20118;
wire v_20119;
wire v_20120;
wire v_20121;
wire v_20122;
wire v_20123;
wire v_20124;
wire v_20125;
wire v_20126;
wire v_20127;
wire v_20128;
wire v_20129;
wire v_20130;
wire v_20131;
wire v_20132;
wire v_20133;
wire v_20134;
wire v_20135;
wire v_20136;
wire v_20137;
wire v_20138;
wire v_20139;
wire v_20140;
wire v_20141;
wire v_20142;
wire v_20143;
wire v_20144;
wire v_20145;
wire v_20146;
wire v_20147;
wire v_20148;
wire v_20149;
wire v_20150;
wire v_20151;
wire v_20152;
wire v_20153;
wire v_20154;
wire v_20155;
wire v_20156;
wire v_20157;
wire v_20158;
wire v_20159;
wire v_20160;
wire v_20161;
wire v_20162;
wire v_20163;
wire v_20164;
wire v_20165;
wire v_20166;
wire v_20167;
wire v_20168;
wire v_20169;
wire v_20170;
wire v_20171;
wire v_20172;
wire v_20173;
wire v_20174;
wire v_20175;
wire v_20176;
wire v_20177;
wire v_20178;
wire v_20179;
wire v_20180;
wire v_20181;
wire v_20182;
wire v_20183;
wire v_20184;
wire v_20185;
wire v_20186;
wire v_20187;
wire v_20188;
wire v_20189;
wire v_20190;
wire v_20191;
wire v_20192;
wire v_20193;
wire v_20194;
wire v_20195;
wire v_20196;
wire v_20197;
wire v_20198;
wire v_20199;
wire v_20200;
wire v_20201;
wire v_20202;
wire v_20203;
wire v_20204;
wire v_20205;
wire v_20206;
wire v_20207;
wire v_20208;
wire v_20209;
wire v_20210;
wire v_20211;
wire v_20212;
wire v_20213;
wire v_20214;
wire v_20215;
wire v_20216;
wire v_20217;
wire v_20218;
wire v_20219;
wire v_20220;
wire v_20221;
wire v_20222;
wire v_20223;
wire v_20224;
wire v_20225;
wire v_20226;
wire v_20227;
wire v_20228;
wire v_20229;
wire v_20230;
wire v_20231;
wire v_20232;
wire v_20233;
wire v_20234;
wire v_20235;
wire v_20236;
wire v_20237;
wire v_20238;
wire v_20239;
wire v_20240;
wire v_20241;
wire v_20242;
wire v_20243;
wire v_20244;
wire v_20245;
wire v_20246;
wire v_20247;
wire v_20248;
wire v_20249;
wire v_20250;
wire v_20251;
wire v_20252;
wire v_20253;
wire v_20254;
wire v_20255;
wire v_20256;
wire v_20257;
wire v_20258;
wire v_20259;
wire v_20260;
wire v_20261;
wire v_20262;
wire v_20263;
wire v_20264;
wire v_20265;
wire v_20266;
wire v_20267;
wire v_20268;
wire v_20269;
wire v_20270;
wire v_20271;
wire v_20272;
wire v_20273;
wire v_20274;
wire v_20275;
wire v_20276;
wire v_20277;
wire v_20278;
wire v_20279;
wire v_20280;
wire v_20281;
wire v_20282;
wire v_20283;
wire v_20284;
wire v_20285;
wire v_20286;
wire v_20287;
wire v_20288;
wire v_20289;
wire v_20290;
wire v_20291;
wire v_20292;
wire v_20293;
wire v_20294;
wire v_20295;
wire v_20296;
wire v_20297;
wire v_20298;
wire v_20299;
wire v_20300;
wire v_20301;
wire v_20302;
wire v_20303;
wire v_20304;
wire v_20306;
wire v_20307;
wire v_20308;
wire v_20309;
wire v_20310;
wire v_20311;
wire v_20312;
wire v_20313;
wire v_20314;
wire v_20315;
wire v_20316;
wire v_20317;
wire v_20318;
wire v_20319;
wire v_20320;
wire v_20321;
wire v_20322;
wire v_20323;
wire v_20324;
wire v_20325;
wire v_20326;
wire v_20327;
wire v_20328;
wire v_20329;
wire v_20330;
wire v_20331;
wire v_20332;
wire v_20333;
wire v_20334;
wire v_20335;
wire v_20336;
wire v_20337;
wire v_20338;
wire v_20339;
wire v_20340;
wire v_20341;
wire v_20342;
wire v_20343;
wire v_20344;
wire v_20345;
wire v_20346;
wire v_20347;
wire v_20348;
wire v_20349;
wire v_20350;
wire v_20351;
wire v_20352;
wire v_20353;
wire v_20354;
wire v_20355;
wire v_20356;
wire v_20357;
wire v_20358;
wire v_20359;
wire v_20360;
wire v_20361;
wire v_20362;
wire v_20363;
wire v_20364;
wire v_20365;
wire v_20366;
wire v_20367;
wire v_20368;
wire v_20369;
wire v_20370;
wire v_20371;
wire v_20372;
wire v_20373;
wire v_20374;
wire v_20375;
wire v_20376;
wire v_20377;
wire v_20378;
wire v_20379;
wire v_20380;
wire v_20381;
wire v_20382;
wire v_20383;
wire v_20384;
wire v_20385;
wire v_20386;
wire v_20387;
wire v_20388;
wire v_20389;
wire v_20390;
wire v_20391;
wire v_20392;
wire v_20393;
wire v_20394;
wire v_20395;
wire v_20396;
wire v_20397;
wire v_20398;
wire v_20399;
wire v_20400;
wire v_20401;
wire v_20402;
wire v_20403;
wire v_20404;
wire v_20405;
wire v_20406;
wire v_20407;
wire v_20408;
wire v_20409;
wire v_20410;
wire v_20411;
wire v_20412;
wire v_20413;
wire v_20414;
wire v_20415;
wire v_20416;
wire v_20417;
wire v_20418;
wire v_20419;
wire v_20420;
wire v_20421;
wire v_20422;
wire v_20423;
wire v_20424;
wire v_20425;
wire v_20426;
wire v_20427;
wire v_20428;
wire v_20429;
wire v_20430;
wire v_20431;
wire v_20432;
wire v_20433;
wire v_20434;
wire v_20435;
wire v_20436;
wire v_20437;
wire v_20438;
wire v_20439;
wire v_20440;
wire v_20441;
wire v_20442;
wire v_20443;
wire v_20444;
wire v_20445;
wire v_20446;
wire v_20447;
wire v_20448;
wire v_20449;
wire v_20450;
wire v_20451;
wire v_20452;
wire v_20453;
wire v_20454;
wire v_20455;
wire v_20456;
wire v_20457;
wire v_20458;
wire v_20459;
wire v_20460;
wire v_20461;
wire v_20462;
wire v_20463;
wire v_20464;
wire v_20465;
wire v_20466;
wire v_20467;
wire v_20468;
wire v_20469;
wire v_20470;
wire v_20471;
wire v_20472;
wire v_20473;
wire v_20474;
wire v_20475;
wire v_20476;
wire v_20477;
wire v_20478;
wire v_20479;
wire v_20480;
wire v_20481;
wire v_20482;
wire v_20483;
wire v_20484;
wire v_20485;
wire v_20486;
wire v_20487;
wire v_20488;
wire v_20489;
wire v_20490;
wire v_20491;
wire v_20492;
wire v_20493;
wire v_20494;
wire v_20495;
wire v_20496;
wire v_20497;
wire v_20498;
wire v_20499;
wire v_20500;
wire v_20501;
wire v_20502;
wire v_20503;
wire v_20504;
wire v_20505;
wire v_20506;
wire v_20507;
wire v_20508;
wire v_20509;
wire v_20510;
wire v_20511;
wire v_20512;
wire v_20513;
wire v_20514;
wire v_20515;
wire v_20516;
wire v_20517;
wire v_20518;
wire v_20519;
wire v_20520;
wire v_20521;
wire v_20522;
wire v_20523;
wire v_20524;
wire v_20525;
wire v_20526;
wire v_20527;
wire v_20528;
wire v_20529;
wire v_20530;
wire v_20531;
wire v_20532;
wire v_20533;
wire v_20534;
wire v_20535;
wire v_20536;
wire v_20537;
wire v_20538;
wire v_20539;
wire v_20540;
wire v_20541;
wire v_20542;
wire v_20543;
wire v_20544;
wire v_20545;
wire v_20546;
wire v_20547;
wire v_20549;
wire v_20550;
wire v_20551;
wire v_20552;
wire v_20553;
wire v_20554;
wire v_20555;
wire v_20556;
wire v_20557;
wire v_20558;
wire v_20559;
wire v_20560;
wire v_20561;
wire v_20562;
wire v_20563;
wire v_20564;
wire v_20565;
wire v_20566;
wire v_20567;
wire v_20568;
wire v_20569;
wire v_20570;
wire v_20571;
wire v_20572;
wire v_20573;
wire v_20574;
wire v_20575;
wire v_20576;
wire v_20577;
wire v_20578;
wire v_20579;
wire v_20580;
wire v_20581;
wire v_20582;
wire v_20583;
wire v_20584;
wire v_20585;
wire v_20586;
wire v_20587;
wire v_20588;
wire v_20589;
wire v_20590;
wire v_20591;
wire v_20592;
wire v_20593;
wire v_20594;
wire v_20595;
wire v_20596;
wire v_20597;
wire v_20598;
wire v_20599;
wire v_20600;
wire v_20601;
wire v_20602;
wire v_20603;
wire v_20604;
wire v_20605;
wire v_20606;
wire v_20607;
wire v_20608;
wire v_20609;
wire v_20610;
wire v_20611;
wire v_20612;
wire v_20613;
wire v_20614;
wire v_20615;
wire v_20616;
wire v_20617;
wire v_20618;
wire v_20619;
wire v_20620;
wire v_20621;
wire v_20622;
wire v_20623;
wire v_20624;
wire v_20625;
wire v_20626;
wire v_20627;
wire v_20628;
wire v_20629;
wire v_20630;
wire v_20631;
wire v_20632;
wire v_20633;
wire v_20634;
wire v_20635;
wire v_20636;
wire v_20637;
wire v_20638;
wire v_20639;
wire v_20640;
wire v_20641;
wire v_20642;
wire v_20643;
wire v_20644;
wire v_20645;
wire v_20646;
wire v_20647;
wire v_20648;
wire v_20649;
wire v_20650;
wire v_20651;
wire v_20652;
wire v_20653;
wire v_20654;
wire v_20655;
wire v_20656;
wire v_20657;
wire v_20658;
wire v_20659;
wire v_20660;
wire v_20661;
wire v_20662;
wire v_20663;
wire v_20664;
wire v_20665;
wire v_20666;
wire v_20667;
wire v_20668;
wire v_20669;
wire v_20670;
wire v_20671;
wire v_20672;
wire v_20673;
wire v_20674;
wire v_20675;
wire v_20676;
wire v_20677;
wire v_20678;
wire v_20679;
wire v_20680;
wire v_20681;
wire v_20682;
wire v_20683;
wire v_20684;
wire v_20685;
wire v_20686;
wire v_20687;
wire v_20688;
wire v_20689;
wire v_20690;
wire v_20691;
wire v_20692;
wire v_20693;
wire v_20694;
wire v_20695;
wire v_20696;
wire v_20697;
wire v_20698;
wire v_20699;
wire v_20700;
wire v_20701;
wire v_20702;
wire v_20703;
wire v_20704;
wire v_20705;
wire v_20706;
wire v_20707;
wire v_20708;
wire v_20709;
wire v_20710;
wire v_20711;
wire v_20712;
wire v_20713;
wire v_20714;
wire v_20715;
wire v_20716;
wire v_20717;
wire v_20718;
wire v_20719;
wire v_20720;
wire v_20721;
wire v_20722;
wire v_20723;
wire v_20724;
wire v_20725;
wire v_20726;
wire v_20727;
wire v_20728;
wire v_20729;
wire v_20730;
wire v_20731;
wire v_20732;
wire v_20733;
wire v_20734;
wire v_20735;
wire v_20736;
wire v_20737;
wire v_20738;
wire v_20739;
wire v_20740;
wire v_20741;
wire v_20742;
wire v_20743;
wire v_20744;
wire v_20745;
wire v_20746;
wire v_20747;
wire v_20748;
wire v_20749;
wire v_20750;
wire v_20751;
wire v_20752;
wire v_20753;
wire v_20754;
wire v_20755;
wire v_20756;
wire v_20757;
wire v_20758;
wire v_20759;
wire v_20760;
wire v_20761;
wire v_20762;
wire v_20763;
wire v_20764;
wire v_20765;
wire v_20766;
wire v_20767;
wire v_20768;
wire v_20769;
wire v_20770;
wire v_20771;
wire v_20772;
wire v_20773;
wire v_20774;
wire v_20775;
wire v_20776;
wire v_20777;
wire v_20778;
wire v_20779;
wire v_20780;
wire v_20781;
wire v_20782;
wire v_20783;
wire v_20784;
wire v_20785;
wire v_20786;
wire v_20787;
wire v_20788;
wire v_20789;
wire v_20790;
wire v_20791;
wire v_20792;
wire v_20793;
wire v_20794;
wire v_20795;
wire v_20796;
wire v_20797;
wire v_20798;
wire v_20799;
wire v_20800;
wire v_20801;
wire v_20802;
wire v_20803;
wire v_20804;
wire v_20805;
wire v_20806;
wire v_20807;
wire v_20808;
wire v_20809;
wire v_20810;
wire v_20811;
wire v_20812;
wire v_20813;
wire v_20814;
wire v_20815;
wire v_20816;
wire v_20817;
wire v_20818;
wire v_20819;
wire v_20820;
wire v_20821;
wire v_20822;
wire v_20823;
wire v_20824;
wire v_20825;
wire v_20826;
wire v_20827;
wire v_20828;
wire v_20829;
wire v_20830;
wire v_20831;
wire v_20832;
wire v_20833;
wire v_20834;
wire v_20835;
wire v_20836;
wire v_20837;
wire v_20838;
wire v_20839;
wire v_20840;
wire v_20841;
wire v_20842;
wire v_20843;
wire v_20844;
wire v_20845;
wire v_20846;
wire v_20847;
wire v_20848;
wire v_20849;
wire v_20850;
wire v_20851;
wire v_20852;
wire v_20853;
wire v_20854;
wire v_20855;
wire v_20856;
wire v_20857;
wire v_20858;
wire v_20859;
wire v_20860;
wire v_20861;
wire v_20862;
wire v_20863;
wire v_20864;
wire v_20865;
wire v_20866;
wire v_20867;
wire v_20868;
wire v_20869;
wire v_20870;
wire v_20871;
wire v_20872;
wire v_20873;
wire v_20874;
wire v_20875;
wire v_20876;
wire v_20877;
wire v_20878;
wire v_20879;
wire v_20880;
wire v_20881;
wire v_20882;
wire v_20883;
wire v_20884;
wire v_20885;
wire v_20886;
wire v_20887;
wire v_20888;
wire v_20889;
wire v_20890;
wire v_20891;
wire v_20892;
wire v_20893;
wire v_20894;
wire v_20895;
wire v_20896;
wire v_20897;
wire v_20898;
wire v_20899;
wire v_20900;
wire v_20901;
wire v_20902;
wire v_20903;
wire v_20904;
wire v_20905;
wire v_20906;
wire v_20907;
wire v_20908;
wire v_20909;
wire v_20910;
wire v_20911;
wire v_20912;
wire v_20913;
wire v_20914;
wire v_20915;
wire v_20916;
wire v_20917;
wire v_20918;
wire v_20919;
wire v_20920;
wire v_20921;
wire v_20922;
wire v_20923;
wire v_20924;
wire v_20925;
wire v_20926;
wire v_20927;
wire v_20928;
wire v_20929;
wire v_20930;
wire v_20931;
wire v_20932;
wire v_20933;
wire v_20934;
wire v_20935;
wire v_20936;
wire v_20937;
wire v_20938;
wire v_20939;
wire v_20941;
wire v_20942;
wire v_20943;
wire v_20944;
wire v_20945;
wire v_20946;
wire v_20947;
wire v_20948;
wire v_20949;
wire v_20950;
wire v_20951;
wire v_20952;
wire v_20953;
wire v_20954;
wire v_20955;
wire v_20956;
wire v_20957;
wire v_20958;
wire v_20959;
wire v_20960;
wire v_20961;
wire v_20962;
wire v_20963;
wire v_20964;
wire v_20965;
wire v_20966;
wire v_20967;
wire v_20968;
wire v_20969;
wire v_20970;
wire v_20971;
wire v_20972;
wire v_20973;
wire v_20974;
wire v_20975;
wire v_20976;
wire v_20977;
wire v_20978;
wire v_20979;
wire v_20980;
wire v_20981;
wire v_20982;
wire v_20983;
wire v_20984;
wire v_20985;
wire v_20986;
wire v_20987;
wire v_20988;
wire v_20989;
wire v_20990;
wire v_20991;
wire v_20992;
wire v_20993;
wire v_20994;
wire v_20995;
wire v_20996;
wire v_20997;
wire v_20998;
wire v_20999;
wire v_21000;
wire v_21001;
wire v_21002;
wire v_21003;
wire v_21004;
wire v_21005;
wire v_21006;
wire v_21007;
wire v_21008;
wire v_21009;
wire v_21010;
wire v_21011;
wire v_21012;
wire v_21013;
wire v_21014;
wire v_21015;
wire v_21016;
wire v_21017;
wire v_21018;
wire v_21019;
wire v_21020;
wire v_21021;
wire v_21022;
wire v_21023;
wire v_21024;
wire v_21025;
wire v_21026;
wire v_21027;
wire v_21028;
wire v_21029;
wire v_21030;
wire v_21031;
wire v_21032;
wire v_21033;
wire v_21035;
wire v_21037;
wire v_21038;
wire v_21039;
wire v_21041;
wire v_21042;
wire v_21043;
wire v_21045;
wire v_21046;
wire v_21047;
wire v_21049;
wire v_21050;
wire v_21052;
wire v_21053;
wire v_21054;
wire v_21056;
wire v_21057;
wire v_21058;
wire v_21060;
wire v_21061;
wire v_21062;
wire v_21064;
wire v_21065;
wire v_21066;
wire v_21068;
wire v_21069;
wire v_21070;
wire v_21072;
wire v_21073;
wire v_21074;
wire v_21076;
wire v_21077;
wire v_21078;
wire v_21080;
wire v_21081;
wire v_21082;
wire v_21084;
wire v_21085;
wire v_21086;
wire v_21088;
wire v_21089;
wire v_21090;
wire v_21092;
wire v_21093;
wire v_21094;
wire v_21096;
wire v_21097;
wire v_21098;
wire v_21100;
wire v_21101;
wire v_21102;
wire v_21103;
wire v_21104;
wire v_21105;
wire v_21106;
wire v_21107;
wire v_21108;
wire v_21109;
wire v_21110;
wire v_21111;
wire v_21112;
wire v_21113;
wire v_21114;
wire v_21115;
wire v_21116;
wire v_21117;
wire v_21118;
wire v_21119;
wire v_21120;
wire v_21121;
wire v_21122;
wire v_21123;
wire v_21124;
wire v_21125;
wire v_21126;
wire v_21127;
wire v_21128;
wire v_21129;
wire v_21130;
wire v_21131;
wire v_21132;
wire v_21133;
wire v_21134;
wire v_21135;
wire v_21136;
wire v_21137;
wire v_21138;
wire v_21139;
wire v_21140;
wire v_21141;
wire v_21142;
wire v_21143;
wire v_21144;
wire v_21145;
wire v_21146;
wire v_21147;
wire v_21148;
wire v_21149;
wire v_21150;
wire v_21151;
wire v_21152;
wire v_21153;
wire v_21154;
wire v_21155;
wire v_21156;
wire v_21157;
wire v_21158;
wire v_21159;
wire v_21160;
wire v_21161;
wire v_21162;
wire v_21163;
wire v_21164;
wire v_21165;
wire v_21166;
wire v_21167;
wire v_21168;
wire v_21169;
wire v_21170;
wire v_21171;
wire v_21172;
wire v_21173;
wire v_21174;
wire v_21175;
wire v_21176;
wire v_21177;
wire v_21178;
wire v_21179;
wire v_21180;
wire v_21181;
wire v_21182;
wire v_21183;
wire v_21184;
wire v_21185;
wire v_21186;
wire v_21187;
wire v_21188;
wire v_21189;
wire v_21190;
wire v_21191;
wire v_21192;
wire v_21193;
wire v_21194;
wire v_21195;
wire v_21196;
wire v_21197;
wire v_21198;
wire v_21199;
wire v_21200;
wire v_21201;
wire v_21202;
wire v_21203;
wire v_21204;
wire v_21205;
wire v_21206;
wire v_21207;
wire v_21208;
wire v_21209;
wire v_21210;
wire v_21211;
wire v_21212;
wire v_21213;
wire v_21214;
wire v_21215;
wire v_21216;
wire v_21217;
wire v_21218;
wire v_21219;
wire v_21220;
wire v_21221;
wire v_21222;
wire v_21223;
wire v_21224;
wire v_21225;
wire v_21226;
wire v_21227;
wire v_21228;
wire v_21229;
wire v_21230;
wire v_21231;
wire v_21232;
wire v_21233;
wire v_21234;
wire v_21235;
wire v_21236;
wire v_21237;
wire v_21238;
wire v_21239;
wire v_21240;
wire v_21241;
wire v_21242;
wire v_21243;
wire v_21244;
wire v_21245;
wire v_21246;
wire v_21247;
wire v_21248;
wire v_21249;
wire v_21250;
wire v_21251;
wire v_21252;
wire v_21253;
wire v_21254;
wire v_21255;
wire v_21256;
wire v_21257;
wire v_21258;
wire v_21259;
wire v_21260;
wire v_21261;
wire v_21262;
wire v_21263;
wire v_21264;
wire v_21265;
wire v_21266;
wire v_21267;
wire v_21268;
wire v_21269;
wire v_21270;
wire v_21271;
wire v_21272;
wire v_21273;
wire v_21274;
wire v_21275;
wire v_21276;
wire v_21277;
wire v_21278;
wire v_21279;
wire v_21280;
wire v_21281;
wire v_21282;
wire v_21283;
wire v_21284;
wire v_21285;
wire v_21286;
wire v_21287;
wire v_21288;
wire v_21289;
wire v_21290;
wire v_21291;
wire v_21292;
wire v_21293;
wire v_21295;
wire v_21296;
wire v_21297;
wire v_21298;
wire v_21299;
wire v_21300;
wire v_21301;
wire v_21302;
wire v_21303;
wire v_21304;
wire v_21305;
wire v_21306;
wire v_21307;
wire v_21308;
wire v_21309;
wire v_21310;
wire v_21311;
wire v_21312;
wire v_21313;
wire v_21314;
wire v_21315;
wire v_21316;
wire v_21317;
wire v_21318;
wire v_21319;
wire v_21320;
wire v_21321;
wire v_21322;
wire v_21323;
wire v_21324;
wire v_21325;
wire v_21326;
wire v_21327;
wire v_21328;
wire v_21329;
wire v_21330;
wire v_21331;
wire v_21332;
wire v_21333;
wire v_21334;
wire v_21335;
wire v_21336;
wire v_21337;
wire v_21338;
wire v_21339;
wire v_21340;
wire v_21341;
wire v_21342;
wire v_21343;
wire v_21344;
wire v_21345;
wire v_21346;
wire v_21347;
wire v_21348;
wire v_21349;
wire v_21350;
wire v_21351;
wire v_21352;
wire v_21353;
wire v_21354;
wire v_21355;
wire v_21356;
wire v_21357;
wire v_21358;
wire v_21359;
wire v_21360;
wire v_21361;
wire v_21362;
wire v_21363;
wire v_21364;
wire v_21365;
wire v_21366;
wire v_21367;
wire v_21368;
wire v_21369;
wire v_21370;
wire v_21371;
wire v_21372;
wire v_21373;
wire v_21374;
wire v_21375;
wire v_21376;
wire v_21377;
wire v_21378;
wire v_21379;
wire v_21380;
wire v_21381;
wire v_21382;
wire v_21383;
wire v_21384;
wire v_21385;
wire v_21386;
wire v_21387;
wire v_21388;
wire v_21389;
wire v_21390;
wire v_21391;
wire v_21392;
wire v_21393;
wire v_21394;
wire v_21395;
wire v_21396;
wire v_21397;
wire v_21398;
wire v_21399;
wire v_21400;
wire v_21401;
wire v_21402;
wire v_21403;
wire v_21404;
wire v_21405;
wire v_21406;
wire v_21407;
wire v_21408;
wire v_21409;
wire v_21410;
wire v_21411;
wire v_21412;
wire v_21413;
wire v_21414;
wire v_21415;
wire v_21416;
wire v_21417;
wire v_21418;
wire v_21419;
wire v_21420;
wire v_21421;
wire v_21422;
wire v_21423;
wire v_21424;
wire v_21425;
wire v_21426;
wire v_21427;
wire v_21428;
wire v_21429;
wire v_21430;
wire v_21431;
wire v_21432;
wire v_21433;
wire v_21434;
wire v_21435;
wire v_21436;
wire v_21437;
wire v_21438;
wire v_21439;
wire v_21440;
wire v_21441;
wire v_21442;
wire v_21443;
wire v_21444;
wire v_21445;
wire v_21446;
wire v_21447;
wire v_21448;
wire v_21449;
wire v_21450;
wire v_21451;
wire v_21452;
wire v_21453;
wire v_21454;
wire v_21455;
wire v_21456;
wire v_21457;
wire v_21458;
wire v_21459;
wire v_21460;
wire v_21461;
wire v_21462;
wire v_21463;
wire v_21464;
wire v_21465;
wire v_21466;
wire v_21467;
wire v_21468;
wire v_21469;
wire v_21470;
wire v_21471;
wire v_21472;
wire v_21473;
wire v_21474;
wire v_21475;
wire v_21476;
wire v_21477;
wire v_21478;
wire v_21479;
wire v_21480;
wire v_21481;
wire v_21482;
wire v_21483;
wire v_21484;
wire v_21485;
wire v_21486;
wire v_21487;
wire v_21488;
wire v_21489;
wire v_21490;
wire v_21491;
wire v_21492;
wire v_21493;
wire v_21494;
wire v_21495;
wire v_21496;
wire v_21497;
wire v_21498;
wire v_21499;
wire v_21500;
wire v_21501;
wire v_21502;
wire v_21503;
wire v_21504;
wire v_21505;
wire v_21506;
wire v_21507;
wire v_21508;
wire v_21509;
wire v_21510;
wire v_21511;
wire v_21512;
wire v_21513;
wire v_21514;
wire v_21515;
wire v_21516;
wire v_21517;
wire v_21518;
wire v_21519;
wire v_21520;
wire v_21521;
wire v_21522;
wire v_21523;
wire v_21524;
wire v_21525;
wire v_21526;
wire v_21527;
wire v_21528;
wire v_21529;
wire v_21530;
wire v_21531;
wire v_21532;
wire v_21533;
wire v_21534;
wire v_21535;
wire v_21536;
wire v_21538;
wire v_21539;
wire v_21540;
wire v_21541;
wire v_21542;
wire v_21543;
wire v_21544;
wire v_21545;
wire v_21546;
wire v_21547;
wire v_21548;
wire v_21549;
wire v_21550;
wire v_21551;
wire v_21552;
wire v_21553;
wire v_21554;
wire v_21555;
wire v_21556;
wire v_21557;
wire v_21558;
wire v_21559;
wire v_21560;
wire v_21561;
wire v_21562;
wire v_21563;
wire v_21564;
wire v_21565;
wire v_21566;
wire v_21567;
wire v_21568;
wire v_21569;
wire v_21570;
wire v_21571;
wire v_21572;
wire v_21573;
wire v_21574;
wire v_21575;
wire v_21576;
wire v_21577;
wire v_21578;
wire v_21579;
wire v_21580;
wire v_21581;
wire v_21582;
wire v_21583;
wire v_21584;
wire v_21585;
wire v_21586;
wire v_21587;
wire v_21588;
wire v_21589;
wire v_21590;
wire v_21591;
wire v_21592;
wire v_21593;
wire v_21594;
wire v_21595;
wire v_21596;
wire v_21597;
wire v_21598;
wire v_21599;
wire v_21600;
wire v_21601;
wire v_21602;
wire v_21603;
wire v_21604;
wire v_21605;
wire v_21606;
wire v_21607;
wire v_21608;
wire v_21609;
wire v_21610;
wire v_21611;
wire v_21612;
wire v_21613;
wire v_21614;
wire v_21615;
wire v_21616;
wire v_21617;
wire v_21618;
wire v_21619;
wire v_21620;
wire v_21621;
wire v_21622;
wire v_21623;
wire v_21624;
wire v_21625;
wire v_21626;
wire v_21627;
wire v_21628;
wire v_21629;
wire v_21630;
wire v_21631;
wire v_21632;
wire v_21633;
wire v_21634;
wire v_21635;
wire v_21636;
wire v_21637;
wire v_21638;
wire v_21639;
wire v_21640;
wire v_21641;
wire v_21642;
wire v_21643;
wire v_21644;
wire v_21645;
wire v_21646;
wire v_21647;
wire v_21648;
wire v_21649;
wire v_21650;
wire v_21651;
wire v_21652;
wire v_21653;
wire v_21654;
wire v_21655;
wire v_21656;
wire v_21657;
wire v_21658;
wire v_21659;
wire v_21660;
wire v_21661;
wire v_21662;
wire v_21663;
wire v_21664;
wire v_21665;
wire v_21666;
wire v_21667;
wire v_21668;
wire v_21669;
wire v_21670;
wire v_21671;
wire v_21672;
wire v_21673;
wire v_21674;
wire v_21675;
wire v_21676;
wire v_21677;
wire v_21678;
wire v_21679;
wire v_21680;
wire v_21681;
wire v_21682;
wire v_21683;
wire v_21684;
wire v_21685;
wire v_21686;
wire v_21687;
wire v_21688;
wire v_21689;
wire v_21690;
wire v_21691;
wire v_21692;
wire v_21693;
wire v_21694;
wire v_21695;
wire v_21696;
wire v_21697;
wire v_21698;
wire v_21699;
wire v_21700;
wire v_21701;
wire v_21702;
wire v_21703;
wire v_21704;
wire v_21705;
wire v_21706;
wire v_21707;
wire v_21708;
wire v_21709;
wire v_21710;
wire v_21711;
wire v_21712;
wire v_21713;
wire v_21714;
wire v_21715;
wire v_21716;
wire v_21717;
wire v_21718;
wire v_21719;
wire v_21720;
wire v_21721;
wire v_21722;
wire v_21723;
wire v_21724;
wire v_21725;
wire v_21726;
wire v_21727;
wire v_21728;
wire v_21729;
wire v_21730;
wire v_21731;
wire v_21732;
wire v_21733;
wire v_21734;
wire v_21735;
wire v_21736;
wire v_21737;
wire v_21738;
wire v_21739;
wire v_21740;
wire v_21741;
wire v_21742;
wire v_21743;
wire v_21744;
wire v_21745;
wire v_21746;
wire v_21747;
wire v_21748;
wire v_21749;
wire v_21750;
wire v_21751;
wire v_21752;
wire v_21753;
wire v_21754;
wire v_21755;
wire v_21756;
wire v_21757;
wire v_21758;
wire v_21759;
wire v_21760;
wire v_21761;
wire v_21762;
wire v_21763;
wire v_21764;
wire v_21765;
wire v_21766;
wire v_21767;
wire v_21768;
wire v_21769;
wire v_21770;
wire v_21771;
wire v_21772;
wire v_21773;
wire v_21774;
wire v_21775;
wire v_21776;
wire v_21777;
wire v_21778;
wire v_21779;
wire v_21781;
wire v_21782;
wire v_21783;
wire v_21784;
wire v_21785;
wire v_21786;
wire v_21787;
wire v_21788;
wire v_21789;
wire v_21790;
wire v_21791;
wire v_21792;
wire v_21793;
wire v_21794;
wire v_21795;
wire v_21796;
wire v_21797;
wire v_21798;
wire v_21799;
wire v_21800;
wire v_21801;
wire v_21802;
wire v_21803;
wire v_21804;
wire v_21805;
wire v_21806;
wire v_21807;
wire v_21808;
wire v_21809;
wire v_21810;
wire v_21811;
wire v_21812;
wire v_21813;
wire v_21814;
wire v_21815;
wire v_21816;
wire v_21817;
wire v_21818;
wire v_21819;
wire v_21820;
wire v_21821;
wire v_21822;
wire v_21823;
wire v_21824;
wire v_21825;
wire v_21826;
wire v_21827;
wire v_21828;
wire v_21829;
wire v_21830;
wire v_21831;
wire v_21832;
wire v_21833;
wire v_21834;
wire v_21835;
wire v_21836;
wire v_21837;
wire v_21838;
wire v_21839;
wire v_21840;
wire v_21841;
wire v_21842;
wire v_21843;
wire v_21844;
wire v_21845;
wire v_21846;
wire v_21847;
wire v_21848;
wire v_21849;
wire v_21850;
wire v_21851;
wire v_21852;
wire v_21853;
wire v_21854;
wire v_21855;
wire v_21856;
wire v_21857;
wire v_21858;
wire v_21859;
wire v_21860;
wire v_21861;
wire v_21862;
wire v_21863;
wire v_21864;
wire v_21865;
wire v_21866;
wire v_21867;
wire v_21868;
wire v_21869;
wire v_21870;
wire v_21871;
wire v_21872;
wire v_21873;
wire v_21874;
wire v_21875;
wire v_21876;
wire v_21877;
wire v_21878;
wire v_21879;
wire v_21880;
wire v_21881;
wire v_21882;
wire v_21883;
wire v_21884;
wire v_21885;
wire v_21886;
wire v_21887;
wire v_21888;
wire v_21889;
wire v_21890;
wire v_21891;
wire v_21892;
wire v_21893;
wire v_21894;
wire v_21895;
wire v_21896;
wire v_21897;
wire v_21898;
wire v_21899;
wire v_21900;
wire v_21901;
wire v_21902;
wire v_21903;
wire v_21904;
wire v_21905;
wire v_21906;
wire v_21907;
wire v_21908;
wire v_21909;
wire v_21910;
wire v_21911;
wire v_21912;
wire v_21913;
wire v_21914;
wire v_21915;
wire v_21916;
wire v_21917;
wire v_21918;
wire v_21919;
wire v_21920;
wire v_21921;
wire v_21922;
wire v_21923;
wire v_21924;
wire v_21925;
wire v_21926;
wire v_21927;
wire v_21928;
wire v_21929;
wire v_21930;
wire v_21931;
wire v_21932;
wire v_21933;
wire v_21934;
wire v_21935;
wire v_21936;
wire v_21937;
wire v_21938;
wire v_21939;
wire v_21940;
wire v_21941;
wire v_21942;
wire v_21943;
wire v_21944;
wire v_21945;
wire v_21946;
wire v_21947;
wire v_21948;
wire v_21949;
wire v_21950;
wire v_21951;
wire v_21952;
wire v_21953;
wire v_21954;
wire v_21955;
wire v_21956;
wire v_21957;
wire v_21958;
wire v_21959;
wire v_21960;
wire v_21961;
wire v_21962;
wire v_21963;
wire v_21964;
wire v_21965;
wire v_21966;
wire v_21967;
wire v_21968;
wire v_21969;
wire v_21970;
wire v_21971;
wire v_21972;
wire v_21973;
wire v_21974;
wire v_21975;
wire v_21976;
wire v_21977;
wire v_21978;
wire v_21979;
wire v_21980;
wire v_21981;
wire v_21982;
wire v_21983;
wire v_21984;
wire v_21985;
wire v_21986;
wire v_21987;
wire v_21988;
wire v_21989;
wire v_21990;
wire v_21991;
wire v_21992;
wire v_21993;
wire v_21994;
wire v_21995;
wire v_21996;
wire v_21997;
wire v_21998;
wire v_21999;
wire v_22000;
wire v_22001;
wire v_22002;
wire v_22003;
wire v_22004;
wire v_22005;
wire v_22006;
wire v_22007;
wire v_22008;
wire v_22009;
wire v_22010;
wire v_22011;
wire v_22012;
wire v_22013;
wire v_22014;
wire v_22015;
wire v_22016;
wire v_22017;
wire v_22018;
wire v_22019;
wire v_22020;
wire v_22021;
wire v_22022;
wire v_22024;
wire v_22025;
wire v_22026;
wire v_22027;
wire v_22028;
wire v_22029;
wire v_22030;
wire v_22031;
wire v_22032;
wire v_22033;
wire v_22034;
wire v_22035;
wire v_22036;
wire v_22037;
wire v_22038;
wire v_22039;
wire v_22040;
wire v_22041;
wire v_22042;
wire v_22043;
wire v_22044;
wire v_22045;
wire v_22046;
wire v_22047;
wire v_22048;
wire v_22049;
wire v_22050;
wire v_22051;
wire v_22052;
wire v_22053;
wire v_22054;
wire v_22055;
wire v_22056;
wire v_22057;
wire v_22058;
wire v_22059;
wire v_22060;
wire v_22061;
wire v_22062;
wire v_22063;
wire v_22064;
wire v_22065;
wire v_22066;
wire v_22067;
wire v_22068;
wire v_22069;
wire v_22070;
wire v_22071;
wire v_22072;
wire v_22073;
wire v_22074;
wire v_22075;
wire v_22076;
wire v_22077;
wire v_22078;
wire v_22079;
wire v_22080;
wire v_22081;
wire v_22082;
wire v_22083;
wire v_22084;
wire v_22085;
wire v_22086;
wire v_22087;
wire v_22088;
wire v_22089;
wire v_22090;
wire v_22091;
wire v_22092;
wire v_22093;
wire v_22094;
wire v_22095;
wire v_22096;
wire v_22097;
wire v_22098;
wire v_22099;
wire v_22100;
wire v_22101;
wire v_22102;
wire v_22103;
wire v_22104;
wire v_22105;
wire v_22106;
wire v_22107;
wire v_22108;
wire v_22109;
wire v_22110;
wire v_22111;
wire v_22112;
wire v_22113;
wire v_22114;
wire v_22115;
wire v_22116;
wire v_22117;
wire v_22118;
wire v_22119;
wire v_22120;
wire v_22121;
wire v_22122;
wire v_22123;
wire v_22124;
wire v_22125;
wire v_22126;
wire v_22127;
wire v_22128;
wire v_22129;
wire v_22130;
wire v_22131;
wire v_22132;
wire v_22133;
wire v_22134;
wire v_22135;
wire v_22136;
wire v_22137;
wire v_22138;
wire v_22139;
wire v_22140;
wire v_22141;
wire v_22142;
wire v_22143;
wire v_22144;
wire v_22145;
wire v_22146;
wire v_22147;
wire v_22148;
wire v_22149;
wire v_22150;
wire v_22151;
wire v_22152;
wire v_22153;
wire v_22154;
wire v_22155;
wire v_22156;
wire v_22157;
wire v_22158;
wire v_22159;
wire v_22160;
wire v_22161;
wire v_22162;
wire v_22163;
wire v_22164;
wire v_22165;
wire v_22166;
wire v_22167;
wire v_22168;
wire v_22169;
wire v_22170;
wire v_22171;
wire v_22172;
wire v_22173;
wire v_22174;
wire v_22175;
wire v_22176;
wire v_22177;
wire v_22178;
wire v_22179;
wire v_22180;
wire v_22181;
wire v_22182;
wire v_22183;
wire v_22184;
wire v_22185;
wire v_22186;
wire v_22187;
wire v_22188;
wire v_22189;
wire v_22190;
wire v_22191;
wire v_22192;
wire v_22193;
wire v_22194;
wire v_22195;
wire v_22196;
wire v_22197;
wire v_22198;
wire v_22199;
wire v_22200;
wire v_22201;
wire v_22202;
wire v_22203;
wire v_22204;
wire v_22205;
wire v_22206;
wire v_22207;
wire v_22208;
wire v_22209;
wire v_22210;
wire v_22211;
wire v_22212;
wire v_22213;
wire v_22214;
wire v_22215;
wire v_22216;
wire v_22217;
wire v_22218;
wire v_22219;
wire v_22220;
wire v_22221;
wire v_22222;
wire v_22223;
wire v_22224;
wire v_22225;
wire v_22226;
wire v_22227;
wire v_22228;
wire v_22229;
wire v_22230;
wire v_22231;
wire v_22232;
wire v_22233;
wire v_22234;
wire v_22235;
wire v_22236;
wire v_22237;
wire v_22238;
wire v_22239;
wire v_22240;
wire v_22241;
wire v_22242;
wire v_22243;
wire v_22244;
wire v_22245;
wire v_22246;
wire v_22247;
wire v_22248;
wire v_22249;
wire v_22250;
wire v_22251;
wire v_22252;
wire v_22253;
wire v_22254;
wire v_22255;
wire v_22256;
wire v_22257;
wire v_22258;
wire v_22259;
wire v_22260;
wire v_22261;
wire v_22262;
wire v_22263;
wire v_22264;
wire v_22265;
wire v_22267;
wire v_22268;
wire v_22269;
wire v_22270;
wire v_22271;
wire v_22272;
wire v_22273;
wire v_22274;
wire v_22275;
wire v_22276;
wire v_22277;
wire v_22278;
wire v_22279;
wire v_22280;
wire v_22281;
wire v_22282;
wire v_22283;
wire v_22284;
wire v_22285;
wire v_22286;
wire v_22287;
wire v_22288;
wire v_22289;
wire v_22290;
wire v_22291;
wire v_22292;
wire v_22293;
wire v_22294;
wire v_22295;
wire v_22296;
wire v_22297;
wire v_22298;
wire v_22299;
wire v_22300;
wire v_22301;
wire v_22302;
wire v_22303;
wire v_22304;
wire v_22305;
wire v_22306;
wire v_22307;
wire v_22308;
wire v_22309;
wire v_22310;
wire v_22311;
wire v_22312;
wire v_22313;
wire v_22314;
wire v_22315;
wire v_22316;
wire v_22317;
wire v_22318;
wire v_22319;
wire v_22320;
wire v_22321;
wire v_22322;
wire v_22323;
wire v_22324;
wire v_22325;
wire v_22326;
wire v_22327;
wire v_22328;
wire v_22329;
wire v_22330;
wire v_22331;
wire v_22332;
wire v_22333;
wire v_22334;
wire v_22335;
wire v_22336;
wire v_22337;
wire v_22338;
wire v_22339;
wire v_22340;
wire v_22341;
wire v_22342;
wire v_22343;
wire v_22344;
wire v_22345;
wire v_22346;
wire v_22347;
wire v_22348;
wire v_22349;
wire v_22350;
wire v_22351;
wire v_22352;
wire v_22353;
wire v_22354;
wire v_22355;
wire v_22356;
wire v_22357;
wire v_22358;
wire v_22359;
wire v_22360;
wire v_22361;
wire v_22362;
wire v_22363;
wire v_22364;
wire v_22365;
wire v_22366;
wire v_22367;
wire v_22368;
wire v_22369;
wire v_22370;
wire v_22371;
wire v_22372;
wire v_22373;
wire v_22374;
wire v_22375;
wire v_22376;
wire v_22377;
wire v_22378;
wire v_22379;
wire v_22380;
wire v_22381;
wire v_22382;
wire v_22383;
wire v_22384;
wire v_22385;
wire v_22386;
wire v_22387;
wire v_22388;
wire v_22389;
wire v_22390;
wire v_22391;
wire v_22392;
wire v_22393;
wire v_22394;
wire v_22395;
wire v_22396;
wire v_22397;
wire v_22398;
wire v_22399;
wire v_22400;
wire v_22401;
wire v_22402;
wire v_22403;
wire v_22404;
wire v_22405;
wire v_22406;
wire v_22407;
wire v_22408;
wire v_22409;
wire v_22410;
wire v_22411;
wire v_22412;
wire v_22413;
wire v_22414;
wire v_22415;
wire v_22416;
wire v_22417;
wire v_22418;
wire v_22419;
wire v_22420;
wire v_22421;
wire v_22422;
wire v_22423;
wire v_22424;
wire v_22425;
wire v_22426;
wire v_22427;
wire v_22428;
wire v_22429;
wire v_22430;
wire v_22431;
wire v_22432;
wire v_22433;
wire v_22434;
wire v_22435;
wire v_22436;
wire v_22437;
wire v_22438;
wire v_22439;
wire v_22440;
wire v_22441;
wire v_22442;
wire v_22443;
wire v_22444;
wire v_22445;
wire v_22446;
wire v_22447;
wire v_22448;
wire v_22449;
wire v_22450;
wire v_22451;
wire v_22452;
wire v_22453;
wire v_22454;
wire v_22455;
wire v_22456;
wire v_22457;
wire v_22458;
wire v_22459;
wire v_22460;
wire v_22461;
wire v_22462;
wire v_22463;
wire v_22464;
wire v_22465;
wire v_22466;
wire v_22467;
wire v_22468;
wire v_22469;
wire v_22470;
wire v_22471;
wire v_22472;
wire v_22473;
wire v_22474;
wire v_22475;
wire v_22476;
wire v_22477;
wire v_22478;
wire v_22479;
wire v_22480;
wire v_22481;
wire v_22482;
wire v_22483;
wire v_22484;
wire v_22485;
wire v_22486;
wire v_22487;
wire v_22488;
wire v_22489;
wire v_22490;
wire v_22491;
wire v_22492;
wire v_22493;
wire v_22494;
wire v_22495;
wire v_22496;
wire v_22497;
wire v_22498;
wire v_22499;
wire v_22500;
wire v_22501;
wire v_22502;
wire v_22503;
wire v_22504;
wire v_22505;
wire v_22506;
wire v_22507;
wire v_22508;
wire v_22510;
wire v_22511;
wire v_22512;
wire v_22513;
wire v_22514;
wire v_22515;
wire v_22516;
wire v_22517;
wire v_22518;
wire v_22519;
wire v_22520;
wire v_22521;
wire v_22522;
wire v_22523;
wire v_22524;
wire v_22525;
wire v_22526;
wire v_22527;
wire v_22528;
wire v_22529;
wire v_22530;
wire v_22531;
wire v_22532;
wire v_22533;
wire v_22534;
wire v_22535;
wire v_22536;
wire v_22537;
wire v_22538;
wire v_22539;
wire v_22540;
wire v_22541;
wire v_22542;
wire v_22543;
wire v_22544;
wire v_22545;
wire v_22546;
wire v_22547;
wire v_22548;
wire v_22549;
wire v_22550;
wire v_22551;
wire v_22552;
wire v_22553;
wire v_22554;
wire v_22555;
wire v_22556;
wire v_22557;
wire v_22558;
wire v_22559;
wire v_22560;
wire v_22561;
wire v_22562;
wire v_22563;
wire v_22564;
wire v_22565;
wire v_22566;
wire v_22567;
wire v_22568;
wire v_22569;
wire v_22570;
wire v_22571;
wire v_22572;
wire v_22573;
wire v_22574;
wire v_22575;
wire v_22576;
wire v_22577;
wire v_22578;
wire v_22579;
wire v_22580;
wire v_22581;
wire v_22582;
wire v_22583;
wire v_22584;
wire v_22585;
wire v_22586;
wire v_22587;
wire v_22588;
wire v_22589;
wire v_22590;
wire v_22591;
wire v_22592;
wire v_22593;
wire v_22594;
wire v_22595;
wire v_22596;
wire v_22597;
wire v_22598;
wire v_22599;
wire v_22600;
wire v_22601;
wire v_22602;
wire v_22603;
wire v_22604;
wire v_22605;
wire v_22606;
wire v_22607;
wire v_22608;
wire v_22609;
wire v_22610;
wire v_22611;
wire v_22612;
wire v_22613;
wire v_22614;
wire v_22615;
wire v_22616;
wire v_22617;
wire v_22618;
wire v_22619;
wire v_22620;
wire v_22621;
wire v_22622;
wire v_22623;
wire v_22624;
wire v_22625;
wire v_22626;
wire v_22627;
wire v_22628;
wire v_22629;
wire v_22630;
wire v_22631;
wire v_22632;
wire v_22633;
wire v_22634;
wire v_22635;
wire v_22636;
wire v_22637;
wire v_22638;
wire v_22639;
wire v_22640;
wire v_22641;
wire v_22642;
wire v_22643;
wire v_22644;
wire v_22645;
wire v_22646;
wire v_22647;
wire v_22648;
wire v_22649;
wire v_22650;
wire v_22651;
wire v_22652;
wire v_22653;
wire v_22654;
wire v_22655;
wire v_22656;
wire v_22657;
wire v_22658;
wire v_22659;
wire v_22660;
wire v_22661;
wire v_22662;
wire v_22663;
wire v_22664;
wire v_22665;
wire v_22666;
wire v_22667;
wire v_22668;
wire v_22669;
wire v_22670;
wire v_22671;
wire v_22672;
wire v_22673;
wire v_22674;
wire v_22675;
wire v_22676;
wire v_22677;
wire v_22678;
wire v_22679;
wire v_22680;
wire v_22681;
wire v_22682;
wire v_22683;
wire v_22684;
wire v_22685;
wire v_22686;
wire v_22687;
wire v_22688;
wire v_22689;
wire v_22690;
wire v_22691;
wire v_22692;
wire v_22693;
wire v_22694;
wire v_22695;
wire v_22696;
wire v_22697;
wire v_22698;
wire v_22699;
wire v_22700;
wire v_22701;
wire v_22702;
wire v_22703;
wire v_22704;
wire v_22705;
wire v_22706;
wire v_22707;
wire v_22708;
wire v_22709;
wire v_22710;
wire v_22711;
wire v_22712;
wire v_22713;
wire v_22714;
wire v_22715;
wire v_22716;
wire v_22717;
wire v_22718;
wire v_22719;
wire v_22720;
wire v_22721;
wire v_22722;
wire v_22723;
wire v_22724;
wire v_22725;
wire v_22726;
wire v_22727;
wire v_22728;
wire v_22729;
wire v_22730;
wire v_22731;
wire v_22732;
wire v_22733;
wire v_22734;
wire v_22735;
wire v_22736;
wire v_22737;
wire v_22738;
wire v_22739;
wire v_22740;
wire v_22741;
wire v_22742;
wire v_22743;
wire v_22744;
wire v_22745;
wire v_22746;
wire v_22747;
wire v_22748;
wire v_22749;
wire v_22750;
wire v_22751;
wire v_22753;
wire v_22754;
wire v_22755;
wire v_22756;
wire v_22757;
wire v_22758;
wire v_22759;
wire v_22760;
wire v_22761;
wire v_22762;
wire v_22763;
wire v_22764;
wire v_22765;
wire v_22766;
wire v_22767;
wire v_22768;
wire v_22769;
wire v_22770;
wire v_22771;
wire v_22772;
wire v_22773;
wire v_22774;
wire v_22775;
wire v_22776;
wire v_22777;
wire v_22778;
wire v_22779;
wire v_22780;
wire v_22781;
wire v_22782;
wire v_22783;
wire v_22784;
wire v_22785;
wire v_22786;
wire v_22787;
wire v_22788;
wire v_22789;
wire v_22790;
wire v_22791;
wire v_22792;
wire v_22793;
wire v_22794;
wire v_22795;
wire v_22796;
wire v_22797;
wire v_22798;
wire v_22799;
wire v_22800;
wire v_22801;
wire v_22802;
wire v_22803;
wire v_22804;
wire v_22805;
wire v_22806;
wire v_22807;
wire v_22808;
wire v_22809;
wire v_22810;
wire v_22811;
wire v_22812;
wire v_22813;
wire v_22814;
wire v_22815;
wire v_22816;
wire v_22817;
wire v_22818;
wire v_22819;
wire v_22820;
wire v_22821;
wire v_22822;
wire v_22823;
wire v_22824;
wire v_22825;
wire v_22826;
wire v_22827;
wire v_22828;
wire v_22829;
wire v_22830;
wire v_22831;
wire v_22832;
wire v_22833;
wire v_22834;
wire v_22835;
wire v_22836;
wire v_22837;
wire v_22838;
wire v_22839;
wire v_22840;
wire v_22841;
wire v_22842;
wire v_22843;
wire v_22844;
wire v_22845;
wire v_22846;
wire v_22847;
wire v_22848;
wire v_22849;
wire v_22850;
wire v_22851;
wire v_22852;
wire v_22853;
wire v_22854;
wire v_22855;
wire v_22856;
wire v_22857;
wire v_22858;
wire v_22859;
wire v_22860;
wire v_22861;
wire v_22862;
wire v_22863;
wire v_22864;
wire v_22865;
wire v_22866;
wire v_22867;
wire v_22868;
wire v_22869;
wire v_22870;
wire v_22871;
wire v_22872;
wire v_22873;
wire v_22874;
wire v_22875;
wire v_22876;
wire v_22877;
wire v_22878;
wire v_22879;
wire v_22880;
wire v_22881;
wire v_22882;
wire v_22883;
wire v_22884;
wire v_22885;
wire v_22886;
wire v_22887;
wire v_22888;
wire v_22889;
wire v_22890;
wire v_22891;
wire v_22892;
wire v_22893;
wire v_22894;
wire v_22895;
wire v_22896;
wire v_22897;
wire v_22898;
wire v_22899;
wire v_22900;
wire v_22901;
wire v_22902;
wire v_22903;
wire v_22904;
wire v_22905;
wire v_22906;
wire v_22907;
wire v_22908;
wire v_22909;
wire v_22910;
wire v_22911;
wire v_22912;
wire v_22913;
wire v_22914;
wire v_22915;
wire v_22916;
wire v_22917;
wire v_22918;
wire v_22919;
wire v_22920;
wire v_22921;
wire v_22922;
wire v_22923;
wire v_22924;
wire v_22925;
wire v_22926;
wire v_22927;
wire v_22928;
wire v_22929;
wire v_22930;
wire v_22931;
wire v_22932;
wire v_22933;
wire v_22934;
wire v_22935;
wire v_22936;
wire v_22937;
wire v_22938;
wire v_22939;
wire v_22940;
wire v_22941;
wire v_22942;
wire v_22943;
wire v_22944;
wire v_22945;
wire v_22946;
wire v_22947;
wire v_22948;
wire v_22949;
wire v_22950;
wire v_22951;
wire v_22952;
wire v_22953;
wire v_22954;
wire v_22955;
wire v_22956;
wire v_22957;
wire v_22958;
wire v_22959;
wire v_22960;
wire v_22961;
wire v_22962;
wire v_22963;
wire v_22964;
wire v_22965;
wire v_22966;
wire v_22967;
wire v_22968;
wire v_22969;
wire v_22970;
wire v_22971;
wire v_22972;
wire v_22973;
wire v_22974;
wire v_22975;
wire v_22976;
wire v_22977;
wire v_22978;
wire v_22979;
wire v_22980;
wire v_22981;
wire v_22982;
wire v_22983;
wire v_22984;
wire v_22985;
wire v_22986;
wire v_22987;
wire v_22988;
wire v_22989;
wire v_22990;
wire v_22991;
wire v_22992;
wire v_22993;
wire v_22994;
wire v_22996;
wire v_22997;
wire v_22998;
wire v_22999;
wire v_23000;
wire v_23001;
wire v_23002;
wire v_23003;
wire v_23004;
wire v_23005;
wire v_23006;
wire v_23007;
wire v_23008;
wire v_23009;
wire v_23010;
wire v_23011;
wire v_23012;
wire v_23013;
wire v_23014;
wire v_23015;
wire v_23016;
wire v_23017;
wire v_23018;
wire v_23019;
wire v_23020;
wire v_23021;
wire v_23022;
wire v_23023;
wire v_23024;
wire v_23025;
wire v_23026;
wire v_23027;
wire v_23028;
wire v_23029;
wire v_23030;
wire v_23031;
wire v_23032;
wire v_23033;
wire v_23034;
wire v_23035;
wire v_23036;
wire v_23037;
wire v_23038;
wire v_23039;
wire v_23040;
wire v_23041;
wire v_23042;
wire v_23043;
wire v_23044;
wire v_23045;
wire v_23046;
wire v_23047;
wire v_23048;
wire v_23049;
wire v_23050;
wire v_23051;
wire v_23052;
wire v_23053;
wire v_23054;
wire v_23055;
wire v_23056;
wire v_23057;
wire v_23058;
wire v_23059;
wire v_23060;
wire v_23061;
wire v_23062;
wire v_23063;
wire v_23064;
wire v_23065;
wire v_23066;
wire v_23067;
wire v_23068;
wire v_23069;
wire v_23070;
wire v_23071;
wire v_23072;
wire v_23073;
wire v_23074;
wire v_23075;
wire v_23076;
wire v_23077;
wire v_23078;
wire v_23079;
wire v_23080;
wire v_23081;
wire v_23082;
wire v_23083;
wire v_23084;
wire v_23085;
wire v_23086;
wire v_23087;
wire v_23088;
wire v_23089;
wire v_23090;
wire v_23091;
wire v_23092;
wire v_23093;
wire v_23094;
wire v_23095;
wire v_23096;
wire v_23097;
wire v_23098;
wire v_23099;
wire v_23100;
wire v_23101;
wire v_23102;
wire v_23103;
wire v_23104;
wire v_23105;
wire v_23106;
wire v_23107;
wire v_23108;
wire v_23109;
wire v_23110;
wire v_23111;
wire v_23112;
wire v_23113;
wire v_23114;
wire v_23115;
wire v_23116;
wire v_23117;
wire v_23118;
wire v_23119;
wire v_23120;
wire v_23121;
wire v_23122;
wire v_23123;
wire v_23124;
wire v_23125;
wire v_23126;
wire v_23127;
wire v_23128;
wire v_23129;
wire v_23130;
wire v_23131;
wire v_23132;
wire v_23133;
wire v_23134;
wire v_23135;
wire v_23136;
wire v_23137;
wire v_23138;
wire v_23139;
wire v_23140;
wire v_23141;
wire v_23142;
wire v_23143;
wire v_23144;
wire v_23145;
wire v_23146;
wire v_23147;
wire v_23148;
wire v_23149;
wire v_23150;
wire v_23151;
wire v_23152;
wire v_23153;
wire v_23154;
wire v_23155;
wire v_23156;
wire v_23157;
wire v_23158;
wire v_23159;
wire v_23160;
wire v_23161;
wire v_23162;
wire v_23163;
wire v_23164;
wire v_23165;
wire v_23166;
wire v_23167;
wire v_23168;
wire v_23169;
wire v_23170;
wire v_23171;
wire v_23172;
wire v_23173;
wire v_23174;
wire v_23175;
wire v_23176;
wire v_23177;
wire v_23178;
wire v_23179;
wire v_23180;
wire v_23181;
wire v_23182;
wire v_23183;
wire v_23184;
wire v_23185;
wire v_23186;
wire v_23187;
wire v_23188;
wire v_23189;
wire v_23190;
wire v_23191;
wire v_23192;
wire v_23193;
wire v_23194;
wire v_23195;
wire v_23196;
wire v_23197;
wire v_23198;
wire v_23199;
wire v_23200;
wire v_23201;
wire v_23202;
wire v_23203;
wire v_23204;
wire v_23205;
wire v_23206;
wire v_23207;
wire v_23208;
wire v_23209;
wire v_23210;
wire v_23211;
wire v_23212;
wire v_23213;
wire v_23214;
wire v_23215;
wire v_23216;
wire v_23217;
wire v_23218;
wire v_23219;
wire v_23220;
wire v_23221;
wire v_23222;
wire v_23223;
wire v_23224;
wire v_23225;
wire v_23226;
wire v_23227;
wire v_23228;
wire v_23229;
wire v_23230;
wire v_23231;
wire v_23232;
wire v_23233;
wire v_23234;
wire v_23235;
wire v_23236;
wire v_23237;
wire v_23239;
wire v_23240;
wire v_23241;
wire v_23242;
wire v_23243;
wire v_23244;
wire v_23245;
wire v_23246;
wire v_23247;
wire v_23248;
wire v_23249;
wire v_23250;
wire v_23251;
wire v_23252;
wire v_23253;
wire v_23254;
wire v_23255;
wire v_23256;
wire v_23257;
wire v_23258;
wire v_23259;
wire v_23260;
wire v_23261;
wire v_23262;
wire v_23263;
wire v_23264;
wire v_23265;
wire v_23266;
wire v_23267;
wire v_23268;
wire v_23269;
wire v_23270;
wire v_23271;
wire v_23272;
wire v_23273;
wire v_23274;
wire v_23275;
wire v_23276;
wire v_23277;
wire v_23278;
wire v_23279;
wire v_23280;
wire v_23281;
wire v_23282;
wire v_23283;
wire v_23284;
wire v_23285;
wire v_23286;
wire v_23287;
wire v_23288;
wire v_23289;
wire v_23290;
wire v_23291;
wire v_23292;
wire v_23293;
wire v_23294;
wire v_23295;
wire v_23296;
wire v_23297;
wire v_23298;
wire v_23299;
wire v_23300;
wire v_23301;
wire v_23302;
wire v_23303;
wire v_23304;
wire v_23305;
wire v_23306;
wire v_23307;
wire v_23308;
wire v_23309;
wire v_23310;
wire v_23311;
wire v_23312;
wire v_23313;
wire v_23314;
wire v_23315;
wire v_23316;
wire v_23317;
wire v_23318;
wire v_23319;
wire v_23320;
wire v_23321;
wire v_23322;
wire v_23323;
wire v_23324;
wire v_23325;
wire v_23326;
wire v_23327;
wire v_23328;
wire v_23329;
wire v_23330;
wire v_23331;
wire v_23332;
wire v_23333;
wire v_23334;
wire v_23335;
wire v_23336;
wire v_23337;
wire v_23338;
wire v_23339;
wire v_23340;
wire v_23341;
wire v_23342;
wire v_23343;
wire v_23344;
wire v_23345;
wire v_23346;
wire v_23347;
wire v_23348;
wire v_23349;
wire v_23350;
wire v_23351;
wire v_23352;
wire v_23353;
wire v_23354;
wire v_23355;
wire v_23356;
wire v_23357;
wire v_23358;
wire v_23359;
wire v_23360;
wire v_23361;
wire v_23362;
wire v_23363;
wire v_23364;
wire v_23365;
wire v_23366;
wire v_23367;
wire v_23368;
wire v_23369;
wire v_23370;
wire v_23371;
wire v_23372;
wire v_23373;
wire v_23374;
wire v_23375;
wire v_23376;
wire v_23377;
wire v_23378;
wire v_23379;
wire v_23380;
wire v_23381;
wire v_23382;
wire v_23383;
wire v_23384;
wire v_23385;
wire v_23386;
wire v_23387;
wire v_23388;
wire v_23389;
wire v_23390;
wire v_23391;
wire v_23392;
wire v_23393;
wire v_23394;
wire v_23395;
wire v_23396;
wire v_23397;
wire v_23398;
wire v_23399;
wire v_23400;
wire v_23401;
wire v_23402;
wire v_23403;
wire v_23404;
wire v_23405;
wire v_23406;
wire v_23407;
wire v_23408;
wire v_23409;
wire v_23410;
wire v_23411;
wire v_23412;
wire v_23413;
wire v_23414;
wire v_23415;
wire v_23416;
wire v_23417;
wire v_23418;
wire v_23419;
wire v_23420;
wire v_23421;
wire v_23422;
wire v_23423;
wire v_23424;
wire v_23425;
wire v_23426;
wire v_23427;
wire v_23428;
wire v_23429;
wire v_23430;
wire v_23431;
wire v_23432;
wire v_23433;
wire v_23434;
wire v_23435;
wire v_23436;
wire v_23437;
wire v_23438;
wire v_23439;
wire v_23440;
wire v_23441;
wire v_23442;
wire v_23443;
wire v_23444;
wire v_23445;
wire v_23446;
wire v_23447;
wire v_23448;
wire v_23449;
wire v_23450;
wire v_23451;
wire v_23452;
wire v_23453;
wire v_23454;
wire v_23455;
wire v_23456;
wire v_23457;
wire v_23458;
wire v_23459;
wire v_23460;
wire v_23461;
wire v_23462;
wire v_23463;
wire v_23464;
wire v_23465;
wire v_23466;
wire v_23467;
wire v_23468;
wire v_23469;
wire v_23470;
wire v_23471;
wire v_23472;
wire v_23473;
wire v_23474;
wire v_23475;
wire v_23476;
wire v_23477;
wire v_23478;
wire v_23479;
wire v_23480;
wire v_23482;
wire v_23483;
wire v_23484;
wire v_23485;
wire v_23486;
wire v_23487;
wire v_23488;
wire v_23489;
wire v_23490;
wire v_23491;
wire v_23492;
wire v_23493;
wire v_23494;
wire v_23495;
wire v_23496;
wire v_23497;
wire v_23498;
wire v_23499;
wire v_23500;
wire v_23501;
wire v_23502;
wire v_23503;
wire v_23504;
wire v_23505;
wire v_23506;
wire v_23507;
wire v_23508;
wire v_23509;
wire v_23510;
wire v_23511;
wire v_23512;
wire v_23513;
wire v_23514;
wire v_23515;
wire v_23516;
wire v_23517;
wire v_23518;
wire v_23519;
wire v_23520;
wire v_23521;
wire v_23522;
wire v_23523;
wire v_23524;
wire v_23525;
wire v_23526;
wire v_23527;
wire v_23528;
wire v_23529;
wire v_23530;
wire v_23531;
wire v_23532;
wire v_23533;
wire v_23534;
wire v_23535;
wire v_23536;
wire v_23537;
wire v_23538;
wire v_23539;
wire v_23540;
wire v_23541;
wire v_23542;
wire v_23543;
wire v_23544;
wire v_23545;
wire v_23546;
wire v_23547;
wire v_23548;
wire v_23549;
wire v_23550;
wire v_23551;
wire v_23552;
wire v_23553;
wire v_23554;
wire v_23555;
wire v_23556;
wire v_23557;
wire v_23558;
wire v_23559;
wire v_23560;
wire v_23561;
wire v_23562;
wire v_23563;
wire v_23564;
wire v_23565;
wire v_23566;
wire v_23567;
wire v_23568;
wire v_23569;
wire v_23570;
wire v_23571;
wire v_23572;
wire v_23573;
wire v_23574;
wire v_23575;
wire v_23576;
wire v_23577;
wire v_23578;
wire v_23579;
wire v_23580;
wire v_23581;
wire v_23582;
wire v_23583;
wire v_23584;
wire v_23585;
wire v_23586;
wire v_23587;
wire v_23588;
wire v_23589;
wire v_23590;
wire v_23591;
wire v_23592;
wire v_23593;
wire v_23594;
wire v_23595;
wire v_23596;
wire v_23597;
wire v_23598;
wire v_23599;
wire v_23600;
wire v_23601;
wire v_23602;
wire v_23603;
wire v_23604;
wire v_23605;
wire v_23606;
wire v_23607;
wire v_23608;
wire v_23609;
wire v_23610;
wire v_23611;
wire v_23612;
wire v_23613;
wire v_23614;
wire v_23615;
wire v_23616;
wire v_23617;
wire v_23618;
wire v_23619;
wire v_23620;
wire v_23621;
wire v_23622;
wire v_23623;
wire v_23624;
wire v_23625;
wire v_23626;
wire v_23627;
wire v_23628;
wire v_23629;
wire v_23630;
wire v_23631;
wire v_23632;
wire v_23633;
wire v_23634;
wire v_23635;
wire v_23636;
wire v_23637;
wire v_23638;
wire v_23639;
wire v_23640;
wire v_23641;
wire v_23642;
wire v_23643;
wire v_23644;
wire v_23645;
wire v_23646;
wire v_23647;
wire v_23648;
wire v_23649;
wire v_23650;
wire v_23651;
wire v_23652;
wire v_23653;
wire v_23654;
wire v_23655;
wire v_23656;
wire v_23657;
wire v_23658;
wire v_23659;
wire v_23660;
wire v_23661;
wire v_23662;
wire v_23663;
wire v_23664;
wire v_23665;
wire v_23666;
wire v_23667;
wire v_23668;
wire v_23669;
wire v_23670;
wire v_23671;
wire v_23672;
wire v_23673;
wire v_23674;
wire v_23675;
wire v_23676;
wire v_23677;
wire v_23678;
wire v_23679;
wire v_23680;
wire v_23681;
wire v_23682;
wire v_23683;
wire v_23684;
wire v_23685;
wire v_23686;
wire v_23687;
wire v_23688;
wire v_23689;
wire v_23690;
wire v_23691;
wire v_23692;
wire v_23693;
wire v_23694;
wire v_23695;
wire v_23696;
wire v_23697;
wire v_23698;
wire v_23699;
wire v_23700;
wire v_23701;
wire v_23702;
wire v_23703;
wire v_23704;
wire v_23705;
wire v_23706;
wire v_23707;
wire v_23708;
wire v_23709;
wire v_23710;
wire v_23711;
wire v_23712;
wire v_23713;
wire v_23714;
wire v_23715;
wire v_23716;
wire v_23717;
wire v_23718;
wire v_23719;
wire v_23720;
wire v_23721;
wire v_23722;
wire v_23723;
wire v_23725;
wire v_23726;
wire v_23727;
wire v_23728;
wire v_23729;
wire v_23730;
wire v_23731;
wire v_23732;
wire v_23733;
wire v_23734;
wire v_23735;
wire v_23736;
wire v_23737;
wire v_23738;
wire v_23739;
wire v_23740;
wire v_23741;
wire v_23742;
wire v_23743;
wire v_23744;
wire v_23745;
wire v_23746;
wire v_23747;
wire v_23748;
wire v_23749;
wire v_23750;
wire v_23751;
wire v_23752;
wire v_23753;
wire v_23754;
wire v_23755;
wire v_23756;
wire v_23757;
wire v_23758;
wire v_23759;
wire v_23760;
wire v_23761;
wire v_23762;
wire v_23763;
wire v_23764;
wire v_23765;
wire v_23766;
wire v_23767;
wire v_23768;
wire v_23769;
wire v_23770;
wire v_23771;
wire v_23772;
wire v_23773;
wire v_23774;
wire v_23775;
wire v_23776;
wire v_23777;
wire v_23778;
wire v_23779;
wire v_23780;
wire v_23781;
wire v_23782;
wire v_23783;
wire v_23784;
wire v_23785;
wire v_23786;
wire v_23787;
wire v_23788;
wire v_23789;
wire v_23790;
wire v_23791;
wire v_23792;
wire v_23793;
wire v_23794;
wire v_23795;
wire v_23796;
wire v_23797;
wire v_23798;
wire v_23799;
wire v_23800;
wire v_23801;
wire v_23802;
wire v_23803;
wire v_23804;
wire v_23805;
wire v_23806;
wire v_23807;
wire v_23808;
wire v_23809;
wire v_23810;
wire v_23811;
wire v_23812;
wire v_23813;
wire v_23814;
wire v_23815;
wire v_23816;
wire v_23817;
wire v_23818;
wire v_23819;
wire v_23820;
wire v_23821;
wire v_23822;
wire v_23823;
wire v_23824;
wire v_23825;
wire v_23826;
wire v_23827;
wire v_23828;
wire v_23829;
wire v_23830;
wire v_23831;
wire v_23832;
wire v_23833;
wire v_23834;
wire v_23835;
wire v_23836;
wire v_23837;
wire v_23838;
wire v_23839;
wire v_23840;
wire v_23841;
wire v_23842;
wire v_23843;
wire v_23844;
wire v_23845;
wire v_23846;
wire v_23847;
wire v_23848;
wire v_23849;
wire v_23850;
wire v_23851;
wire v_23852;
wire v_23853;
wire v_23854;
wire v_23855;
wire v_23856;
wire v_23857;
wire v_23858;
wire v_23859;
wire v_23860;
wire v_23861;
wire v_23862;
wire v_23863;
wire v_23864;
wire v_23865;
wire v_23866;
wire v_23867;
wire v_23868;
wire v_23869;
wire v_23870;
wire v_23871;
wire v_23872;
wire v_23873;
wire v_23874;
wire v_23875;
wire v_23876;
wire v_23877;
wire v_23878;
wire v_23879;
wire v_23880;
wire v_23881;
wire v_23882;
wire v_23883;
wire v_23884;
wire v_23885;
wire v_23886;
wire v_23887;
wire v_23888;
wire v_23889;
wire v_23890;
wire v_23891;
wire v_23892;
wire v_23893;
wire v_23894;
wire v_23895;
wire v_23896;
wire v_23897;
wire v_23898;
wire v_23899;
wire v_23900;
wire v_23901;
wire v_23902;
wire v_23903;
wire v_23904;
wire v_23905;
wire v_23906;
wire v_23907;
wire v_23908;
wire v_23909;
wire v_23910;
wire v_23911;
wire v_23912;
wire v_23913;
wire v_23914;
wire v_23915;
wire v_23916;
wire v_23917;
wire v_23918;
wire v_23919;
wire v_23920;
wire v_23921;
wire v_23922;
wire v_23923;
wire v_23924;
wire v_23925;
wire v_23926;
wire v_23927;
wire v_23928;
wire v_23929;
wire v_23930;
wire v_23931;
wire v_23932;
wire v_23933;
wire v_23934;
wire v_23935;
wire v_23936;
wire v_23937;
wire v_23938;
wire v_23939;
wire v_23940;
wire v_23941;
wire v_23942;
wire v_23943;
wire v_23944;
wire v_23945;
wire v_23946;
wire v_23947;
wire v_23948;
wire v_23949;
wire v_23950;
wire v_23951;
wire v_23952;
wire v_23953;
wire v_23954;
wire v_23955;
wire v_23956;
wire v_23957;
wire v_23958;
wire v_23959;
wire v_23960;
wire v_23961;
wire v_23962;
wire v_23963;
wire v_23964;
wire v_23965;
wire v_23966;
wire v_23968;
wire v_23969;
wire v_23970;
wire v_23971;
wire v_23972;
wire v_23973;
wire v_23974;
wire v_23975;
wire v_23976;
wire v_23977;
wire v_23978;
wire v_23979;
wire v_23980;
wire v_23981;
wire v_23982;
wire v_23983;
wire v_23984;
wire v_23985;
wire v_23986;
wire v_23987;
wire v_23988;
wire v_23989;
wire v_23990;
wire v_23991;
wire v_23992;
wire v_23993;
wire v_23994;
wire v_23995;
wire v_23996;
wire v_23997;
wire v_23998;
wire v_23999;
wire v_24000;
wire v_24001;
wire v_24002;
wire v_24003;
wire v_24004;
wire v_24005;
wire v_24006;
wire v_24007;
wire v_24008;
wire v_24009;
wire v_24010;
wire v_24011;
wire v_24012;
wire v_24013;
wire v_24014;
wire v_24015;
wire v_24016;
wire v_24017;
wire v_24018;
wire v_24019;
wire v_24020;
wire v_24021;
wire v_24022;
wire v_24023;
wire v_24024;
wire v_24025;
wire v_24026;
wire v_24027;
wire v_24028;
wire v_24029;
wire v_24030;
wire v_24031;
wire v_24032;
wire v_24033;
wire v_24034;
wire v_24035;
wire v_24036;
wire v_24037;
wire v_24038;
wire v_24039;
wire v_24040;
wire v_24041;
wire v_24042;
wire v_24043;
wire v_24044;
wire v_24045;
wire v_24046;
wire v_24047;
wire v_24048;
wire v_24049;
wire v_24050;
wire v_24051;
wire v_24052;
wire v_24053;
wire v_24054;
wire v_24055;
wire v_24056;
wire v_24057;
wire v_24058;
wire v_24059;
wire v_24060;
wire v_24061;
wire v_24062;
wire v_24063;
wire v_24064;
wire v_24065;
wire v_24066;
wire v_24067;
wire v_24068;
wire v_24069;
wire v_24070;
wire v_24071;
wire v_24072;
wire v_24073;
wire v_24074;
wire v_24075;
wire v_24076;
wire v_24077;
wire v_24078;
wire v_24079;
wire v_24080;
wire v_24081;
wire v_24082;
wire v_24083;
wire v_24084;
wire v_24085;
wire v_24086;
wire v_24087;
wire v_24088;
wire v_24089;
wire v_24090;
wire v_24091;
wire v_24092;
wire v_24093;
wire v_24094;
wire v_24095;
wire v_24096;
wire v_24097;
wire v_24098;
wire v_24099;
wire v_24100;
wire v_24101;
wire v_24102;
wire v_24103;
wire v_24104;
wire v_24105;
wire v_24106;
wire v_24107;
wire v_24108;
wire v_24109;
wire v_24110;
wire v_24111;
wire v_24112;
wire v_24113;
wire v_24114;
wire v_24115;
wire v_24116;
wire v_24117;
wire v_24118;
wire v_24119;
wire v_24120;
wire v_24121;
wire v_24122;
wire v_24123;
wire v_24124;
wire v_24125;
wire v_24126;
wire v_24127;
wire v_24128;
wire v_24129;
wire v_24130;
wire v_24131;
wire v_24132;
wire v_24133;
wire v_24134;
wire v_24135;
wire v_24136;
wire v_24137;
wire v_24138;
wire v_24139;
wire v_24140;
wire v_24141;
wire v_24142;
wire v_24143;
wire v_24144;
wire v_24145;
wire v_24146;
wire v_24147;
wire v_24148;
wire v_24149;
wire v_24150;
wire v_24151;
wire v_24152;
wire v_24153;
wire v_24154;
wire v_24155;
wire v_24156;
wire v_24157;
wire v_24158;
wire v_24159;
wire v_24160;
wire v_24161;
wire v_24162;
wire v_24163;
wire v_24164;
wire v_24165;
wire v_24166;
wire v_24167;
wire v_24168;
wire v_24169;
wire v_24170;
wire v_24171;
wire v_24172;
wire v_24173;
wire v_24174;
wire v_24175;
wire v_24176;
wire v_24177;
wire v_24178;
wire v_24179;
wire v_24180;
wire v_24181;
wire v_24182;
wire v_24183;
wire v_24184;
wire v_24185;
wire v_24186;
wire v_24187;
wire v_24188;
wire v_24189;
wire v_24190;
wire v_24191;
wire v_24192;
wire v_24193;
wire v_24194;
wire v_24195;
wire v_24196;
wire v_24197;
wire v_24198;
wire v_24199;
wire v_24200;
wire v_24201;
wire v_24202;
wire v_24203;
wire v_24204;
wire v_24205;
wire v_24206;
wire v_24207;
wire v_24208;
wire v_24209;
wire v_24211;
wire v_24212;
wire v_24213;
wire v_24214;
wire v_24215;
wire v_24216;
wire v_24217;
wire v_24218;
wire v_24219;
wire v_24220;
wire v_24221;
wire v_24222;
wire v_24223;
wire v_24224;
wire v_24225;
wire v_24226;
wire v_24227;
wire v_24228;
wire v_24229;
wire v_24230;
wire v_24231;
wire v_24232;
wire v_24233;
wire v_24234;
wire v_24235;
wire v_24236;
wire v_24237;
wire v_24238;
wire v_24239;
wire v_24240;
wire v_24241;
wire v_24242;
wire v_24243;
wire v_24244;
wire v_24245;
wire v_24246;
wire v_24247;
wire v_24248;
wire v_24249;
wire v_24250;
wire v_24251;
wire v_24252;
wire v_24253;
wire v_24254;
wire v_24255;
wire v_24256;
wire v_24257;
wire v_24258;
wire v_24259;
wire v_24260;
wire v_24261;
wire v_24262;
wire v_24263;
wire v_24264;
wire v_24265;
wire v_24266;
wire v_24267;
wire v_24268;
wire v_24269;
wire v_24270;
wire v_24271;
wire v_24272;
wire v_24273;
wire v_24274;
wire v_24275;
wire v_24276;
wire v_24277;
wire v_24278;
wire v_24279;
wire v_24280;
wire v_24281;
wire v_24282;
wire v_24283;
wire v_24284;
wire v_24285;
wire v_24286;
wire v_24287;
wire v_24288;
wire v_24289;
wire v_24290;
wire v_24291;
wire v_24292;
wire v_24293;
wire v_24294;
wire v_24295;
wire v_24296;
wire v_24297;
wire v_24298;
wire v_24299;
wire v_24300;
wire v_24301;
wire v_24302;
wire v_24303;
wire v_24304;
wire v_24305;
wire v_24306;
wire v_24307;
wire v_24308;
wire v_24309;
wire v_24310;
wire v_24311;
wire v_24312;
wire v_24313;
wire v_24314;
wire v_24315;
wire v_24316;
wire v_24317;
wire v_24318;
wire v_24319;
wire v_24320;
wire v_24321;
wire v_24322;
wire v_24323;
wire v_24324;
wire v_24325;
wire v_24326;
wire v_24327;
wire v_24328;
wire v_24329;
wire v_24330;
wire v_24331;
wire v_24332;
wire v_24333;
wire v_24334;
wire v_24335;
wire v_24336;
wire v_24337;
wire v_24338;
wire v_24339;
wire v_24340;
wire v_24341;
wire v_24342;
wire v_24343;
wire v_24344;
wire v_24345;
wire v_24346;
wire v_24347;
wire v_24348;
wire v_24349;
wire v_24350;
wire v_24351;
wire v_24352;
wire v_24353;
wire v_24354;
wire v_24355;
wire v_24356;
wire v_24357;
wire v_24358;
wire v_24359;
wire v_24360;
wire v_24361;
wire v_24362;
wire v_24363;
wire v_24364;
wire v_24365;
wire v_24366;
wire v_24367;
wire v_24368;
wire v_24369;
wire v_24370;
wire v_24371;
wire v_24372;
wire v_24373;
wire v_24374;
wire v_24375;
wire v_24376;
wire v_24377;
wire v_24378;
wire v_24379;
wire v_24380;
wire v_24381;
wire v_24382;
wire v_24383;
wire v_24384;
wire v_24385;
wire v_24386;
wire v_24387;
wire v_24388;
wire v_24389;
wire v_24390;
wire v_24391;
wire v_24392;
wire v_24393;
wire v_24394;
wire v_24395;
wire v_24396;
wire v_24397;
wire v_24398;
wire v_24399;
wire v_24400;
wire v_24401;
wire v_24402;
wire v_24403;
wire v_24404;
wire v_24405;
wire v_24406;
wire v_24407;
wire v_24408;
wire v_24409;
wire v_24410;
wire v_24411;
wire v_24412;
wire v_24413;
wire v_24414;
wire v_24415;
wire v_24416;
wire v_24417;
wire v_24418;
wire v_24419;
wire v_24420;
wire v_24421;
wire v_24422;
wire v_24423;
wire v_24424;
wire v_24425;
wire v_24426;
wire v_24427;
wire v_24428;
wire v_24429;
wire v_24430;
wire v_24431;
wire v_24432;
wire v_24433;
wire v_24434;
wire v_24435;
wire v_24436;
wire v_24437;
wire v_24438;
wire v_24439;
wire v_24440;
wire v_24441;
wire v_24442;
wire v_24443;
wire v_24444;
wire v_24445;
wire v_24446;
wire v_24447;
wire v_24448;
wire v_24449;
wire v_24450;
wire v_24451;
wire v_24452;
wire v_24454;
wire v_24455;
wire v_24456;
wire v_24457;
wire v_24458;
wire v_24459;
wire v_24460;
wire v_24461;
wire v_24462;
wire v_24463;
wire v_24464;
wire v_24465;
wire v_24466;
wire v_24467;
wire v_24468;
wire v_24469;
wire v_24470;
wire v_24471;
wire v_24472;
wire v_24473;
wire v_24474;
wire v_24475;
wire v_24476;
wire v_24477;
wire v_24478;
wire v_24479;
wire v_24480;
wire v_24481;
wire v_24482;
wire v_24483;
wire v_24484;
wire v_24485;
wire v_24486;
wire v_24487;
wire v_24488;
wire v_24489;
wire v_24490;
wire v_24491;
wire v_24492;
wire v_24493;
wire v_24494;
wire v_24495;
wire v_24496;
wire v_24497;
wire v_24498;
wire v_24499;
wire v_24500;
wire v_24501;
wire v_24502;
wire v_24503;
wire v_24504;
wire v_24505;
wire v_24506;
wire v_24507;
wire v_24508;
wire v_24509;
wire v_24510;
wire v_24511;
wire v_24512;
wire v_24513;
wire v_24514;
wire v_24515;
wire v_24516;
wire v_24517;
wire v_24518;
wire v_24519;
wire v_24520;
wire v_24521;
wire v_24522;
wire v_24523;
wire v_24524;
wire v_24525;
wire v_24526;
wire v_24527;
wire v_24528;
wire v_24529;
wire v_24530;
wire v_24531;
wire v_24532;
wire v_24533;
wire v_24534;
wire v_24535;
wire v_24536;
wire v_24537;
wire v_24538;
wire v_24539;
wire v_24540;
wire v_24541;
wire v_24542;
wire v_24543;
wire v_24544;
wire v_24545;
wire v_24546;
wire v_24547;
wire v_24548;
wire v_24549;
wire v_24550;
wire v_24551;
wire v_24552;
wire v_24553;
wire v_24554;
wire v_24555;
wire v_24556;
wire v_24557;
wire v_24558;
wire v_24559;
wire v_24560;
wire v_24561;
wire v_24562;
wire v_24563;
wire v_24564;
wire v_24565;
wire v_24566;
wire v_24567;
wire v_24568;
wire v_24569;
wire v_24570;
wire v_24571;
wire v_24572;
wire v_24573;
wire v_24574;
wire v_24575;
wire v_24576;
wire v_24577;
wire v_24578;
wire v_24579;
wire v_24580;
wire v_24581;
wire v_24582;
wire v_24583;
wire v_24584;
wire v_24585;
wire v_24586;
wire v_24587;
wire v_24588;
wire v_24589;
wire v_24590;
wire v_24591;
wire v_24592;
wire v_24593;
wire v_24594;
wire v_24595;
wire v_24596;
wire v_24597;
wire v_24598;
wire v_24599;
wire v_24600;
wire v_24601;
wire v_24602;
wire v_24603;
wire v_24604;
wire v_24605;
wire v_24606;
wire v_24607;
wire v_24608;
wire v_24609;
wire v_24610;
wire v_24611;
wire v_24612;
wire v_24613;
wire v_24614;
wire v_24615;
wire v_24616;
wire v_24617;
wire v_24618;
wire v_24619;
wire v_24620;
wire v_24621;
wire v_24622;
wire v_24623;
wire v_24624;
wire v_24625;
wire v_24626;
wire v_24627;
wire v_24628;
wire v_24629;
wire v_24630;
wire v_24631;
wire v_24632;
wire v_24633;
wire v_24634;
wire v_24635;
wire v_24636;
wire v_24637;
wire v_24638;
wire v_24639;
wire v_24640;
wire v_24641;
wire v_24642;
wire v_24643;
wire v_24644;
wire v_24645;
wire v_24646;
wire v_24647;
wire v_24648;
wire v_24649;
wire v_24650;
wire v_24651;
wire v_24652;
wire v_24653;
wire v_24654;
wire v_24655;
wire v_24656;
wire v_24657;
wire v_24658;
wire v_24659;
wire v_24660;
wire v_24661;
wire v_24662;
wire v_24663;
wire v_24664;
wire v_24665;
wire v_24666;
wire v_24667;
wire v_24668;
wire v_24669;
wire v_24670;
wire v_24671;
wire v_24672;
wire v_24673;
wire v_24674;
wire v_24675;
wire v_24676;
wire v_24677;
wire v_24678;
wire v_24679;
wire v_24680;
wire v_24681;
wire v_24682;
wire v_24683;
wire v_24684;
wire v_24685;
wire v_24686;
wire v_24687;
wire v_24688;
wire v_24689;
wire v_24690;
wire v_24691;
wire v_24692;
wire v_24693;
wire v_24694;
wire v_24695;
wire v_24697;
wire v_24698;
wire v_24699;
wire v_24700;
wire v_24701;
wire v_24702;
wire v_24703;
wire v_24704;
wire v_24705;
wire v_24706;
wire v_24707;
wire v_24708;
wire v_24709;
wire v_24710;
wire v_24711;
wire v_24712;
wire v_24713;
wire v_24714;
wire v_24715;
wire v_24716;
wire v_24717;
wire v_24718;
wire v_24719;
wire v_24720;
wire v_24721;
wire v_24722;
wire v_24723;
wire v_24724;
wire v_24725;
wire v_24726;
wire v_24727;
wire v_24728;
wire v_24729;
wire v_24730;
wire v_24731;
wire v_24732;
wire v_24733;
wire v_24734;
wire v_24735;
wire v_24736;
wire v_24737;
wire v_24738;
wire v_24739;
wire v_24740;
wire v_24741;
wire v_24742;
wire v_24743;
wire v_24744;
wire v_24745;
wire v_24746;
wire v_24747;
wire v_24748;
wire v_24749;
wire v_24750;
wire v_24751;
wire v_24752;
wire v_24753;
wire v_24754;
wire v_24755;
wire v_24756;
wire v_24757;
wire v_24758;
wire v_24759;
wire v_24760;
wire v_24761;
wire v_24762;
wire v_24763;
wire v_24764;
wire v_24765;
wire v_24766;
wire v_24767;
wire v_24768;
wire v_24769;
wire v_24770;
wire v_24771;
wire v_24772;
wire v_24773;
wire v_24774;
wire v_24775;
wire v_24776;
wire v_24777;
wire v_24778;
wire v_24779;
wire v_24780;
wire v_24781;
wire v_24782;
wire v_24783;
wire v_24784;
wire v_24785;
wire v_24786;
wire v_24787;
wire v_24788;
wire v_24789;
wire v_24790;
wire v_24791;
wire v_24792;
wire v_24793;
wire v_24794;
wire v_24795;
wire v_24796;
wire v_24797;
wire v_24798;
wire v_24799;
wire v_24800;
wire v_24801;
wire v_24802;
wire v_24803;
wire v_24804;
wire v_24805;
wire v_24806;
wire v_24807;
wire v_24808;
wire v_24809;
wire v_24810;
wire v_24811;
wire v_24812;
wire v_24813;
wire v_24814;
wire v_24815;
wire v_24816;
wire v_24817;
wire v_24818;
wire v_24819;
wire v_24820;
wire v_24821;
wire v_24822;
wire v_24823;
wire v_24824;
wire v_24825;
wire v_24826;
wire v_24827;
wire v_24828;
wire v_24829;
wire v_24830;
wire v_24831;
wire v_24832;
wire v_24833;
wire v_24834;
wire v_24835;
wire v_24836;
wire v_24837;
wire v_24838;
wire v_24839;
wire v_24840;
wire v_24841;
wire v_24842;
wire v_24843;
wire v_24844;
wire v_24845;
wire v_24846;
wire v_24847;
wire v_24848;
wire v_24849;
wire v_24850;
wire v_24851;
wire v_24852;
wire v_24853;
wire v_24854;
wire v_24855;
wire v_24856;
wire v_24857;
wire v_24858;
wire v_24859;
wire v_24860;
wire v_24861;
wire v_24862;
wire v_24863;
wire v_24864;
wire v_24865;
wire v_24866;
wire v_24867;
wire v_24868;
wire v_24869;
wire v_24870;
wire v_24871;
wire v_24872;
wire v_24873;
wire v_24874;
wire v_24875;
wire v_24876;
wire v_24877;
wire v_24878;
wire v_24879;
wire v_24880;
wire v_24881;
wire v_24882;
wire v_24883;
wire v_24884;
wire v_24885;
wire v_24886;
wire v_24887;
wire v_24888;
wire v_24889;
wire v_24890;
wire v_24891;
wire v_24892;
wire v_24893;
wire v_24894;
wire v_24895;
wire v_24896;
wire v_24897;
wire v_24898;
wire v_24899;
wire v_24900;
wire v_24901;
wire v_24902;
wire v_24903;
wire v_24904;
wire v_24905;
wire v_24906;
wire v_24907;
wire v_24908;
wire v_24909;
wire v_24910;
wire v_24911;
wire v_24912;
wire v_24913;
wire v_24914;
wire v_24915;
wire v_24916;
wire v_24917;
wire v_24918;
wire v_24919;
wire v_24920;
wire v_24921;
wire v_24922;
wire v_24923;
wire v_24924;
wire v_24925;
wire v_24926;
wire v_24927;
wire v_24928;
wire v_24929;
wire v_24930;
wire v_24931;
wire v_24932;
wire v_24933;
wire v_24934;
wire v_24935;
wire v_24936;
wire v_24937;
wire v_24938;
wire v_24939;
wire v_24940;
wire v_24941;
wire v_24942;
wire v_24943;
wire v_24944;
wire v_24945;
wire v_24946;
wire v_24947;
wire v_24948;
wire v_24949;
wire v_24950;
wire v_24951;
wire v_24952;
wire v_24953;
wire v_24954;
wire v_24955;
wire v_24956;
wire v_24957;
wire v_24958;
wire v_24959;
wire v_24960;
wire v_24961;
wire v_24962;
wire v_24963;
wire v_24964;
wire v_24965;
wire v_24966;
wire v_24967;
wire v_24968;
wire v_24969;
wire v_24970;
wire v_24971;
wire v_24972;
wire v_24973;
wire v_24974;
wire v_24975;
wire v_24976;
wire v_24977;
wire v_24978;
wire v_24979;
wire v_24980;
wire v_24981;
wire v_24982;
wire v_24983;
wire v_24984;
wire v_24985;
wire v_24986;
wire v_24987;
wire v_24988;
wire v_24989;
wire v_24990;
wire v_24991;
wire v_24992;
wire v_24993;
wire v_24994;
wire v_24995;
wire v_24996;
wire v_24997;
wire v_24998;
wire v_24999;
wire v_25000;
wire v_25001;
wire v_25002;
wire v_25003;
wire v_25004;
wire v_25005;
wire v_25006;
wire v_25007;
wire v_25008;
wire v_25009;
wire v_25010;
wire v_25011;
wire v_25012;
wire v_25013;
wire v_25014;
wire v_25015;
wire v_25016;
wire v_25017;
wire v_25018;
wire v_25019;
wire v_25020;
wire v_25021;
wire v_25022;
wire v_25023;
wire v_25024;
wire v_25025;
wire v_25026;
wire v_25027;
wire v_25028;
wire v_25029;
wire v_25030;
wire v_25031;
wire v_25032;
wire v_25033;
wire v_25034;
wire v_25035;
wire v_25036;
wire v_25037;
wire v_25038;
wire v_25039;
wire v_25040;
wire v_25041;
wire v_25042;
wire v_25043;
wire v_25044;
wire v_25045;
wire v_25046;
wire v_25047;
wire v_25048;
wire v_25049;
wire v_25050;
wire v_25051;
wire v_25052;
wire v_25053;
wire v_25054;
wire v_25055;
wire v_25056;
wire v_25057;
wire v_25058;
wire v_25059;
wire v_25060;
wire v_25061;
wire v_25062;
wire v_25063;
wire v_25064;
wire v_25065;
wire v_25066;
wire v_25067;
wire v_25068;
wire v_25069;
wire v_25070;
wire v_25071;
wire v_25072;
wire v_25073;
wire v_25074;
wire v_25075;
wire v_25076;
wire v_25077;
wire v_25078;
wire v_25079;
wire v_25080;
wire v_25081;
wire v_25082;
wire v_25083;
wire v_25084;
wire v_25085;
wire v_25086;
wire v_25087;
wire v_25089;
wire v_25090;
wire v_25091;
wire v_25092;
wire v_25093;
wire v_25094;
wire v_25095;
wire v_25096;
wire v_25097;
wire v_25098;
wire v_25099;
wire v_25100;
wire v_25101;
wire v_25102;
wire v_25103;
wire v_25104;
wire v_25105;
wire v_25106;
wire v_25107;
wire v_25108;
wire v_25109;
wire v_25110;
wire v_25111;
wire v_25112;
wire v_25113;
wire v_25114;
wire v_25115;
wire v_25116;
wire v_25117;
wire v_25118;
wire v_25119;
wire v_25120;
wire v_25121;
wire v_25122;
wire v_25123;
wire v_25124;
wire v_25125;
wire v_25126;
wire v_25127;
wire v_25128;
wire v_25129;
wire v_25130;
wire v_25131;
wire v_25132;
wire v_25133;
wire v_25134;
wire v_25135;
wire v_25136;
wire v_25137;
wire v_25138;
wire v_25139;
wire v_25140;
wire v_25141;
wire v_25142;
wire v_25143;
wire v_25144;
wire v_25145;
wire v_25146;
wire v_25147;
wire v_25148;
wire v_25149;
wire v_25150;
wire v_25151;
wire v_25152;
wire v_25153;
wire v_25154;
wire v_25155;
wire v_25156;
wire v_25157;
wire v_25158;
wire v_25159;
wire v_25160;
wire v_25161;
wire v_25162;
wire v_25163;
wire v_25164;
wire v_25165;
wire v_25166;
wire v_25167;
wire v_25168;
wire v_25169;
wire v_25170;
wire v_25171;
wire v_25172;
wire v_25173;
wire v_25174;
wire v_25175;
wire v_25176;
wire v_25177;
wire v_25178;
wire v_25179;
wire v_25180;
wire v_25181;
wire v_25183;
wire v_25185;
wire v_25186;
wire v_25187;
wire v_25189;
wire v_25190;
wire v_25191;
wire v_25193;
wire v_25194;
wire v_25195;
wire v_25197;
wire v_25198;
wire v_25200;
wire v_25201;
wire v_25202;
wire v_25204;
wire v_25205;
wire v_25206;
wire v_25208;
wire v_25209;
wire v_25210;
wire v_25212;
wire v_25213;
wire v_25214;
wire v_25216;
wire v_25217;
wire v_25218;
wire v_25220;
wire v_25221;
wire v_25222;
wire v_25224;
wire v_25225;
wire v_25226;
wire v_25228;
wire v_25229;
wire v_25230;
wire v_25232;
wire v_25233;
wire v_25234;
wire v_25236;
wire v_25237;
wire v_25238;
wire v_25240;
wire v_25241;
wire v_25242;
wire v_25244;
wire v_25245;
wire v_25246;
wire v_25248;
wire v_25249;
wire v_25250;
wire v_25251;
wire v_25252;
wire v_25253;
wire v_25254;
wire v_25255;
wire v_25256;
wire v_25257;
wire v_25258;
wire v_25259;
wire v_25260;
wire v_25261;
wire v_25262;
wire v_25263;
wire v_25264;
wire v_25265;
wire v_25266;
wire v_25267;
wire v_25268;
wire v_25269;
wire v_25270;
wire v_25271;
wire v_25272;
wire v_25273;
wire v_25274;
wire v_25275;
wire v_25276;
wire v_25277;
wire v_25278;
wire v_25279;
wire v_25280;
wire v_25281;
wire v_25282;
wire v_25283;
wire v_25284;
wire v_25285;
wire v_25286;
wire v_25287;
wire v_25288;
wire v_25289;
wire v_25290;
wire v_25291;
wire v_25292;
wire v_25293;
wire v_25294;
wire v_25295;
wire v_25296;
wire v_25297;
wire v_25298;
wire v_25299;
wire v_25300;
wire v_25301;
wire v_25302;
wire v_25303;
wire v_25304;
wire v_25305;
wire v_25306;
wire v_25307;
wire v_25308;
wire v_25309;
wire v_25310;
wire v_25311;
wire v_25312;
wire v_25313;
wire v_25314;
wire v_25315;
wire v_25316;
wire v_25317;
wire v_25318;
wire v_25319;
wire v_25320;
wire v_25321;
wire v_25322;
wire v_25323;
wire v_25324;
wire v_25325;
wire v_25326;
wire v_25327;
wire v_25328;
wire v_25329;
wire v_25330;
wire v_25331;
wire v_25332;
wire v_25333;
wire v_25334;
wire v_25335;
wire v_25336;
wire v_25337;
wire v_25338;
wire v_25339;
wire v_25340;
wire v_25341;
wire v_25342;
wire v_25343;
wire v_25344;
wire v_25345;
wire v_25346;
wire v_25347;
wire v_25348;
wire v_25349;
wire v_25350;
wire v_25351;
wire v_25352;
wire v_25353;
wire v_25354;
wire v_25355;
wire v_25356;
wire v_25357;
wire v_25358;
wire v_25359;
wire v_25360;
wire v_25361;
wire v_25362;
wire v_25363;
wire v_25364;
wire v_25365;
wire v_25366;
wire v_25367;
wire v_25368;
wire v_25369;
wire v_25370;
wire v_25371;
wire v_25372;
wire v_25373;
wire v_25374;
wire v_25375;
wire v_25376;
wire v_25377;
wire v_25378;
wire v_25379;
wire v_25380;
wire v_25381;
wire v_25382;
wire v_25383;
wire v_25384;
wire v_25385;
wire v_25386;
wire v_25387;
wire v_25388;
wire v_25389;
wire v_25390;
wire v_25391;
wire v_25392;
wire v_25393;
wire v_25394;
wire v_25395;
wire v_25396;
wire v_25397;
wire v_25398;
wire v_25399;
wire v_25400;
wire v_25401;
wire v_25402;
wire v_25403;
wire v_25404;
wire v_25405;
wire v_25406;
wire v_25407;
wire v_25408;
wire v_25409;
wire v_25410;
wire v_25411;
wire v_25412;
wire v_25413;
wire v_25414;
wire v_25415;
wire v_25416;
wire v_25417;
wire v_25418;
wire v_25419;
wire v_25420;
wire v_25421;
wire v_25422;
wire v_25423;
wire v_25424;
wire v_25425;
wire v_25426;
wire v_25427;
wire v_25428;
wire v_25429;
wire v_25430;
wire v_25431;
wire v_25432;
wire v_25433;
wire v_25434;
wire v_25435;
wire v_25436;
wire v_25437;
wire v_25438;
wire v_25439;
wire v_25440;
wire v_25441;
wire v_25443;
wire v_25444;
wire v_25445;
wire v_25446;
wire v_25447;
wire v_25448;
wire v_25449;
wire v_25450;
wire v_25451;
wire v_25452;
wire v_25453;
wire v_25454;
wire v_25455;
wire v_25456;
wire v_25457;
wire v_25458;
wire v_25459;
wire v_25460;
wire v_25461;
wire v_25462;
wire v_25463;
wire v_25464;
wire v_25465;
wire v_25466;
wire v_25467;
wire v_25468;
wire v_25469;
wire v_25470;
wire v_25471;
wire v_25472;
wire v_25473;
wire v_25474;
wire v_25475;
wire v_25476;
wire v_25477;
wire v_25478;
wire v_25479;
wire v_25480;
wire v_25481;
wire v_25482;
wire v_25483;
wire v_25484;
wire v_25485;
wire v_25486;
wire v_25487;
wire v_25488;
wire v_25489;
wire v_25490;
wire v_25491;
wire v_25492;
wire v_25493;
wire v_25494;
wire v_25495;
wire v_25496;
wire v_25497;
wire v_25498;
wire v_25499;
wire v_25500;
wire v_25501;
wire v_25502;
wire v_25503;
wire v_25504;
wire v_25505;
wire v_25506;
wire v_25507;
wire v_25508;
wire v_25509;
wire v_25510;
wire v_25511;
wire v_25512;
wire v_25513;
wire v_25514;
wire v_25515;
wire v_25516;
wire v_25517;
wire v_25518;
wire v_25519;
wire v_25520;
wire v_25521;
wire v_25522;
wire v_25523;
wire v_25524;
wire v_25525;
wire v_25526;
wire v_25527;
wire v_25528;
wire v_25529;
wire v_25530;
wire v_25531;
wire v_25532;
wire v_25533;
wire v_25534;
wire v_25535;
wire v_25536;
wire v_25537;
wire v_25538;
wire v_25539;
wire v_25540;
wire v_25541;
wire v_25542;
wire v_25543;
wire v_25544;
wire v_25545;
wire v_25546;
wire v_25547;
wire v_25548;
wire v_25549;
wire v_25550;
wire v_25551;
wire v_25552;
wire v_25553;
wire v_25554;
wire v_25555;
wire v_25556;
wire v_25557;
wire v_25558;
wire v_25559;
wire v_25560;
wire v_25561;
wire v_25562;
wire v_25563;
wire v_25564;
wire v_25565;
wire v_25566;
wire v_25567;
wire v_25568;
wire v_25569;
wire v_25570;
wire v_25571;
wire v_25572;
wire v_25573;
wire v_25574;
wire v_25575;
wire v_25576;
wire v_25577;
wire v_25578;
wire v_25579;
wire v_25580;
wire v_25581;
wire v_25582;
wire v_25583;
wire v_25584;
wire v_25585;
wire v_25586;
wire v_25587;
wire v_25588;
wire v_25589;
wire v_25590;
wire v_25591;
wire v_25592;
wire v_25593;
wire v_25594;
wire v_25595;
wire v_25596;
wire v_25597;
wire v_25598;
wire v_25599;
wire v_25600;
wire v_25601;
wire v_25602;
wire v_25603;
wire v_25604;
wire v_25605;
wire v_25606;
wire v_25607;
wire v_25608;
wire v_25609;
wire v_25610;
wire v_25611;
wire v_25612;
wire v_25613;
wire v_25614;
wire v_25615;
wire v_25616;
wire v_25617;
wire v_25618;
wire v_25619;
wire v_25620;
wire v_25621;
wire v_25622;
wire v_25623;
wire v_25624;
wire v_25625;
wire v_25626;
wire v_25627;
wire v_25628;
wire v_25629;
wire v_25630;
wire v_25631;
wire v_25632;
wire v_25633;
wire v_25634;
wire v_25635;
wire v_25636;
wire v_25637;
wire v_25638;
wire v_25639;
wire v_25640;
wire v_25641;
wire v_25642;
wire v_25643;
wire v_25644;
wire v_25645;
wire v_25646;
wire v_25647;
wire v_25648;
wire v_25649;
wire v_25650;
wire v_25651;
wire v_25652;
wire v_25653;
wire v_25654;
wire v_25655;
wire v_25656;
wire v_25657;
wire v_25658;
wire v_25659;
wire v_25660;
wire v_25661;
wire v_25662;
wire v_25663;
wire v_25664;
wire v_25665;
wire v_25666;
wire v_25667;
wire v_25668;
wire v_25669;
wire v_25670;
wire v_25671;
wire v_25672;
wire v_25673;
wire v_25674;
wire v_25675;
wire v_25676;
wire v_25677;
wire v_25678;
wire v_25679;
wire v_25680;
wire v_25681;
wire v_25682;
wire v_25683;
wire v_25684;
wire v_25686;
wire v_25687;
wire v_25688;
wire v_25689;
wire v_25690;
wire v_25691;
wire v_25692;
wire v_25693;
wire v_25694;
wire v_25695;
wire v_25696;
wire v_25697;
wire v_25698;
wire v_25699;
wire v_25700;
wire v_25701;
wire v_25702;
wire v_25703;
wire v_25704;
wire v_25705;
wire v_25706;
wire v_25707;
wire v_25708;
wire v_25709;
wire v_25710;
wire v_25711;
wire v_25712;
wire v_25713;
wire v_25714;
wire v_25715;
wire v_25716;
wire v_25717;
wire v_25718;
wire v_25719;
wire v_25720;
wire v_25721;
wire v_25722;
wire v_25723;
wire v_25724;
wire v_25725;
wire v_25726;
wire v_25727;
wire v_25728;
wire v_25729;
wire v_25730;
wire v_25731;
wire v_25732;
wire v_25733;
wire v_25734;
wire v_25735;
wire v_25736;
wire v_25737;
wire v_25738;
wire v_25739;
wire v_25740;
wire v_25741;
wire v_25742;
wire v_25743;
wire v_25744;
wire v_25745;
wire v_25746;
wire v_25747;
wire v_25748;
wire v_25749;
wire v_25750;
wire v_25751;
wire v_25752;
wire v_25753;
wire v_25754;
wire v_25755;
wire v_25756;
wire v_25757;
wire v_25758;
wire v_25759;
wire v_25760;
wire v_25761;
wire v_25762;
wire v_25763;
wire v_25764;
wire v_25765;
wire v_25766;
wire v_25767;
wire v_25768;
wire v_25769;
wire v_25770;
wire v_25771;
wire v_25772;
wire v_25773;
wire v_25774;
wire v_25775;
wire v_25776;
wire v_25777;
wire v_25778;
wire v_25779;
wire v_25780;
wire v_25781;
wire v_25782;
wire v_25783;
wire v_25784;
wire v_25785;
wire v_25786;
wire v_25787;
wire v_25788;
wire v_25789;
wire v_25790;
wire v_25791;
wire v_25792;
wire v_25793;
wire v_25794;
wire v_25795;
wire v_25796;
wire v_25797;
wire v_25798;
wire v_25799;
wire v_25800;
wire v_25801;
wire v_25802;
wire v_25803;
wire v_25804;
wire v_25805;
wire v_25806;
wire v_25807;
wire v_25808;
wire v_25809;
wire v_25810;
wire v_25811;
wire v_25812;
wire v_25813;
wire v_25814;
wire v_25815;
wire v_25816;
wire v_25817;
wire v_25818;
wire v_25819;
wire v_25820;
wire v_25821;
wire v_25822;
wire v_25823;
wire v_25824;
wire v_25825;
wire v_25826;
wire v_25827;
wire v_25828;
wire v_25829;
wire v_25830;
wire v_25831;
wire v_25832;
wire v_25833;
wire v_25834;
wire v_25835;
wire v_25836;
wire v_25837;
wire v_25838;
wire v_25839;
wire v_25840;
wire v_25841;
wire v_25842;
wire v_25843;
wire v_25844;
wire v_25845;
wire v_25846;
wire v_25847;
wire v_25848;
wire v_25849;
wire v_25850;
wire v_25851;
wire v_25852;
wire v_25853;
wire v_25854;
wire v_25855;
wire v_25856;
wire v_25857;
wire v_25858;
wire v_25859;
wire v_25860;
wire v_25861;
wire v_25862;
wire v_25863;
wire v_25864;
wire v_25865;
wire v_25866;
wire v_25867;
wire v_25868;
wire v_25869;
wire v_25870;
wire v_25871;
wire v_25872;
wire v_25873;
wire v_25874;
wire v_25875;
wire v_25876;
wire v_25877;
wire v_25878;
wire v_25879;
wire v_25880;
wire v_25881;
wire v_25882;
wire v_25883;
wire v_25884;
wire v_25885;
wire v_25886;
wire v_25887;
wire v_25888;
wire v_25889;
wire v_25890;
wire v_25891;
wire v_25892;
wire v_25893;
wire v_25894;
wire v_25895;
wire v_25896;
wire v_25897;
wire v_25898;
wire v_25899;
wire v_25900;
wire v_25901;
wire v_25902;
wire v_25903;
wire v_25904;
wire v_25905;
wire v_25906;
wire v_25907;
wire v_25908;
wire v_25909;
wire v_25910;
wire v_25911;
wire v_25912;
wire v_25913;
wire v_25914;
wire v_25915;
wire v_25916;
wire v_25917;
wire v_25918;
wire v_25919;
wire v_25920;
wire v_25921;
wire v_25922;
wire v_25923;
wire v_25924;
wire v_25925;
wire v_25926;
wire v_25927;
wire v_25929;
wire v_25930;
wire v_25931;
wire v_25932;
wire v_25933;
wire v_25934;
wire v_25935;
wire v_25936;
wire v_25937;
wire v_25938;
wire v_25939;
wire v_25940;
wire v_25941;
wire v_25942;
wire v_25943;
wire v_25944;
wire v_25945;
wire v_25946;
wire v_25947;
wire v_25948;
wire v_25949;
wire v_25950;
wire v_25951;
wire v_25952;
wire v_25953;
wire v_25954;
wire v_25955;
wire v_25956;
wire v_25957;
wire v_25958;
wire v_25959;
wire v_25960;
wire v_25961;
wire v_25962;
wire v_25963;
wire v_25964;
wire v_25965;
wire v_25966;
wire v_25967;
wire v_25968;
wire v_25969;
wire v_25970;
wire v_25971;
wire v_25972;
wire v_25973;
wire v_25974;
wire v_25975;
wire v_25976;
wire v_25977;
wire v_25978;
wire v_25979;
wire v_25980;
wire v_25981;
wire v_25982;
wire v_25983;
wire v_25984;
wire v_25985;
wire v_25986;
wire v_25987;
wire v_25988;
wire v_25989;
wire v_25990;
wire v_25991;
wire v_25992;
wire v_25993;
wire v_25994;
wire v_25995;
wire v_25996;
wire v_25997;
wire v_25998;
wire v_25999;
wire v_26000;
wire v_26001;
wire v_26002;
wire v_26003;
wire v_26004;
wire v_26005;
wire v_26006;
wire v_26007;
wire v_26008;
wire v_26009;
wire v_26010;
wire v_26011;
wire v_26012;
wire v_26013;
wire v_26014;
wire v_26015;
wire v_26016;
wire v_26017;
wire v_26018;
wire v_26019;
wire v_26020;
wire v_26021;
wire v_26022;
wire v_26023;
wire v_26024;
wire v_26025;
wire v_26026;
wire v_26027;
wire v_26028;
wire v_26029;
wire v_26030;
wire v_26031;
wire v_26032;
wire v_26033;
wire v_26034;
wire v_26035;
wire v_26036;
wire v_26037;
wire v_26038;
wire v_26039;
wire v_26040;
wire v_26041;
wire v_26042;
wire v_26043;
wire v_26044;
wire v_26045;
wire v_26046;
wire v_26047;
wire v_26048;
wire v_26049;
wire v_26050;
wire v_26051;
wire v_26052;
wire v_26053;
wire v_26054;
wire v_26055;
wire v_26056;
wire v_26057;
wire v_26058;
wire v_26059;
wire v_26060;
wire v_26061;
wire v_26062;
wire v_26063;
wire v_26064;
wire v_26065;
wire v_26066;
wire v_26067;
wire v_26068;
wire v_26069;
wire v_26070;
wire v_26071;
wire v_26072;
wire v_26073;
wire v_26074;
wire v_26075;
wire v_26076;
wire v_26077;
wire v_26078;
wire v_26079;
wire v_26080;
wire v_26081;
wire v_26082;
wire v_26083;
wire v_26084;
wire v_26085;
wire v_26086;
wire v_26087;
wire v_26088;
wire v_26089;
wire v_26090;
wire v_26091;
wire v_26092;
wire v_26093;
wire v_26094;
wire v_26095;
wire v_26096;
wire v_26097;
wire v_26098;
wire v_26099;
wire v_26100;
wire v_26101;
wire v_26102;
wire v_26103;
wire v_26104;
wire v_26105;
wire v_26106;
wire v_26107;
wire v_26108;
wire v_26109;
wire v_26110;
wire v_26111;
wire v_26112;
wire v_26113;
wire v_26114;
wire v_26115;
wire v_26116;
wire v_26117;
wire v_26118;
wire v_26119;
wire v_26120;
wire v_26121;
wire v_26122;
wire v_26123;
wire v_26124;
wire v_26125;
wire v_26126;
wire v_26127;
wire v_26128;
wire v_26129;
wire v_26130;
wire v_26131;
wire v_26132;
wire v_26133;
wire v_26134;
wire v_26135;
wire v_26136;
wire v_26137;
wire v_26138;
wire v_26139;
wire v_26140;
wire v_26141;
wire v_26142;
wire v_26143;
wire v_26144;
wire v_26145;
wire v_26146;
wire v_26147;
wire v_26148;
wire v_26149;
wire v_26150;
wire v_26151;
wire v_26152;
wire v_26153;
wire v_26154;
wire v_26155;
wire v_26156;
wire v_26157;
wire v_26158;
wire v_26159;
wire v_26160;
wire v_26161;
wire v_26162;
wire v_26163;
wire v_26164;
wire v_26165;
wire v_26166;
wire v_26167;
wire v_26168;
wire v_26169;
wire v_26170;
wire v_26172;
wire v_26173;
wire v_26174;
wire v_26175;
wire v_26176;
wire v_26177;
wire v_26178;
wire v_26179;
wire v_26180;
wire v_26181;
wire v_26182;
wire v_26183;
wire v_26184;
wire v_26185;
wire v_26186;
wire v_26187;
wire v_26188;
wire v_26189;
wire v_26190;
wire v_26191;
wire v_26192;
wire v_26193;
wire v_26194;
wire v_26195;
wire v_26196;
wire v_26197;
wire v_26198;
wire v_26199;
wire v_26200;
wire v_26201;
wire v_26202;
wire v_26203;
wire v_26204;
wire v_26205;
wire v_26206;
wire v_26207;
wire v_26208;
wire v_26209;
wire v_26210;
wire v_26211;
wire v_26212;
wire v_26213;
wire v_26214;
wire v_26215;
wire v_26216;
wire v_26217;
wire v_26218;
wire v_26219;
wire v_26220;
wire v_26221;
wire v_26222;
wire v_26223;
wire v_26224;
wire v_26225;
wire v_26226;
wire v_26227;
wire v_26228;
wire v_26229;
wire v_26230;
wire v_26231;
wire v_26232;
wire v_26233;
wire v_26234;
wire v_26235;
wire v_26236;
wire v_26237;
wire v_26238;
wire v_26239;
wire v_26240;
wire v_26241;
wire v_26242;
wire v_26243;
wire v_26244;
wire v_26245;
wire v_26246;
wire v_26247;
wire v_26248;
wire v_26249;
wire v_26250;
wire v_26251;
wire v_26252;
wire v_26253;
wire v_26254;
wire v_26255;
wire v_26256;
wire v_26257;
wire v_26258;
wire v_26259;
wire v_26260;
wire v_26261;
wire v_26262;
wire v_26263;
wire v_26264;
wire v_26265;
wire v_26266;
wire v_26267;
wire v_26268;
wire v_26269;
wire v_26270;
wire v_26271;
wire v_26272;
wire v_26273;
wire v_26274;
wire v_26275;
wire v_26276;
wire v_26277;
wire v_26278;
wire v_26279;
wire v_26280;
wire v_26281;
wire v_26282;
wire v_26283;
wire v_26284;
wire v_26285;
wire v_26286;
wire v_26287;
wire v_26288;
wire v_26289;
wire v_26290;
wire v_26291;
wire v_26292;
wire v_26293;
wire v_26294;
wire v_26295;
wire v_26296;
wire v_26297;
wire v_26298;
wire v_26299;
wire v_26300;
wire v_26301;
wire v_26302;
wire v_26303;
wire v_26304;
wire v_26305;
wire v_26306;
wire v_26307;
wire v_26308;
wire v_26309;
wire v_26310;
wire v_26311;
wire v_26312;
wire v_26313;
wire v_26314;
wire v_26315;
wire v_26316;
wire v_26317;
wire v_26318;
wire v_26319;
wire v_26320;
wire v_26321;
wire v_26322;
wire v_26323;
wire v_26324;
wire v_26325;
wire v_26326;
wire v_26327;
wire v_26328;
wire v_26329;
wire v_26330;
wire v_26331;
wire v_26332;
wire v_26333;
wire v_26334;
wire v_26335;
wire v_26336;
wire v_26337;
wire v_26338;
wire v_26339;
wire v_26340;
wire v_26341;
wire v_26342;
wire v_26343;
wire v_26344;
wire v_26345;
wire v_26346;
wire v_26347;
wire v_26348;
wire v_26349;
wire v_26350;
wire v_26351;
wire v_26352;
wire v_26353;
wire v_26354;
wire v_26355;
wire v_26356;
wire v_26357;
wire v_26358;
wire v_26359;
wire v_26360;
wire v_26361;
wire v_26362;
wire v_26363;
wire v_26364;
wire v_26365;
wire v_26366;
wire v_26367;
wire v_26368;
wire v_26369;
wire v_26370;
wire v_26371;
wire v_26372;
wire v_26373;
wire v_26374;
wire v_26375;
wire v_26376;
wire v_26377;
wire v_26378;
wire v_26379;
wire v_26380;
wire v_26381;
wire v_26382;
wire v_26383;
wire v_26384;
wire v_26385;
wire v_26386;
wire v_26387;
wire v_26388;
wire v_26389;
wire v_26390;
wire v_26391;
wire v_26392;
wire v_26393;
wire v_26394;
wire v_26395;
wire v_26396;
wire v_26397;
wire v_26398;
wire v_26399;
wire v_26400;
wire v_26401;
wire v_26402;
wire v_26403;
wire v_26404;
wire v_26405;
wire v_26406;
wire v_26407;
wire v_26408;
wire v_26409;
wire v_26410;
wire v_26411;
wire v_26412;
wire v_26413;
wire v_26415;
wire v_26416;
wire v_26417;
wire v_26418;
wire v_26419;
wire v_26420;
wire v_26421;
wire v_26422;
wire v_26423;
wire v_26424;
wire v_26425;
wire v_26426;
wire v_26427;
wire v_26428;
wire v_26429;
wire v_26430;
wire v_26431;
wire v_26432;
wire v_26433;
wire v_26434;
wire v_26435;
wire v_26436;
wire v_26437;
wire v_26438;
wire v_26439;
wire v_26440;
wire v_26441;
wire v_26442;
wire v_26443;
wire v_26444;
wire v_26445;
wire v_26446;
wire v_26447;
wire v_26448;
wire v_26449;
wire v_26450;
wire v_26451;
wire v_26452;
wire v_26453;
wire v_26454;
wire v_26455;
wire v_26456;
wire v_26457;
wire v_26458;
wire v_26459;
wire v_26460;
wire v_26461;
wire v_26462;
wire v_26463;
wire v_26464;
wire v_26465;
wire v_26466;
wire v_26467;
wire v_26468;
wire v_26469;
wire v_26470;
wire v_26471;
wire v_26472;
wire v_26473;
wire v_26474;
wire v_26475;
wire v_26476;
wire v_26477;
wire v_26478;
wire v_26479;
wire v_26480;
wire v_26481;
wire v_26482;
wire v_26483;
wire v_26484;
wire v_26485;
wire v_26486;
wire v_26487;
wire v_26488;
wire v_26489;
wire v_26490;
wire v_26491;
wire v_26492;
wire v_26493;
wire v_26494;
wire v_26495;
wire v_26496;
wire v_26497;
wire v_26498;
wire v_26499;
wire v_26500;
wire v_26501;
wire v_26502;
wire v_26503;
wire v_26504;
wire v_26505;
wire v_26506;
wire v_26507;
wire v_26508;
wire v_26509;
wire v_26510;
wire v_26511;
wire v_26512;
wire v_26513;
wire v_26514;
wire v_26515;
wire v_26516;
wire v_26517;
wire v_26518;
wire v_26519;
wire v_26520;
wire v_26521;
wire v_26522;
wire v_26523;
wire v_26524;
wire v_26525;
wire v_26526;
wire v_26527;
wire v_26528;
wire v_26529;
wire v_26530;
wire v_26531;
wire v_26532;
wire v_26533;
wire v_26534;
wire v_26535;
wire v_26536;
wire v_26537;
wire v_26538;
wire v_26539;
wire v_26540;
wire v_26541;
wire v_26542;
wire v_26543;
wire v_26544;
wire v_26545;
wire v_26546;
wire v_26547;
wire v_26548;
wire v_26549;
wire v_26550;
wire v_26551;
wire v_26552;
wire v_26553;
wire v_26554;
wire v_26555;
wire v_26556;
wire v_26557;
wire v_26558;
wire v_26559;
wire v_26560;
wire v_26561;
wire v_26562;
wire v_26563;
wire v_26564;
wire v_26565;
wire v_26566;
wire v_26567;
wire v_26568;
wire v_26569;
wire v_26570;
wire v_26571;
wire v_26572;
wire v_26573;
wire v_26574;
wire v_26575;
wire v_26576;
wire v_26577;
wire v_26578;
wire v_26579;
wire v_26580;
wire v_26581;
wire v_26582;
wire v_26583;
wire v_26584;
wire v_26585;
wire v_26586;
wire v_26587;
wire v_26588;
wire v_26589;
wire v_26590;
wire v_26591;
wire v_26592;
wire v_26593;
wire v_26594;
wire v_26595;
wire v_26596;
wire v_26597;
wire v_26598;
wire v_26599;
wire v_26600;
wire v_26601;
wire v_26602;
wire v_26603;
wire v_26604;
wire v_26605;
wire v_26606;
wire v_26607;
wire v_26608;
wire v_26609;
wire v_26610;
wire v_26611;
wire v_26612;
wire v_26613;
wire v_26614;
wire v_26615;
wire v_26616;
wire v_26617;
wire v_26618;
wire v_26619;
wire v_26620;
wire v_26621;
wire v_26622;
wire v_26623;
wire v_26624;
wire v_26625;
wire v_26626;
wire v_26627;
wire v_26628;
wire v_26629;
wire v_26630;
wire v_26631;
wire v_26632;
wire v_26633;
wire v_26634;
wire v_26635;
wire v_26636;
wire v_26637;
wire v_26638;
wire v_26639;
wire v_26640;
wire v_26641;
wire v_26642;
wire v_26643;
wire v_26644;
wire v_26645;
wire v_26646;
wire v_26647;
wire v_26648;
wire v_26649;
wire v_26650;
wire v_26651;
wire v_26652;
wire v_26653;
wire v_26654;
wire v_26655;
wire v_26656;
wire v_26658;
wire v_26659;
wire v_26660;
wire v_26661;
wire v_26662;
wire v_26663;
wire v_26664;
wire v_26665;
wire v_26666;
wire v_26667;
wire v_26668;
wire v_26669;
wire v_26670;
wire v_26671;
wire v_26672;
wire v_26673;
wire v_26674;
wire v_26675;
wire v_26676;
wire v_26677;
wire v_26678;
wire v_26679;
wire v_26680;
wire v_26681;
wire v_26682;
wire v_26683;
wire v_26684;
wire v_26685;
wire v_26686;
wire v_26687;
wire v_26688;
wire v_26689;
wire v_26690;
wire v_26691;
wire v_26692;
wire v_26693;
wire v_26694;
wire v_26695;
wire v_26696;
wire v_26697;
wire v_26698;
wire v_26699;
wire v_26700;
wire v_26701;
wire v_26702;
wire v_26703;
wire v_26704;
wire v_26705;
wire v_26706;
wire v_26707;
wire v_26708;
wire v_26709;
wire v_26710;
wire v_26711;
wire v_26712;
wire v_26713;
wire v_26714;
wire v_26715;
wire v_26716;
wire v_26717;
wire v_26718;
wire v_26719;
wire v_26720;
wire v_26721;
wire v_26722;
wire v_26723;
wire v_26724;
wire v_26725;
wire v_26726;
wire v_26727;
wire v_26728;
wire v_26729;
wire v_26730;
wire v_26731;
wire v_26732;
wire v_26733;
wire v_26734;
wire v_26735;
wire v_26736;
wire v_26737;
wire v_26738;
wire v_26739;
wire v_26740;
wire v_26741;
wire v_26742;
wire v_26743;
wire v_26744;
wire v_26745;
wire v_26746;
wire v_26747;
wire v_26748;
wire v_26749;
wire v_26750;
wire v_26751;
wire v_26752;
wire v_26753;
wire v_26754;
wire v_26755;
wire v_26756;
wire v_26757;
wire v_26758;
wire v_26759;
wire v_26760;
wire v_26761;
wire v_26762;
wire v_26763;
wire v_26764;
wire v_26765;
wire v_26766;
wire v_26767;
wire v_26768;
wire v_26769;
wire v_26770;
wire v_26771;
wire v_26772;
wire v_26773;
wire v_26774;
wire v_26775;
wire v_26776;
wire v_26777;
wire v_26778;
wire v_26779;
wire v_26780;
wire v_26781;
wire v_26782;
wire v_26783;
wire v_26784;
wire v_26785;
wire v_26786;
wire v_26787;
wire v_26788;
wire v_26789;
wire v_26790;
wire v_26791;
wire v_26792;
wire v_26793;
wire v_26794;
wire v_26795;
wire v_26796;
wire v_26797;
wire v_26798;
wire v_26799;
wire v_26800;
wire v_26801;
wire v_26802;
wire v_26803;
wire v_26804;
wire v_26805;
wire v_26806;
wire v_26807;
wire v_26808;
wire v_26809;
wire v_26810;
wire v_26811;
wire v_26812;
wire v_26813;
wire v_26814;
wire v_26815;
wire v_26816;
wire v_26817;
wire v_26818;
wire v_26819;
wire v_26820;
wire v_26821;
wire v_26822;
wire v_26823;
wire v_26824;
wire v_26825;
wire v_26826;
wire v_26827;
wire v_26828;
wire v_26829;
wire v_26830;
wire v_26831;
wire v_26832;
wire v_26833;
wire v_26834;
wire v_26835;
wire v_26836;
wire v_26837;
wire v_26838;
wire v_26839;
wire v_26840;
wire v_26841;
wire v_26842;
wire v_26843;
wire v_26844;
wire v_26845;
wire v_26846;
wire v_26847;
wire v_26848;
wire v_26849;
wire v_26850;
wire v_26851;
wire v_26852;
wire v_26853;
wire v_26854;
wire v_26855;
wire v_26856;
wire v_26857;
wire v_26858;
wire v_26859;
wire v_26860;
wire v_26861;
wire v_26862;
wire v_26863;
wire v_26864;
wire v_26865;
wire v_26866;
wire v_26867;
wire v_26868;
wire v_26869;
wire v_26870;
wire v_26871;
wire v_26872;
wire v_26873;
wire v_26874;
wire v_26875;
wire v_26876;
wire v_26877;
wire v_26878;
wire v_26879;
wire v_26880;
wire v_26881;
wire v_26882;
wire v_26883;
wire v_26884;
wire v_26885;
wire v_26886;
wire v_26887;
wire v_26888;
wire v_26889;
wire v_26890;
wire v_26891;
wire v_26892;
wire v_26893;
wire v_26894;
wire v_26895;
wire v_26896;
wire v_26897;
wire v_26898;
wire v_26899;
wire v_26901;
wire v_26902;
wire v_26903;
wire v_26904;
wire v_26905;
wire v_26906;
wire v_26907;
wire v_26908;
wire v_26909;
wire v_26910;
wire v_26911;
wire v_26912;
wire v_26913;
wire v_26914;
wire v_26915;
wire v_26916;
wire v_26917;
wire v_26918;
wire v_26919;
wire v_26920;
wire v_26921;
wire v_26922;
wire v_26923;
wire v_26924;
wire v_26925;
wire v_26926;
wire v_26927;
wire v_26928;
wire v_26929;
wire v_26930;
wire v_26931;
wire v_26932;
wire v_26933;
wire v_26934;
wire v_26935;
wire v_26936;
wire v_26937;
wire v_26938;
wire v_26939;
wire v_26940;
wire v_26941;
wire v_26942;
wire v_26943;
wire v_26944;
wire v_26945;
wire v_26946;
wire v_26947;
wire v_26948;
wire v_26949;
wire v_26950;
wire v_26951;
wire v_26952;
wire v_26953;
wire v_26954;
wire v_26955;
wire v_26956;
wire v_26957;
wire v_26958;
wire v_26959;
wire v_26960;
wire v_26961;
wire v_26962;
wire v_26963;
wire v_26964;
wire v_26965;
wire v_26966;
wire v_26967;
wire v_26968;
wire v_26969;
wire v_26970;
wire v_26971;
wire v_26972;
wire v_26973;
wire v_26974;
wire v_26975;
wire v_26976;
wire v_26977;
wire v_26978;
wire v_26979;
wire v_26980;
wire v_26981;
wire v_26982;
wire v_26983;
wire v_26984;
wire v_26985;
wire v_26986;
wire v_26987;
wire v_26988;
wire v_26989;
wire v_26990;
wire v_26991;
wire v_26992;
wire v_26993;
wire v_26994;
wire v_26995;
wire v_26996;
wire v_26997;
wire v_26998;
wire v_26999;
wire v_27000;
wire v_27001;
wire v_27002;
wire v_27003;
wire v_27004;
wire v_27005;
wire v_27006;
wire v_27007;
wire v_27008;
wire v_27009;
wire v_27010;
wire v_27011;
wire v_27012;
wire v_27013;
wire v_27014;
wire v_27015;
wire v_27016;
wire v_27017;
wire v_27018;
wire v_27019;
wire v_27020;
wire v_27021;
wire v_27022;
wire v_27023;
wire v_27024;
wire v_27025;
wire v_27026;
wire v_27027;
wire v_27028;
wire v_27029;
wire v_27030;
wire v_27031;
wire v_27032;
wire v_27033;
wire v_27034;
wire v_27035;
wire v_27036;
wire v_27037;
wire v_27038;
wire v_27039;
wire v_27040;
wire v_27041;
wire v_27042;
wire v_27043;
wire v_27044;
wire v_27045;
wire v_27046;
wire v_27047;
wire v_27048;
wire v_27049;
wire v_27050;
wire v_27051;
wire v_27052;
wire v_27053;
wire v_27054;
wire v_27055;
wire v_27056;
wire v_27057;
wire v_27058;
wire v_27059;
wire v_27060;
wire v_27061;
wire v_27062;
wire v_27063;
wire v_27064;
wire v_27065;
wire v_27066;
wire v_27067;
wire v_27068;
wire v_27069;
wire v_27070;
wire v_27071;
wire v_27072;
wire v_27073;
wire v_27074;
wire v_27075;
wire v_27076;
wire v_27077;
wire v_27078;
wire v_27079;
wire v_27080;
wire v_27081;
wire v_27082;
wire v_27083;
wire v_27084;
wire v_27085;
wire v_27086;
wire v_27087;
wire v_27088;
wire v_27089;
wire v_27090;
wire v_27091;
wire v_27092;
wire v_27093;
wire v_27094;
wire v_27095;
wire v_27096;
wire v_27097;
wire v_27098;
wire v_27099;
wire v_27100;
wire v_27101;
wire v_27102;
wire v_27103;
wire v_27104;
wire v_27105;
wire v_27106;
wire v_27107;
wire v_27108;
wire v_27109;
wire v_27110;
wire v_27111;
wire v_27112;
wire v_27113;
wire v_27114;
wire v_27115;
wire v_27116;
wire v_27117;
wire v_27118;
wire v_27119;
wire v_27120;
wire v_27121;
wire v_27122;
wire v_27123;
wire v_27124;
wire v_27125;
wire v_27126;
wire v_27127;
wire v_27128;
wire v_27129;
wire v_27130;
wire v_27131;
wire v_27132;
wire v_27133;
wire v_27134;
wire v_27135;
wire v_27136;
wire v_27137;
wire v_27138;
wire v_27139;
wire v_27140;
wire v_27141;
wire v_27142;
wire v_27144;
wire v_27145;
wire v_27146;
wire v_27147;
wire v_27148;
wire v_27149;
wire v_27150;
wire v_27151;
wire v_27152;
wire v_27153;
wire v_27154;
wire v_27155;
wire v_27156;
wire v_27157;
wire v_27158;
wire v_27159;
wire v_27160;
wire v_27161;
wire v_27162;
wire v_27163;
wire v_27164;
wire v_27165;
wire v_27166;
wire v_27167;
wire v_27168;
wire v_27169;
wire v_27170;
wire v_27171;
wire v_27172;
wire v_27173;
wire v_27174;
wire v_27175;
wire v_27176;
wire v_27177;
wire v_27178;
wire v_27179;
wire v_27180;
wire v_27181;
wire v_27182;
wire v_27183;
wire v_27184;
wire v_27185;
wire v_27186;
wire v_27187;
wire v_27188;
wire v_27189;
wire v_27190;
wire v_27191;
wire v_27192;
wire v_27193;
wire v_27194;
wire v_27195;
wire v_27196;
wire v_27197;
wire v_27198;
wire v_27199;
wire v_27200;
wire v_27201;
wire v_27202;
wire v_27203;
wire v_27204;
wire v_27205;
wire v_27206;
wire v_27207;
wire v_27208;
wire v_27209;
wire v_27210;
wire v_27211;
wire v_27212;
wire v_27213;
wire v_27214;
wire v_27215;
wire v_27216;
wire v_27217;
wire v_27218;
wire v_27219;
wire v_27220;
wire v_27221;
wire v_27222;
wire v_27223;
wire v_27224;
wire v_27225;
wire v_27226;
wire v_27227;
wire v_27228;
wire v_27229;
wire v_27230;
wire v_27231;
wire v_27232;
wire v_27233;
wire v_27234;
wire v_27235;
wire v_27236;
wire v_27237;
wire v_27238;
wire v_27239;
wire v_27240;
wire v_27241;
wire v_27242;
wire v_27243;
wire v_27244;
wire v_27245;
wire v_27246;
wire v_27247;
wire v_27248;
wire v_27249;
wire v_27250;
wire v_27251;
wire v_27252;
wire v_27253;
wire v_27254;
wire v_27255;
wire v_27256;
wire v_27257;
wire v_27258;
wire v_27259;
wire v_27260;
wire v_27261;
wire v_27262;
wire v_27263;
wire v_27264;
wire v_27265;
wire v_27266;
wire v_27267;
wire v_27268;
wire v_27269;
wire v_27270;
wire v_27271;
wire v_27272;
wire v_27273;
wire v_27274;
wire v_27275;
wire v_27276;
wire v_27277;
wire v_27278;
wire v_27279;
wire v_27280;
wire v_27281;
wire v_27282;
wire v_27283;
wire v_27284;
wire v_27285;
wire v_27286;
wire v_27287;
wire v_27288;
wire v_27289;
wire v_27290;
wire v_27291;
wire v_27292;
wire v_27293;
wire v_27294;
wire v_27295;
wire v_27296;
wire v_27297;
wire v_27298;
wire v_27299;
wire v_27300;
wire v_27301;
wire v_27302;
wire v_27303;
wire v_27304;
wire v_27305;
wire v_27306;
wire v_27307;
wire v_27308;
wire v_27309;
wire v_27310;
wire v_27311;
wire v_27312;
wire v_27313;
wire v_27314;
wire v_27315;
wire v_27316;
wire v_27317;
wire v_27318;
wire v_27319;
wire v_27320;
wire v_27321;
wire v_27322;
wire v_27323;
wire v_27324;
wire v_27325;
wire v_27326;
wire v_27327;
wire v_27328;
wire v_27329;
wire v_27330;
wire v_27331;
wire v_27332;
wire v_27333;
wire v_27334;
wire v_27335;
wire v_27336;
wire v_27337;
wire v_27338;
wire v_27339;
wire v_27340;
wire v_27341;
wire v_27342;
wire v_27343;
wire v_27344;
wire v_27345;
wire v_27346;
wire v_27347;
wire v_27348;
wire v_27349;
wire v_27350;
wire v_27351;
wire v_27352;
wire v_27353;
wire v_27354;
wire v_27355;
wire v_27356;
wire v_27357;
wire v_27358;
wire v_27359;
wire v_27360;
wire v_27361;
wire v_27362;
wire v_27363;
wire v_27364;
wire v_27365;
wire v_27366;
wire v_27367;
wire v_27368;
wire v_27369;
wire v_27370;
wire v_27371;
wire v_27372;
wire v_27373;
wire v_27374;
wire v_27375;
wire v_27376;
wire v_27377;
wire v_27378;
wire v_27379;
wire v_27380;
wire v_27381;
wire v_27382;
wire v_27383;
wire v_27384;
wire v_27385;
wire v_27387;
wire v_27388;
wire v_27389;
wire v_27390;
wire v_27391;
wire v_27392;
wire v_27393;
wire v_27394;
wire v_27395;
wire v_27396;
wire v_27397;
wire v_27398;
wire v_27399;
wire v_27400;
wire v_27401;
wire v_27402;
wire v_27403;
wire v_27404;
wire v_27405;
wire v_27406;
wire v_27407;
wire v_27408;
wire v_27409;
wire v_27410;
wire v_27411;
wire v_27412;
wire v_27413;
wire v_27414;
wire v_27415;
wire v_27416;
wire v_27417;
wire v_27418;
wire v_27419;
wire v_27420;
wire v_27421;
wire v_27422;
wire v_27423;
wire v_27424;
wire v_27425;
wire v_27426;
wire v_27427;
wire v_27428;
wire v_27429;
wire v_27430;
wire v_27431;
wire v_27432;
wire v_27433;
wire v_27434;
wire v_27435;
wire v_27436;
wire v_27437;
wire v_27438;
wire v_27439;
wire v_27440;
wire v_27441;
wire v_27442;
wire v_27443;
wire v_27444;
wire v_27445;
wire v_27446;
wire v_27447;
wire v_27448;
wire v_27449;
wire v_27450;
wire v_27451;
wire v_27452;
wire v_27453;
wire v_27454;
wire v_27455;
wire v_27456;
wire v_27457;
wire v_27458;
wire v_27459;
wire v_27460;
wire v_27461;
wire v_27462;
wire v_27463;
wire v_27464;
wire v_27465;
wire v_27466;
wire v_27467;
wire v_27468;
wire v_27469;
wire v_27470;
wire v_27471;
wire v_27472;
wire v_27473;
wire v_27474;
wire v_27475;
wire v_27476;
wire v_27477;
wire v_27478;
wire v_27479;
wire v_27480;
wire v_27481;
wire v_27482;
wire v_27483;
wire v_27484;
wire v_27485;
wire v_27486;
wire v_27487;
wire v_27488;
wire v_27489;
wire v_27490;
wire v_27491;
wire v_27492;
wire v_27493;
wire v_27494;
wire v_27495;
wire v_27496;
wire v_27497;
wire v_27498;
wire v_27499;
wire v_27500;
wire v_27501;
wire v_27502;
wire v_27503;
wire v_27504;
wire v_27505;
wire v_27506;
wire v_27507;
wire v_27508;
wire v_27509;
wire v_27510;
wire v_27511;
wire v_27512;
wire v_27513;
wire v_27514;
wire v_27515;
wire v_27516;
wire v_27517;
wire v_27518;
wire v_27519;
wire v_27520;
wire v_27521;
wire v_27522;
wire v_27523;
wire v_27524;
wire v_27525;
wire v_27526;
wire v_27527;
wire v_27528;
wire v_27529;
wire v_27530;
wire v_27531;
wire v_27532;
wire v_27533;
wire v_27534;
wire v_27535;
wire v_27536;
wire v_27537;
wire v_27538;
wire v_27539;
wire v_27540;
wire v_27541;
wire v_27542;
wire v_27543;
wire v_27544;
wire v_27545;
wire v_27546;
wire v_27547;
wire v_27548;
wire v_27549;
wire v_27550;
wire v_27551;
wire v_27552;
wire v_27553;
wire v_27554;
wire v_27555;
wire v_27556;
wire v_27557;
wire v_27558;
wire v_27559;
wire v_27560;
wire v_27561;
wire v_27562;
wire v_27563;
wire v_27564;
wire v_27565;
wire v_27566;
wire v_27567;
wire v_27568;
wire v_27569;
wire v_27570;
wire v_27571;
wire v_27572;
wire v_27573;
wire v_27574;
wire v_27575;
wire v_27576;
wire v_27577;
wire v_27578;
wire v_27579;
wire v_27580;
wire v_27581;
wire v_27582;
wire v_27583;
wire v_27584;
wire v_27585;
wire v_27586;
wire v_27587;
wire v_27588;
wire v_27589;
wire v_27590;
wire v_27591;
wire v_27592;
wire v_27593;
wire v_27594;
wire v_27595;
wire v_27596;
wire v_27597;
wire v_27598;
wire v_27599;
wire v_27600;
wire v_27601;
wire v_27602;
wire v_27603;
wire v_27604;
wire v_27605;
wire v_27606;
wire v_27607;
wire v_27608;
wire v_27609;
wire v_27610;
wire v_27611;
wire v_27612;
wire v_27613;
wire v_27614;
wire v_27615;
wire v_27616;
wire v_27617;
wire v_27618;
wire v_27619;
wire v_27620;
wire v_27621;
wire v_27622;
wire v_27623;
wire v_27624;
wire v_27625;
wire v_27626;
wire v_27627;
wire v_27628;
wire v_27630;
wire v_27631;
wire v_27632;
wire v_27633;
wire v_27634;
wire v_27635;
wire v_27636;
wire v_27637;
wire v_27638;
wire v_27639;
wire v_27640;
wire v_27641;
wire v_27642;
wire v_27643;
wire v_27644;
wire v_27645;
wire v_27646;
wire v_27647;
wire v_27648;
wire v_27649;
wire v_27650;
wire v_27651;
wire v_27652;
wire v_27653;
wire v_27654;
wire v_27655;
wire v_27656;
wire v_27657;
wire v_27658;
wire v_27659;
wire v_27660;
wire v_27661;
wire v_27662;
wire v_27663;
wire v_27664;
wire v_27665;
wire v_27666;
wire v_27667;
wire v_27668;
wire v_27669;
wire v_27670;
wire v_27671;
wire v_27672;
wire v_27673;
wire v_27674;
wire v_27675;
wire v_27676;
wire v_27677;
wire v_27678;
wire v_27679;
wire v_27680;
wire v_27681;
wire v_27682;
wire v_27683;
wire v_27684;
wire v_27685;
wire v_27686;
wire v_27687;
wire v_27688;
wire v_27689;
wire v_27690;
wire v_27691;
wire v_27692;
wire v_27693;
wire v_27694;
wire v_27695;
wire v_27696;
wire v_27697;
wire v_27698;
wire v_27699;
wire v_27700;
wire v_27701;
wire v_27702;
wire v_27703;
wire v_27704;
wire v_27705;
wire v_27706;
wire v_27707;
wire v_27708;
wire v_27709;
wire v_27710;
wire v_27711;
wire v_27712;
wire v_27713;
wire v_27714;
wire v_27715;
wire v_27716;
wire v_27717;
wire v_27718;
wire v_27719;
wire v_27720;
wire v_27721;
wire v_27722;
wire v_27723;
wire v_27724;
wire v_27725;
wire v_27726;
wire v_27727;
wire v_27728;
wire v_27729;
wire v_27730;
wire v_27731;
wire v_27732;
wire v_27733;
wire v_27734;
wire v_27735;
wire v_27736;
wire v_27737;
wire v_27738;
wire v_27739;
wire v_27740;
wire v_27741;
wire v_27742;
wire v_27743;
wire v_27744;
wire v_27745;
wire v_27746;
wire v_27747;
wire v_27748;
wire v_27749;
wire v_27750;
wire v_27751;
wire v_27752;
wire v_27753;
wire v_27754;
wire v_27755;
wire v_27756;
wire v_27757;
wire v_27758;
wire v_27759;
wire v_27760;
wire v_27761;
wire v_27762;
wire v_27763;
wire v_27764;
wire v_27765;
wire v_27766;
wire v_27767;
wire v_27768;
wire v_27769;
wire v_27770;
wire v_27771;
wire v_27772;
wire v_27773;
wire v_27774;
wire v_27775;
wire v_27776;
wire v_27777;
wire v_27778;
wire v_27779;
wire v_27780;
wire v_27781;
wire v_27782;
wire v_27783;
wire v_27784;
wire v_27785;
wire v_27786;
wire v_27787;
wire v_27788;
wire v_27789;
wire v_27790;
wire v_27791;
wire v_27792;
wire v_27793;
wire v_27794;
wire v_27795;
wire v_27796;
wire v_27797;
wire v_27798;
wire v_27799;
wire v_27800;
wire v_27801;
wire v_27802;
wire v_27803;
wire v_27804;
wire v_27805;
wire v_27806;
wire v_27807;
wire v_27808;
wire v_27809;
wire v_27810;
wire v_27811;
wire v_27812;
wire v_27813;
wire v_27814;
wire v_27815;
wire v_27816;
wire v_27817;
wire v_27818;
wire v_27819;
wire v_27820;
wire v_27821;
wire v_27822;
wire v_27823;
wire v_27824;
wire v_27825;
wire v_27826;
wire v_27827;
wire v_27828;
wire v_27829;
wire v_27830;
wire v_27831;
wire v_27832;
wire v_27833;
wire v_27834;
wire v_27835;
wire v_27836;
wire v_27837;
wire v_27838;
wire v_27839;
wire v_27840;
wire v_27841;
wire v_27842;
wire v_27843;
wire v_27844;
wire v_27845;
wire v_27846;
wire v_27847;
wire v_27848;
wire v_27849;
wire v_27850;
wire v_27851;
wire v_27852;
wire v_27853;
wire v_27854;
wire v_27855;
wire v_27856;
wire v_27857;
wire v_27858;
wire v_27859;
wire v_27860;
wire v_27861;
wire v_27862;
wire v_27863;
wire v_27864;
wire v_27865;
wire v_27866;
wire v_27867;
wire v_27868;
wire v_27869;
wire v_27870;
wire v_27871;
wire v_27873;
wire v_27874;
wire v_27875;
wire v_27876;
wire v_27877;
wire v_27878;
wire v_27879;
wire v_27880;
wire v_27881;
wire v_27882;
wire v_27883;
wire v_27884;
wire v_27885;
wire v_27886;
wire v_27887;
wire v_27888;
wire v_27889;
wire v_27890;
wire v_27891;
wire v_27892;
wire v_27893;
wire v_27894;
wire v_27895;
wire v_27896;
wire v_27897;
wire v_27898;
wire v_27899;
wire v_27900;
wire v_27901;
wire v_27902;
wire v_27903;
wire v_27904;
wire v_27905;
wire v_27906;
wire v_27907;
wire v_27908;
wire v_27909;
wire v_27910;
wire v_27911;
wire v_27912;
wire v_27913;
wire v_27914;
wire v_27915;
wire v_27916;
wire v_27917;
wire v_27918;
wire v_27919;
wire v_27920;
wire v_27921;
wire v_27922;
wire v_27923;
wire v_27924;
wire v_27925;
wire v_27926;
wire v_27927;
wire v_27928;
wire v_27929;
wire v_27930;
wire v_27931;
wire v_27932;
wire v_27933;
wire v_27934;
wire v_27935;
wire v_27936;
wire v_27937;
wire v_27938;
wire v_27939;
wire v_27940;
wire v_27941;
wire v_27942;
wire v_27943;
wire v_27944;
wire v_27945;
wire v_27946;
wire v_27947;
wire v_27948;
wire v_27949;
wire v_27950;
wire v_27951;
wire v_27952;
wire v_27953;
wire v_27954;
wire v_27955;
wire v_27956;
wire v_27957;
wire v_27958;
wire v_27959;
wire v_27960;
wire v_27961;
wire v_27962;
wire v_27963;
wire v_27964;
wire v_27965;
wire v_27966;
wire v_27967;
wire v_27968;
wire v_27969;
wire v_27970;
wire v_27971;
wire v_27972;
wire v_27973;
wire v_27974;
wire v_27975;
wire v_27976;
wire v_27977;
wire v_27978;
wire v_27979;
wire v_27980;
wire v_27981;
wire v_27982;
wire v_27983;
wire v_27984;
wire v_27985;
wire v_27986;
wire v_27987;
wire v_27988;
wire v_27989;
wire v_27990;
wire v_27991;
wire v_27992;
wire v_27993;
wire v_27994;
wire v_27995;
wire v_27996;
wire v_27997;
wire v_27998;
wire v_27999;
wire v_28000;
wire v_28001;
wire v_28002;
wire v_28003;
wire v_28004;
wire v_28005;
wire v_28006;
wire v_28007;
wire v_28008;
wire v_28009;
wire v_28010;
wire v_28011;
wire v_28012;
wire v_28013;
wire v_28014;
wire v_28015;
wire v_28016;
wire v_28017;
wire v_28018;
wire v_28019;
wire v_28020;
wire v_28021;
wire v_28022;
wire v_28023;
wire v_28024;
wire v_28025;
wire v_28026;
wire v_28027;
wire v_28028;
wire v_28029;
wire v_28030;
wire v_28031;
wire v_28032;
wire v_28033;
wire v_28034;
wire v_28035;
wire v_28036;
wire v_28037;
wire v_28038;
wire v_28039;
wire v_28040;
wire v_28041;
wire v_28042;
wire v_28043;
wire v_28044;
wire v_28045;
wire v_28046;
wire v_28047;
wire v_28048;
wire v_28049;
wire v_28050;
wire v_28051;
wire v_28052;
wire v_28053;
wire v_28054;
wire v_28055;
wire v_28056;
wire v_28057;
wire v_28058;
wire v_28059;
wire v_28060;
wire v_28061;
wire v_28062;
wire v_28063;
wire v_28064;
wire v_28065;
wire v_28066;
wire v_28067;
wire v_28068;
wire v_28069;
wire v_28070;
wire v_28071;
wire v_28072;
wire v_28073;
wire v_28074;
wire v_28075;
wire v_28076;
wire v_28077;
wire v_28078;
wire v_28079;
wire v_28080;
wire v_28081;
wire v_28082;
wire v_28083;
wire v_28084;
wire v_28085;
wire v_28086;
wire v_28087;
wire v_28088;
wire v_28089;
wire v_28090;
wire v_28091;
wire v_28092;
wire v_28093;
wire v_28094;
wire v_28095;
wire v_28096;
wire v_28097;
wire v_28098;
wire v_28099;
wire v_28100;
wire v_28101;
wire v_28102;
wire v_28103;
wire v_28104;
wire v_28105;
wire v_28106;
wire v_28107;
wire v_28108;
wire v_28109;
wire v_28110;
wire v_28111;
wire v_28112;
wire v_28113;
wire v_28114;
wire v_28116;
wire v_28117;
wire v_28118;
wire v_28119;
wire v_28120;
wire v_28121;
wire v_28122;
wire v_28123;
wire v_28124;
wire v_28125;
wire v_28126;
wire v_28127;
wire v_28128;
wire v_28129;
wire v_28130;
wire v_28131;
wire v_28132;
wire v_28133;
wire v_28134;
wire v_28135;
wire v_28136;
wire v_28137;
wire v_28138;
wire v_28139;
wire v_28140;
wire v_28141;
wire v_28142;
wire v_28143;
wire v_28144;
wire v_28145;
wire v_28146;
wire v_28147;
wire v_28148;
wire v_28149;
wire v_28150;
wire v_28151;
wire v_28152;
wire v_28153;
wire v_28154;
wire v_28155;
wire v_28156;
wire v_28157;
wire v_28158;
wire v_28159;
wire v_28160;
wire v_28161;
wire v_28162;
wire v_28163;
wire v_28164;
wire v_28165;
wire v_28166;
wire v_28167;
wire v_28168;
wire v_28169;
wire v_28170;
wire v_28171;
wire v_28172;
wire v_28173;
wire v_28174;
wire v_28175;
wire v_28176;
wire v_28177;
wire v_28178;
wire v_28179;
wire v_28180;
wire v_28181;
wire v_28182;
wire v_28183;
wire v_28184;
wire v_28185;
wire v_28186;
wire v_28187;
wire v_28188;
wire v_28189;
wire v_28190;
wire v_28191;
wire v_28192;
wire v_28193;
wire v_28194;
wire v_28195;
wire v_28196;
wire v_28197;
wire v_28198;
wire v_28199;
wire v_28200;
wire v_28201;
wire v_28202;
wire v_28203;
wire v_28204;
wire v_28205;
wire v_28206;
wire v_28207;
wire v_28208;
wire v_28209;
wire v_28210;
wire v_28211;
wire v_28212;
wire v_28213;
wire v_28214;
wire v_28215;
wire v_28216;
wire v_28217;
wire v_28218;
wire v_28219;
wire v_28220;
wire v_28221;
wire v_28222;
wire v_28223;
wire v_28224;
wire v_28225;
wire v_28226;
wire v_28227;
wire v_28228;
wire v_28229;
wire v_28230;
wire v_28231;
wire v_28232;
wire v_28233;
wire v_28234;
wire v_28235;
wire v_28236;
wire v_28237;
wire v_28238;
wire v_28239;
wire v_28240;
wire v_28241;
wire v_28242;
wire v_28243;
wire v_28244;
wire v_28245;
wire v_28246;
wire v_28247;
wire v_28248;
wire v_28249;
wire v_28250;
wire v_28251;
wire v_28252;
wire v_28253;
wire v_28254;
wire v_28255;
wire v_28256;
wire v_28257;
wire v_28258;
wire v_28259;
wire v_28260;
wire v_28261;
wire v_28262;
wire v_28263;
wire v_28264;
wire v_28265;
wire v_28266;
wire v_28267;
wire v_28268;
wire v_28269;
wire v_28270;
wire v_28271;
wire v_28272;
wire v_28273;
wire v_28274;
wire v_28275;
wire v_28276;
wire v_28277;
wire v_28278;
wire v_28279;
wire v_28280;
wire v_28281;
wire v_28282;
wire v_28283;
wire v_28284;
wire v_28285;
wire v_28286;
wire v_28287;
wire v_28288;
wire v_28289;
wire v_28290;
wire v_28291;
wire v_28292;
wire v_28293;
wire v_28294;
wire v_28295;
wire v_28296;
wire v_28297;
wire v_28298;
wire v_28299;
wire v_28300;
wire v_28301;
wire v_28302;
wire v_28303;
wire v_28304;
wire v_28305;
wire v_28306;
wire v_28307;
wire v_28308;
wire v_28309;
wire v_28310;
wire v_28311;
wire v_28312;
wire v_28313;
wire v_28314;
wire v_28315;
wire v_28316;
wire v_28317;
wire v_28318;
wire v_28319;
wire v_28320;
wire v_28321;
wire v_28322;
wire v_28323;
wire v_28324;
wire v_28325;
wire v_28326;
wire v_28327;
wire v_28328;
wire v_28329;
wire v_28330;
wire v_28331;
wire v_28332;
wire v_28333;
wire v_28334;
wire v_28335;
wire v_28336;
wire v_28337;
wire v_28338;
wire v_28339;
wire v_28340;
wire v_28341;
wire v_28342;
wire v_28343;
wire v_28344;
wire v_28345;
wire v_28346;
wire v_28347;
wire v_28348;
wire v_28349;
wire v_28350;
wire v_28351;
wire v_28352;
wire v_28353;
wire v_28354;
wire v_28355;
wire v_28356;
wire v_28357;
wire v_28359;
wire v_28360;
wire v_28361;
wire v_28362;
wire v_28363;
wire v_28364;
wire v_28365;
wire v_28366;
wire v_28367;
wire v_28368;
wire v_28369;
wire v_28370;
wire v_28371;
wire v_28372;
wire v_28373;
wire v_28374;
wire v_28375;
wire v_28376;
wire v_28377;
wire v_28378;
wire v_28379;
wire v_28380;
wire v_28381;
wire v_28382;
wire v_28383;
wire v_28384;
wire v_28385;
wire v_28386;
wire v_28387;
wire v_28388;
wire v_28389;
wire v_28390;
wire v_28391;
wire v_28392;
wire v_28393;
wire v_28394;
wire v_28395;
wire v_28396;
wire v_28397;
wire v_28398;
wire v_28399;
wire v_28400;
wire v_28401;
wire v_28402;
wire v_28403;
wire v_28404;
wire v_28405;
wire v_28406;
wire v_28407;
wire v_28408;
wire v_28409;
wire v_28410;
wire v_28411;
wire v_28412;
wire v_28413;
wire v_28414;
wire v_28415;
wire v_28416;
wire v_28417;
wire v_28418;
wire v_28419;
wire v_28420;
wire v_28421;
wire v_28422;
wire v_28423;
wire v_28424;
wire v_28425;
wire v_28426;
wire v_28427;
wire v_28428;
wire v_28429;
wire v_28430;
wire v_28431;
wire v_28432;
wire v_28433;
wire v_28434;
wire v_28435;
wire v_28436;
wire v_28437;
wire v_28438;
wire v_28439;
wire v_28440;
wire v_28441;
wire v_28442;
wire v_28443;
wire v_28444;
wire v_28445;
wire v_28446;
wire v_28447;
wire v_28448;
wire v_28449;
wire v_28450;
wire v_28451;
wire v_28452;
wire v_28453;
wire v_28454;
wire v_28455;
wire v_28456;
wire v_28457;
wire v_28458;
wire v_28459;
wire v_28460;
wire v_28461;
wire v_28462;
wire v_28463;
wire v_28464;
wire v_28465;
wire v_28466;
wire v_28467;
wire v_28468;
wire v_28469;
wire v_28470;
wire v_28471;
wire v_28472;
wire v_28473;
wire v_28474;
wire v_28475;
wire v_28476;
wire v_28477;
wire v_28478;
wire v_28479;
wire v_28480;
wire v_28481;
wire v_28482;
wire v_28483;
wire v_28484;
wire v_28485;
wire v_28486;
wire v_28487;
wire v_28488;
wire v_28489;
wire v_28490;
wire v_28491;
wire v_28492;
wire v_28493;
wire v_28494;
wire v_28495;
wire v_28496;
wire v_28497;
wire v_28498;
wire v_28499;
wire v_28500;
wire v_28501;
wire v_28502;
wire v_28503;
wire v_28504;
wire v_28505;
wire v_28506;
wire v_28507;
wire v_28508;
wire v_28509;
wire v_28510;
wire v_28511;
wire v_28512;
wire v_28513;
wire v_28514;
wire v_28515;
wire v_28516;
wire v_28517;
wire v_28518;
wire v_28519;
wire v_28520;
wire v_28521;
wire v_28522;
wire v_28523;
wire v_28524;
wire v_28525;
wire v_28526;
wire v_28527;
wire v_28528;
wire v_28529;
wire v_28530;
wire v_28531;
wire v_28532;
wire v_28533;
wire v_28534;
wire v_28535;
wire v_28536;
wire v_28537;
wire v_28538;
wire v_28539;
wire v_28540;
wire v_28541;
wire v_28542;
wire v_28543;
wire v_28544;
wire v_28545;
wire v_28546;
wire v_28547;
wire v_28548;
wire v_28549;
wire v_28550;
wire v_28551;
wire v_28552;
wire v_28553;
wire v_28554;
wire v_28555;
wire v_28556;
wire v_28557;
wire v_28558;
wire v_28559;
wire v_28560;
wire v_28561;
wire v_28562;
wire v_28563;
wire v_28564;
wire v_28565;
wire v_28566;
wire v_28567;
wire v_28568;
wire v_28569;
wire v_28570;
wire v_28571;
wire v_28572;
wire v_28573;
wire v_28574;
wire v_28575;
wire v_28576;
wire v_28577;
wire v_28578;
wire v_28579;
wire v_28580;
wire v_28581;
wire v_28582;
wire v_28583;
wire v_28584;
wire v_28585;
wire v_28586;
wire v_28587;
wire v_28588;
wire v_28589;
wire v_28590;
wire v_28591;
wire v_28592;
wire v_28593;
wire v_28594;
wire v_28595;
wire v_28596;
wire v_28597;
wire v_28598;
wire v_28599;
wire v_28600;
wire v_28602;
wire v_28603;
wire v_28604;
wire v_28605;
wire v_28606;
wire v_28607;
wire v_28608;
wire v_28609;
wire v_28610;
wire v_28611;
wire v_28612;
wire v_28613;
wire v_28614;
wire v_28615;
wire v_28616;
wire v_28617;
wire v_28618;
wire v_28619;
wire v_28620;
wire v_28621;
wire v_28622;
wire v_28623;
wire v_28624;
wire v_28625;
wire v_28626;
wire v_28627;
wire v_28628;
wire v_28629;
wire v_28630;
wire v_28631;
wire v_28632;
wire v_28633;
wire v_28634;
wire v_28635;
wire v_28636;
wire v_28637;
wire v_28638;
wire v_28639;
wire v_28640;
wire v_28641;
wire v_28642;
wire v_28643;
wire v_28644;
wire v_28645;
wire v_28646;
wire v_28647;
wire v_28648;
wire v_28649;
wire v_28650;
wire v_28651;
wire v_28652;
wire v_28653;
wire v_28654;
wire v_28655;
wire v_28656;
wire v_28657;
wire v_28658;
wire v_28659;
wire v_28660;
wire v_28661;
wire v_28662;
wire v_28663;
wire v_28664;
wire v_28665;
wire v_28666;
wire v_28667;
wire v_28668;
wire v_28669;
wire v_28670;
wire v_28671;
wire v_28672;
wire v_28673;
wire v_28674;
wire v_28675;
wire v_28676;
wire v_28677;
wire v_28678;
wire v_28679;
wire v_28680;
wire v_28681;
wire v_28682;
wire v_28683;
wire v_28684;
wire v_28685;
wire v_28686;
wire v_28687;
wire v_28688;
wire v_28689;
wire v_28690;
wire v_28691;
wire v_28692;
wire v_28693;
wire v_28694;
wire v_28695;
wire v_28696;
wire v_28697;
wire v_28698;
wire v_28699;
wire v_28700;
wire v_28701;
wire v_28702;
wire v_28703;
wire v_28704;
wire v_28705;
wire v_28706;
wire v_28707;
wire v_28708;
wire v_28709;
wire v_28710;
wire v_28711;
wire v_28712;
wire v_28713;
wire v_28714;
wire v_28715;
wire v_28716;
wire v_28717;
wire v_28718;
wire v_28719;
wire v_28720;
wire v_28721;
wire v_28722;
wire v_28723;
wire v_28724;
wire v_28725;
wire v_28726;
wire v_28727;
wire v_28728;
wire v_28729;
wire v_28730;
wire v_28731;
wire v_28732;
wire v_28733;
wire v_28734;
wire v_28735;
wire v_28736;
wire v_28737;
wire v_28738;
wire v_28739;
wire v_28740;
wire v_28741;
wire v_28742;
wire v_28743;
wire v_28744;
wire v_28745;
wire v_28746;
wire v_28747;
wire v_28748;
wire v_28749;
wire v_28750;
wire v_28751;
wire v_28752;
wire v_28753;
wire v_28754;
wire v_28755;
wire v_28756;
wire v_28757;
wire v_28758;
wire v_28759;
wire v_28760;
wire v_28761;
wire v_28762;
wire v_28763;
wire v_28764;
wire v_28765;
wire v_28766;
wire v_28767;
wire v_28768;
wire v_28769;
wire v_28770;
wire v_28771;
wire v_28772;
wire v_28773;
wire v_28774;
wire v_28775;
wire v_28776;
wire v_28777;
wire v_28778;
wire v_28779;
wire v_28780;
wire v_28781;
wire v_28782;
wire v_28783;
wire v_28784;
wire v_28785;
wire v_28786;
wire v_28787;
wire v_28788;
wire v_28789;
wire v_28790;
wire v_28791;
wire v_28792;
wire v_28793;
wire v_28794;
wire v_28795;
wire v_28796;
wire v_28797;
wire v_28798;
wire v_28799;
wire v_28800;
wire v_28801;
wire v_28802;
wire v_28803;
wire v_28804;
wire v_28805;
wire v_28806;
wire v_28807;
wire v_28808;
wire v_28809;
wire v_28810;
wire v_28811;
wire v_28812;
wire v_28813;
wire v_28814;
wire v_28815;
wire v_28816;
wire v_28817;
wire v_28818;
wire v_28819;
wire v_28820;
wire v_28821;
wire v_28822;
wire v_28823;
wire v_28824;
wire v_28825;
wire v_28826;
wire v_28827;
wire v_28828;
wire v_28829;
wire v_28830;
wire v_28831;
wire v_28832;
wire v_28833;
wire v_28834;
wire v_28835;
wire v_28836;
wire v_28837;
wire v_28838;
wire v_28839;
wire v_28840;
wire v_28841;
wire v_28842;
wire v_28843;
wire v_28845;
wire v_28846;
wire v_28847;
wire v_28848;
wire v_28849;
wire v_28850;
wire v_28851;
wire v_28852;
wire v_28853;
wire v_28854;
wire v_28855;
wire v_28856;
wire v_28857;
wire v_28858;
wire v_28859;
wire v_28860;
wire v_28861;
wire v_28862;
wire v_28863;
wire v_28864;
wire v_28865;
wire v_28866;
wire v_28867;
wire v_28868;
wire v_28869;
wire v_28870;
wire v_28871;
wire v_28872;
wire v_28873;
wire v_28874;
wire v_28875;
wire v_28876;
wire v_28877;
wire v_28878;
wire v_28879;
wire v_28880;
wire v_28881;
wire v_28882;
wire v_28883;
wire v_28884;
wire v_28885;
wire v_28886;
wire v_28887;
wire v_28888;
wire v_28889;
wire v_28890;
wire v_28891;
wire v_28892;
wire v_28893;
wire v_28894;
wire v_28895;
wire v_28896;
wire v_28897;
wire v_28898;
wire v_28899;
wire v_28900;
wire v_28901;
wire v_28902;
wire v_28903;
wire v_28904;
wire v_28905;
wire v_28906;
wire v_28907;
wire v_28908;
wire v_28909;
wire v_28910;
wire v_28911;
wire v_28912;
wire v_28913;
wire v_28914;
wire v_28915;
wire v_28916;
wire v_28917;
wire v_28918;
wire v_28919;
wire v_28920;
wire v_28921;
wire v_28922;
wire v_28923;
wire v_28924;
wire v_28925;
wire v_28926;
wire v_28927;
wire v_28928;
wire v_28929;
wire v_28930;
wire v_28931;
wire v_28932;
wire v_28933;
wire v_28934;
wire v_28935;
wire v_28936;
wire v_28937;
wire v_28938;
wire v_28939;
wire v_28940;
wire v_28941;
wire v_28942;
wire v_28943;
wire v_28944;
wire v_28945;
wire v_28946;
wire v_28947;
wire v_28948;
wire v_28949;
wire v_28950;
wire v_28951;
wire v_28952;
wire v_28953;
wire v_28954;
wire v_28955;
wire v_28956;
wire v_28957;
wire v_28958;
wire v_28959;
wire v_28960;
wire v_28961;
wire v_28962;
wire v_28963;
wire v_28964;
wire v_28965;
wire v_28966;
wire v_28967;
wire v_28968;
wire v_28969;
wire v_28970;
wire v_28971;
wire v_28972;
wire v_28973;
wire v_28974;
wire v_28975;
wire v_28976;
wire v_28977;
wire v_28978;
wire v_28979;
wire v_28980;
wire v_28981;
wire v_28982;
wire v_28983;
wire v_28984;
wire v_28985;
wire v_28986;
wire v_28987;
wire v_28988;
wire v_28989;
wire v_28990;
wire v_28991;
wire v_28992;
wire v_28993;
wire v_28994;
wire v_28995;
wire v_28996;
wire v_28997;
wire v_28998;
wire v_28999;
wire v_29000;
wire v_29001;
wire v_29002;
wire v_29003;
wire v_29004;
wire v_29005;
wire v_29006;
wire v_29007;
wire v_29008;
wire v_29009;
wire v_29010;
wire v_29011;
wire v_29012;
wire v_29013;
wire v_29014;
wire v_29015;
wire v_29016;
wire v_29017;
wire v_29018;
wire v_29019;
wire v_29020;
wire v_29021;
wire v_29022;
wire v_29023;
wire v_29024;
wire v_29025;
wire v_29026;
wire v_29027;
wire v_29028;
wire v_29029;
wire v_29030;
wire v_29031;
wire v_29032;
wire v_29033;
wire v_29034;
wire v_29035;
wire v_29036;
wire v_29037;
wire v_29038;
wire v_29039;
wire v_29040;
wire v_29041;
wire v_29042;
wire v_29043;
wire v_29044;
wire v_29045;
wire v_29046;
wire v_29047;
wire v_29048;
wire v_29049;
wire v_29050;
wire v_29051;
wire v_29052;
wire v_29053;
wire v_29054;
wire v_29055;
wire v_29056;
wire v_29057;
wire v_29058;
wire v_29059;
wire v_29060;
wire v_29061;
wire v_29062;
wire v_29063;
wire v_29064;
wire v_29065;
wire v_29066;
wire v_29067;
wire v_29068;
wire v_29069;
wire v_29070;
wire v_29071;
wire v_29072;
wire v_29073;
wire v_29074;
wire v_29075;
wire v_29076;
wire v_29077;
wire v_29078;
wire v_29079;
wire v_29080;
wire v_29081;
wire v_29082;
wire v_29083;
wire v_29084;
wire v_29085;
wire v_29086;
wire v_29087;
wire v_29088;
wire v_29089;
wire v_29090;
wire v_29091;
wire v_29092;
wire v_29093;
wire v_29094;
wire v_29095;
wire v_29096;
wire v_29097;
wire v_29098;
wire v_29099;
wire v_29100;
wire v_29101;
wire v_29102;
wire v_29103;
wire v_29104;
wire v_29105;
wire v_29106;
wire v_29107;
wire v_29108;
wire v_29109;
wire v_29110;
wire v_29111;
wire v_29112;
wire v_29113;
wire v_29114;
wire v_29115;
wire v_29116;
wire v_29117;
wire v_29118;
wire v_29119;
wire v_29120;
wire v_29121;
wire v_29122;
wire v_29123;
wire v_29124;
wire v_29125;
wire v_29126;
wire v_29127;
wire v_29128;
wire v_29129;
wire v_29130;
wire v_29131;
wire v_29132;
wire v_29133;
wire v_29134;
wire v_29135;
wire v_29136;
wire v_29137;
wire v_29138;
wire v_29139;
wire v_29140;
wire v_29141;
wire v_29142;
wire v_29143;
wire v_29144;
wire v_29145;
wire v_29146;
wire v_29147;
wire v_29148;
wire v_29149;
wire v_29150;
wire v_29151;
wire v_29152;
wire v_29153;
wire v_29154;
wire v_29155;
wire v_29156;
wire v_29157;
wire v_29158;
wire v_29159;
wire v_29160;
wire v_29161;
wire v_29162;
wire v_29163;
wire v_29164;
wire v_29165;
wire v_29166;
wire v_29167;
wire v_29168;
wire v_29169;
wire v_29170;
wire v_29171;
wire v_29172;
wire v_29173;
wire v_29174;
wire v_29175;
wire v_29176;
wire v_29177;
wire v_29178;
wire v_29179;
wire v_29180;
wire v_29181;
wire v_29182;
wire v_29183;
wire v_29184;
wire v_29185;
wire v_29186;
wire v_29187;
wire v_29188;
wire v_29189;
wire v_29190;
wire v_29191;
wire v_29192;
wire v_29193;
wire v_29194;
wire v_29195;
wire v_29196;
wire v_29197;
wire v_29198;
wire v_29199;
wire v_29200;
wire v_29201;
wire v_29202;
wire v_29203;
wire v_29204;
wire v_29205;
wire v_29206;
wire v_29207;
wire v_29208;
wire v_29209;
wire v_29210;
wire v_29211;
wire v_29212;
wire v_29213;
wire v_29214;
wire v_29215;
wire v_29216;
wire v_29217;
wire v_29218;
wire v_29219;
wire v_29220;
wire v_29221;
wire v_29222;
wire v_29223;
wire v_29224;
wire v_29225;
wire v_29226;
wire v_29227;
wire v_29228;
wire v_29229;
wire v_29230;
wire v_29231;
wire v_29232;
wire v_29233;
wire v_29234;
wire v_29235;
wire v_29237;
wire v_29238;
wire v_29239;
wire v_29240;
wire v_29241;
wire v_29242;
wire v_29243;
wire v_29244;
wire v_29245;
wire v_29246;
wire v_29247;
wire v_29248;
wire v_29249;
wire v_29250;
wire v_29251;
wire v_29252;
wire v_29253;
wire v_29254;
wire v_29255;
wire v_29256;
wire v_29257;
wire v_29258;
wire v_29259;
wire v_29260;
wire v_29261;
wire v_29262;
wire v_29263;
wire v_29264;
wire v_29265;
wire v_29266;
wire v_29267;
wire v_29268;
wire v_29269;
wire v_29270;
wire v_29271;
wire v_29272;
wire v_29273;
wire v_29274;
wire v_29275;
wire v_29276;
wire v_29277;
wire v_29278;
wire v_29279;
wire v_29280;
wire v_29281;
wire v_29282;
wire v_29283;
wire v_29284;
wire v_29285;
wire v_29286;
wire v_29287;
wire v_29288;
wire v_29289;
wire v_29290;
wire v_29291;
wire v_29292;
wire v_29293;
wire v_29294;
wire v_29295;
wire v_29296;
wire v_29297;
wire v_29298;
wire v_29299;
wire v_29300;
wire v_29301;
wire v_29302;
wire v_29303;
wire v_29304;
wire v_29305;
wire v_29306;
wire v_29307;
wire v_29308;
wire v_29309;
wire v_29310;
wire v_29311;
wire v_29312;
wire v_29313;
wire v_29314;
wire v_29315;
wire v_29316;
wire v_29317;
wire v_29318;
wire v_29319;
wire v_29320;
wire v_29321;
wire v_29322;
wire v_29323;
wire v_29324;
wire v_29325;
wire v_29326;
wire v_29327;
wire v_29328;
wire v_29329;
wire v_29331;
wire v_29333;
wire v_29334;
wire v_29335;
wire v_29337;
wire v_29338;
wire v_29339;
wire v_29341;
wire v_29342;
wire v_29343;
wire v_29345;
wire v_29346;
wire v_29348;
wire v_29349;
wire v_29350;
wire v_29352;
wire v_29353;
wire v_29354;
wire v_29356;
wire v_29357;
wire v_29358;
wire v_29360;
wire v_29361;
wire v_29362;
wire v_29364;
wire v_29365;
wire v_29366;
wire v_29368;
wire v_29369;
wire v_29370;
wire v_29372;
wire v_29373;
wire v_29374;
wire v_29376;
wire v_29377;
wire v_29378;
wire v_29380;
wire v_29381;
wire v_29382;
wire v_29384;
wire v_29385;
wire v_29386;
wire v_29388;
wire v_29389;
wire v_29390;
wire v_29392;
wire v_29393;
wire v_29394;
wire v_29396;
wire v_29397;
wire v_29398;
wire v_29399;
wire v_29400;
wire v_29401;
wire v_29402;
wire v_29403;
wire v_29404;
wire v_29405;
wire v_29406;
wire v_29407;
wire v_29408;
wire v_29409;
wire v_29410;
wire v_29411;
wire v_29412;
wire v_29413;
wire v_29414;
wire v_29415;
wire v_29416;
wire v_29417;
wire v_29418;
wire v_29419;
wire v_29420;
wire v_29421;
wire v_29422;
wire v_29423;
wire v_29424;
wire v_29425;
wire v_29426;
wire v_29427;
wire v_29428;
wire v_29429;
wire v_29430;
wire v_29431;
wire v_29432;
wire v_29433;
wire v_29434;
wire v_29435;
wire v_29436;
wire v_29437;
wire v_29438;
wire v_29439;
wire v_29440;
wire v_29441;
wire v_29442;
wire v_29443;
wire v_29444;
wire v_29445;
wire v_29446;
wire v_29447;
wire v_29448;
wire v_29449;
wire v_29450;
wire v_29451;
wire v_29452;
wire v_29453;
wire v_29454;
wire v_29455;
wire v_29456;
wire v_29457;
wire v_29458;
wire v_29459;
wire v_29460;
wire v_29461;
wire v_29462;
wire v_29463;
wire v_29464;
wire v_29465;
wire v_29466;
wire v_29467;
wire v_29468;
wire v_29469;
wire v_29470;
wire v_29471;
wire v_29472;
wire v_29473;
wire v_29474;
wire v_29475;
wire v_29476;
wire v_29477;
wire v_29478;
wire v_29479;
wire v_29480;
wire v_29481;
wire v_29482;
wire v_29483;
wire v_29484;
wire v_29485;
wire v_29486;
wire v_29487;
wire v_29488;
wire v_29489;
wire v_29490;
wire v_29491;
wire v_29492;
wire v_29493;
wire v_29494;
wire v_29495;
wire v_29496;
wire v_29497;
wire v_29498;
wire v_29499;
wire v_29500;
wire v_29501;
wire v_29502;
wire v_29503;
wire v_29504;
wire v_29505;
wire v_29506;
wire v_29507;
wire v_29508;
wire v_29509;
wire v_29510;
wire v_29511;
wire v_29512;
wire v_29513;
wire v_29514;
wire v_29515;
wire v_29516;
wire v_29517;
wire v_29518;
wire v_29519;
wire v_29520;
wire v_29521;
wire v_29522;
wire v_29523;
wire v_29524;
wire v_29525;
wire v_29526;
wire v_29527;
wire v_29528;
wire v_29529;
wire v_29530;
wire v_29531;
wire v_29532;
wire v_29533;
wire v_29534;
wire v_29535;
wire v_29536;
wire v_29537;
wire v_29538;
wire v_29539;
wire v_29540;
wire v_29541;
wire v_29542;
wire v_29543;
wire v_29544;
wire v_29545;
wire v_29546;
wire v_29547;
wire v_29548;
wire v_29549;
wire v_29550;
wire v_29551;
wire v_29552;
wire v_29553;
wire v_29554;
wire v_29555;
wire v_29556;
wire v_29557;
wire v_29558;
wire v_29559;
wire v_29560;
wire v_29561;
wire v_29562;
wire v_29563;
wire v_29564;
wire v_29565;
wire v_29566;
wire v_29567;
wire v_29568;
wire v_29569;
wire v_29570;
wire v_29571;
wire v_29572;
wire v_29573;
wire v_29574;
wire v_29575;
wire v_29576;
wire v_29577;
wire v_29578;
wire v_29579;
wire v_29580;
wire v_29581;
wire v_29582;
wire v_29583;
wire v_29584;
wire v_29585;
wire v_29586;
wire v_29587;
wire v_29588;
wire v_29589;
wire v_29591;
wire v_29592;
wire v_29593;
wire v_29594;
wire v_29595;
wire v_29596;
wire v_29597;
wire v_29598;
wire v_29599;
wire v_29600;
wire v_29601;
wire v_29602;
wire v_29603;
wire v_29604;
wire v_29605;
wire v_29606;
wire v_29607;
wire v_29608;
wire v_29609;
wire v_29610;
wire v_29611;
wire v_29612;
wire v_29613;
wire v_29614;
wire v_29615;
wire v_29616;
wire v_29617;
wire v_29618;
wire v_29619;
wire v_29620;
wire v_29621;
wire v_29622;
wire v_29623;
wire v_29624;
wire v_29625;
wire v_29626;
wire v_29627;
wire v_29628;
wire v_29629;
wire v_29630;
wire v_29631;
wire v_29632;
wire v_29633;
wire v_29634;
wire v_29635;
wire v_29636;
wire v_29637;
wire v_29638;
wire v_29639;
wire v_29640;
wire v_29641;
wire v_29642;
wire v_29643;
wire v_29644;
wire v_29645;
wire v_29646;
wire v_29647;
wire v_29648;
wire v_29649;
wire v_29650;
wire v_29651;
wire v_29652;
wire v_29653;
wire v_29654;
wire v_29655;
wire v_29656;
wire v_29657;
wire v_29658;
wire v_29659;
wire v_29660;
wire v_29661;
wire v_29662;
wire v_29663;
wire v_29664;
wire v_29665;
wire v_29666;
wire v_29667;
wire v_29668;
wire v_29669;
wire v_29670;
wire v_29671;
wire v_29672;
wire v_29673;
wire v_29674;
wire v_29675;
wire v_29676;
wire v_29677;
wire v_29678;
wire v_29679;
wire v_29680;
wire v_29681;
wire v_29682;
wire v_29683;
wire v_29684;
wire v_29685;
wire v_29686;
wire v_29687;
wire v_29688;
wire v_29689;
wire v_29690;
wire v_29691;
wire v_29692;
wire v_29693;
wire v_29694;
wire v_29695;
wire v_29696;
wire v_29697;
wire v_29698;
wire v_29699;
wire v_29700;
wire v_29701;
wire v_29702;
wire v_29703;
wire v_29704;
wire v_29705;
wire v_29706;
wire v_29707;
wire v_29708;
wire v_29709;
wire v_29710;
wire v_29711;
wire v_29712;
wire v_29713;
wire v_29714;
wire v_29715;
wire v_29716;
wire v_29717;
wire v_29718;
wire v_29719;
wire v_29720;
wire v_29721;
wire v_29722;
wire v_29723;
wire v_29724;
wire v_29725;
wire v_29726;
wire v_29727;
wire v_29728;
wire v_29729;
wire v_29730;
wire v_29731;
wire v_29732;
wire v_29733;
wire v_29734;
wire v_29735;
wire v_29736;
wire v_29737;
wire v_29738;
wire v_29739;
wire v_29740;
wire v_29741;
wire v_29742;
wire v_29743;
wire v_29744;
wire v_29745;
wire v_29746;
wire v_29747;
wire v_29748;
wire v_29749;
wire v_29750;
wire v_29751;
wire v_29752;
wire v_29753;
wire v_29754;
wire v_29755;
wire v_29756;
wire v_29757;
wire v_29758;
wire v_29759;
wire v_29760;
wire v_29761;
wire v_29762;
wire v_29763;
wire v_29764;
wire v_29765;
wire v_29766;
wire v_29767;
wire v_29768;
wire v_29769;
wire v_29770;
wire v_29771;
wire v_29772;
wire v_29773;
wire v_29774;
wire v_29775;
wire v_29776;
wire v_29777;
wire v_29778;
wire v_29779;
wire v_29780;
wire v_29781;
wire v_29782;
wire v_29783;
wire v_29784;
wire v_29785;
wire v_29786;
wire v_29787;
wire v_29788;
wire v_29789;
wire v_29790;
wire v_29791;
wire v_29792;
wire v_29793;
wire v_29794;
wire v_29795;
wire v_29796;
wire v_29797;
wire v_29798;
wire v_29799;
wire v_29800;
wire v_29801;
wire v_29802;
wire v_29803;
wire v_29804;
wire v_29805;
wire v_29806;
wire v_29807;
wire v_29808;
wire v_29809;
wire v_29810;
wire v_29811;
wire v_29812;
wire v_29813;
wire v_29814;
wire v_29815;
wire v_29816;
wire v_29817;
wire v_29818;
wire v_29819;
wire v_29820;
wire v_29821;
wire v_29822;
wire v_29823;
wire v_29824;
wire v_29825;
wire v_29826;
wire v_29827;
wire v_29828;
wire v_29829;
wire v_29830;
wire v_29831;
wire v_29832;
wire v_29834;
wire v_29835;
wire v_29836;
wire v_29837;
wire v_29838;
wire v_29839;
wire v_29840;
wire v_29841;
wire v_29842;
wire v_29843;
wire v_29844;
wire v_29845;
wire v_29846;
wire v_29847;
wire v_29848;
wire v_29849;
wire v_29850;
wire v_29851;
wire v_29852;
wire v_29853;
wire v_29854;
wire v_29855;
wire v_29856;
wire v_29857;
wire v_29858;
wire v_29859;
wire v_29860;
wire v_29861;
wire v_29862;
wire v_29863;
wire v_29864;
wire v_29865;
wire v_29866;
wire v_29867;
wire v_29868;
wire v_29869;
wire v_29870;
wire v_29871;
wire v_29872;
wire v_29873;
wire v_29874;
wire v_29875;
wire v_29876;
wire v_29877;
wire v_29878;
wire v_29879;
wire v_29880;
wire v_29881;
wire v_29882;
wire v_29883;
wire v_29884;
wire v_29885;
wire v_29886;
wire v_29887;
wire v_29888;
wire v_29889;
wire v_29890;
wire v_29891;
wire v_29892;
wire v_29893;
wire v_29894;
wire v_29895;
wire v_29896;
wire v_29897;
wire v_29898;
wire v_29899;
wire v_29900;
wire v_29901;
wire v_29902;
wire v_29903;
wire v_29904;
wire v_29905;
wire v_29906;
wire v_29907;
wire v_29908;
wire v_29909;
wire v_29910;
wire v_29911;
wire v_29912;
wire v_29913;
wire v_29914;
wire v_29915;
wire v_29916;
wire v_29917;
wire v_29918;
wire v_29919;
wire v_29920;
wire v_29921;
wire v_29922;
wire v_29923;
wire v_29924;
wire v_29925;
wire v_29926;
wire v_29927;
wire v_29928;
wire v_29929;
wire v_29930;
wire v_29931;
wire v_29932;
wire v_29933;
wire v_29934;
wire v_29935;
wire v_29936;
wire v_29937;
wire v_29938;
wire v_29939;
wire v_29940;
wire v_29941;
wire v_29942;
wire v_29943;
wire v_29944;
wire v_29945;
wire v_29946;
wire v_29947;
wire v_29948;
wire v_29949;
wire v_29950;
wire v_29951;
wire v_29952;
wire v_29953;
wire v_29954;
wire v_29955;
wire v_29956;
wire v_29957;
wire v_29958;
wire v_29959;
wire v_29960;
wire v_29961;
wire v_29962;
wire v_29963;
wire v_29964;
wire v_29965;
wire v_29966;
wire v_29967;
wire v_29968;
wire v_29969;
wire v_29970;
wire v_29971;
wire v_29972;
wire v_29973;
wire v_29974;
wire v_29975;
wire v_29976;
wire v_29977;
wire v_29978;
wire v_29979;
wire v_29980;
wire v_29981;
wire v_29982;
wire v_29983;
wire v_29984;
wire v_29985;
wire v_29986;
wire v_29987;
wire v_29988;
wire v_29989;
wire v_29990;
wire v_29991;
wire v_29992;
wire v_29993;
wire v_29994;
wire v_29995;
wire v_29996;
wire v_29997;
wire v_29998;
wire v_29999;
wire v_30000;
wire v_30001;
wire v_30002;
wire v_30003;
wire v_30004;
wire v_30005;
wire v_30006;
wire v_30007;
wire v_30008;
wire v_30009;
wire v_30010;
wire v_30011;
wire v_30012;
wire v_30013;
wire v_30014;
wire v_30015;
wire v_30016;
wire v_30017;
wire v_30018;
wire v_30019;
wire v_30020;
wire v_30021;
wire v_30022;
wire v_30023;
wire v_30024;
wire v_30025;
wire v_30026;
wire v_30027;
wire v_30028;
wire v_30029;
wire v_30030;
wire v_30031;
wire v_30032;
wire v_30033;
wire v_30034;
wire v_30035;
wire v_30036;
wire v_30037;
wire v_30038;
wire v_30039;
wire v_30040;
wire v_30041;
wire v_30042;
wire v_30043;
wire v_30044;
wire v_30045;
wire v_30046;
wire v_30047;
wire v_30048;
wire v_30049;
wire v_30050;
wire v_30051;
wire v_30052;
wire v_30053;
wire v_30054;
wire v_30055;
wire v_30056;
wire v_30057;
wire v_30058;
wire v_30059;
wire v_30060;
wire v_30061;
wire v_30062;
wire v_30063;
wire v_30064;
wire v_30065;
wire v_30066;
wire v_30067;
wire v_30068;
wire v_30069;
wire v_30070;
wire v_30071;
wire v_30072;
wire v_30073;
wire v_30074;
wire v_30075;
wire v_30077;
wire v_30078;
wire v_30079;
wire v_30080;
wire v_30081;
wire v_30082;
wire v_30083;
wire v_30084;
wire v_30085;
wire v_30086;
wire v_30087;
wire v_30088;
wire v_30089;
wire v_30090;
wire v_30091;
wire v_30092;
wire v_30093;
wire v_30094;
wire v_30095;
wire v_30096;
wire v_30097;
wire v_30098;
wire v_30099;
wire v_30100;
wire v_30101;
wire v_30102;
wire v_30103;
wire v_30104;
wire v_30105;
wire v_30106;
wire v_30107;
wire v_30108;
wire v_30109;
wire v_30110;
wire v_30111;
wire v_30112;
wire v_30113;
wire v_30114;
wire v_30115;
wire v_30116;
wire v_30117;
wire v_30118;
wire v_30119;
wire v_30120;
wire v_30121;
wire v_30122;
wire v_30123;
wire v_30124;
wire v_30125;
wire v_30126;
wire v_30127;
wire v_30128;
wire v_30129;
wire v_30130;
wire v_30131;
wire v_30132;
wire v_30133;
wire v_30134;
wire v_30135;
wire v_30136;
wire v_30137;
wire v_30138;
wire v_30139;
wire v_30140;
wire v_30141;
wire v_30142;
wire v_30143;
wire v_30144;
wire v_30145;
wire v_30146;
wire v_30147;
wire v_30148;
wire v_30149;
wire v_30150;
wire v_30151;
wire v_30152;
wire v_30153;
wire v_30154;
wire v_30155;
wire v_30156;
wire v_30157;
wire v_30158;
wire v_30159;
wire v_30160;
wire v_30161;
wire v_30162;
wire v_30163;
wire v_30164;
wire v_30165;
wire v_30166;
wire v_30167;
wire v_30168;
wire v_30169;
wire v_30170;
wire v_30171;
wire v_30172;
wire v_30173;
wire v_30174;
wire v_30175;
wire v_30176;
wire v_30177;
wire v_30178;
wire v_30179;
wire v_30180;
wire v_30181;
wire v_30182;
wire v_30183;
wire v_30184;
wire v_30185;
wire v_30186;
wire v_30187;
wire v_30188;
wire v_30189;
wire v_30190;
wire v_30191;
wire v_30192;
wire v_30193;
wire v_30194;
wire v_30195;
wire v_30196;
wire v_30197;
wire v_30198;
wire v_30199;
wire v_30200;
wire v_30201;
wire v_30202;
wire v_30203;
wire v_30204;
wire v_30205;
wire v_30206;
wire v_30207;
wire v_30208;
wire v_30209;
wire v_30210;
wire v_30211;
wire v_30212;
wire v_30213;
wire v_30214;
wire v_30215;
wire v_30216;
wire v_30217;
wire v_30218;
wire v_30219;
wire v_30220;
wire v_30221;
wire v_30222;
wire v_30223;
wire v_30224;
wire v_30225;
wire v_30226;
wire v_30227;
wire v_30228;
wire v_30229;
wire v_30230;
wire v_30231;
wire v_30232;
wire v_30233;
wire v_30234;
wire v_30235;
wire v_30236;
wire v_30237;
wire v_30238;
wire v_30239;
wire v_30240;
wire v_30241;
wire v_30242;
wire v_30243;
wire v_30244;
wire v_30245;
wire v_30246;
wire v_30247;
wire v_30248;
wire v_30249;
wire v_30250;
wire v_30251;
wire v_30252;
wire v_30253;
wire v_30254;
wire v_30255;
wire v_30256;
wire v_30257;
wire v_30258;
wire v_30259;
wire v_30260;
wire v_30261;
wire v_30262;
wire v_30263;
wire v_30264;
wire v_30265;
wire v_30266;
wire v_30267;
wire v_30268;
wire v_30269;
wire v_30270;
wire v_30271;
wire v_30272;
wire v_30273;
wire v_30274;
wire v_30275;
wire v_30276;
wire v_30277;
wire v_30278;
wire v_30279;
wire v_30280;
wire v_30281;
wire v_30282;
wire v_30283;
wire v_30284;
wire v_30285;
wire v_30286;
wire v_30287;
wire v_30288;
wire v_30289;
wire v_30290;
wire v_30291;
wire v_30292;
wire v_30293;
wire v_30294;
wire v_30295;
wire v_30296;
wire v_30297;
wire v_30298;
wire v_30299;
wire v_30300;
wire v_30301;
wire v_30302;
wire v_30303;
wire v_30304;
wire v_30305;
wire v_30306;
wire v_30307;
wire v_30308;
wire v_30309;
wire v_30310;
wire v_30311;
wire v_30312;
wire v_30313;
wire v_30314;
wire v_30315;
wire v_30316;
wire v_30317;
wire v_30318;
wire v_30320;
wire v_30321;
wire v_30322;
wire v_30323;
wire v_30324;
wire v_30325;
wire v_30326;
wire v_30327;
wire v_30328;
wire v_30329;
wire v_30330;
wire v_30331;
wire v_30332;
wire v_30333;
wire v_30334;
wire v_30335;
wire v_30336;
wire v_30337;
wire v_30338;
wire v_30339;
wire v_30340;
wire v_30341;
wire v_30342;
wire v_30343;
wire v_30344;
wire v_30345;
wire v_30346;
wire v_30347;
wire v_30348;
wire v_30349;
wire v_30350;
wire v_30351;
wire v_30352;
wire v_30353;
wire v_30354;
wire v_30355;
wire v_30356;
wire v_30357;
wire v_30358;
wire v_30359;
wire v_30360;
wire v_30361;
wire v_30362;
wire v_30363;
wire v_30364;
wire v_30365;
wire v_30366;
wire v_30367;
wire v_30368;
wire v_30369;
wire v_30370;
wire v_30371;
wire v_30372;
wire v_30373;
wire v_30374;
wire v_30375;
wire v_30376;
wire v_30377;
wire v_30378;
wire v_30379;
wire v_30380;
wire v_30381;
wire v_30382;
wire v_30383;
wire v_30384;
wire v_30385;
wire v_30386;
wire v_30387;
wire v_30388;
wire v_30389;
wire v_30390;
wire v_30391;
wire v_30392;
wire v_30393;
wire v_30394;
wire v_30395;
wire v_30396;
wire v_30397;
wire v_30398;
wire v_30399;
wire v_30400;
wire v_30401;
wire v_30402;
wire v_30403;
wire v_30404;
wire v_30405;
wire v_30406;
wire v_30407;
wire v_30408;
wire v_30409;
wire v_30410;
wire v_30411;
wire v_30412;
wire v_30413;
wire v_30414;
wire v_30415;
wire v_30416;
wire v_30417;
wire v_30418;
wire v_30419;
wire v_30420;
wire v_30421;
wire v_30422;
wire v_30423;
wire v_30424;
wire v_30425;
wire v_30426;
wire v_30427;
wire v_30428;
wire v_30429;
wire v_30430;
wire v_30431;
wire v_30432;
wire v_30433;
wire v_30434;
wire v_30435;
wire v_30436;
wire v_30437;
wire v_30438;
wire v_30439;
wire v_30440;
wire v_30441;
wire v_30442;
wire v_30443;
wire v_30444;
wire v_30445;
wire v_30446;
wire v_30447;
wire v_30448;
wire v_30449;
wire v_30450;
wire v_30451;
wire v_30452;
wire v_30453;
wire v_30454;
wire v_30455;
wire v_30456;
wire v_30457;
wire v_30458;
wire v_30459;
wire v_30460;
wire v_30461;
wire v_30462;
wire v_30463;
wire v_30464;
wire v_30465;
wire v_30466;
wire v_30467;
wire v_30468;
wire v_30469;
wire v_30470;
wire v_30471;
wire v_30472;
wire v_30473;
wire v_30474;
wire v_30475;
wire v_30476;
wire v_30477;
wire v_30478;
wire v_30479;
wire v_30480;
wire v_30481;
wire v_30482;
wire v_30483;
wire v_30484;
wire v_30485;
wire v_30486;
wire v_30487;
wire v_30488;
wire v_30489;
wire v_30490;
wire v_30491;
wire v_30492;
wire v_30493;
wire v_30494;
wire v_30495;
wire v_30496;
wire v_30497;
wire v_30498;
wire v_30499;
wire v_30500;
wire v_30501;
wire v_30502;
wire v_30503;
wire v_30504;
wire v_30505;
wire v_30506;
wire v_30507;
wire v_30508;
wire v_30509;
wire v_30510;
wire v_30511;
wire v_30512;
wire v_30513;
wire v_30514;
wire v_30515;
wire v_30516;
wire v_30517;
wire v_30518;
wire v_30519;
wire v_30520;
wire v_30521;
wire v_30522;
wire v_30523;
wire v_30524;
wire v_30525;
wire v_30526;
wire v_30527;
wire v_30528;
wire v_30529;
wire v_30530;
wire v_30531;
wire v_30532;
wire v_30533;
wire v_30534;
wire v_30535;
wire v_30536;
wire v_30537;
wire v_30538;
wire v_30539;
wire v_30540;
wire v_30541;
wire v_30542;
wire v_30543;
wire v_30544;
wire v_30545;
wire v_30546;
wire v_30547;
wire v_30548;
wire v_30549;
wire v_30550;
wire v_30551;
wire v_30552;
wire v_30553;
wire v_30554;
wire v_30555;
wire v_30556;
wire v_30557;
wire v_30558;
wire v_30559;
wire v_30560;
wire v_30561;
wire v_30563;
wire v_30564;
wire v_30565;
wire v_30566;
wire v_30567;
wire v_30568;
wire v_30569;
wire v_30570;
wire v_30571;
wire v_30572;
wire v_30573;
wire v_30574;
wire v_30575;
wire v_30576;
wire v_30577;
wire v_30578;
wire v_30579;
wire v_30580;
wire v_30581;
wire v_30582;
wire v_30583;
wire v_30584;
wire v_30585;
wire v_30586;
wire v_30587;
wire v_30588;
wire v_30589;
wire v_30590;
wire v_30591;
wire v_30592;
wire v_30593;
wire v_30594;
wire v_30595;
wire v_30596;
wire v_30597;
wire v_30598;
wire v_30599;
wire v_30600;
wire v_30601;
wire v_30602;
wire v_30603;
wire v_30604;
wire v_30605;
wire v_30606;
wire v_30607;
wire v_30608;
wire v_30609;
wire v_30610;
wire v_30611;
wire v_30612;
wire v_30613;
wire v_30614;
wire v_30615;
wire v_30616;
wire v_30617;
wire v_30618;
wire v_30619;
wire v_30620;
wire v_30621;
wire v_30622;
wire v_30623;
wire v_30624;
wire v_30625;
wire v_30626;
wire v_30627;
wire v_30628;
wire v_30629;
wire v_30630;
wire v_30631;
wire v_30632;
wire v_30633;
wire v_30634;
wire v_30635;
wire v_30636;
wire v_30637;
wire v_30638;
wire v_30639;
wire v_30640;
wire v_30641;
wire v_30642;
wire v_30643;
wire v_30644;
wire v_30645;
wire v_30646;
wire v_30647;
wire v_30648;
wire v_30649;
wire v_30650;
wire v_30651;
wire v_30652;
wire v_30653;
wire v_30654;
wire v_30655;
wire v_30656;
wire v_30657;
wire v_30658;
wire v_30659;
wire v_30660;
wire v_30661;
wire v_30662;
wire v_30663;
wire v_30664;
wire v_30665;
wire v_30666;
wire v_30667;
wire v_30668;
wire v_30669;
wire v_30670;
wire v_30671;
wire v_30672;
wire v_30673;
wire v_30674;
wire v_30675;
wire v_30676;
wire v_30677;
wire v_30678;
wire v_30679;
wire v_30680;
wire v_30681;
wire v_30682;
wire v_30683;
wire v_30684;
wire v_30685;
wire v_30686;
wire v_30687;
wire v_30688;
wire v_30689;
wire v_30690;
wire v_30691;
wire v_30692;
wire v_30693;
wire v_30694;
wire v_30695;
wire v_30696;
wire v_30697;
wire v_30698;
wire v_30699;
wire v_30700;
wire v_30701;
wire v_30702;
wire v_30703;
wire v_30704;
wire v_30705;
wire v_30706;
wire v_30707;
wire v_30708;
wire v_30709;
wire v_30710;
wire v_30711;
wire v_30712;
wire v_30713;
wire v_30714;
wire v_30715;
wire v_30716;
wire v_30717;
wire v_30718;
wire v_30719;
wire v_30720;
wire v_30721;
wire v_30722;
wire v_30723;
wire v_30724;
wire v_30725;
wire v_30726;
wire v_30727;
wire v_30728;
wire v_30729;
wire v_30730;
wire v_30731;
wire v_30732;
wire v_30733;
wire v_30734;
wire v_30735;
wire v_30736;
wire v_30737;
wire v_30738;
wire v_30739;
wire v_30740;
wire v_30741;
wire v_30742;
wire v_30743;
wire v_30744;
wire v_30745;
wire v_30746;
wire v_30747;
wire v_30748;
wire v_30749;
wire v_30750;
wire v_30751;
wire v_30752;
wire v_30753;
wire v_30754;
wire v_30755;
wire v_30756;
wire v_30757;
wire v_30758;
wire v_30759;
wire v_30760;
wire v_30761;
wire v_30762;
wire v_30763;
wire v_30764;
wire v_30765;
wire v_30766;
wire v_30767;
wire v_30768;
wire v_30769;
wire v_30770;
wire v_30771;
wire v_30772;
wire v_30773;
wire v_30774;
wire v_30775;
wire v_30776;
wire v_30777;
wire v_30778;
wire v_30779;
wire v_30780;
wire v_30781;
wire v_30782;
wire v_30783;
wire v_30784;
wire v_30785;
wire v_30786;
wire v_30787;
wire v_30788;
wire v_30789;
wire v_30790;
wire v_30791;
wire v_30792;
wire v_30793;
wire v_30794;
wire v_30795;
wire v_30796;
wire v_30797;
wire v_30798;
wire v_30799;
wire v_30800;
wire v_30801;
wire v_30802;
wire v_30803;
wire v_30804;
wire v_30806;
wire v_30807;
wire v_30808;
wire v_30809;
wire v_30810;
wire v_30811;
wire v_30812;
wire v_30813;
wire v_30814;
wire v_30815;
wire v_30816;
wire v_30817;
wire v_30818;
wire v_30819;
wire v_30820;
wire v_30821;
wire v_30822;
wire v_30823;
wire v_30824;
wire v_30825;
wire v_30826;
wire v_30827;
wire v_30828;
wire v_30829;
wire v_30830;
wire v_30831;
wire v_30832;
wire v_30833;
wire v_30834;
wire v_30835;
wire v_30836;
wire v_30837;
wire v_30838;
wire v_30839;
wire v_30840;
wire v_30841;
wire v_30842;
wire v_30843;
wire v_30844;
wire v_30845;
wire v_30846;
wire v_30847;
wire v_30848;
wire v_30849;
wire v_30850;
wire v_30851;
wire v_30852;
wire v_30853;
wire v_30854;
wire v_30855;
wire v_30856;
wire v_30857;
wire v_30858;
wire v_30859;
wire v_30860;
wire v_30861;
wire v_30862;
wire v_30863;
wire v_30864;
wire v_30865;
wire v_30866;
wire v_30867;
wire v_30868;
wire v_30869;
wire v_30870;
wire v_30871;
wire v_30872;
wire v_30873;
wire v_30874;
wire v_30875;
wire v_30876;
wire v_30877;
wire v_30878;
wire v_30879;
wire v_30880;
wire v_30881;
wire v_30882;
wire v_30883;
wire v_30884;
wire v_30885;
wire v_30886;
wire v_30887;
wire v_30888;
wire v_30889;
wire v_30890;
wire v_30891;
wire v_30892;
wire v_30893;
wire v_30894;
wire v_30895;
wire v_30896;
wire v_30897;
wire v_30898;
wire v_30899;
wire v_30900;
wire v_30901;
wire v_30902;
wire v_30903;
wire v_30904;
wire v_30905;
wire v_30906;
wire v_30907;
wire v_30908;
wire v_30909;
wire v_30910;
wire v_30911;
wire v_30912;
wire v_30913;
wire v_30914;
wire v_30915;
wire v_30916;
wire v_30917;
wire v_30918;
wire v_30919;
wire v_30920;
wire v_30921;
wire v_30922;
wire v_30923;
wire v_30924;
wire v_30925;
wire v_30926;
wire v_30927;
wire v_30928;
wire v_30929;
wire v_30930;
wire v_30931;
wire v_30932;
wire v_30933;
wire v_30934;
wire v_30935;
wire v_30936;
wire v_30937;
wire v_30938;
wire v_30939;
wire v_30940;
wire v_30941;
wire v_30942;
wire v_30943;
wire v_30944;
wire v_30945;
wire v_30946;
wire v_30947;
wire v_30948;
wire v_30949;
wire v_30950;
wire v_30951;
wire v_30952;
wire v_30953;
wire v_30954;
wire v_30955;
wire v_30956;
wire v_30957;
wire v_30958;
wire v_30959;
wire v_30960;
wire v_30961;
wire v_30962;
wire v_30963;
wire v_30964;
wire v_30965;
wire v_30966;
wire v_30967;
wire v_30968;
wire v_30969;
wire v_30970;
wire v_30971;
wire v_30972;
wire v_30973;
wire v_30974;
wire v_30975;
wire v_30976;
wire v_30977;
wire v_30978;
wire v_30979;
wire v_30980;
wire v_30981;
wire v_30982;
wire v_30983;
wire v_30984;
wire v_30985;
wire v_30986;
wire v_30987;
wire v_30988;
wire v_30989;
wire v_30990;
wire v_30991;
wire v_30992;
wire v_30993;
wire v_30994;
wire v_30995;
wire v_30996;
wire v_30997;
wire v_30998;
wire v_30999;
wire v_31000;
wire v_31001;
wire v_31002;
wire v_31003;
wire v_31004;
wire v_31005;
wire v_31006;
wire v_31007;
wire v_31008;
wire v_31009;
wire v_31010;
wire v_31011;
wire v_31012;
wire v_31013;
wire v_31014;
wire v_31015;
wire v_31016;
wire v_31017;
wire v_31018;
wire v_31019;
wire v_31020;
wire v_31021;
wire v_31022;
wire v_31023;
wire v_31024;
wire v_31025;
wire v_31026;
wire v_31027;
wire v_31028;
wire v_31029;
wire v_31030;
wire v_31031;
wire v_31032;
wire v_31033;
wire v_31034;
wire v_31035;
wire v_31036;
wire v_31037;
wire v_31038;
wire v_31039;
wire v_31040;
wire v_31041;
wire v_31042;
wire v_31043;
wire v_31044;
wire v_31045;
wire v_31046;
wire v_31047;
wire v_31049;
wire v_31050;
wire v_31051;
wire v_31052;
wire v_31053;
wire v_31054;
wire v_31055;
wire v_31056;
wire v_31057;
wire v_31058;
wire v_31059;
wire v_31060;
wire v_31061;
wire v_31062;
wire v_31063;
wire v_31064;
wire v_31065;
wire v_31066;
wire v_31067;
wire v_31068;
wire v_31069;
wire v_31070;
wire v_31071;
wire v_31072;
wire v_31073;
wire v_31074;
wire v_31075;
wire v_31076;
wire v_31077;
wire v_31078;
wire v_31079;
wire v_31080;
wire v_31081;
wire v_31082;
wire v_31083;
wire v_31084;
wire v_31085;
wire v_31086;
wire v_31087;
wire v_31088;
wire v_31089;
wire v_31090;
wire v_31091;
wire v_31092;
wire v_31093;
wire v_31094;
wire v_31095;
wire v_31096;
wire v_31097;
wire v_31098;
wire v_31099;
wire v_31100;
wire v_31101;
wire v_31102;
wire v_31103;
wire v_31104;
wire v_31105;
wire v_31106;
wire v_31107;
wire v_31108;
wire v_31109;
wire v_31110;
wire v_31111;
wire v_31112;
wire v_31113;
wire v_31114;
wire v_31115;
wire v_31116;
wire v_31117;
wire v_31118;
wire v_31119;
wire v_31120;
wire v_31121;
wire v_31122;
wire v_31123;
wire v_31124;
wire v_31125;
wire v_31126;
wire v_31127;
wire v_31128;
wire v_31129;
wire v_31130;
wire v_31131;
wire v_31132;
wire v_31133;
wire v_31134;
wire v_31135;
wire v_31136;
wire v_31137;
wire v_31138;
wire v_31139;
wire v_31140;
wire v_31141;
wire v_31142;
wire v_31143;
wire v_31144;
wire v_31145;
wire v_31146;
wire v_31147;
wire v_31148;
wire v_31149;
wire v_31150;
wire v_31151;
wire v_31152;
wire v_31153;
wire v_31154;
wire v_31155;
wire v_31156;
wire v_31157;
wire v_31158;
wire v_31159;
wire v_31160;
wire v_31161;
wire v_31162;
wire v_31163;
wire v_31164;
wire v_31165;
wire v_31166;
wire v_31167;
wire v_31168;
wire v_31169;
wire v_31170;
wire v_31171;
wire v_31172;
wire v_31173;
wire v_31174;
wire v_31175;
wire v_31176;
wire v_31177;
wire v_31178;
wire v_31179;
wire v_31180;
wire v_31181;
wire v_31182;
wire v_31183;
wire v_31184;
wire v_31185;
wire v_31186;
wire v_31187;
wire v_31188;
wire v_31189;
wire v_31190;
wire v_31191;
wire v_31192;
wire v_31193;
wire v_31194;
wire v_31195;
wire v_31196;
wire v_31197;
wire v_31198;
wire v_31199;
wire v_31200;
wire v_31201;
wire v_31202;
wire v_31203;
wire v_31204;
wire v_31205;
wire v_31206;
wire v_31207;
wire v_31208;
wire v_31209;
wire v_31210;
wire v_31211;
wire v_31212;
wire v_31213;
wire v_31214;
wire v_31215;
wire v_31216;
wire v_31217;
wire v_31218;
wire v_31219;
wire v_31220;
wire v_31221;
wire v_31222;
wire v_31223;
wire v_31224;
wire v_31225;
wire v_31226;
wire v_31227;
wire v_31228;
wire v_31229;
wire v_31230;
wire v_31231;
wire v_31232;
wire v_31233;
wire v_31234;
wire v_31235;
wire v_31236;
wire v_31237;
wire v_31238;
wire v_31239;
wire v_31240;
wire v_31241;
wire v_31242;
wire v_31243;
wire v_31244;
wire v_31245;
wire v_31246;
wire v_31247;
wire v_31248;
wire v_31249;
wire v_31250;
wire v_31251;
wire v_31252;
wire v_31253;
wire v_31254;
wire v_31255;
wire v_31256;
wire v_31257;
wire v_31258;
wire v_31259;
wire v_31260;
wire v_31261;
wire v_31262;
wire v_31263;
wire v_31264;
wire v_31265;
wire v_31266;
wire v_31267;
wire v_31268;
wire v_31269;
wire v_31270;
wire v_31271;
wire v_31272;
wire v_31273;
wire v_31274;
wire v_31275;
wire v_31276;
wire v_31277;
wire v_31278;
wire v_31279;
wire v_31280;
wire v_31281;
wire v_31282;
wire v_31283;
wire v_31284;
wire v_31285;
wire v_31286;
wire v_31287;
wire v_31288;
wire v_31289;
wire v_31290;
wire v_31292;
wire v_31293;
wire v_31294;
wire v_31295;
wire v_31296;
wire v_31297;
wire v_31298;
wire v_31299;
wire v_31300;
wire v_31301;
wire v_31302;
wire v_31303;
wire v_31304;
wire v_31305;
wire v_31306;
wire v_31307;
wire v_31308;
wire v_31309;
wire v_31310;
wire v_31311;
wire v_31312;
wire v_31313;
wire v_31314;
wire v_31315;
wire v_31316;
wire v_31317;
wire v_31318;
wire v_31319;
wire v_31320;
wire v_31321;
wire v_31322;
wire v_31323;
wire v_31324;
wire v_31325;
wire v_31326;
wire v_31327;
wire v_31328;
wire v_31329;
wire v_31330;
wire v_31331;
wire v_31332;
wire v_31333;
wire v_31334;
wire v_31335;
wire v_31336;
wire v_31337;
wire v_31338;
wire v_31339;
wire v_31340;
wire v_31341;
wire v_31342;
wire v_31343;
wire v_31344;
wire v_31345;
wire v_31346;
wire v_31347;
wire v_31348;
wire v_31349;
wire v_31350;
wire v_31351;
wire v_31352;
wire v_31353;
wire v_31354;
wire v_31355;
wire v_31356;
wire v_31357;
wire v_31358;
wire v_31359;
wire v_31360;
wire v_31361;
wire v_31362;
wire v_31363;
wire v_31364;
wire v_31365;
wire v_31366;
wire v_31367;
wire v_31368;
wire v_31369;
wire v_31370;
wire v_31371;
wire v_31372;
wire v_31373;
wire v_31374;
wire v_31375;
wire v_31376;
wire v_31377;
wire v_31378;
wire v_31379;
wire v_31380;
wire v_31381;
wire v_31382;
wire v_31383;
wire v_31384;
wire v_31385;
wire v_31386;
wire v_31387;
wire v_31388;
wire v_31389;
wire v_31390;
wire v_31391;
wire v_31392;
wire v_31393;
wire v_31394;
wire v_31395;
wire v_31396;
wire v_31397;
wire v_31398;
wire v_31399;
wire v_31400;
wire v_31401;
wire v_31402;
wire v_31403;
wire v_31404;
wire v_31405;
wire v_31406;
wire v_31407;
wire v_31408;
wire v_31409;
wire v_31410;
wire v_31411;
wire v_31412;
wire v_31413;
wire v_31414;
wire v_31415;
wire v_31416;
wire v_31417;
wire v_31418;
wire v_31419;
wire v_31420;
wire v_31421;
wire v_31422;
wire v_31423;
wire v_31424;
wire v_31425;
wire v_31426;
wire v_31427;
wire v_31428;
wire v_31429;
wire v_31430;
wire v_31431;
wire v_31432;
wire v_31433;
wire v_31434;
wire v_31435;
wire v_31436;
wire v_31437;
wire v_31438;
wire v_31439;
wire v_31440;
wire v_31441;
wire v_31442;
wire v_31443;
wire v_31444;
wire v_31445;
wire v_31446;
wire v_31447;
wire v_31448;
wire v_31449;
wire v_31450;
wire v_31451;
wire v_31452;
wire v_31453;
wire v_31454;
wire v_31455;
wire v_31456;
wire v_31457;
wire v_31458;
wire v_31459;
wire v_31460;
wire v_31461;
wire v_31462;
wire v_31463;
wire v_31464;
wire v_31465;
wire v_31466;
wire v_31467;
wire v_31468;
wire v_31469;
wire v_31470;
wire v_31471;
wire v_31472;
wire v_31473;
wire v_31474;
wire v_31475;
wire v_31476;
wire v_31477;
wire v_31478;
wire v_31479;
wire v_31480;
wire v_31481;
wire v_31482;
wire v_31483;
wire v_31484;
wire v_31485;
wire v_31486;
wire v_31487;
wire v_31488;
wire v_31489;
wire v_31490;
wire v_31491;
wire v_31492;
wire v_31493;
wire v_31494;
wire v_31495;
wire v_31496;
wire v_31497;
wire v_31498;
wire v_31499;
wire v_31500;
wire v_31501;
wire v_31502;
wire v_31503;
wire v_31504;
wire v_31505;
wire v_31506;
wire v_31507;
wire v_31508;
wire v_31509;
wire v_31510;
wire v_31511;
wire v_31512;
wire v_31513;
wire v_31514;
wire v_31515;
wire v_31516;
wire v_31517;
wire v_31518;
wire v_31519;
wire v_31520;
wire v_31521;
wire v_31522;
wire v_31523;
wire v_31524;
wire v_31525;
wire v_31526;
wire v_31527;
wire v_31528;
wire v_31529;
wire v_31530;
wire v_31531;
wire v_31532;
wire v_31533;
wire v_31535;
wire v_31536;
wire v_31537;
wire v_31538;
wire v_31539;
wire v_31540;
wire v_31541;
wire v_31542;
wire v_31543;
wire v_31544;
wire v_31545;
wire v_31546;
wire v_31547;
wire v_31548;
wire v_31549;
wire v_31550;
wire v_31551;
wire v_31552;
wire v_31553;
wire v_31554;
wire v_31555;
wire v_31556;
wire v_31557;
wire v_31558;
wire v_31559;
wire v_31560;
wire v_31561;
wire v_31562;
wire v_31563;
wire v_31564;
wire v_31565;
wire v_31566;
wire v_31567;
wire v_31568;
wire v_31569;
wire v_31570;
wire v_31571;
wire v_31572;
wire v_31573;
wire v_31574;
wire v_31575;
wire v_31576;
wire v_31577;
wire v_31578;
wire v_31579;
wire v_31580;
wire v_31581;
wire v_31582;
wire v_31583;
wire v_31584;
wire v_31585;
wire v_31586;
wire v_31587;
wire v_31588;
wire v_31589;
wire v_31590;
wire v_31591;
wire v_31592;
wire v_31593;
wire v_31594;
wire v_31595;
wire v_31596;
wire v_31597;
wire v_31598;
wire v_31599;
wire v_31600;
wire v_31601;
wire v_31602;
wire v_31603;
wire v_31604;
wire v_31605;
wire v_31606;
wire v_31607;
wire v_31608;
wire v_31609;
wire v_31610;
wire v_31611;
wire v_31612;
wire v_31613;
wire v_31614;
wire v_31615;
wire v_31616;
wire v_31617;
wire v_31618;
wire v_31619;
wire v_31620;
wire v_31621;
wire v_31622;
wire v_31623;
wire v_31624;
wire v_31625;
wire v_31626;
wire v_31627;
wire v_31628;
wire v_31629;
wire v_31630;
wire v_31631;
wire v_31632;
wire v_31633;
wire v_31634;
wire v_31635;
wire v_31636;
wire v_31637;
wire v_31638;
wire v_31639;
wire v_31640;
wire v_31641;
wire v_31642;
wire v_31643;
wire v_31644;
wire v_31645;
wire v_31646;
wire v_31647;
wire v_31648;
wire v_31649;
wire v_31650;
wire v_31651;
wire v_31652;
wire v_31653;
wire v_31654;
wire v_31655;
wire v_31656;
wire v_31657;
wire v_31658;
wire v_31659;
wire v_31660;
wire v_31661;
wire v_31662;
wire v_31663;
wire v_31664;
wire v_31665;
wire v_31666;
wire v_31667;
wire v_31668;
wire v_31669;
wire v_31670;
wire v_31671;
wire v_31672;
wire v_31673;
wire v_31674;
wire v_31675;
wire v_31676;
wire v_31677;
wire v_31678;
wire v_31679;
wire v_31680;
wire v_31681;
wire v_31682;
wire v_31683;
wire v_31684;
wire v_31685;
wire v_31686;
wire v_31687;
wire v_31688;
wire v_31689;
wire v_31690;
wire v_31691;
wire v_31692;
wire v_31693;
wire v_31694;
wire v_31695;
wire v_31696;
wire v_31697;
wire v_31698;
wire v_31699;
wire v_31700;
wire v_31701;
wire v_31702;
wire v_31703;
wire v_31704;
wire v_31705;
wire v_31706;
wire v_31707;
wire v_31708;
wire v_31709;
wire v_31710;
wire v_31711;
wire v_31712;
wire v_31713;
wire v_31714;
wire v_31715;
wire v_31716;
wire v_31717;
wire v_31718;
wire v_31719;
wire v_31720;
wire v_31721;
wire v_31722;
wire v_31723;
wire v_31724;
wire v_31725;
wire v_31726;
wire v_31727;
wire v_31728;
wire v_31729;
wire v_31730;
wire v_31731;
wire v_31732;
wire v_31733;
wire v_31734;
wire v_31735;
wire v_31736;
wire v_31737;
wire v_31738;
wire v_31739;
wire v_31740;
wire v_31741;
wire v_31742;
wire v_31743;
wire v_31744;
wire v_31745;
wire v_31746;
wire v_31747;
wire v_31748;
wire v_31749;
wire v_31750;
wire v_31751;
wire v_31752;
wire v_31753;
wire v_31754;
wire v_31755;
wire v_31756;
wire v_31757;
wire v_31758;
wire v_31759;
wire v_31760;
wire v_31761;
wire v_31762;
wire v_31763;
wire v_31764;
wire v_31765;
wire v_31766;
wire v_31767;
wire v_31768;
wire v_31769;
wire v_31770;
wire v_31771;
wire v_31772;
wire v_31773;
wire v_31774;
wire v_31775;
wire v_31776;
wire v_31778;
wire v_31779;
wire v_31780;
wire v_31781;
wire v_31782;
wire v_31783;
wire v_31784;
wire v_31785;
wire v_31786;
wire v_31787;
wire v_31788;
wire v_31789;
wire v_31790;
wire v_31791;
wire v_31792;
wire v_31793;
wire v_31794;
wire v_31795;
wire v_31796;
wire v_31797;
wire v_31798;
wire v_31799;
wire v_31800;
wire v_31801;
wire v_31802;
wire v_31803;
wire v_31804;
wire v_31805;
wire v_31806;
wire v_31807;
wire v_31808;
wire v_31809;
wire v_31810;
wire v_31811;
wire v_31812;
wire v_31813;
wire v_31814;
wire v_31815;
wire v_31816;
wire v_31817;
wire v_31818;
wire v_31819;
wire v_31820;
wire v_31821;
wire v_31822;
wire v_31823;
wire v_31824;
wire v_31825;
wire v_31826;
wire v_31827;
wire v_31828;
wire v_31829;
wire v_31830;
wire v_31831;
wire v_31832;
wire v_31833;
wire v_31834;
wire v_31835;
wire v_31836;
wire v_31837;
wire v_31838;
wire v_31839;
wire v_31840;
wire v_31841;
wire v_31842;
wire v_31843;
wire v_31844;
wire v_31845;
wire v_31846;
wire v_31847;
wire v_31848;
wire v_31849;
wire v_31850;
wire v_31851;
wire v_31852;
wire v_31853;
wire v_31854;
wire v_31855;
wire v_31856;
wire v_31857;
wire v_31858;
wire v_31859;
wire v_31860;
wire v_31861;
wire v_31862;
wire v_31863;
wire v_31864;
wire v_31865;
wire v_31866;
wire v_31867;
wire v_31868;
wire v_31869;
wire v_31870;
wire v_31871;
wire v_31872;
wire v_31873;
wire v_31874;
wire v_31875;
wire v_31876;
wire v_31877;
wire v_31878;
wire v_31879;
wire v_31880;
wire v_31881;
wire v_31882;
wire v_31883;
wire v_31884;
wire v_31885;
wire v_31886;
wire v_31887;
wire v_31888;
wire v_31889;
wire v_31890;
wire v_31891;
wire v_31892;
wire v_31893;
wire v_31894;
wire v_31895;
wire v_31896;
wire v_31897;
wire v_31898;
wire v_31899;
wire v_31900;
wire v_31901;
wire v_31902;
wire v_31903;
wire v_31904;
wire v_31905;
wire v_31906;
wire v_31907;
wire v_31908;
wire v_31909;
wire v_31910;
wire v_31911;
wire v_31912;
wire v_31913;
wire v_31914;
wire v_31915;
wire v_31916;
wire v_31917;
wire v_31918;
wire v_31919;
wire v_31920;
wire v_31921;
wire v_31922;
wire v_31923;
wire v_31924;
wire v_31925;
wire v_31926;
wire v_31927;
wire v_31928;
wire v_31929;
wire v_31930;
wire v_31931;
wire v_31932;
wire v_31933;
wire v_31934;
wire v_31935;
wire v_31936;
wire v_31937;
wire v_31938;
wire v_31939;
wire v_31940;
wire v_31941;
wire v_31942;
wire v_31943;
wire v_31944;
wire v_31945;
wire v_31946;
wire v_31947;
wire v_31948;
wire v_31949;
wire v_31950;
wire v_31951;
wire v_31952;
wire v_31953;
wire v_31954;
wire v_31955;
wire v_31956;
wire v_31957;
wire v_31958;
wire v_31959;
wire v_31960;
wire v_31961;
wire v_31962;
wire v_31963;
wire v_31964;
wire v_31965;
wire v_31966;
wire v_31967;
wire v_31968;
wire v_31969;
wire v_31970;
wire v_31971;
wire v_31972;
wire v_31973;
wire v_31974;
wire v_31975;
wire v_31976;
wire v_31977;
wire v_31978;
wire v_31979;
wire v_31980;
wire v_31981;
wire v_31982;
wire v_31983;
wire v_31984;
wire v_31985;
wire v_31986;
wire v_31987;
wire v_31988;
wire v_31989;
wire v_31990;
wire v_31991;
wire v_31992;
wire v_31993;
wire v_31994;
wire v_31995;
wire v_31996;
wire v_31997;
wire v_31998;
wire v_31999;
wire v_32000;
wire v_32001;
wire v_32002;
wire v_32003;
wire v_32004;
wire v_32005;
wire v_32006;
wire v_32007;
wire v_32008;
wire v_32009;
wire v_32010;
wire v_32011;
wire v_32012;
wire v_32013;
wire v_32014;
wire v_32015;
wire v_32016;
wire v_32017;
wire v_32018;
wire v_32019;
wire v_32021;
wire v_32022;
wire v_32023;
wire v_32024;
wire v_32025;
wire v_32026;
wire v_32027;
wire v_32028;
wire v_32029;
wire v_32030;
wire v_32031;
wire v_32032;
wire v_32033;
wire v_32034;
wire v_32035;
wire v_32036;
wire v_32037;
wire v_32038;
wire v_32039;
wire v_32040;
wire v_32041;
wire v_32042;
wire v_32043;
wire v_32044;
wire v_32045;
wire v_32046;
wire v_32047;
wire v_32048;
wire v_32049;
wire v_32050;
wire v_32051;
wire v_32052;
wire v_32053;
wire v_32054;
wire v_32055;
wire v_32056;
wire v_32057;
wire v_32058;
wire v_32059;
wire v_32060;
wire v_32061;
wire v_32062;
wire v_32063;
wire v_32064;
wire v_32065;
wire v_32066;
wire v_32067;
wire v_32068;
wire v_32069;
wire v_32070;
wire v_32071;
wire v_32072;
wire v_32073;
wire v_32074;
wire v_32075;
wire v_32076;
wire v_32077;
wire v_32078;
wire v_32079;
wire v_32080;
wire v_32081;
wire v_32082;
wire v_32083;
wire v_32084;
wire v_32085;
wire v_32086;
wire v_32087;
wire v_32088;
wire v_32089;
wire v_32090;
wire v_32091;
wire v_32092;
wire v_32093;
wire v_32094;
wire v_32095;
wire v_32096;
wire v_32097;
wire v_32098;
wire v_32099;
wire v_32100;
wire v_32101;
wire v_32102;
wire v_32103;
wire v_32104;
wire v_32105;
wire v_32106;
wire v_32107;
wire v_32108;
wire v_32109;
wire v_32110;
wire v_32111;
wire v_32112;
wire v_32113;
wire v_32114;
wire v_32115;
wire v_32116;
wire v_32117;
wire v_32118;
wire v_32119;
wire v_32120;
wire v_32121;
wire v_32122;
wire v_32123;
wire v_32124;
wire v_32125;
wire v_32126;
wire v_32127;
wire v_32128;
wire v_32129;
wire v_32130;
wire v_32131;
wire v_32132;
wire v_32133;
wire v_32134;
wire v_32135;
wire v_32136;
wire v_32137;
wire v_32138;
wire v_32139;
wire v_32140;
wire v_32141;
wire v_32142;
wire v_32143;
wire v_32144;
wire v_32145;
wire v_32146;
wire v_32147;
wire v_32148;
wire v_32149;
wire v_32150;
wire v_32151;
wire v_32152;
wire v_32153;
wire v_32154;
wire v_32155;
wire v_32156;
wire v_32157;
wire v_32158;
wire v_32159;
wire v_32160;
wire v_32161;
wire v_32162;
wire v_32163;
wire v_32164;
wire v_32165;
wire v_32166;
wire v_32167;
wire v_32168;
wire v_32169;
wire v_32170;
wire v_32171;
wire v_32172;
wire v_32173;
wire v_32174;
wire v_32175;
wire v_32176;
wire v_32177;
wire v_32178;
wire v_32179;
wire v_32180;
wire v_32181;
wire v_32182;
wire v_32183;
wire v_32184;
wire v_32185;
wire v_32186;
wire v_32187;
wire v_32188;
wire v_32189;
wire v_32190;
wire v_32191;
wire v_32192;
wire v_32193;
wire v_32194;
wire v_32195;
wire v_32196;
wire v_32197;
wire v_32198;
wire v_32199;
wire v_32200;
wire v_32201;
wire v_32202;
wire v_32203;
wire v_32204;
wire v_32205;
wire v_32206;
wire v_32207;
wire v_32208;
wire v_32209;
wire v_32210;
wire v_32211;
wire v_32212;
wire v_32213;
wire v_32214;
wire v_32215;
wire v_32216;
wire v_32217;
wire v_32218;
wire v_32219;
wire v_32220;
wire v_32221;
wire v_32222;
wire v_32223;
wire v_32224;
wire v_32225;
wire v_32226;
wire v_32227;
wire v_32228;
wire v_32229;
wire v_32230;
wire v_32231;
wire v_32232;
wire v_32233;
wire v_32234;
wire v_32235;
wire v_32236;
wire v_32237;
wire v_32238;
wire v_32239;
wire v_32240;
wire v_32241;
wire v_32242;
wire v_32243;
wire v_32244;
wire v_32245;
wire v_32246;
wire v_32247;
wire v_32248;
wire v_32249;
wire v_32250;
wire v_32251;
wire v_32252;
wire v_32253;
wire v_32254;
wire v_32255;
wire v_32256;
wire v_32257;
wire v_32258;
wire v_32259;
wire v_32260;
wire v_32261;
wire v_32262;
wire v_32264;
wire v_32265;
wire v_32266;
wire v_32267;
wire v_32268;
wire v_32269;
wire v_32270;
wire v_32271;
wire v_32272;
wire v_32273;
wire v_32274;
wire v_32275;
wire v_32276;
wire v_32277;
wire v_32278;
wire v_32279;
wire v_32280;
wire v_32281;
wire v_32282;
wire v_32283;
wire v_32284;
wire v_32285;
wire v_32286;
wire v_32287;
wire v_32288;
wire v_32289;
wire v_32290;
wire v_32291;
wire v_32292;
wire v_32293;
wire v_32294;
wire v_32295;
wire v_32296;
wire v_32297;
wire v_32298;
wire v_32299;
wire v_32300;
wire v_32301;
wire v_32302;
wire v_32303;
wire v_32304;
wire v_32305;
wire v_32306;
wire v_32307;
wire v_32308;
wire v_32309;
wire v_32310;
wire v_32311;
wire v_32312;
wire v_32313;
wire v_32314;
wire v_32315;
wire v_32316;
wire v_32317;
wire v_32318;
wire v_32319;
wire v_32320;
wire v_32321;
wire v_32322;
wire v_32323;
wire v_32324;
wire v_32325;
wire v_32326;
wire v_32327;
wire v_32328;
wire v_32329;
wire v_32330;
wire v_32331;
wire v_32332;
wire v_32333;
wire v_32334;
wire v_32335;
wire v_32336;
wire v_32337;
wire v_32338;
wire v_32339;
wire v_32340;
wire v_32341;
wire v_32342;
wire v_32343;
wire v_32344;
wire v_32345;
wire v_32346;
wire v_32347;
wire v_32348;
wire v_32349;
wire v_32350;
wire v_32351;
wire v_32352;
wire v_32353;
wire v_32354;
wire v_32355;
wire v_32356;
wire v_32357;
wire v_32358;
wire v_32359;
wire v_32360;
wire v_32361;
wire v_32362;
wire v_32363;
wire v_32364;
wire v_32365;
wire v_32366;
wire v_32367;
wire v_32368;
wire v_32369;
wire v_32370;
wire v_32371;
wire v_32372;
wire v_32373;
wire v_32374;
wire v_32375;
wire v_32376;
wire v_32377;
wire v_32378;
wire v_32379;
wire v_32380;
wire v_32381;
wire v_32382;
wire v_32383;
wire v_32384;
wire v_32385;
wire v_32386;
wire v_32387;
wire v_32388;
wire v_32389;
wire v_32390;
wire v_32391;
wire v_32392;
wire v_32393;
wire v_32394;
wire v_32395;
wire v_32396;
wire v_32397;
wire v_32398;
wire v_32399;
wire v_32400;
wire v_32401;
wire v_32402;
wire v_32403;
wire v_32404;
wire v_32405;
wire v_32406;
wire v_32407;
wire v_32408;
wire v_32409;
wire v_32410;
wire v_32411;
wire v_32412;
wire v_32413;
wire v_32414;
wire v_32415;
wire v_32416;
wire v_32417;
wire v_32418;
wire v_32419;
wire v_32420;
wire v_32421;
wire v_32422;
wire v_32423;
wire v_32424;
wire v_32425;
wire v_32426;
wire v_32427;
wire v_32428;
wire v_32429;
wire v_32430;
wire v_32431;
wire v_32432;
wire v_32433;
wire v_32434;
wire v_32435;
wire v_32436;
wire v_32437;
wire v_32438;
wire v_32439;
wire v_32440;
wire v_32441;
wire v_32442;
wire v_32443;
wire v_32444;
wire v_32445;
wire v_32446;
wire v_32447;
wire v_32448;
wire v_32449;
wire v_32450;
wire v_32451;
wire v_32452;
wire v_32453;
wire v_32454;
wire v_32455;
wire v_32456;
wire v_32457;
wire v_32458;
wire v_32459;
wire v_32460;
wire v_32461;
wire v_32462;
wire v_32463;
wire v_32464;
wire v_32465;
wire v_32466;
wire v_32467;
wire v_32468;
wire v_32469;
wire v_32470;
wire v_32471;
wire v_32472;
wire v_32473;
wire v_32474;
wire v_32475;
wire v_32476;
wire v_32477;
wire v_32478;
wire v_32479;
wire v_32480;
wire v_32481;
wire v_32482;
wire v_32483;
wire v_32484;
wire v_32485;
wire v_32486;
wire v_32487;
wire v_32488;
wire v_32489;
wire v_32490;
wire v_32491;
wire v_32492;
wire v_32493;
wire v_32494;
wire v_32495;
wire v_32496;
wire v_32497;
wire v_32498;
wire v_32499;
wire v_32500;
wire v_32501;
wire v_32502;
wire v_32503;
wire v_32504;
wire v_32505;
wire v_32507;
wire v_32508;
wire v_32509;
wire v_32510;
wire v_32511;
wire v_32512;
wire v_32513;
wire v_32514;
wire v_32515;
wire v_32516;
wire v_32517;
wire v_32518;
wire v_32519;
wire v_32520;
wire v_32521;
wire v_32522;
wire v_32523;
wire v_32524;
wire v_32525;
wire v_32526;
wire v_32527;
wire v_32528;
wire v_32529;
wire v_32530;
wire v_32531;
wire v_32532;
wire v_32533;
wire v_32534;
wire v_32535;
wire v_32536;
wire v_32537;
wire v_32538;
wire v_32539;
wire v_32540;
wire v_32541;
wire v_32542;
wire v_32543;
wire v_32544;
wire v_32545;
wire v_32546;
wire v_32547;
wire v_32548;
wire v_32549;
wire v_32550;
wire v_32551;
wire v_32552;
wire v_32553;
wire v_32554;
wire v_32555;
wire v_32556;
wire v_32557;
wire v_32558;
wire v_32559;
wire v_32560;
wire v_32561;
wire v_32562;
wire v_32563;
wire v_32564;
wire v_32565;
wire v_32566;
wire v_32567;
wire v_32568;
wire v_32569;
wire v_32570;
wire v_32571;
wire v_32572;
wire v_32573;
wire v_32574;
wire v_32575;
wire v_32576;
wire v_32577;
wire v_32578;
wire v_32579;
wire v_32580;
wire v_32581;
wire v_32582;
wire v_32583;
wire v_32584;
wire v_32585;
wire v_32586;
wire v_32587;
wire v_32588;
wire v_32589;
wire v_32590;
wire v_32591;
wire v_32592;
wire v_32593;
wire v_32594;
wire v_32595;
wire v_32596;
wire v_32597;
wire v_32598;
wire v_32599;
wire v_32600;
wire v_32601;
wire v_32602;
wire v_32603;
wire v_32604;
wire v_32605;
wire v_32606;
wire v_32607;
wire v_32608;
wire v_32609;
wire v_32610;
wire v_32611;
wire v_32612;
wire v_32613;
wire v_32614;
wire v_32615;
wire v_32616;
wire v_32617;
wire v_32618;
wire v_32619;
wire v_32620;
wire v_32621;
wire v_32622;
wire v_32623;
wire v_32624;
wire v_32625;
wire v_32626;
wire v_32627;
wire v_32628;
wire v_32629;
wire v_32630;
wire v_32631;
wire v_32632;
wire v_32633;
wire v_32634;
wire v_32635;
wire v_32636;
wire v_32637;
wire v_32638;
wire v_32639;
wire v_32640;
wire v_32641;
wire v_32642;
wire v_32643;
wire v_32644;
wire v_32645;
wire v_32646;
wire v_32647;
wire v_32648;
wire v_32649;
wire v_32650;
wire v_32651;
wire v_32652;
wire v_32653;
wire v_32654;
wire v_32655;
wire v_32656;
wire v_32657;
wire v_32658;
wire v_32659;
wire v_32660;
wire v_32661;
wire v_32662;
wire v_32663;
wire v_32664;
wire v_32665;
wire v_32666;
wire v_32667;
wire v_32668;
wire v_32669;
wire v_32670;
wire v_32671;
wire v_32672;
wire v_32673;
wire v_32674;
wire v_32675;
wire v_32676;
wire v_32677;
wire v_32678;
wire v_32679;
wire v_32680;
wire v_32681;
wire v_32682;
wire v_32683;
wire v_32684;
wire v_32685;
wire v_32686;
wire v_32687;
wire v_32688;
wire v_32689;
wire v_32690;
wire v_32691;
wire v_32692;
wire v_32693;
wire v_32694;
wire v_32695;
wire v_32696;
wire v_32697;
wire v_32698;
wire v_32699;
wire v_32700;
wire v_32701;
wire v_32702;
wire v_32703;
wire v_32704;
wire v_32705;
wire v_32706;
wire v_32707;
wire v_32708;
wire v_32709;
wire v_32710;
wire v_32711;
wire v_32712;
wire v_32713;
wire v_32714;
wire v_32715;
wire v_32716;
wire v_32717;
wire v_32718;
wire v_32719;
wire v_32720;
wire v_32721;
wire v_32722;
wire v_32723;
wire v_32724;
wire v_32725;
wire v_32726;
wire v_32727;
wire v_32728;
wire v_32729;
wire v_32730;
wire v_32731;
wire v_32732;
wire v_32733;
wire v_32734;
wire v_32735;
wire v_32736;
wire v_32737;
wire v_32738;
wire v_32739;
wire v_32740;
wire v_32741;
wire v_32742;
wire v_32743;
wire v_32744;
wire v_32745;
wire v_32746;
wire v_32747;
wire v_32748;
wire v_32750;
wire v_32751;
wire v_32752;
wire v_32753;
wire v_32754;
wire v_32755;
wire v_32756;
wire v_32757;
wire v_32758;
wire v_32759;
wire v_32760;
wire v_32761;
wire v_32762;
wire v_32763;
wire v_32764;
wire v_32765;
wire v_32766;
wire v_32767;
wire v_32768;
wire v_32769;
wire v_32770;
wire v_32771;
wire v_32772;
wire v_32773;
wire v_32774;
wire v_32775;
wire v_32776;
wire v_32777;
wire v_32778;
wire v_32779;
wire v_32780;
wire v_32781;
wire v_32782;
wire v_32783;
wire v_32784;
wire v_32785;
wire v_32786;
wire v_32787;
wire v_32788;
wire v_32789;
wire v_32790;
wire v_32791;
wire v_32792;
wire v_32793;
wire v_32794;
wire v_32795;
wire v_32796;
wire v_32797;
wire v_32798;
wire v_32799;
wire v_32800;
wire v_32801;
wire v_32802;
wire v_32803;
wire v_32804;
wire v_32805;
wire v_32806;
wire v_32807;
wire v_32808;
wire v_32809;
wire v_32810;
wire v_32811;
wire v_32812;
wire v_32813;
wire v_32814;
wire v_32815;
wire v_32816;
wire v_32817;
wire v_32818;
wire v_32819;
wire v_32820;
wire v_32821;
wire v_32822;
wire v_32823;
wire v_32824;
wire v_32825;
wire v_32826;
wire v_32827;
wire v_32828;
wire v_32829;
wire v_32830;
wire v_32831;
wire v_32832;
wire v_32833;
wire v_32834;
wire v_32835;
wire v_32836;
wire v_32837;
wire v_32838;
wire v_32839;
wire v_32840;
wire v_32841;
wire v_32842;
wire v_32843;
wire v_32844;
wire v_32845;
wire v_32846;
wire v_32847;
wire v_32848;
wire v_32849;
wire v_32850;
wire v_32851;
wire v_32852;
wire v_32853;
wire v_32854;
wire v_32855;
wire v_32856;
wire v_32857;
wire v_32858;
wire v_32859;
wire v_32860;
wire v_32861;
wire v_32862;
wire v_32863;
wire v_32864;
wire v_32865;
wire v_32866;
wire v_32867;
wire v_32868;
wire v_32869;
wire v_32870;
wire v_32871;
wire v_32872;
wire v_32873;
wire v_32874;
wire v_32875;
wire v_32876;
wire v_32877;
wire v_32878;
wire v_32879;
wire v_32880;
wire v_32881;
wire v_32882;
wire v_32883;
wire v_32884;
wire v_32885;
wire v_32886;
wire v_32887;
wire v_32888;
wire v_32889;
wire v_32890;
wire v_32891;
wire v_32892;
wire v_32893;
wire v_32894;
wire v_32895;
wire v_32896;
wire v_32897;
wire v_32898;
wire v_32899;
wire v_32900;
wire v_32901;
wire v_32902;
wire v_32903;
wire v_32904;
wire v_32905;
wire v_32906;
wire v_32907;
wire v_32908;
wire v_32909;
wire v_32910;
wire v_32911;
wire v_32912;
wire v_32913;
wire v_32914;
wire v_32915;
wire v_32916;
wire v_32917;
wire v_32918;
wire v_32919;
wire v_32920;
wire v_32921;
wire v_32922;
wire v_32923;
wire v_32924;
wire v_32925;
wire v_32926;
wire v_32927;
wire v_32928;
wire v_32929;
wire v_32930;
wire v_32931;
wire v_32932;
wire v_32933;
wire v_32934;
wire v_32935;
wire v_32936;
wire v_32937;
wire v_32938;
wire v_32939;
wire v_32940;
wire v_32941;
wire v_32942;
wire v_32943;
wire v_32944;
wire v_32945;
wire v_32946;
wire v_32947;
wire v_32948;
wire v_32949;
wire v_32950;
wire v_32951;
wire v_32952;
wire v_32953;
wire v_32954;
wire v_32955;
wire v_32956;
wire v_32957;
wire v_32958;
wire v_32959;
wire v_32960;
wire v_32961;
wire v_32962;
wire v_32963;
wire v_32964;
wire v_32965;
wire v_32966;
wire v_32967;
wire v_32968;
wire v_32969;
wire v_32970;
wire v_32971;
wire v_32972;
wire v_32973;
wire v_32974;
wire v_32975;
wire v_32976;
wire v_32977;
wire v_32978;
wire v_32979;
wire v_32980;
wire v_32981;
wire v_32982;
wire v_32983;
wire v_32984;
wire v_32985;
wire v_32986;
wire v_32987;
wire v_32988;
wire v_32989;
wire v_32990;
wire v_32991;
wire v_32993;
wire v_32994;
wire v_32995;
wire v_32996;
wire v_32997;
wire v_32998;
wire v_32999;
wire v_33000;
wire v_33001;
wire v_33002;
wire v_33003;
wire v_33004;
wire v_33005;
wire v_33006;
wire v_33007;
wire v_33008;
wire v_33009;
wire v_33010;
wire v_33011;
wire v_33012;
wire v_33013;
wire v_33014;
wire v_33015;
wire v_33016;
wire v_33017;
wire v_33018;
wire v_33019;
wire v_33020;
wire v_33021;
wire v_33022;
wire v_33023;
wire v_33024;
wire v_33025;
wire v_33026;
wire v_33027;
wire v_33028;
wire v_33029;
wire v_33030;
wire v_33031;
wire v_33032;
wire v_33033;
wire v_33034;
wire v_33035;
wire v_33036;
wire v_33037;
wire v_33038;
wire v_33039;
wire v_33040;
wire v_33041;
wire v_33042;
wire v_33043;
wire v_33044;
wire v_33045;
wire v_33046;
wire v_33047;
wire v_33048;
wire v_33049;
wire v_33050;
wire v_33051;
wire v_33052;
wire v_33053;
wire v_33054;
wire v_33055;
wire v_33056;
wire v_33057;
wire v_33058;
wire v_33059;
wire v_33060;
wire v_33061;
wire v_33062;
wire v_33063;
wire v_33064;
wire v_33065;
wire v_33066;
wire v_33067;
wire v_33068;
wire v_33069;
wire v_33070;
wire v_33071;
wire v_33072;
wire v_33073;
wire v_33074;
wire v_33075;
wire v_33076;
wire v_33077;
wire v_33078;
wire v_33079;
wire v_33080;
wire v_33081;
wire v_33082;
wire v_33083;
wire v_33084;
wire v_33085;
wire v_33086;
wire v_33087;
wire v_33088;
wire v_33089;
wire v_33090;
wire v_33091;
wire v_33092;
wire v_33093;
wire v_33094;
wire v_33095;
wire v_33096;
wire v_33097;
wire v_33098;
wire v_33099;
wire v_33100;
wire v_33101;
wire v_33102;
wire v_33103;
wire v_33104;
wire v_33105;
wire v_33106;
wire v_33107;
wire v_33108;
wire v_33109;
wire v_33110;
wire v_33111;
wire v_33112;
wire v_33113;
wire v_33114;
wire v_33115;
wire v_33116;
wire v_33117;
wire v_33118;
wire v_33119;
wire v_33120;
wire v_33121;
wire v_33122;
wire v_33123;
wire v_33124;
wire v_33125;
wire v_33126;
wire v_33127;
wire v_33128;
wire v_33129;
wire v_33130;
wire v_33131;
wire v_33132;
wire v_33133;
wire v_33134;
wire v_33135;
wire v_33136;
wire v_33137;
wire v_33138;
wire v_33139;
wire v_33140;
wire v_33141;
wire v_33142;
wire v_33143;
wire v_33144;
wire v_33145;
wire v_33146;
wire v_33147;
wire v_33148;
wire v_33149;
wire v_33150;
wire v_33151;
wire v_33152;
wire v_33153;
wire v_33154;
wire v_33155;
wire v_33156;
wire v_33157;
wire v_33158;
wire v_33159;
wire v_33160;
wire v_33161;
wire v_33162;
wire v_33163;
wire v_33164;
wire v_33165;
wire v_33166;
wire v_33167;
wire v_33168;
wire v_33169;
wire v_33170;
wire v_33171;
wire v_33172;
wire v_33173;
wire v_33174;
wire v_33175;
wire v_33176;
wire v_33177;
wire v_33178;
wire v_33179;
wire v_33180;
wire v_33181;
wire v_33182;
wire v_33183;
wire v_33184;
wire v_33185;
wire v_33186;
wire v_33187;
wire v_33188;
wire v_33189;
wire v_33190;
wire v_33191;
wire v_33192;
wire v_33193;
wire v_33194;
wire v_33195;
wire v_33196;
wire v_33197;
wire v_33198;
wire v_33199;
wire v_33200;
wire v_33201;
wire v_33202;
wire v_33203;
wire v_33204;
wire v_33205;
wire v_33206;
wire v_33207;
wire v_33208;
wire v_33209;
wire v_33210;
wire v_33211;
wire v_33212;
wire v_33213;
wire v_33214;
wire v_33215;
wire v_33216;
wire v_33217;
wire v_33218;
wire v_33219;
wire v_33220;
wire v_33221;
wire v_33222;
wire v_33223;
wire v_33224;
wire v_33225;
wire v_33226;
wire v_33227;
wire v_33228;
wire v_33229;
wire v_33230;
wire v_33231;
wire v_33232;
wire v_33233;
wire v_33234;
wire v_33235;
wire v_33236;
wire v_33237;
wire v_33238;
wire v_33239;
wire v_33240;
wire v_33241;
wire v_33242;
wire v_33243;
wire v_33244;
wire v_33245;
wire v_33246;
wire v_33247;
wire v_33248;
wire v_33249;
wire v_33250;
wire v_33251;
wire v_33252;
wire v_33253;
wire v_33254;
wire v_33255;
wire v_33256;
wire v_33257;
wire v_33258;
wire v_33259;
wire v_33260;
wire v_33261;
wire v_33262;
wire v_33263;
wire v_33264;
wire v_33265;
wire v_33266;
wire v_33267;
wire v_33268;
wire v_33269;
wire v_33270;
wire v_33271;
wire v_33272;
wire v_33273;
wire v_33274;
wire v_33275;
wire v_33276;
wire v_33277;
wire v_33278;
wire v_33279;
wire v_33280;
wire v_33281;
wire v_33282;
wire v_33283;
wire v_33284;
wire v_33285;
wire v_33286;
wire v_33287;
wire v_33288;
wire v_33289;
wire v_33290;
wire v_33291;
wire v_33292;
wire v_33293;
wire v_33294;
wire v_33295;
wire v_33296;
wire v_33297;
wire v_33298;
wire v_33299;
wire v_33300;
wire v_33301;
wire v_33302;
wire v_33303;
wire v_33304;
wire v_33305;
wire v_33306;
wire v_33307;
wire v_33308;
wire v_33309;
wire v_33310;
wire v_33311;
wire v_33312;
wire v_33313;
wire v_33314;
wire v_33315;
wire v_33316;
wire v_33317;
wire v_33318;
wire v_33319;
wire v_33320;
wire v_33321;
wire v_33322;
wire v_33323;
wire v_33324;
wire v_33325;
wire v_33326;
wire v_33327;
wire v_33328;
wire v_33329;
wire v_33330;
wire v_33331;
wire v_33332;
wire v_33333;
wire v_33334;
wire v_33335;
wire v_33336;
wire v_33337;
wire v_33338;
wire v_33339;
wire v_33340;
wire v_33341;
wire v_33342;
wire v_33343;
wire v_33344;
wire v_33345;
wire v_33346;
wire v_33347;
wire v_33348;
wire v_33349;
wire v_33350;
wire v_33351;
wire v_33352;
wire v_33353;
wire v_33354;
wire v_33355;
wire v_33356;
wire v_33357;
wire v_33358;
wire v_33359;
wire v_33360;
wire v_33361;
wire v_33362;
wire v_33363;
wire v_33364;
wire v_33365;
wire v_33366;
wire v_33367;
wire v_33368;
wire v_33369;
wire v_33370;
wire v_33371;
wire v_33372;
wire v_33373;
wire v_33374;
wire v_33375;
wire v_33376;
wire v_33377;
wire v_33378;
wire v_33379;
wire v_33380;
wire v_33381;
wire v_33382;
wire v_33383;
wire v_33385;
wire v_33386;
wire v_33387;
wire v_33388;
wire v_33389;
wire v_33390;
wire v_33391;
wire v_33392;
wire v_33393;
wire v_33394;
wire v_33395;
wire v_33396;
wire v_33397;
wire v_33398;
wire v_33399;
wire v_33400;
wire v_33401;
wire v_33402;
wire v_33403;
wire v_33404;
wire v_33405;
wire v_33406;
wire v_33407;
wire v_33408;
wire v_33409;
wire v_33410;
wire v_33411;
wire v_33412;
wire v_33413;
wire v_33414;
wire v_33415;
wire v_33416;
wire v_33417;
wire v_33418;
wire v_33419;
wire v_33420;
wire v_33421;
wire v_33422;
wire v_33423;
wire v_33424;
wire v_33425;
wire v_33426;
wire v_33427;
wire v_33428;
wire v_33429;
wire v_33430;
wire v_33431;
wire v_33432;
wire v_33433;
wire v_33434;
wire v_33435;
wire v_33436;
wire v_33437;
wire v_33438;
wire v_33439;
wire v_33440;
wire v_33441;
wire v_33442;
wire v_33443;
wire v_33444;
wire v_33445;
wire v_33446;
wire v_33447;
wire v_33448;
wire v_33449;
wire v_33450;
wire v_33451;
wire v_33452;
wire v_33453;
wire v_33454;
wire v_33455;
wire v_33456;
wire v_33457;
wire v_33458;
wire v_33459;
wire v_33460;
wire v_33461;
wire v_33462;
wire v_33463;
wire v_33464;
wire v_33465;
wire v_33466;
wire v_33467;
wire v_33468;
wire v_33469;
wire v_33470;
wire v_33471;
wire v_33472;
wire v_33473;
wire v_33474;
wire v_33475;
wire v_33476;
wire v_33477;
wire v_33479;
wire v_33481;
wire v_33482;
wire v_33483;
wire v_33485;
wire v_33486;
wire v_33487;
wire v_33489;
wire v_33490;
wire v_33491;
wire v_33493;
wire v_33494;
wire v_33496;
wire v_33497;
wire v_33498;
wire v_33500;
wire v_33501;
wire v_33502;
wire v_33504;
wire v_33505;
wire v_33506;
wire v_33508;
wire v_33509;
wire v_33510;
wire v_33512;
wire v_33513;
wire v_33514;
wire v_33516;
wire v_33517;
wire v_33518;
wire v_33520;
wire v_33521;
wire v_33522;
wire v_33524;
wire v_33525;
wire v_33526;
wire v_33528;
wire v_33529;
wire v_33530;
wire v_33532;
wire v_33533;
wire v_33534;
wire v_33536;
wire v_33537;
wire v_33538;
wire v_33540;
wire v_33541;
wire v_33542;
wire v_33544;
wire v_33545;
wire v_33546;
wire v_33547;
wire v_33548;
wire v_33549;
wire v_33550;
wire v_33551;
wire v_33552;
wire v_33553;
wire v_33554;
wire v_33555;
wire v_33556;
wire v_33557;
wire v_33558;
wire v_33559;
wire v_33560;
wire v_33561;
wire v_33562;
wire v_33563;
wire v_33564;
wire v_33565;
wire v_33566;
wire v_33567;
wire v_33568;
wire v_33569;
wire v_33570;
wire v_33571;
wire v_33572;
wire v_33573;
wire v_33574;
wire v_33575;
wire v_33576;
wire v_33577;
wire v_33578;
wire v_33579;
wire v_33580;
wire v_33581;
wire v_33582;
wire v_33583;
wire v_33584;
wire v_33585;
wire v_33586;
wire v_33587;
wire v_33588;
wire v_33589;
wire v_33590;
wire v_33591;
wire v_33592;
wire v_33593;
wire v_33594;
wire v_33595;
wire v_33596;
wire v_33597;
wire v_33598;
wire v_33599;
wire v_33600;
wire v_33601;
wire v_33602;
wire v_33603;
wire v_33604;
wire v_33605;
wire v_33606;
wire v_33607;
wire v_33608;
wire v_33609;
wire v_33610;
wire v_33611;
wire v_33612;
wire v_33613;
wire v_33614;
wire v_33615;
wire v_33616;
wire v_33617;
wire v_33618;
wire v_33619;
wire v_33620;
wire v_33621;
wire v_33622;
wire v_33623;
wire v_33624;
wire v_33625;
wire v_33626;
wire v_33627;
wire v_33628;
wire v_33629;
wire v_33630;
wire v_33631;
wire v_33632;
wire v_33633;
wire v_33634;
wire v_33635;
wire v_33636;
wire v_33637;
wire v_33638;
wire v_33639;
wire v_33640;
wire v_33641;
wire v_33642;
wire v_33643;
wire v_33644;
wire v_33645;
wire v_33646;
wire v_33647;
wire v_33648;
wire v_33649;
wire v_33650;
wire v_33651;
wire v_33652;
wire v_33653;
wire v_33654;
wire v_33655;
wire v_33656;
wire v_33657;
wire v_33658;
wire v_33659;
wire v_33660;
wire v_33661;
wire v_33662;
wire v_33663;
wire v_33664;
wire v_33665;
wire v_33666;
wire v_33667;
wire v_33668;
wire v_33669;
wire v_33670;
wire v_33671;
wire v_33672;
wire v_33673;
wire v_33674;
wire v_33675;
wire v_33676;
wire v_33677;
wire v_33678;
wire v_33679;
wire v_33680;
wire v_33681;
wire v_33682;
wire v_33683;
wire v_33684;
wire v_33685;
wire v_33686;
wire v_33687;
wire v_33688;
wire v_33689;
wire v_33690;
wire v_33691;
wire v_33692;
wire v_33693;
wire v_33694;
wire v_33695;
wire v_33696;
wire v_33697;
wire v_33698;
wire v_33699;
wire v_33700;
wire v_33701;
wire v_33702;
wire v_33703;
wire v_33704;
wire v_33705;
wire v_33706;
wire v_33707;
wire v_33708;
wire v_33709;
wire v_33710;
wire v_33711;
wire v_33712;
wire v_33713;
wire v_33714;
wire v_33715;
wire v_33716;
wire v_33717;
wire v_33718;
wire v_33719;
wire v_33720;
wire v_33721;
wire v_33722;
wire v_33723;
wire v_33724;
wire v_33725;
wire v_33726;
wire v_33727;
wire v_33728;
wire v_33729;
wire v_33730;
wire v_33731;
wire v_33732;
wire v_33733;
wire v_33734;
wire v_33735;
wire v_33736;
wire v_33737;
wire v_33739;
wire v_33740;
wire v_33741;
wire v_33742;
wire v_33743;
wire v_33744;
wire v_33745;
wire v_33746;
wire v_33747;
wire v_33748;
wire v_33749;
wire v_33750;
wire v_33751;
wire v_33752;
wire v_33753;
wire v_33754;
wire v_33755;
wire v_33756;
wire v_33757;
wire v_33758;
wire v_33759;
wire v_33760;
wire v_33761;
wire v_33762;
wire v_33763;
wire v_33764;
wire v_33765;
wire v_33766;
wire v_33767;
wire v_33768;
wire v_33769;
wire v_33770;
wire v_33771;
wire v_33772;
wire v_33773;
wire v_33774;
wire v_33775;
wire v_33776;
wire v_33777;
wire v_33778;
wire v_33779;
wire v_33780;
wire v_33781;
wire v_33782;
wire v_33783;
wire v_33784;
wire v_33785;
wire v_33786;
wire v_33787;
wire v_33788;
wire v_33789;
wire v_33790;
wire v_33791;
wire v_33792;
wire v_33793;
wire v_33794;
wire v_33795;
wire v_33796;
wire v_33797;
wire v_33798;
wire v_33799;
wire v_33800;
wire v_33801;
wire v_33802;
wire v_33803;
wire v_33804;
wire v_33805;
wire v_33806;
wire v_33807;
wire v_33808;
wire v_33809;
wire v_33810;
wire v_33811;
wire v_33812;
wire v_33813;
wire v_33814;
wire v_33815;
wire v_33816;
wire v_33817;
wire v_33818;
wire v_33819;
wire v_33820;
wire v_33821;
wire v_33822;
wire v_33823;
wire v_33824;
wire v_33825;
wire v_33826;
wire v_33827;
wire v_33828;
wire v_33829;
wire v_33830;
wire v_33831;
wire v_33832;
wire v_33833;
wire v_33834;
wire v_33835;
wire v_33836;
wire v_33837;
wire v_33838;
wire v_33839;
wire v_33840;
wire v_33841;
wire v_33842;
wire v_33843;
wire v_33844;
wire v_33845;
wire v_33846;
wire v_33847;
wire v_33848;
wire v_33849;
wire v_33850;
wire v_33851;
wire v_33852;
wire v_33853;
wire v_33854;
wire v_33855;
wire v_33856;
wire v_33857;
wire v_33858;
wire v_33859;
wire v_33860;
wire v_33861;
wire v_33862;
wire v_33863;
wire v_33864;
wire v_33865;
wire v_33866;
wire v_33867;
wire v_33868;
wire v_33869;
wire v_33870;
wire v_33871;
wire v_33872;
wire v_33873;
wire v_33874;
wire v_33875;
wire v_33876;
wire v_33877;
wire v_33878;
wire v_33879;
wire v_33880;
wire v_33881;
wire v_33882;
wire v_33883;
wire v_33884;
wire v_33885;
wire v_33886;
wire v_33887;
wire v_33888;
wire v_33889;
wire v_33890;
wire v_33891;
wire v_33892;
wire v_33893;
wire v_33894;
wire v_33895;
wire v_33896;
wire v_33897;
wire v_33898;
wire v_33899;
wire v_33900;
wire v_33901;
wire v_33902;
wire v_33903;
wire v_33904;
wire v_33905;
wire v_33906;
wire v_33907;
wire v_33908;
wire v_33909;
wire v_33910;
wire v_33911;
wire v_33912;
wire v_33913;
wire v_33914;
wire v_33915;
wire v_33916;
wire v_33917;
wire v_33918;
wire v_33919;
wire v_33920;
wire v_33921;
wire v_33922;
wire v_33923;
wire v_33924;
wire v_33925;
wire v_33926;
wire v_33927;
wire v_33928;
wire v_33929;
wire v_33930;
wire v_33931;
wire v_33932;
wire v_33933;
wire v_33934;
wire v_33935;
wire v_33936;
wire v_33937;
wire v_33938;
wire v_33939;
wire v_33940;
wire v_33941;
wire v_33942;
wire v_33943;
wire v_33944;
wire v_33945;
wire v_33946;
wire v_33947;
wire v_33948;
wire v_33949;
wire v_33950;
wire v_33951;
wire v_33952;
wire v_33953;
wire v_33954;
wire v_33955;
wire v_33956;
wire v_33957;
wire v_33958;
wire v_33959;
wire v_33960;
wire v_33961;
wire v_33962;
wire v_33963;
wire v_33964;
wire v_33965;
wire v_33966;
wire v_33967;
wire v_33968;
wire v_33969;
wire v_33970;
wire v_33971;
wire v_33972;
wire v_33973;
wire v_33974;
wire v_33975;
wire v_33976;
wire v_33977;
wire v_33978;
wire v_33979;
wire v_33980;
wire v_33982;
wire v_33983;
wire v_33984;
wire v_33985;
wire v_33986;
wire v_33987;
wire v_33988;
wire v_33989;
wire v_33990;
wire v_33991;
wire v_33992;
wire v_33993;
wire v_33994;
wire v_33995;
wire v_33996;
wire v_33997;
wire v_33998;
wire v_33999;
wire v_34000;
wire v_34001;
wire v_34002;
wire v_34003;
wire v_34004;
wire v_34005;
wire v_34006;
wire v_34007;
wire v_34008;
wire v_34009;
wire v_34010;
wire v_34011;
wire v_34012;
wire v_34013;
wire v_34014;
wire v_34015;
wire v_34016;
wire v_34017;
wire v_34018;
wire v_34019;
wire v_34020;
wire v_34021;
wire v_34022;
wire v_34023;
wire v_34024;
wire v_34025;
wire v_34026;
wire v_34027;
wire v_34028;
wire v_34029;
wire v_34030;
wire v_34031;
wire v_34032;
wire v_34033;
wire v_34034;
wire v_34035;
wire v_34036;
wire v_34037;
wire v_34038;
wire v_34039;
wire v_34040;
wire v_34041;
wire v_34042;
wire v_34043;
wire v_34044;
wire v_34045;
wire v_34046;
wire v_34047;
wire v_34048;
wire v_34049;
wire v_34050;
wire v_34051;
wire v_34052;
wire v_34053;
wire v_34054;
wire v_34055;
wire v_34056;
wire v_34057;
wire v_34058;
wire v_34059;
wire v_34060;
wire v_34061;
wire v_34062;
wire v_34063;
wire v_34064;
wire v_34065;
wire v_34066;
wire v_34067;
wire v_34068;
wire v_34069;
wire v_34070;
wire v_34071;
wire v_34072;
wire v_34073;
wire v_34074;
wire v_34075;
wire v_34076;
wire v_34077;
wire v_34078;
wire v_34079;
wire v_34080;
wire v_34081;
wire v_34082;
wire v_34083;
wire v_34084;
wire v_34085;
wire v_34086;
wire v_34087;
wire v_34088;
wire v_34089;
wire v_34090;
wire v_34091;
wire v_34092;
wire v_34093;
wire v_34094;
wire v_34095;
wire v_34096;
wire v_34097;
wire v_34098;
wire v_34099;
wire v_34100;
wire v_34101;
wire v_34102;
wire v_34103;
wire v_34104;
wire v_34105;
wire v_34106;
wire v_34107;
wire v_34108;
wire v_34109;
wire v_34110;
wire v_34111;
wire v_34112;
wire v_34113;
wire v_34114;
wire v_34115;
wire v_34116;
wire v_34117;
wire v_34118;
wire v_34119;
wire v_34120;
wire v_34121;
wire v_34122;
wire v_34123;
wire v_34124;
wire v_34125;
wire v_34126;
wire v_34127;
wire v_34128;
wire v_34129;
wire v_34130;
wire v_34131;
wire v_34132;
wire v_34133;
wire v_34134;
wire v_34135;
wire v_34136;
wire v_34137;
wire v_34138;
wire v_34139;
wire v_34140;
wire v_34141;
wire v_34142;
wire v_34143;
wire v_34144;
wire v_34145;
wire v_34146;
wire v_34147;
wire v_34148;
wire v_34149;
wire v_34150;
wire v_34151;
wire v_34152;
wire v_34153;
wire v_34154;
wire v_34155;
wire v_34156;
wire v_34157;
wire v_34158;
wire v_34159;
wire v_34160;
wire v_34161;
wire v_34162;
wire v_34163;
wire v_34164;
wire v_34165;
wire v_34166;
wire v_34167;
wire v_34168;
wire v_34169;
wire v_34170;
wire v_34171;
wire v_34172;
wire v_34173;
wire v_34174;
wire v_34175;
wire v_34176;
wire v_34177;
wire v_34178;
wire v_34179;
wire v_34180;
wire v_34181;
wire v_34182;
wire v_34183;
wire v_34184;
wire v_34185;
wire v_34186;
wire v_34187;
wire v_34188;
wire v_34189;
wire v_34190;
wire v_34191;
wire v_34192;
wire v_34193;
wire v_34194;
wire v_34195;
wire v_34196;
wire v_34197;
wire v_34198;
wire v_34199;
wire v_34200;
wire v_34201;
wire v_34202;
wire v_34203;
wire v_34204;
wire v_34205;
wire v_34206;
wire v_34207;
wire v_34208;
wire v_34209;
wire v_34210;
wire v_34211;
wire v_34212;
wire v_34213;
wire v_34214;
wire v_34215;
wire v_34216;
wire v_34217;
wire v_34218;
wire v_34219;
wire v_34220;
wire v_34221;
wire v_34222;
wire v_34223;
wire v_34225;
wire v_34226;
wire v_34227;
wire v_34228;
wire v_34229;
wire v_34230;
wire v_34231;
wire v_34232;
wire v_34233;
wire v_34234;
wire v_34235;
wire v_34236;
wire v_34237;
wire v_34238;
wire v_34239;
wire v_34240;
wire v_34241;
wire v_34242;
wire v_34243;
wire v_34244;
wire v_34245;
wire v_34246;
wire v_34247;
wire v_34248;
wire v_34249;
wire v_34250;
wire v_34251;
wire v_34252;
wire v_34253;
wire v_34254;
wire v_34255;
wire v_34256;
wire v_34257;
wire v_34258;
wire v_34259;
wire v_34260;
wire v_34261;
wire v_34262;
wire v_34263;
wire v_34264;
wire v_34265;
wire v_34266;
wire v_34267;
wire v_34268;
wire v_34269;
wire v_34270;
wire v_34271;
wire v_34272;
wire v_34273;
wire v_34274;
wire v_34275;
wire v_34276;
wire v_34277;
wire v_34278;
wire v_34279;
wire v_34280;
wire v_34281;
wire v_34282;
wire v_34283;
wire v_34284;
wire v_34285;
wire v_34286;
wire v_34287;
wire v_34288;
wire v_34289;
wire v_34290;
wire v_34291;
wire v_34292;
wire v_34293;
wire v_34294;
wire v_34295;
wire v_34296;
wire v_34297;
wire v_34298;
wire v_34299;
wire v_34300;
wire v_34301;
wire v_34302;
wire v_34303;
wire v_34304;
wire v_34305;
wire v_34306;
wire v_34307;
wire v_34308;
wire v_34309;
wire v_34310;
wire v_34311;
wire v_34312;
wire v_34313;
wire v_34314;
wire v_34315;
wire v_34316;
wire v_34317;
wire v_34318;
wire v_34319;
wire v_34320;
wire v_34321;
wire v_34322;
wire v_34323;
wire v_34324;
wire v_34325;
wire v_34326;
wire v_34327;
wire v_34328;
wire v_34329;
wire v_34330;
wire v_34331;
wire v_34332;
wire v_34333;
wire v_34334;
wire v_34335;
wire v_34336;
wire v_34337;
wire v_34338;
wire v_34339;
wire v_34340;
wire v_34341;
wire v_34342;
wire v_34343;
wire v_34344;
wire v_34345;
wire v_34346;
wire v_34347;
wire v_34348;
wire v_34349;
wire v_34350;
wire v_34351;
wire v_34352;
wire v_34353;
wire v_34354;
wire v_34355;
wire v_34356;
wire v_34357;
wire v_34358;
wire v_34359;
wire v_34360;
wire v_34361;
wire v_34362;
wire v_34363;
wire v_34364;
wire v_34365;
wire v_34366;
wire v_34367;
wire v_34368;
wire v_34369;
wire v_34370;
wire v_34371;
wire v_34372;
wire v_34373;
wire v_34374;
wire v_34375;
wire v_34376;
wire v_34377;
wire v_34378;
wire v_34379;
wire v_34380;
wire v_34381;
wire v_34382;
wire v_34383;
wire v_34384;
wire v_34385;
wire v_34386;
wire v_34387;
wire v_34388;
wire v_34389;
wire v_34390;
wire v_34391;
wire v_34392;
wire v_34393;
wire v_34394;
wire v_34395;
wire v_34396;
wire v_34397;
wire v_34398;
wire v_34399;
wire v_34400;
wire v_34401;
wire v_34402;
wire v_34403;
wire v_34404;
wire v_34405;
wire v_34406;
wire v_34407;
wire v_34408;
wire v_34409;
wire v_34410;
wire v_34411;
wire v_34412;
wire v_34413;
wire v_34414;
wire v_34415;
wire v_34416;
wire v_34417;
wire v_34418;
wire v_34419;
wire v_34420;
wire v_34421;
wire v_34422;
wire v_34423;
wire v_34424;
wire v_34425;
wire v_34426;
wire v_34427;
wire v_34428;
wire v_34429;
wire v_34430;
wire v_34431;
wire v_34432;
wire v_34433;
wire v_34434;
wire v_34435;
wire v_34436;
wire v_34437;
wire v_34438;
wire v_34439;
wire v_34440;
wire v_34441;
wire v_34442;
wire v_34443;
wire v_34444;
wire v_34445;
wire v_34446;
wire v_34447;
wire v_34448;
wire v_34449;
wire v_34450;
wire v_34451;
wire v_34452;
wire v_34453;
wire v_34454;
wire v_34455;
wire v_34456;
wire v_34457;
wire v_34458;
wire v_34459;
wire v_34460;
wire v_34461;
wire v_34462;
wire v_34463;
wire v_34464;
wire v_34465;
wire v_34466;
wire v_34468;
wire v_34469;
wire v_34470;
wire v_34471;
wire v_34472;
wire v_34473;
wire v_34474;
wire v_34475;
wire v_34476;
wire v_34477;
wire v_34478;
wire v_34479;
wire v_34480;
wire v_34481;
wire v_34482;
wire v_34483;
wire v_34484;
wire v_34485;
wire v_34486;
wire v_34487;
wire v_34488;
wire v_34489;
wire v_34490;
wire v_34491;
wire v_34492;
wire v_34493;
wire v_34494;
wire v_34495;
wire v_34496;
wire v_34497;
wire v_34498;
wire v_34499;
wire v_34500;
wire v_34501;
wire v_34502;
wire v_34503;
wire v_34504;
wire v_34505;
wire v_34506;
wire v_34507;
wire v_34508;
wire v_34509;
wire v_34510;
wire v_34511;
wire v_34512;
wire v_34513;
wire v_34514;
wire v_34515;
wire v_34516;
wire v_34517;
wire v_34518;
wire v_34519;
wire v_34520;
wire v_34521;
wire v_34522;
wire v_34523;
wire v_34524;
wire v_34525;
wire v_34526;
wire v_34527;
wire v_34528;
wire v_34529;
wire v_34530;
wire v_34531;
wire v_34532;
wire v_34533;
wire v_34534;
wire v_34535;
wire v_34536;
wire v_34537;
wire v_34538;
wire v_34539;
wire v_34540;
wire v_34541;
wire v_34542;
wire v_34543;
wire v_34544;
wire v_34545;
wire v_34546;
wire v_34547;
wire v_34548;
wire v_34549;
wire v_34550;
wire v_34551;
wire v_34552;
wire v_34553;
wire v_34554;
wire v_34555;
wire v_34556;
wire v_34557;
wire v_34558;
wire v_34559;
wire v_34560;
wire v_34561;
wire v_34562;
wire v_34563;
wire v_34564;
wire v_34565;
wire v_34566;
wire v_34567;
wire v_34568;
wire v_34569;
wire v_34570;
wire v_34571;
wire v_34572;
wire v_34573;
wire v_34574;
wire v_34575;
wire v_34576;
wire v_34577;
wire v_34578;
wire v_34579;
wire v_34580;
wire v_34581;
wire v_34582;
wire v_34583;
wire v_34584;
wire v_34585;
wire v_34586;
wire v_34587;
wire v_34588;
wire v_34589;
wire v_34590;
wire v_34591;
wire v_34592;
wire v_34593;
wire v_34594;
wire v_34595;
wire v_34596;
wire v_34597;
wire v_34598;
wire v_34599;
wire v_34600;
wire v_34601;
wire v_34602;
wire v_34603;
wire v_34604;
wire v_34605;
wire v_34606;
wire v_34607;
wire v_34608;
wire v_34609;
wire v_34610;
wire v_34611;
wire v_34612;
wire v_34613;
wire v_34614;
wire v_34615;
wire v_34616;
wire v_34617;
wire v_34618;
wire v_34619;
wire v_34620;
wire v_34621;
wire v_34622;
wire v_34623;
wire v_34624;
wire v_34625;
wire v_34626;
wire v_34627;
wire v_34628;
wire v_34629;
wire v_34630;
wire v_34631;
wire v_34632;
wire v_34633;
wire v_34634;
wire v_34635;
wire v_34636;
wire v_34637;
wire v_34638;
wire v_34639;
wire v_34640;
wire v_34641;
wire v_34642;
wire v_34643;
wire v_34644;
wire v_34645;
wire v_34646;
wire v_34647;
wire v_34648;
wire v_34649;
wire v_34650;
wire v_34651;
wire v_34652;
wire v_34653;
wire v_34654;
wire v_34655;
wire v_34656;
wire v_34657;
wire v_34658;
wire v_34659;
wire v_34660;
wire v_34661;
wire v_34662;
wire v_34663;
wire v_34664;
wire v_34665;
wire v_34666;
wire v_34667;
wire v_34668;
wire v_34669;
wire v_34670;
wire v_34671;
wire v_34672;
wire v_34673;
wire v_34674;
wire v_34675;
wire v_34676;
wire v_34677;
wire v_34678;
wire v_34679;
wire v_34680;
wire v_34681;
wire v_34682;
wire v_34683;
wire v_34684;
wire v_34685;
wire v_34686;
wire v_34687;
wire v_34688;
wire v_34689;
wire v_34690;
wire v_34691;
wire v_34692;
wire v_34693;
wire v_34694;
wire v_34695;
wire v_34696;
wire v_34697;
wire v_34698;
wire v_34699;
wire v_34700;
wire v_34701;
wire v_34702;
wire v_34703;
wire v_34704;
wire v_34705;
wire v_34706;
wire v_34707;
wire v_34708;
wire v_34709;
wire v_34711;
wire v_34712;
wire v_34713;
wire v_34714;
wire v_34715;
wire v_34716;
wire v_34717;
wire v_34718;
wire v_34719;
wire v_34720;
wire v_34721;
wire v_34722;
wire v_34723;
wire v_34724;
wire v_34725;
wire v_34726;
wire v_34727;
wire v_34728;
wire v_34729;
wire v_34730;
wire v_34731;
wire v_34732;
wire v_34733;
wire v_34734;
wire v_34735;
wire v_34736;
wire v_34737;
wire v_34738;
wire v_34739;
wire v_34740;
wire v_34741;
wire v_34742;
wire v_34743;
wire v_34744;
wire v_34745;
wire v_34746;
wire v_34747;
wire v_34748;
wire v_34749;
wire v_34750;
wire v_34751;
wire v_34752;
wire v_34753;
wire v_34754;
wire v_34755;
wire v_34756;
wire v_34757;
wire v_34758;
wire v_34759;
wire v_34760;
wire v_34761;
wire v_34762;
wire v_34763;
wire v_34764;
wire v_34765;
wire v_34766;
wire v_34767;
wire v_34768;
wire v_34769;
wire v_34770;
wire v_34771;
wire v_34772;
wire v_34773;
wire v_34774;
wire v_34775;
wire v_34776;
wire v_34777;
wire v_34778;
wire v_34779;
wire v_34780;
wire v_34781;
wire v_34782;
wire v_34783;
wire v_34784;
wire v_34785;
wire v_34786;
wire v_34787;
wire v_34788;
wire v_34789;
wire v_34790;
wire v_34791;
wire v_34792;
wire v_34793;
wire v_34794;
wire v_34795;
wire v_34796;
wire v_34797;
wire v_34798;
wire v_34799;
wire v_34800;
wire v_34801;
wire v_34802;
wire v_34803;
wire v_34804;
wire v_34805;
wire v_34806;
wire v_34807;
wire v_34808;
wire v_34809;
wire v_34810;
wire v_34811;
wire v_34812;
wire v_34813;
wire v_34814;
wire v_34815;
wire v_34816;
wire v_34817;
wire v_34818;
wire v_34819;
wire v_34820;
wire v_34821;
wire v_34822;
wire v_34823;
wire v_34824;
wire v_34825;
wire v_34826;
wire v_34827;
wire v_34828;
wire v_34829;
wire v_34830;
wire v_34831;
wire v_34832;
wire v_34833;
wire v_34834;
wire v_34835;
wire v_34836;
wire v_34837;
wire v_34838;
wire v_34839;
wire v_34840;
wire v_34841;
wire v_34842;
wire v_34843;
wire v_34844;
wire v_34845;
wire v_34846;
wire v_34847;
wire v_34848;
wire v_34849;
wire v_34850;
wire v_34851;
wire v_34852;
wire v_34853;
wire v_34854;
wire v_34855;
wire v_34856;
wire v_34857;
wire v_34858;
wire v_34859;
wire v_34860;
wire v_34861;
wire v_34862;
wire v_34863;
wire v_34864;
wire v_34865;
wire v_34866;
wire v_34867;
wire v_34868;
wire v_34869;
wire v_34870;
wire v_34871;
wire v_34872;
wire v_34873;
wire v_34874;
wire v_34875;
wire v_34876;
wire v_34877;
wire v_34878;
wire v_34879;
wire v_34880;
wire v_34881;
wire v_34882;
wire v_34883;
wire v_34884;
wire v_34885;
wire v_34886;
wire v_34887;
wire v_34888;
wire v_34889;
wire v_34890;
wire v_34891;
wire v_34892;
wire v_34893;
wire v_34894;
wire v_34895;
wire v_34896;
wire v_34897;
wire v_34898;
wire v_34899;
wire v_34900;
wire v_34901;
wire v_34902;
wire v_34903;
wire v_34904;
wire v_34905;
wire v_34906;
wire v_34907;
wire v_34908;
wire v_34909;
wire v_34910;
wire v_34911;
wire v_34912;
wire v_34913;
wire v_34914;
wire v_34915;
wire v_34916;
wire v_34917;
wire v_34918;
wire v_34919;
wire v_34920;
wire v_34921;
wire v_34922;
wire v_34923;
wire v_34924;
wire v_34925;
wire v_34926;
wire v_34927;
wire v_34928;
wire v_34929;
wire v_34930;
wire v_34931;
wire v_34932;
wire v_34933;
wire v_34934;
wire v_34935;
wire v_34936;
wire v_34937;
wire v_34938;
wire v_34939;
wire v_34940;
wire v_34941;
wire v_34942;
wire v_34943;
wire v_34944;
wire v_34945;
wire v_34946;
wire v_34947;
wire v_34948;
wire v_34949;
wire v_34950;
wire v_34951;
wire v_34952;
wire v_34954;
wire v_34955;
wire v_34956;
wire v_34957;
wire v_34958;
wire v_34959;
wire v_34960;
wire v_34961;
wire v_34962;
wire v_34963;
wire v_34964;
wire v_34965;
wire v_34966;
wire v_34967;
wire v_34968;
wire v_34969;
wire v_34970;
wire v_34971;
wire v_34972;
wire v_34973;
wire v_34974;
wire v_34975;
wire v_34976;
wire v_34977;
wire v_34978;
wire v_34979;
wire v_34980;
wire v_34981;
wire v_34982;
wire v_34983;
wire v_34984;
wire v_34985;
wire v_34986;
wire v_34987;
wire v_34988;
wire v_34989;
wire v_34990;
wire v_34991;
wire v_34992;
wire v_34993;
wire v_34994;
wire v_34995;
wire v_34996;
wire v_34997;
wire v_34998;
wire v_34999;
wire v_35000;
wire v_35001;
wire v_35002;
wire v_35003;
wire v_35004;
wire v_35005;
wire v_35006;
wire v_35007;
wire v_35008;
wire v_35009;
wire v_35010;
wire v_35011;
wire v_35012;
wire v_35013;
wire v_35014;
wire v_35015;
wire v_35016;
wire v_35017;
wire v_35018;
wire v_35019;
wire v_35020;
wire v_35021;
wire v_35022;
wire v_35023;
wire v_35024;
wire v_35025;
wire v_35026;
wire v_35027;
wire v_35028;
wire v_35029;
wire v_35030;
wire v_35031;
wire v_35032;
wire v_35033;
wire v_35034;
wire v_35035;
wire v_35036;
wire v_35037;
wire v_35038;
wire v_35039;
wire v_35040;
wire v_35041;
wire v_35042;
wire v_35043;
wire v_35044;
wire v_35045;
wire v_35046;
wire v_35047;
wire v_35048;
wire v_35049;
wire v_35050;
wire v_35051;
wire v_35052;
wire v_35053;
wire v_35054;
wire v_35055;
wire v_35056;
wire v_35057;
wire v_35058;
wire v_35059;
wire v_35060;
wire v_35061;
wire v_35062;
wire v_35063;
wire v_35064;
wire v_35065;
wire v_35066;
wire v_35067;
wire v_35068;
wire v_35069;
wire v_35070;
wire v_35071;
wire v_35072;
wire v_35073;
wire v_35074;
wire v_35075;
wire v_35076;
wire v_35077;
wire v_35078;
wire v_35079;
wire v_35080;
wire v_35081;
wire v_35082;
wire v_35083;
wire v_35084;
wire v_35085;
wire v_35086;
wire v_35087;
wire v_35088;
wire v_35089;
wire v_35090;
wire v_35091;
wire v_35092;
wire v_35093;
wire v_35094;
wire v_35095;
wire v_35096;
wire v_35097;
wire v_35098;
wire v_35099;
wire v_35100;
wire v_35101;
wire v_35102;
wire v_35103;
wire v_35104;
wire v_35105;
wire v_35106;
wire v_35107;
wire v_35108;
wire v_35109;
wire v_35110;
wire v_35111;
wire v_35112;
wire v_35113;
wire v_35114;
wire v_35115;
wire v_35116;
wire v_35117;
wire v_35118;
wire v_35119;
wire v_35120;
wire v_35121;
wire v_35122;
wire v_35123;
wire v_35124;
wire v_35125;
wire v_35126;
wire v_35127;
wire v_35128;
wire v_35129;
wire v_35130;
wire v_35131;
wire v_35132;
wire v_35133;
wire v_35134;
wire v_35135;
wire v_35136;
wire v_35137;
wire v_35138;
wire v_35139;
wire v_35140;
wire v_35141;
wire v_35142;
wire v_35143;
wire v_35144;
wire v_35145;
wire v_35146;
wire v_35147;
wire v_35148;
wire v_35149;
wire v_35150;
wire v_35151;
wire v_35152;
wire v_35153;
wire v_35154;
wire v_35155;
wire v_35156;
wire v_35157;
wire v_35158;
wire v_35159;
wire v_35160;
wire v_35161;
wire v_35162;
wire v_35163;
wire v_35164;
wire v_35165;
wire v_35166;
wire v_35167;
wire v_35168;
wire v_35169;
wire v_35170;
wire v_35171;
wire v_35172;
wire v_35173;
wire v_35174;
wire v_35175;
wire v_35176;
wire v_35177;
wire v_35178;
wire v_35179;
wire v_35180;
wire v_35181;
wire v_35182;
wire v_35183;
wire v_35184;
wire v_35185;
wire v_35186;
wire v_35187;
wire v_35188;
wire v_35189;
wire v_35190;
wire v_35191;
wire v_35192;
wire v_35193;
wire v_35194;
wire v_35195;
wire v_35197;
wire v_35198;
wire v_35199;
wire v_35200;
wire v_35201;
wire v_35202;
wire v_35203;
wire v_35204;
wire v_35205;
wire v_35206;
wire v_35207;
wire v_35208;
wire v_35209;
wire v_35210;
wire v_35211;
wire v_35212;
wire v_35213;
wire v_35214;
wire v_35215;
wire v_35216;
wire v_35217;
wire v_35218;
wire v_35219;
wire v_35220;
wire v_35221;
wire v_35222;
wire v_35223;
wire v_35224;
wire v_35225;
wire v_35226;
wire v_35227;
wire v_35228;
wire v_35229;
wire v_35230;
wire v_35231;
wire v_35232;
wire v_35233;
wire v_35234;
wire v_35235;
wire v_35236;
wire v_35237;
wire v_35238;
wire v_35239;
wire v_35240;
wire v_35241;
wire v_35242;
wire v_35243;
wire v_35244;
wire v_35245;
wire v_35246;
wire v_35247;
wire v_35248;
wire v_35249;
wire v_35250;
wire v_35251;
wire v_35252;
wire v_35253;
wire v_35254;
wire v_35255;
wire v_35256;
wire v_35257;
wire v_35258;
wire v_35259;
wire v_35260;
wire v_35261;
wire v_35262;
wire v_35263;
wire v_35264;
wire v_35265;
wire v_35266;
wire v_35267;
wire v_35268;
wire v_35269;
wire v_35270;
wire v_35271;
wire v_35272;
wire v_35273;
wire v_35274;
wire v_35275;
wire v_35276;
wire v_35277;
wire v_35278;
wire v_35279;
wire v_35280;
wire v_35281;
wire v_35282;
wire v_35283;
wire v_35284;
wire v_35285;
wire v_35286;
wire v_35287;
wire v_35288;
wire v_35289;
wire v_35290;
wire v_35291;
wire v_35292;
wire v_35293;
wire v_35294;
wire v_35295;
wire v_35296;
wire v_35297;
wire v_35298;
wire v_35299;
wire v_35300;
wire v_35301;
wire v_35302;
wire v_35303;
wire v_35304;
wire v_35305;
wire v_35306;
wire v_35307;
wire v_35308;
wire v_35309;
wire v_35310;
wire v_35311;
wire v_35312;
wire v_35313;
wire v_35314;
wire v_35315;
wire v_35316;
wire v_35317;
wire v_35318;
wire v_35319;
wire v_35320;
wire v_35321;
wire v_35322;
wire v_35323;
wire v_35324;
wire v_35325;
wire v_35326;
wire v_35327;
wire v_35328;
wire v_35329;
wire v_35330;
wire v_35331;
wire v_35332;
wire v_35333;
wire v_35334;
wire v_35335;
wire v_35336;
wire v_35337;
wire v_35338;
wire v_35339;
wire v_35340;
wire v_35341;
wire v_35342;
wire v_35343;
wire v_35344;
wire v_35345;
wire v_35346;
wire v_35347;
wire v_35348;
wire v_35349;
wire v_35350;
wire v_35351;
wire v_35352;
wire v_35353;
wire v_35354;
wire v_35355;
wire v_35356;
wire v_35357;
wire v_35358;
wire v_35359;
wire v_35360;
wire v_35361;
wire v_35362;
wire v_35363;
wire v_35364;
wire v_35365;
wire v_35366;
wire v_35367;
wire v_35368;
wire v_35369;
wire v_35370;
wire v_35371;
wire v_35372;
wire v_35373;
wire v_35374;
wire v_35375;
wire v_35376;
wire v_35377;
wire v_35378;
wire v_35379;
wire v_35380;
wire v_35381;
wire v_35382;
wire v_35383;
wire v_35384;
wire v_35385;
wire v_35386;
wire v_35387;
wire v_35388;
wire v_35389;
wire v_35390;
wire v_35391;
wire v_35392;
wire v_35393;
wire v_35394;
wire v_35395;
wire v_35396;
wire v_35397;
wire v_35398;
wire v_35399;
wire v_35400;
wire v_35401;
wire v_35402;
wire v_35403;
wire v_35404;
wire v_35405;
wire v_35406;
wire v_35407;
wire v_35408;
wire v_35409;
wire v_35410;
wire v_35411;
wire v_35412;
wire v_35413;
wire v_35414;
wire v_35415;
wire v_35416;
wire v_35417;
wire v_35418;
wire v_35419;
wire v_35420;
wire v_35421;
wire v_35422;
wire v_35423;
wire v_35424;
wire v_35425;
wire v_35426;
wire v_35427;
wire v_35428;
wire v_35429;
wire v_35430;
wire v_35431;
wire v_35432;
wire v_35433;
wire v_35434;
wire v_35435;
wire v_35436;
wire v_35437;
wire v_35438;
wire v_35440;
wire v_35441;
wire v_35442;
wire v_35443;
wire v_35444;
wire v_35445;
wire v_35446;
wire v_35447;
wire v_35448;
wire v_35449;
wire v_35450;
wire v_35451;
wire v_35452;
wire v_35453;
wire v_35454;
wire v_35455;
wire v_35456;
wire v_35457;
wire v_35458;
wire v_35459;
wire v_35460;
wire v_35461;
wire v_35462;
wire v_35463;
wire v_35464;
wire v_35465;
wire v_35466;
wire v_35467;
wire v_35468;
wire v_35469;
wire v_35470;
wire v_35471;
wire v_35472;
wire v_35473;
wire v_35474;
wire v_35475;
wire v_35476;
wire v_35477;
wire v_35478;
wire v_35479;
wire v_35480;
wire v_35481;
wire v_35482;
wire v_35483;
wire v_35484;
wire v_35485;
wire v_35486;
wire v_35487;
wire v_35488;
wire v_35489;
wire v_35490;
wire v_35491;
wire v_35492;
wire v_35493;
wire v_35494;
wire v_35495;
wire v_35496;
wire v_35497;
wire v_35498;
wire v_35499;
wire v_35500;
wire v_35501;
wire v_35502;
wire v_35503;
wire v_35504;
wire v_35505;
wire v_35506;
wire v_35507;
wire v_35508;
wire v_35509;
wire v_35510;
wire v_35511;
wire v_35512;
wire v_35513;
wire v_35514;
wire v_35515;
wire v_35516;
wire v_35517;
wire v_35518;
wire v_35519;
wire v_35520;
wire v_35521;
wire v_35522;
wire v_35523;
wire v_35524;
wire v_35525;
wire v_35526;
wire v_35527;
wire v_35528;
wire v_35529;
wire v_35530;
wire v_35531;
wire v_35532;
wire v_35533;
wire v_35534;
wire v_35535;
wire v_35536;
wire v_35537;
wire v_35538;
wire v_35539;
wire v_35540;
wire v_35541;
wire v_35542;
wire v_35543;
wire v_35544;
wire v_35545;
wire v_35546;
wire v_35547;
wire v_35548;
wire v_35549;
wire v_35550;
wire v_35551;
wire v_35552;
wire v_35553;
wire v_35554;
wire v_35555;
wire v_35556;
wire v_35557;
wire v_35558;
wire v_35559;
wire v_35560;
wire v_35561;
wire v_35562;
wire v_35563;
wire v_35564;
wire v_35565;
wire v_35566;
wire v_35567;
wire v_35568;
wire v_35569;
wire v_35570;
wire v_35571;
wire v_35572;
wire v_35573;
wire v_35574;
wire v_35575;
wire v_35576;
wire v_35577;
wire v_35578;
wire v_35579;
wire v_35580;
wire v_35581;
wire v_35582;
wire v_35583;
wire v_35584;
wire v_35585;
wire v_35586;
wire v_35587;
wire v_35588;
wire v_35589;
wire v_35590;
wire v_35591;
wire v_35592;
wire v_35593;
wire v_35594;
wire v_35595;
wire v_35596;
wire v_35597;
wire v_35598;
wire v_35599;
wire v_35600;
wire v_35601;
wire v_35602;
wire v_35603;
wire v_35604;
wire v_35605;
wire v_35606;
wire v_35607;
wire v_35608;
wire v_35609;
wire v_35610;
wire v_35611;
wire v_35612;
wire v_35613;
wire v_35614;
wire v_35615;
wire v_35616;
wire v_35617;
wire v_35618;
wire v_35619;
wire v_35620;
wire v_35621;
wire v_35622;
wire v_35623;
wire v_35624;
wire v_35625;
wire v_35626;
wire v_35627;
wire v_35628;
wire v_35629;
wire v_35630;
wire v_35631;
wire v_35632;
wire v_35633;
wire v_35634;
wire v_35635;
wire v_35636;
wire v_35637;
wire v_35638;
wire v_35639;
wire v_35640;
wire v_35641;
wire v_35642;
wire v_35643;
wire v_35644;
wire v_35645;
wire v_35646;
wire v_35647;
wire v_35648;
wire v_35649;
wire v_35650;
wire v_35651;
wire v_35652;
wire v_35653;
wire v_35654;
wire v_35655;
wire v_35656;
wire v_35657;
wire v_35658;
wire v_35659;
wire v_35660;
wire v_35661;
wire v_35662;
wire v_35663;
wire v_35664;
wire v_35665;
wire v_35666;
wire v_35667;
wire v_35668;
wire v_35669;
wire v_35670;
wire v_35671;
wire v_35672;
wire v_35673;
wire v_35674;
wire v_35675;
wire v_35676;
wire v_35677;
wire v_35678;
wire v_35679;
wire v_35680;
wire v_35681;
wire v_35683;
wire v_35684;
wire v_35685;
wire v_35686;
wire v_35687;
wire v_35688;
wire v_35689;
wire v_35690;
wire v_35691;
wire v_35692;
wire v_35693;
wire v_35694;
wire v_35695;
wire v_35696;
wire v_35697;
wire v_35698;
wire v_35699;
wire v_35700;
wire v_35701;
wire v_35702;
wire v_35703;
wire v_35704;
wire v_35705;
wire v_35706;
wire v_35707;
wire v_35708;
wire v_35709;
wire v_35710;
wire v_35711;
wire v_35712;
wire v_35713;
wire v_35714;
wire v_35715;
wire v_35716;
wire v_35717;
wire v_35718;
wire v_35719;
wire v_35720;
wire v_35721;
wire v_35722;
wire v_35723;
wire v_35724;
wire v_35725;
wire v_35726;
wire v_35727;
wire v_35728;
wire v_35729;
wire v_35730;
wire v_35731;
wire v_35732;
wire v_35733;
wire v_35734;
wire v_35735;
wire v_35736;
wire v_35737;
wire v_35738;
wire v_35739;
wire v_35740;
wire v_35741;
wire v_35742;
wire v_35743;
wire v_35744;
wire v_35745;
wire v_35746;
wire v_35747;
wire v_35748;
wire v_35749;
wire v_35750;
wire v_35751;
wire v_35752;
wire v_35753;
wire v_35754;
wire v_35755;
wire v_35756;
wire v_35757;
wire v_35758;
wire v_35759;
wire v_35760;
wire v_35761;
wire v_35762;
wire v_35763;
wire v_35764;
wire v_35765;
wire v_35766;
wire v_35767;
wire v_35768;
wire v_35769;
wire v_35770;
wire v_35771;
wire v_35772;
wire v_35773;
wire v_35774;
wire v_35775;
wire v_35776;
wire v_35777;
wire v_35778;
wire v_35779;
wire v_35780;
wire v_35781;
wire v_35782;
wire v_35783;
wire v_35784;
wire v_35785;
wire v_35786;
wire v_35787;
wire v_35788;
wire v_35789;
wire v_35790;
wire v_35791;
wire v_35792;
wire v_35793;
wire v_35794;
wire v_35795;
wire v_35796;
wire v_35797;
wire v_35798;
wire v_35799;
wire v_35800;
wire v_35801;
wire v_35802;
wire v_35803;
wire v_35804;
wire v_35805;
wire v_35806;
wire v_35807;
wire v_35808;
wire v_35809;
wire v_35810;
wire v_35811;
wire v_35812;
wire v_35813;
wire v_35814;
wire v_35815;
wire v_35816;
wire v_35817;
wire v_35818;
wire v_35819;
wire v_35820;
wire v_35821;
wire v_35822;
wire v_35823;
wire v_35824;
wire v_35825;
wire v_35826;
wire v_35827;
wire v_35828;
wire v_35829;
wire v_35830;
wire v_35831;
wire v_35832;
wire v_35833;
wire v_35834;
wire v_35835;
wire v_35836;
wire v_35837;
wire v_35838;
wire v_35839;
wire v_35840;
wire v_35841;
wire v_35842;
wire v_35843;
wire v_35844;
wire v_35845;
wire v_35846;
wire v_35847;
wire v_35848;
wire v_35849;
wire v_35850;
wire v_35851;
wire v_35852;
wire v_35853;
wire v_35854;
wire v_35855;
wire v_35856;
wire v_35857;
wire v_35858;
wire v_35859;
wire v_35860;
wire v_35861;
wire v_35862;
wire v_35863;
wire v_35864;
wire v_35865;
wire v_35866;
wire v_35867;
wire v_35868;
wire v_35869;
wire v_35870;
wire v_35871;
wire v_35872;
wire v_35873;
wire v_35874;
wire v_35875;
wire v_35876;
wire v_35877;
wire v_35878;
wire v_35879;
wire v_35880;
wire v_35881;
wire v_35882;
wire v_35883;
wire v_35884;
wire v_35885;
wire v_35886;
wire v_35887;
wire v_35888;
wire v_35889;
wire v_35890;
wire v_35891;
wire v_35892;
wire v_35893;
wire v_35894;
wire v_35895;
wire v_35896;
wire v_35897;
wire v_35898;
wire v_35899;
wire v_35900;
wire v_35901;
wire v_35902;
wire v_35903;
wire v_35904;
wire v_35905;
wire v_35906;
wire v_35907;
wire v_35908;
wire v_35909;
wire v_35910;
wire v_35911;
wire v_35912;
wire v_35913;
wire v_35914;
wire v_35915;
wire v_35916;
wire v_35917;
wire v_35918;
wire v_35919;
wire v_35920;
wire v_35921;
wire v_35922;
wire v_35923;
wire v_35924;
wire v_35926;
wire v_35927;
wire v_35928;
wire v_35929;
wire v_35930;
wire v_35931;
wire v_35932;
wire v_35933;
wire v_35934;
wire v_35935;
wire v_35936;
wire v_35937;
wire v_35938;
wire v_35939;
wire v_35940;
wire v_35941;
wire v_35942;
wire v_35943;
wire v_35944;
wire v_35945;
wire v_35946;
wire v_35947;
wire v_35948;
wire v_35949;
wire v_35950;
wire v_35951;
wire v_35952;
wire v_35953;
wire v_35954;
wire v_35955;
wire v_35956;
wire v_35957;
wire v_35958;
wire v_35959;
wire v_35960;
wire v_35961;
wire v_35962;
wire v_35963;
wire v_35964;
wire v_35965;
wire v_35966;
wire v_35967;
wire v_35968;
wire v_35969;
wire v_35970;
wire v_35971;
wire v_35972;
wire v_35973;
wire v_35974;
wire v_35975;
wire v_35976;
wire v_35977;
wire v_35978;
wire v_35979;
wire v_35980;
wire v_35981;
wire v_35982;
wire v_35983;
wire v_35984;
wire v_35985;
wire v_35986;
wire v_35987;
wire v_35988;
wire v_35989;
wire v_35990;
wire v_35991;
wire v_35992;
wire v_35993;
wire v_35994;
wire v_35995;
wire v_35996;
wire v_35997;
wire v_35998;
wire v_35999;
wire v_36000;
wire v_36001;
wire v_36002;
wire v_36003;
wire v_36004;
wire v_36005;
wire v_36006;
wire v_36007;
wire v_36008;
wire v_36009;
wire v_36010;
wire v_36011;
wire v_36012;
wire v_36013;
wire v_36014;
wire v_36015;
wire v_36016;
wire v_36017;
wire v_36018;
wire v_36019;
wire v_36020;
wire v_36021;
wire v_36022;
wire v_36023;
wire v_36024;
wire v_36025;
wire v_36026;
wire v_36027;
wire v_36028;
wire v_36029;
wire v_36030;
wire v_36031;
wire v_36032;
wire v_36033;
wire v_36034;
wire v_36035;
wire v_36036;
wire v_36037;
wire v_36038;
wire v_36039;
wire v_36040;
wire v_36041;
wire v_36042;
wire v_36043;
wire v_36044;
wire v_36045;
wire v_36046;
wire v_36047;
wire v_36048;
wire v_36049;
wire v_36050;
wire v_36051;
wire v_36052;
wire v_36053;
wire v_36054;
wire v_36055;
wire v_36056;
wire v_36057;
wire v_36058;
wire v_36059;
wire v_36060;
wire v_36061;
wire v_36062;
wire v_36063;
wire v_36064;
wire v_36065;
wire v_36066;
wire v_36067;
wire v_36068;
wire v_36069;
wire v_36070;
wire v_36071;
wire v_36072;
wire v_36073;
wire v_36074;
wire v_36075;
wire v_36076;
wire v_36077;
wire v_36078;
wire v_36079;
wire v_36080;
wire v_36081;
wire v_36082;
wire v_36083;
wire v_36084;
wire v_36085;
wire v_36086;
wire v_36087;
wire v_36088;
wire v_36089;
wire v_36090;
wire v_36091;
wire v_36092;
wire v_36093;
wire v_36094;
wire v_36095;
wire v_36096;
wire v_36097;
wire v_36098;
wire v_36099;
wire v_36100;
wire v_36101;
wire v_36102;
wire v_36103;
wire v_36104;
wire v_36105;
wire v_36106;
wire v_36107;
wire v_36108;
wire v_36109;
wire v_36110;
wire v_36111;
wire v_36112;
wire v_36113;
wire v_36114;
wire v_36115;
wire v_36116;
wire v_36117;
wire v_36118;
wire v_36119;
wire v_36120;
wire v_36121;
wire v_36122;
wire v_36123;
wire v_36124;
wire v_36125;
wire v_36126;
wire v_36127;
wire v_36128;
wire v_36129;
wire v_36130;
wire v_36131;
wire v_36132;
wire v_36133;
wire v_36134;
wire v_36135;
wire v_36136;
wire v_36137;
wire v_36138;
wire v_36139;
wire v_36140;
wire v_36141;
wire v_36142;
wire v_36143;
wire v_36144;
wire v_36145;
wire v_36146;
wire v_36147;
wire v_36148;
wire v_36149;
wire v_36150;
wire v_36151;
wire v_36152;
wire v_36153;
wire v_36154;
wire v_36155;
wire v_36156;
wire v_36157;
wire v_36158;
wire v_36159;
wire v_36160;
wire v_36161;
wire v_36162;
wire v_36163;
wire v_36164;
wire v_36165;
wire v_36166;
wire v_36167;
wire v_36169;
wire v_36170;
wire v_36171;
wire v_36172;
wire v_36173;
wire v_36174;
wire v_36175;
wire v_36176;
wire v_36177;
wire v_36178;
wire v_36179;
wire v_36180;
wire v_36181;
wire v_36182;
wire v_36183;
wire v_36184;
wire v_36185;
wire v_36186;
wire v_36187;
wire v_36188;
wire v_36189;
wire v_36190;
wire v_36191;
wire v_36192;
wire v_36193;
wire v_36194;
wire v_36195;
wire v_36196;
wire v_36197;
wire v_36198;
wire v_36199;
wire v_36200;
wire v_36201;
wire v_36202;
wire v_36203;
wire v_36204;
wire v_36205;
wire v_36206;
wire v_36207;
wire v_36208;
wire v_36209;
wire v_36210;
wire v_36211;
wire v_36212;
wire v_36213;
wire v_36214;
wire v_36215;
wire v_36216;
wire v_36217;
wire v_36218;
wire v_36219;
wire v_36220;
wire v_36221;
wire v_36222;
wire v_36223;
wire v_36224;
wire v_36225;
wire v_36226;
wire v_36227;
wire v_36228;
wire v_36229;
wire v_36230;
wire v_36231;
wire v_36232;
wire v_36233;
wire v_36234;
wire v_36235;
wire v_36236;
wire v_36237;
wire v_36238;
wire v_36239;
wire v_36240;
wire v_36241;
wire v_36242;
wire v_36243;
wire v_36244;
wire v_36245;
wire v_36246;
wire v_36247;
wire v_36248;
wire v_36249;
wire v_36250;
wire v_36251;
wire v_36252;
wire v_36253;
wire v_36254;
wire v_36255;
wire v_36256;
wire v_36257;
wire v_36258;
wire v_36259;
wire v_36260;
wire v_36261;
wire v_36262;
wire v_36263;
wire v_36264;
wire v_36265;
wire v_36266;
wire v_36267;
wire v_36268;
wire v_36269;
wire v_36270;
wire v_36271;
wire v_36272;
wire v_36273;
wire v_36274;
wire v_36275;
wire v_36276;
wire v_36277;
wire v_36278;
wire v_36279;
wire v_36280;
wire v_36281;
wire v_36282;
wire v_36283;
wire v_36284;
wire v_36285;
wire v_36286;
wire v_36287;
wire v_36288;
wire v_36289;
wire v_36290;
wire v_36291;
wire v_36292;
wire v_36293;
wire v_36294;
wire v_36295;
wire v_36296;
wire v_36297;
wire v_36298;
wire v_36299;
wire v_36300;
wire v_36301;
wire v_36302;
wire v_36303;
wire v_36304;
wire v_36305;
wire v_36306;
wire v_36307;
wire v_36308;
wire v_36309;
wire v_36310;
wire v_36311;
wire v_36312;
wire v_36313;
wire v_36314;
wire v_36315;
wire v_36316;
wire v_36317;
wire v_36318;
wire v_36319;
wire v_36320;
wire v_36321;
wire v_36322;
wire v_36323;
wire v_36324;
wire v_36325;
wire v_36326;
wire v_36327;
wire v_36328;
wire v_36329;
wire v_36330;
wire v_36331;
wire v_36332;
wire v_36333;
wire v_36334;
wire v_36335;
wire v_36336;
wire v_36337;
wire v_36338;
wire v_36339;
wire v_36340;
wire v_36341;
wire v_36342;
wire v_36343;
wire v_36344;
wire v_36345;
wire v_36346;
wire v_36347;
wire v_36348;
wire v_36349;
wire v_36350;
wire v_36351;
wire v_36352;
wire v_36353;
wire v_36354;
wire v_36355;
wire v_36356;
wire v_36357;
wire v_36358;
wire v_36359;
wire v_36360;
wire v_36361;
wire v_36362;
wire v_36363;
wire v_36364;
wire v_36365;
wire v_36366;
wire v_36367;
wire v_36368;
wire v_36369;
wire v_36370;
wire v_36371;
wire v_36372;
wire v_36373;
wire v_36374;
wire v_36375;
wire v_36376;
wire v_36377;
wire v_36378;
wire v_36379;
wire v_36380;
wire v_36381;
wire v_36382;
wire v_36383;
wire v_36384;
wire v_36385;
wire v_36386;
wire v_36387;
wire v_36388;
wire v_36389;
wire v_36390;
wire v_36391;
wire v_36392;
wire v_36393;
wire v_36394;
wire v_36395;
wire v_36396;
wire v_36397;
wire v_36398;
wire v_36399;
wire v_36400;
wire v_36401;
wire v_36402;
wire v_36403;
wire v_36404;
wire v_36405;
wire v_36406;
wire v_36407;
wire v_36408;
wire v_36409;
wire v_36410;
wire v_36412;
wire v_36413;
wire v_36414;
wire v_36415;
wire v_36416;
wire v_36417;
wire v_36418;
wire v_36419;
wire v_36420;
wire v_36421;
wire v_36422;
wire v_36423;
wire v_36424;
wire v_36425;
wire v_36426;
wire v_36427;
wire v_36428;
wire v_36429;
wire v_36430;
wire v_36431;
wire v_36432;
wire v_36433;
wire v_36434;
wire v_36435;
wire v_36436;
wire v_36437;
wire v_36438;
wire v_36439;
wire v_36440;
wire v_36441;
wire v_36442;
wire v_36443;
wire v_36444;
wire v_36445;
wire v_36446;
wire v_36447;
wire v_36448;
wire v_36449;
wire v_36450;
wire v_36451;
wire v_36452;
wire v_36453;
wire v_36454;
wire v_36455;
wire v_36456;
wire v_36457;
wire v_36458;
wire v_36459;
wire v_36460;
wire v_36461;
wire v_36462;
wire v_36463;
wire v_36464;
wire v_36465;
wire v_36466;
wire v_36467;
wire v_36468;
wire v_36469;
wire v_36470;
wire v_36471;
wire v_36472;
wire v_36473;
wire v_36474;
wire v_36475;
wire v_36476;
wire v_36477;
wire v_36478;
wire v_36479;
wire v_36480;
wire v_36481;
wire v_36482;
wire v_36483;
wire v_36484;
wire v_36485;
wire v_36486;
wire v_36487;
wire v_36488;
wire v_36489;
wire v_36490;
wire v_36491;
wire v_36492;
wire v_36493;
wire v_36494;
wire v_36495;
wire v_36496;
wire v_36497;
wire v_36498;
wire v_36499;
wire v_36500;
wire v_36501;
wire v_36502;
wire v_36503;
wire v_36504;
wire v_36505;
wire v_36506;
wire v_36507;
wire v_36508;
wire v_36509;
wire v_36510;
wire v_36511;
wire v_36512;
wire v_36513;
wire v_36514;
wire v_36515;
wire v_36516;
wire v_36517;
wire v_36518;
wire v_36519;
wire v_36520;
wire v_36521;
wire v_36522;
wire v_36523;
wire v_36524;
wire v_36525;
wire v_36526;
wire v_36527;
wire v_36528;
wire v_36529;
wire v_36530;
wire v_36531;
wire v_36532;
wire v_36533;
wire v_36534;
wire v_36535;
wire v_36536;
wire v_36537;
wire v_36538;
wire v_36539;
wire v_36540;
wire v_36541;
wire v_36542;
wire v_36543;
wire v_36544;
wire v_36545;
wire v_36546;
wire v_36547;
wire v_36548;
wire v_36549;
wire v_36550;
wire v_36551;
wire v_36552;
wire v_36553;
wire v_36554;
wire v_36555;
wire v_36556;
wire v_36557;
wire v_36558;
wire v_36559;
wire v_36560;
wire v_36561;
wire v_36562;
wire v_36563;
wire v_36564;
wire v_36565;
wire v_36566;
wire v_36567;
wire v_36568;
wire v_36569;
wire v_36570;
wire v_36571;
wire v_36572;
wire v_36573;
wire v_36574;
wire v_36575;
wire v_36576;
wire v_36577;
wire v_36578;
wire v_36579;
wire v_36580;
wire v_36581;
wire v_36582;
wire v_36583;
wire v_36584;
wire v_36585;
wire v_36586;
wire v_36587;
wire v_36588;
wire v_36589;
wire v_36590;
wire v_36591;
wire v_36592;
wire v_36593;
wire v_36594;
wire v_36595;
wire v_36596;
wire v_36597;
wire v_36598;
wire v_36599;
wire v_36600;
wire v_36601;
wire v_36602;
wire v_36603;
wire v_36604;
wire v_36605;
wire v_36606;
wire v_36607;
wire v_36608;
wire v_36609;
wire v_36610;
wire v_36611;
wire v_36612;
wire v_36613;
wire v_36614;
wire v_36615;
wire v_36616;
wire v_36617;
wire v_36618;
wire v_36619;
wire v_36620;
wire v_36621;
wire v_36622;
wire v_36623;
wire v_36624;
wire v_36625;
wire v_36626;
wire v_36627;
wire v_36628;
wire v_36629;
wire v_36630;
wire v_36631;
wire v_36632;
wire v_36633;
wire v_36634;
wire v_36635;
wire v_36636;
wire v_36637;
wire v_36638;
wire v_36639;
wire v_36640;
wire v_36641;
wire v_36642;
wire v_36643;
wire v_36644;
wire v_36645;
wire v_36646;
wire v_36647;
wire v_36648;
wire v_36649;
wire v_36650;
wire v_36651;
wire v_36652;
wire v_36653;
wire v_36655;
wire v_36656;
wire v_36657;
wire v_36658;
wire v_36659;
wire v_36660;
wire v_36661;
wire v_36662;
wire v_36663;
wire v_36664;
wire v_36665;
wire v_36666;
wire v_36667;
wire v_36668;
wire v_36669;
wire v_36670;
wire v_36671;
wire v_36672;
wire v_36673;
wire v_36674;
wire v_36675;
wire v_36676;
wire v_36677;
wire v_36678;
wire v_36679;
wire v_36680;
wire v_36681;
wire v_36682;
wire v_36683;
wire v_36684;
wire v_36685;
wire v_36686;
wire v_36687;
wire v_36688;
wire v_36689;
wire v_36690;
wire v_36691;
wire v_36692;
wire v_36693;
wire v_36694;
wire v_36695;
wire v_36696;
wire v_36697;
wire v_36698;
wire v_36699;
wire v_36700;
wire v_36701;
wire v_36702;
wire v_36703;
wire v_36704;
wire v_36705;
wire v_36706;
wire v_36707;
wire v_36708;
wire v_36709;
wire v_36710;
wire v_36711;
wire v_36712;
wire v_36713;
wire v_36714;
wire v_36715;
wire v_36716;
wire v_36717;
wire v_36718;
wire v_36719;
wire v_36720;
wire v_36721;
wire v_36722;
wire v_36723;
wire v_36724;
wire v_36725;
wire v_36726;
wire v_36727;
wire v_36728;
wire v_36729;
wire v_36730;
wire v_36731;
wire v_36732;
wire v_36733;
wire v_36734;
wire v_36735;
wire v_36736;
wire v_36737;
wire v_36738;
wire v_36739;
wire v_36740;
wire v_36741;
wire v_36742;
wire v_36743;
wire v_36744;
wire v_36745;
wire v_36746;
wire v_36747;
wire v_36748;
wire v_36749;
wire v_36750;
wire v_36751;
wire v_36752;
wire v_36753;
wire v_36754;
wire v_36755;
wire v_36756;
wire v_36757;
wire v_36758;
wire v_36759;
wire v_36760;
wire v_36761;
wire v_36762;
wire v_36763;
wire v_36764;
wire v_36765;
wire v_36766;
wire v_36767;
wire v_36768;
wire v_36769;
wire v_36770;
wire v_36771;
wire v_36772;
wire v_36773;
wire v_36774;
wire v_36775;
wire v_36776;
wire v_36777;
wire v_36778;
wire v_36779;
wire v_36780;
wire v_36781;
wire v_36782;
wire v_36783;
wire v_36784;
wire v_36785;
wire v_36786;
wire v_36787;
wire v_36788;
wire v_36789;
wire v_36790;
wire v_36791;
wire v_36792;
wire v_36793;
wire v_36794;
wire v_36795;
wire v_36796;
wire v_36797;
wire v_36798;
wire v_36799;
wire v_36800;
wire v_36801;
wire v_36802;
wire v_36803;
wire v_36804;
wire v_36805;
wire v_36806;
wire v_36807;
wire v_36808;
wire v_36809;
wire v_36810;
wire v_36811;
wire v_36812;
wire v_36813;
wire v_36814;
wire v_36815;
wire v_36816;
wire v_36817;
wire v_36818;
wire v_36819;
wire v_36820;
wire v_36821;
wire v_36822;
wire v_36823;
wire v_36824;
wire v_36825;
wire v_36826;
wire v_36827;
wire v_36828;
wire v_36829;
wire v_36830;
wire v_36831;
wire v_36832;
wire v_36833;
wire v_36834;
wire v_36835;
wire v_36836;
wire v_36837;
wire v_36838;
wire v_36839;
wire v_36840;
wire v_36841;
wire v_36842;
wire v_36843;
wire v_36844;
wire v_36845;
wire v_36846;
wire v_36847;
wire v_36848;
wire v_36849;
wire v_36850;
wire v_36851;
wire v_36852;
wire v_36853;
wire v_36854;
wire v_36855;
wire v_36856;
wire v_36857;
wire v_36858;
wire v_36859;
wire v_36860;
wire v_36861;
wire v_36862;
wire v_36863;
wire v_36864;
wire v_36865;
wire v_36866;
wire v_36867;
wire v_36868;
wire v_36869;
wire v_36870;
wire v_36871;
wire v_36872;
wire v_36873;
wire v_36874;
wire v_36875;
wire v_36876;
wire v_36877;
wire v_36878;
wire v_36879;
wire v_36880;
wire v_36881;
wire v_36882;
wire v_36883;
wire v_36884;
wire v_36885;
wire v_36886;
wire v_36887;
wire v_36888;
wire v_36889;
wire v_36890;
wire v_36891;
wire v_36892;
wire v_36893;
wire v_36894;
wire v_36895;
wire v_36896;
wire v_36898;
wire v_36899;
wire v_36900;
wire v_36901;
wire v_36902;
wire v_36903;
wire v_36904;
wire v_36905;
wire v_36906;
wire v_36907;
wire v_36908;
wire v_36909;
wire v_36910;
wire v_36911;
wire v_36912;
wire v_36913;
wire v_36914;
wire v_36915;
wire v_36916;
wire v_36917;
wire v_36918;
wire v_36919;
wire v_36920;
wire v_36921;
wire v_36922;
wire v_36923;
wire v_36924;
wire v_36925;
wire v_36926;
wire v_36927;
wire v_36928;
wire v_36929;
wire v_36930;
wire v_36931;
wire v_36932;
wire v_36933;
wire v_36934;
wire v_36935;
wire v_36936;
wire v_36937;
wire v_36938;
wire v_36939;
wire v_36940;
wire v_36941;
wire v_36942;
wire v_36943;
wire v_36944;
wire v_36945;
wire v_36946;
wire v_36947;
wire v_36948;
wire v_36949;
wire v_36950;
wire v_36951;
wire v_36952;
wire v_36953;
wire v_36954;
wire v_36955;
wire v_36956;
wire v_36957;
wire v_36958;
wire v_36959;
wire v_36960;
wire v_36961;
wire v_36962;
wire v_36963;
wire v_36964;
wire v_36965;
wire v_36966;
wire v_36967;
wire v_36968;
wire v_36969;
wire v_36970;
wire v_36971;
wire v_36972;
wire v_36973;
wire v_36974;
wire v_36975;
wire v_36976;
wire v_36977;
wire v_36978;
wire v_36979;
wire v_36980;
wire v_36981;
wire v_36982;
wire v_36983;
wire v_36984;
wire v_36985;
wire v_36986;
wire v_36987;
wire v_36988;
wire v_36989;
wire v_36990;
wire v_36991;
wire v_36992;
wire v_36993;
wire v_36994;
wire v_36995;
wire v_36996;
wire v_36997;
wire v_36998;
wire v_36999;
wire v_37000;
wire v_37001;
wire v_37002;
wire v_37003;
wire v_37004;
wire v_37005;
wire v_37006;
wire v_37007;
wire v_37008;
wire v_37009;
wire v_37010;
wire v_37011;
wire v_37012;
wire v_37013;
wire v_37014;
wire v_37015;
wire v_37016;
wire v_37017;
wire v_37018;
wire v_37019;
wire v_37020;
wire v_37021;
wire v_37022;
wire v_37023;
wire v_37024;
wire v_37025;
wire v_37026;
wire v_37027;
wire v_37028;
wire v_37029;
wire v_37030;
wire v_37031;
wire v_37032;
wire v_37033;
wire v_37034;
wire v_37035;
wire v_37036;
wire v_37037;
wire v_37038;
wire v_37039;
wire v_37040;
wire v_37041;
wire v_37042;
wire v_37043;
wire v_37044;
wire v_37045;
wire v_37046;
wire v_37047;
wire v_37048;
wire v_37049;
wire v_37050;
wire v_37051;
wire v_37052;
wire v_37053;
wire v_37054;
wire v_37055;
wire v_37056;
wire v_37057;
wire v_37058;
wire v_37059;
wire v_37060;
wire v_37061;
wire v_37062;
wire v_37063;
wire v_37064;
wire v_37065;
wire v_37066;
wire v_37067;
wire v_37068;
wire v_37069;
wire v_37070;
wire v_37071;
wire v_37072;
wire v_37073;
wire v_37074;
wire v_37075;
wire v_37076;
wire v_37077;
wire v_37078;
wire v_37079;
wire v_37080;
wire v_37081;
wire v_37082;
wire v_37083;
wire v_37084;
wire v_37085;
wire v_37086;
wire v_37087;
wire v_37088;
wire v_37089;
wire v_37090;
wire v_37091;
wire v_37092;
wire v_37093;
wire v_37094;
wire v_37095;
wire v_37096;
wire v_37097;
wire v_37098;
wire v_37099;
wire v_37100;
wire v_37101;
wire v_37102;
wire v_37103;
wire v_37104;
wire v_37105;
wire v_37106;
wire v_37107;
wire v_37108;
wire v_37109;
wire v_37110;
wire v_37111;
wire v_37112;
wire v_37113;
wire v_37114;
wire v_37115;
wire v_37116;
wire v_37117;
wire v_37118;
wire v_37119;
wire v_37120;
wire v_37121;
wire v_37122;
wire v_37123;
wire v_37124;
wire v_37125;
wire v_37126;
wire v_37127;
wire v_37128;
wire v_37129;
wire v_37130;
wire v_37131;
wire v_37132;
wire v_37133;
wire v_37134;
wire v_37135;
wire v_37136;
wire v_37137;
wire v_37138;
wire v_37139;
wire v_37141;
wire v_37142;
wire v_37143;
wire v_37144;
wire v_37145;
wire v_37146;
wire v_37147;
wire v_37148;
wire v_37149;
wire v_37150;
wire v_37151;
wire v_37152;
wire v_37153;
wire v_37154;
wire v_37155;
wire v_37156;
wire v_37157;
wire v_37158;
wire v_37159;
wire v_37160;
wire v_37161;
wire v_37162;
wire v_37163;
wire v_37164;
wire v_37165;
wire v_37166;
wire v_37167;
wire v_37168;
wire v_37169;
wire v_37170;
wire v_37171;
wire v_37172;
wire v_37173;
wire v_37174;
wire v_37175;
wire v_37176;
wire v_37177;
wire v_37178;
wire v_37179;
wire v_37180;
wire v_37181;
wire v_37182;
wire v_37183;
wire v_37184;
wire v_37185;
wire v_37186;
wire v_37187;
wire v_37188;
wire v_37189;
wire v_37190;
wire v_37191;
wire v_37192;
wire v_37193;
wire v_37194;
wire v_37195;
wire v_37196;
wire v_37197;
wire v_37198;
wire v_37199;
wire v_37200;
wire v_37201;
wire v_37202;
wire v_37203;
wire v_37204;
wire v_37205;
wire v_37206;
wire v_37207;
wire v_37208;
wire v_37209;
wire v_37210;
wire v_37211;
wire v_37212;
wire v_37213;
wire v_37214;
wire v_37215;
wire v_37216;
wire v_37217;
wire v_37218;
wire v_37219;
wire v_37220;
wire v_37221;
wire v_37222;
wire v_37223;
wire v_37224;
wire v_37225;
wire v_37226;
wire v_37227;
wire v_37228;
wire v_37229;
wire v_37230;
wire v_37231;
wire v_37232;
wire v_37233;
wire v_37234;
wire v_37235;
wire v_37236;
wire v_37237;
wire v_37238;
wire v_37239;
wire v_37240;
wire v_37241;
wire v_37242;
wire v_37243;
wire v_37244;
wire v_37245;
wire v_37246;
wire v_37247;
wire v_37248;
wire v_37249;
wire v_37250;
wire v_37251;
wire v_37252;
wire v_37253;
wire v_37254;
wire v_37255;
wire v_37256;
wire v_37257;
wire v_37258;
wire v_37259;
wire v_37260;
wire v_37261;
wire v_37262;
wire v_37263;
wire v_37264;
wire v_37265;
wire v_37266;
wire v_37267;
wire v_37268;
wire v_37269;
wire v_37270;
wire v_37271;
wire v_37272;
wire v_37273;
wire v_37274;
wire v_37275;
wire v_37276;
wire v_37277;
wire v_37278;
wire v_37279;
wire v_37280;
wire v_37281;
wire v_37282;
wire v_37283;
wire v_37284;
wire v_37285;
wire v_37286;
wire v_37287;
wire v_37288;
wire v_37289;
wire v_37290;
wire v_37291;
wire v_37292;
wire v_37293;
wire v_37294;
wire v_37295;
wire v_37296;
wire v_37297;
wire v_37298;
wire v_37299;
wire v_37300;
wire v_37301;
wire v_37302;
wire v_37303;
wire v_37304;
wire v_37305;
wire v_37306;
wire v_37307;
wire v_37308;
wire v_37309;
wire v_37310;
wire v_37311;
wire v_37312;
wire v_37313;
wire v_37314;
wire v_37315;
wire v_37316;
wire v_37317;
wire v_37318;
wire v_37319;
wire v_37320;
wire v_37321;
wire v_37322;
wire v_37323;
wire v_37324;
wire v_37325;
wire v_37326;
wire v_37327;
wire v_37328;
wire v_37329;
wire v_37330;
wire v_37331;
wire v_37332;
wire v_37333;
wire v_37334;
wire v_37335;
wire v_37336;
wire v_37337;
wire v_37338;
wire v_37339;
wire v_37340;
wire v_37341;
wire v_37342;
wire v_37343;
wire v_37344;
wire v_37345;
wire v_37346;
wire v_37347;
wire v_37348;
wire v_37349;
wire v_37350;
wire v_37351;
wire v_37352;
wire v_37353;
wire v_37354;
wire v_37355;
wire v_37356;
wire v_37357;
wire v_37358;
wire v_37359;
wire v_37360;
wire v_37361;
wire v_37362;
wire v_37363;
wire v_37364;
wire v_37365;
wire v_37366;
wire v_37367;
wire v_37368;
wire v_37369;
wire v_37370;
wire v_37371;
wire v_37372;
wire v_37373;
wire v_37374;
wire v_37375;
wire v_37376;
wire v_37377;
wire v_37378;
wire v_37379;
wire v_37380;
wire v_37381;
wire v_37382;
wire v_37383;
wire v_37384;
wire v_37385;
wire v_37386;
wire v_37387;
wire v_37388;
wire v_37389;
wire v_37390;
wire v_37391;
wire v_37392;
wire v_37393;
wire v_37394;
wire v_37395;
wire v_37396;
wire v_37397;
wire v_37398;
wire v_37399;
wire v_37400;
wire v_37401;
wire v_37402;
wire v_37403;
wire v_37404;
wire v_37405;
wire v_37406;
wire v_37407;
wire v_37408;
wire v_37409;
wire v_37410;
wire v_37411;
wire v_37412;
wire v_37413;
wire v_37414;
wire v_37415;
wire v_37416;
wire v_37417;
wire v_37418;
wire v_37419;
wire v_37420;
wire v_37421;
wire v_37422;
wire v_37423;
wire v_37424;
wire v_37425;
wire v_37426;
wire v_37427;
wire v_37428;
wire v_37429;
wire v_37430;
wire v_37431;
wire v_37432;
wire v_37433;
wire v_37434;
wire v_37435;
wire v_37436;
wire v_37437;
wire v_37438;
wire v_37439;
wire v_37440;
wire v_37441;
wire v_37442;
wire v_37443;
wire v_37444;
wire v_37445;
wire v_37446;
wire v_37447;
wire v_37448;
wire v_37449;
wire v_37450;
wire v_37451;
wire v_37452;
wire v_37453;
wire v_37454;
wire v_37455;
wire v_37456;
wire v_37457;
wire v_37458;
wire v_37459;
wire v_37460;
wire v_37461;
wire v_37462;
wire v_37463;
wire v_37464;
wire v_37465;
wire v_37466;
wire v_37467;
wire v_37468;
wire v_37469;
wire v_37470;
wire v_37471;
wire v_37472;
wire v_37473;
wire v_37474;
wire v_37475;
wire v_37476;
wire v_37477;
wire v_37478;
wire v_37479;
wire v_37480;
wire v_37481;
wire v_37482;
wire v_37483;
wire v_37484;
wire v_37485;
wire v_37486;
wire v_37487;
wire v_37488;
wire v_37489;
wire v_37490;
wire v_37491;
wire v_37492;
wire v_37493;
wire v_37494;
wire v_37495;
wire v_37496;
wire v_37497;
wire v_37498;
wire v_37499;
wire v_37500;
wire v_37501;
wire v_37502;
wire v_37503;
wire v_37504;
wire v_37505;
wire v_37506;
wire v_37507;
wire v_37508;
wire v_37509;
wire v_37510;
wire v_37511;
wire v_37512;
wire v_37513;
wire v_37514;
wire v_37515;
wire v_37516;
wire v_37517;
wire v_37518;
wire v_37519;
wire v_37520;
wire v_37521;
wire v_37522;
wire v_37523;
wire v_37524;
wire v_37525;
wire v_37526;
wire v_37527;
wire v_37528;
wire v_37529;
wire v_37530;
wire v_37531;
wire v_37533;
wire v_37534;
wire v_37535;
wire v_37536;
wire v_37537;
wire v_37538;
wire v_37539;
wire v_37540;
wire v_37541;
wire v_37542;
wire v_37543;
wire v_37544;
wire v_37545;
wire v_37546;
wire v_37547;
wire v_37548;
wire v_37549;
wire v_37550;
wire v_37551;
wire v_37552;
wire v_37553;
wire v_37554;
wire v_37555;
wire v_37556;
wire v_37557;
wire v_37558;
wire v_37559;
wire v_37560;
wire v_37561;
wire v_37562;
wire v_37563;
wire v_37564;
wire v_37565;
wire v_37566;
wire v_37567;
wire v_37568;
wire v_37569;
wire v_37570;
wire v_37571;
wire v_37572;
wire v_37573;
wire v_37574;
wire v_37575;
wire v_37576;
wire v_37577;
wire v_37578;
wire v_37579;
wire v_37580;
wire v_37581;
wire v_37582;
wire v_37583;
wire v_37584;
wire v_37585;
wire v_37586;
wire v_37587;
wire v_37588;
wire v_37589;
wire v_37590;
wire v_37591;
wire v_37592;
wire v_37593;
wire v_37594;
wire v_37595;
wire v_37596;
wire v_37597;
wire v_37598;
wire v_37599;
wire v_37600;
wire v_37601;
wire v_37602;
wire v_37603;
wire v_37604;
wire v_37605;
wire v_37606;
wire v_37607;
wire v_37608;
wire v_37609;
wire v_37610;
wire v_37611;
wire v_37612;
wire v_37613;
wire v_37614;
wire v_37615;
wire v_37616;
wire v_37617;
wire v_37618;
wire v_37619;
wire v_37620;
wire v_37621;
wire v_37622;
wire v_37623;
wire v_37624;
wire v_37625;
wire v_37627;
wire v_37629;
wire v_37630;
wire v_37631;
wire v_37633;
wire v_37634;
wire v_37635;
wire v_37637;
wire v_37638;
wire v_37639;
wire v_37641;
wire v_37642;
wire v_37644;
wire v_37645;
wire v_37646;
wire v_37648;
wire v_37649;
wire v_37650;
wire v_37652;
wire v_37653;
wire v_37654;
wire v_37656;
wire v_37657;
wire v_37658;
wire v_37660;
wire v_37661;
wire v_37662;
wire v_37664;
wire v_37665;
wire v_37666;
wire v_37668;
wire v_37669;
wire v_37670;
wire v_37672;
wire v_37673;
wire v_37674;
wire v_37676;
wire v_37677;
wire v_37678;
wire v_37680;
wire v_37681;
wire v_37682;
wire v_37684;
wire v_37685;
wire v_37686;
wire v_37688;
wire v_37689;
wire v_37690;
wire v_37692;
wire v_37693;
wire v_37694;
wire v_37695;
wire v_37696;
wire v_37697;
wire v_37698;
wire v_37699;
wire v_37700;
wire v_37701;
wire v_37702;
wire v_37703;
wire v_37704;
wire v_37705;
wire v_37706;
wire v_37707;
wire v_37708;
wire v_37709;
wire v_37710;
wire v_37711;
wire v_37712;
wire v_37713;
wire v_37714;
wire v_37715;
wire v_37716;
wire v_37717;
wire v_37718;
wire v_37719;
wire v_37720;
wire v_37721;
wire v_37722;
wire v_37723;
wire v_37724;
wire v_37725;
wire v_37726;
wire v_37727;
wire v_37728;
wire v_37729;
wire v_37730;
wire v_37731;
wire v_37732;
wire v_37733;
wire v_37734;
wire v_37735;
wire v_37736;
wire v_37737;
wire v_37738;
wire v_37739;
wire v_37740;
wire v_37741;
wire v_37742;
wire v_37743;
wire v_37744;
wire v_37745;
wire v_37746;
wire v_37747;
wire v_37748;
wire v_37749;
wire v_37750;
wire v_37751;
wire v_37752;
wire v_37753;
wire v_37754;
wire v_37755;
wire v_37756;
wire v_37757;
wire v_37758;
wire v_37759;
wire v_37760;
wire v_37761;
wire v_37762;
wire v_37763;
wire v_37764;
wire v_37765;
wire v_37766;
wire v_37767;
wire v_37768;
wire v_37769;
wire v_37770;
wire v_37771;
wire v_37772;
wire v_37773;
wire v_37774;
wire v_37775;
wire v_37776;
wire v_37777;
wire v_37778;
wire v_37779;
wire v_37780;
wire v_37781;
wire v_37782;
wire v_37783;
wire v_37784;
wire v_37785;
wire v_37786;
wire v_37787;
wire v_37788;
wire v_37789;
wire v_37790;
wire v_37791;
wire v_37792;
wire v_37793;
wire v_37794;
wire v_37795;
wire v_37796;
wire v_37797;
wire v_37798;
wire v_37799;
wire v_37800;
wire v_37801;
wire v_37802;
wire v_37803;
wire v_37804;
wire v_37805;
wire v_37806;
wire v_37807;
wire v_37808;
wire v_37809;
wire v_37810;
wire v_37811;
wire v_37812;
wire v_37813;
wire v_37814;
wire v_37815;
wire v_37816;
wire v_37817;
wire v_37818;
wire v_37819;
wire v_37820;
wire v_37821;
wire v_37822;
wire v_37823;
wire v_37824;
wire v_37825;
wire v_37826;
wire v_37827;
wire v_37828;
wire v_37829;
wire v_37830;
wire v_37831;
wire v_37832;
wire v_37833;
wire v_37834;
wire v_37835;
wire v_37836;
wire v_37837;
wire v_37838;
wire v_37839;
wire v_37840;
wire v_37841;
wire v_37842;
wire v_37843;
wire v_37844;
wire v_37845;
wire v_37846;
wire v_37847;
wire v_37848;
wire v_37849;
wire v_37850;
wire v_37851;
wire v_37852;
wire v_37853;
wire v_37854;
wire v_37855;
wire v_37856;
wire v_37857;
wire v_37858;
wire v_37859;
wire v_37860;
wire v_37861;
wire v_37862;
wire v_37863;
wire v_37864;
wire v_37865;
wire v_37866;
wire v_37867;
wire v_37868;
wire v_37869;
wire v_37870;
wire v_37871;
wire v_37872;
wire v_37873;
wire v_37874;
wire v_37875;
wire v_37876;
wire v_37877;
wire v_37878;
wire v_37879;
wire v_37880;
wire v_37881;
wire v_37882;
wire v_37883;
wire v_37884;
wire v_37885;
wire v_37887;
wire v_37888;
wire v_37889;
wire v_37890;
wire v_37891;
wire v_37892;
wire v_37893;
wire v_37894;
wire v_37895;
wire v_37896;
wire v_37897;
wire v_37898;
wire v_37899;
wire v_37900;
wire v_37901;
wire v_37902;
wire v_37903;
wire v_37904;
wire v_37905;
wire v_37906;
wire v_37907;
wire v_37908;
wire v_37909;
wire v_37910;
wire v_37911;
wire v_37912;
wire v_37913;
wire v_37914;
wire v_37915;
wire v_37916;
wire v_37917;
wire v_37918;
wire v_37919;
wire v_37920;
wire v_37921;
wire v_37922;
wire v_37923;
wire v_37924;
wire v_37925;
wire v_37926;
wire v_37927;
wire v_37928;
wire v_37929;
wire v_37930;
wire v_37931;
wire v_37932;
wire v_37933;
wire v_37934;
wire v_37935;
wire v_37936;
wire v_37937;
wire v_37938;
wire v_37939;
wire v_37940;
wire v_37941;
wire v_37942;
wire v_37943;
wire v_37944;
wire v_37945;
wire v_37946;
wire v_37947;
wire v_37948;
wire v_37949;
wire v_37950;
wire v_37951;
wire v_37952;
wire v_37953;
wire v_37954;
wire v_37955;
wire v_37956;
wire v_37957;
wire v_37958;
wire v_37959;
wire v_37960;
wire v_37961;
wire v_37962;
wire v_37963;
wire v_37964;
wire v_37965;
wire v_37966;
wire v_37967;
wire v_37968;
wire v_37969;
wire v_37970;
wire v_37971;
wire v_37972;
wire v_37973;
wire v_37974;
wire v_37975;
wire v_37976;
wire v_37977;
wire v_37978;
wire v_37979;
wire v_37980;
wire v_37981;
wire v_37982;
wire v_37983;
wire v_37984;
wire v_37985;
wire v_37986;
wire v_37987;
wire v_37988;
wire v_37989;
wire v_37990;
wire v_37991;
wire v_37992;
wire v_37993;
wire v_37994;
wire v_37995;
wire v_37996;
wire v_37997;
wire v_37998;
wire v_37999;
wire v_38000;
wire v_38001;
wire v_38002;
wire v_38003;
wire v_38004;
wire v_38005;
wire v_38006;
wire v_38007;
wire v_38008;
wire v_38009;
wire v_38010;
wire v_38011;
wire v_38012;
wire v_38013;
wire v_38014;
wire v_38015;
wire v_38016;
wire v_38017;
wire v_38018;
wire v_38019;
wire v_38020;
wire v_38021;
wire v_38022;
wire v_38023;
wire v_38024;
wire v_38025;
wire v_38026;
wire v_38027;
wire v_38028;
wire v_38029;
wire v_38030;
wire v_38031;
wire v_38032;
wire v_38033;
wire v_38034;
wire v_38035;
wire v_38036;
wire v_38037;
wire v_38038;
wire v_38039;
wire v_38040;
wire v_38041;
wire v_38042;
wire v_38043;
wire v_38044;
wire v_38045;
wire v_38046;
wire v_38047;
wire v_38048;
wire v_38049;
wire v_38050;
wire v_38051;
wire v_38052;
wire v_38053;
wire v_38054;
wire v_38055;
wire v_38056;
wire v_38057;
wire v_38058;
wire v_38059;
wire v_38060;
wire v_38061;
wire v_38062;
wire v_38063;
wire v_38064;
wire v_38065;
wire v_38066;
wire v_38067;
wire v_38068;
wire v_38069;
wire v_38070;
wire v_38071;
wire v_38072;
wire v_38073;
wire v_38074;
wire v_38075;
wire v_38076;
wire v_38077;
wire v_38078;
wire v_38079;
wire v_38080;
wire v_38081;
wire v_38082;
wire v_38083;
wire v_38084;
wire v_38085;
wire v_38086;
wire v_38087;
wire v_38088;
wire v_38089;
wire v_38090;
wire v_38091;
wire v_38092;
wire v_38093;
wire v_38094;
wire v_38095;
wire v_38096;
wire v_38097;
wire v_38098;
wire v_38099;
wire v_38100;
wire v_38101;
wire v_38102;
wire v_38103;
wire v_38104;
wire v_38105;
wire v_38106;
wire v_38107;
wire v_38108;
wire v_38109;
wire v_38110;
wire v_38111;
wire v_38112;
wire v_38113;
wire v_38114;
wire v_38115;
wire v_38116;
wire v_38117;
wire v_38118;
wire v_38119;
wire v_38120;
wire v_38121;
wire v_38122;
wire v_38123;
wire v_38124;
wire v_38125;
wire v_38126;
wire v_38127;
wire v_38128;
wire v_38130;
wire v_38131;
wire v_38132;
wire v_38133;
wire v_38134;
wire v_38135;
wire v_38136;
wire v_38137;
wire v_38138;
wire v_38139;
wire v_38140;
wire v_38141;
wire v_38142;
wire v_38143;
wire v_38144;
wire v_38145;
wire v_38146;
wire v_38147;
wire v_38148;
wire v_38149;
wire v_38150;
wire v_38151;
wire v_38152;
wire v_38153;
wire v_38154;
wire v_38155;
wire v_38156;
wire v_38157;
wire v_38158;
wire v_38159;
wire v_38160;
wire v_38161;
wire v_38162;
wire v_38163;
wire v_38164;
wire v_38165;
wire v_38166;
wire v_38167;
wire v_38168;
wire v_38169;
wire v_38170;
wire v_38171;
wire v_38172;
wire v_38173;
wire v_38174;
wire v_38175;
wire v_38176;
wire v_38177;
wire v_38178;
wire v_38179;
wire v_38180;
wire v_38181;
wire v_38182;
wire v_38183;
wire v_38184;
wire v_38185;
wire v_38186;
wire v_38187;
wire v_38188;
wire v_38189;
wire v_38190;
wire v_38191;
wire v_38192;
wire v_38193;
wire v_38194;
wire v_38195;
wire v_38196;
wire v_38197;
wire v_38198;
wire v_38199;
wire v_38200;
wire v_38201;
wire v_38202;
wire v_38203;
wire v_38204;
wire v_38205;
wire v_38206;
wire v_38207;
wire v_38208;
wire v_38209;
wire v_38210;
wire v_38211;
wire v_38212;
wire v_38213;
wire v_38214;
wire v_38215;
wire v_38216;
wire v_38217;
wire v_38218;
wire v_38219;
wire v_38220;
wire v_38221;
wire v_38222;
wire v_38223;
wire v_38224;
wire v_38225;
wire v_38226;
wire v_38227;
wire v_38228;
wire v_38229;
wire v_38230;
wire v_38231;
wire v_38232;
wire v_38233;
wire v_38234;
wire v_38235;
wire v_38236;
wire v_38237;
wire v_38238;
wire v_38239;
wire v_38240;
wire v_38241;
wire v_38242;
wire v_38243;
wire v_38244;
wire v_38245;
wire v_38246;
wire v_38247;
wire v_38248;
wire v_38249;
wire v_38250;
wire v_38251;
wire v_38252;
wire v_38253;
wire v_38254;
wire v_38255;
wire v_38256;
wire v_38257;
wire v_38258;
wire v_38259;
wire v_38260;
wire v_38261;
wire v_38262;
wire v_38263;
wire v_38264;
wire v_38265;
wire v_38266;
wire v_38267;
wire v_38268;
wire v_38269;
wire v_38270;
wire v_38271;
wire v_38272;
wire v_38273;
wire v_38274;
wire v_38275;
wire v_38276;
wire v_38277;
wire v_38278;
wire v_38279;
wire v_38280;
wire v_38281;
wire v_38282;
wire v_38283;
wire v_38284;
wire v_38285;
wire v_38286;
wire v_38287;
wire v_38288;
wire v_38289;
wire v_38290;
wire v_38291;
wire v_38292;
wire v_38293;
wire v_38294;
wire v_38295;
wire v_38296;
wire v_38297;
wire v_38298;
wire v_38299;
wire v_38300;
wire v_38301;
wire v_38302;
wire v_38303;
wire v_38304;
wire v_38305;
wire v_38306;
wire v_38307;
wire v_38308;
wire v_38309;
wire v_38310;
wire v_38311;
wire v_38312;
wire v_38313;
wire v_38314;
wire v_38315;
wire v_38316;
wire v_38317;
wire v_38318;
wire v_38319;
wire v_38320;
wire v_38321;
wire v_38322;
wire v_38323;
wire v_38324;
wire v_38325;
wire v_38326;
wire v_38327;
wire v_38328;
wire v_38329;
wire v_38330;
wire v_38331;
wire v_38332;
wire v_38333;
wire v_38334;
wire v_38335;
wire v_38336;
wire v_38337;
wire v_38338;
wire v_38339;
wire v_38340;
wire v_38341;
wire v_38342;
wire v_38343;
wire v_38344;
wire v_38345;
wire v_38346;
wire v_38347;
wire v_38348;
wire v_38349;
wire v_38350;
wire v_38351;
wire v_38352;
wire v_38353;
wire v_38354;
wire v_38355;
wire v_38356;
wire v_38357;
wire v_38358;
wire v_38359;
wire v_38360;
wire v_38361;
wire v_38362;
wire v_38363;
wire v_38364;
wire v_38365;
wire v_38366;
wire v_38367;
wire v_38368;
wire v_38369;
wire v_38370;
wire v_38371;
wire v_38373;
wire v_38374;
wire v_38375;
wire v_38376;
wire v_38377;
wire v_38378;
wire v_38379;
wire v_38380;
wire v_38381;
wire v_38382;
wire v_38383;
wire v_38384;
wire v_38385;
wire v_38386;
wire v_38387;
wire v_38388;
wire v_38389;
wire v_38390;
wire v_38391;
wire v_38392;
wire v_38393;
wire v_38394;
wire v_38395;
wire v_38396;
wire v_38397;
wire v_38398;
wire v_38399;
wire v_38400;
wire v_38401;
wire v_38402;
wire v_38403;
wire v_38404;
wire v_38405;
wire v_38406;
wire v_38407;
wire v_38408;
wire v_38409;
wire v_38410;
wire v_38411;
wire v_38412;
wire v_38413;
wire v_38414;
wire v_38415;
wire v_38416;
wire v_38417;
wire v_38418;
wire v_38419;
wire v_38420;
wire v_38421;
wire v_38422;
wire v_38423;
wire v_38424;
wire v_38425;
wire v_38426;
wire v_38427;
wire v_38428;
wire v_38429;
wire v_38430;
wire v_38431;
wire v_38432;
wire v_38433;
wire v_38434;
wire v_38435;
wire v_38436;
wire v_38437;
wire v_38438;
wire v_38439;
wire v_38440;
wire v_38441;
wire v_38442;
wire v_38443;
wire v_38444;
wire v_38445;
wire v_38446;
wire v_38447;
wire v_38448;
wire v_38449;
wire v_38450;
wire v_38451;
wire v_38452;
wire v_38453;
wire v_38454;
wire v_38455;
wire v_38456;
wire v_38457;
wire v_38458;
wire v_38459;
wire v_38460;
wire v_38461;
wire v_38462;
wire v_38463;
wire v_38464;
wire v_38465;
wire v_38466;
wire v_38467;
wire v_38468;
wire v_38469;
wire v_38470;
wire v_38471;
wire v_38472;
wire v_38473;
wire v_38474;
wire v_38475;
wire v_38476;
wire v_38477;
wire v_38478;
wire v_38479;
wire v_38480;
wire v_38481;
wire v_38482;
wire v_38483;
wire v_38484;
wire v_38485;
wire v_38486;
wire v_38487;
wire v_38488;
wire v_38489;
wire v_38490;
wire v_38491;
wire v_38492;
wire v_38493;
wire v_38494;
wire v_38495;
wire v_38496;
wire v_38497;
wire v_38498;
wire v_38499;
wire v_38500;
wire v_38501;
wire v_38502;
wire v_38503;
wire v_38504;
wire v_38505;
wire v_38506;
wire v_38507;
wire v_38508;
wire v_38509;
wire v_38510;
wire v_38511;
wire v_38512;
wire v_38513;
wire v_38514;
wire v_38515;
wire v_38516;
wire v_38517;
wire v_38518;
wire v_38519;
wire v_38520;
wire v_38521;
wire v_38522;
wire v_38523;
wire v_38524;
wire v_38525;
wire v_38526;
wire v_38527;
wire v_38528;
wire v_38529;
wire v_38530;
wire v_38531;
wire v_38532;
wire v_38533;
wire v_38534;
wire v_38535;
wire v_38536;
wire v_38537;
wire v_38538;
wire v_38539;
wire v_38540;
wire v_38541;
wire v_38542;
wire v_38543;
wire v_38544;
wire v_38545;
wire v_38546;
wire v_38547;
wire v_38548;
wire v_38549;
wire v_38550;
wire v_38551;
wire v_38552;
wire v_38553;
wire v_38554;
wire v_38555;
wire v_38556;
wire v_38557;
wire v_38558;
wire v_38559;
wire v_38560;
wire v_38561;
wire v_38562;
wire v_38563;
wire v_38564;
wire v_38565;
wire v_38566;
wire v_38567;
wire v_38568;
wire v_38569;
wire v_38570;
wire v_38571;
wire v_38572;
wire v_38573;
wire v_38574;
wire v_38575;
wire v_38576;
wire v_38577;
wire v_38578;
wire v_38579;
wire v_38580;
wire v_38581;
wire v_38582;
wire v_38583;
wire v_38584;
wire v_38585;
wire v_38586;
wire v_38587;
wire v_38588;
wire v_38589;
wire v_38590;
wire v_38591;
wire v_38592;
wire v_38593;
wire v_38594;
wire v_38595;
wire v_38596;
wire v_38597;
wire v_38598;
wire v_38599;
wire v_38600;
wire v_38601;
wire v_38602;
wire v_38603;
wire v_38604;
wire v_38605;
wire v_38606;
wire v_38607;
wire v_38608;
wire v_38609;
wire v_38610;
wire v_38611;
wire v_38612;
wire v_38613;
wire v_38614;
wire v_38616;
wire v_38617;
wire v_38618;
wire v_38619;
wire v_38620;
wire v_38621;
wire v_38622;
wire v_38623;
wire v_38624;
wire v_38625;
wire v_38626;
wire v_38627;
wire v_38628;
wire v_38629;
wire v_38630;
wire v_38631;
wire v_38632;
wire v_38633;
wire v_38634;
wire v_38635;
wire v_38636;
wire v_38637;
wire v_38638;
wire v_38639;
wire v_38640;
wire v_38641;
wire v_38642;
wire v_38643;
wire v_38644;
wire v_38645;
wire v_38646;
wire v_38647;
wire v_38648;
wire v_38649;
wire v_38650;
wire v_38651;
wire v_38652;
wire v_38653;
wire v_38654;
wire v_38655;
wire v_38656;
wire v_38657;
wire v_38658;
wire v_38659;
wire v_38660;
wire v_38661;
wire v_38662;
wire v_38663;
wire v_38664;
wire v_38665;
wire v_38666;
wire v_38667;
wire v_38668;
wire v_38669;
wire v_38670;
wire v_38671;
wire v_38672;
wire v_38673;
wire v_38674;
wire v_38675;
wire v_38676;
wire v_38677;
wire v_38678;
wire v_38679;
wire v_38680;
wire v_38681;
wire v_38682;
wire v_38683;
wire v_38684;
wire v_38685;
wire v_38686;
wire v_38687;
wire v_38688;
wire v_38689;
wire v_38690;
wire v_38691;
wire v_38692;
wire v_38693;
wire v_38694;
wire v_38695;
wire v_38696;
wire v_38697;
wire v_38698;
wire v_38699;
wire v_38700;
wire v_38701;
wire v_38702;
wire v_38703;
wire v_38704;
wire v_38705;
wire v_38706;
wire v_38707;
wire v_38708;
wire v_38709;
wire v_38710;
wire v_38711;
wire v_38712;
wire v_38713;
wire v_38714;
wire v_38715;
wire v_38716;
wire v_38717;
wire v_38718;
wire v_38719;
wire v_38720;
wire v_38721;
wire v_38722;
wire v_38723;
wire v_38724;
wire v_38725;
wire v_38726;
wire v_38727;
wire v_38728;
wire v_38729;
wire v_38730;
wire v_38731;
wire v_38732;
wire v_38733;
wire v_38734;
wire v_38735;
wire v_38736;
wire v_38737;
wire v_38738;
wire v_38739;
wire v_38740;
wire v_38741;
wire v_38742;
wire v_38743;
wire v_38744;
wire v_38745;
wire v_38746;
wire v_38747;
wire v_38748;
wire v_38749;
wire v_38750;
wire v_38751;
wire v_38752;
wire v_38753;
wire v_38754;
wire v_38755;
wire v_38756;
wire v_38757;
wire v_38758;
wire v_38759;
wire v_38760;
wire v_38761;
wire v_38762;
wire v_38763;
wire v_38764;
wire v_38765;
wire v_38766;
wire v_38767;
wire v_38768;
wire v_38769;
wire v_38770;
wire v_38771;
wire v_38772;
wire v_38773;
wire v_38774;
wire v_38775;
wire v_38776;
wire v_38777;
wire v_38778;
wire v_38779;
wire v_38780;
wire v_38781;
wire v_38782;
wire v_38783;
wire v_38784;
wire v_38785;
wire v_38786;
wire v_38787;
wire v_38788;
wire v_38789;
wire v_38790;
wire v_38791;
wire v_38792;
wire v_38793;
wire v_38794;
wire v_38795;
wire v_38796;
wire v_38797;
wire v_38798;
wire v_38799;
wire v_38800;
wire v_38801;
wire v_38802;
wire v_38803;
wire v_38804;
wire v_38805;
wire v_38806;
wire v_38807;
wire v_38808;
wire v_38809;
wire v_38810;
wire v_38811;
wire v_38812;
wire v_38813;
wire v_38814;
wire v_38815;
wire v_38816;
wire v_38817;
wire v_38818;
wire v_38819;
wire v_38820;
wire v_38821;
wire v_38822;
wire v_38823;
wire v_38824;
wire v_38825;
wire v_38826;
wire v_38827;
wire v_38828;
wire v_38829;
wire v_38830;
wire v_38831;
wire v_38832;
wire v_38833;
wire v_38834;
wire v_38835;
wire v_38836;
wire v_38837;
wire v_38838;
wire v_38839;
wire v_38840;
wire v_38841;
wire v_38842;
wire v_38843;
wire v_38844;
wire v_38845;
wire v_38846;
wire v_38847;
wire v_38848;
wire v_38849;
wire v_38850;
wire v_38851;
wire v_38852;
wire v_38853;
wire v_38854;
wire v_38855;
wire v_38856;
wire v_38857;
wire v_38859;
wire v_38860;
wire v_38861;
wire v_38862;
wire v_38863;
wire v_38864;
wire v_38865;
wire v_38866;
wire v_38867;
wire v_38868;
wire v_38869;
wire v_38870;
wire v_38871;
wire v_38872;
wire v_38873;
wire v_38874;
wire v_38875;
wire v_38876;
wire v_38877;
wire v_38878;
wire v_38879;
wire v_38880;
wire v_38881;
wire v_38882;
wire v_38883;
wire v_38884;
wire v_38885;
wire v_38886;
wire v_38887;
wire v_38888;
wire v_38889;
wire v_38890;
wire v_38891;
wire v_38892;
wire v_38893;
wire v_38894;
wire v_38895;
wire v_38896;
wire v_38897;
wire v_38898;
wire v_38899;
wire v_38900;
wire v_38901;
wire v_38902;
wire v_38903;
wire v_38904;
wire v_38905;
wire v_38906;
wire v_38907;
wire v_38908;
wire v_38909;
wire v_38910;
wire v_38911;
wire v_38912;
wire v_38913;
wire v_38914;
wire v_38915;
wire v_38916;
wire v_38917;
wire v_38918;
wire v_38919;
wire v_38920;
wire v_38921;
wire v_38922;
wire v_38923;
wire v_38924;
wire v_38925;
wire v_38926;
wire v_38927;
wire v_38928;
wire v_38929;
wire v_38930;
wire v_38931;
wire v_38932;
wire v_38933;
wire v_38934;
wire v_38935;
wire v_38936;
wire v_38937;
wire v_38938;
wire v_38939;
wire v_38940;
wire v_38941;
wire v_38942;
wire v_38943;
wire v_38944;
wire v_38945;
wire v_38946;
wire v_38947;
wire v_38948;
wire v_38949;
wire v_38950;
wire v_38951;
wire v_38952;
wire v_38953;
wire v_38954;
wire v_38955;
wire v_38956;
wire v_38957;
wire v_38958;
wire v_38959;
wire v_38960;
wire v_38961;
wire v_38962;
wire v_38963;
wire v_38964;
wire v_38965;
wire v_38966;
wire v_38967;
wire v_38968;
wire v_38969;
wire v_38970;
wire v_38971;
wire v_38972;
wire v_38973;
wire v_38974;
wire v_38975;
wire v_38976;
wire v_38977;
wire v_38978;
wire v_38979;
wire v_38980;
wire v_38981;
wire v_38982;
wire v_38983;
wire v_38984;
wire v_38985;
wire v_38986;
wire v_38987;
wire v_38988;
wire v_38989;
wire v_38990;
wire v_38991;
wire v_38992;
wire v_38993;
wire v_38994;
wire v_38995;
wire v_38996;
wire v_38997;
wire v_38998;
wire v_38999;
wire v_39000;
wire v_39001;
wire v_39002;
wire v_39003;
wire v_39004;
wire v_39005;
wire v_39006;
wire v_39007;
wire v_39008;
wire v_39009;
wire v_39010;
wire v_39011;
wire v_39012;
wire v_39013;
wire v_39014;
wire v_39015;
wire v_39016;
wire v_39017;
wire v_39018;
wire v_39019;
wire v_39020;
wire v_39021;
wire v_39022;
wire v_39023;
wire v_39024;
wire v_39025;
wire v_39026;
wire v_39027;
wire v_39028;
wire v_39029;
wire v_39030;
wire v_39031;
wire v_39032;
wire v_39033;
wire v_39034;
wire v_39035;
wire v_39036;
wire v_39037;
wire v_39038;
wire v_39039;
wire v_39040;
wire v_39041;
wire v_39042;
wire v_39043;
wire v_39044;
wire v_39045;
wire v_39046;
wire v_39047;
wire v_39048;
wire v_39049;
wire v_39050;
wire v_39051;
wire v_39052;
wire v_39053;
wire v_39054;
wire v_39055;
wire v_39056;
wire v_39057;
wire v_39058;
wire v_39059;
wire v_39060;
wire v_39061;
wire v_39062;
wire v_39063;
wire v_39064;
wire v_39065;
wire v_39066;
wire v_39067;
wire v_39068;
wire v_39069;
wire v_39070;
wire v_39071;
wire v_39072;
wire v_39073;
wire v_39074;
wire v_39075;
wire v_39076;
wire v_39077;
wire v_39078;
wire v_39079;
wire v_39080;
wire v_39081;
wire v_39082;
wire v_39083;
wire v_39084;
wire v_39085;
wire v_39086;
wire v_39087;
wire v_39088;
wire v_39089;
wire v_39090;
wire v_39091;
wire v_39092;
wire v_39093;
wire v_39094;
wire v_39095;
wire v_39096;
wire v_39097;
wire v_39098;
wire v_39099;
wire v_39100;
wire v_39102;
wire v_39103;
wire v_39104;
wire v_39105;
wire v_39106;
wire v_39107;
wire v_39108;
wire v_39109;
wire v_39110;
wire v_39111;
wire v_39112;
wire v_39113;
wire v_39114;
wire v_39115;
wire v_39116;
wire v_39117;
wire v_39118;
wire v_39119;
wire v_39120;
wire v_39121;
wire v_39122;
wire v_39123;
wire v_39124;
wire v_39125;
wire v_39126;
wire v_39127;
wire v_39128;
wire v_39129;
wire v_39130;
wire v_39131;
wire v_39132;
wire v_39133;
wire v_39134;
wire v_39135;
wire v_39136;
wire v_39137;
wire v_39138;
wire v_39139;
wire v_39140;
wire v_39141;
wire v_39142;
wire v_39143;
wire v_39144;
wire v_39145;
wire v_39146;
wire v_39147;
wire v_39148;
wire v_39149;
wire v_39150;
wire v_39151;
wire v_39152;
wire v_39153;
wire v_39154;
wire v_39155;
wire v_39156;
wire v_39157;
wire v_39158;
wire v_39159;
wire v_39160;
wire v_39161;
wire v_39162;
wire v_39163;
wire v_39164;
wire v_39165;
wire v_39166;
wire v_39167;
wire v_39168;
wire v_39169;
wire v_39170;
wire v_39171;
wire v_39172;
wire v_39173;
wire v_39174;
wire v_39175;
wire v_39176;
wire v_39177;
wire v_39178;
wire v_39179;
wire v_39180;
wire v_39181;
wire v_39182;
wire v_39183;
wire v_39184;
wire v_39185;
wire v_39186;
wire v_39187;
wire v_39188;
wire v_39189;
wire v_39190;
wire v_39191;
wire v_39192;
wire v_39193;
wire v_39194;
wire v_39195;
wire v_39196;
wire v_39197;
wire v_39198;
wire v_39199;
wire v_39200;
wire v_39201;
wire v_39202;
wire v_39203;
wire v_39204;
wire v_39205;
wire v_39206;
wire v_39207;
wire v_39208;
wire v_39209;
wire v_39210;
wire v_39211;
wire v_39212;
wire v_39213;
wire v_39214;
wire v_39215;
wire v_39216;
wire v_39217;
wire v_39218;
wire v_39219;
wire v_39220;
wire v_39221;
wire v_39222;
wire v_39223;
wire v_39224;
wire v_39225;
wire v_39226;
wire v_39227;
wire v_39228;
wire v_39229;
wire v_39230;
wire v_39231;
wire v_39232;
wire v_39233;
wire v_39234;
wire v_39235;
wire v_39236;
wire v_39237;
wire v_39238;
wire v_39239;
wire v_39240;
wire v_39241;
wire v_39242;
wire v_39243;
wire v_39244;
wire v_39245;
wire v_39246;
wire v_39247;
wire v_39248;
wire v_39249;
wire v_39250;
wire v_39251;
wire v_39252;
wire v_39253;
wire v_39254;
wire v_39255;
wire v_39256;
wire v_39257;
wire v_39258;
wire v_39259;
wire v_39260;
wire v_39261;
wire v_39262;
wire v_39263;
wire v_39264;
wire v_39265;
wire v_39266;
wire v_39267;
wire v_39268;
wire v_39269;
wire v_39270;
wire v_39271;
wire v_39272;
wire v_39273;
wire v_39274;
wire v_39275;
wire v_39276;
wire v_39277;
wire v_39278;
wire v_39279;
wire v_39280;
wire v_39281;
wire v_39282;
wire v_39283;
wire v_39284;
wire v_39285;
wire v_39286;
wire v_39287;
wire v_39288;
wire v_39289;
wire v_39290;
wire v_39291;
wire v_39292;
wire v_39293;
wire v_39294;
wire v_39295;
wire v_39296;
wire v_39297;
wire v_39298;
wire v_39299;
wire v_39300;
wire v_39301;
wire v_39302;
wire v_39303;
wire v_39304;
wire v_39305;
wire v_39306;
wire v_39307;
wire v_39308;
wire v_39309;
wire v_39310;
wire v_39311;
wire v_39312;
wire v_39313;
wire v_39314;
wire v_39315;
wire v_39316;
wire v_39317;
wire v_39318;
wire v_39319;
wire v_39320;
wire v_39321;
wire v_39322;
wire v_39323;
wire v_39324;
wire v_39325;
wire v_39326;
wire v_39327;
wire v_39328;
wire v_39329;
wire v_39330;
wire v_39331;
wire v_39332;
wire v_39333;
wire v_39334;
wire v_39335;
wire v_39336;
wire v_39337;
wire v_39338;
wire v_39339;
wire v_39340;
wire v_39341;
wire v_39342;
wire v_39343;
wire v_39345;
wire v_39346;
wire v_39347;
wire v_39348;
wire v_39349;
wire v_39350;
wire v_39351;
wire v_39352;
wire v_39353;
wire v_39354;
wire v_39355;
wire v_39356;
wire v_39357;
wire v_39358;
wire v_39359;
wire v_39360;
wire v_39361;
wire v_39362;
wire v_39363;
wire v_39364;
wire v_39365;
wire v_39366;
wire v_39367;
wire v_39368;
wire v_39369;
wire v_39370;
wire v_39371;
wire v_39372;
wire v_39373;
wire v_39374;
wire v_39375;
wire v_39376;
wire v_39377;
wire v_39378;
wire v_39379;
wire v_39380;
wire v_39381;
wire v_39382;
wire v_39383;
wire v_39384;
wire v_39385;
wire v_39386;
wire v_39387;
wire v_39388;
wire v_39389;
wire v_39390;
wire v_39391;
wire v_39392;
wire v_39393;
wire v_39394;
wire v_39395;
wire v_39396;
wire v_39397;
wire v_39398;
wire v_39399;
wire v_39400;
wire v_39401;
wire v_39402;
wire v_39403;
wire v_39404;
wire v_39405;
wire v_39406;
wire v_39407;
wire v_39408;
wire v_39409;
wire v_39410;
wire v_39411;
wire v_39412;
wire v_39413;
wire v_39414;
wire v_39415;
wire v_39416;
wire v_39417;
wire v_39418;
wire v_39419;
wire v_39420;
wire v_39421;
wire v_39422;
wire v_39423;
wire v_39424;
wire v_39425;
wire v_39426;
wire v_39427;
wire v_39428;
wire v_39429;
wire v_39430;
wire v_39431;
wire v_39432;
wire v_39433;
wire v_39434;
wire v_39435;
wire v_39436;
wire v_39437;
wire v_39438;
wire v_39439;
wire v_39440;
wire v_39441;
wire v_39442;
wire v_39443;
wire v_39444;
wire v_39445;
wire v_39446;
wire v_39447;
wire v_39448;
wire v_39449;
wire v_39450;
wire v_39451;
wire v_39452;
wire v_39453;
wire v_39454;
wire v_39455;
wire v_39456;
wire v_39457;
wire v_39458;
wire v_39459;
wire v_39460;
wire v_39461;
wire v_39462;
wire v_39463;
wire v_39464;
wire v_39465;
wire v_39466;
wire v_39467;
wire v_39468;
wire v_39469;
wire v_39470;
wire v_39471;
wire v_39472;
wire v_39473;
wire v_39474;
wire v_39475;
wire v_39476;
wire v_39477;
wire v_39478;
wire v_39479;
wire v_39480;
wire v_39481;
wire v_39482;
wire v_39483;
wire v_39484;
wire v_39485;
wire v_39486;
wire v_39487;
wire v_39488;
wire v_39489;
wire v_39490;
wire v_39491;
wire v_39492;
wire v_39493;
wire v_39494;
wire v_39495;
wire v_39496;
wire v_39497;
wire v_39498;
wire v_39499;
wire v_39500;
wire v_39501;
wire v_39502;
wire v_39503;
wire v_39504;
wire v_39505;
wire v_39506;
wire v_39507;
wire v_39508;
wire v_39509;
wire v_39510;
wire v_39511;
wire v_39512;
wire v_39513;
wire v_39514;
wire v_39515;
wire v_39516;
wire v_39517;
wire v_39518;
wire v_39519;
wire v_39520;
wire v_39521;
wire v_39522;
wire v_39523;
wire v_39524;
wire v_39525;
wire v_39526;
wire v_39527;
wire v_39528;
wire v_39529;
wire v_39530;
wire v_39531;
wire v_39532;
wire v_39533;
wire v_39534;
wire v_39535;
wire v_39536;
wire v_39537;
wire v_39538;
wire v_39539;
wire v_39540;
wire v_39541;
wire v_39542;
wire v_39543;
wire v_39544;
wire v_39545;
wire v_39546;
wire v_39547;
wire v_39548;
wire v_39549;
wire v_39550;
wire v_39551;
wire v_39552;
wire v_39553;
wire v_39554;
wire v_39555;
wire v_39556;
wire v_39557;
wire v_39558;
wire v_39559;
wire v_39560;
wire v_39561;
wire v_39562;
wire v_39563;
wire v_39564;
wire v_39565;
wire v_39566;
wire v_39567;
wire v_39568;
wire v_39569;
wire v_39570;
wire v_39571;
wire v_39572;
wire v_39573;
wire v_39574;
wire v_39575;
wire v_39576;
wire v_39577;
wire v_39578;
wire v_39579;
wire v_39580;
wire v_39581;
wire v_39582;
wire v_39583;
wire v_39584;
wire v_39585;
wire v_39586;
wire v_39588;
wire v_39589;
wire v_39590;
wire v_39591;
wire v_39592;
wire v_39593;
wire v_39594;
wire v_39595;
wire v_39596;
wire v_39597;
wire v_39598;
wire v_39599;
wire v_39600;
wire v_39601;
wire v_39602;
wire v_39603;
wire v_39604;
wire v_39605;
wire v_39606;
wire v_39607;
wire v_39608;
wire v_39609;
wire v_39610;
wire v_39611;
wire v_39612;
wire v_39613;
wire v_39614;
wire v_39615;
wire v_39616;
wire v_39617;
wire v_39618;
wire v_39619;
wire v_39620;
wire v_39621;
wire v_39622;
wire v_39623;
wire v_39624;
wire v_39625;
wire v_39626;
wire v_39627;
wire v_39628;
wire v_39629;
wire v_39630;
wire v_39631;
wire v_39632;
wire v_39633;
wire v_39634;
wire v_39635;
wire v_39636;
wire v_39637;
wire v_39638;
wire v_39639;
wire v_39640;
wire v_39641;
wire v_39642;
wire v_39643;
wire v_39644;
wire v_39645;
wire v_39646;
wire v_39647;
wire v_39648;
wire v_39649;
wire v_39650;
wire v_39651;
wire v_39652;
wire v_39653;
wire v_39654;
wire v_39655;
wire v_39656;
wire v_39657;
wire v_39658;
wire v_39659;
wire v_39660;
wire v_39661;
wire v_39662;
wire v_39663;
wire v_39664;
wire v_39665;
wire v_39666;
wire v_39667;
wire v_39668;
wire v_39669;
wire v_39670;
wire v_39671;
wire v_39672;
wire v_39673;
wire v_39674;
wire v_39675;
wire v_39676;
wire v_39677;
wire v_39678;
wire v_39679;
wire v_39680;
wire v_39681;
wire v_39682;
wire v_39683;
wire v_39684;
wire v_39685;
wire v_39686;
wire v_39687;
wire v_39688;
wire v_39689;
wire v_39690;
wire v_39691;
wire v_39692;
wire v_39693;
wire v_39694;
wire v_39695;
wire v_39696;
wire v_39697;
wire v_39698;
wire v_39699;
wire v_39700;
wire v_39701;
wire v_39702;
wire v_39703;
wire v_39704;
wire v_39705;
wire v_39706;
wire v_39707;
wire v_39708;
wire v_39709;
wire v_39710;
wire v_39711;
wire v_39712;
wire v_39713;
wire v_39714;
wire v_39715;
wire v_39716;
wire v_39717;
wire v_39718;
wire v_39719;
wire v_39720;
wire v_39721;
wire v_39722;
wire v_39723;
wire v_39724;
wire v_39725;
wire v_39726;
wire v_39727;
wire v_39728;
wire v_39729;
wire v_39730;
wire v_39731;
wire v_39732;
wire v_39733;
wire v_39734;
wire v_39735;
wire v_39736;
wire v_39737;
wire v_39738;
wire v_39739;
wire v_39740;
wire v_39741;
wire v_39742;
wire v_39743;
wire v_39744;
wire v_39745;
wire v_39746;
wire v_39747;
wire v_39748;
wire v_39749;
wire v_39750;
wire v_39751;
wire v_39752;
wire v_39753;
wire v_39754;
wire v_39755;
wire v_39756;
wire v_39757;
wire v_39758;
wire v_39759;
wire v_39760;
wire v_39761;
wire v_39762;
wire v_39763;
wire v_39764;
wire v_39765;
wire v_39766;
wire v_39767;
wire v_39768;
wire v_39769;
wire v_39770;
wire v_39771;
wire v_39772;
wire v_39773;
wire v_39774;
wire v_39775;
wire v_39776;
wire v_39777;
wire v_39778;
wire v_39779;
wire v_39780;
wire v_39781;
wire v_39782;
wire v_39783;
wire v_39784;
wire v_39785;
wire v_39786;
wire v_39787;
wire v_39788;
wire v_39789;
wire v_39790;
wire v_39791;
wire v_39792;
wire v_39793;
wire v_39794;
wire v_39795;
wire v_39796;
wire v_39797;
wire v_39798;
wire v_39799;
wire v_39800;
wire v_39801;
wire v_39802;
wire v_39803;
wire v_39804;
wire v_39805;
wire v_39806;
wire v_39807;
wire v_39808;
wire v_39809;
wire v_39810;
wire v_39811;
wire v_39812;
wire v_39813;
wire v_39814;
wire v_39815;
wire v_39816;
wire v_39817;
wire v_39818;
wire v_39819;
wire v_39820;
wire v_39821;
wire v_39822;
wire v_39823;
wire v_39824;
wire v_39825;
wire v_39826;
wire v_39827;
wire v_39828;
wire v_39829;
wire v_39831;
wire v_39832;
wire v_39833;
wire v_39834;
wire v_39835;
wire v_39836;
wire v_39837;
wire v_39838;
wire v_39839;
wire v_39840;
wire v_39841;
wire v_39842;
wire v_39843;
wire v_39844;
wire v_39845;
wire v_39846;
wire v_39847;
wire v_39848;
wire v_39849;
wire v_39850;
wire v_39851;
wire v_39852;
wire v_39853;
wire v_39854;
wire v_39855;
wire v_39856;
wire v_39857;
wire v_39858;
wire v_39859;
wire v_39860;
wire v_39861;
wire v_39862;
wire v_39863;
wire v_39864;
wire v_39865;
wire v_39866;
wire v_39867;
wire v_39868;
wire v_39869;
wire v_39870;
wire v_39871;
wire v_39872;
wire v_39873;
wire v_39874;
wire v_39875;
wire v_39876;
wire v_39877;
wire v_39878;
wire v_39879;
wire v_39880;
wire v_39881;
wire v_39882;
wire v_39883;
wire v_39884;
wire v_39885;
wire v_39886;
wire v_39887;
wire v_39888;
wire v_39889;
wire v_39890;
wire v_39891;
wire v_39892;
wire v_39893;
wire v_39894;
wire v_39895;
wire v_39896;
wire v_39897;
wire v_39898;
wire v_39899;
wire v_39900;
wire v_39901;
wire v_39902;
wire v_39903;
wire v_39904;
wire v_39905;
wire v_39906;
wire v_39907;
wire v_39908;
wire v_39909;
wire v_39910;
wire v_39911;
wire v_39912;
wire v_39913;
wire v_39914;
wire v_39915;
wire v_39916;
wire v_39917;
wire v_39918;
wire v_39919;
wire v_39920;
wire v_39921;
wire v_39922;
wire v_39923;
wire v_39924;
wire v_39925;
wire v_39926;
wire v_39927;
wire v_39928;
wire v_39929;
wire v_39930;
wire v_39931;
wire v_39932;
wire v_39933;
wire v_39934;
wire v_39935;
wire v_39936;
wire v_39937;
wire v_39938;
wire v_39939;
wire v_39940;
wire v_39941;
wire v_39942;
wire v_39943;
wire v_39944;
wire v_39945;
wire v_39946;
wire v_39947;
wire v_39948;
wire v_39949;
wire v_39950;
wire v_39951;
wire v_39952;
wire v_39953;
wire v_39954;
wire v_39955;
wire v_39956;
wire v_39957;
wire v_39958;
wire v_39959;
wire v_39960;
wire v_39961;
wire v_39962;
wire v_39963;
wire v_39964;
wire v_39965;
wire v_39966;
wire v_39967;
wire v_39968;
wire v_39969;
wire v_39970;
wire v_39971;
wire v_39972;
wire v_39973;
wire v_39974;
wire v_39975;
wire v_39976;
wire v_39977;
wire v_39978;
wire v_39979;
wire v_39980;
wire v_39981;
wire v_39982;
wire v_39983;
wire v_39984;
wire v_39985;
wire v_39986;
wire v_39987;
wire v_39988;
wire v_39989;
wire v_39990;
wire v_39991;
wire v_39992;
wire v_39993;
wire v_39994;
wire v_39995;
wire v_39996;
wire v_39997;
wire v_39998;
wire v_39999;
wire v_40000;
wire v_40001;
wire v_40002;
wire v_40003;
wire v_40004;
wire v_40005;
wire v_40006;
wire v_40007;
wire v_40008;
wire v_40009;
wire v_40010;
wire v_40011;
wire v_40012;
wire v_40013;
wire v_40014;
wire v_40015;
wire v_40016;
wire v_40017;
wire v_40018;
wire v_40019;
wire v_40020;
wire v_40021;
wire v_40022;
wire v_40023;
wire v_40024;
wire v_40025;
wire v_40026;
wire v_40027;
wire v_40028;
wire v_40029;
wire v_40030;
wire v_40031;
wire v_40032;
wire v_40033;
wire v_40034;
wire v_40035;
wire v_40036;
wire v_40037;
wire v_40038;
wire v_40039;
wire v_40040;
wire v_40041;
wire v_40042;
wire v_40043;
wire v_40044;
wire v_40045;
wire v_40046;
wire v_40047;
wire v_40048;
wire v_40049;
wire v_40050;
wire v_40051;
wire v_40052;
wire v_40053;
wire v_40054;
wire v_40055;
wire v_40056;
wire v_40057;
wire v_40058;
wire v_40059;
wire v_40060;
wire v_40061;
wire v_40062;
wire v_40063;
wire v_40064;
wire v_40065;
wire v_40066;
wire v_40067;
wire v_40068;
wire v_40069;
wire v_40070;
wire v_40071;
wire v_40072;
wire v_40074;
wire v_40075;
wire v_40076;
wire v_40077;
wire v_40078;
wire v_40079;
wire v_40080;
wire v_40081;
wire v_40082;
wire v_40083;
wire v_40084;
wire v_40085;
wire v_40086;
wire v_40087;
wire v_40088;
wire v_40089;
wire v_40090;
wire v_40091;
wire v_40092;
wire v_40093;
wire v_40094;
wire v_40095;
wire v_40096;
wire v_40097;
wire v_40098;
wire v_40099;
wire v_40100;
wire v_40101;
wire v_40102;
wire v_40103;
wire v_40104;
wire v_40105;
wire v_40106;
wire v_40107;
wire v_40108;
wire v_40109;
wire v_40110;
wire v_40111;
wire v_40112;
wire v_40113;
wire v_40114;
wire v_40115;
wire v_40116;
wire v_40117;
wire v_40118;
wire v_40119;
wire v_40120;
wire v_40121;
wire v_40122;
wire v_40123;
wire v_40124;
wire v_40125;
wire v_40126;
wire v_40127;
wire v_40128;
wire v_40129;
wire v_40130;
wire v_40131;
wire v_40132;
wire v_40133;
wire v_40134;
wire v_40135;
wire v_40136;
wire v_40137;
wire v_40138;
wire v_40139;
wire v_40140;
wire v_40141;
wire v_40142;
wire v_40143;
wire v_40144;
wire v_40145;
wire v_40146;
wire v_40147;
wire v_40148;
wire v_40149;
wire v_40150;
wire v_40151;
wire v_40152;
wire v_40153;
wire v_40154;
wire v_40155;
wire v_40156;
wire v_40157;
wire v_40158;
wire v_40159;
wire v_40160;
wire v_40161;
wire v_40162;
wire v_40163;
wire v_40164;
wire v_40165;
wire v_40166;
wire v_40167;
wire v_40168;
wire v_40169;
wire v_40170;
wire v_40171;
wire v_40172;
wire v_40173;
wire v_40174;
wire v_40175;
wire v_40176;
wire v_40177;
wire v_40178;
wire v_40179;
wire v_40180;
wire v_40181;
wire v_40182;
wire v_40183;
wire v_40184;
wire v_40185;
wire v_40186;
wire v_40187;
wire v_40188;
wire v_40189;
wire v_40190;
wire v_40191;
wire v_40192;
wire v_40193;
wire v_40194;
wire v_40195;
wire v_40196;
wire v_40197;
wire v_40198;
wire v_40199;
wire v_40200;
wire v_40201;
wire v_40202;
wire v_40203;
wire v_40204;
wire v_40205;
wire v_40206;
wire v_40207;
wire v_40208;
wire v_40209;
wire v_40210;
wire v_40211;
wire v_40212;
wire v_40213;
wire v_40214;
wire v_40215;
wire v_40216;
wire v_40217;
wire v_40218;
wire v_40219;
wire v_40220;
wire v_40221;
wire v_40222;
wire v_40223;
wire v_40224;
wire v_40225;
wire v_40226;
wire v_40227;
wire v_40228;
wire v_40229;
wire v_40230;
wire v_40231;
wire v_40232;
wire v_40233;
wire v_40234;
wire v_40235;
wire v_40236;
wire v_40237;
wire v_40238;
wire v_40239;
wire v_40240;
wire v_40241;
wire v_40242;
wire v_40243;
wire v_40244;
wire v_40245;
wire v_40246;
wire v_40247;
wire v_40248;
wire v_40249;
wire v_40250;
wire v_40251;
wire v_40252;
wire v_40253;
wire v_40254;
wire v_40255;
wire v_40256;
wire v_40257;
wire v_40258;
wire v_40259;
wire v_40260;
wire v_40261;
wire v_40262;
wire v_40263;
wire v_40264;
wire v_40265;
wire v_40266;
wire v_40267;
wire v_40268;
wire v_40269;
wire v_40270;
wire v_40271;
wire v_40272;
wire v_40273;
wire v_40274;
wire v_40275;
wire v_40276;
wire v_40277;
wire v_40278;
wire v_40279;
wire v_40280;
wire v_40281;
wire v_40282;
wire v_40283;
wire v_40284;
wire v_40285;
wire v_40286;
wire v_40287;
wire v_40288;
wire v_40289;
wire v_40290;
wire v_40291;
wire v_40292;
wire v_40293;
wire v_40294;
wire v_40295;
wire v_40296;
wire v_40297;
wire v_40298;
wire v_40299;
wire v_40300;
wire v_40301;
wire v_40302;
wire v_40303;
wire v_40304;
wire v_40305;
wire v_40306;
wire v_40307;
wire v_40308;
wire v_40309;
wire v_40310;
wire v_40311;
wire v_40312;
wire v_40313;
wire v_40314;
wire v_40315;
wire v_40317;
wire v_40318;
wire v_40319;
wire v_40320;
wire v_40321;
wire v_40322;
wire v_40323;
wire v_40324;
wire v_40325;
wire v_40326;
wire v_40327;
wire v_40328;
wire v_40329;
wire v_40330;
wire v_40331;
wire v_40332;
wire v_40333;
wire v_40334;
wire v_40335;
wire v_40336;
wire v_40337;
wire v_40338;
wire v_40339;
wire v_40340;
wire v_40341;
wire v_40342;
wire v_40343;
wire v_40344;
wire v_40345;
wire v_40346;
wire v_40347;
wire v_40348;
wire v_40349;
wire v_40350;
wire v_40351;
wire v_40352;
wire v_40353;
wire v_40354;
wire v_40355;
wire v_40356;
wire v_40357;
wire v_40358;
wire v_40359;
wire v_40360;
wire v_40361;
wire v_40362;
wire v_40363;
wire v_40364;
wire v_40365;
wire v_40366;
wire v_40367;
wire v_40368;
wire v_40369;
wire v_40370;
wire v_40371;
wire v_40372;
wire v_40373;
wire v_40374;
wire v_40375;
wire v_40376;
wire v_40377;
wire v_40378;
wire v_40379;
wire v_40380;
wire v_40381;
wire v_40382;
wire v_40383;
wire v_40384;
wire v_40385;
wire v_40386;
wire v_40387;
wire v_40388;
wire v_40389;
wire v_40390;
wire v_40391;
wire v_40392;
wire v_40393;
wire v_40394;
wire v_40395;
wire v_40396;
wire v_40397;
wire v_40398;
wire v_40399;
wire v_40400;
wire v_40401;
wire v_40402;
wire v_40403;
wire v_40404;
wire v_40405;
wire v_40406;
wire v_40407;
wire v_40408;
wire v_40409;
wire v_40410;
wire v_40411;
wire v_40412;
wire v_40413;
wire v_40414;
wire v_40415;
wire v_40416;
wire v_40417;
wire v_40418;
wire v_40419;
wire v_40420;
wire v_40421;
wire v_40422;
wire v_40423;
wire v_40424;
wire v_40425;
wire v_40426;
wire v_40427;
wire v_40428;
wire v_40429;
wire v_40430;
wire v_40431;
wire v_40432;
wire v_40433;
wire v_40434;
wire v_40435;
wire v_40436;
wire v_40437;
wire v_40438;
wire v_40439;
wire v_40440;
wire v_40441;
wire v_40442;
wire v_40443;
wire v_40444;
wire v_40445;
wire v_40446;
wire v_40447;
wire v_40448;
wire v_40449;
wire v_40450;
wire v_40451;
wire v_40452;
wire v_40453;
wire v_40454;
wire v_40455;
wire v_40456;
wire v_40457;
wire v_40458;
wire v_40459;
wire v_40460;
wire v_40461;
wire v_40462;
wire v_40463;
wire v_40464;
wire v_40465;
wire v_40466;
wire v_40467;
wire v_40468;
wire v_40469;
wire v_40470;
wire v_40471;
wire v_40472;
wire v_40473;
wire v_40474;
wire v_40475;
wire v_40476;
wire v_40477;
wire v_40478;
wire v_40479;
wire v_40480;
wire v_40481;
wire v_40482;
wire v_40483;
wire v_40484;
wire v_40485;
wire v_40486;
wire v_40487;
wire v_40488;
wire v_40489;
wire v_40490;
wire v_40491;
wire v_40492;
wire v_40493;
wire v_40494;
wire v_40495;
wire v_40496;
wire v_40497;
wire v_40498;
wire v_40499;
wire v_40500;
wire v_40501;
wire v_40502;
wire v_40503;
wire v_40504;
wire v_40505;
wire v_40506;
wire v_40507;
wire v_40508;
wire v_40509;
wire v_40510;
wire v_40511;
wire v_40512;
wire v_40513;
wire v_40514;
wire v_40515;
wire v_40516;
wire v_40517;
wire v_40518;
wire v_40519;
wire v_40520;
wire v_40521;
wire v_40522;
wire v_40523;
wire v_40524;
wire v_40525;
wire v_40526;
wire v_40527;
wire v_40528;
wire v_40529;
wire v_40530;
wire v_40531;
wire v_40532;
wire v_40533;
wire v_40534;
wire v_40535;
wire v_40536;
wire v_40537;
wire v_40538;
wire v_40539;
wire v_40540;
wire v_40541;
wire v_40542;
wire v_40543;
wire v_40544;
wire v_40545;
wire v_40546;
wire v_40547;
wire v_40548;
wire v_40549;
wire v_40550;
wire v_40551;
wire v_40552;
wire v_40553;
wire v_40554;
wire v_40555;
wire v_40556;
wire v_40557;
wire v_40558;
wire v_40560;
wire v_40561;
wire v_40562;
wire v_40563;
wire v_40564;
wire v_40565;
wire v_40566;
wire v_40567;
wire v_40568;
wire v_40569;
wire v_40570;
wire v_40571;
wire v_40572;
wire v_40573;
wire v_40574;
wire v_40575;
wire v_40576;
wire v_40577;
wire v_40578;
wire v_40579;
wire v_40580;
wire v_40581;
wire v_40582;
wire v_40583;
wire v_40584;
wire v_40585;
wire v_40586;
wire v_40587;
wire v_40588;
wire v_40589;
wire v_40590;
wire v_40591;
wire v_40592;
wire v_40593;
wire v_40594;
wire v_40595;
wire v_40596;
wire v_40597;
wire v_40598;
wire v_40599;
wire v_40600;
wire v_40601;
wire v_40602;
wire v_40603;
wire v_40604;
wire v_40605;
wire v_40606;
wire v_40607;
wire v_40608;
wire v_40609;
wire v_40610;
wire v_40611;
wire v_40612;
wire v_40613;
wire v_40614;
wire v_40615;
wire v_40616;
wire v_40617;
wire v_40618;
wire v_40619;
wire v_40620;
wire v_40621;
wire v_40622;
wire v_40623;
wire v_40624;
wire v_40625;
wire v_40626;
wire v_40627;
wire v_40628;
wire v_40629;
wire v_40630;
wire v_40631;
wire v_40632;
wire v_40633;
wire v_40634;
wire v_40635;
wire v_40636;
wire v_40637;
wire v_40638;
wire v_40639;
wire v_40640;
wire v_40641;
wire v_40642;
wire v_40643;
wire v_40644;
wire v_40645;
wire v_40646;
wire v_40647;
wire v_40648;
wire v_40649;
wire v_40650;
wire v_40651;
wire v_40652;
wire v_40653;
wire v_40654;
wire v_40655;
wire v_40656;
wire v_40657;
wire v_40658;
wire v_40659;
wire v_40660;
wire v_40661;
wire v_40662;
wire v_40663;
wire v_40664;
wire v_40665;
wire v_40666;
wire v_40667;
wire v_40668;
wire v_40669;
wire v_40670;
wire v_40671;
wire v_40672;
wire v_40673;
wire v_40674;
wire v_40675;
wire v_40676;
wire v_40677;
wire v_40678;
wire v_40679;
wire v_40680;
wire v_40681;
wire v_40682;
wire v_40683;
wire v_40684;
wire v_40685;
wire v_40686;
wire v_40687;
wire v_40688;
wire v_40689;
wire v_40690;
wire v_40691;
wire v_40692;
wire v_40693;
wire v_40694;
wire v_40695;
wire v_40696;
wire v_40697;
wire v_40698;
wire v_40699;
wire v_40700;
wire v_40701;
wire v_40702;
wire v_40703;
wire v_40704;
wire v_40705;
wire v_40706;
wire v_40707;
wire v_40708;
wire v_40709;
wire v_40710;
wire v_40711;
wire v_40712;
wire v_40713;
wire v_40714;
wire v_40715;
wire v_40716;
wire v_40717;
wire v_40718;
wire v_40719;
wire v_40720;
wire v_40721;
wire v_40722;
wire v_40723;
wire v_40724;
wire v_40725;
wire v_40726;
wire v_40727;
wire v_40728;
wire v_40729;
wire v_40730;
wire v_40731;
wire v_40732;
wire v_40733;
wire v_40734;
wire v_40735;
wire v_40736;
wire v_40737;
wire v_40738;
wire v_40739;
wire v_40740;
wire v_40741;
wire v_40742;
wire v_40743;
wire v_40744;
wire v_40745;
wire v_40746;
wire v_40747;
wire v_40748;
wire v_40749;
wire v_40750;
wire v_40751;
wire v_40752;
wire v_40753;
wire v_40754;
wire v_40755;
wire v_40756;
wire v_40757;
wire v_40758;
wire v_40759;
wire v_40760;
wire v_40761;
wire v_40762;
wire v_40763;
wire v_40764;
wire v_40765;
wire v_40766;
wire v_40767;
wire v_40768;
wire v_40769;
wire v_40770;
wire v_40771;
wire v_40772;
wire v_40773;
wire v_40774;
wire v_40775;
wire v_40776;
wire v_40777;
wire v_40778;
wire v_40779;
wire v_40780;
wire v_40781;
wire v_40782;
wire v_40783;
wire v_40784;
wire v_40785;
wire v_40786;
wire v_40787;
wire v_40788;
wire v_40789;
wire v_40790;
wire v_40791;
wire v_40792;
wire v_40793;
wire v_40794;
wire v_40795;
wire v_40796;
wire v_40797;
wire v_40798;
wire v_40799;
wire v_40800;
wire v_40801;
wire v_40803;
wire v_40804;
wire v_40805;
wire v_40806;
wire v_40807;
wire v_40808;
wire v_40809;
wire v_40810;
wire v_40811;
wire v_40812;
wire v_40813;
wire v_40814;
wire v_40815;
wire v_40816;
wire v_40817;
wire v_40818;
wire v_40819;
wire v_40820;
wire v_40821;
wire v_40822;
wire v_40823;
wire v_40824;
wire v_40825;
wire v_40826;
wire v_40827;
wire v_40828;
wire v_40829;
wire v_40830;
wire v_40831;
wire v_40832;
wire v_40833;
wire v_40834;
wire v_40835;
wire v_40836;
wire v_40837;
wire v_40838;
wire v_40839;
wire v_40840;
wire v_40841;
wire v_40842;
wire v_40843;
wire v_40844;
wire v_40845;
wire v_40846;
wire v_40847;
wire v_40848;
wire v_40849;
wire v_40850;
wire v_40851;
wire v_40852;
wire v_40853;
wire v_40854;
wire v_40855;
wire v_40856;
wire v_40857;
wire v_40858;
wire v_40859;
wire v_40860;
wire v_40861;
wire v_40862;
wire v_40863;
wire v_40864;
wire v_40865;
wire v_40866;
wire v_40867;
wire v_40868;
wire v_40869;
wire v_40870;
wire v_40871;
wire v_40872;
wire v_40873;
wire v_40874;
wire v_40875;
wire v_40876;
wire v_40877;
wire v_40878;
wire v_40879;
wire v_40880;
wire v_40881;
wire v_40882;
wire v_40883;
wire v_40884;
wire v_40885;
wire v_40886;
wire v_40887;
wire v_40888;
wire v_40889;
wire v_40890;
wire v_40891;
wire v_40892;
wire v_40893;
wire v_40894;
wire v_40895;
wire v_40896;
wire v_40897;
wire v_40898;
wire v_40899;
wire v_40900;
wire v_40901;
wire v_40902;
wire v_40903;
wire v_40904;
wire v_40905;
wire v_40906;
wire v_40907;
wire v_40908;
wire v_40909;
wire v_40910;
wire v_40911;
wire v_40912;
wire v_40913;
wire v_40914;
wire v_40915;
wire v_40916;
wire v_40917;
wire v_40918;
wire v_40919;
wire v_40920;
wire v_40921;
wire v_40922;
wire v_40923;
wire v_40924;
wire v_40925;
wire v_40926;
wire v_40927;
wire v_40928;
wire v_40929;
wire v_40930;
wire v_40931;
wire v_40932;
wire v_40933;
wire v_40934;
wire v_40935;
wire v_40936;
wire v_40937;
wire v_40938;
wire v_40939;
wire v_40940;
wire v_40941;
wire v_40942;
wire v_40943;
wire v_40944;
wire v_40945;
wire v_40946;
wire v_40947;
wire v_40948;
wire v_40949;
wire v_40950;
wire v_40951;
wire v_40952;
wire v_40953;
wire v_40954;
wire v_40955;
wire v_40956;
wire v_40957;
wire v_40958;
wire v_40959;
wire v_40960;
wire v_40961;
wire v_40962;
wire v_40963;
wire v_40964;
wire v_40965;
wire v_40966;
wire v_40967;
wire v_40968;
wire v_40969;
wire v_40970;
wire v_40971;
wire v_40972;
wire v_40973;
wire v_40974;
wire v_40975;
wire v_40976;
wire v_40977;
wire v_40978;
wire v_40979;
wire v_40980;
wire v_40981;
wire v_40982;
wire v_40983;
wire v_40984;
wire v_40985;
wire v_40986;
wire v_40987;
wire v_40988;
wire v_40989;
wire v_40990;
wire v_40991;
wire v_40992;
wire v_40993;
wire v_40994;
wire v_40995;
wire v_40996;
wire v_40997;
wire v_40998;
wire v_40999;
wire v_41000;
wire v_41001;
wire v_41002;
wire v_41003;
wire v_41004;
wire v_41005;
wire v_41006;
wire v_41007;
wire v_41008;
wire v_41009;
wire v_41010;
wire v_41011;
wire v_41012;
wire v_41013;
wire v_41014;
wire v_41015;
wire v_41016;
wire v_41017;
wire v_41018;
wire v_41019;
wire v_41020;
wire v_41021;
wire v_41022;
wire v_41023;
wire v_41024;
wire v_41025;
wire v_41026;
wire v_41027;
wire v_41028;
wire v_41029;
wire v_41030;
wire v_41031;
wire v_41032;
wire v_41033;
wire v_41034;
wire v_41035;
wire v_41036;
wire v_41037;
wire v_41038;
wire v_41039;
wire v_41040;
wire v_41041;
wire v_41042;
wire v_41043;
wire v_41044;
wire v_41046;
wire v_41047;
wire v_41048;
wire v_41049;
wire v_41050;
wire v_41051;
wire v_41052;
wire v_41053;
wire v_41054;
wire v_41055;
wire v_41056;
wire v_41057;
wire v_41058;
wire v_41059;
wire v_41060;
wire v_41061;
wire v_41062;
wire v_41063;
wire v_41064;
wire v_41065;
wire v_41066;
wire v_41067;
wire v_41068;
wire v_41069;
wire v_41070;
wire v_41071;
wire v_41072;
wire v_41073;
wire v_41074;
wire v_41075;
wire v_41076;
wire v_41077;
wire v_41078;
wire v_41079;
wire v_41080;
wire v_41081;
wire v_41082;
wire v_41083;
wire v_41084;
wire v_41085;
wire v_41086;
wire v_41087;
wire v_41088;
wire v_41089;
wire v_41090;
wire v_41091;
wire v_41092;
wire v_41093;
wire v_41094;
wire v_41095;
wire v_41096;
wire v_41097;
wire v_41098;
wire v_41099;
wire v_41100;
wire v_41101;
wire v_41102;
wire v_41103;
wire v_41104;
wire v_41105;
wire v_41106;
wire v_41107;
wire v_41108;
wire v_41109;
wire v_41110;
wire v_41111;
wire v_41112;
wire v_41113;
wire v_41114;
wire v_41115;
wire v_41116;
wire v_41117;
wire v_41118;
wire v_41119;
wire v_41120;
wire v_41121;
wire v_41122;
wire v_41123;
wire v_41124;
wire v_41125;
wire v_41126;
wire v_41127;
wire v_41128;
wire v_41129;
wire v_41130;
wire v_41131;
wire v_41132;
wire v_41133;
wire v_41134;
wire v_41135;
wire v_41136;
wire v_41137;
wire v_41138;
wire v_41139;
wire v_41140;
wire v_41141;
wire v_41142;
wire v_41143;
wire v_41144;
wire v_41145;
wire v_41146;
wire v_41147;
wire v_41148;
wire v_41149;
wire v_41150;
wire v_41151;
wire v_41152;
wire v_41153;
wire v_41154;
wire v_41155;
wire v_41156;
wire v_41157;
wire v_41158;
wire v_41159;
wire v_41160;
wire v_41161;
wire v_41162;
wire v_41163;
wire v_41164;
wire v_41165;
wire v_41166;
wire v_41167;
wire v_41168;
wire v_41169;
wire v_41170;
wire v_41171;
wire v_41172;
wire v_41173;
wire v_41174;
wire v_41175;
wire v_41176;
wire v_41177;
wire v_41178;
wire v_41179;
wire v_41180;
wire v_41181;
wire v_41182;
wire v_41183;
wire v_41184;
wire v_41185;
wire v_41186;
wire v_41187;
wire v_41188;
wire v_41189;
wire v_41190;
wire v_41191;
wire v_41192;
wire v_41193;
wire v_41194;
wire v_41195;
wire v_41196;
wire v_41197;
wire v_41198;
wire v_41199;
wire v_41200;
wire v_41201;
wire v_41202;
wire v_41203;
wire v_41204;
wire v_41205;
wire v_41206;
wire v_41207;
wire v_41208;
wire v_41209;
wire v_41210;
wire v_41211;
wire v_41212;
wire v_41213;
wire v_41214;
wire v_41215;
wire v_41216;
wire v_41217;
wire v_41218;
wire v_41219;
wire v_41220;
wire v_41221;
wire v_41222;
wire v_41223;
wire v_41224;
wire v_41225;
wire v_41226;
wire v_41227;
wire v_41228;
wire v_41229;
wire v_41230;
wire v_41231;
wire v_41232;
wire v_41233;
wire v_41234;
wire v_41235;
wire v_41236;
wire v_41237;
wire v_41238;
wire v_41239;
wire v_41240;
wire v_41241;
wire v_41242;
wire v_41243;
wire v_41244;
wire v_41245;
wire v_41246;
wire v_41247;
wire v_41248;
wire v_41249;
wire v_41250;
wire v_41251;
wire v_41252;
wire v_41253;
wire v_41254;
wire v_41255;
wire v_41256;
wire v_41257;
wire v_41258;
wire v_41259;
wire v_41260;
wire v_41261;
wire v_41262;
wire v_41263;
wire v_41264;
wire v_41265;
wire v_41266;
wire v_41267;
wire v_41268;
wire v_41269;
wire v_41270;
wire v_41271;
wire v_41272;
wire v_41273;
wire v_41274;
wire v_41275;
wire v_41276;
wire v_41277;
wire v_41278;
wire v_41279;
wire v_41280;
wire v_41281;
wire v_41282;
wire v_41283;
wire v_41284;
wire v_41285;
wire v_41286;
wire v_41287;
wire v_41289;
wire v_41290;
wire v_41291;
wire v_41292;
wire v_41293;
wire v_41294;
wire v_41295;
wire v_41296;
wire v_41297;
wire v_41298;
wire v_41299;
wire v_41300;
wire v_41301;
wire v_41302;
wire v_41303;
wire v_41304;
wire v_41305;
wire v_41306;
wire v_41307;
wire v_41308;
wire v_41309;
wire v_41310;
wire v_41311;
wire v_41312;
wire v_41313;
wire v_41314;
wire v_41315;
wire v_41316;
wire v_41317;
wire v_41318;
wire v_41319;
wire v_41320;
wire v_41321;
wire v_41322;
wire v_41323;
wire v_41324;
wire v_41325;
wire v_41326;
wire v_41327;
wire v_41328;
wire v_41329;
wire v_41330;
wire v_41331;
wire v_41332;
wire v_41333;
wire v_41334;
wire v_41335;
wire v_41336;
wire v_41337;
wire v_41338;
wire v_41339;
wire v_41340;
wire v_41341;
wire v_41342;
wire v_41343;
wire v_41344;
wire v_41345;
wire v_41346;
wire v_41347;
wire v_41348;
wire v_41349;
wire v_41350;
wire v_41351;
wire v_41352;
wire v_41353;
wire v_41354;
wire v_41355;
wire v_41356;
wire v_41357;
wire v_41358;
wire v_41359;
wire v_41360;
wire v_41361;
wire v_41362;
wire v_41363;
wire v_41364;
wire v_41365;
wire v_41366;
wire v_41367;
wire v_41368;
wire v_41369;
wire v_41370;
wire v_41371;
wire v_41372;
wire v_41373;
wire v_41374;
wire v_41375;
wire v_41376;
wire v_41377;
wire v_41378;
wire v_41379;
wire v_41380;
wire v_41381;
wire v_41382;
wire v_41383;
wire v_41384;
wire v_41385;
wire v_41386;
wire v_41387;
wire v_41388;
wire v_41389;
wire v_41390;
wire v_41391;
wire v_41392;
wire v_41393;
wire v_41394;
wire v_41395;
wire v_41396;
wire v_41397;
wire v_41398;
wire v_41399;
wire v_41400;
wire v_41401;
wire v_41402;
wire v_41403;
wire v_41404;
wire v_41405;
wire v_41406;
wire v_41407;
wire v_41408;
wire v_41409;
wire v_41410;
wire v_41411;
wire v_41412;
wire v_41413;
wire v_41414;
wire v_41415;
wire v_41416;
wire v_41417;
wire v_41418;
wire v_41419;
wire v_41420;
wire v_41421;
wire v_41422;
wire v_41423;
wire v_41424;
wire v_41425;
wire v_41426;
wire v_41427;
wire v_41428;
wire v_41429;
wire v_41430;
wire v_41431;
wire v_41432;
wire v_41433;
wire v_41434;
wire v_41435;
wire v_41436;
wire v_41437;
wire v_41438;
wire v_41439;
wire v_41440;
wire v_41441;
wire v_41442;
wire v_41443;
wire v_41444;
wire v_41445;
wire v_41446;
wire v_41447;
wire v_41448;
wire v_41449;
wire v_41450;
wire v_41451;
wire v_41452;
wire v_41453;
wire v_41454;
wire v_41455;
wire v_41456;
wire v_41457;
wire v_41458;
wire v_41459;
wire v_41460;
wire v_41461;
wire v_41462;
wire v_41463;
wire v_41464;
wire v_41465;
wire v_41466;
wire v_41467;
wire v_41468;
wire v_41469;
wire v_41470;
wire v_41471;
wire v_41472;
wire v_41473;
wire v_41474;
wire v_41475;
wire v_41476;
wire v_41477;
wire v_41478;
wire v_41479;
wire v_41480;
wire v_41481;
wire v_41482;
wire v_41483;
wire v_41484;
wire v_41485;
wire v_41486;
wire v_41487;
wire v_41488;
wire v_41489;
wire v_41490;
wire v_41491;
wire v_41492;
wire v_41493;
wire v_41494;
wire v_41495;
wire v_41496;
wire v_41497;
wire v_41498;
wire v_41499;
wire v_41500;
wire v_41501;
wire v_41502;
wire v_41503;
wire v_41504;
wire v_41505;
wire v_41506;
wire v_41507;
wire v_41508;
wire v_41509;
wire v_41510;
wire v_41511;
wire v_41512;
wire v_41513;
wire v_41514;
wire v_41515;
wire v_41516;
wire v_41517;
wire v_41518;
wire v_41519;
wire v_41520;
wire v_41521;
wire v_41522;
wire v_41523;
wire v_41524;
wire v_41525;
wire v_41526;
wire v_41527;
wire v_41528;
wire v_41529;
wire v_41530;
wire v_41531;
wire v_41532;
wire v_41533;
wire v_41534;
wire v_41535;
wire v_41536;
wire v_41537;
wire v_41538;
wire v_41539;
wire v_41540;
wire v_41541;
wire v_41542;
wire v_41543;
wire v_41544;
wire v_41545;
wire v_41546;
wire v_41547;
wire v_41548;
wire v_41549;
wire v_41550;
wire v_41551;
wire v_41552;
wire v_41553;
wire v_41554;
wire v_41555;
wire v_41556;
wire v_41557;
wire v_41558;
wire v_41559;
wire v_41560;
wire v_41561;
wire v_41562;
wire v_41563;
wire v_41564;
wire v_41565;
wire v_41566;
wire v_41567;
wire v_41568;
wire v_41569;
wire v_41570;
wire v_41571;
wire v_41572;
wire v_41573;
wire v_41574;
wire v_41575;
wire v_41576;
wire v_41577;
wire v_41578;
wire v_41579;
wire v_41580;
wire v_41581;
wire v_41582;
wire v_41583;
wire v_41584;
wire v_41585;
wire v_41586;
wire v_41587;
wire v_41588;
wire v_41589;
wire v_41590;
wire v_41591;
wire v_41592;
wire v_41593;
wire v_41594;
wire v_41595;
wire v_41596;
wire v_41597;
wire v_41598;
wire v_41599;
wire v_41600;
wire v_41601;
wire v_41602;
wire v_41603;
wire v_41604;
wire v_41605;
wire v_41606;
wire v_41607;
wire v_41608;
wire v_41609;
wire v_41610;
wire v_41611;
wire v_41612;
wire v_41613;
wire v_41614;
wire v_41615;
wire v_41616;
wire v_41617;
wire v_41618;
wire v_41619;
wire v_41620;
wire v_41621;
wire v_41622;
wire v_41623;
wire v_41624;
wire v_41625;
wire v_41626;
wire v_41627;
wire v_41628;
wire v_41629;
wire v_41630;
wire v_41631;
wire v_41632;
wire v_41633;
wire v_41634;
wire v_41635;
wire v_41636;
wire v_41637;
wire v_41638;
wire v_41639;
wire v_41640;
wire v_41641;
wire v_41642;
wire v_41643;
wire v_41644;
wire v_41645;
wire v_41646;
wire v_41647;
wire v_41648;
wire v_41649;
wire v_41650;
wire v_41651;
wire v_41652;
wire v_41653;
wire v_41654;
wire v_41655;
wire v_41656;
wire v_41657;
wire v_41658;
wire v_41659;
wire v_41660;
wire v_41661;
wire v_41662;
wire v_41663;
wire v_41664;
wire v_41665;
wire v_41666;
wire v_41667;
wire v_41668;
wire v_41669;
wire v_41670;
wire v_41671;
wire v_41672;
wire v_41673;
wire v_41674;
wire v_41675;
wire v_41676;
wire v_41677;
wire v_41678;
wire v_41679;
wire v_41681;
wire v_41682;
wire v_41683;
wire v_41684;
wire v_41685;
wire v_41686;
wire v_41687;
wire v_41688;
wire v_41689;
wire v_41690;
wire v_41691;
wire v_41692;
wire v_41693;
wire v_41694;
wire v_41695;
wire v_41696;
wire v_41697;
wire v_41698;
wire v_41699;
wire v_41700;
wire v_41701;
wire v_41702;
wire v_41703;
wire v_41704;
wire v_41705;
wire v_41706;
wire v_41707;
wire v_41708;
wire v_41709;
wire v_41710;
wire v_41711;
wire v_41712;
wire v_41713;
wire v_41714;
wire v_41715;
wire v_41716;
wire v_41717;
wire v_41718;
wire v_41719;
wire v_41720;
wire v_41721;
wire v_41722;
wire v_41723;
wire v_41724;
wire v_41725;
wire v_41726;
wire v_41727;
wire v_41728;
wire v_41729;
wire v_41730;
wire v_41731;
wire v_41732;
wire v_41733;
wire v_41734;
wire v_41735;
wire v_41736;
wire v_41737;
wire v_41738;
wire v_41739;
wire v_41740;
wire v_41741;
wire v_41742;
wire v_41743;
wire v_41744;
wire v_41745;
wire v_41746;
wire v_41747;
wire v_41748;
wire v_41749;
wire v_41750;
wire v_41751;
wire v_41752;
wire v_41753;
wire v_41754;
wire v_41755;
wire v_41756;
wire v_41757;
wire v_41758;
wire v_41759;
wire v_41760;
wire v_41761;
wire v_41762;
wire v_41763;
wire v_41764;
wire v_41765;
wire v_41766;
wire v_41767;
wire v_41768;
wire v_41769;
wire v_41770;
wire v_41771;
wire v_41772;
wire v_41773;
wire v_41775;
wire v_41777;
wire v_41778;
wire v_41779;
wire v_41781;
wire v_41782;
wire v_41783;
wire v_41785;
wire v_41786;
wire v_41787;
wire v_41789;
wire v_41790;
wire v_41792;
wire v_41793;
wire v_41794;
wire v_41796;
wire v_41797;
wire v_41798;
wire v_41800;
wire v_41801;
wire v_41802;
wire v_41804;
wire v_41805;
wire v_41806;
wire v_41808;
wire v_41809;
wire v_41810;
wire v_41812;
wire v_41813;
wire v_41814;
wire v_41816;
wire v_41817;
wire v_41818;
wire v_41820;
wire v_41821;
wire v_41822;
wire v_41824;
wire v_41825;
wire v_41826;
wire v_41828;
wire v_41829;
wire v_41830;
wire v_41832;
wire v_41833;
wire v_41834;
wire v_41836;
wire v_41837;
wire v_41838;
wire v_41840;
wire v_41841;
wire v_41842;
wire v_41843;
wire v_41844;
wire v_41845;
wire v_41846;
wire v_41847;
wire v_41848;
wire v_41849;
wire v_41850;
wire v_41851;
wire v_41852;
wire v_41853;
wire v_41854;
wire v_41855;
wire v_41856;
wire v_41857;
wire v_41858;
wire v_41859;
wire v_41860;
wire v_41861;
wire v_41862;
wire v_41863;
wire v_41864;
wire v_41865;
wire v_41866;
wire v_41867;
wire v_41868;
wire v_41869;
wire v_41870;
wire v_41871;
wire v_41872;
wire v_41873;
wire v_41874;
wire v_41875;
wire v_41876;
wire v_41877;
wire v_41878;
wire v_41879;
wire v_41880;
wire v_41881;
wire v_41882;
wire v_41883;
wire v_41884;
wire v_41885;
wire v_41886;
wire v_41887;
wire v_41888;
wire v_41889;
wire v_41890;
wire v_41891;
wire v_41892;
wire v_41893;
wire v_41894;
wire v_41895;
wire v_41896;
wire v_41897;
wire v_41898;
wire v_41899;
wire v_41900;
wire v_41901;
wire v_41902;
wire v_41903;
wire v_41904;
wire v_41905;
wire v_41906;
wire v_41907;
wire v_41908;
wire v_41909;
wire v_41910;
wire v_41911;
wire v_41912;
wire v_41913;
wire v_41914;
wire v_41915;
wire v_41916;
wire v_41917;
wire v_41918;
wire v_41919;
wire v_41920;
wire v_41921;
wire v_41922;
wire v_41923;
wire v_41924;
wire v_41925;
wire v_41926;
wire v_41927;
wire v_41928;
wire v_41929;
wire v_41930;
wire v_41931;
wire v_41932;
wire v_41933;
wire v_41934;
wire v_41935;
wire v_41936;
wire v_41937;
wire v_41938;
wire v_41939;
wire v_41940;
wire v_41941;
wire v_41942;
wire v_41943;
wire v_41944;
wire v_41945;
wire v_41946;
wire v_41947;
wire v_41948;
wire v_41949;
wire v_41950;
wire v_41951;
wire v_41952;
wire v_41953;
wire v_41954;
wire v_41955;
wire v_41956;
wire v_41957;
wire v_41958;
wire v_41959;
wire v_41960;
wire v_41961;
wire v_41962;
wire v_41963;
wire v_41964;
wire v_41965;
wire v_41966;
wire v_41967;
wire v_41968;
wire v_41969;
wire v_41970;
wire v_41971;
wire v_41972;
wire v_41973;
wire v_41974;
wire v_41975;
wire v_41976;
wire v_41977;
wire v_41978;
wire v_41979;
wire v_41980;
wire v_41981;
wire v_41982;
wire v_41983;
wire v_41984;
wire v_41985;
wire v_41986;
wire v_41987;
wire v_41988;
wire v_41989;
wire v_41990;
wire v_41991;
wire v_41992;
wire v_41993;
wire v_41994;
wire v_41995;
wire v_41996;
wire v_41997;
wire v_41998;
wire v_41999;
wire v_42000;
wire v_42001;
wire v_42002;
wire v_42003;
wire v_42004;
wire v_42005;
wire v_42006;
wire v_42007;
wire v_42008;
wire v_42009;
wire v_42010;
wire v_42011;
wire v_42012;
wire v_42013;
wire v_42014;
wire v_42015;
wire v_42016;
wire v_42017;
wire v_42018;
wire v_42019;
wire v_42020;
wire v_42021;
wire v_42022;
wire v_42023;
wire v_42024;
wire v_42025;
wire v_42026;
wire v_42027;
wire v_42028;
wire v_42029;
wire v_42030;
wire v_42031;
wire v_42032;
wire v_42033;
wire v_42035;
wire v_42036;
wire v_42037;
wire v_42038;
wire v_42039;
wire v_42040;
wire v_42041;
wire v_42042;
wire v_42043;
wire v_42044;
wire v_42045;
wire v_42046;
wire v_42047;
wire v_42048;
wire v_42049;
wire v_42050;
wire v_42051;
wire v_42052;
wire v_42053;
wire v_42054;
wire v_42055;
wire v_42056;
wire v_42057;
wire v_42058;
wire v_42059;
wire v_42060;
wire v_42061;
wire v_42062;
wire v_42063;
wire v_42064;
wire v_42065;
wire v_42066;
wire v_42067;
wire v_42068;
wire v_42069;
wire v_42070;
wire v_42071;
wire v_42072;
wire v_42073;
wire v_42074;
wire v_42075;
wire v_42076;
wire v_42077;
wire v_42078;
wire v_42079;
wire v_42080;
wire v_42081;
wire v_42082;
wire v_42083;
wire v_42084;
wire v_42085;
wire v_42086;
wire v_42087;
wire v_42088;
wire v_42089;
wire v_42090;
wire v_42091;
wire v_42092;
wire v_42093;
wire v_42094;
wire v_42095;
wire v_42096;
wire v_42097;
wire v_42098;
wire v_42099;
wire v_42100;
wire v_42101;
wire v_42102;
wire v_42103;
wire v_42104;
wire v_42105;
wire v_42106;
wire v_42107;
wire v_42108;
wire v_42109;
wire v_42110;
wire v_42111;
wire v_42112;
wire v_42113;
wire v_42114;
wire v_42115;
wire v_42116;
wire v_42117;
wire v_42118;
wire v_42119;
wire v_42120;
wire v_42121;
wire v_42122;
wire v_42123;
wire v_42124;
wire v_42125;
wire v_42126;
wire v_42127;
wire v_42128;
wire v_42129;
wire v_42130;
wire v_42131;
wire v_42132;
wire v_42133;
wire v_42134;
wire v_42135;
wire v_42136;
wire v_42137;
wire v_42138;
wire v_42139;
wire v_42140;
wire v_42141;
wire v_42142;
wire v_42143;
wire v_42144;
wire v_42145;
wire v_42146;
wire v_42147;
wire v_42148;
wire v_42149;
wire v_42150;
wire v_42151;
wire v_42152;
wire v_42153;
wire v_42154;
wire v_42155;
wire v_42156;
wire v_42157;
wire v_42158;
wire v_42159;
wire v_42160;
wire v_42161;
wire v_42162;
wire v_42163;
wire v_42164;
wire v_42165;
wire v_42166;
wire v_42167;
wire v_42168;
wire v_42169;
wire v_42170;
wire v_42171;
wire v_42172;
wire v_42173;
wire v_42174;
wire v_42175;
wire v_42176;
wire v_42177;
wire v_42178;
wire v_42179;
wire v_42180;
wire v_42181;
wire v_42182;
wire v_42183;
wire v_42184;
wire v_42185;
wire v_42186;
wire v_42187;
wire v_42188;
wire v_42189;
wire v_42190;
wire v_42191;
wire v_42192;
wire v_42193;
wire v_42194;
wire v_42195;
wire v_42196;
wire v_42197;
wire v_42198;
wire v_42199;
wire v_42200;
wire v_42201;
wire v_42202;
wire v_42203;
wire v_42204;
wire v_42205;
wire v_42206;
wire v_42207;
wire v_42208;
wire v_42209;
wire v_42210;
wire v_42211;
wire v_42212;
wire v_42213;
wire v_42214;
wire v_42215;
wire v_42216;
wire v_42217;
wire v_42218;
wire v_42219;
wire v_42220;
wire v_42221;
wire v_42222;
wire v_42223;
wire v_42224;
wire v_42225;
wire v_42226;
wire v_42227;
wire v_42228;
wire v_42229;
wire v_42230;
wire v_42231;
wire v_42232;
wire v_42233;
wire v_42234;
wire v_42235;
wire v_42236;
wire v_42237;
wire v_42238;
wire v_42239;
wire v_42240;
wire v_42241;
wire v_42242;
wire v_42243;
wire v_42244;
wire v_42245;
wire v_42246;
wire v_42247;
wire v_42248;
wire v_42249;
wire v_42250;
wire v_42251;
wire v_42252;
wire v_42253;
wire v_42254;
wire v_42255;
wire v_42256;
wire v_42257;
wire v_42258;
wire v_42259;
wire v_42260;
wire v_42261;
wire v_42262;
wire v_42263;
wire v_42264;
wire v_42265;
wire v_42266;
wire v_42267;
wire v_42268;
wire v_42269;
wire v_42270;
wire v_42271;
wire v_42272;
wire v_42273;
wire v_42274;
wire v_42275;
wire v_42276;
wire v_42278;
wire v_42279;
wire v_42280;
wire v_42281;
wire v_42282;
wire v_42283;
wire v_42284;
wire v_42285;
wire v_42286;
wire v_42287;
wire v_42288;
wire v_42289;
wire v_42290;
wire v_42291;
wire v_42292;
wire v_42293;
wire v_42294;
wire v_42295;
wire v_42296;
wire v_42297;
wire v_42298;
wire v_42299;
wire v_42300;
wire v_42301;
wire v_42302;
wire v_42303;
wire v_42304;
wire v_42305;
wire v_42306;
wire v_42307;
wire v_42308;
wire v_42309;
wire v_42310;
wire v_42311;
wire v_42312;
wire v_42313;
wire v_42314;
wire v_42315;
wire v_42316;
wire v_42317;
wire v_42318;
wire v_42319;
wire v_42320;
wire v_42321;
wire v_42322;
wire v_42323;
wire v_42324;
wire v_42325;
wire v_42326;
wire v_42327;
wire v_42328;
wire v_42329;
wire v_42330;
wire v_42331;
wire v_42332;
wire v_42333;
wire v_42334;
wire v_42335;
wire v_42336;
wire v_42337;
wire v_42338;
wire v_42339;
wire v_42340;
wire v_42341;
wire v_42342;
wire v_42343;
wire v_42344;
wire v_42345;
wire v_42346;
wire v_42347;
wire v_42348;
wire v_42349;
wire v_42350;
wire v_42351;
wire v_42352;
wire v_42353;
wire v_42354;
wire v_42355;
wire v_42356;
wire v_42357;
wire v_42358;
wire v_42359;
wire v_42360;
wire v_42361;
wire v_42362;
wire v_42363;
wire v_42364;
wire v_42365;
wire v_42366;
wire v_42367;
wire v_42368;
wire v_42369;
wire v_42370;
wire v_42371;
wire v_42372;
wire v_42373;
wire v_42374;
wire v_42375;
wire v_42376;
wire v_42377;
wire v_42378;
wire v_42379;
wire v_42380;
wire v_42381;
wire v_42382;
wire v_42383;
wire v_42384;
wire v_42385;
wire v_42386;
wire v_42387;
wire v_42388;
wire v_42389;
wire v_42390;
wire v_42391;
wire v_42392;
wire v_42393;
wire v_42394;
wire v_42395;
wire v_42396;
wire v_42397;
wire v_42398;
wire v_42399;
wire v_42400;
wire v_42401;
wire v_42402;
wire v_42403;
wire v_42404;
wire v_42405;
wire v_42406;
wire v_42407;
wire v_42408;
wire v_42409;
wire v_42410;
wire v_42411;
wire v_42412;
wire v_42413;
wire v_42414;
wire v_42415;
wire v_42416;
wire v_42417;
wire v_42418;
wire v_42419;
wire v_42420;
wire v_42421;
wire v_42422;
wire v_42423;
wire v_42424;
wire v_42425;
wire v_42426;
wire v_42427;
wire v_42428;
wire v_42429;
wire v_42430;
wire v_42431;
wire v_42432;
wire v_42433;
wire v_42434;
wire v_42435;
wire v_42436;
wire v_42437;
wire v_42438;
wire v_42439;
wire v_42440;
wire v_42441;
wire v_42442;
wire v_42443;
wire v_42444;
wire v_42445;
wire v_42446;
wire v_42447;
wire v_42448;
wire v_42449;
wire v_42450;
wire v_42451;
wire v_42452;
wire v_42453;
wire v_42454;
wire v_42455;
wire v_42456;
wire v_42457;
wire v_42458;
wire v_42459;
wire v_42460;
wire v_42461;
wire v_42462;
wire v_42463;
wire v_42464;
wire v_42465;
wire v_42466;
wire v_42467;
wire v_42468;
wire v_42469;
wire v_42470;
wire v_42471;
wire v_42472;
wire v_42473;
wire v_42474;
wire v_42475;
wire v_42476;
wire v_42477;
wire v_42478;
wire v_42479;
wire v_42480;
wire v_42481;
wire v_42482;
wire v_42483;
wire v_42484;
wire v_42485;
wire v_42486;
wire v_42487;
wire v_42488;
wire v_42489;
wire v_42490;
wire v_42491;
wire v_42492;
wire v_42493;
wire v_42494;
wire v_42495;
wire v_42496;
wire v_42497;
wire v_42498;
wire v_42499;
wire v_42500;
wire v_42501;
wire v_42502;
wire v_42503;
wire v_42504;
wire v_42505;
wire v_42506;
wire v_42507;
wire v_42508;
wire v_42509;
wire v_42510;
wire v_42511;
wire v_42512;
wire v_42513;
wire v_42514;
wire v_42515;
wire v_42516;
wire v_42517;
wire v_42518;
wire v_42519;
wire v_42521;
wire v_42522;
wire v_42523;
wire v_42524;
wire v_42525;
wire v_42526;
wire v_42527;
wire v_42528;
wire v_42529;
wire v_42530;
wire v_42531;
wire v_42532;
wire v_42533;
wire v_42534;
wire v_42535;
wire v_42536;
wire v_42537;
wire v_42538;
wire v_42539;
wire v_42540;
wire v_42541;
wire v_42542;
wire v_42543;
wire v_42544;
wire v_42545;
wire v_42546;
wire v_42547;
wire v_42548;
wire v_42549;
wire v_42550;
wire v_42551;
wire v_42552;
wire v_42553;
wire v_42554;
wire v_42555;
wire v_42556;
wire v_42557;
wire v_42558;
wire v_42559;
wire v_42560;
wire v_42561;
wire v_42562;
wire v_42563;
wire v_42564;
wire v_42565;
wire v_42566;
wire v_42567;
wire v_42568;
wire v_42569;
wire v_42570;
wire v_42571;
wire v_42572;
wire v_42573;
wire v_42574;
wire v_42575;
wire v_42576;
wire v_42577;
wire v_42578;
wire v_42579;
wire v_42580;
wire v_42581;
wire v_42582;
wire v_42583;
wire v_42584;
wire v_42585;
wire v_42586;
wire v_42587;
wire v_42588;
wire v_42589;
wire v_42590;
wire v_42591;
wire v_42592;
wire v_42593;
wire v_42594;
wire v_42595;
wire v_42596;
wire v_42597;
wire v_42598;
wire v_42599;
wire v_42600;
wire v_42601;
wire v_42602;
wire v_42603;
wire v_42604;
wire v_42605;
wire v_42606;
wire v_42607;
wire v_42608;
wire v_42609;
wire v_42610;
wire v_42611;
wire v_42612;
wire v_42613;
wire v_42614;
wire v_42615;
wire v_42616;
wire v_42617;
wire v_42618;
wire v_42619;
wire v_42620;
wire v_42621;
wire v_42622;
wire v_42623;
wire v_42624;
wire v_42625;
wire v_42626;
wire v_42627;
wire v_42628;
wire v_42629;
wire v_42630;
wire v_42631;
wire v_42632;
wire v_42633;
wire v_42634;
wire v_42635;
wire v_42636;
wire v_42637;
wire v_42638;
wire v_42639;
wire v_42640;
wire v_42641;
wire v_42642;
wire v_42643;
wire v_42644;
wire v_42645;
wire v_42646;
wire v_42647;
wire v_42648;
wire v_42649;
wire v_42650;
wire v_42651;
wire v_42652;
wire v_42653;
wire v_42654;
wire v_42655;
wire v_42656;
wire v_42657;
wire v_42658;
wire v_42659;
wire v_42660;
wire v_42661;
wire v_42662;
wire v_42663;
wire v_42664;
wire v_42665;
wire v_42666;
wire v_42667;
wire v_42668;
wire v_42669;
wire v_42670;
wire v_42671;
wire v_42672;
wire v_42673;
wire v_42674;
wire v_42675;
wire v_42676;
wire v_42677;
wire v_42678;
wire v_42679;
wire v_42680;
wire v_42681;
wire v_42682;
wire v_42683;
wire v_42684;
wire v_42685;
wire v_42686;
wire v_42687;
wire v_42688;
wire v_42689;
wire v_42690;
wire v_42691;
wire v_42692;
wire v_42693;
wire v_42694;
wire v_42695;
wire v_42696;
wire v_42697;
wire v_42698;
wire v_42699;
wire v_42700;
wire v_42701;
wire v_42702;
wire v_42703;
wire v_42704;
wire v_42705;
wire v_42706;
wire v_42707;
wire v_42708;
wire v_42709;
wire v_42710;
wire v_42711;
wire v_42712;
wire v_42713;
wire v_42714;
wire v_42715;
wire v_42716;
wire v_42717;
wire v_42718;
wire v_42719;
wire v_42720;
wire v_42721;
wire v_42722;
wire v_42723;
wire v_42724;
wire v_42725;
wire v_42726;
wire v_42727;
wire v_42728;
wire v_42729;
wire v_42730;
wire v_42731;
wire v_42732;
wire v_42733;
wire v_42734;
wire v_42735;
wire v_42736;
wire v_42737;
wire v_42738;
wire v_42739;
wire v_42740;
wire v_42741;
wire v_42742;
wire v_42743;
wire v_42744;
wire v_42745;
wire v_42746;
wire v_42747;
wire v_42748;
wire v_42749;
wire v_42750;
wire v_42751;
wire v_42752;
wire v_42753;
wire v_42754;
wire v_42755;
wire v_42756;
wire v_42757;
wire v_42758;
wire v_42759;
wire v_42760;
wire v_42761;
wire v_42762;
wire v_42764;
wire v_42765;
wire v_42766;
wire v_42767;
wire v_42768;
wire v_42769;
wire v_42770;
wire v_42771;
wire v_42772;
wire v_42773;
wire v_42774;
wire v_42775;
wire v_42776;
wire v_42777;
wire v_42778;
wire v_42779;
wire v_42780;
wire v_42781;
wire v_42782;
wire v_42783;
wire v_42784;
wire v_42785;
wire v_42786;
wire v_42787;
wire v_42788;
wire v_42789;
wire v_42790;
wire v_42791;
wire v_42792;
wire v_42793;
wire v_42794;
wire v_42795;
wire v_42796;
wire v_42797;
wire v_42798;
wire v_42799;
wire v_42800;
wire v_42801;
wire v_42802;
wire v_42803;
wire v_42804;
wire v_42805;
wire v_42806;
wire v_42807;
wire v_42808;
wire v_42809;
wire v_42810;
wire v_42811;
wire v_42812;
wire v_42813;
wire v_42814;
wire v_42815;
wire v_42816;
wire v_42817;
wire v_42818;
wire v_42819;
wire v_42820;
wire v_42821;
wire v_42822;
wire v_42823;
wire v_42824;
wire v_42825;
wire v_42826;
wire v_42827;
wire v_42828;
wire v_42829;
wire v_42830;
wire v_42831;
wire v_42832;
wire v_42833;
wire v_42834;
wire v_42835;
wire v_42836;
wire v_42837;
wire v_42838;
wire v_42839;
wire v_42840;
wire v_42841;
wire v_42842;
wire v_42843;
wire v_42844;
wire v_42845;
wire v_42846;
wire v_42847;
wire v_42848;
wire v_42849;
wire v_42850;
wire v_42851;
wire v_42852;
wire v_42853;
wire v_42854;
wire v_42855;
wire v_42856;
wire v_42857;
wire v_42858;
wire v_42859;
wire v_42860;
wire v_42861;
wire v_42862;
wire v_42863;
wire v_42864;
wire v_42865;
wire v_42866;
wire v_42867;
wire v_42868;
wire v_42869;
wire v_42870;
wire v_42871;
wire v_42872;
wire v_42873;
wire v_42874;
wire v_42875;
wire v_42876;
wire v_42877;
wire v_42878;
wire v_42879;
wire v_42880;
wire v_42881;
wire v_42882;
wire v_42883;
wire v_42884;
wire v_42885;
wire v_42886;
wire v_42887;
wire v_42888;
wire v_42889;
wire v_42890;
wire v_42891;
wire v_42892;
wire v_42893;
wire v_42894;
wire v_42895;
wire v_42896;
wire v_42897;
wire v_42898;
wire v_42899;
wire v_42900;
wire v_42901;
wire v_42902;
wire v_42903;
wire v_42904;
wire v_42905;
wire v_42906;
wire v_42907;
wire v_42908;
wire v_42909;
wire v_42910;
wire v_42911;
wire v_42912;
wire v_42913;
wire v_42914;
wire v_42915;
wire v_42916;
wire v_42917;
wire v_42918;
wire v_42919;
wire v_42920;
wire v_42921;
wire v_42922;
wire v_42923;
wire v_42924;
wire v_42925;
wire v_42926;
wire v_42927;
wire v_42928;
wire v_42929;
wire v_42930;
wire v_42931;
wire v_42932;
wire v_42933;
wire v_42934;
wire v_42935;
wire v_42936;
wire v_42937;
wire v_42938;
wire v_42939;
wire v_42940;
wire v_42941;
wire v_42942;
wire v_42943;
wire v_42944;
wire v_42945;
wire v_42946;
wire v_42947;
wire v_42948;
wire v_42949;
wire v_42950;
wire v_42951;
wire v_42952;
wire v_42953;
wire v_42954;
wire v_42955;
wire v_42956;
wire v_42957;
wire v_42958;
wire v_42959;
wire v_42960;
wire v_42961;
wire v_42962;
wire v_42963;
wire v_42964;
wire v_42965;
wire v_42966;
wire v_42967;
wire v_42968;
wire v_42969;
wire v_42970;
wire v_42971;
wire v_42972;
wire v_42973;
wire v_42974;
wire v_42975;
wire v_42976;
wire v_42977;
wire v_42978;
wire v_42979;
wire v_42980;
wire v_42981;
wire v_42982;
wire v_42983;
wire v_42984;
wire v_42985;
wire v_42986;
wire v_42987;
wire v_42988;
wire v_42989;
wire v_42990;
wire v_42991;
wire v_42992;
wire v_42993;
wire v_42994;
wire v_42995;
wire v_42996;
wire v_42997;
wire v_42998;
wire v_42999;
wire v_43000;
wire v_43001;
wire v_43002;
wire v_43003;
wire v_43004;
wire v_43005;
wire v_43007;
wire v_43008;
wire v_43009;
wire v_43010;
wire v_43011;
wire v_43012;
wire v_43013;
wire v_43014;
wire v_43015;
wire v_43016;
wire v_43017;
wire v_43018;
wire v_43019;
wire v_43020;
wire v_43021;
wire v_43022;
wire v_43023;
wire v_43024;
wire v_43025;
wire v_43026;
wire v_43027;
wire v_43028;
wire v_43029;
wire v_43030;
wire v_43031;
wire v_43032;
wire v_43033;
wire v_43034;
wire v_43035;
wire v_43036;
wire v_43037;
wire v_43038;
wire v_43039;
wire v_43040;
wire v_43041;
wire v_43042;
wire v_43043;
wire v_43044;
wire v_43045;
wire v_43046;
wire v_43047;
wire v_43048;
wire v_43049;
wire v_43050;
wire v_43051;
wire v_43052;
wire v_43053;
wire v_43054;
wire v_43055;
wire v_43056;
wire v_43057;
wire v_43058;
wire v_43059;
wire v_43060;
wire v_43061;
wire v_43062;
wire v_43063;
wire v_43064;
wire v_43065;
wire v_43066;
wire v_43067;
wire v_43068;
wire v_43069;
wire v_43070;
wire v_43071;
wire v_43072;
wire v_43073;
wire v_43074;
wire v_43075;
wire v_43076;
wire v_43077;
wire v_43078;
wire v_43079;
wire v_43080;
wire v_43081;
wire v_43082;
wire v_43083;
wire v_43084;
wire v_43085;
wire v_43086;
wire v_43087;
wire v_43088;
wire v_43089;
wire v_43090;
wire v_43091;
wire v_43092;
wire v_43093;
wire v_43094;
wire v_43095;
wire v_43096;
wire v_43097;
wire v_43098;
wire v_43099;
wire v_43100;
wire v_43101;
wire v_43102;
wire v_43103;
wire v_43104;
wire v_43105;
wire v_43106;
wire v_43107;
wire v_43108;
wire v_43109;
wire v_43110;
wire v_43111;
wire v_43112;
wire v_43113;
wire v_43114;
wire v_43115;
wire v_43116;
wire v_43117;
wire v_43118;
wire v_43119;
wire v_43120;
wire v_43121;
wire v_43122;
wire v_43123;
wire v_43124;
wire v_43125;
wire v_43126;
wire v_43127;
wire v_43128;
wire v_43129;
wire v_43130;
wire v_43131;
wire v_43132;
wire v_43133;
wire v_43134;
wire v_43135;
wire v_43136;
wire v_43137;
wire v_43138;
wire v_43139;
wire v_43140;
wire v_43141;
wire v_43142;
wire v_43143;
wire v_43144;
wire v_43145;
wire v_43146;
wire v_43147;
wire v_43148;
wire v_43149;
wire v_43150;
wire v_43151;
wire v_43152;
wire v_43153;
wire v_43154;
wire v_43155;
wire v_43156;
wire v_43157;
wire v_43158;
wire v_43159;
wire v_43160;
wire v_43161;
wire v_43162;
wire v_43163;
wire v_43164;
wire v_43165;
wire v_43166;
wire v_43167;
wire v_43168;
wire v_43169;
wire v_43170;
wire v_43171;
wire v_43172;
wire v_43173;
wire v_43174;
wire v_43175;
wire v_43176;
wire v_43177;
wire v_43178;
wire v_43179;
wire v_43180;
wire v_43181;
wire v_43182;
wire v_43183;
wire v_43184;
wire v_43185;
wire v_43186;
wire v_43187;
wire v_43188;
wire v_43189;
wire v_43190;
wire v_43191;
wire v_43192;
wire v_43193;
wire v_43194;
wire v_43195;
wire v_43196;
wire v_43197;
wire v_43198;
wire v_43199;
wire v_43200;
wire v_43201;
wire v_43202;
wire v_43203;
wire v_43204;
wire v_43205;
wire v_43206;
wire v_43207;
wire v_43208;
wire v_43209;
wire v_43210;
wire v_43211;
wire v_43212;
wire v_43213;
wire v_43214;
wire v_43215;
wire v_43216;
wire v_43217;
wire v_43218;
wire v_43219;
wire v_43220;
wire v_43221;
wire v_43222;
wire v_43223;
wire v_43224;
wire v_43225;
wire v_43226;
wire v_43227;
wire v_43228;
wire v_43229;
wire v_43230;
wire v_43231;
wire v_43232;
wire v_43233;
wire v_43234;
wire v_43235;
wire v_43236;
wire v_43237;
wire v_43238;
wire v_43239;
wire v_43240;
wire v_43241;
wire v_43242;
wire v_43243;
wire v_43244;
wire v_43245;
wire v_43246;
wire v_43247;
wire v_43248;
wire v_43250;
wire v_43251;
wire v_43252;
wire v_43253;
wire v_43254;
wire v_43255;
wire v_43256;
wire v_43257;
wire v_43258;
wire v_43259;
wire v_43260;
wire v_43261;
wire v_43262;
wire v_43263;
wire v_43264;
wire v_43265;
wire v_43266;
wire v_43267;
wire v_43268;
wire v_43269;
wire v_43270;
wire v_43271;
wire v_43272;
wire v_43273;
wire v_43274;
wire v_43275;
wire v_43276;
wire v_43277;
wire v_43278;
wire v_43279;
wire v_43280;
wire v_43281;
wire v_43282;
wire v_43283;
wire v_43284;
wire v_43285;
wire v_43286;
wire v_43287;
wire v_43288;
wire v_43289;
wire v_43290;
wire v_43291;
wire v_43292;
wire v_43293;
wire v_43294;
wire v_43295;
wire v_43296;
wire v_43297;
wire v_43298;
wire v_43299;
wire v_43300;
wire v_43301;
wire v_43302;
wire v_43303;
wire v_43304;
wire v_43305;
wire v_43306;
wire v_43307;
wire v_43308;
wire v_43309;
wire v_43310;
wire v_43311;
wire v_43312;
wire v_43313;
wire v_43314;
wire v_43315;
wire v_43316;
wire v_43317;
wire v_43318;
wire v_43319;
wire v_43320;
wire v_43321;
wire v_43322;
wire v_43323;
wire v_43324;
wire v_43325;
wire v_43326;
wire v_43327;
wire v_43328;
wire v_43329;
wire v_43330;
wire v_43331;
wire v_43332;
wire v_43333;
wire v_43334;
wire v_43335;
wire v_43336;
wire v_43337;
wire v_43338;
wire v_43339;
wire v_43340;
wire v_43341;
wire v_43342;
wire v_43343;
wire v_43344;
wire v_43345;
wire v_43346;
wire v_43347;
wire v_43348;
wire v_43349;
wire v_43350;
wire v_43351;
wire v_43352;
wire v_43353;
wire v_43354;
wire v_43355;
wire v_43356;
wire v_43357;
wire v_43358;
wire v_43359;
wire v_43360;
wire v_43361;
wire v_43362;
wire v_43363;
wire v_43364;
wire v_43365;
wire v_43366;
wire v_43367;
wire v_43368;
wire v_43369;
wire v_43370;
wire v_43371;
wire v_43372;
wire v_43373;
wire v_43374;
wire v_43375;
wire v_43376;
wire v_43377;
wire v_43378;
wire v_43379;
wire v_43380;
wire v_43381;
wire v_43382;
wire v_43383;
wire v_43384;
wire v_43385;
wire v_43386;
wire v_43387;
wire v_43388;
wire v_43389;
wire v_43390;
wire v_43391;
wire v_43392;
wire v_43393;
wire v_43394;
wire v_43395;
wire v_43396;
wire v_43397;
wire v_43398;
wire v_43399;
wire v_43400;
wire v_43401;
wire v_43402;
wire v_43403;
wire v_43404;
wire v_43405;
wire v_43406;
wire v_43407;
wire v_43408;
wire v_43409;
wire v_43410;
wire v_43411;
wire v_43412;
wire v_43413;
wire v_43414;
wire v_43415;
wire v_43416;
wire v_43417;
wire v_43418;
wire v_43419;
wire v_43420;
wire v_43421;
wire v_43422;
wire v_43423;
wire v_43424;
wire v_43425;
wire v_43426;
wire v_43427;
wire v_43428;
wire v_43429;
wire v_43430;
wire v_43431;
wire v_43432;
wire v_43433;
wire v_43434;
wire v_43435;
wire v_43436;
wire v_43437;
wire v_43438;
wire v_43439;
wire v_43440;
wire v_43441;
wire v_43442;
wire v_43443;
wire v_43444;
wire v_43445;
wire v_43446;
wire v_43447;
wire v_43448;
wire v_43449;
wire v_43450;
wire v_43451;
wire v_43452;
wire v_43453;
wire v_43454;
wire v_43455;
wire v_43456;
wire v_43457;
wire v_43458;
wire v_43459;
wire v_43460;
wire v_43461;
wire v_43462;
wire v_43463;
wire v_43464;
wire v_43465;
wire v_43466;
wire v_43467;
wire v_43468;
wire v_43469;
wire v_43470;
wire v_43471;
wire v_43472;
wire v_43473;
wire v_43474;
wire v_43475;
wire v_43476;
wire v_43477;
wire v_43478;
wire v_43479;
wire v_43480;
wire v_43481;
wire v_43482;
wire v_43483;
wire v_43484;
wire v_43485;
wire v_43486;
wire v_43487;
wire v_43488;
wire v_43489;
wire v_43490;
wire v_43491;
wire v_43493;
wire v_43494;
wire v_43495;
wire v_43496;
wire v_43497;
wire v_43498;
wire v_43499;
wire v_43500;
wire v_43501;
wire v_43502;
wire v_43503;
wire v_43504;
wire v_43505;
wire v_43506;
wire v_43507;
wire v_43508;
wire v_43509;
wire v_43510;
wire v_43511;
wire v_43512;
wire v_43513;
wire v_43514;
wire v_43515;
wire v_43516;
wire v_43517;
wire v_43518;
wire v_43519;
wire v_43520;
wire v_43521;
wire v_43522;
wire v_43523;
wire v_43524;
wire v_43525;
wire v_43526;
wire v_43527;
wire v_43528;
wire v_43529;
wire v_43530;
wire v_43531;
wire v_43532;
wire v_43533;
wire v_43534;
wire v_43535;
wire v_43536;
wire v_43537;
wire v_43538;
wire v_43539;
wire v_43540;
wire v_43541;
wire v_43542;
wire v_43543;
wire v_43544;
wire v_43545;
wire v_43546;
wire v_43547;
wire v_43548;
wire v_43549;
wire v_43550;
wire v_43551;
wire v_43552;
wire v_43553;
wire v_43554;
wire v_43555;
wire v_43556;
wire v_43557;
wire v_43558;
wire v_43559;
wire v_43560;
wire v_43561;
wire v_43562;
wire v_43563;
wire v_43564;
wire v_43565;
wire v_43566;
wire v_43567;
wire v_43568;
wire v_43569;
wire v_43570;
wire v_43571;
wire v_43572;
wire v_43573;
wire v_43574;
wire v_43575;
wire v_43576;
wire v_43577;
wire v_43578;
wire v_43579;
wire v_43580;
wire v_43581;
wire v_43582;
wire v_43583;
wire v_43584;
wire v_43585;
wire v_43586;
wire v_43587;
wire v_43588;
wire v_43589;
wire v_43590;
wire v_43591;
wire v_43592;
wire v_43593;
wire v_43594;
wire v_43595;
wire v_43596;
wire v_43597;
wire v_43598;
wire v_43599;
wire v_43600;
wire v_43601;
wire v_43602;
wire v_43603;
wire v_43604;
wire v_43605;
wire v_43606;
wire v_43607;
wire v_43608;
wire v_43609;
wire v_43610;
wire v_43611;
wire v_43612;
wire v_43613;
wire v_43614;
wire v_43615;
wire v_43616;
wire v_43617;
wire v_43618;
wire v_43619;
wire v_43620;
wire v_43621;
wire v_43622;
wire v_43623;
wire v_43624;
wire v_43625;
wire v_43626;
wire v_43627;
wire v_43628;
wire v_43629;
wire v_43630;
wire v_43631;
wire v_43632;
wire v_43633;
wire v_43634;
wire v_43635;
wire v_43636;
wire v_43637;
wire v_43638;
wire v_43639;
wire v_43640;
wire v_43641;
wire v_43642;
wire v_43643;
wire v_43644;
wire v_43645;
wire v_43646;
wire v_43647;
wire v_43648;
wire v_43649;
wire v_43650;
wire v_43651;
wire v_43652;
wire v_43653;
wire v_43654;
wire v_43655;
wire v_43656;
wire v_43657;
wire v_43658;
wire v_43659;
wire v_43660;
wire v_43661;
wire v_43662;
wire v_43663;
wire v_43664;
wire v_43665;
wire v_43666;
wire v_43667;
wire v_43668;
wire v_43669;
wire v_43670;
wire v_43671;
wire v_43672;
wire v_43673;
wire v_43674;
wire v_43675;
wire v_43676;
wire v_43677;
wire v_43678;
wire v_43679;
wire v_43680;
wire v_43681;
wire v_43682;
wire v_43683;
wire v_43684;
wire v_43685;
wire v_43686;
wire v_43687;
wire v_43688;
wire v_43689;
wire v_43690;
wire v_43691;
wire v_43692;
wire v_43693;
wire v_43694;
wire v_43695;
wire v_43696;
wire v_43697;
wire v_43698;
wire v_43699;
wire v_43700;
wire v_43701;
wire v_43702;
wire v_43703;
wire v_43704;
wire v_43705;
wire v_43706;
wire v_43707;
wire v_43708;
wire v_43709;
wire v_43710;
wire v_43711;
wire v_43712;
wire v_43713;
wire v_43714;
wire v_43715;
wire v_43716;
wire v_43717;
wire v_43718;
wire v_43719;
wire v_43720;
wire v_43721;
wire v_43722;
wire v_43723;
wire v_43724;
wire v_43725;
wire v_43726;
wire v_43727;
wire v_43728;
wire v_43729;
wire v_43730;
wire v_43731;
wire v_43732;
wire v_43733;
wire v_43734;
wire v_43736;
wire v_43737;
wire v_43738;
wire v_43739;
wire v_43740;
wire v_43741;
wire v_43742;
wire v_43743;
wire v_43744;
wire v_43745;
wire v_43746;
wire v_43747;
wire v_43748;
wire v_43749;
wire v_43750;
wire v_43751;
wire v_43752;
wire v_43753;
wire v_43754;
wire v_43755;
wire v_43756;
wire v_43757;
wire v_43758;
wire v_43759;
wire v_43760;
wire v_43761;
wire v_43762;
wire v_43763;
wire v_43764;
wire v_43765;
wire v_43766;
wire v_43767;
wire v_43768;
wire v_43769;
wire v_43770;
wire v_43771;
wire v_43772;
wire v_43773;
wire v_43774;
wire v_43775;
wire v_43776;
wire v_43777;
wire v_43778;
wire v_43779;
wire v_43780;
wire v_43781;
wire v_43782;
wire v_43783;
wire v_43784;
wire v_43785;
wire v_43786;
wire v_43787;
wire v_43788;
wire v_43789;
wire v_43790;
wire v_43791;
wire v_43792;
wire v_43793;
wire v_43794;
wire v_43795;
wire v_43796;
wire v_43797;
wire v_43798;
wire v_43799;
wire v_43800;
wire v_43801;
wire v_43802;
wire v_43803;
wire v_43804;
wire v_43805;
wire v_43806;
wire v_43807;
wire v_43808;
wire v_43809;
wire v_43810;
wire v_43811;
wire v_43812;
wire v_43813;
wire v_43814;
wire v_43815;
wire v_43816;
wire v_43817;
wire v_43818;
wire v_43819;
wire v_43820;
wire v_43821;
wire v_43822;
wire v_43823;
wire v_43824;
wire v_43825;
wire v_43826;
wire v_43827;
wire v_43828;
wire v_43829;
wire v_43830;
wire v_43831;
wire v_43832;
wire v_43833;
wire v_43834;
wire v_43835;
wire v_43836;
wire v_43837;
wire v_43838;
wire v_43839;
wire v_43840;
wire v_43841;
wire v_43842;
wire v_43843;
wire v_43844;
wire v_43845;
wire v_43846;
wire v_43847;
wire v_43848;
wire v_43849;
wire v_43850;
wire v_43851;
wire v_43852;
wire v_43853;
wire v_43854;
wire v_43855;
wire v_43856;
wire v_43857;
wire v_43858;
wire v_43859;
wire v_43860;
wire v_43861;
wire v_43862;
wire v_43863;
wire v_43864;
wire v_43865;
wire v_43866;
wire v_43867;
wire v_43868;
wire v_43869;
wire v_43870;
wire v_43871;
wire v_43872;
wire v_43873;
wire v_43874;
wire v_43875;
wire v_43876;
wire v_43877;
wire v_43878;
wire v_43879;
wire v_43880;
wire v_43881;
wire v_43882;
wire v_43883;
wire v_43884;
wire v_43885;
wire v_43886;
wire v_43887;
wire v_43888;
wire v_43889;
wire v_43890;
wire v_43891;
wire v_43892;
wire v_43893;
wire v_43894;
wire v_43895;
wire v_43896;
wire v_43897;
wire v_43898;
wire v_43899;
wire v_43900;
wire v_43901;
wire v_43902;
wire v_43903;
wire v_43904;
wire v_43905;
wire v_43906;
wire v_43907;
wire v_43908;
wire v_43909;
wire v_43910;
wire v_43911;
wire v_43912;
wire v_43913;
wire v_43914;
wire v_43915;
wire v_43916;
wire v_43917;
wire v_43918;
wire v_43919;
wire v_43920;
wire v_43921;
wire v_43922;
wire v_43923;
wire v_43924;
wire v_43925;
wire v_43926;
wire v_43927;
wire v_43928;
wire v_43929;
wire v_43930;
wire v_43931;
wire v_43932;
wire v_43933;
wire v_43934;
wire v_43935;
wire v_43936;
wire v_43937;
wire v_43938;
wire v_43939;
wire v_43940;
wire v_43941;
wire v_43942;
wire v_43943;
wire v_43944;
wire v_43945;
wire v_43946;
wire v_43947;
wire v_43948;
wire v_43949;
wire v_43950;
wire v_43951;
wire v_43952;
wire v_43953;
wire v_43954;
wire v_43955;
wire v_43956;
wire v_43957;
wire v_43958;
wire v_43959;
wire v_43960;
wire v_43961;
wire v_43962;
wire v_43963;
wire v_43964;
wire v_43965;
wire v_43966;
wire v_43967;
wire v_43968;
wire v_43969;
wire v_43970;
wire v_43971;
wire v_43972;
wire v_43973;
wire v_43974;
wire v_43975;
wire v_43976;
wire v_43977;
wire v_43979;
wire v_43980;
wire v_43981;
wire v_43982;
wire v_43983;
wire v_43984;
wire v_43985;
wire v_43986;
wire v_43987;
wire v_43988;
wire v_43989;
wire v_43990;
wire v_43991;
wire v_43992;
wire v_43993;
wire v_43994;
wire v_43995;
wire v_43996;
wire v_43997;
wire v_43998;
wire v_43999;
wire v_44000;
wire v_44001;
wire v_44002;
wire v_44003;
wire v_44004;
wire v_44005;
wire v_44006;
wire v_44007;
wire v_44008;
wire v_44009;
wire v_44010;
wire v_44011;
wire v_44012;
wire v_44013;
wire v_44014;
wire v_44015;
wire v_44016;
wire v_44017;
wire v_44018;
wire v_44019;
wire v_44020;
wire v_44021;
wire v_44022;
wire v_44023;
wire v_44024;
wire v_44025;
wire v_44026;
wire v_44027;
wire v_44028;
wire v_44029;
wire v_44030;
wire v_44031;
wire v_44032;
wire v_44033;
wire v_44034;
wire v_44035;
wire v_44036;
wire v_44037;
wire v_44038;
wire v_44039;
wire v_44040;
wire v_44041;
wire v_44042;
wire v_44043;
wire v_44044;
wire v_44045;
wire v_44046;
wire v_44047;
wire v_44048;
wire v_44049;
wire v_44050;
wire v_44051;
wire v_44052;
wire v_44053;
wire v_44054;
wire v_44055;
wire v_44056;
wire v_44057;
wire v_44058;
wire v_44059;
wire v_44060;
wire v_44061;
wire v_44062;
wire v_44063;
wire v_44064;
wire v_44065;
wire v_44066;
wire v_44067;
wire v_44068;
wire v_44069;
wire v_44070;
wire v_44071;
wire v_44072;
wire v_44073;
wire v_44074;
wire v_44075;
wire v_44076;
wire v_44077;
wire v_44078;
wire v_44079;
wire v_44080;
wire v_44081;
wire v_44082;
wire v_44083;
wire v_44084;
wire v_44085;
wire v_44086;
wire v_44087;
wire v_44088;
wire v_44089;
wire v_44090;
wire v_44091;
wire v_44092;
wire v_44093;
wire v_44094;
wire v_44095;
wire v_44096;
wire v_44097;
wire v_44098;
wire v_44099;
wire v_44100;
wire v_44101;
wire v_44102;
wire v_44103;
wire v_44104;
wire v_44105;
wire v_44106;
wire v_44107;
wire v_44108;
wire v_44109;
wire v_44110;
wire v_44111;
wire v_44112;
wire v_44113;
wire v_44114;
wire v_44115;
wire v_44116;
wire v_44117;
wire v_44118;
wire v_44119;
wire v_44120;
wire v_44121;
wire v_44122;
wire v_44123;
wire v_44124;
wire v_44125;
wire v_44126;
wire v_44127;
wire v_44128;
wire v_44129;
wire v_44130;
wire v_44131;
wire v_44132;
wire v_44133;
wire v_44134;
wire v_44135;
wire v_44136;
wire v_44137;
wire v_44138;
wire v_44139;
wire v_44140;
wire v_44141;
wire v_44142;
wire v_44143;
wire v_44144;
wire v_44145;
wire v_44146;
wire v_44147;
wire v_44148;
wire v_44149;
wire v_44150;
wire v_44151;
wire v_44152;
wire v_44153;
wire v_44154;
wire v_44155;
wire v_44156;
wire v_44157;
wire v_44158;
wire v_44159;
wire v_44160;
wire v_44161;
wire v_44162;
wire v_44163;
wire v_44164;
wire v_44165;
wire v_44166;
wire v_44167;
wire v_44168;
wire v_44169;
wire v_44170;
wire v_44171;
wire v_44172;
wire v_44173;
wire v_44174;
wire v_44175;
wire v_44176;
wire v_44177;
wire v_44178;
wire v_44179;
wire v_44180;
wire v_44181;
wire v_44182;
wire v_44183;
wire v_44184;
wire v_44185;
wire v_44186;
wire v_44187;
wire v_44188;
wire v_44189;
wire v_44190;
wire v_44191;
wire v_44192;
wire v_44193;
wire v_44194;
wire v_44195;
wire v_44196;
wire v_44197;
wire v_44198;
wire v_44199;
wire v_44200;
wire v_44201;
wire v_44202;
wire v_44203;
wire v_44204;
wire v_44205;
wire v_44206;
wire v_44207;
wire v_44208;
wire v_44209;
wire v_44210;
wire v_44211;
wire v_44212;
wire v_44213;
wire v_44214;
wire v_44215;
wire v_44216;
wire v_44217;
wire v_44218;
wire v_44219;
wire v_44220;
wire v_44222;
wire v_44223;
wire v_44224;
wire v_44225;
wire v_44226;
wire v_44227;
wire v_44228;
wire v_44229;
wire v_44230;
wire v_44231;
wire v_44232;
wire v_44233;
wire v_44234;
wire v_44235;
wire v_44236;
wire v_44237;
wire v_44238;
wire v_44239;
wire v_44240;
wire v_44241;
wire v_44242;
wire v_44243;
wire v_44244;
wire v_44245;
wire v_44246;
wire v_44247;
wire v_44248;
wire v_44249;
wire v_44250;
wire v_44251;
wire v_44252;
wire v_44253;
wire v_44254;
wire v_44255;
wire v_44256;
wire v_44257;
wire v_44258;
wire v_44259;
wire v_44260;
wire v_44261;
wire v_44262;
wire v_44263;
wire v_44264;
wire v_44265;
wire v_44266;
wire v_44267;
wire v_44268;
wire v_44269;
wire v_44270;
wire v_44271;
wire v_44272;
wire v_44273;
wire v_44274;
wire v_44275;
wire v_44276;
wire v_44277;
wire v_44278;
wire v_44279;
wire v_44280;
wire v_44281;
wire v_44282;
wire v_44283;
wire v_44284;
wire v_44285;
wire v_44286;
wire v_44287;
wire v_44288;
wire v_44289;
wire v_44290;
wire v_44291;
wire v_44292;
wire v_44293;
wire v_44294;
wire v_44295;
wire v_44296;
wire v_44297;
wire v_44298;
wire v_44299;
wire v_44300;
wire v_44301;
wire v_44302;
wire v_44303;
wire v_44304;
wire v_44305;
wire v_44306;
wire v_44307;
wire v_44308;
wire v_44309;
wire v_44310;
wire v_44311;
wire v_44312;
wire v_44313;
wire v_44314;
wire v_44315;
wire v_44316;
wire v_44317;
wire v_44318;
wire v_44319;
wire v_44320;
wire v_44321;
wire v_44322;
wire v_44323;
wire v_44324;
wire v_44325;
wire v_44326;
wire v_44327;
wire v_44328;
wire v_44329;
wire v_44330;
wire v_44331;
wire v_44332;
wire v_44333;
wire v_44334;
wire v_44335;
wire v_44336;
wire v_44337;
wire v_44338;
wire v_44339;
wire v_44340;
wire v_44341;
wire v_44342;
wire v_44343;
wire v_44344;
wire v_44345;
wire v_44346;
wire v_44347;
wire v_44348;
wire v_44349;
wire v_44350;
wire v_44351;
wire v_44352;
wire v_44353;
wire v_44354;
wire v_44355;
wire v_44356;
wire v_44357;
wire v_44358;
wire v_44359;
wire v_44360;
wire v_44361;
wire v_44362;
wire v_44363;
wire v_44364;
wire v_44365;
wire v_44366;
wire v_44367;
wire v_44368;
wire v_44369;
wire v_44370;
wire v_44371;
wire v_44372;
wire v_44373;
wire v_44374;
wire v_44375;
wire v_44376;
wire v_44377;
wire v_44378;
wire v_44379;
wire v_44380;
wire v_44381;
wire v_44382;
wire v_44383;
wire v_44384;
wire v_44385;
wire v_44386;
wire v_44387;
wire v_44388;
wire v_44389;
wire v_44390;
wire v_44391;
wire v_44392;
wire v_44393;
wire v_44394;
wire v_44395;
wire v_44396;
wire v_44397;
wire v_44398;
wire v_44399;
wire v_44400;
wire v_44401;
wire v_44402;
wire v_44403;
wire v_44404;
wire v_44405;
wire v_44406;
wire v_44407;
wire v_44408;
wire v_44409;
wire v_44410;
wire v_44411;
wire v_44412;
wire v_44413;
wire v_44414;
wire v_44415;
wire v_44416;
wire v_44417;
wire v_44418;
wire v_44419;
wire v_44420;
wire v_44421;
wire v_44422;
wire v_44423;
wire v_44424;
wire v_44425;
wire v_44426;
wire v_44427;
wire v_44428;
wire v_44429;
wire v_44430;
wire v_44431;
wire v_44432;
wire v_44433;
wire v_44434;
wire v_44435;
wire v_44436;
wire v_44437;
wire v_44438;
wire v_44439;
wire v_44440;
wire v_44441;
wire v_44442;
wire v_44443;
wire v_44444;
wire v_44445;
wire v_44446;
wire v_44447;
wire v_44448;
wire v_44449;
wire v_44450;
wire v_44451;
wire v_44452;
wire v_44453;
wire v_44454;
wire v_44455;
wire v_44456;
wire v_44457;
wire v_44458;
wire v_44459;
wire v_44460;
wire v_44461;
wire v_44462;
wire v_44463;
wire v_44465;
wire v_44466;
wire v_44467;
wire v_44468;
wire v_44469;
wire v_44470;
wire v_44471;
wire v_44472;
wire v_44473;
wire v_44474;
wire v_44475;
wire v_44476;
wire v_44477;
wire v_44478;
wire v_44479;
wire v_44480;
wire v_44481;
wire v_44482;
wire v_44483;
wire v_44484;
wire v_44485;
wire v_44486;
wire v_44487;
wire v_44488;
wire v_44489;
wire v_44490;
wire v_44491;
wire v_44492;
wire v_44493;
wire v_44494;
wire v_44495;
wire v_44496;
wire v_44497;
wire v_44498;
wire v_44499;
wire v_44500;
wire v_44501;
wire v_44502;
wire v_44503;
wire v_44504;
wire v_44505;
wire v_44506;
wire v_44507;
wire v_44508;
wire v_44509;
wire v_44510;
wire v_44511;
wire v_44512;
wire v_44513;
wire v_44514;
wire v_44515;
wire v_44516;
wire v_44517;
wire v_44518;
wire v_44519;
wire v_44520;
wire v_44521;
wire v_44522;
wire v_44523;
wire v_44524;
wire v_44525;
wire v_44526;
wire v_44527;
wire v_44528;
wire v_44529;
wire v_44530;
wire v_44531;
wire v_44532;
wire v_44533;
wire v_44534;
wire v_44535;
wire v_44536;
wire v_44537;
wire v_44538;
wire v_44539;
wire v_44540;
wire v_44541;
wire v_44542;
wire v_44543;
wire v_44544;
wire v_44545;
wire v_44546;
wire v_44547;
wire v_44548;
wire v_44549;
wire v_44550;
wire v_44551;
wire v_44552;
wire v_44553;
wire v_44554;
wire v_44555;
wire v_44556;
wire v_44557;
wire v_44558;
wire v_44559;
wire v_44560;
wire v_44561;
wire v_44562;
wire v_44563;
wire v_44564;
wire v_44565;
wire v_44566;
wire v_44567;
wire v_44568;
wire v_44569;
wire v_44570;
wire v_44571;
wire v_44572;
wire v_44573;
wire v_44574;
wire v_44575;
wire v_44576;
wire v_44577;
wire v_44578;
wire v_44579;
wire v_44580;
wire v_44581;
wire v_44582;
wire v_44583;
wire v_44584;
wire v_44585;
wire v_44586;
wire v_44587;
wire v_44588;
wire v_44589;
wire v_44590;
wire v_44591;
wire v_44592;
wire v_44593;
wire v_44594;
wire v_44595;
wire v_44596;
wire v_44597;
wire v_44598;
wire v_44599;
wire v_44600;
wire v_44601;
wire v_44602;
wire v_44603;
wire v_44604;
wire v_44605;
wire v_44606;
wire v_44607;
wire v_44608;
wire v_44609;
wire v_44610;
wire v_44611;
wire v_44612;
wire v_44613;
wire v_44614;
wire v_44615;
wire v_44616;
wire v_44617;
wire v_44618;
wire v_44619;
wire v_44620;
wire v_44621;
wire v_44622;
wire v_44623;
wire v_44624;
wire v_44625;
wire v_44626;
wire v_44627;
wire v_44628;
wire v_44629;
wire v_44630;
wire v_44631;
wire v_44632;
wire v_44633;
wire v_44634;
wire v_44635;
wire v_44636;
wire v_44637;
wire v_44638;
wire v_44639;
wire v_44640;
wire v_44641;
wire v_44642;
wire v_44643;
wire v_44644;
wire v_44645;
wire v_44646;
wire v_44647;
wire v_44648;
wire v_44649;
wire v_44650;
wire v_44651;
wire v_44652;
wire v_44653;
wire v_44654;
wire v_44655;
wire v_44656;
wire v_44657;
wire v_44658;
wire v_44659;
wire v_44660;
wire v_44661;
wire v_44662;
wire v_44663;
wire v_44664;
wire v_44665;
wire v_44666;
wire v_44667;
wire v_44668;
wire v_44669;
wire v_44670;
wire v_44671;
wire v_44672;
wire v_44673;
wire v_44674;
wire v_44675;
wire v_44676;
wire v_44677;
wire v_44678;
wire v_44679;
wire v_44680;
wire v_44681;
wire v_44682;
wire v_44683;
wire v_44684;
wire v_44685;
wire v_44686;
wire v_44687;
wire v_44688;
wire v_44689;
wire v_44690;
wire v_44691;
wire v_44692;
wire v_44693;
wire v_44694;
wire v_44695;
wire v_44696;
wire v_44697;
wire v_44698;
wire v_44699;
wire v_44700;
wire v_44701;
wire v_44702;
wire v_44703;
wire v_44704;
wire v_44705;
wire v_44706;
wire v_44708;
wire v_44709;
wire v_44710;
wire v_44711;
wire v_44712;
wire v_44713;
wire v_44714;
wire v_44715;
wire v_44716;
wire v_44717;
wire v_44718;
wire v_44719;
wire v_44720;
wire v_44721;
wire v_44722;
wire v_44723;
wire v_44724;
wire v_44725;
wire v_44726;
wire v_44727;
wire v_44728;
wire v_44729;
wire v_44730;
wire v_44731;
wire v_44732;
wire v_44733;
wire v_44734;
wire v_44735;
wire v_44736;
wire v_44737;
wire v_44738;
wire v_44739;
wire v_44740;
wire v_44741;
wire v_44742;
wire v_44743;
wire v_44744;
wire v_44745;
wire v_44746;
wire v_44747;
wire v_44748;
wire v_44749;
wire v_44750;
wire v_44751;
wire v_44752;
wire v_44753;
wire v_44754;
wire v_44755;
wire v_44756;
wire v_44757;
wire v_44758;
wire v_44759;
wire v_44760;
wire v_44761;
wire v_44762;
wire v_44763;
wire v_44764;
wire v_44765;
wire v_44766;
wire v_44767;
wire v_44768;
wire v_44769;
wire v_44770;
wire v_44771;
wire v_44772;
wire v_44773;
wire v_44774;
wire v_44775;
wire v_44776;
wire v_44777;
wire v_44778;
wire v_44779;
wire v_44780;
wire v_44781;
wire v_44782;
wire v_44783;
wire v_44784;
wire v_44785;
wire v_44786;
wire v_44787;
wire v_44788;
wire v_44789;
wire v_44790;
wire v_44791;
wire v_44792;
wire v_44793;
wire v_44794;
wire v_44795;
wire v_44796;
wire v_44797;
wire v_44798;
wire v_44799;
wire v_44800;
wire v_44801;
wire v_44802;
wire v_44803;
wire v_44804;
wire v_44805;
wire v_44806;
wire v_44807;
wire v_44808;
wire v_44809;
wire v_44810;
wire v_44811;
wire v_44812;
wire v_44813;
wire v_44814;
wire v_44815;
wire v_44816;
wire v_44817;
wire v_44818;
wire v_44819;
wire v_44820;
wire v_44821;
wire v_44822;
wire v_44823;
wire v_44824;
wire v_44825;
wire v_44826;
wire v_44827;
wire v_44828;
wire v_44829;
wire v_44830;
wire v_44831;
wire v_44832;
wire v_44833;
wire v_44834;
wire v_44835;
wire v_44836;
wire v_44837;
wire v_44838;
wire v_44839;
wire v_44840;
wire v_44841;
wire v_44842;
wire v_44843;
wire v_44844;
wire v_44845;
wire v_44846;
wire v_44847;
wire v_44848;
wire v_44849;
wire v_44850;
wire v_44851;
wire v_44852;
wire v_44853;
wire v_44854;
wire v_44855;
wire v_44856;
wire v_44857;
wire v_44858;
wire v_44859;
wire v_44860;
wire v_44861;
wire v_44862;
wire v_44863;
wire v_44864;
wire v_44865;
wire v_44866;
wire v_44867;
wire v_44868;
wire v_44869;
wire v_44870;
wire v_44871;
wire v_44872;
wire v_44873;
wire v_44874;
wire v_44875;
wire v_44876;
wire v_44877;
wire v_44878;
wire v_44879;
wire v_44880;
wire v_44881;
wire v_44882;
wire v_44883;
wire v_44884;
wire v_44885;
wire v_44886;
wire v_44887;
wire v_44888;
wire v_44889;
wire v_44890;
wire v_44891;
wire v_44892;
wire v_44893;
wire v_44894;
wire v_44895;
wire v_44896;
wire v_44897;
wire v_44898;
wire v_44899;
wire v_44900;
wire v_44901;
wire v_44902;
wire v_44903;
wire v_44904;
wire v_44905;
wire v_44906;
wire v_44907;
wire v_44908;
wire v_44909;
wire v_44910;
wire v_44911;
wire v_44912;
wire v_44913;
wire v_44914;
wire v_44915;
wire v_44916;
wire v_44917;
wire v_44918;
wire v_44919;
wire v_44920;
wire v_44921;
wire v_44922;
wire v_44923;
wire v_44924;
wire v_44925;
wire v_44926;
wire v_44927;
wire v_44928;
wire v_44929;
wire v_44930;
wire v_44931;
wire v_44932;
wire v_44933;
wire v_44934;
wire v_44935;
wire v_44936;
wire v_44937;
wire v_44938;
wire v_44939;
wire v_44940;
wire v_44941;
wire v_44942;
wire v_44943;
wire v_44944;
wire v_44945;
wire v_44946;
wire v_44947;
wire v_44948;
wire v_44949;
wire v_44951;
wire v_44952;
wire v_44953;
wire v_44954;
wire v_44955;
wire v_44956;
wire v_44957;
wire v_44958;
wire v_44959;
wire v_44960;
wire v_44961;
wire v_44962;
wire v_44963;
wire v_44964;
wire v_44965;
wire v_44966;
wire v_44967;
wire v_44968;
wire v_44969;
wire v_44970;
wire v_44971;
wire v_44972;
wire v_44973;
wire v_44974;
wire v_44975;
wire v_44976;
wire v_44977;
wire v_44978;
wire v_44979;
wire v_44980;
wire v_44981;
wire v_44982;
wire v_44983;
wire v_44984;
wire v_44985;
wire v_44986;
wire v_44987;
wire v_44988;
wire v_44989;
wire v_44990;
wire v_44991;
wire v_44992;
wire v_44993;
wire v_44994;
wire v_44995;
wire v_44996;
wire v_44997;
wire v_44998;
wire v_44999;
wire v_45000;
wire v_45001;
wire v_45002;
wire v_45003;
wire v_45004;
wire v_45005;
wire v_45006;
wire v_45007;
wire v_45008;
wire v_45009;
wire v_45010;
wire v_45011;
wire v_45012;
wire v_45013;
wire v_45014;
wire v_45015;
wire v_45016;
wire v_45017;
wire v_45018;
wire v_45019;
wire v_45020;
wire v_45021;
wire v_45022;
wire v_45023;
wire v_45024;
wire v_45025;
wire v_45026;
wire v_45027;
wire v_45028;
wire v_45029;
wire v_45030;
wire v_45031;
wire v_45032;
wire v_45033;
wire v_45034;
wire v_45035;
wire v_45036;
wire v_45037;
wire v_45038;
wire v_45039;
wire v_45040;
wire v_45041;
wire v_45042;
wire v_45043;
wire v_45044;
wire v_45045;
wire v_45046;
wire v_45047;
wire v_45048;
wire v_45049;
wire v_45050;
wire v_45051;
wire v_45052;
wire v_45053;
wire v_45054;
wire v_45055;
wire v_45056;
wire v_45057;
wire v_45058;
wire v_45059;
wire v_45060;
wire v_45061;
wire v_45062;
wire v_45063;
wire v_45064;
wire v_45065;
wire v_45066;
wire v_45067;
wire v_45068;
wire v_45069;
wire v_45070;
wire v_45071;
wire v_45072;
wire v_45073;
wire v_45074;
wire v_45075;
wire v_45076;
wire v_45077;
wire v_45078;
wire v_45079;
wire v_45080;
wire v_45081;
wire v_45082;
wire v_45083;
wire v_45084;
wire v_45085;
wire v_45086;
wire v_45087;
wire v_45088;
wire v_45089;
wire v_45090;
wire v_45091;
wire v_45092;
wire v_45093;
wire v_45094;
wire v_45095;
wire v_45096;
wire v_45097;
wire v_45098;
wire v_45099;
wire v_45100;
wire v_45101;
wire v_45102;
wire v_45103;
wire v_45104;
wire v_45105;
wire v_45106;
wire v_45107;
wire v_45108;
wire v_45109;
wire v_45110;
wire v_45111;
wire v_45112;
wire v_45113;
wire v_45114;
wire v_45115;
wire v_45116;
wire v_45117;
wire v_45118;
wire v_45119;
wire v_45120;
wire v_45121;
wire v_45122;
wire v_45123;
wire v_45124;
wire v_45125;
wire v_45126;
wire v_45127;
wire v_45128;
wire v_45129;
wire v_45130;
wire v_45131;
wire v_45132;
wire v_45133;
wire v_45134;
wire v_45135;
wire v_45136;
wire v_45137;
wire v_45138;
wire v_45139;
wire v_45140;
wire v_45141;
wire v_45142;
wire v_45143;
wire v_45144;
wire v_45145;
wire v_45146;
wire v_45147;
wire v_45148;
wire v_45149;
wire v_45150;
wire v_45151;
wire v_45152;
wire v_45153;
wire v_45154;
wire v_45155;
wire v_45156;
wire v_45157;
wire v_45158;
wire v_45159;
wire v_45160;
wire v_45161;
wire v_45162;
wire v_45163;
wire v_45164;
wire v_45165;
wire v_45166;
wire v_45167;
wire v_45168;
wire v_45169;
wire v_45170;
wire v_45171;
wire v_45172;
wire v_45173;
wire v_45174;
wire v_45175;
wire v_45176;
wire v_45177;
wire v_45178;
wire v_45179;
wire v_45180;
wire v_45181;
wire v_45182;
wire v_45183;
wire v_45184;
wire v_45185;
wire v_45186;
wire v_45187;
wire v_45188;
wire v_45189;
wire v_45190;
wire v_45191;
wire v_45192;
wire v_45194;
wire v_45195;
wire v_45196;
wire v_45197;
wire v_45198;
wire v_45199;
wire v_45200;
wire v_45201;
wire v_45202;
wire v_45203;
wire v_45204;
wire v_45205;
wire v_45206;
wire v_45207;
wire v_45208;
wire v_45209;
wire v_45210;
wire v_45211;
wire v_45212;
wire v_45213;
wire v_45214;
wire v_45215;
wire v_45216;
wire v_45217;
wire v_45218;
wire v_45219;
wire v_45220;
wire v_45221;
wire v_45222;
wire v_45223;
wire v_45224;
wire v_45225;
wire v_45226;
wire v_45227;
wire v_45228;
wire v_45229;
wire v_45230;
wire v_45231;
wire v_45232;
wire v_45233;
wire v_45234;
wire v_45235;
wire v_45236;
wire v_45237;
wire v_45238;
wire v_45239;
wire v_45240;
wire v_45241;
wire v_45242;
wire v_45243;
wire v_45244;
wire v_45245;
wire v_45246;
wire v_45247;
wire v_45248;
wire v_45249;
wire v_45250;
wire v_45251;
wire v_45252;
wire v_45253;
wire v_45254;
wire v_45255;
wire v_45256;
wire v_45257;
wire v_45258;
wire v_45259;
wire v_45260;
wire v_45261;
wire v_45262;
wire v_45263;
wire v_45264;
wire v_45265;
wire v_45266;
wire v_45267;
wire v_45268;
wire v_45269;
wire v_45270;
wire v_45271;
wire v_45272;
wire v_45273;
wire v_45274;
wire v_45275;
wire v_45276;
wire v_45277;
wire v_45278;
wire v_45279;
wire v_45280;
wire v_45281;
wire v_45282;
wire v_45283;
wire v_45284;
wire v_45285;
wire v_45286;
wire v_45287;
wire v_45288;
wire v_45289;
wire v_45290;
wire v_45291;
wire v_45292;
wire v_45293;
wire v_45294;
wire v_45295;
wire v_45296;
wire v_45297;
wire v_45298;
wire v_45299;
wire v_45300;
wire v_45301;
wire v_45302;
wire v_45303;
wire v_45304;
wire v_45305;
wire v_45306;
wire v_45307;
wire v_45308;
wire v_45309;
wire v_45310;
wire v_45311;
wire v_45312;
wire v_45313;
wire v_45314;
wire v_45315;
wire v_45316;
wire v_45317;
wire v_45318;
wire v_45319;
wire v_45320;
wire v_45321;
wire v_45322;
wire v_45323;
wire v_45324;
wire v_45325;
wire v_45326;
wire v_45327;
wire v_45328;
wire v_45329;
wire v_45330;
wire v_45331;
wire v_45332;
wire v_45333;
wire v_45334;
wire v_45335;
wire v_45336;
wire v_45337;
wire v_45338;
wire v_45339;
wire v_45340;
wire v_45341;
wire v_45342;
wire v_45343;
wire v_45344;
wire v_45345;
wire v_45346;
wire v_45347;
wire v_45348;
wire v_45349;
wire v_45350;
wire v_45351;
wire v_45352;
wire v_45353;
wire v_45354;
wire v_45355;
wire v_45356;
wire v_45357;
wire v_45358;
wire v_45359;
wire v_45360;
wire v_45361;
wire v_45362;
wire v_45363;
wire v_45364;
wire v_45365;
wire v_45366;
wire v_45367;
wire v_45368;
wire v_45369;
wire v_45370;
wire v_45371;
wire v_45372;
wire v_45373;
wire v_45374;
wire v_45375;
wire v_45376;
wire v_45377;
wire v_45378;
wire v_45379;
wire v_45380;
wire v_45381;
wire v_45382;
wire v_45383;
wire v_45384;
wire v_45385;
wire v_45386;
wire v_45387;
wire v_45388;
wire v_45389;
wire v_45390;
wire v_45391;
wire v_45392;
wire v_45393;
wire v_45394;
wire v_45395;
wire v_45396;
wire v_45397;
wire v_45398;
wire v_45399;
wire v_45400;
wire v_45401;
wire v_45402;
wire v_45403;
wire v_45404;
wire v_45405;
wire v_45406;
wire v_45407;
wire v_45408;
wire v_45409;
wire v_45410;
wire v_45411;
wire v_45412;
wire v_45413;
wire v_45414;
wire v_45415;
wire v_45416;
wire v_45417;
wire v_45418;
wire v_45419;
wire v_45420;
wire v_45421;
wire v_45422;
wire v_45423;
wire v_45424;
wire v_45425;
wire v_45426;
wire v_45427;
wire v_45428;
wire v_45429;
wire v_45430;
wire v_45431;
wire v_45432;
wire v_45433;
wire v_45434;
wire v_45435;
wire v_45437;
wire v_45438;
wire v_45439;
wire v_45440;
wire v_45441;
wire v_45442;
wire v_45443;
wire v_45444;
wire v_45445;
wire v_45446;
wire v_45447;
wire v_45448;
wire v_45449;
wire v_45450;
wire v_45451;
wire v_45452;
wire v_45453;
wire v_45454;
wire v_45455;
wire v_45456;
wire v_45457;
wire v_45458;
wire v_45459;
wire v_45460;
wire v_45461;
wire v_45462;
wire v_45463;
wire v_45464;
wire v_45465;
wire v_45466;
wire v_45467;
wire v_45468;
wire v_45469;
wire v_45470;
wire v_45471;
wire v_45472;
wire v_45473;
wire v_45474;
wire v_45475;
wire v_45476;
wire v_45477;
wire v_45478;
wire v_45479;
wire v_45480;
wire v_45481;
wire v_45482;
wire v_45483;
wire v_45484;
wire v_45485;
wire v_45486;
wire v_45487;
wire v_45488;
wire v_45489;
wire v_45490;
wire v_45491;
wire v_45492;
wire v_45493;
wire v_45494;
wire v_45495;
wire v_45496;
wire v_45497;
wire v_45498;
wire v_45499;
wire v_45500;
wire v_45501;
wire v_45502;
wire v_45503;
wire v_45504;
wire v_45505;
wire v_45506;
wire v_45507;
wire v_45508;
wire v_45509;
wire v_45510;
wire v_45511;
wire v_45512;
wire v_45513;
wire v_45514;
wire v_45515;
wire v_45516;
wire v_45517;
wire v_45518;
wire v_45519;
wire v_45520;
wire v_45521;
wire v_45522;
wire v_45523;
wire v_45524;
wire v_45525;
wire v_45526;
wire v_45527;
wire v_45528;
wire v_45529;
wire v_45530;
wire v_45531;
wire v_45532;
wire v_45533;
wire v_45534;
wire v_45535;
wire v_45536;
wire v_45537;
wire v_45538;
wire v_45539;
wire v_45540;
wire v_45541;
wire v_45542;
wire v_45543;
wire v_45544;
wire v_45545;
wire v_45546;
wire v_45547;
wire v_45548;
wire v_45549;
wire v_45550;
wire v_45551;
wire v_45552;
wire v_45553;
wire v_45554;
wire v_45555;
wire v_45556;
wire v_45557;
wire v_45558;
wire v_45559;
wire v_45560;
wire v_45561;
wire v_45562;
wire v_45563;
wire v_45564;
wire v_45565;
wire v_45566;
wire v_45567;
wire v_45568;
wire v_45569;
wire v_45570;
wire v_45571;
wire v_45572;
wire v_45573;
wire v_45574;
wire v_45575;
wire v_45576;
wire v_45577;
wire v_45578;
wire v_45579;
wire v_45580;
wire v_45581;
wire v_45582;
wire v_45583;
wire v_45584;
wire v_45585;
wire v_45586;
wire v_45587;
wire v_45588;
wire v_45589;
wire v_45590;
wire v_45591;
wire v_45592;
wire v_45593;
wire v_45594;
wire v_45595;
wire v_45596;
wire v_45597;
wire v_45598;
wire v_45599;
wire v_45600;
wire v_45601;
wire v_45602;
wire v_45603;
wire v_45604;
wire v_45605;
wire v_45606;
wire v_45607;
wire v_45608;
wire v_45609;
wire v_45610;
wire v_45611;
wire v_45612;
wire v_45613;
wire v_45614;
wire v_45615;
wire v_45616;
wire v_45617;
wire v_45618;
wire v_45619;
wire v_45620;
wire v_45621;
wire v_45622;
wire v_45623;
wire v_45624;
wire v_45625;
wire v_45626;
wire v_45627;
wire v_45628;
wire v_45629;
wire v_45630;
wire v_45631;
wire v_45632;
wire v_45633;
wire v_45634;
wire v_45635;
wire v_45636;
wire v_45637;
wire v_45638;
wire v_45639;
wire v_45640;
wire v_45641;
wire v_45642;
wire v_45643;
wire v_45644;
wire v_45645;
wire v_45646;
wire v_45647;
wire v_45648;
wire v_45649;
wire v_45650;
wire v_45651;
wire v_45652;
wire v_45653;
wire v_45654;
wire v_45655;
wire v_45656;
wire v_45657;
wire v_45658;
wire v_45659;
wire v_45660;
wire v_45661;
wire v_45662;
wire v_45663;
wire v_45664;
wire v_45665;
wire v_45666;
wire v_45667;
wire v_45668;
wire v_45669;
wire v_45670;
wire v_45671;
wire v_45672;
wire v_45673;
wire v_45674;
wire v_45675;
wire v_45676;
wire v_45677;
wire v_45678;
wire v_45679;
wire v_45680;
wire v_45681;
wire v_45682;
wire v_45683;
wire v_45684;
wire v_45685;
wire v_45686;
wire v_45687;
wire v_45688;
wire v_45689;
wire v_45690;
wire v_45691;
wire v_45692;
wire v_45693;
wire v_45694;
wire v_45695;
wire v_45696;
wire v_45697;
wire v_45698;
wire v_45699;
wire v_45700;
wire v_45701;
wire v_45702;
wire v_45703;
wire v_45704;
wire v_45705;
wire v_45706;
wire v_45707;
wire v_45708;
wire v_45709;
wire v_45710;
wire v_45711;
wire v_45712;
wire v_45713;
wire v_45714;
wire v_45715;
wire v_45716;
wire v_45717;
wire v_45718;
wire v_45719;
wire v_45720;
wire v_45721;
wire v_45722;
wire v_45723;
wire v_45724;
wire v_45725;
wire v_45726;
wire v_45727;
wire v_45728;
wire v_45729;
wire v_45730;
wire v_45731;
wire v_45732;
wire v_45733;
wire v_45734;
wire v_45735;
wire v_45736;
wire v_45737;
wire v_45738;
wire v_45739;
wire v_45740;
wire v_45741;
wire v_45742;
wire v_45743;
wire v_45744;
wire v_45745;
wire v_45746;
wire v_45747;
wire v_45748;
wire v_45749;
wire v_45750;
wire v_45751;
wire v_45752;
wire v_45753;
wire v_45754;
wire v_45755;
wire v_45756;
wire v_45757;
wire v_45758;
wire v_45759;
wire v_45760;
wire v_45761;
wire v_45762;
wire v_45763;
wire v_45764;
wire v_45765;
wire v_45766;
wire v_45767;
wire v_45768;
wire v_45769;
wire v_45770;
wire v_45771;
wire v_45772;
wire v_45773;
wire v_45774;
wire v_45775;
wire v_45776;
wire v_45777;
wire v_45778;
wire v_45779;
wire v_45780;
wire v_45781;
wire v_45782;
wire v_45783;
wire v_45784;
wire v_45785;
wire v_45786;
wire v_45787;
wire v_45788;
wire v_45789;
wire v_45790;
wire v_45791;
wire v_45792;
wire v_45793;
wire v_45794;
wire v_45795;
wire v_45796;
wire v_45797;
wire v_45798;
wire v_45799;
wire v_45800;
wire v_45801;
wire v_45802;
wire v_45803;
wire v_45804;
wire v_45805;
wire v_45806;
wire v_45807;
wire v_45808;
wire v_45809;
wire v_45810;
wire v_45811;
wire v_45812;
wire v_45813;
wire v_45814;
wire v_45815;
wire v_45816;
wire v_45817;
wire v_45818;
wire v_45819;
wire v_45820;
wire v_45821;
wire v_45822;
wire v_45823;
wire v_45824;
wire v_45825;
wire v_45826;
wire v_45827;
wire v_45829;
wire v_45830;
wire v_45831;
wire v_45832;
wire v_45833;
wire v_45834;
wire v_45835;
wire v_45836;
wire v_45837;
wire v_45838;
wire v_45839;
wire v_45840;
wire v_45841;
wire v_45842;
wire v_45843;
wire v_45844;
wire v_45845;
wire v_45846;
wire v_45847;
wire v_45848;
wire v_45849;
wire v_45850;
wire v_45851;
wire v_45852;
wire v_45853;
wire v_45854;
wire v_45855;
wire v_45856;
wire v_45857;
wire v_45858;
wire v_45859;
wire v_45860;
wire v_45861;
wire v_45862;
wire v_45863;
wire v_45864;
wire v_45865;
wire v_45866;
wire v_45867;
wire v_45868;
wire v_45869;
wire v_45870;
wire v_45871;
wire v_45872;
wire v_45873;
wire v_45874;
wire v_45875;
wire v_45876;
wire v_45877;
wire v_45878;
wire v_45879;
wire v_45880;
wire v_45881;
wire v_45882;
wire v_45883;
wire v_45884;
wire v_45885;
wire v_45886;
wire v_45887;
wire v_45888;
wire v_45889;
wire v_45890;
wire v_45891;
wire v_45892;
wire v_45893;
wire v_45894;
wire v_45895;
wire v_45896;
wire v_45897;
wire v_45898;
wire v_45899;
wire v_45900;
wire v_45901;
wire v_45902;
wire v_45903;
wire v_45904;
wire v_45905;
wire v_45906;
wire v_45907;
wire v_45908;
wire v_45909;
wire v_45910;
wire v_45911;
wire v_45912;
wire v_45913;
wire v_45914;
wire v_45915;
wire v_45916;
wire v_45917;
wire v_45918;
wire v_45919;
wire v_45920;
wire v_45921;
wire v_45923;
wire v_45925;
wire v_45926;
wire v_45927;
wire v_45929;
wire v_45930;
wire v_45931;
wire v_45933;
wire v_45934;
wire v_45935;
wire v_45937;
wire v_45938;
wire v_45940;
wire v_45941;
wire v_45942;
wire v_45944;
wire v_45945;
wire v_45946;
wire v_45948;
wire v_45949;
wire v_45950;
wire v_45952;
wire v_45953;
wire v_45954;
wire v_45956;
wire v_45957;
wire v_45958;
wire v_45960;
wire v_45961;
wire v_45962;
wire v_45964;
wire v_45965;
wire v_45966;
wire v_45968;
wire v_45969;
wire v_45970;
wire v_45972;
wire v_45973;
wire v_45974;
wire v_45976;
wire v_45977;
wire v_45978;
wire v_45980;
wire v_45981;
wire v_45982;
wire v_45984;
wire v_45985;
wire v_45986;
wire v_45988;
wire v_45989;
wire v_45990;
wire v_45991;
wire v_45992;
wire v_45993;
wire v_45994;
wire v_45995;
wire v_45996;
wire v_45997;
wire v_45998;
wire v_45999;
wire v_46000;
wire v_46001;
wire v_46002;
wire v_46003;
wire v_46004;
wire v_46005;
wire v_46006;
wire v_46007;
wire v_46008;
wire v_46009;
wire v_46010;
wire v_46011;
wire v_46012;
wire v_46013;
wire v_46014;
wire v_46015;
wire v_46016;
wire v_46017;
wire v_46018;
wire v_46019;
wire v_46020;
wire v_46021;
wire v_46022;
wire v_46023;
wire v_46024;
wire v_46025;
wire v_46026;
wire v_46027;
wire v_46028;
wire v_46029;
wire v_46030;
wire v_46031;
wire v_46032;
wire v_46033;
wire v_46034;
wire v_46035;
wire v_46036;
wire v_46037;
wire v_46038;
wire v_46039;
wire v_46040;
wire v_46041;
wire v_46042;
wire v_46043;
wire v_46044;
wire v_46045;
wire v_46046;
wire v_46047;
wire v_46048;
wire v_46049;
wire v_46050;
wire v_46051;
wire v_46052;
wire v_46053;
wire v_46054;
wire v_46055;
wire v_46056;
wire v_46057;
wire v_46058;
wire v_46059;
wire v_46060;
wire v_46061;
wire v_46062;
wire v_46063;
wire v_46064;
wire v_46065;
wire v_46066;
wire v_46067;
wire v_46068;
wire v_46069;
wire v_46070;
wire v_46071;
wire v_46072;
wire v_46073;
wire v_46074;
wire v_46075;
wire v_46076;
wire v_46077;
wire v_46078;
wire v_46079;
wire v_46080;
wire v_46081;
wire v_46082;
wire v_46083;
wire v_46084;
wire v_46085;
wire v_46086;
wire v_46087;
wire v_46088;
wire v_46089;
wire v_46090;
wire v_46091;
wire v_46092;
wire v_46093;
wire v_46094;
wire v_46095;
wire v_46096;
wire v_46097;
wire v_46098;
wire v_46099;
wire v_46100;
wire v_46101;
wire v_46102;
wire v_46103;
wire v_46104;
wire v_46105;
wire v_46106;
wire v_46107;
wire v_46108;
wire v_46109;
wire v_46110;
wire v_46111;
wire v_46112;
wire v_46113;
wire v_46114;
wire v_46115;
wire v_46116;
wire v_46117;
wire v_46118;
wire v_46119;
wire v_46120;
wire v_46121;
wire v_46122;
wire v_46123;
wire v_46124;
wire v_46125;
wire v_46126;
wire v_46127;
wire v_46128;
wire v_46129;
wire v_46130;
wire v_46131;
wire v_46132;
wire v_46133;
wire v_46134;
wire v_46135;
wire v_46136;
wire v_46137;
wire v_46138;
wire v_46139;
wire v_46140;
wire v_46141;
wire v_46142;
wire v_46143;
wire v_46144;
wire v_46145;
wire v_46146;
wire v_46147;
wire v_46148;
wire v_46149;
wire v_46150;
wire v_46151;
wire v_46152;
wire v_46153;
wire v_46154;
wire v_46155;
wire v_46156;
wire v_46157;
wire v_46158;
wire v_46159;
wire v_46160;
wire v_46161;
wire v_46162;
wire v_46163;
wire v_46164;
wire v_46165;
wire v_46166;
wire v_46167;
wire v_46168;
wire v_46169;
wire v_46170;
wire v_46171;
wire v_46172;
wire v_46173;
wire v_46174;
wire v_46175;
wire v_46176;
wire v_46177;
wire v_46178;
wire v_46179;
wire v_46180;
wire v_46181;
wire v_46183;
wire v_46184;
wire v_46185;
wire v_46186;
wire v_46187;
wire v_46188;
wire v_46189;
wire v_46190;
wire v_46191;
wire v_46192;
wire v_46193;
wire v_46194;
wire v_46195;
wire v_46196;
wire v_46197;
wire v_46198;
wire v_46199;
wire v_46200;
wire v_46201;
wire v_46202;
wire v_46203;
wire v_46204;
wire v_46205;
wire v_46206;
wire v_46207;
wire v_46208;
wire v_46209;
wire v_46210;
wire v_46211;
wire v_46212;
wire v_46213;
wire v_46214;
wire v_46215;
wire v_46216;
wire v_46217;
wire v_46218;
wire v_46219;
wire v_46220;
wire v_46221;
wire v_46222;
wire v_46223;
wire v_46224;
wire v_46225;
wire v_46226;
wire v_46227;
wire v_46228;
wire v_46229;
wire v_46230;
wire v_46231;
wire v_46232;
wire v_46233;
wire v_46234;
wire v_46235;
wire v_46236;
wire v_46237;
wire v_46238;
wire v_46239;
wire v_46240;
wire v_46241;
wire v_46242;
wire v_46243;
wire v_46244;
wire v_46245;
wire v_46246;
wire v_46247;
wire v_46248;
wire v_46249;
wire v_46250;
wire v_46251;
wire v_46252;
wire v_46253;
wire v_46254;
wire v_46255;
wire v_46256;
wire v_46257;
wire v_46258;
wire v_46259;
wire v_46260;
wire v_46261;
wire v_46262;
wire v_46263;
wire v_46264;
wire v_46265;
wire v_46266;
wire v_46267;
wire v_46268;
wire v_46269;
wire v_46270;
wire v_46271;
wire v_46272;
wire v_46273;
wire v_46274;
wire v_46275;
wire v_46276;
wire v_46277;
wire v_46278;
wire v_46279;
wire v_46280;
wire v_46281;
wire v_46282;
wire v_46283;
wire v_46284;
wire v_46285;
wire v_46286;
wire v_46287;
wire v_46288;
wire v_46289;
wire v_46290;
wire v_46291;
wire v_46292;
wire v_46293;
wire v_46294;
wire v_46295;
wire v_46296;
wire v_46297;
wire v_46298;
wire v_46299;
wire v_46300;
wire v_46301;
wire v_46302;
wire v_46303;
wire v_46304;
wire v_46305;
wire v_46306;
wire v_46307;
wire v_46308;
wire v_46309;
wire v_46310;
wire v_46311;
wire v_46312;
wire v_46313;
wire v_46314;
wire v_46315;
wire v_46316;
wire v_46317;
wire v_46318;
wire v_46319;
wire v_46320;
wire v_46321;
wire v_46322;
wire v_46323;
wire v_46324;
wire v_46325;
wire v_46326;
wire v_46327;
wire v_46328;
wire v_46329;
wire v_46330;
wire v_46331;
wire v_46332;
wire v_46333;
wire v_46334;
wire v_46335;
wire v_46336;
wire v_46337;
wire v_46338;
wire v_46339;
wire v_46340;
wire v_46341;
wire v_46342;
wire v_46343;
wire v_46344;
wire v_46345;
wire v_46346;
wire v_46347;
wire v_46348;
wire v_46349;
wire v_46350;
wire v_46351;
wire v_46352;
wire v_46353;
wire v_46354;
wire v_46355;
wire v_46356;
wire v_46357;
wire v_46358;
wire v_46359;
wire v_46360;
wire v_46361;
wire v_46362;
wire v_46363;
wire v_46364;
wire v_46365;
wire v_46366;
wire v_46367;
wire v_46368;
wire v_46369;
wire v_46370;
wire v_46371;
wire v_46372;
wire v_46373;
wire v_46374;
wire v_46375;
wire v_46376;
wire v_46377;
wire v_46378;
wire v_46379;
wire v_46380;
wire v_46381;
wire v_46382;
wire v_46383;
wire v_46384;
wire v_46385;
wire v_46386;
wire v_46387;
wire v_46388;
wire v_46389;
wire v_46390;
wire v_46391;
wire v_46392;
wire v_46393;
wire v_46394;
wire v_46395;
wire v_46396;
wire v_46397;
wire v_46398;
wire v_46399;
wire v_46400;
wire v_46401;
wire v_46402;
wire v_46403;
wire v_46404;
wire v_46405;
wire v_46406;
wire v_46407;
wire v_46408;
wire v_46409;
wire v_46410;
wire v_46411;
wire v_46412;
wire v_46413;
wire v_46414;
wire v_46415;
wire v_46416;
wire v_46417;
wire v_46418;
wire v_46419;
wire v_46420;
wire v_46421;
wire v_46422;
wire v_46423;
wire v_46424;
wire v_46426;
wire v_46427;
wire v_46428;
wire v_46429;
wire v_46430;
wire v_46431;
wire v_46432;
wire v_46433;
wire v_46434;
wire v_46435;
wire v_46436;
wire v_46437;
wire v_46438;
wire v_46439;
wire v_46440;
wire v_46441;
wire v_46442;
wire v_46443;
wire v_46444;
wire v_46445;
wire v_46446;
wire v_46447;
wire v_46448;
wire v_46449;
wire v_46450;
wire v_46451;
wire v_46452;
wire v_46453;
wire v_46454;
wire v_46455;
wire v_46456;
wire v_46457;
wire v_46458;
wire v_46459;
wire v_46460;
wire v_46461;
wire v_46462;
wire v_46463;
wire v_46464;
wire v_46465;
wire v_46466;
wire v_46467;
wire v_46468;
wire v_46469;
wire v_46470;
wire v_46471;
wire v_46472;
wire v_46473;
wire v_46474;
wire v_46475;
wire v_46476;
wire v_46477;
wire v_46478;
wire v_46479;
wire v_46480;
wire v_46481;
wire v_46482;
wire v_46483;
wire v_46484;
wire v_46485;
wire v_46486;
wire v_46487;
wire v_46488;
wire v_46489;
wire v_46490;
wire v_46491;
wire v_46492;
wire v_46493;
wire v_46494;
wire v_46495;
wire v_46496;
wire v_46497;
wire v_46498;
wire v_46499;
wire v_46500;
wire v_46501;
wire v_46502;
wire v_46503;
wire v_46504;
wire v_46505;
wire v_46506;
wire v_46507;
wire v_46508;
wire v_46509;
wire v_46510;
wire v_46511;
wire v_46512;
wire v_46513;
wire v_46514;
wire v_46515;
wire v_46516;
wire v_46517;
wire v_46518;
wire v_46519;
wire v_46520;
wire v_46521;
wire v_46522;
wire v_46523;
wire v_46524;
wire v_46525;
wire v_46526;
wire v_46527;
wire v_46528;
wire v_46529;
wire v_46530;
wire v_46531;
wire v_46532;
wire v_46533;
wire v_46534;
wire v_46535;
wire v_46536;
wire v_46537;
wire v_46538;
wire v_46539;
wire v_46540;
wire v_46541;
wire v_46542;
wire v_46543;
wire v_46544;
wire v_46545;
wire v_46546;
wire v_46547;
wire v_46548;
wire v_46549;
wire v_46550;
wire v_46551;
wire v_46552;
wire v_46553;
wire v_46554;
wire v_46555;
wire v_46556;
wire v_46557;
wire v_46558;
wire v_46559;
wire v_46560;
wire v_46561;
wire v_46562;
wire v_46563;
wire v_46564;
wire v_46565;
wire v_46566;
wire v_46567;
wire v_46568;
wire v_46569;
wire v_46570;
wire v_46571;
wire v_46572;
wire v_46573;
wire v_46574;
wire v_46575;
wire v_46576;
wire v_46577;
wire v_46578;
wire v_46579;
wire v_46580;
wire v_46581;
wire v_46582;
wire v_46583;
wire v_46584;
wire v_46585;
wire v_46586;
wire v_46587;
wire v_46588;
wire v_46589;
wire v_46590;
wire v_46591;
wire v_46592;
wire v_46593;
wire v_46594;
wire v_46595;
wire v_46596;
wire v_46597;
wire v_46598;
wire v_46599;
wire v_46600;
wire v_46601;
wire v_46602;
wire v_46603;
wire v_46604;
wire v_46605;
wire v_46606;
wire v_46607;
wire v_46608;
wire v_46609;
wire v_46610;
wire v_46611;
wire v_46612;
wire v_46613;
wire v_46614;
wire v_46615;
wire v_46616;
wire v_46617;
wire v_46618;
wire v_46619;
wire v_46620;
wire v_46621;
wire v_46622;
wire v_46623;
wire v_46624;
wire v_46625;
wire v_46626;
wire v_46627;
wire v_46628;
wire v_46629;
wire v_46630;
wire v_46631;
wire v_46632;
wire v_46633;
wire v_46634;
wire v_46635;
wire v_46636;
wire v_46637;
wire v_46638;
wire v_46639;
wire v_46640;
wire v_46641;
wire v_46642;
wire v_46643;
wire v_46644;
wire v_46645;
wire v_46646;
wire v_46647;
wire v_46648;
wire v_46649;
wire v_46650;
wire v_46651;
wire v_46652;
wire v_46653;
wire v_46654;
wire v_46655;
wire v_46656;
wire v_46657;
wire v_46658;
wire v_46659;
wire v_46660;
wire v_46661;
wire v_46662;
wire v_46663;
wire v_46664;
wire v_46665;
wire v_46666;
wire v_46667;
wire v_46669;
wire v_46670;
wire v_46671;
wire v_46672;
wire v_46673;
wire v_46674;
wire v_46675;
wire v_46676;
wire v_46677;
wire v_46678;
wire v_46679;
wire v_46680;
wire v_46681;
wire v_46682;
wire v_46683;
wire v_46684;
wire v_46685;
wire v_46686;
wire v_46687;
wire v_46688;
wire v_46689;
wire v_46690;
wire v_46691;
wire v_46692;
wire v_46693;
wire v_46694;
wire v_46695;
wire v_46696;
wire v_46697;
wire v_46698;
wire v_46699;
wire v_46700;
wire v_46701;
wire v_46702;
wire v_46703;
wire v_46704;
wire v_46705;
wire v_46706;
wire v_46707;
wire v_46708;
wire v_46709;
wire v_46710;
wire v_46711;
wire v_46712;
wire v_46713;
wire v_46714;
wire v_46715;
wire v_46716;
wire v_46717;
wire v_46718;
wire v_46719;
wire v_46720;
wire v_46721;
wire v_46722;
wire v_46723;
wire v_46724;
wire v_46725;
wire v_46726;
wire v_46727;
wire v_46728;
wire v_46729;
wire v_46730;
wire v_46731;
wire v_46732;
wire v_46733;
wire v_46734;
wire v_46735;
wire v_46736;
wire v_46737;
wire v_46738;
wire v_46739;
wire v_46740;
wire v_46741;
wire v_46742;
wire v_46743;
wire v_46744;
wire v_46745;
wire v_46746;
wire v_46747;
wire v_46748;
wire v_46749;
wire v_46750;
wire v_46751;
wire v_46752;
wire v_46753;
wire v_46754;
wire v_46755;
wire v_46756;
wire v_46757;
wire v_46758;
wire v_46759;
wire v_46760;
wire v_46761;
wire v_46762;
wire v_46763;
wire v_46764;
wire v_46765;
wire v_46766;
wire v_46767;
wire v_46768;
wire v_46769;
wire v_46770;
wire v_46771;
wire v_46772;
wire v_46773;
wire v_46774;
wire v_46775;
wire v_46776;
wire v_46777;
wire v_46778;
wire v_46779;
wire v_46780;
wire v_46781;
wire v_46782;
wire v_46783;
wire v_46784;
wire v_46785;
wire v_46786;
wire v_46787;
wire v_46788;
wire v_46789;
wire v_46790;
wire v_46791;
wire v_46792;
wire v_46793;
wire v_46794;
wire v_46795;
wire v_46796;
wire v_46797;
wire v_46798;
wire v_46799;
wire v_46800;
wire v_46801;
wire v_46802;
wire v_46803;
wire v_46804;
wire v_46805;
wire v_46806;
wire v_46807;
wire v_46808;
wire v_46809;
wire v_46810;
wire v_46811;
wire v_46812;
wire v_46813;
wire v_46814;
wire v_46815;
wire v_46816;
wire v_46817;
wire v_46818;
wire v_46819;
wire v_46820;
wire v_46821;
wire v_46822;
wire v_46823;
wire v_46824;
wire v_46825;
wire v_46826;
wire v_46827;
wire v_46828;
wire v_46829;
wire v_46830;
wire v_46831;
wire v_46832;
wire v_46833;
wire v_46834;
wire v_46835;
wire v_46836;
wire v_46837;
wire v_46838;
wire v_46839;
wire v_46840;
wire v_46841;
wire v_46842;
wire v_46843;
wire v_46844;
wire v_46845;
wire v_46846;
wire v_46847;
wire v_46848;
wire v_46849;
wire v_46850;
wire v_46851;
wire v_46852;
wire v_46853;
wire v_46854;
wire v_46855;
wire v_46856;
wire v_46857;
wire v_46858;
wire v_46859;
wire v_46860;
wire v_46861;
wire v_46862;
wire v_46863;
wire v_46864;
wire v_46865;
wire v_46866;
wire v_46867;
wire v_46868;
wire v_46869;
wire v_46870;
wire v_46871;
wire v_46872;
wire v_46873;
wire v_46874;
wire v_46875;
wire v_46876;
wire v_46877;
wire v_46878;
wire v_46879;
wire v_46880;
wire v_46881;
wire v_46882;
wire v_46883;
wire v_46884;
wire v_46885;
wire v_46886;
wire v_46887;
wire v_46888;
wire v_46889;
wire v_46890;
wire v_46891;
wire v_46892;
wire v_46893;
wire v_46894;
wire v_46895;
wire v_46896;
wire v_46897;
wire v_46898;
wire v_46899;
wire v_46900;
wire v_46901;
wire v_46902;
wire v_46903;
wire v_46904;
wire v_46905;
wire v_46906;
wire v_46907;
wire v_46908;
wire v_46909;
wire v_46910;
wire v_46912;
wire v_46913;
wire v_46914;
wire v_46915;
wire v_46916;
wire v_46917;
wire v_46918;
wire v_46919;
wire v_46920;
wire v_46921;
wire v_46922;
wire v_46923;
wire v_46924;
wire v_46925;
wire v_46926;
wire v_46927;
wire v_46928;
wire v_46929;
wire v_46930;
wire v_46931;
wire v_46932;
wire v_46933;
wire v_46934;
wire v_46935;
wire v_46936;
wire v_46937;
wire v_46938;
wire v_46939;
wire v_46940;
wire v_46941;
wire v_46942;
wire v_46943;
wire v_46944;
wire v_46945;
wire v_46946;
wire v_46947;
wire v_46948;
wire v_46949;
wire v_46950;
wire v_46951;
wire v_46952;
wire v_46953;
wire v_46954;
wire v_46955;
wire v_46956;
wire v_46957;
wire v_46958;
wire v_46959;
wire v_46960;
wire v_46961;
wire v_46962;
wire v_46963;
wire v_46964;
wire v_46965;
wire v_46966;
wire v_46967;
wire v_46968;
wire v_46969;
wire v_46970;
wire v_46971;
wire v_46972;
wire v_46973;
wire v_46974;
wire v_46975;
wire v_46976;
wire v_46977;
wire v_46978;
wire v_46979;
wire v_46980;
wire v_46981;
wire v_46982;
wire v_46983;
wire v_46984;
wire v_46985;
wire v_46986;
wire v_46987;
wire v_46988;
wire v_46989;
wire v_46990;
wire v_46991;
wire v_46992;
wire v_46993;
wire v_46994;
wire v_46995;
wire v_46996;
wire v_46997;
wire v_46998;
wire v_46999;
wire v_47000;
wire v_47001;
wire v_47002;
wire v_47003;
wire v_47004;
wire v_47005;
wire v_47006;
wire v_47007;
wire v_47008;
wire v_47009;
wire v_47010;
wire v_47011;
wire v_47012;
wire v_47013;
wire v_47014;
wire v_47015;
wire v_47016;
wire v_47017;
wire v_47018;
wire v_47019;
wire v_47020;
wire v_47021;
wire v_47022;
wire v_47023;
wire v_47024;
wire v_47025;
wire v_47026;
wire v_47027;
wire v_47028;
wire v_47029;
wire v_47030;
wire v_47031;
wire v_47032;
wire v_47033;
wire v_47034;
wire v_47035;
wire v_47036;
wire v_47037;
wire v_47038;
wire v_47039;
wire v_47040;
wire v_47041;
wire v_47042;
wire v_47043;
wire v_47044;
wire v_47045;
wire v_47046;
wire v_47047;
wire v_47048;
wire v_47049;
wire v_47050;
wire v_47051;
wire v_47052;
wire v_47053;
wire v_47054;
wire v_47055;
wire v_47056;
wire v_47057;
wire v_47058;
wire v_47059;
wire v_47060;
wire v_47061;
wire v_47062;
wire v_47063;
wire v_47064;
wire v_47065;
wire v_47066;
wire v_47067;
wire v_47068;
wire v_47069;
wire v_47070;
wire v_47071;
wire v_47072;
wire v_47073;
wire v_47074;
wire v_47075;
wire v_47076;
wire v_47077;
wire v_47078;
wire v_47079;
wire v_47080;
wire v_47081;
wire v_47082;
wire v_47083;
wire v_47084;
wire v_47085;
wire v_47086;
wire v_47087;
wire v_47088;
wire v_47089;
wire v_47090;
wire v_47091;
wire v_47092;
wire v_47093;
wire v_47094;
wire v_47095;
wire v_47096;
wire v_47097;
wire v_47098;
wire v_47099;
wire v_47100;
wire v_47101;
wire v_47102;
wire v_47103;
wire v_47104;
wire v_47105;
wire v_47106;
wire v_47107;
wire v_47108;
wire v_47109;
wire v_47110;
wire v_47111;
wire v_47112;
wire v_47113;
wire v_47114;
wire v_47115;
wire v_47116;
wire v_47117;
wire v_47118;
wire v_47119;
wire v_47120;
wire v_47121;
wire v_47122;
wire v_47123;
wire v_47124;
wire v_47125;
wire v_47126;
wire v_47127;
wire v_47128;
wire v_47129;
wire v_47130;
wire v_47131;
wire v_47132;
wire v_47133;
wire v_47134;
wire v_47135;
wire v_47136;
wire v_47137;
wire v_47138;
wire v_47139;
wire v_47140;
wire v_47141;
wire v_47142;
wire v_47143;
wire v_47144;
wire v_47145;
wire v_47146;
wire v_47147;
wire v_47148;
wire v_47149;
wire v_47150;
wire v_47151;
wire v_47152;
wire v_47153;
wire v_47155;
wire v_47156;
wire v_47157;
wire v_47158;
wire v_47159;
wire v_47160;
wire v_47161;
wire v_47162;
wire v_47163;
wire v_47164;
wire v_47165;
wire v_47166;
wire v_47167;
wire v_47168;
wire v_47169;
wire v_47170;
wire v_47171;
wire v_47172;
wire v_47173;
wire v_47174;
wire v_47175;
wire v_47176;
wire v_47177;
wire v_47178;
wire v_47179;
wire v_47180;
wire v_47181;
wire v_47182;
wire v_47183;
wire v_47184;
wire v_47185;
wire v_47186;
wire v_47187;
wire v_47188;
wire v_47189;
wire v_47190;
wire v_47191;
wire v_47192;
wire v_47193;
wire v_47194;
wire v_47195;
wire v_47196;
wire v_47197;
wire v_47198;
wire v_47199;
wire v_47200;
wire v_47201;
wire v_47202;
wire v_47203;
wire v_47204;
wire v_47205;
wire v_47206;
wire v_47207;
wire v_47208;
wire v_47209;
wire v_47210;
wire v_47211;
wire v_47212;
wire v_47213;
wire v_47214;
wire v_47215;
wire v_47216;
wire v_47217;
wire v_47218;
wire v_47219;
wire v_47220;
wire v_47221;
wire v_47222;
wire v_47223;
wire v_47224;
wire v_47225;
wire v_47226;
wire v_47227;
wire v_47228;
wire v_47229;
wire v_47230;
wire v_47231;
wire v_47232;
wire v_47233;
wire v_47234;
wire v_47235;
wire v_47236;
wire v_47237;
wire v_47238;
wire v_47239;
wire v_47240;
wire v_47241;
wire v_47242;
wire v_47243;
wire v_47244;
wire v_47245;
wire v_47246;
wire v_47247;
wire v_47248;
wire v_47249;
wire v_47250;
wire v_47251;
wire v_47252;
wire v_47253;
wire v_47254;
wire v_47255;
wire v_47256;
wire v_47257;
wire v_47258;
wire v_47259;
wire v_47260;
wire v_47261;
wire v_47262;
wire v_47263;
wire v_47264;
wire v_47265;
wire v_47266;
wire v_47267;
wire v_47268;
wire v_47269;
wire v_47270;
wire v_47271;
wire v_47272;
wire v_47273;
wire v_47274;
wire v_47275;
wire v_47276;
wire v_47277;
wire v_47278;
wire v_47279;
wire v_47280;
wire v_47281;
wire v_47282;
wire v_47283;
wire v_47284;
wire v_47285;
wire v_47286;
wire v_47287;
wire v_47288;
wire v_47289;
wire v_47290;
wire v_47291;
wire v_47292;
wire v_47293;
wire v_47294;
wire v_47295;
wire v_47296;
wire v_47297;
wire v_47298;
wire v_47299;
wire v_47300;
wire v_47301;
wire v_47302;
wire v_47303;
wire v_47304;
wire v_47305;
wire v_47306;
wire v_47307;
wire v_47308;
wire v_47309;
wire v_47310;
wire v_47311;
wire v_47312;
wire v_47313;
wire v_47314;
wire v_47315;
wire v_47316;
wire v_47317;
wire v_47318;
wire v_47319;
wire v_47320;
wire v_47321;
wire v_47322;
wire v_47323;
wire v_47324;
wire v_47325;
wire v_47326;
wire v_47327;
wire v_47328;
wire v_47329;
wire v_47330;
wire v_47331;
wire v_47332;
wire v_47333;
wire v_47334;
wire v_47335;
wire v_47336;
wire v_47337;
wire v_47338;
wire v_47339;
wire v_47340;
wire v_47341;
wire v_47342;
wire v_47343;
wire v_47344;
wire v_47345;
wire v_47346;
wire v_47347;
wire v_47348;
wire v_47349;
wire v_47350;
wire v_47351;
wire v_47352;
wire v_47353;
wire v_47354;
wire v_47355;
wire v_47356;
wire v_47357;
wire v_47358;
wire v_47359;
wire v_47360;
wire v_47361;
wire v_47362;
wire v_47363;
wire v_47364;
wire v_47365;
wire v_47366;
wire v_47367;
wire v_47368;
wire v_47369;
wire v_47370;
wire v_47371;
wire v_47372;
wire v_47373;
wire v_47374;
wire v_47375;
wire v_47376;
wire v_47377;
wire v_47378;
wire v_47379;
wire v_47380;
wire v_47381;
wire v_47382;
wire v_47383;
wire v_47384;
wire v_47385;
wire v_47386;
wire v_47387;
wire v_47388;
wire v_47389;
wire v_47390;
wire v_47391;
wire v_47392;
wire v_47393;
wire v_47394;
wire v_47395;
wire v_47396;
wire v_47398;
wire v_47399;
wire v_47400;
wire v_47401;
wire v_47402;
wire v_47403;
wire v_47404;
wire v_47405;
wire v_47406;
wire v_47407;
wire v_47408;
wire v_47409;
wire v_47410;
wire v_47411;
wire v_47412;
wire v_47413;
wire v_47414;
wire v_47415;
wire v_47416;
wire v_47417;
wire v_47418;
wire v_47419;
wire v_47420;
wire v_47421;
wire v_47422;
wire v_47423;
wire v_47424;
wire v_47425;
wire v_47426;
wire v_47427;
wire v_47428;
wire v_47429;
wire v_47430;
wire v_47431;
wire v_47432;
wire v_47433;
wire v_47434;
wire v_47435;
wire v_47436;
wire v_47437;
wire v_47438;
wire v_47439;
wire v_47440;
wire v_47441;
wire v_47442;
wire v_47443;
wire v_47444;
wire v_47445;
wire v_47446;
wire v_47447;
wire v_47448;
wire v_47449;
wire v_47450;
wire v_47451;
wire v_47452;
wire v_47453;
wire v_47454;
wire v_47455;
wire v_47456;
wire v_47457;
wire v_47458;
wire v_47459;
wire v_47460;
wire v_47461;
wire v_47462;
wire v_47463;
wire v_47464;
wire v_47465;
wire v_47466;
wire v_47467;
wire v_47468;
wire v_47469;
wire v_47470;
wire v_47471;
wire v_47472;
wire v_47473;
wire v_47474;
wire v_47475;
wire v_47476;
wire v_47477;
wire v_47478;
wire v_47479;
wire v_47480;
wire v_47481;
wire v_47482;
wire v_47483;
wire v_47484;
wire v_47485;
wire v_47486;
wire v_47487;
wire v_47488;
wire v_47489;
wire v_47490;
wire v_47491;
wire v_47492;
wire v_47493;
wire v_47494;
wire v_47495;
wire v_47496;
wire v_47497;
wire v_47498;
wire v_47499;
wire v_47500;
wire v_47501;
wire v_47502;
wire v_47503;
wire v_47504;
wire v_47505;
wire v_47506;
wire v_47507;
wire v_47508;
wire v_47509;
wire v_47510;
wire v_47511;
wire v_47512;
wire v_47513;
wire v_47514;
wire v_47515;
wire v_47516;
wire v_47517;
wire v_47518;
wire v_47519;
wire v_47520;
wire v_47521;
wire v_47522;
wire v_47523;
wire v_47524;
wire v_47525;
wire v_47526;
wire v_47527;
wire v_47528;
wire v_47529;
wire v_47530;
wire v_47531;
wire v_47532;
wire v_47533;
wire v_47534;
wire v_47535;
wire v_47536;
wire v_47537;
wire v_47538;
wire v_47539;
wire v_47540;
wire v_47541;
wire v_47542;
wire v_47543;
wire v_47544;
wire v_47545;
wire v_47546;
wire v_47547;
wire v_47548;
wire v_47549;
wire v_47550;
wire v_47551;
wire v_47552;
wire v_47553;
wire v_47554;
wire v_47555;
wire v_47556;
wire v_47557;
wire v_47558;
wire v_47559;
wire v_47560;
wire v_47561;
wire v_47562;
wire v_47563;
wire v_47564;
wire v_47565;
wire v_47566;
wire v_47567;
wire v_47568;
wire v_47569;
wire v_47570;
wire v_47571;
wire v_47572;
wire v_47573;
wire v_47574;
wire v_47575;
wire v_47576;
wire v_47577;
wire v_47578;
wire v_47579;
wire v_47580;
wire v_47581;
wire v_47582;
wire v_47583;
wire v_47584;
wire v_47585;
wire v_47586;
wire v_47587;
wire v_47588;
wire v_47589;
wire v_47590;
wire v_47591;
wire v_47592;
wire v_47593;
wire v_47594;
wire v_47595;
wire v_47596;
wire v_47597;
wire v_47598;
wire v_47599;
wire v_47600;
wire v_47601;
wire v_47602;
wire v_47603;
wire v_47604;
wire v_47605;
wire v_47606;
wire v_47607;
wire v_47608;
wire v_47609;
wire v_47610;
wire v_47611;
wire v_47612;
wire v_47613;
wire v_47614;
wire v_47615;
wire v_47616;
wire v_47617;
wire v_47618;
wire v_47619;
wire v_47620;
wire v_47621;
wire v_47622;
wire v_47623;
wire v_47624;
wire v_47625;
wire v_47626;
wire v_47627;
wire v_47628;
wire v_47629;
wire v_47630;
wire v_47631;
wire v_47632;
wire v_47633;
wire v_47634;
wire v_47635;
wire v_47636;
wire v_47637;
wire v_47638;
wire v_47639;
wire v_47641;
wire v_47642;
wire v_47643;
wire v_47644;
wire v_47645;
wire v_47646;
wire v_47647;
wire v_47648;
wire v_47649;
wire v_47650;
wire v_47651;
wire v_47652;
wire v_47653;
wire v_47654;
wire v_47655;
wire v_47656;
wire v_47657;
wire v_47658;
wire v_47659;
wire v_47660;
wire v_47661;
wire v_47662;
wire v_47663;
wire v_47664;
wire v_47665;
wire v_47666;
wire v_47667;
wire v_47668;
wire v_47669;
wire v_47670;
wire v_47671;
wire v_47672;
wire v_47673;
wire v_47674;
wire v_47675;
wire v_47676;
wire v_47677;
wire v_47678;
wire v_47679;
wire v_47680;
wire v_47681;
wire v_47682;
wire v_47683;
wire v_47684;
wire v_47685;
wire v_47686;
wire v_47687;
wire v_47688;
wire v_47689;
wire v_47690;
wire v_47691;
wire v_47692;
wire v_47693;
wire v_47694;
wire v_47695;
wire v_47696;
wire v_47697;
wire v_47698;
wire v_47699;
wire v_47700;
wire v_47701;
wire v_47702;
wire v_47703;
wire v_47704;
wire v_47705;
wire v_47706;
wire v_47707;
wire v_47708;
wire v_47709;
wire v_47710;
wire v_47711;
wire v_47712;
wire v_47713;
wire v_47714;
wire v_47715;
wire v_47716;
wire v_47717;
wire v_47718;
wire v_47719;
wire v_47720;
wire v_47721;
wire v_47722;
wire v_47723;
wire v_47724;
wire v_47725;
wire v_47726;
wire v_47727;
wire v_47728;
wire v_47729;
wire v_47730;
wire v_47731;
wire v_47732;
wire v_47733;
wire v_47734;
wire v_47735;
wire v_47736;
wire v_47737;
wire v_47738;
wire v_47739;
wire v_47740;
wire v_47741;
wire v_47742;
wire v_47743;
wire v_47744;
wire v_47745;
wire v_47746;
wire v_47747;
wire v_47748;
wire v_47749;
wire v_47750;
wire v_47751;
wire v_47752;
wire v_47753;
wire v_47754;
wire v_47755;
wire v_47756;
wire v_47757;
wire v_47758;
wire v_47759;
wire v_47760;
wire v_47761;
wire v_47762;
wire v_47763;
wire v_47764;
wire v_47765;
wire v_47766;
wire v_47767;
wire v_47768;
wire v_47769;
wire v_47770;
wire v_47771;
wire v_47772;
wire v_47773;
wire v_47774;
wire v_47775;
wire v_47776;
wire v_47777;
wire v_47778;
wire v_47779;
wire v_47780;
wire v_47781;
wire v_47782;
wire v_47783;
wire v_47784;
wire v_47785;
wire v_47786;
wire v_47787;
wire v_47788;
wire v_47789;
wire v_47790;
wire v_47791;
wire v_47792;
wire v_47793;
wire v_47794;
wire v_47795;
wire v_47796;
wire v_47797;
wire v_47798;
wire v_47799;
wire v_47800;
wire v_47801;
wire v_47802;
wire v_47803;
wire v_47804;
wire v_47805;
wire v_47806;
wire v_47807;
wire v_47808;
wire v_47809;
wire v_47810;
wire v_47811;
wire v_47812;
wire v_47813;
wire v_47814;
wire v_47815;
wire v_47816;
wire v_47817;
wire v_47818;
wire v_47819;
wire v_47820;
wire v_47821;
wire v_47822;
wire v_47823;
wire v_47824;
wire v_47825;
wire v_47826;
wire v_47827;
wire v_47828;
wire v_47829;
wire v_47830;
wire v_47831;
wire v_47832;
wire v_47833;
wire v_47834;
wire v_47835;
wire v_47836;
wire v_47837;
wire v_47838;
wire v_47839;
wire v_47840;
wire v_47841;
wire v_47842;
wire v_47843;
wire v_47844;
wire v_47845;
wire v_47846;
wire v_47847;
wire v_47848;
wire v_47849;
wire v_47850;
wire v_47851;
wire v_47852;
wire v_47853;
wire v_47854;
wire v_47855;
wire v_47856;
wire v_47857;
wire v_47858;
wire v_47859;
wire v_47860;
wire v_47861;
wire v_47862;
wire v_47863;
wire v_47864;
wire v_47865;
wire v_47866;
wire v_47867;
wire v_47868;
wire v_47869;
wire v_47870;
wire v_47871;
wire v_47872;
wire v_47873;
wire v_47874;
wire v_47875;
wire v_47876;
wire v_47877;
wire v_47878;
wire v_47879;
wire v_47880;
wire v_47881;
wire v_47882;
wire v_47884;
wire v_47885;
wire v_47886;
wire v_47887;
wire v_47888;
wire v_47889;
wire v_47890;
wire v_47891;
wire v_47892;
wire v_47893;
wire v_47894;
wire v_47895;
wire v_47896;
wire v_47897;
wire v_47898;
wire v_47899;
wire v_47900;
wire v_47901;
wire v_47902;
wire v_47903;
wire v_47904;
wire v_47905;
wire v_47906;
wire v_47907;
wire v_47908;
wire v_47909;
wire v_47910;
wire v_47911;
wire v_47912;
wire v_47913;
wire v_47914;
wire v_47915;
wire v_47916;
wire v_47917;
wire v_47918;
wire v_47919;
wire v_47920;
wire v_47921;
wire v_47922;
wire v_47923;
wire v_47924;
wire v_47925;
wire v_47926;
wire v_47927;
wire v_47928;
wire v_47929;
wire v_47930;
wire v_47931;
wire v_47932;
wire v_47933;
wire v_47934;
wire v_47935;
wire v_47936;
wire v_47937;
wire v_47938;
wire v_47939;
wire v_47940;
wire v_47941;
wire v_47942;
wire v_47943;
wire v_47944;
wire v_47945;
wire v_47946;
wire v_47947;
wire v_47948;
wire v_47949;
wire v_47950;
wire v_47951;
wire v_47952;
wire v_47953;
wire v_47954;
wire v_47955;
wire v_47956;
wire v_47957;
wire v_47958;
wire v_47959;
wire v_47960;
wire v_47961;
wire v_47962;
wire v_47963;
wire v_47964;
wire v_47965;
wire v_47966;
wire v_47967;
wire v_47968;
wire v_47969;
wire v_47970;
wire v_47971;
wire v_47972;
wire v_47973;
wire v_47974;
wire v_47975;
wire v_47976;
wire v_47977;
wire v_47978;
wire v_47979;
wire v_47980;
wire v_47981;
wire v_47982;
wire v_47983;
wire v_47984;
wire v_47985;
wire v_47986;
wire v_47987;
wire v_47988;
wire v_47989;
wire v_47990;
wire v_47991;
wire v_47992;
wire v_47993;
wire v_47994;
wire v_47995;
wire v_47996;
wire v_47997;
wire v_47998;
wire v_47999;
wire v_48000;
wire v_48001;
wire v_48002;
wire v_48003;
wire v_48004;
wire v_48005;
wire v_48006;
wire v_48007;
wire v_48008;
wire v_48009;
wire v_48010;
wire v_48011;
wire v_48012;
wire v_48013;
wire v_48014;
wire v_48015;
wire v_48016;
wire v_48017;
wire v_48018;
wire v_48019;
wire v_48020;
wire v_48021;
wire v_48022;
wire v_48023;
wire v_48024;
wire v_48025;
wire v_48026;
wire v_48027;
wire v_48028;
wire v_48029;
wire v_48030;
wire v_48031;
wire v_48032;
wire v_48033;
wire v_48034;
wire v_48035;
wire v_48036;
wire v_48037;
wire v_48038;
wire v_48039;
wire v_48040;
wire v_48041;
wire v_48042;
wire v_48043;
wire v_48044;
wire v_48045;
wire v_48046;
wire v_48047;
wire v_48048;
wire v_48049;
wire v_48050;
wire v_48051;
wire v_48052;
wire v_48053;
wire v_48054;
wire v_48055;
wire v_48056;
wire v_48057;
wire v_48058;
wire v_48059;
wire v_48060;
wire v_48061;
wire v_48062;
wire v_48063;
wire v_48064;
wire v_48065;
wire v_48066;
wire v_48067;
wire v_48068;
wire v_48069;
wire v_48070;
wire v_48071;
wire v_48072;
wire v_48073;
wire v_48074;
wire v_48075;
wire v_48076;
wire v_48077;
wire v_48078;
wire v_48079;
wire v_48080;
wire v_48081;
wire v_48082;
wire v_48083;
wire v_48084;
wire v_48085;
wire v_48086;
wire v_48087;
wire v_48088;
wire v_48089;
wire v_48090;
wire v_48091;
wire v_48092;
wire v_48093;
wire v_48094;
wire v_48095;
wire v_48096;
wire v_48097;
wire v_48098;
wire v_48099;
wire v_48100;
wire v_48101;
wire v_48102;
wire v_48103;
wire v_48104;
wire v_48105;
wire v_48106;
wire v_48107;
wire v_48108;
wire v_48109;
wire v_48110;
wire v_48111;
wire v_48112;
wire v_48113;
wire v_48114;
wire v_48115;
wire v_48116;
wire v_48117;
wire v_48118;
wire v_48119;
wire v_48120;
wire v_48121;
wire v_48122;
wire v_48123;
wire v_48124;
wire v_48125;
wire v_48127;
wire v_48128;
wire v_48129;
wire v_48130;
wire v_48131;
wire v_48132;
wire v_48133;
wire v_48134;
wire v_48135;
wire v_48136;
wire v_48137;
wire v_48138;
wire v_48139;
wire v_48140;
wire v_48141;
wire v_48142;
wire v_48143;
wire v_48144;
wire v_48145;
wire v_48146;
wire v_48147;
wire v_48148;
wire v_48149;
wire v_48150;
wire v_48151;
wire v_48152;
wire v_48153;
wire v_48154;
wire v_48155;
wire v_48156;
wire v_48157;
wire v_48158;
wire v_48159;
wire v_48160;
wire v_48161;
wire v_48162;
wire v_48163;
wire v_48164;
wire v_48165;
wire v_48166;
wire v_48167;
wire v_48168;
wire v_48169;
wire v_48170;
wire v_48171;
wire v_48172;
wire v_48173;
wire v_48174;
wire v_48175;
wire v_48176;
wire v_48177;
wire v_48178;
wire v_48179;
wire v_48180;
wire v_48181;
wire v_48182;
wire v_48183;
wire v_48184;
wire v_48185;
wire v_48186;
wire v_48187;
wire v_48188;
wire v_48189;
wire v_48190;
wire v_48191;
wire v_48192;
wire v_48193;
wire v_48194;
wire v_48195;
wire v_48196;
wire v_48197;
wire v_48198;
wire v_48199;
wire v_48200;
wire v_48201;
wire v_48202;
wire v_48203;
wire v_48204;
wire v_48205;
wire v_48206;
wire v_48207;
wire v_48208;
wire v_48209;
wire v_48210;
wire v_48211;
wire v_48212;
wire v_48213;
wire v_48214;
wire v_48215;
wire v_48216;
wire v_48217;
wire v_48218;
wire v_48219;
wire v_48220;
wire v_48221;
wire v_48222;
wire v_48223;
wire v_48224;
wire v_48225;
wire v_48226;
wire v_48227;
wire v_48228;
wire v_48229;
wire v_48230;
wire v_48231;
wire v_48232;
wire v_48233;
wire v_48234;
wire v_48235;
wire v_48236;
wire v_48237;
wire v_48238;
wire v_48239;
wire v_48240;
wire v_48241;
wire v_48242;
wire v_48243;
wire v_48244;
wire v_48245;
wire v_48246;
wire v_48247;
wire v_48248;
wire v_48249;
wire v_48250;
wire v_48251;
wire v_48252;
wire v_48253;
wire v_48254;
wire v_48255;
wire v_48256;
wire v_48257;
wire v_48258;
wire v_48259;
wire v_48260;
wire v_48261;
wire v_48262;
wire v_48263;
wire v_48264;
wire v_48265;
wire v_48266;
wire v_48267;
wire v_48268;
wire v_48269;
wire v_48270;
wire v_48271;
wire v_48272;
wire v_48273;
wire v_48274;
wire v_48275;
wire v_48276;
wire v_48277;
wire v_48278;
wire v_48279;
wire v_48280;
wire v_48281;
wire v_48282;
wire v_48283;
wire v_48284;
wire v_48285;
wire v_48286;
wire v_48287;
wire v_48288;
wire v_48289;
wire v_48290;
wire v_48291;
wire v_48292;
wire v_48293;
wire v_48294;
wire v_48295;
wire v_48296;
wire v_48297;
wire v_48298;
wire v_48299;
wire v_48300;
wire v_48301;
wire v_48302;
wire v_48303;
wire v_48304;
wire v_48305;
wire v_48306;
wire v_48307;
wire v_48308;
wire v_48309;
wire v_48310;
wire v_48311;
wire v_48312;
wire v_48313;
wire v_48314;
wire v_48315;
wire v_48316;
wire v_48317;
wire v_48318;
wire v_48319;
wire v_48320;
wire v_48321;
wire v_48322;
wire v_48323;
wire v_48324;
wire v_48325;
wire v_48326;
wire v_48327;
wire v_48328;
wire v_48329;
wire v_48330;
wire v_48331;
wire v_48332;
wire v_48333;
wire v_48334;
wire v_48335;
wire v_48336;
wire v_48337;
wire v_48338;
wire v_48339;
wire v_48340;
wire v_48341;
wire v_48342;
wire v_48343;
wire v_48344;
wire v_48345;
wire v_48346;
wire v_48347;
wire v_48348;
wire v_48349;
wire v_48350;
wire v_48351;
wire v_48352;
wire v_48353;
wire v_48354;
wire v_48355;
wire v_48356;
wire v_48357;
wire v_48358;
wire v_48359;
wire v_48360;
wire v_48361;
wire v_48362;
wire v_48363;
wire v_48364;
wire v_48365;
wire v_48366;
wire v_48367;
wire v_48368;
wire v_48370;
wire v_48371;
wire v_48372;
wire v_48373;
wire v_48374;
wire v_48375;
wire v_48376;
wire v_48377;
wire v_48378;
wire v_48379;
wire v_48380;
wire v_48381;
wire v_48382;
wire v_48383;
wire v_48384;
wire v_48385;
wire v_48386;
wire v_48387;
wire v_48388;
wire v_48389;
wire v_48390;
wire v_48391;
wire v_48392;
wire v_48393;
wire v_48394;
wire v_48395;
wire v_48396;
wire v_48397;
wire v_48398;
wire v_48399;
wire v_48400;
wire v_48401;
wire v_48402;
wire v_48403;
wire v_48404;
wire v_48405;
wire v_48406;
wire v_48407;
wire v_48408;
wire v_48409;
wire v_48410;
wire v_48411;
wire v_48412;
wire v_48413;
wire v_48414;
wire v_48415;
wire v_48416;
wire v_48417;
wire v_48418;
wire v_48419;
wire v_48420;
wire v_48421;
wire v_48422;
wire v_48423;
wire v_48424;
wire v_48425;
wire v_48426;
wire v_48427;
wire v_48428;
wire v_48429;
wire v_48430;
wire v_48431;
wire v_48432;
wire v_48433;
wire v_48434;
wire v_48435;
wire v_48436;
wire v_48437;
wire v_48438;
wire v_48439;
wire v_48440;
wire v_48441;
wire v_48442;
wire v_48443;
wire v_48444;
wire v_48445;
wire v_48446;
wire v_48447;
wire v_48448;
wire v_48449;
wire v_48450;
wire v_48451;
wire v_48452;
wire v_48453;
wire v_48454;
wire v_48455;
wire v_48456;
wire v_48457;
wire v_48458;
wire v_48459;
wire v_48460;
wire v_48461;
wire v_48462;
wire v_48463;
wire v_48464;
wire v_48465;
wire v_48466;
wire v_48467;
wire v_48468;
wire v_48469;
wire v_48470;
wire v_48471;
wire v_48472;
wire v_48473;
wire v_48474;
wire v_48475;
wire v_48476;
wire v_48477;
wire v_48478;
wire v_48479;
wire v_48480;
wire v_48481;
wire v_48482;
wire v_48483;
wire v_48484;
wire v_48485;
wire v_48486;
wire v_48487;
wire v_48488;
wire v_48489;
wire v_48490;
wire v_48491;
wire v_48492;
wire v_48493;
wire v_48494;
wire v_48495;
wire v_48496;
wire v_48497;
wire v_48498;
wire v_48499;
wire v_48500;
wire v_48501;
wire v_48502;
wire v_48503;
wire v_48504;
wire v_48505;
wire v_48506;
wire v_48507;
wire v_48508;
wire v_48509;
wire v_48510;
wire v_48511;
wire v_48512;
wire v_48513;
wire v_48514;
wire v_48515;
wire v_48516;
wire v_48517;
wire v_48518;
wire v_48519;
wire v_48520;
wire v_48521;
wire v_48522;
wire v_48523;
wire v_48524;
wire v_48525;
wire v_48526;
wire v_48527;
wire v_48528;
wire v_48529;
wire v_48530;
wire v_48531;
wire v_48532;
wire v_48533;
wire v_48534;
wire v_48535;
wire v_48536;
wire v_48537;
wire v_48538;
wire v_48539;
wire v_48540;
wire v_48541;
wire v_48542;
wire v_48543;
wire v_48544;
wire v_48545;
wire v_48546;
wire v_48547;
wire v_48548;
wire v_48549;
wire v_48550;
wire v_48551;
wire v_48552;
wire v_48553;
wire v_48554;
wire v_48555;
wire v_48556;
wire v_48557;
wire v_48558;
wire v_48559;
wire v_48560;
wire v_48561;
wire v_48562;
wire v_48563;
wire v_48564;
wire v_48565;
wire v_48566;
wire v_48567;
wire v_48568;
wire v_48569;
wire v_48570;
wire v_48571;
wire v_48572;
wire v_48573;
wire v_48574;
wire v_48575;
wire v_48576;
wire v_48577;
wire v_48578;
wire v_48579;
wire v_48580;
wire v_48581;
wire v_48582;
wire v_48583;
wire v_48584;
wire v_48585;
wire v_48586;
wire v_48587;
wire v_48588;
wire v_48589;
wire v_48590;
wire v_48591;
wire v_48592;
wire v_48593;
wire v_48594;
wire v_48595;
wire v_48596;
wire v_48597;
wire v_48598;
wire v_48599;
wire v_48600;
wire v_48601;
wire v_48602;
wire v_48603;
wire v_48604;
wire v_48605;
wire v_48606;
wire v_48607;
wire v_48608;
wire v_48609;
wire v_48610;
wire v_48611;
wire v_48613;
wire v_48614;
wire v_48615;
wire v_48616;
wire v_48617;
wire v_48618;
wire v_48619;
wire v_48620;
wire v_48621;
wire v_48622;
wire v_48623;
wire v_48624;
wire v_48625;
wire v_48626;
wire v_48627;
wire v_48628;
wire v_48629;
wire v_48630;
wire v_48631;
wire v_48632;
wire v_48633;
wire v_48634;
wire v_48635;
wire v_48636;
wire v_48637;
wire v_48638;
wire v_48639;
wire v_48640;
wire v_48641;
wire v_48642;
wire v_48643;
wire v_48644;
wire v_48645;
wire v_48646;
wire v_48647;
wire v_48648;
wire v_48649;
wire v_48650;
wire v_48651;
wire v_48652;
wire v_48653;
wire v_48654;
wire v_48655;
wire v_48656;
wire v_48657;
wire v_48658;
wire v_48659;
wire v_48660;
wire v_48661;
wire v_48662;
wire v_48663;
wire v_48664;
wire v_48665;
wire v_48666;
wire v_48667;
wire v_48668;
wire v_48669;
wire v_48670;
wire v_48671;
wire v_48672;
wire v_48673;
wire v_48674;
wire v_48675;
wire v_48676;
wire v_48677;
wire v_48678;
wire v_48679;
wire v_48680;
wire v_48681;
wire v_48682;
wire v_48683;
wire v_48684;
wire v_48685;
wire v_48686;
wire v_48687;
wire v_48688;
wire v_48689;
wire v_48690;
wire v_48691;
wire v_48692;
wire v_48693;
wire v_48694;
wire v_48695;
wire v_48696;
wire v_48697;
wire v_48698;
wire v_48699;
wire v_48700;
wire v_48701;
wire v_48702;
wire v_48703;
wire v_48704;
wire v_48705;
wire v_48706;
wire v_48707;
wire v_48708;
wire v_48709;
wire v_48710;
wire v_48711;
wire v_48712;
wire v_48713;
wire v_48714;
wire v_48715;
wire v_48716;
wire v_48717;
wire v_48718;
wire v_48719;
wire v_48720;
wire v_48721;
wire v_48722;
wire v_48723;
wire v_48724;
wire v_48725;
wire v_48726;
wire v_48727;
wire v_48728;
wire v_48729;
wire v_48730;
wire v_48731;
wire v_48732;
wire v_48733;
wire v_48734;
wire v_48735;
wire v_48736;
wire v_48737;
wire v_48738;
wire v_48739;
wire v_48740;
wire v_48741;
wire v_48742;
wire v_48743;
wire v_48744;
wire v_48745;
wire v_48746;
wire v_48747;
wire v_48748;
wire v_48749;
wire v_48750;
wire v_48751;
wire v_48752;
wire v_48753;
wire v_48754;
wire v_48755;
wire v_48756;
wire v_48757;
wire v_48758;
wire v_48759;
wire v_48760;
wire v_48761;
wire v_48762;
wire v_48763;
wire v_48764;
wire v_48765;
wire v_48766;
wire v_48767;
wire v_48768;
wire v_48769;
wire v_48770;
wire v_48771;
wire v_48772;
wire v_48773;
wire v_48774;
wire v_48775;
wire v_48776;
wire v_48777;
wire v_48778;
wire v_48779;
wire v_48780;
wire v_48781;
wire v_48782;
wire v_48783;
wire v_48784;
wire v_48785;
wire v_48786;
wire v_48787;
wire v_48788;
wire v_48789;
wire v_48790;
wire v_48791;
wire v_48792;
wire v_48793;
wire v_48794;
wire v_48795;
wire v_48796;
wire v_48797;
wire v_48798;
wire v_48799;
wire v_48800;
wire v_48801;
wire v_48802;
wire v_48803;
wire v_48804;
wire v_48805;
wire v_48806;
wire v_48807;
wire v_48808;
wire v_48809;
wire v_48810;
wire v_48811;
wire v_48812;
wire v_48813;
wire v_48814;
wire v_48815;
wire v_48816;
wire v_48817;
wire v_48818;
wire v_48819;
wire v_48820;
wire v_48821;
wire v_48822;
wire v_48823;
wire v_48824;
wire v_48825;
wire v_48826;
wire v_48827;
wire v_48828;
wire v_48829;
wire v_48830;
wire v_48831;
wire v_48832;
wire v_48833;
wire v_48834;
wire v_48835;
wire v_48836;
wire v_48837;
wire v_48838;
wire v_48839;
wire v_48840;
wire v_48841;
wire v_48842;
wire v_48843;
wire v_48844;
wire v_48845;
wire v_48846;
wire v_48847;
wire v_48848;
wire v_48849;
wire v_48850;
wire v_48851;
wire v_48852;
wire v_48853;
wire v_48854;
wire v_48856;
wire v_48857;
wire v_48858;
wire v_48859;
wire v_48860;
wire v_48861;
wire v_48862;
wire v_48863;
wire v_48864;
wire v_48865;
wire v_48866;
wire v_48867;
wire v_48868;
wire v_48869;
wire v_48870;
wire v_48871;
wire v_48872;
wire v_48873;
wire v_48874;
wire v_48875;
wire v_48876;
wire v_48877;
wire v_48878;
wire v_48879;
wire v_48880;
wire v_48881;
wire v_48882;
wire v_48883;
wire v_48884;
wire v_48885;
wire v_48886;
wire v_48887;
wire v_48888;
wire v_48889;
wire v_48890;
wire v_48891;
wire v_48892;
wire v_48893;
wire v_48894;
wire v_48895;
wire v_48896;
wire v_48897;
wire v_48898;
wire v_48899;
wire v_48900;
wire v_48901;
wire v_48902;
wire v_48903;
wire v_48904;
wire v_48905;
wire v_48906;
wire v_48907;
wire v_48908;
wire v_48909;
wire v_48910;
wire v_48911;
wire v_48912;
wire v_48913;
wire v_48914;
wire v_48915;
wire v_48916;
wire v_48917;
wire v_48918;
wire v_48919;
wire v_48920;
wire v_48921;
wire v_48922;
wire v_48923;
wire v_48924;
wire v_48925;
wire v_48926;
wire v_48927;
wire v_48928;
wire v_48929;
wire v_48930;
wire v_48931;
wire v_48932;
wire v_48933;
wire v_48934;
wire v_48935;
wire v_48936;
wire v_48937;
wire v_48938;
wire v_48939;
wire v_48940;
wire v_48941;
wire v_48942;
wire v_48943;
wire v_48944;
wire v_48945;
wire v_48946;
wire v_48947;
wire v_48948;
wire v_48949;
wire v_48950;
wire v_48951;
wire v_48952;
wire v_48953;
wire v_48954;
wire v_48955;
wire v_48956;
wire v_48957;
wire v_48958;
wire v_48959;
wire v_48960;
wire v_48961;
wire v_48962;
wire v_48963;
wire v_48964;
wire v_48965;
wire v_48966;
wire v_48967;
wire v_48968;
wire v_48969;
wire v_48970;
wire v_48971;
wire v_48972;
wire v_48973;
wire v_48974;
wire v_48975;
wire v_48976;
wire v_48977;
wire v_48978;
wire v_48979;
wire v_48980;
wire v_48981;
wire v_48982;
wire v_48983;
wire v_48984;
wire v_48985;
wire v_48986;
wire v_48987;
wire v_48988;
wire v_48989;
wire v_48990;
wire v_48991;
wire v_48992;
wire v_48993;
wire v_48994;
wire v_48995;
wire v_48996;
wire v_48997;
wire v_48998;
wire v_48999;
wire v_49000;
wire v_49001;
wire v_49002;
wire v_49003;
wire v_49004;
wire v_49005;
wire v_49006;
wire v_49007;
wire v_49008;
wire v_49009;
wire v_49010;
wire v_49011;
wire v_49012;
wire v_49013;
wire v_49014;
wire v_49015;
wire v_49016;
wire v_49017;
wire v_49018;
wire v_49019;
wire v_49020;
wire v_49021;
wire v_49022;
wire v_49023;
wire v_49024;
wire v_49025;
wire v_49026;
wire v_49027;
wire v_49028;
wire v_49029;
wire v_49030;
wire v_49031;
wire v_49032;
wire v_49033;
wire v_49034;
wire v_49035;
wire v_49036;
wire v_49037;
wire v_49038;
wire v_49039;
wire v_49040;
wire v_49041;
wire v_49042;
wire v_49043;
wire v_49044;
wire v_49045;
wire v_49046;
wire v_49047;
wire v_49048;
wire v_49049;
wire v_49050;
wire v_49051;
wire v_49052;
wire v_49053;
wire v_49054;
wire v_49055;
wire v_49056;
wire v_49057;
wire v_49058;
wire v_49059;
wire v_49060;
wire v_49061;
wire v_49062;
wire v_49063;
wire v_49064;
wire v_49065;
wire v_49066;
wire v_49067;
wire v_49068;
wire v_49069;
wire v_49070;
wire v_49071;
wire v_49072;
wire v_49073;
wire v_49074;
wire v_49075;
wire v_49076;
wire v_49077;
wire v_49078;
wire v_49079;
wire v_49080;
wire v_49081;
wire v_49082;
wire v_49083;
wire v_49084;
wire v_49085;
wire v_49086;
wire v_49087;
wire v_49088;
wire v_49089;
wire v_49090;
wire v_49091;
wire v_49092;
wire v_49093;
wire v_49094;
wire v_49095;
wire v_49096;
wire v_49097;
wire v_49099;
wire v_49100;
wire v_49101;
wire v_49102;
wire v_49103;
wire v_49104;
wire v_49105;
wire v_49106;
wire v_49107;
wire v_49108;
wire v_49109;
wire v_49110;
wire v_49111;
wire v_49112;
wire v_49113;
wire v_49114;
wire v_49115;
wire v_49116;
wire v_49117;
wire v_49118;
wire v_49119;
wire v_49120;
wire v_49121;
wire v_49122;
wire v_49123;
wire v_49124;
wire v_49125;
wire v_49126;
wire v_49127;
wire v_49128;
wire v_49129;
wire v_49130;
wire v_49131;
wire v_49132;
wire v_49133;
wire v_49134;
wire v_49135;
wire v_49136;
wire v_49137;
wire v_49138;
wire v_49139;
wire v_49140;
wire v_49141;
wire v_49142;
wire v_49143;
wire v_49144;
wire v_49145;
wire v_49146;
wire v_49147;
wire v_49148;
wire v_49149;
wire v_49150;
wire v_49151;
wire v_49152;
wire v_49153;
wire v_49154;
wire v_49155;
wire v_49156;
wire v_49157;
wire v_49158;
wire v_49159;
wire v_49160;
wire v_49161;
wire v_49162;
wire v_49163;
wire v_49164;
wire v_49165;
wire v_49166;
wire v_49167;
wire v_49168;
wire v_49169;
wire v_49170;
wire v_49171;
wire v_49172;
wire v_49173;
wire v_49174;
wire v_49175;
wire v_49176;
wire v_49177;
wire v_49178;
wire v_49179;
wire v_49180;
wire v_49181;
wire v_49182;
wire v_49183;
wire v_49184;
wire v_49185;
wire v_49186;
wire v_49187;
wire v_49188;
wire v_49189;
wire v_49190;
wire v_49191;
wire v_49192;
wire v_49193;
wire v_49194;
wire v_49195;
wire v_49196;
wire v_49197;
wire v_49198;
wire v_49199;
wire v_49200;
wire v_49201;
wire v_49202;
wire v_49203;
wire v_49204;
wire v_49205;
wire v_49206;
wire v_49207;
wire v_49208;
wire v_49209;
wire v_49210;
wire v_49211;
wire v_49212;
wire v_49213;
wire v_49214;
wire v_49215;
wire v_49216;
wire v_49217;
wire v_49218;
wire v_49219;
wire v_49220;
wire v_49221;
wire v_49222;
wire v_49223;
wire v_49224;
wire v_49225;
wire v_49226;
wire v_49227;
wire v_49228;
wire v_49229;
wire v_49230;
wire v_49231;
wire v_49232;
wire v_49233;
wire v_49234;
wire v_49235;
wire v_49236;
wire v_49237;
wire v_49238;
wire v_49239;
wire v_49240;
wire v_49241;
wire v_49242;
wire v_49243;
wire v_49244;
wire v_49245;
wire v_49246;
wire v_49247;
wire v_49248;
wire v_49249;
wire v_49250;
wire v_49251;
wire v_49252;
wire v_49253;
wire v_49254;
wire v_49255;
wire v_49256;
wire v_49257;
wire v_49258;
wire v_49259;
wire v_49260;
wire v_49261;
wire v_49262;
wire v_49263;
wire v_49264;
wire v_49265;
wire v_49266;
wire v_49267;
wire v_49268;
wire v_49269;
wire v_49270;
wire v_49271;
wire v_49272;
wire v_49273;
wire v_49274;
wire v_49275;
wire v_49276;
wire v_49277;
wire v_49278;
wire v_49279;
wire v_49280;
wire v_49281;
wire v_49282;
wire v_49283;
wire v_49284;
wire v_49285;
wire v_49286;
wire v_49287;
wire v_49288;
wire v_49289;
wire v_49290;
wire v_49291;
wire v_49292;
wire v_49293;
wire v_49294;
wire v_49295;
wire v_49296;
wire v_49297;
wire v_49298;
wire v_49299;
wire v_49300;
wire v_49301;
wire v_49302;
wire v_49303;
wire v_49304;
wire v_49305;
wire v_49306;
wire v_49307;
wire v_49308;
wire v_49309;
wire v_49310;
wire v_49311;
wire v_49312;
wire v_49313;
wire v_49314;
wire v_49315;
wire v_49316;
wire v_49317;
wire v_49318;
wire v_49319;
wire v_49320;
wire v_49321;
wire v_49322;
wire v_49323;
wire v_49324;
wire v_49325;
wire v_49326;
wire v_49327;
wire v_49328;
wire v_49329;
wire v_49330;
wire v_49331;
wire v_49332;
wire v_49333;
wire v_49334;
wire v_49335;
wire v_49336;
wire v_49337;
wire v_49338;
wire v_49339;
wire v_49340;
wire v_49342;
wire v_49343;
wire v_49344;
wire v_49345;
wire v_49346;
wire v_49347;
wire v_49348;
wire v_49349;
wire v_49350;
wire v_49351;
wire v_49352;
wire v_49353;
wire v_49354;
wire v_49355;
wire v_49356;
wire v_49357;
wire v_49358;
wire v_49359;
wire v_49360;
wire v_49361;
wire v_49362;
wire v_49363;
wire v_49364;
wire v_49365;
wire v_49366;
wire v_49367;
wire v_49368;
wire v_49369;
wire v_49370;
wire v_49371;
wire v_49372;
wire v_49373;
wire v_49374;
wire v_49375;
wire v_49376;
wire v_49377;
wire v_49378;
wire v_49379;
wire v_49380;
wire v_49381;
wire v_49382;
wire v_49383;
wire v_49384;
wire v_49385;
wire v_49386;
wire v_49387;
wire v_49388;
wire v_49389;
wire v_49390;
wire v_49391;
wire v_49392;
wire v_49393;
wire v_49394;
wire v_49395;
wire v_49396;
wire v_49397;
wire v_49398;
wire v_49399;
wire v_49400;
wire v_49401;
wire v_49402;
wire v_49403;
wire v_49404;
wire v_49405;
wire v_49406;
wire v_49407;
wire v_49408;
wire v_49409;
wire v_49410;
wire v_49411;
wire v_49412;
wire v_49413;
wire v_49414;
wire v_49415;
wire v_49416;
wire v_49417;
wire v_49418;
wire v_49419;
wire v_49420;
wire v_49421;
wire v_49422;
wire v_49423;
wire v_49424;
wire v_49425;
wire v_49426;
wire v_49427;
wire v_49428;
wire v_49429;
wire v_49430;
wire v_49431;
wire v_49432;
wire v_49433;
wire v_49434;
wire v_49435;
wire v_49436;
wire v_49437;
wire v_49438;
wire v_49439;
wire v_49440;
wire v_49441;
wire v_49442;
wire v_49443;
wire v_49444;
wire v_49445;
wire v_49446;
wire v_49447;
wire v_49448;
wire v_49449;
wire v_49450;
wire v_49451;
wire v_49452;
wire v_49453;
wire v_49454;
wire v_49455;
wire v_49456;
wire v_49457;
wire v_49458;
wire v_49459;
wire v_49460;
wire v_49461;
wire v_49462;
wire v_49463;
wire v_49464;
wire v_49465;
wire v_49466;
wire v_49467;
wire v_49468;
wire v_49469;
wire v_49470;
wire v_49471;
wire v_49472;
wire v_49473;
wire v_49474;
wire v_49475;
wire v_49476;
wire v_49477;
wire v_49478;
wire v_49479;
wire v_49480;
wire v_49481;
wire v_49482;
wire v_49483;
wire v_49484;
wire v_49485;
wire v_49486;
wire v_49487;
wire v_49488;
wire v_49489;
wire v_49490;
wire v_49491;
wire v_49492;
wire v_49493;
wire v_49494;
wire v_49495;
wire v_49496;
wire v_49497;
wire v_49498;
wire v_49499;
wire v_49500;
wire v_49501;
wire v_49502;
wire v_49503;
wire v_49504;
wire v_49505;
wire v_49506;
wire v_49507;
wire v_49508;
wire v_49509;
wire v_49510;
wire v_49511;
wire v_49512;
wire v_49513;
wire v_49514;
wire v_49515;
wire v_49516;
wire v_49517;
wire v_49518;
wire v_49519;
wire v_49520;
wire v_49521;
wire v_49522;
wire v_49523;
wire v_49524;
wire v_49525;
wire v_49526;
wire v_49527;
wire v_49528;
wire v_49529;
wire v_49530;
wire v_49531;
wire v_49532;
wire v_49533;
wire v_49534;
wire v_49535;
wire v_49536;
wire v_49537;
wire v_49538;
wire v_49539;
wire v_49540;
wire v_49541;
wire v_49542;
wire v_49543;
wire v_49544;
wire v_49545;
wire v_49546;
wire v_49547;
wire v_49548;
wire v_49549;
wire v_49550;
wire v_49551;
wire v_49552;
wire v_49553;
wire v_49554;
wire v_49555;
wire v_49556;
wire v_49557;
wire v_49558;
wire v_49559;
wire v_49560;
wire v_49561;
wire v_49562;
wire v_49563;
wire v_49564;
wire v_49565;
wire v_49566;
wire v_49567;
wire v_49568;
wire v_49569;
wire v_49570;
wire v_49571;
wire v_49572;
wire v_49573;
wire v_49574;
wire v_49575;
wire v_49576;
wire v_49577;
wire v_49578;
wire v_49579;
wire v_49580;
wire v_49581;
wire v_49582;
wire v_49583;
wire v_49585;
wire v_49586;
wire v_49587;
wire v_49588;
wire v_49589;
wire v_49590;
wire v_49591;
wire v_49592;
wire v_49593;
wire v_49594;
wire v_49595;
wire v_49596;
wire v_49597;
wire v_49598;
wire v_49599;
wire v_49600;
wire v_49601;
wire v_49602;
wire v_49603;
wire v_49604;
wire v_49605;
wire v_49606;
wire v_49607;
wire v_49608;
wire v_49609;
wire v_49610;
wire v_49611;
wire v_49612;
wire v_49613;
wire v_49614;
wire v_49615;
wire v_49616;
wire v_49617;
wire v_49618;
wire v_49619;
wire v_49620;
wire v_49621;
wire v_49622;
wire v_49623;
wire v_49624;
wire v_49625;
wire v_49626;
wire v_49627;
wire v_49628;
wire v_49629;
wire v_49630;
wire v_49631;
wire v_49632;
wire v_49633;
wire v_49634;
wire v_49635;
wire v_49636;
wire v_49637;
wire v_49638;
wire v_49639;
wire v_49640;
wire v_49641;
wire v_49642;
wire v_49643;
wire v_49644;
wire v_49645;
wire v_49646;
wire v_49647;
wire v_49648;
wire v_49649;
wire v_49650;
wire v_49651;
wire v_49652;
wire v_49653;
wire v_49654;
wire v_49655;
wire v_49656;
wire v_49657;
wire v_49658;
wire v_49659;
wire v_49660;
wire v_49661;
wire v_49662;
wire v_49663;
wire v_49664;
wire v_49665;
wire v_49666;
wire v_49667;
wire v_49668;
wire v_49669;
wire v_49670;
wire v_49671;
wire v_49672;
wire v_49673;
wire v_49674;
wire v_49675;
wire v_49676;
wire v_49677;
wire v_49678;
wire v_49679;
wire v_49680;
wire v_49681;
wire v_49682;
wire v_49683;
wire v_49684;
wire v_49685;
wire v_49686;
wire v_49687;
wire v_49688;
wire v_49689;
wire v_49690;
wire v_49691;
wire v_49692;
wire v_49693;
wire v_49694;
wire v_49695;
wire v_49696;
wire v_49697;
wire v_49698;
wire v_49699;
wire v_49700;
wire v_49701;
wire v_49702;
wire v_49703;
wire v_49704;
wire v_49705;
wire v_49706;
wire v_49707;
wire v_49708;
wire v_49709;
wire v_49710;
wire v_49711;
wire v_49712;
wire v_49713;
wire v_49714;
wire v_49715;
wire v_49716;
wire v_49717;
wire v_49718;
wire v_49719;
wire v_49720;
wire v_49721;
wire v_49722;
wire v_49723;
wire v_49724;
wire v_49725;
wire v_49726;
wire v_49727;
wire v_49728;
wire v_49729;
wire v_49730;
wire v_49731;
wire v_49732;
wire v_49733;
wire v_49734;
wire v_49735;
wire v_49736;
wire v_49737;
wire v_49738;
wire v_49739;
wire v_49740;
wire v_49741;
wire v_49742;
wire v_49743;
wire v_49744;
wire v_49745;
wire v_49746;
wire v_49747;
wire v_49748;
wire v_49749;
wire v_49750;
wire v_49751;
wire v_49752;
wire v_49753;
wire v_49754;
wire v_49755;
wire v_49756;
wire v_49757;
wire v_49758;
wire v_49759;
wire v_49760;
wire v_49761;
wire v_49762;
wire v_49763;
wire v_49764;
wire v_49765;
wire v_49766;
wire v_49767;
wire v_49768;
wire v_49769;
wire v_49770;
wire v_49771;
wire v_49772;
wire v_49773;
wire v_49774;
wire v_49775;
wire v_49776;
wire v_49777;
wire v_49778;
wire v_49779;
wire v_49780;
wire v_49781;
wire v_49782;
wire v_49783;
wire v_49784;
wire v_49785;
wire v_49786;
wire v_49787;
wire v_49788;
wire v_49789;
wire v_49790;
wire v_49791;
wire v_49792;
wire v_49793;
wire v_49794;
wire v_49795;
wire v_49796;
wire v_49797;
wire v_49798;
wire v_49799;
wire v_49800;
wire v_49801;
wire v_49802;
wire v_49803;
wire v_49804;
wire v_49805;
wire v_49806;
wire v_49807;
wire v_49808;
wire v_49809;
wire v_49810;
wire v_49811;
wire v_49812;
wire v_49813;
wire v_49814;
wire v_49815;
wire v_49816;
wire v_49817;
wire v_49818;
wire v_49819;
wire v_49820;
wire v_49821;
wire v_49822;
wire v_49823;
wire v_49824;
wire v_49825;
wire v_49826;
wire v_49827;
wire v_49828;
wire v_49829;
wire v_49830;
wire v_49831;
wire v_49832;
wire v_49833;
wire v_49834;
wire v_49835;
wire v_49836;
wire v_49837;
wire v_49838;
wire v_49839;
wire v_49840;
wire v_49841;
wire v_49842;
wire v_49843;
wire v_49844;
wire v_49845;
wire v_49846;
wire v_49847;
wire v_49848;
wire v_49849;
wire v_49850;
wire v_49851;
wire v_49852;
wire v_49853;
wire v_49854;
wire v_49855;
wire v_49856;
wire v_49857;
wire v_49858;
wire v_49859;
wire v_49860;
wire v_49861;
wire v_49862;
wire v_49863;
wire v_49864;
wire v_49865;
wire v_49866;
wire v_49867;
wire v_49868;
wire v_49869;
wire v_49870;
wire v_49871;
wire v_49872;
wire v_49873;
wire v_49874;
wire v_49875;
wire v_49876;
wire v_49877;
wire v_49878;
wire v_49879;
wire v_49880;
wire v_49881;
wire v_49882;
wire v_49883;
wire v_49884;
wire v_49885;
wire v_49886;
wire v_49887;
wire v_49888;
wire v_49889;
wire v_49890;
wire v_49891;
wire v_49892;
wire v_49893;
wire v_49894;
wire v_49895;
wire v_49896;
wire v_49897;
wire v_49898;
wire v_49899;
wire v_49900;
wire v_49901;
wire v_49902;
wire v_49903;
wire v_49904;
wire v_49905;
wire v_49906;
wire v_49907;
wire v_49908;
wire v_49909;
wire v_49910;
wire v_49911;
wire v_49912;
wire v_49913;
wire v_49914;
wire v_49915;
wire v_49916;
wire v_49917;
wire v_49918;
wire v_49919;
wire v_49920;
wire v_49921;
wire v_49922;
wire v_49923;
wire v_49924;
wire v_49925;
wire v_49926;
wire v_49927;
wire v_49928;
wire v_49929;
wire v_49930;
wire v_49931;
wire v_49932;
wire v_49933;
wire v_49934;
wire v_49935;
wire v_49936;
wire v_49937;
wire v_49938;
wire v_49939;
wire v_49940;
wire v_49941;
wire v_49942;
wire v_49943;
wire v_49944;
wire v_49945;
wire v_49946;
wire v_49947;
wire v_49948;
wire v_49949;
wire v_49950;
wire v_49951;
wire v_49952;
wire v_49953;
wire v_49954;
wire v_49955;
wire v_49956;
wire v_49957;
wire v_49958;
wire v_49959;
wire v_49960;
wire v_49961;
wire v_49962;
wire v_49963;
wire v_49964;
wire v_49965;
wire v_49966;
wire v_49967;
wire v_49968;
wire v_49969;
wire v_49970;
wire v_49971;
wire v_49972;
wire v_49973;
wire v_49974;
wire v_49975;
wire v_49977;
wire v_49978;
wire v_49979;
wire v_49980;
wire v_49981;
wire v_49982;
wire v_49983;
wire v_49984;
wire v_49985;
wire v_49986;
wire v_49987;
wire v_49988;
wire v_49989;
wire v_49990;
wire v_49991;
wire v_49992;
wire v_49993;
wire v_49994;
wire v_49995;
wire v_49996;
wire v_49997;
wire v_49998;
wire v_49999;
wire v_50000;
wire v_50001;
wire v_50002;
wire v_50003;
wire v_50004;
wire v_50005;
wire v_50006;
wire v_50007;
wire v_50008;
wire v_50009;
wire v_50010;
wire v_50011;
wire v_50012;
wire v_50013;
wire v_50014;
wire v_50015;
wire v_50016;
wire v_50017;
wire v_50018;
wire v_50019;
wire v_50020;
wire v_50021;
wire v_50022;
wire v_50023;
wire v_50024;
wire v_50025;
wire v_50026;
wire v_50027;
wire v_50028;
wire v_50029;
wire v_50030;
wire v_50031;
wire v_50032;
wire v_50033;
wire v_50034;
wire v_50035;
wire v_50036;
wire v_50037;
wire v_50038;
wire v_50039;
wire v_50040;
wire v_50041;
wire v_50042;
wire v_50043;
wire v_50044;
wire v_50045;
wire v_50046;
wire v_50047;
wire v_50048;
wire v_50049;
wire v_50050;
wire v_50051;
wire v_50052;
wire v_50053;
wire v_50054;
wire v_50055;
wire v_50056;
wire v_50057;
wire v_50058;
wire v_50059;
wire v_50060;
wire v_50061;
wire v_50062;
wire v_50063;
wire v_50064;
wire v_50065;
wire v_50066;
wire v_50067;
wire v_50068;
wire v_50069;
wire v_50071;
wire v_50073;
wire v_50074;
wire v_50075;
wire v_50077;
wire v_50078;
wire v_50079;
wire v_50081;
wire v_50082;
wire v_50083;
wire v_50085;
wire v_50086;
wire v_50088;
wire v_50089;
wire v_50090;
wire v_50092;
wire v_50093;
wire v_50094;
wire v_50096;
wire v_50097;
wire v_50098;
wire v_50100;
wire v_50101;
wire v_50102;
wire v_50104;
wire v_50105;
wire v_50106;
wire v_50108;
wire v_50109;
wire v_50110;
wire v_50112;
wire v_50113;
wire v_50114;
wire v_50116;
wire v_50117;
wire v_50118;
wire v_50120;
wire v_50121;
wire v_50122;
wire v_50124;
wire v_50125;
wire v_50126;
wire v_50128;
wire v_50129;
wire v_50130;
wire v_50132;
wire v_50133;
wire v_50134;
wire v_50136;
wire v_50137;
wire v_50138;
wire v_50139;
wire v_50140;
wire v_50141;
wire v_50142;
wire v_50143;
wire v_50144;
wire v_50145;
wire v_50146;
wire v_50147;
wire v_50148;
wire v_50149;
wire v_50150;
wire v_50151;
wire v_50152;
wire v_50153;
wire v_50154;
wire v_50155;
wire v_50156;
wire v_50157;
wire v_50158;
wire v_50159;
wire v_50160;
wire v_50161;
wire v_50162;
wire v_50163;
wire v_50164;
wire v_50165;
wire v_50166;
wire v_50167;
wire v_50168;
wire v_50169;
wire v_50170;
wire v_50171;
wire v_50172;
wire v_50173;
wire v_50174;
wire v_50175;
wire v_50176;
wire v_50177;
wire v_50178;
wire v_50179;
wire v_50180;
wire v_50181;
wire v_50182;
wire v_50183;
wire v_50184;
wire v_50185;
wire v_50186;
wire v_50187;
wire v_50188;
wire v_50189;
wire v_50190;
wire v_50191;
wire v_50192;
wire v_50193;
wire v_50194;
wire v_50195;
wire v_50196;
wire v_50197;
wire v_50198;
wire v_50199;
wire v_50200;
wire v_50201;
wire v_50202;
wire v_50203;
wire v_50204;
wire v_50205;
wire v_50206;
wire v_50207;
wire v_50208;
wire v_50209;
wire v_50210;
wire v_50211;
wire v_50212;
wire v_50213;
wire v_50214;
wire v_50215;
wire v_50216;
wire v_50217;
wire v_50218;
wire v_50219;
wire v_50220;
wire v_50221;
wire v_50222;
wire v_50223;
wire v_50224;
wire v_50225;
wire v_50226;
wire v_50227;
wire v_50228;
wire v_50229;
wire v_50230;
wire v_50231;
wire v_50232;
wire v_50233;
wire v_50234;
wire v_50235;
wire v_50236;
wire v_50237;
wire v_50238;
wire v_50239;
wire v_50240;
wire v_50241;
wire v_50242;
wire v_50243;
wire v_50244;
wire v_50245;
wire v_50246;
wire v_50247;
wire v_50248;
wire v_50249;
wire v_50250;
wire v_50251;
wire v_50252;
wire v_50253;
wire v_50254;
wire v_50255;
wire v_50256;
wire v_50257;
wire v_50258;
wire v_50259;
wire v_50260;
wire v_50261;
wire v_50262;
wire v_50263;
wire v_50264;
wire v_50265;
wire v_50266;
wire v_50267;
wire v_50268;
wire v_50269;
wire v_50270;
wire v_50271;
wire v_50272;
wire v_50273;
wire v_50274;
wire v_50275;
wire v_50276;
wire v_50277;
wire v_50278;
wire v_50279;
wire v_50280;
wire v_50281;
wire v_50282;
wire v_50283;
wire v_50284;
wire v_50285;
wire v_50286;
wire v_50287;
wire v_50288;
wire v_50289;
wire v_50290;
wire v_50291;
wire v_50292;
wire v_50293;
wire v_50294;
wire v_50295;
wire v_50296;
wire v_50297;
wire v_50298;
wire v_50299;
wire v_50300;
wire v_50301;
wire v_50302;
wire v_50303;
wire v_50304;
wire v_50305;
wire v_50306;
wire v_50307;
wire v_50308;
wire v_50309;
wire v_50310;
wire v_50311;
wire v_50312;
wire v_50313;
wire v_50314;
wire v_50315;
wire v_50316;
wire v_50317;
wire v_50318;
wire v_50319;
wire v_50320;
wire v_50321;
wire v_50322;
wire v_50323;
wire v_50324;
wire v_50325;
wire v_50326;
wire v_50327;
wire v_50328;
wire v_50329;
wire v_50331;
wire v_50332;
wire v_50333;
wire v_50334;
wire v_50335;
wire v_50336;
wire v_50337;
wire v_50338;
wire v_50339;
wire v_50340;
wire v_50341;
wire v_50342;
wire v_50343;
wire v_50344;
wire v_50345;
wire v_50346;
wire v_50347;
wire v_50348;
wire v_50349;
wire v_50350;
wire v_50351;
wire v_50352;
wire v_50353;
wire v_50354;
wire v_50355;
wire v_50356;
wire v_50357;
wire v_50358;
wire v_50359;
wire v_50360;
wire v_50361;
wire v_50362;
wire v_50363;
wire v_50364;
wire v_50365;
wire v_50366;
wire v_50367;
wire v_50368;
wire v_50369;
wire v_50370;
wire v_50371;
wire v_50372;
wire v_50373;
wire v_50374;
wire v_50375;
wire v_50376;
wire v_50377;
wire v_50378;
wire v_50379;
wire v_50380;
wire v_50381;
wire v_50382;
wire v_50383;
wire v_50384;
wire v_50385;
wire v_50386;
wire v_50387;
wire v_50388;
wire v_50389;
wire v_50390;
wire v_50391;
wire v_50392;
wire v_50393;
wire v_50394;
wire v_50395;
wire v_50396;
wire v_50397;
wire v_50398;
wire v_50399;
wire v_50400;
wire v_50401;
wire v_50402;
wire v_50403;
wire v_50404;
wire v_50405;
wire v_50406;
wire v_50407;
wire v_50408;
wire v_50409;
wire v_50410;
wire v_50411;
wire v_50412;
wire v_50413;
wire v_50414;
wire v_50415;
wire v_50416;
wire v_50417;
wire v_50418;
wire v_50419;
wire v_50420;
wire v_50421;
wire v_50422;
wire v_50423;
wire v_50424;
wire v_50425;
wire v_50426;
wire v_50427;
wire v_50428;
wire v_50429;
wire v_50430;
wire v_50431;
wire v_50432;
wire v_50433;
wire v_50434;
wire v_50435;
wire v_50436;
wire v_50437;
wire v_50438;
wire v_50439;
wire v_50440;
wire v_50441;
wire v_50442;
wire v_50443;
wire v_50444;
wire v_50445;
wire v_50446;
wire v_50447;
wire v_50448;
wire v_50449;
wire v_50450;
wire v_50451;
wire v_50452;
wire v_50453;
wire v_50454;
wire v_50455;
wire v_50456;
wire v_50457;
wire v_50458;
wire v_50459;
wire v_50460;
wire v_50461;
wire v_50462;
wire v_50463;
wire v_50464;
wire v_50465;
wire v_50466;
wire v_50467;
wire v_50468;
wire v_50469;
wire v_50470;
wire v_50471;
wire v_50472;
wire v_50473;
wire v_50474;
wire v_50475;
wire v_50476;
wire v_50477;
wire v_50478;
wire v_50479;
wire v_50480;
wire v_50481;
wire v_50482;
wire v_50483;
wire v_50484;
wire v_50485;
wire v_50486;
wire v_50487;
wire v_50488;
wire v_50489;
wire v_50490;
wire v_50491;
wire v_50492;
wire v_50493;
wire v_50494;
wire v_50495;
wire v_50496;
wire v_50497;
wire v_50498;
wire v_50499;
wire v_50500;
wire v_50501;
wire v_50502;
wire v_50503;
wire v_50504;
wire v_50505;
wire v_50506;
wire v_50507;
wire v_50508;
wire v_50509;
wire v_50510;
wire v_50511;
wire v_50512;
wire v_50513;
wire v_50514;
wire v_50515;
wire v_50516;
wire v_50517;
wire v_50518;
wire v_50519;
wire v_50520;
wire v_50521;
wire v_50522;
wire v_50523;
wire v_50524;
wire v_50525;
wire v_50526;
wire v_50527;
wire v_50528;
wire v_50529;
wire v_50530;
wire v_50531;
wire v_50532;
wire v_50533;
wire v_50534;
wire v_50535;
wire v_50536;
wire v_50537;
wire v_50538;
wire v_50539;
wire v_50540;
wire v_50541;
wire v_50542;
wire v_50543;
wire v_50544;
wire v_50545;
wire v_50546;
wire v_50547;
wire v_50548;
wire v_50549;
wire v_50550;
wire v_50551;
wire v_50552;
wire v_50553;
wire v_50554;
wire v_50555;
wire v_50556;
wire v_50557;
wire v_50558;
wire v_50559;
wire v_50560;
wire v_50561;
wire v_50562;
wire v_50563;
wire v_50564;
wire v_50565;
wire v_50566;
wire v_50567;
wire v_50568;
wire v_50569;
wire v_50570;
wire v_50571;
wire v_50572;
wire v_50574;
wire v_50575;
wire v_50576;
wire v_50577;
wire v_50578;
wire v_50579;
wire v_50580;
wire v_50581;
wire v_50582;
wire v_50583;
wire v_50584;
wire v_50585;
wire v_50586;
wire v_50587;
wire v_50588;
wire v_50589;
wire v_50590;
wire v_50591;
wire v_50592;
wire v_50593;
wire v_50594;
wire v_50595;
wire v_50596;
wire v_50597;
wire v_50598;
wire v_50599;
wire v_50600;
wire v_50601;
wire v_50602;
wire v_50603;
wire v_50604;
wire v_50605;
wire v_50606;
wire v_50607;
wire v_50608;
wire v_50609;
wire v_50610;
wire v_50611;
wire v_50612;
wire v_50613;
wire v_50614;
wire v_50615;
wire v_50616;
wire v_50617;
wire v_50618;
wire v_50619;
wire v_50620;
wire v_50621;
wire v_50622;
wire v_50623;
wire v_50624;
wire v_50625;
wire v_50626;
wire v_50627;
wire v_50628;
wire v_50629;
wire v_50630;
wire v_50631;
wire v_50632;
wire v_50633;
wire v_50634;
wire v_50635;
wire v_50636;
wire v_50637;
wire v_50638;
wire v_50639;
wire v_50640;
wire v_50641;
wire v_50642;
wire v_50643;
wire v_50644;
wire v_50645;
wire v_50646;
wire v_50647;
wire v_50648;
wire v_50649;
wire v_50650;
wire v_50651;
wire v_50652;
wire v_50653;
wire v_50654;
wire v_50655;
wire v_50656;
wire v_50657;
wire v_50658;
wire v_50659;
wire v_50660;
wire v_50661;
wire v_50662;
wire v_50663;
wire v_50664;
wire v_50665;
wire v_50666;
wire v_50667;
wire v_50668;
wire v_50669;
wire v_50670;
wire v_50671;
wire v_50672;
wire v_50673;
wire v_50674;
wire v_50675;
wire v_50676;
wire v_50677;
wire v_50678;
wire v_50679;
wire v_50680;
wire v_50681;
wire v_50682;
wire v_50683;
wire v_50684;
wire v_50685;
wire v_50686;
wire v_50687;
wire v_50688;
wire v_50689;
wire v_50690;
wire v_50691;
wire v_50692;
wire v_50693;
wire v_50694;
wire v_50695;
wire v_50696;
wire v_50697;
wire v_50698;
wire v_50699;
wire v_50700;
wire v_50701;
wire v_50702;
wire v_50703;
wire v_50704;
wire v_50705;
wire v_50706;
wire v_50707;
wire v_50708;
wire v_50709;
wire v_50710;
wire v_50711;
wire v_50712;
wire v_50713;
wire v_50714;
wire v_50715;
wire v_50716;
wire v_50717;
wire v_50718;
wire v_50719;
wire v_50720;
wire v_50721;
wire v_50722;
wire v_50723;
wire v_50724;
wire v_50725;
wire v_50726;
wire v_50727;
wire v_50728;
wire v_50729;
wire v_50730;
wire v_50731;
wire v_50732;
wire v_50733;
wire v_50734;
wire v_50735;
wire v_50736;
wire v_50737;
wire v_50738;
wire v_50739;
wire v_50740;
wire v_50741;
wire v_50742;
wire v_50743;
wire v_50744;
wire v_50745;
wire v_50746;
wire v_50747;
wire v_50748;
wire v_50749;
wire v_50750;
wire v_50751;
wire v_50752;
wire v_50753;
wire v_50754;
wire v_50755;
wire v_50756;
wire v_50757;
wire v_50758;
wire v_50759;
wire v_50760;
wire v_50761;
wire v_50762;
wire v_50763;
wire v_50764;
wire v_50765;
wire v_50766;
wire v_50767;
wire v_50768;
wire v_50769;
wire v_50770;
wire v_50771;
wire v_50772;
wire v_50773;
wire v_50774;
wire v_50775;
wire v_50776;
wire v_50777;
wire v_50778;
wire v_50779;
wire v_50780;
wire v_50781;
wire v_50782;
wire v_50783;
wire v_50784;
wire v_50785;
wire v_50786;
wire v_50787;
wire v_50788;
wire v_50789;
wire v_50790;
wire v_50791;
wire v_50792;
wire v_50793;
wire v_50794;
wire v_50795;
wire v_50796;
wire v_50797;
wire v_50798;
wire v_50799;
wire v_50800;
wire v_50801;
wire v_50802;
wire v_50803;
wire v_50804;
wire v_50805;
wire v_50806;
wire v_50807;
wire v_50808;
wire v_50809;
wire v_50810;
wire v_50811;
wire v_50812;
wire v_50813;
wire v_50814;
wire v_50815;
wire v_50817;
wire v_50818;
wire v_50819;
wire v_50820;
wire v_50821;
wire v_50822;
wire v_50823;
wire v_50824;
wire v_50825;
wire v_50826;
wire v_50827;
wire v_50828;
wire v_50829;
wire v_50830;
wire v_50831;
wire v_50832;
wire v_50833;
wire v_50834;
wire v_50835;
wire v_50836;
wire v_50837;
wire v_50838;
wire v_50839;
wire v_50840;
wire v_50841;
wire v_50842;
wire v_50843;
wire v_50844;
wire v_50845;
wire v_50846;
wire v_50847;
wire v_50848;
wire v_50849;
wire v_50850;
wire v_50851;
wire v_50852;
wire v_50853;
wire v_50854;
wire v_50855;
wire v_50856;
wire v_50857;
wire v_50858;
wire v_50859;
wire v_50860;
wire v_50861;
wire v_50862;
wire v_50863;
wire v_50864;
wire v_50865;
wire v_50866;
wire v_50867;
wire v_50868;
wire v_50869;
wire v_50870;
wire v_50871;
wire v_50872;
wire v_50873;
wire v_50874;
wire v_50875;
wire v_50876;
wire v_50877;
wire v_50878;
wire v_50879;
wire v_50880;
wire v_50881;
wire v_50882;
wire v_50883;
wire v_50884;
wire v_50885;
wire v_50886;
wire v_50887;
wire v_50888;
wire v_50889;
wire v_50890;
wire v_50891;
wire v_50892;
wire v_50893;
wire v_50894;
wire v_50895;
wire v_50896;
wire v_50897;
wire v_50898;
wire v_50899;
wire v_50900;
wire v_50901;
wire v_50902;
wire v_50903;
wire v_50904;
wire v_50905;
wire v_50906;
wire v_50907;
wire v_50908;
wire v_50909;
wire v_50910;
wire v_50911;
wire v_50912;
wire v_50913;
wire v_50914;
wire v_50915;
wire v_50916;
wire v_50917;
wire v_50918;
wire v_50919;
wire v_50920;
wire v_50921;
wire v_50922;
wire v_50923;
wire v_50924;
wire v_50925;
wire v_50926;
wire v_50927;
wire v_50928;
wire v_50929;
wire v_50930;
wire v_50931;
wire v_50932;
wire v_50933;
wire v_50934;
wire v_50935;
wire v_50936;
wire v_50937;
wire v_50938;
wire v_50939;
wire v_50940;
wire v_50941;
wire v_50942;
wire v_50943;
wire v_50944;
wire v_50945;
wire v_50946;
wire v_50947;
wire v_50948;
wire v_50949;
wire v_50950;
wire v_50951;
wire v_50952;
wire v_50953;
wire v_50954;
wire v_50955;
wire v_50956;
wire v_50957;
wire v_50958;
wire v_50959;
wire v_50960;
wire v_50961;
wire v_50962;
wire v_50963;
wire v_50964;
wire v_50965;
wire v_50966;
wire v_50967;
wire v_50968;
wire v_50969;
wire v_50970;
wire v_50971;
wire v_50972;
wire v_50973;
wire v_50974;
wire v_50975;
wire v_50976;
wire v_50977;
wire v_50978;
wire v_50979;
wire v_50980;
wire v_50981;
wire v_50982;
wire v_50983;
wire v_50984;
wire v_50985;
wire v_50986;
wire v_50987;
wire v_50988;
wire v_50989;
wire v_50990;
wire v_50991;
wire v_50992;
wire v_50993;
wire v_50994;
wire v_50995;
wire v_50996;
wire v_50997;
wire v_50998;
wire v_50999;
wire v_51000;
wire v_51001;
wire v_51002;
wire v_51003;
wire v_51004;
wire v_51005;
wire v_51006;
wire v_51007;
wire v_51008;
wire v_51009;
wire v_51010;
wire v_51011;
wire v_51012;
wire v_51013;
wire v_51014;
wire v_51015;
wire v_51016;
wire v_51017;
wire v_51018;
wire v_51019;
wire v_51020;
wire v_51021;
wire v_51022;
wire v_51023;
wire v_51024;
wire v_51025;
wire v_51026;
wire v_51027;
wire v_51028;
wire v_51029;
wire v_51030;
wire v_51031;
wire v_51032;
wire v_51033;
wire v_51034;
wire v_51035;
wire v_51036;
wire v_51037;
wire v_51038;
wire v_51039;
wire v_51040;
wire v_51041;
wire v_51042;
wire v_51043;
wire v_51044;
wire v_51045;
wire v_51046;
wire v_51047;
wire v_51048;
wire v_51049;
wire v_51050;
wire v_51051;
wire v_51052;
wire v_51053;
wire v_51054;
wire v_51055;
wire v_51056;
wire v_51057;
wire v_51058;
wire v_51060;
wire v_51061;
wire v_51062;
wire v_51063;
wire v_51064;
wire v_51065;
wire v_51066;
wire v_51067;
wire v_51068;
wire v_51069;
wire v_51070;
wire v_51071;
wire v_51072;
wire v_51073;
wire v_51074;
wire v_51075;
wire v_51076;
wire v_51077;
wire v_51078;
wire v_51079;
wire v_51080;
wire v_51081;
wire v_51082;
wire v_51083;
wire v_51084;
wire v_51085;
wire v_51086;
wire v_51087;
wire v_51088;
wire v_51089;
wire v_51090;
wire v_51091;
wire v_51092;
wire v_51093;
wire v_51094;
wire v_51095;
wire v_51096;
wire v_51097;
wire v_51098;
wire v_51099;
wire v_51100;
wire v_51101;
wire v_51102;
wire v_51103;
wire v_51104;
wire v_51105;
wire v_51106;
wire v_51107;
wire v_51108;
wire v_51109;
wire v_51110;
wire v_51111;
wire v_51112;
wire v_51113;
wire v_51114;
wire v_51115;
wire v_51116;
wire v_51117;
wire v_51118;
wire v_51119;
wire v_51120;
wire v_51121;
wire v_51122;
wire v_51123;
wire v_51124;
wire v_51125;
wire v_51126;
wire v_51127;
wire v_51128;
wire v_51129;
wire v_51130;
wire v_51131;
wire v_51132;
wire v_51133;
wire v_51134;
wire v_51135;
wire v_51136;
wire v_51137;
wire v_51138;
wire v_51139;
wire v_51140;
wire v_51141;
wire v_51142;
wire v_51143;
wire v_51144;
wire v_51145;
wire v_51146;
wire v_51147;
wire v_51148;
wire v_51149;
wire v_51150;
wire v_51151;
wire v_51152;
wire v_51153;
wire v_51154;
wire v_51155;
wire v_51156;
wire v_51157;
wire v_51158;
wire v_51159;
wire v_51160;
wire v_51161;
wire v_51162;
wire v_51163;
wire v_51164;
wire v_51165;
wire v_51166;
wire v_51167;
wire v_51168;
wire v_51169;
wire v_51170;
wire v_51171;
wire v_51172;
wire v_51173;
wire v_51174;
wire v_51175;
wire v_51176;
wire v_51177;
wire v_51178;
wire v_51179;
wire v_51180;
wire v_51181;
wire v_51182;
wire v_51183;
wire v_51184;
wire v_51185;
wire v_51186;
wire v_51187;
wire v_51188;
wire v_51189;
wire v_51190;
wire v_51191;
wire v_51192;
wire v_51193;
wire v_51194;
wire v_51195;
wire v_51196;
wire v_51197;
wire v_51198;
wire v_51199;
wire v_51200;
wire v_51201;
wire v_51202;
wire v_51203;
wire v_51204;
wire v_51205;
wire v_51206;
wire v_51207;
wire v_51208;
wire v_51209;
wire v_51210;
wire v_51211;
wire v_51212;
wire v_51213;
wire v_51214;
wire v_51215;
wire v_51216;
wire v_51217;
wire v_51218;
wire v_51219;
wire v_51220;
wire v_51221;
wire v_51222;
wire v_51223;
wire v_51224;
wire v_51225;
wire v_51226;
wire v_51227;
wire v_51228;
wire v_51229;
wire v_51230;
wire v_51231;
wire v_51232;
wire v_51233;
wire v_51234;
wire v_51235;
wire v_51236;
wire v_51237;
wire v_51238;
wire v_51239;
wire v_51240;
wire v_51241;
wire v_51242;
wire v_51243;
wire v_51244;
wire v_51245;
wire v_51246;
wire v_51247;
wire v_51248;
wire v_51249;
wire v_51250;
wire v_51251;
wire v_51252;
wire v_51253;
wire v_51254;
wire v_51255;
wire v_51256;
wire v_51257;
wire v_51258;
wire v_51259;
wire v_51260;
wire v_51261;
wire v_51262;
wire v_51263;
wire v_51264;
wire v_51265;
wire v_51266;
wire v_51267;
wire v_51268;
wire v_51269;
wire v_51270;
wire v_51271;
wire v_51272;
wire v_51273;
wire v_51274;
wire v_51275;
wire v_51276;
wire v_51277;
wire v_51278;
wire v_51279;
wire v_51280;
wire v_51281;
wire v_51282;
wire v_51283;
wire v_51284;
wire v_51285;
wire v_51286;
wire v_51287;
wire v_51288;
wire v_51289;
wire v_51290;
wire v_51291;
wire v_51292;
wire v_51293;
wire v_51294;
wire v_51295;
wire v_51296;
wire v_51297;
wire v_51298;
wire v_51299;
wire v_51300;
wire v_51301;
wire v_51303;
wire v_51304;
wire v_51305;
wire v_51306;
wire v_51307;
wire v_51308;
wire v_51309;
wire v_51310;
wire v_51311;
wire v_51312;
wire v_51313;
wire v_51314;
wire v_51315;
wire v_51316;
wire v_51317;
wire v_51318;
wire v_51319;
wire v_51320;
wire v_51321;
wire v_51322;
wire v_51323;
wire v_51324;
wire v_51325;
wire v_51326;
wire v_51327;
wire v_51328;
wire v_51329;
wire v_51330;
wire v_51331;
wire v_51332;
wire v_51333;
wire v_51334;
wire v_51335;
wire v_51336;
wire v_51337;
wire v_51338;
wire v_51339;
wire v_51340;
wire v_51341;
wire v_51342;
wire v_51343;
wire v_51344;
wire v_51345;
wire v_51346;
wire v_51347;
wire v_51348;
wire v_51349;
wire v_51350;
wire v_51351;
wire v_51352;
wire v_51353;
wire v_51354;
wire v_51355;
wire v_51356;
wire v_51357;
wire v_51358;
wire v_51359;
wire v_51360;
wire v_51361;
wire v_51362;
wire v_51363;
wire v_51364;
wire v_51365;
wire v_51366;
wire v_51367;
wire v_51368;
wire v_51369;
wire v_51370;
wire v_51371;
wire v_51372;
wire v_51373;
wire v_51374;
wire v_51375;
wire v_51376;
wire v_51377;
wire v_51378;
wire v_51379;
wire v_51380;
wire v_51381;
wire v_51382;
wire v_51383;
wire v_51384;
wire v_51385;
wire v_51386;
wire v_51387;
wire v_51388;
wire v_51389;
wire v_51390;
wire v_51391;
wire v_51392;
wire v_51393;
wire v_51394;
wire v_51395;
wire v_51396;
wire v_51397;
wire v_51398;
wire v_51399;
wire v_51400;
wire v_51401;
wire v_51402;
wire v_51403;
wire v_51404;
wire v_51405;
wire v_51406;
wire v_51407;
wire v_51408;
wire v_51409;
wire v_51410;
wire v_51411;
wire v_51412;
wire v_51413;
wire v_51414;
wire v_51415;
wire v_51416;
wire v_51417;
wire v_51418;
wire v_51419;
wire v_51420;
wire v_51421;
wire v_51422;
wire v_51423;
wire v_51424;
wire v_51425;
wire v_51426;
wire v_51427;
wire v_51428;
wire v_51429;
wire v_51430;
wire v_51431;
wire v_51432;
wire v_51433;
wire v_51434;
wire v_51435;
wire v_51436;
wire v_51437;
wire v_51438;
wire v_51439;
wire v_51440;
wire v_51441;
wire v_51442;
wire v_51443;
wire v_51444;
wire v_51445;
wire v_51446;
wire v_51447;
wire v_51448;
wire v_51449;
wire v_51450;
wire v_51451;
wire v_51452;
wire v_51453;
wire v_51454;
wire v_51455;
wire v_51456;
wire v_51457;
wire v_51458;
wire v_51459;
wire v_51460;
wire v_51461;
wire v_51462;
wire v_51463;
wire v_51464;
wire v_51465;
wire v_51466;
wire v_51467;
wire v_51468;
wire v_51469;
wire v_51470;
wire v_51471;
wire v_51472;
wire v_51473;
wire v_51474;
wire v_51475;
wire v_51476;
wire v_51477;
wire v_51478;
wire v_51479;
wire v_51480;
wire v_51481;
wire v_51482;
wire v_51483;
wire v_51484;
wire v_51485;
wire v_51486;
wire v_51487;
wire v_51488;
wire v_51489;
wire v_51490;
wire v_51491;
wire v_51492;
wire v_51493;
wire v_51494;
wire v_51495;
wire v_51496;
wire v_51497;
wire v_51498;
wire v_51499;
wire v_51500;
wire v_51501;
wire v_51502;
wire v_51503;
wire v_51504;
wire v_51505;
wire v_51506;
wire v_51507;
wire v_51508;
wire v_51509;
wire v_51510;
wire v_51511;
wire v_51512;
wire v_51513;
wire v_51514;
wire v_51515;
wire v_51516;
wire v_51517;
wire v_51518;
wire v_51519;
wire v_51520;
wire v_51521;
wire v_51522;
wire v_51523;
wire v_51524;
wire v_51525;
wire v_51526;
wire v_51527;
wire v_51528;
wire v_51529;
wire v_51530;
wire v_51531;
wire v_51532;
wire v_51533;
wire v_51534;
wire v_51535;
wire v_51536;
wire v_51537;
wire v_51538;
wire v_51539;
wire v_51540;
wire v_51541;
wire v_51542;
wire v_51543;
wire v_51544;
wire v_51546;
wire v_51547;
wire v_51548;
wire v_51549;
wire v_51550;
wire v_51551;
wire v_51552;
wire v_51553;
wire v_51554;
wire v_51555;
wire v_51556;
wire v_51557;
wire v_51558;
wire v_51559;
wire v_51560;
wire v_51561;
wire v_51562;
wire v_51563;
wire v_51564;
wire v_51565;
wire v_51566;
wire v_51567;
wire v_51568;
wire v_51569;
wire v_51570;
wire v_51571;
wire v_51572;
wire v_51573;
wire v_51574;
wire v_51575;
wire v_51576;
wire v_51577;
wire v_51578;
wire v_51579;
wire v_51580;
wire v_51581;
wire v_51582;
wire v_51583;
wire v_51584;
wire v_51585;
wire v_51586;
wire v_51587;
wire v_51588;
wire v_51589;
wire v_51590;
wire v_51591;
wire v_51592;
wire v_51593;
wire v_51594;
wire v_51595;
wire v_51596;
wire v_51597;
wire v_51598;
wire v_51599;
wire v_51600;
wire v_51601;
wire v_51602;
wire v_51603;
wire v_51604;
wire v_51605;
wire v_51606;
wire v_51607;
wire v_51608;
wire v_51609;
wire v_51610;
wire v_51611;
wire v_51612;
wire v_51613;
wire v_51614;
wire v_51615;
wire v_51616;
wire v_51617;
wire v_51618;
wire v_51619;
wire v_51620;
wire v_51621;
wire v_51622;
wire v_51623;
wire v_51624;
wire v_51625;
wire v_51626;
wire v_51627;
wire v_51628;
wire v_51629;
wire v_51630;
wire v_51631;
wire v_51632;
wire v_51633;
wire v_51634;
wire v_51635;
wire v_51636;
wire v_51637;
wire v_51638;
wire v_51639;
wire v_51640;
wire v_51641;
wire v_51642;
wire v_51643;
wire v_51644;
wire v_51645;
wire v_51646;
wire v_51647;
wire v_51648;
wire v_51649;
wire v_51650;
wire v_51651;
wire v_51652;
wire v_51653;
wire v_51654;
wire v_51655;
wire v_51656;
wire v_51657;
wire v_51658;
wire v_51659;
wire v_51660;
wire v_51661;
wire v_51662;
wire v_51663;
wire v_51664;
wire v_51665;
wire v_51666;
wire v_51667;
wire v_51668;
wire v_51669;
wire v_51670;
wire v_51671;
wire v_51672;
wire v_51673;
wire v_51674;
wire v_51675;
wire v_51676;
wire v_51677;
wire v_51678;
wire v_51679;
wire v_51680;
wire v_51681;
wire v_51682;
wire v_51683;
wire v_51684;
wire v_51685;
wire v_51686;
wire v_51687;
wire v_51688;
wire v_51689;
wire v_51690;
wire v_51691;
wire v_51692;
wire v_51693;
wire v_51694;
wire v_51695;
wire v_51696;
wire v_51697;
wire v_51698;
wire v_51699;
wire v_51700;
wire v_51701;
wire v_51702;
wire v_51703;
wire v_51704;
wire v_51705;
wire v_51706;
wire v_51707;
wire v_51708;
wire v_51709;
wire v_51710;
wire v_51711;
wire v_51712;
wire v_51713;
wire v_51714;
wire v_51715;
wire v_51716;
wire v_51717;
wire v_51718;
wire v_51719;
wire v_51720;
wire v_51721;
wire v_51722;
wire v_51723;
wire v_51724;
wire v_51725;
wire v_51726;
wire v_51727;
wire v_51728;
wire v_51729;
wire v_51730;
wire v_51731;
wire v_51732;
wire v_51733;
wire v_51734;
wire v_51735;
wire v_51736;
wire v_51737;
wire v_51738;
wire v_51739;
wire v_51740;
wire v_51741;
wire v_51742;
wire v_51743;
wire v_51744;
wire v_51745;
wire v_51746;
wire v_51747;
wire v_51748;
wire v_51749;
wire v_51750;
wire v_51751;
wire v_51752;
wire v_51753;
wire v_51754;
wire v_51755;
wire v_51756;
wire v_51757;
wire v_51758;
wire v_51759;
wire v_51760;
wire v_51761;
wire v_51762;
wire v_51763;
wire v_51764;
wire v_51765;
wire v_51766;
wire v_51767;
wire v_51768;
wire v_51769;
wire v_51770;
wire v_51771;
wire v_51772;
wire v_51773;
wire v_51774;
wire v_51775;
wire v_51776;
wire v_51777;
wire v_51778;
wire v_51779;
wire v_51780;
wire v_51781;
wire v_51782;
wire v_51783;
wire v_51784;
wire v_51785;
wire v_51786;
wire v_51787;
wire v_51789;
wire v_51790;
wire v_51791;
wire v_51792;
wire v_51793;
wire v_51794;
wire v_51795;
wire v_51796;
wire v_51797;
wire v_51798;
wire v_51799;
wire v_51800;
wire v_51801;
wire v_51802;
wire v_51803;
wire v_51804;
wire v_51805;
wire v_51806;
wire v_51807;
wire v_51808;
wire v_51809;
wire v_51810;
wire v_51811;
wire v_51812;
wire v_51813;
wire v_51814;
wire v_51815;
wire v_51816;
wire v_51817;
wire v_51818;
wire v_51819;
wire v_51820;
wire v_51821;
wire v_51822;
wire v_51823;
wire v_51824;
wire v_51825;
wire v_51826;
wire v_51827;
wire v_51828;
wire v_51829;
wire v_51830;
wire v_51831;
wire v_51832;
wire v_51833;
wire v_51834;
wire v_51835;
wire v_51836;
wire v_51837;
wire v_51838;
wire v_51839;
wire v_51840;
wire v_51841;
wire v_51842;
wire v_51843;
wire v_51844;
wire v_51845;
wire v_51846;
wire v_51847;
wire v_51848;
wire v_51849;
wire v_51850;
wire v_51851;
wire v_51852;
wire v_51853;
wire v_51854;
wire v_51855;
wire v_51856;
wire v_51857;
wire v_51858;
wire v_51859;
wire v_51860;
wire v_51861;
wire v_51862;
wire v_51863;
wire v_51864;
wire v_51865;
wire v_51866;
wire v_51867;
wire v_51868;
wire v_51869;
wire v_51870;
wire v_51871;
wire v_51872;
wire v_51873;
wire v_51874;
wire v_51875;
wire v_51876;
wire v_51877;
wire v_51878;
wire v_51879;
wire v_51880;
wire v_51881;
wire v_51882;
wire v_51883;
wire v_51884;
wire v_51885;
wire v_51886;
wire v_51887;
wire v_51888;
wire v_51889;
wire v_51890;
wire v_51891;
wire v_51892;
wire v_51893;
wire v_51894;
wire v_51895;
wire v_51896;
wire v_51897;
wire v_51898;
wire v_51899;
wire v_51900;
wire v_51901;
wire v_51902;
wire v_51903;
wire v_51904;
wire v_51905;
wire v_51906;
wire v_51907;
wire v_51908;
wire v_51909;
wire v_51910;
wire v_51911;
wire v_51912;
wire v_51913;
wire v_51914;
wire v_51915;
wire v_51916;
wire v_51917;
wire v_51918;
wire v_51919;
wire v_51920;
wire v_51921;
wire v_51922;
wire v_51923;
wire v_51924;
wire v_51925;
wire v_51926;
wire v_51927;
wire v_51928;
wire v_51929;
wire v_51930;
wire v_51931;
wire v_51932;
wire v_51933;
wire v_51934;
wire v_51935;
wire v_51936;
wire v_51937;
wire v_51938;
wire v_51939;
wire v_51940;
wire v_51941;
wire v_51942;
wire v_51943;
wire v_51944;
wire v_51945;
wire v_51946;
wire v_51947;
wire v_51948;
wire v_51949;
wire v_51950;
wire v_51951;
wire v_51952;
wire v_51953;
wire v_51954;
wire v_51955;
wire v_51956;
wire v_51957;
wire v_51958;
wire v_51959;
wire v_51960;
wire v_51961;
wire v_51962;
wire v_51963;
wire v_51964;
wire v_51965;
wire v_51966;
wire v_51967;
wire v_51968;
wire v_51969;
wire v_51970;
wire v_51971;
wire v_51972;
wire v_51973;
wire v_51974;
wire v_51975;
wire v_51976;
wire v_51977;
wire v_51978;
wire v_51979;
wire v_51980;
wire v_51981;
wire v_51982;
wire v_51983;
wire v_51984;
wire v_51985;
wire v_51986;
wire v_51987;
wire v_51988;
wire v_51989;
wire v_51990;
wire v_51991;
wire v_51992;
wire v_51993;
wire v_51994;
wire v_51995;
wire v_51996;
wire v_51997;
wire v_51998;
wire v_51999;
wire v_52000;
wire v_52001;
wire v_52002;
wire v_52003;
wire v_52004;
wire v_52005;
wire v_52006;
wire v_52007;
wire v_52008;
wire v_52009;
wire v_52010;
wire v_52011;
wire v_52012;
wire v_52013;
wire v_52014;
wire v_52015;
wire v_52016;
wire v_52017;
wire v_52018;
wire v_52019;
wire v_52020;
wire v_52021;
wire v_52022;
wire v_52023;
wire v_52024;
wire v_52025;
wire v_52026;
wire v_52027;
wire v_52028;
wire v_52029;
wire v_52030;
wire v_52032;
wire v_52033;
wire v_52034;
wire v_52035;
wire v_52036;
wire v_52037;
wire v_52038;
wire v_52039;
wire v_52040;
wire v_52041;
wire v_52042;
wire v_52043;
wire v_52044;
wire v_52045;
wire v_52046;
wire v_52047;
wire v_52048;
wire v_52049;
wire v_52050;
wire v_52051;
wire v_52052;
wire v_52053;
wire v_52054;
wire v_52055;
wire v_52056;
wire v_52057;
wire v_52058;
wire v_52059;
wire v_52060;
wire v_52061;
wire v_52062;
wire v_52063;
wire v_52064;
wire v_52065;
wire v_52066;
wire v_52067;
wire v_52068;
wire v_52069;
wire v_52070;
wire v_52071;
wire v_52072;
wire v_52073;
wire v_52074;
wire v_52075;
wire v_52076;
wire v_52077;
wire v_52078;
wire v_52079;
wire v_52080;
wire v_52081;
wire v_52082;
wire v_52083;
wire v_52084;
wire v_52085;
wire v_52086;
wire v_52087;
wire v_52088;
wire v_52089;
wire v_52090;
wire v_52091;
wire v_52092;
wire v_52093;
wire v_52094;
wire v_52095;
wire v_52096;
wire v_52097;
wire v_52098;
wire v_52099;
wire v_52100;
wire v_52101;
wire v_52102;
wire v_52103;
wire v_52104;
wire v_52105;
wire v_52106;
wire v_52107;
wire v_52108;
wire v_52109;
wire v_52110;
wire v_52111;
wire v_52112;
wire v_52113;
wire v_52114;
wire v_52115;
wire v_52116;
wire v_52117;
wire v_52118;
wire v_52119;
wire v_52120;
wire v_52121;
wire v_52122;
wire v_52123;
wire v_52124;
wire v_52125;
wire v_52126;
wire v_52127;
wire v_52128;
wire v_52129;
wire v_52130;
wire v_52131;
wire v_52132;
wire v_52133;
wire v_52134;
wire v_52135;
wire v_52136;
wire v_52137;
wire v_52138;
wire v_52139;
wire v_52140;
wire v_52141;
wire v_52142;
wire v_52143;
wire v_52144;
wire v_52145;
wire v_52146;
wire v_52147;
wire v_52148;
wire v_52149;
wire v_52150;
wire v_52151;
wire v_52152;
wire v_52153;
wire v_52154;
wire v_52155;
wire v_52156;
wire v_52157;
wire v_52158;
wire v_52159;
wire v_52160;
wire v_52161;
wire v_52162;
wire v_52163;
wire v_52164;
wire v_52165;
wire v_52166;
wire v_52167;
wire v_52168;
wire v_52169;
wire v_52170;
wire v_52171;
wire v_52172;
wire v_52173;
wire v_52174;
wire v_52175;
wire v_52176;
wire v_52177;
wire v_52178;
wire v_52179;
wire v_52180;
wire v_52181;
wire v_52182;
wire v_52183;
wire v_52184;
wire v_52185;
wire v_52186;
wire v_52187;
wire v_52188;
wire v_52189;
wire v_52190;
wire v_52191;
wire v_52192;
wire v_52193;
wire v_52194;
wire v_52195;
wire v_52196;
wire v_52197;
wire v_52198;
wire v_52199;
wire v_52200;
wire v_52201;
wire v_52202;
wire v_52203;
wire v_52204;
wire v_52205;
wire v_52206;
wire v_52207;
wire v_52208;
wire v_52209;
wire v_52210;
wire v_52211;
wire v_52212;
wire v_52213;
wire v_52214;
wire v_52215;
wire v_52216;
wire v_52217;
wire v_52218;
wire v_52219;
wire v_52220;
wire v_52221;
wire v_52222;
wire v_52223;
wire v_52224;
wire v_52225;
wire v_52226;
wire v_52227;
wire v_52228;
wire v_52229;
wire v_52230;
wire v_52231;
wire v_52232;
wire v_52233;
wire v_52234;
wire v_52235;
wire v_52236;
wire v_52237;
wire v_52238;
wire v_52239;
wire v_52240;
wire v_52241;
wire v_52242;
wire v_52243;
wire v_52244;
wire v_52245;
wire v_52246;
wire v_52247;
wire v_52248;
wire v_52249;
wire v_52250;
wire v_52251;
wire v_52252;
wire v_52253;
wire v_52254;
wire v_52255;
wire v_52256;
wire v_52257;
wire v_52258;
wire v_52259;
wire v_52260;
wire v_52261;
wire v_52262;
wire v_52263;
wire v_52264;
wire v_52265;
wire v_52266;
wire v_52267;
wire v_52268;
wire v_52269;
wire v_52270;
wire v_52271;
wire v_52272;
wire v_52273;
wire v_52275;
wire v_52276;
wire v_52277;
wire v_52278;
wire v_52279;
wire v_52280;
wire v_52281;
wire v_52282;
wire v_52283;
wire v_52284;
wire v_52285;
wire v_52286;
wire v_52287;
wire v_52288;
wire v_52289;
wire v_52290;
wire v_52291;
wire v_52292;
wire v_52293;
wire v_52294;
wire v_52295;
wire v_52296;
wire v_52297;
wire v_52298;
wire v_52299;
wire v_52300;
wire v_52301;
wire v_52302;
wire v_52303;
wire v_52304;
wire v_52305;
wire v_52306;
wire v_52307;
wire v_52308;
wire v_52309;
wire v_52310;
wire v_52311;
wire v_52312;
wire v_52313;
wire v_52314;
wire v_52315;
wire v_52316;
wire v_52317;
wire v_52318;
wire v_52319;
wire v_52320;
wire v_52321;
wire v_52322;
wire v_52323;
wire v_52324;
wire v_52325;
wire v_52326;
wire v_52327;
wire v_52328;
wire v_52329;
wire v_52330;
wire v_52331;
wire v_52332;
wire v_52333;
wire v_52334;
wire v_52335;
wire v_52336;
wire v_52337;
wire v_52338;
wire v_52339;
wire v_52340;
wire v_52341;
wire v_52342;
wire v_52343;
wire v_52344;
wire v_52345;
wire v_52346;
wire v_52347;
wire v_52348;
wire v_52349;
wire v_52350;
wire v_52351;
wire v_52352;
wire v_52353;
wire v_52354;
wire v_52355;
wire v_52356;
wire v_52357;
wire v_52358;
wire v_52359;
wire v_52360;
wire v_52361;
wire v_52362;
wire v_52363;
wire v_52364;
wire v_52365;
wire v_52366;
wire v_52367;
wire v_52368;
wire v_52369;
wire v_52370;
wire v_52371;
wire v_52372;
wire v_52373;
wire v_52374;
wire v_52375;
wire v_52376;
wire v_52377;
wire v_52378;
wire v_52379;
wire v_52380;
wire v_52381;
wire v_52382;
wire v_52383;
wire v_52384;
wire v_52385;
wire v_52386;
wire v_52387;
wire v_52388;
wire v_52389;
wire v_52390;
wire v_52391;
wire v_52392;
wire v_52393;
wire v_52394;
wire v_52395;
wire v_52396;
wire v_52397;
wire v_52398;
wire v_52399;
wire v_52400;
wire v_52401;
wire v_52402;
wire v_52403;
wire v_52404;
wire v_52405;
wire v_52406;
wire v_52407;
wire v_52408;
wire v_52409;
wire v_52410;
wire v_52411;
wire v_52412;
wire v_52413;
wire v_52414;
wire v_52415;
wire v_52416;
wire v_52417;
wire v_52418;
wire v_52419;
wire v_52420;
wire v_52421;
wire v_52422;
wire v_52423;
wire v_52424;
wire v_52425;
wire v_52426;
wire v_52427;
wire v_52428;
wire v_52429;
wire v_52430;
wire v_52431;
wire v_52432;
wire v_52433;
wire v_52434;
wire v_52435;
wire v_52436;
wire v_52437;
wire v_52438;
wire v_52439;
wire v_52440;
wire v_52441;
wire v_52442;
wire v_52443;
wire v_52444;
wire v_52445;
wire v_52446;
wire v_52447;
wire v_52448;
wire v_52449;
wire v_52450;
wire v_52451;
wire v_52452;
wire v_52453;
wire v_52454;
wire v_52455;
wire v_52456;
wire v_52457;
wire v_52458;
wire v_52459;
wire v_52460;
wire v_52461;
wire v_52462;
wire v_52463;
wire v_52464;
wire v_52465;
wire v_52466;
wire v_52467;
wire v_52468;
wire v_52469;
wire v_52470;
wire v_52471;
wire v_52472;
wire v_52473;
wire v_52474;
wire v_52475;
wire v_52476;
wire v_52477;
wire v_52478;
wire v_52479;
wire v_52480;
wire v_52481;
wire v_52482;
wire v_52483;
wire v_52484;
wire v_52485;
wire v_52486;
wire v_52487;
wire v_52488;
wire v_52489;
wire v_52490;
wire v_52491;
wire v_52492;
wire v_52493;
wire v_52494;
wire v_52495;
wire v_52496;
wire v_52497;
wire v_52498;
wire v_52499;
wire v_52500;
wire v_52501;
wire v_52502;
wire v_52503;
wire v_52504;
wire v_52505;
wire v_52506;
wire v_52507;
wire v_52508;
wire v_52509;
wire v_52510;
wire v_52511;
wire v_52512;
wire v_52513;
wire v_52514;
wire v_52515;
wire v_52516;
wire v_52518;
wire v_52519;
wire v_52520;
wire v_52521;
wire v_52522;
wire v_52523;
wire v_52524;
wire v_52525;
wire v_52526;
wire v_52527;
wire v_52528;
wire v_52529;
wire v_52530;
wire v_52531;
wire v_52532;
wire v_52533;
wire v_52534;
wire v_52535;
wire v_52536;
wire v_52537;
wire v_52538;
wire v_52539;
wire v_52540;
wire v_52541;
wire v_52542;
wire v_52543;
wire v_52544;
wire v_52545;
wire v_52546;
wire v_52547;
wire v_52548;
wire v_52549;
wire v_52550;
wire v_52551;
wire v_52552;
wire v_52553;
wire v_52554;
wire v_52555;
wire v_52556;
wire v_52557;
wire v_52558;
wire v_52559;
wire v_52560;
wire v_52561;
wire v_52562;
wire v_52563;
wire v_52564;
wire v_52565;
wire v_52566;
wire v_52567;
wire v_52568;
wire v_52569;
wire v_52570;
wire v_52571;
wire v_52572;
wire v_52573;
wire v_52574;
wire v_52575;
wire v_52576;
wire v_52577;
wire v_52578;
wire v_52579;
wire v_52580;
wire v_52581;
wire v_52582;
wire v_52583;
wire v_52584;
wire v_52585;
wire v_52586;
wire v_52587;
wire v_52588;
wire v_52589;
wire v_52590;
wire v_52591;
wire v_52592;
wire v_52593;
wire v_52594;
wire v_52595;
wire v_52596;
wire v_52597;
wire v_52598;
wire v_52599;
wire v_52600;
wire v_52601;
wire v_52602;
wire v_52603;
wire v_52604;
wire v_52605;
wire v_52606;
wire v_52607;
wire v_52608;
wire v_52609;
wire v_52610;
wire v_52611;
wire v_52612;
wire v_52613;
wire v_52614;
wire v_52615;
wire v_52616;
wire v_52617;
wire v_52618;
wire v_52619;
wire v_52620;
wire v_52621;
wire v_52622;
wire v_52623;
wire v_52624;
wire v_52625;
wire v_52626;
wire v_52627;
wire v_52628;
wire v_52629;
wire v_52630;
wire v_52631;
wire v_52632;
wire v_52633;
wire v_52634;
wire v_52635;
wire v_52636;
wire v_52637;
wire v_52638;
wire v_52639;
wire v_52640;
wire v_52641;
wire v_52642;
wire v_52643;
wire v_52644;
wire v_52645;
wire v_52646;
wire v_52647;
wire v_52648;
wire v_52649;
wire v_52650;
wire v_52651;
wire v_52652;
wire v_52653;
wire v_52654;
wire v_52655;
wire v_52656;
wire v_52657;
wire v_52658;
wire v_52659;
wire v_52660;
wire v_52661;
wire v_52662;
wire v_52663;
wire v_52664;
wire v_52665;
wire v_52666;
wire v_52667;
wire v_52668;
wire v_52669;
wire v_52670;
wire v_52671;
wire v_52672;
wire v_52673;
wire v_52674;
wire v_52675;
wire v_52676;
wire v_52677;
wire v_52678;
wire v_52679;
wire v_52680;
wire v_52681;
wire v_52682;
wire v_52683;
wire v_52684;
wire v_52685;
wire v_52686;
wire v_52687;
wire v_52688;
wire v_52689;
wire v_52690;
wire v_52691;
wire v_52692;
wire v_52693;
wire v_52694;
wire v_52695;
wire v_52696;
wire v_52697;
wire v_52698;
wire v_52699;
wire v_52700;
wire v_52701;
wire v_52702;
wire v_52703;
wire v_52704;
wire v_52705;
wire v_52706;
wire v_52707;
wire v_52708;
wire v_52709;
wire v_52710;
wire v_52711;
wire v_52712;
wire v_52713;
wire v_52714;
wire v_52715;
wire v_52716;
wire v_52717;
wire v_52718;
wire v_52719;
wire v_52720;
wire v_52721;
wire v_52722;
wire v_52723;
wire v_52724;
wire v_52725;
wire v_52726;
wire v_52727;
wire v_52728;
wire v_52729;
wire v_52730;
wire v_52731;
wire v_52732;
wire v_52733;
wire v_52734;
wire v_52735;
wire v_52736;
wire v_52737;
wire v_52738;
wire v_52739;
wire v_52740;
wire v_52741;
wire v_52742;
wire v_52743;
wire v_52744;
wire v_52745;
wire v_52746;
wire v_52747;
wire v_52748;
wire v_52749;
wire v_52750;
wire v_52751;
wire v_52752;
wire v_52753;
wire v_52754;
wire v_52755;
wire v_52756;
wire v_52757;
wire v_52758;
wire v_52759;
wire v_52761;
wire v_52762;
wire v_52763;
wire v_52764;
wire v_52765;
wire v_52766;
wire v_52767;
wire v_52768;
wire v_52769;
wire v_52770;
wire v_52771;
wire v_52772;
wire v_52773;
wire v_52774;
wire v_52775;
wire v_52776;
wire v_52777;
wire v_52778;
wire v_52779;
wire v_52780;
wire v_52781;
wire v_52782;
wire v_52783;
wire v_52784;
wire v_52785;
wire v_52786;
wire v_52787;
wire v_52788;
wire v_52789;
wire v_52790;
wire v_52791;
wire v_52792;
wire v_52793;
wire v_52794;
wire v_52795;
wire v_52796;
wire v_52797;
wire v_52798;
wire v_52799;
wire v_52800;
wire v_52801;
wire v_52802;
wire v_52803;
wire v_52804;
wire v_52805;
wire v_52806;
wire v_52807;
wire v_52808;
wire v_52809;
wire v_52810;
wire v_52811;
wire v_52812;
wire v_52813;
wire v_52814;
wire v_52815;
wire v_52816;
wire v_52817;
wire v_52818;
wire v_52819;
wire v_52820;
wire v_52821;
wire v_52822;
wire v_52823;
wire v_52824;
wire v_52825;
wire v_52826;
wire v_52827;
wire v_52828;
wire v_52829;
wire v_52830;
wire v_52831;
wire v_52832;
wire v_52833;
wire v_52834;
wire v_52835;
wire v_52836;
wire v_52837;
wire v_52838;
wire v_52839;
wire v_52840;
wire v_52841;
wire v_52842;
wire v_52843;
wire v_52844;
wire v_52845;
wire v_52846;
wire v_52847;
wire v_52848;
wire v_52849;
wire v_52850;
wire v_52851;
wire v_52852;
wire v_52853;
wire v_52854;
wire v_52855;
wire v_52856;
wire v_52857;
wire v_52858;
wire v_52859;
wire v_52860;
wire v_52861;
wire v_52862;
wire v_52863;
wire v_52864;
wire v_52865;
wire v_52866;
wire v_52867;
wire v_52868;
wire v_52869;
wire v_52870;
wire v_52871;
wire v_52872;
wire v_52873;
wire v_52874;
wire v_52875;
wire v_52876;
wire v_52877;
wire v_52878;
wire v_52879;
wire v_52880;
wire v_52881;
wire v_52882;
wire v_52883;
wire v_52884;
wire v_52885;
wire v_52886;
wire v_52887;
wire v_52888;
wire v_52889;
wire v_52890;
wire v_52891;
wire v_52892;
wire v_52893;
wire v_52894;
wire v_52895;
wire v_52896;
wire v_52897;
wire v_52898;
wire v_52899;
wire v_52900;
wire v_52901;
wire v_52902;
wire v_52903;
wire v_52904;
wire v_52905;
wire v_52906;
wire v_52907;
wire v_52908;
wire v_52909;
wire v_52910;
wire v_52911;
wire v_52912;
wire v_52913;
wire v_52914;
wire v_52915;
wire v_52916;
wire v_52917;
wire v_52918;
wire v_52919;
wire v_52920;
wire v_52921;
wire v_52922;
wire v_52923;
wire v_52924;
wire v_52925;
wire v_52926;
wire v_52927;
wire v_52928;
wire v_52929;
wire v_52930;
wire v_52931;
wire v_52932;
wire v_52933;
wire v_52934;
wire v_52935;
wire v_52936;
wire v_52937;
wire v_52938;
wire v_52939;
wire v_52940;
wire v_52941;
wire v_52942;
wire v_52943;
wire v_52944;
wire v_52945;
wire v_52946;
wire v_52947;
wire v_52948;
wire v_52949;
wire v_52950;
wire v_52951;
wire v_52952;
wire v_52953;
wire v_52954;
wire v_52955;
wire v_52956;
wire v_52957;
wire v_52958;
wire v_52959;
wire v_52960;
wire v_52961;
wire v_52962;
wire v_52963;
wire v_52964;
wire v_52965;
wire v_52966;
wire v_52967;
wire v_52968;
wire v_52969;
wire v_52970;
wire v_52971;
wire v_52972;
wire v_52973;
wire v_52974;
wire v_52975;
wire v_52976;
wire v_52977;
wire v_52978;
wire v_52979;
wire v_52980;
wire v_52981;
wire v_52982;
wire v_52983;
wire v_52984;
wire v_52985;
wire v_52986;
wire v_52987;
wire v_52988;
wire v_52989;
wire v_52990;
wire v_52991;
wire v_52992;
wire v_52993;
wire v_52994;
wire v_52995;
wire v_52996;
wire v_52997;
wire v_52998;
wire v_52999;
wire v_53000;
wire v_53001;
wire v_53002;
wire v_53004;
wire v_53005;
wire v_53006;
wire v_53007;
wire v_53008;
wire v_53009;
wire v_53010;
wire v_53011;
wire v_53012;
wire v_53013;
wire v_53014;
wire v_53015;
wire v_53016;
wire v_53017;
wire v_53018;
wire v_53019;
wire v_53020;
wire v_53021;
wire v_53022;
wire v_53023;
wire v_53024;
wire v_53025;
wire v_53026;
wire v_53027;
wire v_53028;
wire v_53029;
wire v_53030;
wire v_53031;
wire v_53032;
wire v_53033;
wire v_53034;
wire v_53035;
wire v_53036;
wire v_53037;
wire v_53038;
wire v_53039;
wire v_53040;
wire v_53041;
wire v_53042;
wire v_53043;
wire v_53044;
wire v_53045;
wire v_53046;
wire v_53047;
wire v_53048;
wire v_53049;
wire v_53050;
wire v_53051;
wire v_53052;
wire v_53053;
wire v_53054;
wire v_53055;
wire v_53056;
wire v_53057;
wire v_53058;
wire v_53059;
wire v_53060;
wire v_53061;
wire v_53062;
wire v_53063;
wire v_53064;
wire v_53065;
wire v_53066;
wire v_53067;
wire v_53068;
wire v_53069;
wire v_53070;
wire v_53071;
wire v_53072;
wire v_53073;
wire v_53074;
wire v_53075;
wire v_53076;
wire v_53077;
wire v_53078;
wire v_53079;
wire v_53080;
wire v_53081;
wire v_53082;
wire v_53083;
wire v_53084;
wire v_53085;
wire v_53086;
wire v_53087;
wire v_53088;
wire v_53089;
wire v_53090;
wire v_53091;
wire v_53092;
wire v_53093;
wire v_53094;
wire v_53095;
wire v_53096;
wire v_53097;
wire v_53098;
wire v_53099;
wire v_53100;
wire v_53101;
wire v_53102;
wire v_53103;
wire v_53104;
wire v_53105;
wire v_53106;
wire v_53107;
wire v_53108;
wire v_53109;
wire v_53110;
wire v_53111;
wire v_53112;
wire v_53113;
wire v_53114;
wire v_53115;
wire v_53116;
wire v_53117;
wire v_53118;
wire v_53119;
wire v_53120;
wire v_53121;
wire v_53122;
wire v_53123;
wire v_53124;
wire v_53125;
wire v_53126;
wire v_53127;
wire v_53128;
wire v_53129;
wire v_53130;
wire v_53131;
wire v_53132;
wire v_53133;
wire v_53134;
wire v_53135;
wire v_53136;
wire v_53137;
wire v_53138;
wire v_53139;
wire v_53140;
wire v_53141;
wire v_53142;
wire v_53143;
wire v_53144;
wire v_53145;
wire v_53146;
wire v_53147;
wire v_53148;
wire v_53149;
wire v_53150;
wire v_53151;
wire v_53152;
wire v_53153;
wire v_53154;
wire v_53155;
wire v_53156;
wire v_53157;
wire v_53158;
wire v_53159;
wire v_53160;
wire v_53161;
wire v_53162;
wire v_53163;
wire v_53164;
wire v_53165;
wire v_53166;
wire v_53167;
wire v_53168;
wire v_53169;
wire v_53170;
wire v_53171;
wire v_53172;
wire v_53173;
wire v_53174;
wire v_53175;
wire v_53176;
wire v_53177;
wire v_53178;
wire v_53179;
wire v_53180;
wire v_53181;
wire v_53182;
wire v_53183;
wire v_53184;
wire v_53185;
wire v_53186;
wire v_53187;
wire v_53188;
wire v_53189;
wire v_53190;
wire v_53191;
wire v_53192;
wire v_53193;
wire v_53194;
wire v_53195;
wire v_53196;
wire v_53197;
wire v_53198;
wire v_53199;
wire v_53200;
wire v_53201;
wire v_53202;
wire v_53203;
wire v_53204;
wire v_53205;
wire v_53206;
wire v_53207;
wire v_53208;
wire v_53209;
wire v_53210;
wire v_53211;
wire v_53212;
wire v_53213;
wire v_53214;
wire v_53215;
wire v_53216;
wire v_53217;
wire v_53218;
wire v_53219;
wire v_53220;
wire v_53221;
wire v_53222;
wire v_53223;
wire v_53224;
wire v_53225;
wire v_53226;
wire v_53227;
wire v_53228;
wire v_53229;
wire v_53230;
wire v_53231;
wire v_53232;
wire v_53233;
wire v_53234;
wire v_53235;
wire v_53236;
wire v_53237;
wire v_53238;
wire v_53239;
wire v_53240;
wire v_53241;
wire v_53242;
wire v_53243;
wire v_53244;
wire v_53245;
wire v_53247;
wire v_53248;
wire v_53249;
wire v_53250;
wire v_53251;
wire v_53252;
wire v_53253;
wire v_53254;
wire v_53255;
wire v_53256;
wire v_53257;
wire v_53258;
wire v_53259;
wire v_53260;
wire v_53261;
wire v_53262;
wire v_53263;
wire v_53264;
wire v_53265;
wire v_53266;
wire v_53267;
wire v_53268;
wire v_53269;
wire v_53270;
wire v_53271;
wire v_53272;
wire v_53273;
wire v_53274;
wire v_53275;
wire v_53276;
wire v_53277;
wire v_53278;
wire v_53279;
wire v_53280;
wire v_53281;
wire v_53282;
wire v_53283;
wire v_53284;
wire v_53285;
wire v_53286;
wire v_53287;
wire v_53288;
wire v_53289;
wire v_53290;
wire v_53291;
wire v_53292;
wire v_53293;
wire v_53294;
wire v_53295;
wire v_53296;
wire v_53297;
wire v_53298;
wire v_53299;
wire v_53300;
wire v_53301;
wire v_53302;
wire v_53303;
wire v_53304;
wire v_53305;
wire v_53306;
wire v_53307;
wire v_53308;
wire v_53309;
wire v_53310;
wire v_53311;
wire v_53312;
wire v_53313;
wire v_53314;
wire v_53315;
wire v_53316;
wire v_53317;
wire v_53318;
wire v_53319;
wire v_53320;
wire v_53321;
wire v_53322;
wire v_53323;
wire v_53324;
wire v_53325;
wire v_53326;
wire v_53327;
wire v_53328;
wire v_53329;
wire v_53330;
wire v_53331;
wire v_53332;
wire v_53333;
wire v_53334;
wire v_53335;
wire v_53336;
wire v_53337;
wire v_53338;
wire v_53339;
wire v_53340;
wire v_53341;
wire v_53342;
wire v_53343;
wire v_53344;
wire v_53345;
wire v_53346;
wire v_53347;
wire v_53348;
wire v_53349;
wire v_53350;
wire v_53351;
wire v_53352;
wire v_53353;
wire v_53354;
wire v_53355;
wire v_53356;
wire v_53357;
wire v_53358;
wire v_53359;
wire v_53360;
wire v_53361;
wire v_53362;
wire v_53363;
wire v_53364;
wire v_53365;
wire v_53366;
wire v_53367;
wire v_53368;
wire v_53369;
wire v_53370;
wire v_53371;
wire v_53372;
wire v_53373;
wire v_53374;
wire v_53375;
wire v_53376;
wire v_53377;
wire v_53378;
wire v_53379;
wire v_53380;
wire v_53381;
wire v_53382;
wire v_53383;
wire v_53384;
wire v_53385;
wire v_53386;
wire v_53387;
wire v_53388;
wire v_53389;
wire v_53390;
wire v_53391;
wire v_53392;
wire v_53393;
wire v_53394;
wire v_53395;
wire v_53396;
wire v_53397;
wire v_53398;
wire v_53399;
wire v_53400;
wire v_53401;
wire v_53402;
wire v_53403;
wire v_53404;
wire v_53405;
wire v_53406;
wire v_53407;
wire v_53408;
wire v_53409;
wire v_53410;
wire v_53411;
wire v_53412;
wire v_53413;
wire v_53414;
wire v_53415;
wire v_53416;
wire v_53417;
wire v_53418;
wire v_53419;
wire v_53420;
wire v_53421;
wire v_53422;
wire v_53423;
wire v_53424;
wire v_53425;
wire v_53426;
wire v_53427;
wire v_53428;
wire v_53429;
wire v_53430;
wire v_53431;
wire v_53432;
wire v_53433;
wire v_53434;
wire v_53435;
wire v_53436;
wire v_53437;
wire v_53438;
wire v_53439;
wire v_53440;
wire v_53441;
wire v_53442;
wire v_53443;
wire v_53444;
wire v_53445;
wire v_53446;
wire v_53447;
wire v_53448;
wire v_53449;
wire v_53450;
wire v_53451;
wire v_53452;
wire v_53453;
wire v_53454;
wire v_53455;
wire v_53456;
wire v_53457;
wire v_53458;
wire v_53459;
wire v_53460;
wire v_53461;
wire v_53462;
wire v_53463;
wire v_53464;
wire v_53465;
wire v_53466;
wire v_53467;
wire v_53468;
wire v_53469;
wire v_53470;
wire v_53471;
wire v_53472;
wire v_53473;
wire v_53474;
wire v_53475;
wire v_53476;
wire v_53477;
wire v_53478;
wire v_53479;
wire v_53480;
wire v_53481;
wire v_53482;
wire v_53483;
wire v_53484;
wire v_53485;
wire v_53486;
wire v_53487;
wire v_53488;
wire v_53490;
wire v_53491;
wire v_53492;
wire v_53493;
wire v_53494;
wire v_53495;
wire v_53496;
wire v_53497;
wire v_53498;
wire v_53499;
wire v_53500;
wire v_53501;
wire v_53502;
wire v_53503;
wire v_53504;
wire v_53505;
wire v_53506;
wire v_53507;
wire v_53508;
wire v_53509;
wire v_53510;
wire v_53511;
wire v_53512;
wire v_53513;
wire v_53514;
wire v_53515;
wire v_53516;
wire v_53517;
wire v_53518;
wire v_53519;
wire v_53520;
wire v_53521;
wire v_53522;
wire v_53523;
wire v_53524;
wire v_53525;
wire v_53526;
wire v_53527;
wire v_53528;
wire v_53529;
wire v_53530;
wire v_53531;
wire v_53532;
wire v_53533;
wire v_53534;
wire v_53535;
wire v_53536;
wire v_53537;
wire v_53538;
wire v_53539;
wire v_53540;
wire v_53541;
wire v_53542;
wire v_53543;
wire v_53544;
wire v_53545;
wire v_53546;
wire v_53547;
wire v_53548;
wire v_53549;
wire v_53550;
wire v_53551;
wire v_53552;
wire v_53553;
wire v_53554;
wire v_53555;
wire v_53556;
wire v_53557;
wire v_53558;
wire v_53559;
wire v_53560;
wire v_53561;
wire v_53562;
wire v_53563;
wire v_53564;
wire v_53565;
wire v_53566;
wire v_53567;
wire v_53568;
wire v_53569;
wire v_53570;
wire v_53571;
wire v_53572;
wire v_53573;
wire v_53574;
wire v_53575;
wire v_53576;
wire v_53577;
wire v_53578;
wire v_53579;
wire v_53580;
wire v_53581;
wire v_53582;
wire v_53583;
wire v_53584;
wire v_53585;
wire v_53586;
wire v_53587;
wire v_53588;
wire v_53589;
wire v_53590;
wire v_53591;
wire v_53592;
wire v_53593;
wire v_53594;
wire v_53595;
wire v_53596;
wire v_53597;
wire v_53598;
wire v_53599;
wire v_53600;
wire v_53601;
wire v_53602;
wire v_53603;
wire v_53604;
wire v_53605;
wire v_53606;
wire v_53607;
wire v_53608;
wire v_53609;
wire v_53610;
wire v_53611;
wire v_53612;
wire v_53613;
wire v_53614;
wire v_53615;
wire v_53616;
wire v_53617;
wire v_53618;
wire v_53619;
wire v_53620;
wire v_53621;
wire v_53622;
wire v_53623;
wire v_53624;
wire v_53625;
wire v_53626;
wire v_53627;
wire v_53628;
wire v_53629;
wire v_53630;
wire v_53631;
wire v_53632;
wire v_53633;
wire v_53634;
wire v_53635;
wire v_53636;
wire v_53637;
wire v_53638;
wire v_53639;
wire v_53640;
wire v_53641;
wire v_53642;
wire v_53643;
wire v_53644;
wire v_53645;
wire v_53646;
wire v_53647;
wire v_53648;
wire v_53649;
wire v_53650;
wire v_53651;
wire v_53652;
wire v_53653;
wire v_53654;
wire v_53655;
wire v_53656;
wire v_53657;
wire v_53658;
wire v_53659;
wire v_53660;
wire v_53661;
wire v_53662;
wire v_53663;
wire v_53664;
wire v_53665;
wire v_53666;
wire v_53667;
wire v_53668;
wire v_53669;
wire v_53670;
wire v_53671;
wire v_53672;
wire v_53673;
wire v_53674;
wire v_53675;
wire v_53676;
wire v_53677;
wire v_53678;
wire v_53679;
wire v_53680;
wire v_53681;
wire v_53682;
wire v_53683;
wire v_53684;
wire v_53685;
wire v_53686;
wire v_53687;
wire v_53688;
wire v_53689;
wire v_53690;
wire v_53691;
wire v_53692;
wire v_53693;
wire v_53694;
wire v_53695;
wire v_53696;
wire v_53697;
wire v_53698;
wire v_53699;
wire v_53700;
wire v_53701;
wire v_53702;
wire v_53703;
wire v_53704;
wire v_53705;
wire v_53706;
wire v_53707;
wire v_53708;
wire v_53709;
wire v_53710;
wire v_53711;
wire v_53712;
wire v_53713;
wire v_53714;
wire v_53715;
wire v_53716;
wire v_53717;
wire v_53718;
wire v_53719;
wire v_53720;
wire v_53721;
wire v_53722;
wire v_53723;
wire v_53724;
wire v_53725;
wire v_53726;
wire v_53727;
wire v_53728;
wire v_53729;
wire v_53730;
wire v_53731;
wire v_53733;
wire v_53734;
wire v_53735;
wire v_53736;
wire v_53737;
wire v_53738;
wire v_53739;
wire v_53740;
wire v_53741;
wire v_53742;
wire v_53743;
wire v_53744;
wire v_53745;
wire v_53746;
wire v_53747;
wire v_53748;
wire v_53749;
wire v_53750;
wire v_53751;
wire v_53752;
wire v_53753;
wire v_53754;
wire v_53755;
wire v_53756;
wire v_53757;
wire v_53758;
wire v_53759;
wire v_53760;
wire v_53761;
wire v_53762;
wire v_53763;
wire v_53764;
wire v_53765;
wire v_53766;
wire v_53767;
wire v_53768;
wire v_53769;
wire v_53770;
wire v_53771;
wire v_53772;
wire v_53773;
wire v_53774;
wire v_53775;
wire v_53776;
wire v_53777;
wire v_53778;
wire v_53779;
wire v_53780;
wire v_53781;
wire v_53782;
wire v_53783;
wire v_53784;
wire v_53785;
wire v_53786;
wire v_53787;
wire v_53788;
wire v_53789;
wire v_53790;
wire v_53791;
wire v_53792;
wire v_53793;
wire v_53794;
wire v_53795;
wire v_53796;
wire v_53797;
wire v_53798;
wire v_53799;
wire v_53800;
wire v_53801;
wire v_53802;
wire v_53803;
wire v_53804;
wire v_53805;
wire v_53806;
wire v_53807;
wire v_53808;
wire v_53809;
wire v_53810;
wire v_53811;
wire v_53812;
wire v_53813;
wire v_53814;
wire v_53815;
wire v_53816;
wire v_53817;
wire v_53818;
wire v_53819;
wire v_53820;
wire v_53821;
wire v_53822;
wire v_53823;
wire v_53824;
wire v_53825;
wire v_53826;
wire v_53827;
wire v_53828;
wire v_53829;
wire v_53830;
wire v_53831;
wire v_53832;
wire v_53833;
wire v_53834;
wire v_53835;
wire v_53836;
wire v_53837;
wire v_53838;
wire v_53839;
wire v_53840;
wire v_53841;
wire v_53842;
wire v_53843;
wire v_53844;
wire v_53845;
wire v_53846;
wire v_53847;
wire v_53848;
wire v_53849;
wire v_53850;
wire v_53851;
wire v_53852;
wire v_53853;
wire v_53854;
wire v_53855;
wire v_53856;
wire v_53857;
wire v_53858;
wire v_53859;
wire v_53860;
wire v_53861;
wire v_53862;
wire v_53863;
wire v_53864;
wire v_53865;
wire v_53866;
wire v_53867;
wire v_53868;
wire v_53869;
wire v_53870;
wire v_53871;
wire v_53872;
wire v_53873;
wire v_53874;
wire v_53875;
wire v_53876;
wire v_53877;
wire v_53878;
wire v_53879;
wire v_53880;
wire v_53881;
wire v_53882;
wire v_53883;
wire v_53884;
wire v_53885;
wire v_53886;
wire v_53887;
wire v_53888;
wire v_53889;
wire v_53890;
wire v_53891;
wire v_53892;
wire v_53893;
wire v_53894;
wire v_53895;
wire v_53896;
wire v_53897;
wire v_53898;
wire v_53899;
wire v_53900;
wire v_53901;
wire v_53902;
wire v_53903;
wire v_53904;
wire v_53905;
wire v_53906;
wire v_53907;
wire v_53908;
wire v_53909;
wire v_53910;
wire v_53911;
wire v_53912;
wire v_53913;
wire v_53914;
wire v_53915;
wire v_53916;
wire v_53917;
wire v_53918;
wire v_53919;
wire v_53920;
wire v_53921;
wire v_53922;
wire v_53923;
wire v_53924;
wire v_53925;
wire v_53926;
wire v_53927;
wire v_53928;
wire v_53929;
wire v_53930;
wire v_53931;
wire v_53932;
wire v_53933;
wire v_53934;
wire v_53935;
wire v_53936;
wire v_53937;
wire v_53938;
wire v_53939;
wire v_53940;
wire v_53941;
wire v_53942;
wire v_53943;
wire v_53944;
wire v_53945;
wire v_53946;
wire v_53947;
wire v_53948;
wire v_53949;
wire v_53950;
wire v_53951;
wire v_53952;
wire v_53953;
wire v_53954;
wire v_53955;
wire v_53956;
wire v_53957;
wire v_53958;
wire v_53959;
wire v_53960;
wire v_53961;
wire v_53962;
wire v_53963;
wire v_53964;
wire v_53965;
wire v_53966;
wire v_53967;
wire v_53968;
wire v_53969;
wire v_53970;
wire v_53971;
wire v_53972;
wire v_53973;
wire v_53974;
wire v_53975;
wire v_53976;
wire v_53977;
wire v_53978;
wire v_53979;
wire v_53980;
wire v_53981;
wire v_53982;
wire v_53983;
wire v_53984;
wire v_53985;
wire v_53986;
wire v_53987;
wire v_53988;
wire v_53989;
wire v_53990;
wire v_53991;
wire v_53992;
wire v_53993;
wire v_53994;
wire v_53995;
wire v_53996;
wire v_53997;
wire v_53998;
wire v_53999;
wire v_54000;
wire v_54001;
wire v_54002;
wire v_54003;
wire v_54004;
wire v_54005;
wire v_54006;
wire v_54007;
wire v_54008;
wire v_54009;
wire v_54010;
wire v_54011;
wire v_54012;
wire v_54013;
wire v_54014;
wire v_54015;
wire v_54016;
wire v_54017;
wire v_54018;
wire v_54019;
wire v_54020;
wire v_54021;
wire v_54022;
wire v_54023;
wire v_54024;
wire v_54025;
wire v_54026;
wire v_54027;
wire v_54028;
wire v_54029;
wire v_54030;
wire v_54031;
wire v_54032;
wire v_54033;
wire v_54034;
wire v_54035;
wire v_54036;
wire v_54037;
wire v_54038;
wire v_54039;
wire v_54040;
wire v_54041;
wire v_54042;
wire v_54043;
wire v_54044;
wire v_54045;
wire v_54046;
wire v_54047;
wire v_54048;
wire v_54049;
wire v_54050;
wire v_54051;
wire v_54052;
wire v_54053;
wire v_54054;
wire v_54055;
wire v_54056;
wire v_54057;
wire v_54058;
wire v_54059;
wire v_54060;
wire v_54061;
wire v_54062;
wire v_54063;
wire v_54064;
wire v_54065;
wire v_54066;
wire v_54067;
wire v_54068;
wire v_54069;
wire v_54070;
wire v_54071;
wire v_54072;
wire v_54073;
wire v_54074;
wire v_54075;
wire v_54076;
wire v_54077;
wire v_54078;
wire v_54079;
wire v_54080;
wire v_54081;
wire v_54082;
wire v_54083;
wire v_54084;
wire v_54085;
wire v_54086;
wire v_54087;
wire v_54088;
wire v_54089;
wire v_54090;
wire v_54091;
wire v_54092;
wire v_54093;
wire v_54094;
wire v_54095;
wire v_54096;
wire v_54097;
wire v_54098;
wire v_54099;
wire v_54100;
wire v_54101;
wire v_54102;
wire v_54103;
wire v_54104;
wire v_54105;
wire v_54106;
wire v_54107;
wire v_54108;
wire v_54109;
wire v_54110;
wire v_54111;
wire v_54112;
wire v_54113;
wire v_54114;
wire v_54115;
wire v_54116;
wire v_54117;
wire v_54118;
wire v_54119;
wire v_54120;
wire v_54121;
wire v_54122;
wire v_54123;
wire v_54125;
wire v_54126;
wire v_54127;
wire v_54128;
wire v_54129;
wire v_54130;
wire v_54131;
wire v_54132;
wire v_54133;
wire v_54134;
wire v_54135;
wire v_54136;
wire v_54137;
wire v_54138;
wire v_54139;
wire v_54140;
wire v_54141;
wire v_54142;
wire v_54143;
wire v_54144;
wire v_54145;
wire v_54146;
wire v_54147;
wire v_54148;
wire v_54149;
wire v_54150;
wire v_54151;
wire v_54152;
wire v_54153;
wire v_54154;
wire v_54155;
wire v_54156;
wire v_54157;
wire v_54158;
wire v_54159;
wire v_54160;
wire v_54161;
wire v_54162;
wire v_54163;
wire v_54164;
wire v_54165;
wire v_54166;
wire v_54167;
wire v_54168;
wire v_54169;
wire v_54170;
wire v_54171;
wire v_54172;
wire v_54173;
wire v_54174;
wire v_54175;
wire v_54176;
wire v_54177;
wire v_54178;
wire v_54179;
wire v_54180;
wire v_54181;
wire v_54182;
wire v_54183;
wire v_54184;
wire v_54185;
wire v_54186;
wire v_54187;
wire v_54188;
wire v_54189;
wire v_54190;
wire v_54191;
wire v_54192;
wire v_54193;
wire v_54194;
wire v_54195;
wire v_54196;
wire v_54197;
wire v_54198;
wire v_54199;
wire v_54200;
wire v_54201;
wire v_54202;
wire v_54203;
wire v_54204;
wire v_54205;
wire v_54206;
wire v_54207;
wire v_54208;
wire v_54209;
wire v_54210;
wire v_54211;
wire v_54212;
wire v_54213;
wire v_54214;
wire v_54215;
wire v_54216;
wire v_54217;
wire v_54219;
wire v_54221;
wire v_54222;
wire v_54223;
wire v_54225;
wire v_54226;
wire v_54227;
wire v_54229;
wire v_54230;
wire v_54231;
wire v_54233;
wire v_54234;
wire v_54236;
wire v_54237;
wire v_54238;
wire v_54240;
wire v_54241;
wire v_54242;
wire v_54244;
wire v_54245;
wire v_54246;
wire v_54248;
wire v_54249;
wire v_54250;
wire v_54252;
wire v_54253;
wire v_54254;
wire v_54256;
wire v_54257;
wire v_54258;
wire v_54260;
wire v_54261;
wire v_54262;
wire v_54264;
wire v_54265;
wire v_54266;
wire v_54268;
wire v_54269;
wire v_54270;
wire v_54272;
wire v_54273;
wire v_54274;
wire v_54276;
wire v_54277;
wire v_54278;
wire v_54280;
wire v_54281;
wire v_54282;
wire v_54284;
wire v_54285;
wire v_54286;
wire v_54287;
wire v_54288;
wire v_54289;
wire v_54290;
wire v_54291;
wire v_54292;
wire v_54293;
wire v_54294;
wire v_54295;
wire v_54296;
wire v_54297;
wire v_54298;
wire v_54299;
wire v_54300;
wire v_54301;
wire v_54302;
wire v_54303;
wire v_54304;
wire v_54305;
wire v_54306;
wire v_54307;
wire v_54308;
wire v_54309;
wire v_54310;
wire v_54311;
wire v_54312;
wire v_54313;
wire v_54314;
wire v_54315;
wire v_54316;
wire v_54317;
wire v_54318;
wire v_54319;
wire v_54320;
wire v_54321;
wire v_54322;
wire v_54323;
wire v_54324;
wire v_54325;
wire v_54326;
wire v_54327;
wire v_54328;
wire v_54329;
wire v_54330;
wire v_54331;
wire v_54332;
wire v_54333;
wire v_54334;
wire v_54335;
wire v_54336;
wire v_54337;
wire v_54338;
wire v_54339;
wire v_54340;
wire v_54341;
wire v_54342;
wire v_54343;
wire v_54344;
wire v_54345;
wire v_54346;
wire v_54347;
wire v_54348;
wire v_54349;
wire v_54350;
wire v_54351;
wire v_54352;
wire v_54353;
wire v_54354;
wire v_54355;
wire v_54356;
wire v_54357;
wire v_54358;
wire v_54359;
wire v_54360;
wire v_54361;
wire v_54362;
wire v_54363;
wire v_54364;
wire v_54365;
wire v_54366;
wire v_54367;
wire v_54368;
wire v_54369;
wire v_54370;
wire v_54371;
wire v_54372;
wire v_54373;
wire v_54374;
wire v_54375;
wire v_54376;
wire v_54377;
wire v_54378;
wire v_54379;
wire v_54380;
wire v_54381;
wire v_54382;
wire v_54383;
wire v_54384;
wire v_54385;
wire v_54386;
wire v_54387;
wire v_54388;
wire v_54389;
wire v_54390;
wire v_54391;
wire v_54392;
wire v_54393;
wire v_54394;
wire v_54395;
wire v_54396;
wire v_54397;
wire v_54398;
wire v_54399;
wire v_54400;
wire v_54401;
wire v_54402;
wire v_54403;
wire v_54404;
wire v_54405;
wire v_54406;
wire v_54407;
wire v_54408;
wire v_54409;
wire v_54410;
wire v_54411;
wire v_54412;
wire v_54413;
wire v_54414;
wire v_54415;
wire v_54416;
wire v_54417;
wire v_54418;
wire v_54419;
wire v_54420;
wire v_54421;
wire v_54422;
wire v_54423;
wire v_54424;
wire v_54425;
wire v_54426;
wire v_54427;
wire v_54428;
wire v_54429;
wire v_54430;
wire v_54431;
wire v_54432;
wire v_54433;
wire v_54434;
wire v_54435;
wire v_54436;
wire v_54437;
wire v_54438;
wire v_54439;
wire v_54440;
wire v_54441;
wire v_54442;
wire v_54443;
wire v_54444;
wire v_54445;
wire v_54446;
wire v_54447;
wire v_54448;
wire v_54449;
wire v_54450;
wire v_54451;
wire v_54452;
wire v_54453;
wire v_54454;
wire v_54455;
wire v_54456;
wire v_54457;
wire v_54458;
wire v_54459;
wire v_54460;
wire v_54461;
wire v_54462;
wire v_54463;
wire v_54464;
wire v_54465;
wire v_54466;
wire v_54467;
wire v_54468;
wire v_54469;
wire v_54470;
wire v_54471;
wire v_54472;
wire v_54473;
wire v_54474;
wire v_54475;
wire v_54476;
wire v_54477;
wire v_54479;
wire v_54480;
wire v_54481;
wire v_54482;
wire v_54483;
wire v_54484;
wire v_54485;
wire v_54486;
wire v_54487;
wire v_54488;
wire v_54489;
wire v_54490;
wire v_54491;
wire v_54492;
wire v_54493;
wire v_54494;
wire v_54495;
wire v_54496;
wire v_54497;
wire v_54498;
wire v_54499;
wire v_54500;
wire v_54501;
wire v_54502;
wire v_54503;
wire v_54504;
wire v_54505;
wire v_54506;
wire v_54507;
wire v_54508;
wire v_54509;
wire v_54510;
wire v_54511;
wire v_54512;
wire v_54513;
wire v_54514;
wire v_54515;
wire v_54516;
wire v_54517;
wire v_54518;
wire v_54519;
wire v_54520;
wire v_54521;
wire v_54522;
wire v_54523;
wire v_54524;
wire v_54525;
wire v_54526;
wire v_54527;
wire v_54528;
wire v_54529;
wire v_54530;
wire v_54531;
wire v_54532;
wire v_54533;
wire v_54534;
wire v_54535;
wire v_54536;
wire v_54537;
wire v_54538;
wire v_54539;
wire v_54540;
wire v_54541;
wire v_54542;
wire v_54543;
wire v_54544;
wire v_54545;
wire v_54546;
wire v_54547;
wire v_54548;
wire v_54549;
wire v_54550;
wire v_54551;
wire v_54552;
wire v_54553;
wire v_54554;
wire v_54555;
wire v_54556;
wire v_54557;
wire v_54558;
wire v_54559;
wire v_54560;
wire v_54561;
wire v_54562;
wire v_54563;
wire v_54564;
wire v_54565;
wire v_54566;
wire v_54567;
wire v_54568;
wire v_54569;
wire v_54570;
wire v_54571;
wire v_54572;
wire v_54573;
wire v_54574;
wire v_54575;
wire v_54576;
wire v_54577;
wire v_54578;
wire v_54579;
wire v_54580;
wire v_54581;
wire v_54582;
wire v_54583;
wire v_54584;
wire v_54585;
wire v_54586;
wire v_54587;
wire v_54588;
wire v_54589;
wire v_54590;
wire v_54591;
wire v_54592;
wire v_54593;
wire v_54594;
wire v_54595;
wire v_54596;
wire v_54597;
wire v_54598;
wire v_54599;
wire v_54600;
wire v_54601;
wire v_54602;
wire v_54603;
wire v_54604;
wire v_54605;
wire v_54606;
wire v_54607;
wire v_54608;
wire v_54609;
wire v_54610;
wire v_54611;
wire v_54612;
wire v_54613;
wire v_54614;
wire v_54615;
wire v_54616;
wire v_54617;
wire v_54618;
wire v_54619;
wire v_54620;
wire v_54621;
wire v_54622;
wire v_54623;
wire v_54624;
wire v_54625;
wire v_54626;
wire v_54627;
wire v_54628;
wire v_54629;
wire v_54630;
wire v_54631;
wire v_54632;
wire v_54633;
wire v_54634;
wire v_54635;
wire v_54636;
wire v_54637;
wire v_54638;
wire v_54639;
wire v_54640;
wire v_54641;
wire v_54642;
wire v_54643;
wire v_54644;
wire v_54645;
wire v_54646;
wire v_54647;
wire v_54648;
wire v_54649;
wire v_54650;
wire v_54651;
wire v_54652;
wire v_54653;
wire v_54654;
wire v_54655;
wire v_54656;
wire v_54657;
wire v_54658;
wire v_54659;
wire v_54660;
wire v_54661;
wire v_54662;
wire v_54663;
wire v_54664;
wire v_54665;
wire v_54666;
wire v_54667;
wire v_54668;
wire v_54669;
wire v_54670;
wire v_54671;
wire v_54672;
wire v_54673;
wire v_54674;
wire v_54675;
wire v_54676;
wire v_54677;
wire v_54678;
wire v_54679;
wire v_54680;
wire v_54681;
wire v_54682;
wire v_54683;
wire v_54684;
wire v_54685;
wire v_54686;
wire v_54687;
wire v_54688;
wire v_54689;
wire v_54690;
wire v_54691;
wire v_54692;
wire v_54693;
wire v_54694;
wire v_54695;
wire v_54696;
wire v_54697;
wire v_54698;
wire v_54699;
wire v_54700;
wire v_54701;
wire v_54702;
wire v_54703;
wire v_54704;
wire v_54705;
wire v_54706;
wire v_54707;
wire v_54708;
wire v_54709;
wire v_54710;
wire v_54711;
wire v_54712;
wire v_54713;
wire v_54714;
wire v_54715;
wire v_54716;
wire v_54717;
wire v_54718;
wire v_54719;
wire v_54720;
wire v_54722;
wire v_54723;
wire v_54724;
wire v_54725;
wire v_54726;
wire v_54727;
wire v_54728;
wire v_54729;
wire v_54730;
wire v_54731;
wire v_54732;
wire v_54733;
wire v_54734;
wire v_54735;
wire v_54736;
wire v_54737;
wire v_54738;
wire v_54739;
wire v_54740;
wire v_54741;
wire v_54742;
wire v_54743;
wire v_54744;
wire v_54745;
wire v_54746;
wire v_54747;
wire v_54748;
wire v_54749;
wire v_54750;
wire v_54751;
wire v_54752;
wire v_54753;
wire v_54754;
wire v_54755;
wire v_54756;
wire v_54757;
wire v_54758;
wire v_54759;
wire v_54760;
wire v_54761;
wire v_54762;
wire v_54763;
wire v_54764;
wire v_54765;
wire v_54766;
wire v_54767;
wire v_54768;
wire v_54769;
wire v_54770;
wire v_54771;
wire v_54772;
wire v_54773;
wire v_54774;
wire v_54775;
wire v_54776;
wire v_54777;
wire v_54778;
wire v_54779;
wire v_54780;
wire v_54781;
wire v_54782;
wire v_54783;
wire v_54784;
wire v_54785;
wire v_54786;
wire v_54787;
wire v_54788;
wire v_54789;
wire v_54790;
wire v_54791;
wire v_54792;
wire v_54793;
wire v_54794;
wire v_54795;
wire v_54796;
wire v_54797;
wire v_54798;
wire v_54799;
wire v_54800;
wire v_54801;
wire v_54802;
wire v_54803;
wire v_54804;
wire v_54805;
wire v_54806;
wire v_54807;
wire v_54808;
wire v_54809;
wire v_54810;
wire v_54811;
wire v_54812;
wire v_54813;
wire v_54814;
wire v_54815;
wire v_54816;
wire v_54817;
wire v_54818;
wire v_54819;
wire v_54820;
wire v_54821;
wire v_54822;
wire v_54823;
wire v_54824;
wire v_54825;
wire v_54826;
wire v_54827;
wire v_54828;
wire v_54829;
wire v_54830;
wire v_54831;
wire v_54832;
wire v_54833;
wire v_54834;
wire v_54835;
wire v_54836;
wire v_54837;
wire v_54838;
wire v_54839;
wire v_54840;
wire v_54841;
wire v_54842;
wire v_54843;
wire v_54844;
wire v_54845;
wire v_54846;
wire v_54847;
wire v_54848;
wire v_54849;
wire v_54850;
wire v_54851;
wire v_54852;
wire v_54853;
wire v_54854;
wire v_54855;
wire v_54856;
wire v_54857;
wire v_54858;
wire v_54859;
wire v_54860;
wire v_54861;
wire v_54862;
wire v_54863;
wire v_54864;
wire v_54865;
wire v_54866;
wire v_54867;
wire v_54868;
wire v_54869;
wire v_54870;
wire v_54871;
wire v_54872;
wire v_54873;
wire v_54874;
wire v_54875;
wire v_54876;
wire v_54877;
wire v_54878;
wire v_54879;
wire v_54880;
wire v_54881;
wire v_54882;
wire v_54883;
wire v_54884;
wire v_54885;
wire v_54886;
wire v_54887;
wire v_54888;
wire v_54889;
wire v_54890;
wire v_54891;
wire v_54892;
wire v_54893;
wire v_54894;
wire v_54895;
wire v_54896;
wire v_54897;
wire v_54898;
wire v_54899;
wire v_54900;
wire v_54901;
wire v_54902;
wire v_54903;
wire v_54904;
wire v_54905;
wire v_54906;
wire v_54907;
wire v_54908;
wire v_54909;
wire v_54910;
wire v_54911;
wire v_54912;
wire v_54913;
wire v_54914;
wire v_54915;
wire v_54916;
wire v_54917;
wire v_54918;
wire v_54919;
wire v_54920;
wire v_54921;
wire v_54922;
wire v_54923;
wire v_54924;
wire v_54925;
wire v_54926;
wire v_54927;
wire v_54928;
wire v_54929;
wire v_54930;
wire v_54931;
wire v_54932;
wire v_54933;
wire v_54934;
wire v_54935;
wire v_54936;
wire v_54937;
wire v_54938;
wire v_54939;
wire v_54940;
wire v_54941;
wire v_54942;
wire v_54943;
wire v_54944;
wire v_54945;
wire v_54946;
wire v_54947;
wire v_54948;
wire v_54949;
wire v_54950;
wire v_54951;
wire v_54952;
wire v_54953;
wire v_54954;
wire v_54955;
wire v_54956;
wire v_54957;
wire v_54958;
wire v_54959;
wire v_54960;
wire v_54961;
wire v_54962;
wire v_54963;
wire v_54965;
wire v_54966;
wire v_54967;
wire v_54968;
wire v_54969;
wire v_54970;
wire v_54971;
wire v_54972;
wire v_54973;
wire v_54974;
wire v_54975;
wire v_54976;
wire v_54977;
wire v_54978;
wire v_54979;
wire v_54980;
wire v_54981;
wire v_54982;
wire v_54983;
wire v_54984;
wire v_54985;
wire v_54986;
wire v_54987;
wire v_54988;
wire v_54989;
wire v_54990;
wire v_54991;
wire v_54992;
wire v_54993;
wire v_54994;
wire v_54995;
wire v_54996;
wire v_54997;
wire v_54998;
wire v_54999;
wire v_55000;
wire v_55001;
wire v_55002;
wire v_55003;
wire v_55004;
wire v_55005;
wire v_55006;
wire v_55007;
wire v_55008;
wire v_55009;
wire v_55010;
wire v_55011;
wire v_55012;
wire v_55013;
wire v_55014;
wire v_55015;
wire v_55016;
wire v_55017;
wire v_55018;
wire v_55019;
wire v_55020;
wire v_55021;
wire v_55022;
wire v_55023;
wire v_55024;
wire v_55025;
wire v_55026;
wire v_55027;
wire v_55028;
wire v_55029;
wire v_55030;
wire v_55031;
wire v_55032;
wire v_55033;
wire v_55034;
wire v_55035;
wire v_55036;
wire v_55037;
wire v_55038;
wire v_55039;
wire v_55040;
wire v_55041;
wire v_55042;
wire v_55043;
wire v_55044;
wire v_55045;
wire v_55046;
wire v_55047;
wire v_55048;
wire v_55049;
wire v_55050;
wire v_55051;
wire v_55052;
wire v_55053;
wire v_55054;
wire v_55055;
wire v_55056;
wire v_55057;
wire v_55058;
wire v_55059;
wire v_55060;
wire v_55061;
wire v_55062;
wire v_55063;
wire v_55064;
wire v_55065;
wire v_55066;
wire v_55067;
wire v_55068;
wire v_55069;
wire v_55070;
wire v_55071;
wire v_55072;
wire v_55073;
wire v_55074;
wire v_55075;
wire v_55076;
wire v_55077;
wire v_55078;
wire v_55079;
wire v_55080;
wire v_55081;
wire v_55082;
wire v_55083;
wire v_55084;
wire v_55085;
wire v_55086;
wire v_55087;
wire v_55088;
wire v_55089;
wire v_55090;
wire v_55091;
wire v_55092;
wire v_55093;
wire v_55094;
wire v_55095;
wire v_55096;
wire v_55097;
wire v_55098;
wire v_55099;
wire v_55100;
wire v_55101;
wire v_55102;
wire v_55103;
wire v_55104;
wire v_55105;
wire v_55106;
wire v_55107;
wire v_55108;
wire v_55109;
wire v_55110;
wire v_55111;
wire v_55112;
wire v_55113;
wire v_55114;
wire v_55115;
wire v_55116;
wire v_55117;
wire v_55118;
wire v_55119;
wire v_55120;
wire v_55121;
wire v_55122;
wire v_55123;
wire v_55124;
wire v_55125;
wire v_55126;
wire v_55127;
wire v_55128;
wire v_55129;
wire v_55130;
wire v_55131;
wire v_55132;
wire v_55133;
wire v_55134;
wire v_55135;
wire v_55136;
wire v_55137;
wire v_55138;
wire v_55139;
wire v_55140;
wire v_55141;
wire v_55142;
wire v_55143;
wire v_55144;
wire v_55145;
wire v_55146;
wire v_55147;
wire v_55148;
wire v_55149;
wire v_55150;
wire v_55151;
wire v_55152;
wire v_55153;
wire v_55154;
wire v_55155;
wire v_55156;
wire v_55157;
wire v_55158;
wire v_55159;
wire v_55160;
wire v_55161;
wire v_55162;
wire v_55163;
wire v_55164;
wire v_55165;
wire v_55166;
wire v_55167;
wire v_55168;
wire v_55169;
wire v_55170;
wire v_55171;
wire v_55172;
wire v_55173;
wire v_55174;
wire v_55175;
wire v_55176;
wire v_55177;
wire v_55178;
wire v_55179;
wire v_55180;
wire v_55181;
wire v_55182;
wire v_55183;
wire v_55184;
wire v_55185;
wire v_55186;
wire v_55187;
wire v_55188;
wire v_55189;
wire v_55190;
wire v_55191;
wire v_55192;
wire v_55193;
wire v_55194;
wire v_55195;
wire v_55196;
wire v_55197;
wire v_55198;
wire v_55199;
wire v_55200;
wire v_55201;
wire v_55202;
wire v_55203;
wire v_55204;
wire v_55205;
wire v_55206;
wire v_55208;
wire v_55209;
wire v_55210;
wire v_55211;
wire v_55212;
wire v_55213;
wire v_55214;
wire v_55215;
wire v_55216;
wire v_55217;
wire v_55218;
wire v_55219;
wire v_55220;
wire v_55221;
wire v_55222;
wire v_55223;
wire v_55224;
wire v_55225;
wire v_55226;
wire v_55227;
wire v_55228;
wire v_55229;
wire v_55230;
wire v_55231;
wire v_55232;
wire v_55233;
wire v_55234;
wire v_55235;
wire v_55236;
wire v_55237;
wire v_55238;
wire v_55239;
wire v_55240;
wire v_55241;
wire v_55242;
wire v_55243;
wire v_55244;
wire v_55245;
wire v_55246;
wire v_55247;
wire v_55248;
wire v_55249;
wire v_55250;
wire v_55251;
wire v_55252;
wire v_55253;
wire v_55254;
wire v_55255;
wire v_55256;
wire v_55257;
wire v_55258;
wire v_55259;
wire v_55260;
wire v_55261;
wire v_55262;
wire v_55263;
wire v_55264;
wire v_55265;
wire v_55266;
wire v_55267;
wire v_55268;
wire v_55269;
wire v_55270;
wire v_55271;
wire v_55272;
wire v_55273;
wire v_55274;
wire v_55275;
wire v_55276;
wire v_55277;
wire v_55278;
wire v_55279;
wire v_55280;
wire v_55281;
wire v_55282;
wire v_55283;
wire v_55284;
wire v_55285;
wire v_55286;
wire v_55287;
wire v_55288;
wire v_55289;
wire v_55290;
wire v_55291;
wire v_55292;
wire v_55293;
wire v_55294;
wire v_55295;
wire v_55296;
wire v_55297;
wire v_55298;
wire v_55299;
wire v_55300;
wire v_55301;
wire v_55302;
wire v_55303;
wire v_55304;
wire v_55305;
wire v_55306;
wire v_55307;
wire v_55308;
wire v_55309;
wire v_55310;
wire v_55311;
wire v_55312;
wire v_55313;
wire v_55314;
wire v_55315;
wire v_55316;
wire v_55317;
wire v_55318;
wire v_55319;
wire v_55320;
wire v_55321;
wire v_55322;
wire v_55323;
wire v_55324;
wire v_55325;
wire v_55326;
wire v_55327;
wire v_55328;
wire v_55329;
wire v_55330;
wire v_55331;
wire v_55332;
wire v_55333;
wire v_55334;
wire v_55335;
wire v_55336;
wire v_55337;
wire v_55338;
wire v_55339;
wire v_55340;
wire v_55341;
wire v_55342;
wire v_55343;
wire v_55344;
wire v_55345;
wire v_55346;
wire v_55347;
wire v_55348;
wire v_55349;
wire v_55350;
wire v_55351;
wire v_55352;
wire v_55353;
wire v_55354;
wire v_55355;
wire v_55356;
wire v_55357;
wire v_55358;
wire v_55359;
wire v_55360;
wire v_55361;
wire v_55362;
wire v_55363;
wire v_55364;
wire v_55365;
wire v_55366;
wire v_55367;
wire v_55368;
wire v_55369;
wire v_55370;
wire v_55371;
wire v_55372;
wire v_55373;
wire v_55374;
wire v_55375;
wire v_55376;
wire v_55377;
wire v_55378;
wire v_55379;
wire v_55380;
wire v_55381;
wire v_55382;
wire v_55383;
wire v_55384;
wire v_55385;
wire v_55386;
wire v_55387;
wire v_55388;
wire v_55389;
wire v_55390;
wire v_55391;
wire v_55392;
wire v_55393;
wire v_55394;
wire v_55395;
wire v_55396;
wire v_55397;
wire v_55398;
wire v_55399;
wire v_55400;
wire v_55401;
wire v_55402;
wire v_55403;
wire v_55404;
wire v_55405;
wire v_55406;
wire v_55407;
wire v_55408;
wire v_55409;
wire v_55410;
wire v_55411;
wire v_55412;
wire v_55413;
wire v_55414;
wire v_55415;
wire v_55416;
wire v_55417;
wire v_55418;
wire v_55419;
wire v_55420;
wire v_55421;
wire v_55422;
wire v_55423;
wire v_55424;
wire v_55425;
wire v_55426;
wire v_55427;
wire v_55428;
wire v_55429;
wire v_55430;
wire v_55431;
wire v_55432;
wire v_55433;
wire v_55434;
wire v_55435;
wire v_55436;
wire v_55437;
wire v_55438;
wire v_55439;
wire v_55440;
wire v_55441;
wire v_55442;
wire v_55443;
wire v_55444;
wire v_55445;
wire v_55446;
wire v_55447;
wire v_55448;
wire v_55449;
wire v_55451;
wire v_55452;
wire v_55453;
wire v_55454;
wire v_55455;
wire v_55456;
wire v_55457;
wire v_55458;
wire v_55459;
wire v_55460;
wire v_55461;
wire v_55462;
wire v_55463;
wire v_55464;
wire v_55465;
wire v_55466;
wire v_55467;
wire v_55468;
wire v_55469;
wire v_55470;
wire v_55471;
wire v_55472;
wire v_55473;
wire v_55474;
wire v_55475;
wire v_55476;
wire v_55477;
wire v_55478;
wire v_55479;
wire v_55480;
wire v_55481;
wire v_55482;
wire v_55483;
wire v_55484;
wire v_55485;
wire v_55486;
wire v_55487;
wire v_55488;
wire v_55489;
wire v_55490;
wire v_55491;
wire v_55492;
wire v_55493;
wire v_55494;
wire v_55495;
wire v_55496;
wire v_55497;
wire v_55498;
wire v_55499;
wire v_55500;
wire v_55501;
wire v_55502;
wire v_55503;
wire v_55504;
wire v_55505;
wire v_55506;
wire v_55507;
wire v_55508;
wire v_55509;
wire v_55510;
wire v_55511;
wire v_55512;
wire v_55513;
wire v_55514;
wire v_55515;
wire v_55516;
wire v_55517;
wire v_55518;
wire v_55519;
wire v_55520;
wire v_55521;
wire v_55522;
wire v_55523;
wire v_55524;
wire v_55525;
wire v_55526;
wire v_55527;
wire v_55528;
wire v_55529;
wire v_55530;
wire v_55531;
wire v_55532;
wire v_55533;
wire v_55534;
wire v_55535;
wire v_55536;
wire v_55537;
wire v_55538;
wire v_55539;
wire v_55540;
wire v_55541;
wire v_55542;
wire v_55543;
wire v_55544;
wire v_55545;
wire v_55546;
wire v_55547;
wire v_55548;
wire v_55549;
wire v_55550;
wire v_55551;
wire v_55552;
wire v_55553;
wire v_55554;
wire v_55555;
wire v_55556;
wire v_55557;
wire v_55558;
wire v_55559;
wire v_55560;
wire v_55561;
wire v_55562;
wire v_55563;
wire v_55564;
wire v_55565;
wire v_55566;
wire v_55567;
wire v_55568;
wire v_55569;
wire v_55570;
wire v_55571;
wire v_55572;
wire v_55573;
wire v_55574;
wire v_55575;
wire v_55576;
wire v_55577;
wire v_55578;
wire v_55579;
wire v_55580;
wire v_55581;
wire v_55582;
wire v_55583;
wire v_55584;
wire v_55585;
wire v_55586;
wire v_55587;
wire v_55588;
wire v_55589;
wire v_55590;
wire v_55591;
wire v_55592;
wire v_55593;
wire v_55594;
wire v_55595;
wire v_55596;
wire v_55597;
wire v_55598;
wire v_55599;
wire v_55600;
wire v_55601;
wire v_55602;
wire v_55603;
wire v_55604;
wire v_55605;
wire v_55606;
wire v_55607;
wire v_55608;
wire v_55609;
wire v_55610;
wire v_55611;
wire v_55612;
wire v_55613;
wire v_55614;
wire v_55615;
wire v_55616;
wire v_55617;
wire v_55618;
wire v_55619;
wire v_55620;
wire v_55621;
wire v_55622;
wire v_55623;
wire v_55624;
wire v_55625;
wire v_55626;
wire v_55627;
wire v_55628;
wire v_55629;
wire v_55630;
wire v_55631;
wire v_55632;
wire v_55633;
wire v_55634;
wire v_55635;
wire v_55636;
wire v_55637;
wire v_55638;
wire v_55639;
wire v_55640;
wire v_55641;
wire v_55642;
wire v_55643;
wire v_55644;
wire v_55645;
wire v_55646;
wire v_55647;
wire v_55648;
wire v_55649;
wire v_55650;
wire v_55651;
wire v_55652;
wire v_55653;
wire v_55654;
wire v_55655;
wire v_55656;
wire v_55657;
wire v_55658;
wire v_55659;
wire v_55660;
wire v_55661;
wire v_55662;
wire v_55663;
wire v_55664;
wire v_55665;
wire v_55666;
wire v_55667;
wire v_55668;
wire v_55669;
wire v_55670;
wire v_55671;
wire v_55672;
wire v_55673;
wire v_55674;
wire v_55675;
wire v_55676;
wire v_55677;
wire v_55678;
wire v_55679;
wire v_55680;
wire v_55681;
wire v_55682;
wire v_55683;
wire v_55684;
wire v_55685;
wire v_55686;
wire v_55687;
wire v_55688;
wire v_55689;
wire v_55690;
wire v_55691;
wire v_55692;
wire v_55694;
wire v_55695;
wire v_55696;
wire v_55697;
wire v_55698;
wire v_55699;
wire v_55700;
wire v_55701;
wire v_55702;
wire v_55703;
wire v_55704;
wire v_55705;
wire v_55706;
wire v_55707;
wire v_55708;
wire v_55709;
wire v_55710;
wire v_55711;
wire v_55712;
wire v_55713;
wire v_55714;
wire v_55715;
wire v_55716;
wire v_55717;
wire v_55718;
wire v_55719;
wire v_55720;
wire v_55721;
wire v_55722;
wire v_55723;
wire v_55724;
wire v_55725;
wire v_55726;
wire v_55727;
wire v_55728;
wire v_55729;
wire v_55730;
wire v_55731;
wire v_55732;
wire v_55733;
wire v_55734;
wire v_55735;
wire v_55736;
wire v_55737;
wire v_55738;
wire v_55739;
wire v_55740;
wire v_55741;
wire v_55742;
wire v_55743;
wire v_55744;
wire v_55745;
wire v_55746;
wire v_55747;
wire v_55748;
wire v_55749;
wire v_55750;
wire v_55751;
wire v_55752;
wire v_55753;
wire v_55754;
wire v_55755;
wire v_55756;
wire v_55757;
wire v_55758;
wire v_55759;
wire v_55760;
wire v_55761;
wire v_55762;
wire v_55763;
wire v_55764;
wire v_55765;
wire v_55766;
wire v_55767;
wire v_55768;
wire v_55769;
wire v_55770;
wire v_55771;
wire v_55772;
wire v_55773;
wire v_55774;
wire v_55775;
wire v_55776;
wire v_55777;
wire v_55778;
wire v_55779;
wire v_55780;
wire v_55781;
wire v_55782;
wire v_55783;
wire v_55784;
wire v_55785;
wire v_55786;
wire v_55787;
wire v_55788;
wire v_55789;
wire v_55790;
wire v_55791;
wire v_55792;
wire v_55793;
wire v_55794;
wire v_55795;
wire v_55796;
wire v_55797;
wire v_55798;
wire v_55799;
wire v_55800;
wire v_55801;
wire v_55802;
wire v_55803;
wire v_55804;
wire v_55805;
wire v_55806;
wire v_55807;
wire v_55808;
wire v_55809;
wire v_55810;
wire v_55811;
wire v_55812;
wire v_55813;
wire v_55814;
wire v_55815;
wire v_55816;
wire v_55817;
wire v_55818;
wire v_55819;
wire v_55820;
wire v_55821;
wire v_55822;
wire v_55823;
wire v_55824;
wire v_55825;
wire v_55826;
wire v_55827;
wire v_55828;
wire v_55829;
wire v_55830;
wire v_55831;
wire v_55832;
wire v_55833;
wire v_55834;
wire v_55835;
wire v_55836;
wire v_55837;
wire v_55838;
wire v_55839;
wire v_55840;
wire v_55841;
wire v_55842;
wire v_55843;
wire v_55844;
wire v_55845;
wire v_55846;
wire v_55847;
wire v_55848;
wire v_55849;
wire v_55850;
wire v_55851;
wire v_55852;
wire v_55853;
wire v_55854;
wire v_55855;
wire v_55856;
wire v_55857;
wire v_55858;
wire v_55859;
wire v_55860;
wire v_55861;
wire v_55862;
wire v_55863;
wire v_55864;
wire v_55865;
wire v_55866;
wire v_55867;
wire v_55868;
wire v_55869;
wire v_55870;
wire v_55871;
wire v_55872;
wire v_55873;
wire v_55874;
wire v_55875;
wire v_55876;
wire v_55877;
wire v_55878;
wire v_55879;
wire v_55880;
wire v_55881;
wire v_55882;
wire v_55883;
wire v_55884;
wire v_55885;
wire v_55886;
wire v_55887;
wire v_55888;
wire v_55889;
wire v_55890;
wire v_55891;
wire v_55892;
wire v_55893;
wire v_55894;
wire v_55895;
wire v_55896;
wire v_55897;
wire v_55898;
wire v_55899;
wire v_55900;
wire v_55901;
wire v_55902;
wire v_55903;
wire v_55904;
wire v_55905;
wire v_55906;
wire v_55907;
wire v_55908;
wire v_55909;
wire v_55910;
wire v_55911;
wire v_55912;
wire v_55913;
wire v_55914;
wire v_55915;
wire v_55916;
wire v_55917;
wire v_55918;
wire v_55919;
wire v_55920;
wire v_55921;
wire v_55922;
wire v_55923;
wire v_55924;
wire v_55925;
wire v_55926;
wire v_55927;
wire v_55928;
wire v_55929;
wire v_55930;
wire v_55931;
wire v_55932;
wire v_55933;
wire v_55934;
wire v_55935;
wire v_55937;
wire v_55938;
wire v_55939;
wire v_55940;
wire v_55941;
wire v_55942;
wire v_55943;
wire v_55944;
wire v_55945;
wire v_55946;
wire v_55947;
wire v_55948;
wire v_55949;
wire v_55950;
wire v_55951;
wire v_55952;
wire v_55953;
wire v_55954;
wire v_55955;
wire v_55956;
wire v_55957;
wire v_55958;
wire v_55959;
wire v_55960;
wire v_55961;
wire v_55962;
wire v_55963;
wire v_55964;
wire v_55965;
wire v_55966;
wire v_55967;
wire v_55968;
wire v_55969;
wire v_55970;
wire v_55971;
wire v_55972;
wire v_55973;
wire v_55974;
wire v_55975;
wire v_55976;
wire v_55977;
wire v_55978;
wire v_55979;
wire v_55980;
wire v_55981;
wire v_55982;
wire v_55983;
wire v_55984;
wire v_55985;
wire v_55986;
wire v_55987;
wire v_55988;
wire v_55989;
wire v_55990;
wire v_55991;
wire v_55992;
wire v_55993;
wire v_55994;
wire v_55995;
wire v_55996;
wire v_55997;
wire v_55998;
wire v_55999;
wire v_56000;
wire v_56001;
wire v_56002;
wire v_56003;
wire v_56004;
wire v_56005;
wire v_56006;
wire v_56007;
wire v_56008;
wire v_56009;
wire v_56010;
wire v_56011;
wire v_56012;
wire v_56013;
wire v_56014;
wire v_56015;
wire v_56016;
wire v_56017;
wire v_56018;
wire v_56019;
wire v_56020;
wire v_56021;
wire v_56022;
wire v_56023;
wire v_56024;
wire v_56025;
wire v_56026;
wire v_56027;
wire v_56028;
wire v_56029;
wire v_56030;
wire v_56031;
wire v_56032;
wire v_56033;
wire v_56034;
wire v_56035;
wire v_56036;
wire v_56037;
wire v_56038;
wire v_56039;
wire v_56040;
wire v_56041;
wire v_56042;
wire v_56043;
wire v_56044;
wire v_56045;
wire v_56046;
wire v_56047;
wire v_56048;
wire v_56049;
wire v_56050;
wire v_56051;
wire v_56052;
wire v_56053;
wire v_56054;
wire v_56055;
wire v_56056;
wire v_56057;
wire v_56058;
wire v_56059;
wire v_56060;
wire v_56061;
wire v_56062;
wire v_56063;
wire v_56064;
wire v_56065;
wire v_56066;
wire v_56067;
wire v_56068;
wire v_56069;
wire v_56070;
wire v_56071;
wire v_56072;
wire v_56073;
wire v_56074;
wire v_56075;
wire v_56076;
wire v_56077;
wire v_56078;
wire v_56079;
wire v_56080;
wire v_56081;
wire v_56082;
wire v_56083;
wire v_56084;
wire v_56085;
wire v_56086;
wire v_56087;
wire v_56088;
wire v_56089;
wire v_56090;
wire v_56091;
wire v_56092;
wire v_56093;
wire v_56094;
wire v_56095;
wire v_56096;
wire v_56097;
wire v_56098;
wire v_56099;
wire v_56100;
wire v_56101;
wire v_56102;
wire v_56103;
wire v_56104;
wire v_56105;
wire v_56106;
wire v_56107;
wire v_56108;
wire v_56109;
wire v_56110;
wire v_56111;
wire v_56112;
wire v_56113;
wire v_56114;
wire v_56115;
wire v_56116;
wire v_56117;
wire v_56118;
wire v_56119;
wire v_56120;
wire v_56121;
wire v_56122;
wire v_56123;
wire v_56124;
wire v_56125;
wire v_56126;
wire v_56127;
wire v_56128;
wire v_56129;
wire v_56130;
wire v_56131;
wire v_56132;
wire v_56133;
wire v_56134;
wire v_56135;
wire v_56136;
wire v_56137;
wire v_56138;
wire v_56139;
wire v_56140;
wire v_56141;
wire v_56142;
wire v_56143;
wire v_56144;
wire v_56145;
wire v_56146;
wire v_56147;
wire v_56148;
wire v_56149;
wire v_56150;
wire v_56151;
wire v_56152;
wire v_56153;
wire v_56154;
wire v_56155;
wire v_56156;
wire v_56157;
wire v_56158;
wire v_56159;
wire v_56160;
wire v_56161;
wire v_56162;
wire v_56163;
wire v_56164;
wire v_56165;
wire v_56166;
wire v_56167;
wire v_56168;
wire v_56169;
wire v_56170;
wire v_56171;
wire v_56172;
wire v_56173;
wire v_56174;
wire v_56175;
wire v_56176;
wire v_56177;
wire v_56178;
wire v_56180;
wire v_56181;
wire v_56182;
wire v_56183;
wire v_56184;
wire v_56185;
wire v_56186;
wire v_56187;
wire v_56188;
wire v_56189;
wire v_56190;
wire v_56191;
wire v_56192;
wire v_56193;
wire v_56194;
wire v_56195;
wire v_56196;
wire v_56197;
wire v_56198;
wire v_56199;
wire v_56200;
wire v_56201;
wire v_56202;
wire v_56203;
wire v_56204;
wire v_56205;
wire v_56206;
wire v_56207;
wire v_56208;
wire v_56209;
wire v_56210;
wire v_56211;
wire v_56212;
wire v_56213;
wire v_56214;
wire v_56215;
wire v_56216;
wire v_56217;
wire v_56218;
wire v_56219;
wire v_56220;
wire v_56221;
wire v_56222;
wire v_56223;
wire v_56224;
wire v_56225;
wire v_56226;
wire v_56227;
wire v_56228;
wire v_56229;
wire v_56230;
wire v_56231;
wire v_56232;
wire v_56233;
wire v_56234;
wire v_56235;
wire v_56236;
wire v_56237;
wire v_56238;
wire v_56239;
wire v_56240;
wire v_56241;
wire v_56242;
wire v_56243;
wire v_56244;
wire v_56245;
wire v_56246;
wire v_56247;
wire v_56248;
wire v_56249;
wire v_56250;
wire v_56251;
wire v_56252;
wire v_56253;
wire v_56254;
wire v_56255;
wire v_56256;
wire v_56257;
wire v_56258;
wire v_56259;
wire v_56260;
wire v_56261;
wire v_56262;
wire v_56263;
wire v_56264;
wire v_56265;
wire v_56266;
wire v_56267;
wire v_56268;
wire v_56269;
wire v_56270;
wire v_56271;
wire v_56272;
wire v_56273;
wire v_56274;
wire v_56275;
wire v_56276;
wire v_56277;
wire v_56278;
wire v_56279;
wire v_56280;
wire v_56281;
wire v_56282;
wire v_56283;
wire v_56284;
wire v_56285;
wire v_56286;
wire v_56287;
wire v_56288;
wire v_56289;
wire v_56290;
wire v_56291;
wire v_56292;
wire v_56293;
wire v_56294;
wire v_56295;
wire v_56296;
wire v_56297;
wire v_56298;
wire v_56299;
wire v_56300;
wire v_56301;
wire v_56302;
wire v_56303;
wire v_56304;
wire v_56305;
wire v_56306;
wire v_56307;
wire v_56308;
wire v_56309;
wire v_56310;
wire v_56311;
wire v_56312;
wire v_56313;
wire v_56314;
wire v_56315;
wire v_56316;
wire v_56317;
wire v_56318;
wire v_56319;
wire v_56320;
wire v_56321;
wire v_56322;
wire v_56323;
wire v_56324;
wire v_56325;
wire v_56326;
wire v_56327;
wire v_56328;
wire v_56329;
wire v_56330;
wire v_56331;
wire v_56332;
wire v_56333;
wire v_56334;
wire v_56335;
wire v_56336;
wire v_56337;
wire v_56338;
wire v_56339;
wire v_56340;
wire v_56341;
wire v_56342;
wire v_56343;
wire v_56344;
wire v_56345;
wire v_56346;
wire v_56347;
wire v_56348;
wire v_56349;
wire v_56350;
wire v_56351;
wire v_56352;
wire v_56353;
wire v_56354;
wire v_56355;
wire v_56356;
wire v_56357;
wire v_56358;
wire v_56359;
wire v_56360;
wire v_56361;
wire v_56362;
wire v_56363;
wire v_56364;
wire v_56365;
wire v_56366;
wire v_56367;
wire v_56368;
wire v_56369;
wire v_56370;
wire v_56371;
wire v_56372;
wire v_56373;
wire v_56374;
wire v_56375;
wire v_56376;
wire v_56377;
wire v_56378;
wire v_56379;
wire v_56380;
wire v_56381;
wire v_56382;
wire v_56383;
wire v_56384;
wire v_56385;
wire v_56386;
wire v_56387;
wire v_56388;
wire v_56389;
wire v_56390;
wire v_56391;
wire v_56392;
wire v_56393;
wire v_56394;
wire v_56395;
wire v_56396;
wire v_56397;
wire v_56398;
wire v_56399;
wire v_56400;
wire v_56401;
wire v_56402;
wire v_56403;
wire v_56404;
wire v_56405;
wire v_56406;
wire v_56407;
wire v_56408;
wire v_56409;
wire v_56410;
wire v_56411;
wire v_56412;
wire v_56413;
wire v_56414;
wire v_56415;
wire v_56416;
wire v_56417;
wire v_56418;
wire v_56419;
wire v_56420;
wire v_56421;
wire v_56423;
wire v_56424;
wire v_56425;
wire v_56426;
wire v_56427;
wire v_56428;
wire v_56429;
wire v_56430;
wire v_56431;
wire v_56432;
wire v_56433;
wire v_56434;
wire v_56435;
wire v_56436;
wire v_56437;
wire v_56438;
wire v_56439;
wire v_56440;
wire v_56441;
wire v_56442;
wire v_56443;
wire v_56444;
wire v_56445;
wire v_56446;
wire v_56447;
wire v_56448;
wire v_56449;
wire v_56450;
wire v_56451;
wire v_56452;
wire v_56453;
wire v_56454;
wire v_56455;
wire v_56456;
wire v_56457;
wire v_56458;
wire v_56459;
wire v_56460;
wire v_56461;
wire v_56462;
wire v_56463;
wire v_56464;
wire v_56465;
wire v_56466;
wire v_56467;
wire v_56468;
wire v_56469;
wire v_56470;
wire v_56471;
wire v_56472;
wire v_56473;
wire v_56474;
wire v_56475;
wire v_56476;
wire v_56477;
wire v_56478;
wire v_56479;
wire v_56480;
wire v_56481;
wire v_56482;
wire v_56483;
wire v_56484;
wire v_56485;
wire v_56486;
wire v_56487;
wire v_56488;
wire v_56489;
wire v_56490;
wire v_56491;
wire v_56492;
wire v_56493;
wire v_56494;
wire v_56495;
wire v_56496;
wire v_56497;
wire v_56498;
wire v_56499;
wire v_56500;
wire v_56501;
wire v_56502;
wire v_56503;
wire v_56504;
wire v_56505;
wire v_56506;
wire v_56507;
wire v_56508;
wire v_56509;
wire v_56510;
wire v_56511;
wire v_56512;
wire v_56513;
wire v_56514;
wire v_56515;
wire v_56516;
wire v_56517;
wire v_56518;
wire v_56519;
wire v_56520;
wire v_56521;
wire v_56522;
wire v_56523;
wire v_56524;
wire v_56525;
wire v_56526;
wire v_56527;
wire v_56528;
wire v_56529;
wire v_56530;
wire v_56531;
wire v_56532;
wire v_56533;
wire v_56534;
wire v_56535;
wire v_56536;
wire v_56537;
wire v_56538;
wire v_56539;
wire v_56540;
wire v_56541;
wire v_56542;
wire v_56543;
wire v_56544;
wire v_56545;
wire v_56546;
wire v_56547;
wire v_56548;
wire v_56549;
wire v_56550;
wire v_56551;
wire v_56552;
wire v_56553;
wire v_56554;
wire v_56555;
wire v_56556;
wire v_56557;
wire v_56558;
wire v_56559;
wire v_56560;
wire v_56561;
wire v_56562;
wire v_56563;
wire v_56564;
wire v_56565;
wire v_56566;
wire v_56567;
wire v_56568;
wire v_56569;
wire v_56570;
wire v_56571;
wire v_56572;
wire v_56573;
wire v_56574;
wire v_56575;
wire v_56576;
wire v_56577;
wire v_56578;
wire v_56579;
wire v_56580;
wire v_56581;
wire v_56582;
wire v_56583;
wire v_56584;
wire v_56585;
wire v_56586;
wire v_56587;
wire v_56588;
wire v_56589;
wire v_56590;
wire v_56591;
wire v_56592;
wire v_56593;
wire v_56594;
wire v_56595;
wire v_56596;
wire v_56597;
wire v_56598;
wire v_56599;
wire v_56600;
wire v_56601;
wire v_56602;
wire v_56603;
wire v_56604;
wire v_56605;
wire v_56606;
wire v_56607;
wire v_56608;
wire v_56609;
wire v_56610;
wire v_56611;
wire v_56612;
wire v_56613;
wire v_56614;
wire v_56615;
wire v_56616;
wire v_56617;
wire v_56618;
wire v_56619;
wire v_56620;
wire v_56621;
wire v_56622;
wire v_56623;
wire v_56624;
wire v_56625;
wire v_56626;
wire v_56627;
wire v_56628;
wire v_56629;
wire v_56630;
wire v_56631;
wire v_56632;
wire v_56633;
wire v_56634;
wire v_56635;
wire v_56636;
wire v_56637;
wire v_56638;
wire v_56639;
wire v_56640;
wire v_56641;
wire v_56642;
wire v_56643;
wire v_56644;
wire v_56645;
wire v_56646;
wire v_56647;
wire v_56648;
wire v_56649;
wire v_56650;
wire v_56651;
wire v_56652;
wire v_56653;
wire v_56654;
wire v_56655;
wire v_56656;
wire v_56657;
wire v_56658;
wire v_56659;
wire v_56660;
wire v_56661;
wire v_56662;
wire v_56663;
wire v_56664;
wire v_56666;
wire v_56667;
wire v_56668;
wire v_56669;
wire v_56670;
wire v_56671;
wire v_56672;
wire v_56673;
wire v_56674;
wire v_56675;
wire v_56676;
wire v_56677;
wire v_56678;
wire v_56679;
wire v_56680;
wire v_56681;
wire v_56682;
wire v_56683;
wire v_56684;
wire v_56685;
wire v_56686;
wire v_56687;
wire v_56688;
wire v_56689;
wire v_56690;
wire v_56691;
wire v_56692;
wire v_56693;
wire v_56694;
wire v_56695;
wire v_56696;
wire v_56697;
wire v_56698;
wire v_56699;
wire v_56700;
wire v_56701;
wire v_56702;
wire v_56703;
wire v_56704;
wire v_56705;
wire v_56706;
wire v_56707;
wire v_56708;
wire v_56709;
wire v_56710;
wire v_56711;
wire v_56712;
wire v_56713;
wire v_56714;
wire v_56715;
wire v_56716;
wire v_56717;
wire v_56718;
wire v_56719;
wire v_56720;
wire v_56721;
wire v_56722;
wire v_56723;
wire v_56724;
wire v_56725;
wire v_56726;
wire v_56727;
wire v_56728;
wire v_56729;
wire v_56730;
wire v_56731;
wire v_56732;
wire v_56733;
wire v_56734;
wire v_56735;
wire v_56736;
wire v_56737;
wire v_56738;
wire v_56739;
wire v_56740;
wire v_56741;
wire v_56742;
wire v_56743;
wire v_56744;
wire v_56745;
wire v_56746;
wire v_56747;
wire v_56748;
wire v_56749;
wire v_56750;
wire v_56751;
wire v_56752;
wire v_56753;
wire v_56754;
wire v_56755;
wire v_56756;
wire v_56757;
wire v_56758;
wire v_56759;
wire v_56760;
wire v_56761;
wire v_56762;
wire v_56763;
wire v_56764;
wire v_56765;
wire v_56766;
wire v_56767;
wire v_56768;
wire v_56769;
wire v_56770;
wire v_56771;
wire v_56772;
wire v_56773;
wire v_56774;
wire v_56775;
wire v_56776;
wire v_56777;
wire v_56778;
wire v_56779;
wire v_56780;
wire v_56781;
wire v_56782;
wire v_56783;
wire v_56784;
wire v_56785;
wire v_56786;
wire v_56787;
wire v_56788;
wire v_56789;
wire v_56790;
wire v_56791;
wire v_56792;
wire v_56793;
wire v_56794;
wire v_56795;
wire v_56796;
wire v_56797;
wire v_56798;
wire v_56799;
wire v_56800;
wire v_56801;
wire v_56802;
wire v_56803;
wire v_56804;
wire v_56805;
wire v_56806;
wire v_56807;
wire v_56808;
wire v_56809;
wire v_56810;
wire v_56811;
wire v_56812;
wire v_56813;
wire v_56814;
wire v_56815;
wire v_56816;
wire v_56817;
wire v_56818;
wire v_56819;
wire v_56820;
wire v_56821;
wire v_56822;
wire v_56823;
wire v_56824;
wire v_56825;
wire v_56826;
wire v_56827;
wire v_56828;
wire v_56829;
wire v_56830;
wire v_56831;
wire v_56832;
wire v_56833;
wire v_56834;
wire v_56835;
wire v_56836;
wire v_56837;
wire v_56838;
wire v_56839;
wire v_56840;
wire v_56841;
wire v_56842;
wire v_56843;
wire v_56844;
wire v_56845;
wire v_56846;
wire v_56847;
wire v_56848;
wire v_56849;
wire v_56850;
wire v_56851;
wire v_56852;
wire v_56853;
wire v_56854;
wire v_56855;
wire v_56856;
wire v_56857;
wire v_56858;
wire v_56859;
wire v_56860;
wire v_56861;
wire v_56862;
wire v_56863;
wire v_56864;
wire v_56865;
wire v_56866;
wire v_56867;
wire v_56868;
wire v_56869;
wire v_56870;
wire v_56871;
wire v_56872;
wire v_56873;
wire v_56874;
wire v_56875;
wire v_56876;
wire v_56877;
wire v_56878;
wire v_56879;
wire v_56880;
wire v_56881;
wire v_56882;
wire v_56883;
wire v_56884;
wire v_56885;
wire v_56886;
wire v_56887;
wire v_56888;
wire v_56889;
wire v_56890;
wire v_56891;
wire v_56892;
wire v_56893;
wire v_56894;
wire v_56895;
wire v_56896;
wire v_56897;
wire v_56898;
wire v_56899;
wire v_56900;
wire v_56901;
wire v_56902;
wire v_56903;
wire v_56904;
wire v_56905;
wire v_56906;
wire v_56907;
wire v_56909;
wire v_56910;
wire v_56911;
wire v_56912;
wire v_56913;
wire v_56914;
wire v_56915;
wire v_56916;
wire v_56917;
wire v_56918;
wire v_56919;
wire v_56920;
wire v_56921;
wire v_56922;
wire v_56923;
wire v_56924;
wire v_56925;
wire v_56926;
wire v_56927;
wire v_56928;
wire v_56929;
wire v_56930;
wire v_56931;
wire v_56932;
wire v_56933;
wire v_56934;
wire v_56935;
wire v_56936;
wire v_56937;
wire v_56938;
wire v_56939;
wire v_56940;
wire v_56941;
wire v_56942;
wire v_56943;
wire v_56944;
wire v_56945;
wire v_56946;
wire v_56947;
wire v_56948;
wire v_56949;
wire v_56950;
wire v_56951;
wire v_56952;
wire v_56953;
wire v_56954;
wire v_56955;
wire v_56956;
wire v_56957;
wire v_56958;
wire v_56959;
wire v_56960;
wire v_56961;
wire v_56962;
wire v_56963;
wire v_56964;
wire v_56965;
wire v_56966;
wire v_56967;
wire v_56968;
wire v_56969;
wire v_56970;
wire v_56971;
wire v_56972;
wire v_56973;
wire v_56974;
wire v_56975;
wire v_56976;
wire v_56977;
wire v_56978;
wire v_56979;
wire v_56980;
wire v_56981;
wire v_56982;
wire v_56983;
wire v_56984;
wire v_56985;
wire v_56986;
wire v_56987;
wire v_56988;
wire v_56989;
wire v_56990;
wire v_56991;
wire v_56992;
wire v_56993;
wire v_56994;
wire v_56995;
wire v_56996;
wire v_56997;
wire v_56998;
wire v_56999;
wire v_57000;
wire v_57001;
wire v_57002;
wire v_57003;
wire v_57004;
wire v_57005;
wire v_57006;
wire v_57007;
wire v_57008;
wire v_57009;
wire v_57010;
wire v_57011;
wire v_57012;
wire v_57013;
wire v_57014;
wire v_57015;
wire v_57016;
wire v_57017;
wire v_57018;
wire v_57019;
wire v_57020;
wire v_57021;
wire v_57022;
wire v_57023;
wire v_57024;
wire v_57025;
wire v_57026;
wire v_57027;
wire v_57028;
wire v_57029;
wire v_57030;
wire v_57031;
wire v_57032;
wire v_57033;
wire v_57034;
wire v_57035;
wire v_57036;
wire v_57037;
wire v_57038;
wire v_57039;
wire v_57040;
wire v_57041;
wire v_57042;
wire v_57043;
wire v_57044;
wire v_57045;
wire v_57046;
wire v_57047;
wire v_57048;
wire v_57049;
wire v_57050;
wire v_57051;
wire v_57052;
wire v_57053;
wire v_57054;
wire v_57055;
wire v_57056;
wire v_57057;
wire v_57058;
wire v_57059;
wire v_57060;
wire v_57061;
wire v_57062;
wire v_57063;
wire v_57064;
wire v_57065;
wire v_57066;
wire v_57067;
wire v_57068;
wire v_57069;
wire v_57070;
wire v_57071;
wire v_57072;
wire v_57073;
wire v_57074;
wire v_57075;
wire v_57076;
wire v_57077;
wire v_57078;
wire v_57079;
wire v_57080;
wire v_57081;
wire v_57082;
wire v_57083;
wire v_57084;
wire v_57085;
wire v_57086;
wire v_57087;
wire v_57088;
wire v_57089;
wire v_57090;
wire v_57091;
wire v_57092;
wire v_57093;
wire v_57094;
wire v_57095;
wire v_57096;
wire v_57097;
wire v_57098;
wire v_57099;
wire v_57100;
wire v_57101;
wire v_57102;
wire v_57103;
wire v_57104;
wire v_57105;
wire v_57106;
wire v_57107;
wire v_57108;
wire v_57109;
wire v_57110;
wire v_57111;
wire v_57112;
wire v_57113;
wire v_57114;
wire v_57115;
wire v_57116;
wire v_57117;
wire v_57118;
wire v_57119;
wire v_57120;
wire v_57121;
wire v_57122;
wire v_57123;
wire v_57124;
wire v_57125;
wire v_57126;
wire v_57127;
wire v_57128;
wire v_57129;
wire v_57130;
wire v_57131;
wire v_57132;
wire v_57133;
wire v_57134;
wire v_57135;
wire v_57136;
wire v_57137;
wire v_57138;
wire v_57139;
wire v_57140;
wire v_57141;
wire v_57142;
wire v_57143;
wire v_57144;
wire v_57145;
wire v_57146;
wire v_57147;
wire v_57148;
wire v_57149;
wire v_57150;
wire v_57152;
wire v_57153;
wire v_57154;
wire v_57155;
wire v_57156;
wire v_57157;
wire v_57158;
wire v_57159;
wire v_57160;
wire v_57161;
wire v_57162;
wire v_57163;
wire v_57164;
wire v_57165;
wire v_57166;
wire v_57167;
wire v_57168;
wire v_57169;
wire v_57170;
wire v_57171;
wire v_57172;
wire v_57173;
wire v_57174;
wire v_57175;
wire v_57176;
wire v_57177;
wire v_57178;
wire v_57179;
wire v_57180;
wire v_57181;
wire v_57182;
wire v_57183;
wire v_57184;
wire v_57185;
wire v_57186;
wire v_57187;
wire v_57188;
wire v_57189;
wire v_57190;
wire v_57191;
wire v_57192;
wire v_57193;
wire v_57194;
wire v_57195;
wire v_57196;
wire v_57197;
wire v_57198;
wire v_57199;
wire v_57200;
wire v_57201;
wire v_57202;
wire v_57203;
wire v_57204;
wire v_57205;
wire v_57206;
wire v_57207;
wire v_57208;
wire v_57209;
wire v_57210;
wire v_57211;
wire v_57212;
wire v_57213;
wire v_57214;
wire v_57215;
wire v_57216;
wire v_57217;
wire v_57218;
wire v_57219;
wire v_57220;
wire v_57221;
wire v_57222;
wire v_57223;
wire v_57224;
wire v_57225;
wire v_57226;
wire v_57227;
wire v_57228;
wire v_57229;
wire v_57230;
wire v_57231;
wire v_57232;
wire v_57233;
wire v_57234;
wire v_57235;
wire v_57236;
wire v_57237;
wire v_57238;
wire v_57239;
wire v_57240;
wire v_57241;
wire v_57242;
wire v_57243;
wire v_57244;
wire v_57245;
wire v_57246;
wire v_57247;
wire v_57248;
wire v_57249;
wire v_57250;
wire v_57251;
wire v_57252;
wire v_57253;
wire v_57254;
wire v_57255;
wire v_57256;
wire v_57257;
wire v_57258;
wire v_57259;
wire v_57260;
wire v_57261;
wire v_57262;
wire v_57263;
wire v_57264;
wire v_57265;
wire v_57266;
wire v_57267;
wire v_57268;
wire v_57269;
wire v_57270;
wire v_57271;
wire v_57272;
wire v_57273;
wire v_57274;
wire v_57275;
wire v_57276;
wire v_57277;
wire v_57278;
wire v_57279;
wire v_57280;
wire v_57281;
wire v_57282;
wire v_57283;
wire v_57284;
wire v_57285;
wire v_57286;
wire v_57287;
wire v_57288;
wire v_57289;
wire v_57290;
wire v_57291;
wire v_57292;
wire v_57293;
wire v_57294;
wire v_57295;
wire v_57296;
wire v_57297;
wire v_57298;
wire v_57299;
wire v_57300;
wire v_57301;
wire v_57302;
wire v_57303;
wire v_57304;
wire v_57305;
wire v_57306;
wire v_57307;
wire v_57308;
wire v_57309;
wire v_57310;
wire v_57311;
wire v_57312;
wire v_57313;
wire v_57314;
wire v_57315;
wire v_57316;
wire v_57317;
wire v_57318;
wire v_57319;
wire v_57320;
wire v_57321;
wire v_57322;
wire v_57323;
wire v_57324;
wire v_57325;
wire v_57326;
wire v_57327;
wire v_57328;
wire v_57329;
wire v_57330;
wire v_57331;
wire v_57332;
wire v_57333;
wire v_57334;
wire v_57335;
wire v_57336;
wire v_57337;
wire v_57338;
wire v_57339;
wire v_57340;
wire v_57341;
wire v_57342;
wire v_57343;
wire v_57344;
wire v_57345;
wire v_57346;
wire v_57347;
wire v_57348;
wire v_57349;
wire v_57350;
wire v_57351;
wire v_57352;
wire v_57353;
wire v_57354;
wire v_57355;
wire v_57356;
wire v_57357;
wire v_57358;
wire v_57359;
wire v_57360;
wire v_57361;
wire v_57362;
wire v_57363;
wire v_57364;
wire v_57365;
wire v_57366;
wire v_57367;
wire v_57368;
wire v_57369;
wire v_57370;
wire v_57371;
wire v_57372;
wire v_57373;
wire v_57374;
wire v_57375;
wire v_57376;
wire v_57377;
wire v_57378;
wire v_57379;
wire v_57380;
wire v_57381;
wire v_57382;
wire v_57383;
wire v_57384;
wire v_57385;
wire v_57386;
wire v_57387;
wire v_57388;
wire v_57389;
wire v_57390;
wire v_57391;
wire v_57392;
wire v_57393;
wire v_57395;
wire v_57396;
wire v_57397;
wire v_57398;
wire v_57399;
wire v_57400;
wire v_57401;
wire v_57402;
wire v_57403;
wire v_57404;
wire v_57405;
wire v_57406;
wire v_57407;
wire v_57408;
wire v_57409;
wire v_57410;
wire v_57411;
wire v_57412;
wire v_57413;
wire v_57414;
wire v_57415;
wire v_57416;
wire v_57417;
wire v_57418;
wire v_57419;
wire v_57420;
wire v_57421;
wire v_57422;
wire v_57423;
wire v_57424;
wire v_57425;
wire v_57426;
wire v_57427;
wire v_57428;
wire v_57429;
wire v_57430;
wire v_57431;
wire v_57432;
wire v_57433;
wire v_57434;
wire v_57435;
wire v_57436;
wire v_57437;
wire v_57438;
wire v_57439;
wire v_57440;
wire v_57441;
wire v_57442;
wire v_57443;
wire v_57444;
wire v_57445;
wire v_57446;
wire v_57447;
wire v_57448;
wire v_57449;
wire v_57450;
wire v_57451;
wire v_57452;
wire v_57453;
wire v_57454;
wire v_57455;
wire v_57456;
wire v_57457;
wire v_57458;
wire v_57459;
wire v_57460;
wire v_57461;
wire v_57462;
wire v_57463;
wire v_57464;
wire v_57465;
wire v_57466;
wire v_57467;
wire v_57468;
wire v_57469;
wire v_57470;
wire v_57471;
wire v_57472;
wire v_57473;
wire v_57474;
wire v_57475;
wire v_57476;
wire v_57477;
wire v_57478;
wire v_57479;
wire v_57480;
wire v_57481;
wire v_57482;
wire v_57483;
wire v_57484;
wire v_57485;
wire v_57486;
wire v_57487;
wire v_57488;
wire v_57489;
wire v_57490;
wire v_57491;
wire v_57492;
wire v_57493;
wire v_57494;
wire v_57495;
wire v_57496;
wire v_57497;
wire v_57498;
wire v_57499;
wire v_57500;
wire v_57501;
wire v_57502;
wire v_57503;
wire v_57504;
wire v_57505;
wire v_57506;
wire v_57507;
wire v_57508;
wire v_57509;
wire v_57510;
wire v_57511;
wire v_57512;
wire v_57513;
wire v_57514;
wire v_57515;
wire v_57516;
wire v_57517;
wire v_57518;
wire v_57519;
wire v_57520;
wire v_57521;
wire v_57522;
wire v_57523;
wire v_57524;
wire v_57525;
wire v_57526;
wire v_57527;
wire v_57528;
wire v_57529;
wire v_57530;
wire v_57531;
wire v_57532;
wire v_57533;
wire v_57534;
wire v_57535;
wire v_57536;
wire v_57537;
wire v_57538;
wire v_57539;
wire v_57540;
wire v_57541;
wire v_57542;
wire v_57543;
wire v_57544;
wire v_57545;
wire v_57546;
wire v_57547;
wire v_57548;
wire v_57549;
wire v_57550;
wire v_57551;
wire v_57552;
wire v_57553;
wire v_57554;
wire v_57555;
wire v_57556;
wire v_57557;
wire v_57558;
wire v_57559;
wire v_57560;
wire v_57561;
wire v_57562;
wire v_57563;
wire v_57564;
wire v_57565;
wire v_57566;
wire v_57567;
wire v_57568;
wire v_57569;
wire v_57570;
wire v_57571;
wire v_57572;
wire v_57573;
wire v_57574;
wire v_57575;
wire v_57576;
wire v_57577;
wire v_57578;
wire v_57579;
wire v_57580;
wire v_57581;
wire v_57582;
wire v_57583;
wire v_57584;
wire v_57585;
wire v_57586;
wire v_57587;
wire v_57588;
wire v_57589;
wire v_57590;
wire v_57591;
wire v_57592;
wire v_57593;
wire v_57594;
wire v_57595;
wire v_57596;
wire v_57597;
wire v_57598;
wire v_57599;
wire v_57600;
wire v_57601;
wire v_57602;
wire v_57603;
wire v_57604;
wire v_57605;
wire v_57606;
wire v_57607;
wire v_57608;
wire v_57609;
wire v_57610;
wire v_57611;
wire v_57612;
wire v_57613;
wire v_57614;
wire v_57615;
wire v_57616;
wire v_57617;
wire v_57618;
wire v_57619;
wire v_57620;
wire v_57621;
wire v_57622;
wire v_57623;
wire v_57624;
wire v_57625;
wire v_57626;
wire v_57627;
wire v_57628;
wire v_57629;
wire v_57630;
wire v_57631;
wire v_57632;
wire v_57633;
wire v_57634;
wire v_57635;
wire v_57636;
wire v_57638;
wire v_57639;
wire v_57640;
wire v_57641;
wire v_57642;
wire v_57643;
wire v_57644;
wire v_57645;
wire v_57646;
wire v_57647;
wire v_57648;
wire v_57649;
wire v_57650;
wire v_57651;
wire v_57652;
wire v_57653;
wire v_57654;
wire v_57655;
wire v_57656;
wire v_57657;
wire v_57658;
wire v_57659;
wire v_57660;
wire v_57661;
wire v_57662;
wire v_57663;
wire v_57664;
wire v_57665;
wire v_57666;
wire v_57667;
wire v_57668;
wire v_57669;
wire v_57670;
wire v_57671;
wire v_57672;
wire v_57673;
wire v_57674;
wire v_57675;
wire v_57676;
wire v_57677;
wire v_57678;
wire v_57679;
wire v_57680;
wire v_57681;
wire v_57682;
wire v_57683;
wire v_57684;
wire v_57685;
wire v_57686;
wire v_57687;
wire v_57688;
wire v_57689;
wire v_57690;
wire v_57691;
wire v_57692;
wire v_57693;
wire v_57694;
wire v_57695;
wire v_57696;
wire v_57697;
wire v_57698;
wire v_57699;
wire v_57700;
wire v_57701;
wire v_57702;
wire v_57703;
wire v_57704;
wire v_57705;
wire v_57706;
wire v_57707;
wire v_57708;
wire v_57709;
wire v_57710;
wire v_57711;
wire v_57712;
wire v_57713;
wire v_57714;
wire v_57715;
wire v_57716;
wire v_57717;
wire v_57718;
wire v_57719;
wire v_57720;
wire v_57721;
wire v_57722;
wire v_57723;
wire v_57724;
wire v_57725;
wire v_57726;
wire v_57727;
wire v_57728;
wire v_57729;
wire v_57730;
wire v_57731;
wire v_57732;
wire v_57733;
wire v_57734;
wire v_57735;
wire v_57736;
wire v_57737;
wire v_57738;
wire v_57739;
wire v_57740;
wire v_57741;
wire v_57742;
wire v_57743;
wire v_57744;
wire v_57745;
wire v_57746;
wire v_57747;
wire v_57748;
wire v_57749;
wire v_57750;
wire v_57751;
wire v_57752;
wire v_57753;
wire v_57754;
wire v_57755;
wire v_57756;
wire v_57757;
wire v_57758;
wire v_57759;
wire v_57760;
wire v_57761;
wire v_57762;
wire v_57763;
wire v_57764;
wire v_57765;
wire v_57766;
wire v_57767;
wire v_57768;
wire v_57769;
wire v_57770;
wire v_57771;
wire v_57772;
wire v_57773;
wire v_57774;
wire v_57775;
wire v_57776;
wire v_57777;
wire v_57778;
wire v_57779;
wire v_57780;
wire v_57781;
wire v_57782;
wire v_57783;
wire v_57784;
wire v_57785;
wire v_57786;
wire v_57787;
wire v_57788;
wire v_57789;
wire v_57790;
wire v_57791;
wire v_57792;
wire v_57793;
wire v_57794;
wire v_57795;
wire v_57796;
wire v_57797;
wire v_57798;
wire v_57799;
wire v_57800;
wire v_57801;
wire v_57802;
wire v_57803;
wire v_57804;
wire v_57805;
wire v_57806;
wire v_57807;
wire v_57808;
wire v_57809;
wire v_57810;
wire v_57811;
wire v_57812;
wire v_57813;
wire v_57814;
wire v_57815;
wire v_57816;
wire v_57817;
wire v_57818;
wire v_57819;
wire v_57820;
wire v_57821;
wire v_57822;
wire v_57823;
wire v_57824;
wire v_57825;
wire v_57826;
wire v_57827;
wire v_57828;
wire v_57829;
wire v_57830;
wire v_57831;
wire v_57832;
wire v_57833;
wire v_57834;
wire v_57835;
wire v_57836;
wire v_57837;
wire v_57838;
wire v_57839;
wire v_57840;
wire v_57841;
wire v_57842;
wire v_57843;
wire v_57844;
wire v_57845;
wire v_57846;
wire v_57847;
wire v_57848;
wire v_57849;
wire v_57850;
wire v_57851;
wire v_57852;
wire v_57853;
wire v_57854;
wire v_57855;
wire v_57856;
wire v_57857;
wire v_57858;
wire v_57859;
wire v_57860;
wire v_57861;
wire v_57862;
wire v_57863;
wire v_57864;
wire v_57865;
wire v_57866;
wire v_57867;
wire v_57868;
wire v_57869;
wire v_57870;
wire v_57871;
wire v_57872;
wire v_57873;
wire v_57874;
wire v_57875;
wire v_57876;
wire v_57877;
wire v_57878;
wire v_57879;
wire v_57881;
wire v_57882;
wire v_57883;
wire v_57884;
wire v_57885;
wire v_57886;
wire v_57887;
wire v_57888;
wire v_57889;
wire v_57890;
wire v_57891;
wire v_57892;
wire v_57893;
wire v_57894;
wire v_57895;
wire v_57896;
wire v_57897;
wire v_57898;
wire v_57899;
wire v_57900;
wire v_57901;
wire v_57902;
wire v_57903;
wire v_57904;
wire v_57905;
wire v_57906;
wire v_57907;
wire v_57908;
wire v_57909;
wire v_57910;
wire v_57911;
wire v_57912;
wire v_57913;
wire v_57914;
wire v_57915;
wire v_57916;
wire v_57917;
wire v_57918;
wire v_57919;
wire v_57920;
wire v_57921;
wire v_57922;
wire v_57923;
wire v_57924;
wire v_57925;
wire v_57926;
wire v_57927;
wire v_57928;
wire v_57929;
wire v_57930;
wire v_57931;
wire v_57932;
wire v_57933;
wire v_57934;
wire v_57935;
wire v_57936;
wire v_57937;
wire v_57938;
wire v_57939;
wire v_57940;
wire v_57941;
wire v_57942;
wire v_57943;
wire v_57944;
wire v_57945;
wire v_57946;
wire v_57947;
wire v_57948;
wire v_57949;
wire v_57950;
wire v_57951;
wire v_57952;
wire v_57953;
wire v_57954;
wire v_57955;
wire v_57956;
wire v_57957;
wire v_57958;
wire v_57959;
wire v_57960;
wire v_57961;
wire v_57962;
wire v_57963;
wire v_57964;
wire v_57965;
wire v_57966;
wire v_57967;
wire v_57968;
wire v_57969;
wire v_57970;
wire v_57971;
wire v_57972;
wire v_57973;
wire v_57974;
wire v_57975;
wire v_57976;
wire v_57977;
wire v_57978;
wire v_57979;
wire v_57980;
wire v_57981;
wire v_57982;
wire v_57983;
wire v_57984;
wire v_57985;
wire v_57986;
wire v_57987;
wire v_57988;
wire v_57989;
wire v_57990;
wire v_57991;
wire v_57992;
wire v_57993;
wire v_57994;
wire v_57995;
wire v_57996;
wire v_57997;
wire v_57998;
wire v_57999;
wire v_58000;
wire v_58001;
wire v_58002;
wire v_58003;
wire v_58004;
wire v_58005;
wire v_58006;
wire v_58007;
wire v_58008;
wire v_58009;
wire v_58010;
wire v_58011;
wire v_58012;
wire v_58013;
wire v_58014;
wire v_58015;
wire v_58016;
wire v_58017;
wire v_58018;
wire v_58019;
wire v_58020;
wire v_58021;
wire v_58022;
wire v_58023;
wire v_58024;
wire v_58025;
wire v_58026;
wire v_58027;
wire v_58028;
wire v_58029;
wire v_58030;
wire v_58031;
wire v_58032;
wire v_58033;
wire v_58034;
wire v_58035;
wire v_58036;
wire v_58037;
wire v_58038;
wire v_58039;
wire v_58040;
wire v_58041;
wire v_58042;
wire v_58043;
wire v_58044;
wire v_58045;
wire v_58046;
wire v_58047;
wire v_58048;
wire v_58049;
wire v_58050;
wire v_58051;
wire v_58052;
wire v_58053;
wire v_58054;
wire v_58055;
wire v_58056;
wire v_58057;
wire v_58058;
wire v_58059;
wire v_58060;
wire v_58061;
wire v_58062;
wire v_58063;
wire v_58064;
wire v_58065;
wire v_58066;
wire v_58067;
wire v_58068;
wire v_58069;
wire v_58070;
wire v_58071;
wire v_58072;
wire v_58073;
wire v_58074;
wire v_58075;
wire v_58076;
wire v_58077;
wire v_58078;
wire v_58079;
wire v_58080;
wire v_58081;
wire v_58082;
wire v_58083;
wire v_58084;
wire v_58085;
wire v_58086;
wire v_58087;
wire v_58088;
wire v_58089;
wire v_58090;
wire v_58091;
wire v_58092;
wire v_58093;
wire v_58094;
wire v_58095;
wire v_58096;
wire v_58097;
wire v_58098;
wire v_58099;
wire v_58100;
wire v_58101;
wire v_58102;
wire v_58103;
wire v_58104;
wire v_58105;
wire v_58106;
wire v_58107;
wire v_58108;
wire v_58109;
wire v_58110;
wire v_58111;
wire v_58112;
wire v_58113;
wire v_58114;
wire v_58115;
wire v_58116;
wire v_58117;
wire v_58118;
wire v_58119;
wire v_58120;
wire v_58121;
wire v_58122;
wire v_58123;
wire v_58124;
wire v_58125;
wire v_58126;
wire v_58127;
wire v_58128;
wire v_58129;
wire v_58130;
wire v_58131;
wire v_58132;
wire v_58133;
wire v_58134;
wire v_58135;
wire v_58136;
wire v_58137;
wire v_58138;
wire v_58139;
wire v_58140;
wire v_58141;
wire v_58142;
wire v_58143;
wire v_58144;
wire v_58145;
wire v_58146;
wire v_58147;
wire v_58148;
wire v_58149;
wire v_58150;
wire v_58151;
wire v_58152;
wire v_58153;
wire v_58154;
wire v_58155;
wire v_58156;
wire v_58157;
wire v_58158;
wire v_58159;
wire v_58160;
wire v_58161;
wire v_58162;
wire v_58163;
wire v_58164;
wire v_58165;
wire v_58166;
wire v_58167;
wire v_58168;
wire v_58169;
wire v_58170;
wire v_58171;
wire v_58172;
wire v_58173;
wire v_58174;
wire v_58175;
wire v_58176;
wire v_58177;
wire v_58178;
wire v_58179;
wire v_58180;
wire v_58181;
wire v_58182;
wire v_58183;
wire v_58184;
wire v_58185;
wire v_58186;
wire v_58187;
wire v_58188;
wire v_58189;
wire v_58190;
wire v_58191;
wire v_58192;
wire v_58193;
wire v_58194;
wire v_58195;
wire v_58196;
wire v_58197;
wire v_58198;
wire v_58199;
wire v_58200;
wire v_58201;
wire v_58202;
wire v_58203;
wire v_58204;
wire v_58205;
wire v_58206;
wire v_58207;
wire v_58208;
wire v_58209;
wire v_58210;
wire v_58211;
wire v_58212;
wire v_58213;
wire v_58214;
wire v_58215;
wire v_58216;
wire v_58217;
wire v_58218;
wire v_58219;
wire v_58220;
wire v_58221;
wire v_58222;
wire v_58223;
wire v_58224;
wire v_58225;
wire v_58226;
wire v_58227;
wire v_58228;
wire v_58229;
wire v_58230;
wire v_58231;
wire v_58232;
wire v_58233;
wire v_58234;
wire v_58235;
wire v_58236;
wire v_58237;
wire v_58238;
wire v_58239;
wire v_58240;
wire v_58241;
wire v_58242;
wire v_58243;
wire v_58244;
wire v_58245;
wire v_58246;
wire v_58247;
wire v_58248;
wire v_58249;
wire v_58250;
wire v_58251;
wire v_58252;
wire v_58253;
wire v_58254;
wire v_58255;
wire v_58256;
wire v_58257;
wire v_58258;
wire v_58259;
wire v_58260;
wire v_58261;
wire v_58262;
wire v_58263;
wire v_58264;
wire v_58265;
wire v_58266;
wire v_58267;
wire v_58268;
wire v_58269;
wire v_58270;
wire v_58271;
wire v_58273;
wire v_58274;
wire v_58275;
wire v_58276;
wire v_58277;
wire v_58278;
wire v_58279;
wire v_58280;
wire v_58281;
wire v_58282;
wire v_58283;
wire v_58284;
wire v_58285;
wire v_58286;
wire v_58287;
wire v_58288;
wire v_58289;
wire v_58290;
wire v_58291;
wire v_58292;
wire v_58293;
wire v_58294;
wire v_58295;
wire v_58296;
wire v_58297;
wire v_58298;
wire v_58299;
wire v_58300;
wire v_58301;
wire v_58302;
wire v_58303;
wire v_58304;
wire v_58305;
wire v_58306;
wire v_58307;
wire v_58308;
wire v_58309;
wire v_58310;
wire v_58311;
wire v_58312;
wire v_58313;
wire v_58314;
wire v_58315;
wire v_58316;
wire v_58317;
wire v_58318;
wire v_58319;
wire v_58320;
wire v_58321;
wire v_58322;
wire v_58323;
wire v_58324;
wire v_58325;
wire v_58326;
wire v_58327;
wire v_58328;
wire v_58329;
wire v_58330;
wire v_58331;
wire v_58332;
wire v_58333;
wire v_58334;
wire v_58335;
wire v_58336;
wire v_58337;
wire v_58338;
wire v_58339;
wire v_58340;
wire v_58341;
wire v_58342;
wire v_58343;
wire v_58344;
wire v_58345;
wire v_58346;
wire v_58347;
wire v_58348;
wire v_58349;
wire v_58350;
wire v_58351;
wire v_58352;
wire v_58353;
wire v_58354;
wire v_58355;
wire v_58356;
wire v_58357;
wire v_58358;
wire v_58359;
wire v_58360;
wire v_58361;
wire v_58362;
wire v_58363;
wire v_58364;
wire v_58365;
wire v_58367;
wire v_58369;
wire v_58370;
wire v_58371;
wire v_58373;
wire v_58374;
wire v_58375;
wire v_58377;
wire v_58378;
wire v_58379;
wire v_58381;
wire v_58382;
wire v_58384;
wire v_58385;
wire v_58386;
wire v_58388;
wire v_58389;
wire v_58390;
wire v_58392;
wire v_58393;
wire v_58394;
wire v_58396;
wire v_58397;
wire v_58398;
wire v_58400;
wire v_58401;
wire v_58402;
wire v_58404;
wire v_58405;
wire v_58406;
wire v_58408;
wire v_58409;
wire v_58410;
wire v_58412;
wire v_58413;
wire v_58414;
wire v_58416;
wire v_58417;
wire v_58418;
wire v_58420;
wire v_58421;
wire v_58422;
wire v_58424;
wire v_58425;
wire v_58426;
wire v_58428;
wire v_58429;
wire v_58430;
wire v_58432;
wire v_58433;
wire v_58434;
wire v_58435;
wire v_58436;
wire v_58437;
wire v_58438;
wire v_58439;
wire v_58440;
wire v_58441;
wire v_58442;
wire v_58443;
wire v_58444;
wire v_58445;
wire v_58446;
wire v_58447;
wire v_58448;
wire v_58449;
wire v_58450;
wire v_58451;
wire v_58452;
wire v_58453;
wire v_58454;
wire v_58455;
wire v_58456;
wire v_58457;
wire v_58458;
wire v_58459;
wire v_58460;
wire v_58461;
wire v_58462;
wire v_58463;
wire v_58464;
wire v_58465;
wire v_58466;
wire v_58467;
wire v_58468;
wire v_58469;
wire v_58470;
wire v_58471;
wire v_58472;
wire v_58473;
wire v_58474;
wire v_58475;
wire v_58476;
wire v_58477;
wire v_58478;
wire v_58479;
wire v_58480;
wire v_58481;
wire v_58482;
wire v_58483;
wire v_58484;
wire v_58485;
wire v_58486;
wire v_58487;
wire v_58488;
wire v_58489;
wire v_58490;
wire v_58491;
wire v_58492;
wire v_58493;
wire v_58494;
wire v_58495;
wire v_58496;
wire v_58497;
wire v_58498;
wire v_58499;
wire v_58500;
wire v_58501;
wire v_58502;
wire v_58503;
wire v_58504;
wire v_58505;
wire v_58506;
wire v_58507;
wire v_58508;
wire v_58509;
wire v_58510;
wire v_58511;
wire v_58512;
wire v_58513;
wire v_58514;
wire v_58515;
wire v_58516;
wire v_58517;
wire v_58518;
wire v_58519;
wire v_58520;
wire v_58521;
wire v_58522;
wire v_58523;
wire v_58524;
wire v_58525;
wire v_58526;
wire v_58527;
wire v_58528;
wire v_58529;
wire v_58530;
wire v_58531;
wire v_58532;
wire v_58533;
wire v_58534;
wire v_58535;
wire v_58536;
wire v_58537;
wire v_58538;
wire v_58539;
wire v_58540;
wire v_58541;
wire v_58542;
wire v_58543;
wire v_58544;
wire v_58545;
wire v_58546;
wire v_58547;
wire v_58548;
wire v_58549;
wire v_58550;
wire v_58551;
wire v_58552;
wire v_58553;
wire v_58554;
wire v_58555;
wire v_58556;
wire v_58557;
wire v_58558;
wire v_58559;
wire v_58560;
wire v_58561;
wire v_58562;
wire v_58563;
wire v_58564;
wire v_58565;
wire v_58566;
wire v_58567;
wire v_58568;
wire v_58569;
wire v_58570;
wire v_58571;
wire v_58572;
wire v_58573;
wire v_58574;
wire v_58575;
wire v_58576;
wire v_58577;
wire v_58578;
wire v_58579;
wire v_58580;
wire v_58581;
wire v_58582;
wire v_58583;
wire v_58584;
wire v_58585;
wire v_58586;
wire v_58587;
wire v_58588;
wire v_58589;
wire v_58590;
wire v_58591;
wire v_58592;
wire v_58593;
wire v_58594;
wire v_58595;
wire v_58596;
wire v_58597;
wire v_58598;
wire v_58599;
wire v_58600;
wire v_58601;
wire v_58602;
wire v_58603;
wire v_58604;
wire v_58605;
wire v_58606;
wire v_58607;
wire v_58608;
wire v_58609;
wire v_58610;
wire v_58611;
wire v_58612;
wire v_58613;
wire v_58614;
wire v_58615;
wire v_58616;
wire v_58617;
wire v_58618;
wire v_58619;
wire v_58620;
wire v_58621;
wire v_58622;
wire v_58623;
wire v_58624;
wire v_58625;
wire v_58627;
wire v_58628;
wire v_58629;
wire v_58630;
wire v_58631;
wire v_58632;
wire v_58633;
wire v_58634;
wire v_58635;
wire v_58636;
wire v_58637;
wire v_58638;
wire v_58639;
wire v_58640;
wire v_58641;
wire v_58642;
wire v_58643;
wire v_58644;
wire v_58645;
wire v_58646;
wire v_58647;
wire v_58648;
wire v_58649;
wire v_58650;
wire v_58651;
wire v_58652;
wire v_58653;
wire v_58654;
wire v_58655;
wire v_58656;
wire v_58657;
wire v_58658;
wire v_58659;
wire v_58660;
wire v_58661;
wire v_58662;
wire v_58663;
wire v_58664;
wire v_58665;
wire v_58666;
wire v_58667;
wire v_58668;
wire v_58669;
wire v_58670;
wire v_58671;
wire v_58672;
wire v_58673;
wire v_58674;
wire v_58675;
wire v_58676;
wire v_58677;
wire v_58678;
wire v_58679;
wire v_58680;
wire v_58681;
wire v_58682;
wire v_58683;
wire v_58684;
wire v_58685;
wire v_58686;
wire v_58687;
wire v_58688;
wire v_58689;
wire v_58690;
wire v_58691;
wire v_58692;
wire v_58693;
wire v_58694;
wire v_58695;
wire v_58696;
wire v_58697;
wire v_58698;
wire v_58699;
wire v_58700;
wire v_58701;
wire v_58702;
wire v_58703;
wire v_58704;
wire v_58705;
wire v_58706;
wire v_58707;
wire v_58708;
wire v_58709;
wire v_58710;
wire v_58711;
wire v_58712;
wire v_58713;
wire v_58714;
wire v_58715;
wire v_58716;
wire v_58717;
wire v_58718;
wire v_58719;
wire v_58720;
wire v_58721;
wire v_58722;
wire v_58723;
wire v_58724;
wire v_58725;
wire v_58726;
wire v_58727;
wire v_58728;
wire v_58729;
wire v_58730;
wire v_58731;
wire v_58732;
wire v_58733;
wire v_58734;
wire v_58735;
wire v_58736;
wire v_58737;
wire v_58738;
wire v_58739;
wire v_58740;
wire v_58741;
wire v_58742;
wire v_58743;
wire v_58744;
wire v_58745;
wire v_58746;
wire v_58747;
wire v_58748;
wire v_58749;
wire v_58750;
wire v_58751;
wire v_58752;
wire v_58753;
wire v_58754;
wire v_58755;
wire v_58756;
wire v_58757;
wire v_58758;
wire v_58759;
wire v_58760;
wire v_58761;
wire v_58762;
wire v_58763;
wire v_58764;
wire v_58765;
wire v_58766;
wire v_58767;
wire v_58768;
wire v_58769;
wire v_58770;
wire v_58771;
wire v_58772;
wire v_58773;
wire v_58774;
wire v_58775;
wire v_58776;
wire v_58777;
wire v_58778;
wire v_58779;
wire v_58780;
wire v_58781;
wire v_58782;
wire v_58783;
wire v_58784;
wire v_58785;
wire v_58786;
wire v_58787;
wire v_58788;
wire v_58789;
wire v_58790;
wire v_58791;
wire v_58792;
wire v_58793;
wire v_58794;
wire v_58795;
wire v_58796;
wire v_58797;
wire v_58798;
wire v_58799;
wire v_58800;
wire v_58801;
wire v_58802;
wire v_58803;
wire v_58804;
wire v_58805;
wire v_58806;
wire v_58807;
wire v_58808;
wire v_58809;
wire v_58810;
wire v_58811;
wire v_58812;
wire v_58813;
wire v_58814;
wire v_58815;
wire v_58816;
wire v_58817;
wire v_58818;
wire v_58819;
wire v_58820;
wire v_58821;
wire v_58822;
wire v_58823;
wire v_58824;
wire v_58825;
wire v_58826;
wire v_58827;
wire v_58828;
wire v_58829;
wire v_58830;
wire v_58831;
wire v_58832;
wire v_58833;
wire v_58834;
wire v_58835;
wire v_58836;
wire v_58837;
wire v_58838;
wire v_58839;
wire v_58840;
wire v_58841;
wire v_58842;
wire v_58843;
wire v_58844;
wire v_58845;
wire v_58846;
wire v_58847;
wire v_58848;
wire v_58849;
wire v_58850;
wire v_58851;
wire v_58852;
wire v_58853;
wire v_58854;
wire v_58855;
wire v_58856;
wire v_58857;
wire v_58858;
wire v_58859;
wire v_58860;
wire v_58861;
wire v_58862;
wire v_58863;
wire v_58864;
wire v_58865;
wire v_58866;
wire v_58867;
wire v_58868;
wire v_58870;
wire v_58871;
wire v_58872;
wire v_58873;
wire v_58874;
wire v_58875;
wire v_58876;
wire v_58877;
wire v_58878;
wire v_58879;
wire v_58880;
wire v_58881;
wire v_58882;
wire v_58883;
wire v_58884;
wire v_58885;
wire v_58886;
wire v_58887;
wire v_58888;
wire v_58889;
wire v_58890;
wire v_58891;
wire v_58892;
wire v_58893;
wire v_58894;
wire v_58895;
wire v_58896;
wire v_58897;
wire v_58898;
wire v_58899;
wire v_58900;
wire v_58901;
wire v_58902;
wire v_58903;
wire v_58904;
wire v_58905;
wire v_58906;
wire v_58907;
wire v_58908;
wire v_58909;
wire v_58910;
wire v_58911;
wire v_58912;
wire v_58913;
wire v_58914;
wire v_58915;
wire v_58916;
wire v_58917;
wire v_58918;
wire v_58919;
wire v_58920;
wire v_58921;
wire v_58922;
wire v_58923;
wire v_58924;
wire v_58925;
wire v_58926;
wire v_58927;
wire v_58928;
wire v_58929;
wire v_58930;
wire v_58931;
wire v_58932;
wire v_58933;
wire v_58934;
wire v_58935;
wire v_58936;
wire v_58937;
wire v_58938;
wire v_58939;
wire v_58940;
wire v_58941;
wire v_58942;
wire v_58943;
wire v_58944;
wire v_58945;
wire v_58946;
wire v_58947;
wire v_58948;
wire v_58949;
wire v_58950;
wire v_58951;
wire v_58952;
wire v_58953;
wire v_58954;
wire v_58955;
wire v_58956;
wire v_58957;
wire v_58958;
wire v_58959;
wire v_58960;
wire v_58961;
wire v_58962;
wire v_58963;
wire v_58964;
wire v_58965;
wire v_58966;
wire v_58967;
wire v_58968;
wire v_58969;
wire v_58970;
wire v_58971;
wire v_58972;
wire v_58973;
wire v_58974;
wire v_58975;
wire v_58976;
wire v_58977;
wire v_58978;
wire v_58979;
wire v_58980;
wire v_58981;
wire v_58982;
wire v_58983;
wire v_58984;
wire v_58985;
wire v_58986;
wire v_58987;
wire v_58988;
wire v_58989;
wire v_58990;
wire v_58991;
wire v_58992;
wire v_58993;
wire v_58994;
wire v_58995;
wire v_58996;
wire v_58997;
wire v_58998;
wire v_58999;
wire v_59000;
wire v_59001;
wire v_59002;
wire v_59003;
wire v_59004;
wire v_59005;
wire v_59006;
wire v_59007;
wire v_59008;
wire v_59009;
wire v_59010;
wire v_59011;
wire v_59012;
wire v_59013;
wire v_59014;
wire v_59015;
wire v_59016;
wire v_59017;
wire v_59018;
wire v_59019;
wire v_59020;
wire v_59021;
wire v_59022;
wire v_59023;
wire v_59024;
wire v_59025;
wire v_59026;
wire v_59027;
wire v_59028;
wire v_59029;
wire v_59030;
wire v_59031;
wire v_59032;
wire v_59033;
wire v_59034;
wire v_59035;
wire v_59036;
wire v_59037;
wire v_59038;
wire v_59039;
wire v_59040;
wire v_59041;
wire v_59042;
wire v_59043;
wire v_59044;
wire v_59045;
wire v_59046;
wire v_59047;
wire v_59048;
wire v_59049;
wire v_59050;
wire v_59051;
wire v_59052;
wire v_59053;
wire v_59054;
wire v_59055;
wire v_59056;
wire v_59057;
wire v_59058;
wire v_59059;
wire v_59060;
wire v_59061;
wire v_59062;
wire v_59063;
wire v_59064;
wire v_59065;
wire v_59066;
wire v_59067;
wire v_59068;
wire v_59069;
wire v_59070;
wire v_59071;
wire v_59072;
wire v_59073;
wire v_59074;
wire v_59075;
wire v_59076;
wire v_59077;
wire v_59078;
wire v_59079;
wire v_59080;
wire v_59081;
wire v_59082;
wire v_59083;
wire v_59084;
wire v_59085;
wire v_59086;
wire v_59087;
wire v_59088;
wire v_59089;
wire v_59090;
wire v_59091;
wire v_59092;
wire v_59093;
wire v_59094;
wire v_59095;
wire v_59096;
wire v_59097;
wire v_59098;
wire v_59099;
wire v_59100;
wire v_59101;
wire v_59102;
wire v_59103;
wire v_59104;
wire v_59105;
wire v_59106;
wire v_59107;
wire v_59108;
wire v_59109;
wire v_59110;
wire v_59111;
wire v_59113;
wire v_59114;
wire v_59115;
wire v_59116;
wire v_59117;
wire v_59118;
wire v_59119;
wire v_59120;
wire v_59121;
wire v_59122;
wire v_59123;
wire v_59124;
wire v_59125;
wire v_59126;
wire v_59127;
wire v_59128;
wire v_59129;
wire v_59130;
wire v_59131;
wire v_59132;
wire v_59133;
wire v_59134;
wire v_59135;
wire v_59136;
wire v_59137;
wire v_59138;
wire v_59139;
wire v_59140;
wire v_59141;
wire v_59142;
wire v_59143;
wire v_59144;
wire v_59145;
wire v_59146;
wire v_59147;
wire v_59148;
wire v_59149;
wire v_59150;
wire v_59151;
wire v_59152;
wire v_59153;
wire v_59154;
wire v_59155;
wire v_59156;
wire v_59157;
wire v_59158;
wire v_59159;
wire v_59160;
wire v_59161;
wire v_59162;
wire v_59163;
wire v_59164;
wire v_59165;
wire v_59166;
wire v_59167;
wire v_59168;
wire v_59169;
wire v_59170;
wire v_59171;
wire v_59172;
wire v_59173;
wire v_59174;
wire v_59175;
wire v_59176;
wire v_59177;
wire v_59178;
wire v_59179;
wire v_59180;
wire v_59181;
wire v_59182;
wire v_59183;
wire v_59184;
wire v_59185;
wire v_59186;
wire v_59187;
wire v_59188;
wire v_59189;
wire v_59190;
wire v_59191;
wire v_59192;
wire v_59193;
wire v_59194;
wire v_59195;
wire v_59196;
wire v_59197;
wire v_59198;
wire v_59199;
wire v_59200;
wire v_59201;
wire v_59202;
wire v_59203;
wire v_59204;
wire v_59205;
wire v_59206;
wire v_59207;
wire v_59208;
wire v_59209;
wire v_59210;
wire v_59211;
wire v_59212;
wire v_59213;
wire v_59214;
wire v_59215;
wire v_59216;
wire v_59217;
wire v_59218;
wire v_59219;
wire v_59220;
wire v_59221;
wire v_59222;
wire v_59223;
wire v_59224;
wire v_59225;
wire v_59226;
wire v_59227;
wire v_59228;
wire v_59229;
wire v_59230;
wire v_59231;
wire v_59232;
wire v_59233;
wire v_59234;
wire v_59235;
wire v_59236;
wire v_59237;
wire v_59238;
wire v_59239;
wire v_59240;
wire v_59241;
wire v_59242;
wire v_59243;
wire v_59244;
wire v_59245;
wire v_59246;
wire v_59247;
wire v_59248;
wire v_59249;
wire v_59250;
wire v_59251;
wire v_59252;
wire v_59253;
wire v_59254;
wire v_59255;
wire v_59256;
wire v_59257;
wire v_59258;
wire v_59259;
wire v_59260;
wire v_59261;
wire v_59262;
wire v_59263;
wire v_59264;
wire v_59265;
wire v_59266;
wire v_59267;
wire v_59268;
wire v_59269;
wire v_59270;
wire v_59271;
wire v_59272;
wire v_59273;
wire v_59274;
wire v_59275;
wire v_59276;
wire v_59277;
wire v_59278;
wire v_59279;
wire v_59280;
wire v_59281;
wire v_59282;
wire v_59283;
wire v_59284;
wire v_59285;
wire v_59286;
wire v_59287;
wire v_59288;
wire v_59289;
wire v_59290;
wire v_59291;
wire v_59292;
wire v_59293;
wire v_59294;
wire v_59295;
wire v_59296;
wire v_59297;
wire v_59298;
wire v_59299;
wire v_59300;
wire v_59301;
wire v_59302;
wire v_59303;
wire v_59304;
wire v_59305;
wire v_59306;
wire v_59307;
wire v_59308;
wire v_59309;
wire v_59310;
wire v_59311;
wire v_59312;
wire v_59313;
wire v_59314;
wire v_59315;
wire v_59316;
wire v_59317;
wire v_59318;
wire v_59319;
wire v_59320;
wire v_59321;
wire v_59322;
wire v_59323;
wire v_59324;
wire v_59325;
wire v_59326;
wire v_59327;
wire v_59328;
wire v_59329;
wire v_59330;
wire v_59331;
wire v_59332;
wire v_59333;
wire v_59334;
wire v_59335;
wire v_59336;
wire v_59337;
wire v_59338;
wire v_59339;
wire v_59340;
wire v_59341;
wire v_59342;
wire v_59343;
wire v_59344;
wire v_59345;
wire v_59346;
wire v_59347;
wire v_59348;
wire v_59349;
wire v_59350;
wire v_59351;
wire v_59352;
wire v_59353;
wire v_59354;
wire v_59356;
wire v_59357;
wire v_59358;
wire v_59359;
wire v_59360;
wire v_59361;
wire v_59362;
wire v_59363;
wire v_59364;
wire v_59365;
wire v_59366;
wire v_59367;
wire v_59368;
wire v_59369;
wire v_59370;
wire v_59371;
wire v_59372;
wire v_59373;
wire v_59374;
wire v_59375;
wire v_59376;
wire v_59377;
wire v_59378;
wire v_59379;
wire v_59380;
wire v_59381;
wire v_59382;
wire v_59383;
wire v_59384;
wire v_59385;
wire v_59386;
wire v_59387;
wire v_59388;
wire v_59389;
wire v_59390;
wire v_59391;
wire v_59392;
wire v_59393;
wire v_59394;
wire v_59395;
wire v_59396;
wire v_59397;
wire v_59398;
wire v_59399;
wire v_59400;
wire v_59401;
wire v_59402;
wire v_59403;
wire v_59404;
wire v_59405;
wire v_59406;
wire v_59407;
wire v_59408;
wire v_59409;
wire v_59410;
wire v_59411;
wire v_59412;
wire v_59413;
wire v_59414;
wire v_59415;
wire v_59416;
wire v_59417;
wire v_59418;
wire v_59419;
wire v_59420;
wire v_59421;
wire v_59422;
wire v_59423;
wire v_59424;
wire v_59425;
wire v_59426;
wire v_59427;
wire v_59428;
wire v_59429;
wire v_59430;
wire v_59431;
wire v_59432;
wire v_59433;
wire v_59434;
wire v_59435;
wire v_59436;
wire v_59437;
wire v_59438;
wire v_59439;
wire v_59440;
wire v_59441;
wire v_59442;
wire v_59443;
wire v_59444;
wire v_59445;
wire v_59446;
wire v_59447;
wire v_59448;
wire v_59449;
wire v_59450;
wire v_59451;
wire v_59452;
wire v_59453;
wire v_59454;
wire v_59455;
wire v_59456;
wire v_59457;
wire v_59458;
wire v_59459;
wire v_59460;
wire v_59461;
wire v_59462;
wire v_59463;
wire v_59464;
wire v_59465;
wire v_59466;
wire v_59467;
wire v_59468;
wire v_59469;
wire v_59470;
wire v_59471;
wire v_59472;
wire v_59473;
wire v_59474;
wire v_59475;
wire v_59476;
wire v_59477;
wire v_59478;
wire v_59479;
wire v_59480;
wire v_59481;
wire v_59482;
wire v_59483;
wire v_59484;
wire v_59485;
wire v_59486;
wire v_59487;
wire v_59488;
wire v_59489;
wire v_59490;
wire v_59491;
wire v_59492;
wire v_59493;
wire v_59494;
wire v_59495;
wire v_59496;
wire v_59497;
wire v_59498;
wire v_59499;
wire v_59500;
wire v_59501;
wire v_59502;
wire v_59503;
wire v_59504;
wire v_59505;
wire v_59506;
wire v_59507;
wire v_59508;
wire v_59509;
wire v_59510;
wire v_59511;
wire v_59512;
wire v_59513;
wire v_59514;
wire v_59515;
wire v_59516;
wire v_59517;
wire v_59518;
wire v_59519;
wire v_59520;
wire v_59521;
wire v_59522;
wire v_59523;
wire v_59524;
wire v_59525;
wire v_59526;
wire v_59527;
wire v_59528;
wire v_59529;
wire v_59530;
wire v_59531;
wire v_59532;
wire v_59533;
wire v_59534;
wire v_59535;
wire v_59536;
wire v_59537;
wire v_59538;
wire v_59539;
wire v_59540;
wire v_59541;
wire v_59542;
wire v_59543;
wire v_59544;
wire v_59545;
wire v_59546;
wire v_59547;
wire v_59548;
wire v_59549;
wire v_59550;
wire v_59551;
wire v_59552;
wire v_59553;
wire v_59554;
wire v_59555;
wire v_59556;
wire v_59557;
wire v_59558;
wire v_59559;
wire v_59560;
wire v_59561;
wire v_59562;
wire v_59563;
wire v_59564;
wire v_59565;
wire v_59566;
wire v_59567;
wire v_59568;
wire v_59569;
wire v_59570;
wire v_59571;
wire v_59572;
wire v_59573;
wire v_59574;
wire v_59575;
wire v_59576;
wire v_59577;
wire v_59578;
wire v_59579;
wire v_59580;
wire v_59581;
wire v_59582;
wire v_59583;
wire v_59584;
wire v_59585;
wire v_59586;
wire v_59587;
wire v_59588;
wire v_59589;
wire v_59590;
wire v_59591;
wire v_59592;
wire v_59593;
wire v_59594;
wire v_59595;
wire v_59596;
wire v_59597;
wire v_59599;
wire v_59600;
wire v_59601;
wire v_59602;
wire v_59603;
wire v_59604;
wire v_59605;
wire v_59606;
wire v_59607;
wire v_59608;
wire v_59609;
wire v_59610;
wire v_59611;
wire v_59612;
wire v_59613;
wire v_59614;
wire v_59615;
wire v_59616;
wire v_59617;
wire v_59618;
wire v_59619;
wire v_59620;
wire v_59621;
wire v_59622;
wire v_59623;
wire v_59624;
wire v_59625;
wire v_59626;
wire v_59627;
wire v_59628;
wire v_59629;
wire v_59630;
wire v_59631;
wire v_59632;
wire v_59633;
wire v_59634;
wire v_59635;
wire v_59636;
wire v_59637;
wire v_59638;
wire v_59639;
wire v_59640;
wire v_59641;
wire v_59642;
wire v_59643;
wire v_59644;
wire v_59645;
wire v_59646;
wire v_59647;
wire v_59648;
wire v_59649;
wire v_59650;
wire v_59651;
wire v_59652;
wire v_59653;
wire v_59654;
wire v_59655;
wire v_59656;
wire v_59657;
wire v_59658;
wire v_59659;
wire v_59660;
wire v_59661;
wire v_59662;
wire v_59663;
wire v_59664;
wire v_59665;
wire v_59666;
wire v_59667;
wire v_59668;
wire v_59669;
wire v_59670;
wire v_59671;
wire v_59672;
wire v_59673;
wire v_59674;
wire v_59675;
wire v_59676;
wire v_59677;
wire v_59678;
wire v_59679;
wire v_59680;
wire v_59681;
wire v_59682;
wire v_59683;
wire v_59684;
wire v_59685;
wire v_59686;
wire v_59687;
wire v_59688;
wire v_59689;
wire v_59690;
wire v_59691;
wire v_59692;
wire v_59693;
wire v_59694;
wire v_59695;
wire v_59696;
wire v_59697;
wire v_59698;
wire v_59699;
wire v_59700;
wire v_59701;
wire v_59702;
wire v_59703;
wire v_59704;
wire v_59705;
wire v_59706;
wire v_59707;
wire v_59708;
wire v_59709;
wire v_59710;
wire v_59711;
wire v_59712;
wire v_59713;
wire v_59714;
wire v_59715;
wire v_59716;
wire v_59717;
wire v_59718;
wire v_59719;
wire v_59720;
wire v_59721;
wire v_59722;
wire v_59723;
wire v_59724;
wire v_59725;
wire v_59726;
wire v_59727;
wire v_59728;
wire v_59729;
wire v_59730;
wire v_59731;
wire v_59732;
wire v_59733;
wire v_59734;
wire v_59735;
wire v_59736;
wire v_59737;
wire v_59738;
wire v_59739;
wire v_59740;
wire v_59741;
wire v_59742;
wire v_59743;
wire v_59744;
wire v_59745;
wire v_59746;
wire v_59747;
wire v_59748;
wire v_59749;
wire v_59750;
wire v_59751;
wire v_59752;
wire v_59753;
wire v_59754;
wire v_59755;
wire v_59756;
wire v_59757;
wire v_59758;
wire v_59759;
wire v_59760;
wire v_59761;
wire v_59762;
wire v_59763;
wire v_59764;
wire v_59765;
wire v_59766;
wire v_59767;
wire v_59768;
wire v_59769;
wire v_59770;
wire v_59771;
wire v_59772;
wire v_59773;
wire v_59774;
wire v_59775;
wire v_59776;
wire v_59777;
wire v_59778;
wire v_59779;
wire v_59780;
wire v_59781;
wire v_59782;
wire v_59783;
wire v_59784;
wire v_59785;
wire v_59786;
wire v_59787;
wire v_59788;
wire v_59789;
wire v_59790;
wire v_59791;
wire v_59792;
wire v_59793;
wire v_59794;
wire v_59795;
wire v_59796;
wire v_59797;
wire v_59798;
wire v_59799;
wire v_59800;
wire v_59801;
wire v_59802;
wire v_59803;
wire v_59804;
wire v_59805;
wire v_59806;
wire v_59807;
wire v_59808;
wire v_59809;
wire v_59810;
wire v_59811;
wire v_59812;
wire v_59813;
wire v_59814;
wire v_59815;
wire v_59816;
wire v_59817;
wire v_59818;
wire v_59819;
wire v_59820;
wire v_59821;
wire v_59822;
wire v_59823;
wire v_59824;
wire v_59825;
wire v_59826;
wire v_59827;
wire v_59828;
wire v_59829;
wire v_59830;
wire v_59831;
wire v_59832;
wire v_59833;
wire v_59834;
wire v_59835;
wire v_59836;
wire v_59837;
wire v_59838;
wire v_59839;
wire v_59840;
wire v_59842;
wire v_59843;
wire v_59844;
wire v_59845;
wire v_59846;
wire v_59847;
wire v_59848;
wire v_59849;
wire v_59850;
wire v_59851;
wire v_59852;
wire v_59853;
wire v_59854;
wire v_59855;
wire v_59856;
wire v_59857;
wire v_59858;
wire v_59859;
wire v_59860;
wire v_59861;
wire v_59862;
wire v_59863;
wire v_59864;
wire v_59865;
wire v_59866;
wire v_59867;
wire v_59868;
wire v_59869;
wire v_59870;
wire v_59871;
wire v_59872;
wire v_59873;
wire v_59874;
wire v_59875;
wire v_59876;
wire v_59877;
wire v_59878;
wire v_59879;
wire v_59880;
wire v_59881;
wire v_59882;
wire v_59883;
wire v_59884;
wire v_59885;
wire v_59886;
wire v_59887;
wire v_59888;
wire v_59889;
wire v_59890;
wire v_59891;
wire v_59892;
wire v_59893;
wire v_59894;
wire v_59895;
wire v_59896;
wire v_59897;
wire v_59898;
wire v_59899;
wire v_59900;
wire v_59901;
wire v_59902;
wire v_59903;
wire v_59904;
wire v_59905;
wire v_59906;
wire v_59907;
wire v_59908;
wire v_59909;
wire v_59910;
wire v_59911;
wire v_59912;
wire v_59913;
wire v_59914;
wire v_59915;
wire v_59916;
wire v_59917;
wire v_59918;
wire v_59919;
wire v_59920;
wire v_59921;
wire v_59922;
wire v_59923;
wire v_59924;
wire v_59925;
wire v_59926;
wire v_59927;
wire v_59928;
wire v_59929;
wire v_59930;
wire v_59931;
wire v_59932;
wire v_59933;
wire v_59934;
wire v_59935;
wire v_59936;
wire v_59937;
wire v_59938;
wire v_59939;
wire v_59940;
wire v_59941;
wire v_59942;
wire v_59943;
wire v_59944;
wire v_59945;
wire v_59946;
wire v_59947;
wire v_59948;
wire v_59949;
wire v_59950;
wire v_59951;
wire v_59952;
wire v_59953;
wire v_59954;
wire v_59955;
wire v_59956;
wire v_59957;
wire v_59958;
wire v_59959;
wire v_59960;
wire v_59961;
wire v_59962;
wire v_59963;
wire v_59964;
wire v_59965;
wire v_59966;
wire v_59967;
wire v_59968;
wire v_59969;
wire v_59970;
wire v_59971;
wire v_59972;
wire v_59973;
wire v_59974;
wire v_59975;
wire v_59976;
wire v_59977;
wire v_59978;
wire v_59979;
wire v_59980;
wire v_59981;
wire v_59982;
wire v_59983;
wire v_59984;
wire v_59985;
wire v_59986;
wire v_59987;
wire v_59988;
wire v_59989;
wire v_59990;
wire v_59991;
wire v_59992;
wire v_59993;
wire v_59994;
wire v_59995;
wire v_59996;
wire v_59997;
wire v_59998;
wire v_59999;
wire v_60000;
wire v_60001;
wire v_60002;
wire v_60003;
wire v_60004;
wire v_60005;
wire v_60006;
wire v_60007;
wire v_60008;
wire v_60009;
wire v_60010;
wire v_60011;
wire v_60012;
wire v_60013;
wire v_60014;
wire v_60015;
wire v_60016;
wire v_60017;
wire v_60018;
wire v_60019;
wire v_60020;
wire v_60021;
wire v_60022;
wire v_60023;
wire v_60024;
wire v_60025;
wire v_60026;
wire v_60027;
wire v_60028;
wire v_60029;
wire v_60030;
wire v_60031;
wire v_60032;
wire v_60033;
wire v_60034;
wire v_60035;
wire v_60036;
wire v_60037;
wire v_60038;
wire v_60039;
wire v_60040;
wire v_60041;
wire v_60042;
wire v_60043;
wire v_60044;
wire v_60045;
wire v_60046;
wire v_60047;
wire v_60048;
wire v_60049;
wire v_60050;
wire v_60051;
wire v_60052;
wire v_60053;
wire v_60054;
wire v_60055;
wire v_60056;
wire v_60057;
wire v_60058;
wire v_60059;
wire v_60060;
wire v_60061;
wire v_60062;
wire v_60063;
wire v_60064;
wire v_60065;
wire v_60066;
wire v_60067;
wire v_60068;
wire v_60069;
wire v_60070;
wire v_60071;
wire v_60072;
wire v_60073;
wire v_60074;
wire v_60075;
wire v_60076;
wire v_60077;
wire v_60078;
wire v_60079;
wire v_60080;
wire v_60081;
wire v_60082;
wire v_60083;
wire v_60085;
wire v_60086;
wire v_60087;
wire v_60088;
wire v_60089;
wire v_60090;
wire v_60091;
wire v_60092;
wire v_60093;
wire v_60094;
wire v_60095;
wire v_60096;
wire v_60097;
wire v_60098;
wire v_60099;
wire v_60100;
wire v_60101;
wire v_60102;
wire v_60103;
wire v_60104;
wire v_60105;
wire v_60106;
wire v_60107;
wire v_60108;
wire v_60109;
wire v_60110;
wire v_60111;
wire v_60112;
wire v_60113;
wire v_60114;
wire v_60115;
wire v_60116;
wire v_60117;
wire v_60118;
wire v_60119;
wire v_60120;
wire v_60121;
wire v_60122;
wire v_60123;
wire v_60124;
wire v_60125;
wire v_60126;
wire v_60127;
wire v_60128;
wire v_60129;
wire v_60130;
wire v_60131;
wire v_60132;
wire v_60133;
wire v_60134;
wire v_60135;
wire v_60136;
wire v_60137;
wire v_60138;
wire v_60139;
wire v_60140;
wire v_60141;
wire v_60142;
wire v_60143;
wire v_60144;
wire v_60145;
wire v_60146;
wire v_60147;
wire v_60148;
wire v_60149;
wire v_60150;
wire v_60151;
wire v_60152;
wire v_60153;
wire v_60154;
wire v_60155;
wire v_60156;
wire v_60157;
wire v_60158;
wire v_60159;
wire v_60160;
wire v_60161;
wire v_60162;
wire v_60163;
wire v_60164;
wire v_60165;
wire v_60166;
wire v_60167;
wire v_60168;
wire v_60169;
wire v_60170;
wire v_60171;
wire v_60172;
wire v_60173;
wire v_60174;
wire v_60175;
wire v_60176;
wire v_60177;
wire v_60178;
wire v_60179;
wire v_60180;
wire v_60181;
wire v_60182;
wire v_60183;
wire v_60184;
wire v_60185;
wire v_60186;
wire v_60187;
wire v_60188;
wire v_60189;
wire v_60190;
wire v_60191;
wire v_60192;
wire v_60193;
wire v_60194;
wire v_60195;
wire v_60196;
wire v_60197;
wire v_60198;
wire v_60199;
wire v_60200;
wire v_60201;
wire v_60202;
wire v_60203;
wire v_60204;
wire v_60205;
wire v_60206;
wire v_60207;
wire v_60208;
wire v_60209;
wire v_60210;
wire v_60211;
wire v_60212;
wire v_60213;
wire v_60214;
wire v_60215;
wire v_60216;
wire v_60217;
wire v_60218;
wire v_60219;
wire v_60220;
wire v_60221;
wire v_60222;
wire v_60223;
wire v_60224;
wire v_60225;
wire v_60226;
wire v_60227;
wire v_60228;
wire v_60229;
wire v_60230;
wire v_60231;
wire v_60232;
wire v_60233;
wire v_60234;
wire v_60235;
wire v_60236;
wire v_60237;
wire v_60238;
wire v_60239;
wire v_60240;
wire v_60241;
wire v_60242;
wire v_60243;
wire v_60244;
wire v_60245;
wire v_60246;
wire v_60247;
wire v_60248;
wire v_60249;
wire v_60250;
wire v_60251;
wire v_60252;
wire v_60253;
wire v_60254;
wire v_60255;
wire v_60256;
wire v_60257;
wire v_60258;
wire v_60259;
wire v_60260;
wire v_60261;
wire v_60262;
wire v_60263;
wire v_60264;
wire v_60265;
wire v_60266;
wire v_60267;
wire v_60268;
wire v_60269;
wire v_60270;
wire v_60271;
wire v_60272;
wire v_60273;
wire v_60274;
wire v_60275;
wire v_60276;
wire v_60277;
wire v_60278;
wire v_60279;
wire v_60280;
wire v_60281;
wire v_60282;
wire v_60283;
wire v_60284;
wire v_60285;
wire v_60286;
wire v_60287;
wire v_60288;
wire v_60289;
wire v_60290;
wire v_60291;
wire v_60292;
wire v_60293;
wire v_60294;
wire v_60295;
wire v_60296;
wire v_60297;
wire v_60298;
wire v_60299;
wire v_60300;
wire v_60301;
wire v_60302;
wire v_60303;
wire v_60304;
wire v_60305;
wire v_60306;
wire v_60307;
wire v_60308;
wire v_60309;
wire v_60310;
wire v_60311;
wire v_60312;
wire v_60313;
wire v_60314;
wire v_60315;
wire v_60316;
wire v_60317;
wire v_60318;
wire v_60319;
wire v_60320;
wire v_60321;
wire v_60322;
wire v_60323;
wire v_60324;
wire v_60325;
wire v_60326;
wire v_60328;
wire v_60329;
wire v_60330;
wire v_60331;
wire v_60332;
wire v_60333;
wire v_60334;
wire v_60335;
wire v_60336;
wire v_60337;
wire v_60338;
wire v_60339;
wire v_60340;
wire v_60341;
wire v_60342;
wire v_60343;
wire v_60344;
wire v_60345;
wire v_60346;
wire v_60347;
wire v_60348;
wire v_60349;
wire v_60350;
wire v_60351;
wire v_60352;
wire v_60353;
wire v_60354;
wire v_60355;
wire v_60356;
wire v_60357;
wire v_60358;
wire v_60359;
wire v_60360;
wire v_60361;
wire v_60362;
wire v_60363;
wire v_60364;
wire v_60365;
wire v_60366;
wire v_60367;
wire v_60368;
wire v_60369;
wire v_60370;
wire v_60371;
wire v_60372;
wire v_60373;
wire v_60374;
wire v_60375;
wire v_60376;
wire v_60377;
wire v_60378;
wire v_60379;
wire v_60380;
wire v_60381;
wire v_60382;
wire v_60383;
wire v_60384;
wire v_60385;
wire v_60386;
wire v_60387;
wire v_60388;
wire v_60389;
wire v_60390;
wire v_60391;
wire v_60392;
wire v_60393;
wire v_60394;
wire v_60395;
wire v_60396;
wire v_60397;
wire v_60398;
wire v_60399;
wire v_60400;
wire v_60401;
wire v_60402;
wire v_60403;
wire v_60404;
wire v_60405;
wire v_60406;
wire v_60407;
wire v_60408;
wire v_60409;
wire v_60410;
wire v_60411;
wire v_60412;
wire v_60413;
wire v_60414;
wire v_60415;
wire v_60416;
wire v_60417;
wire v_60418;
wire v_60419;
wire v_60420;
wire v_60421;
wire v_60422;
wire v_60423;
wire v_60424;
wire v_60425;
wire v_60426;
wire v_60427;
wire v_60428;
wire v_60429;
wire v_60430;
wire v_60431;
wire v_60432;
wire v_60433;
wire v_60434;
wire v_60435;
wire v_60436;
wire v_60437;
wire v_60438;
wire v_60439;
wire v_60440;
wire v_60441;
wire v_60442;
wire v_60443;
wire v_60444;
wire v_60445;
wire v_60446;
wire v_60447;
wire v_60448;
wire v_60449;
wire v_60450;
wire v_60451;
wire v_60452;
wire v_60453;
wire v_60454;
wire v_60455;
wire v_60456;
wire v_60457;
wire v_60458;
wire v_60459;
wire v_60460;
wire v_60461;
wire v_60462;
wire v_60463;
wire v_60464;
wire v_60465;
wire v_60466;
wire v_60467;
wire v_60468;
wire v_60469;
wire v_60470;
wire v_60471;
wire v_60472;
wire v_60473;
wire v_60474;
wire v_60475;
wire v_60476;
wire v_60477;
wire v_60478;
wire v_60479;
wire v_60480;
wire v_60481;
wire v_60482;
wire v_60483;
wire v_60484;
wire v_60485;
wire v_60486;
wire v_60487;
wire v_60488;
wire v_60489;
wire v_60490;
wire v_60491;
wire v_60492;
wire v_60493;
wire v_60494;
wire v_60495;
wire v_60496;
wire v_60497;
wire v_60498;
wire v_60499;
wire v_60500;
wire v_60501;
wire v_60502;
wire v_60503;
wire v_60504;
wire v_60505;
wire v_60506;
wire v_60507;
wire v_60508;
wire v_60509;
wire v_60510;
wire v_60511;
wire v_60512;
wire v_60513;
wire v_60514;
wire v_60515;
wire v_60516;
wire v_60517;
wire v_60518;
wire v_60519;
wire v_60520;
wire v_60521;
wire v_60522;
wire v_60523;
wire v_60524;
wire v_60525;
wire v_60526;
wire v_60527;
wire v_60528;
wire v_60529;
wire v_60530;
wire v_60531;
wire v_60532;
wire v_60533;
wire v_60534;
wire v_60535;
wire v_60536;
wire v_60537;
wire v_60538;
wire v_60539;
wire v_60540;
wire v_60541;
wire v_60542;
wire v_60543;
wire v_60544;
wire v_60545;
wire v_60546;
wire v_60547;
wire v_60548;
wire v_60549;
wire v_60550;
wire v_60551;
wire v_60552;
wire v_60553;
wire v_60554;
wire v_60555;
wire v_60556;
wire v_60557;
wire v_60558;
wire v_60559;
wire v_60560;
wire v_60561;
wire v_60562;
wire v_60563;
wire v_60564;
wire v_60565;
wire v_60566;
wire v_60567;
wire v_60568;
wire v_60569;
wire v_60571;
wire v_60572;
wire v_60573;
wire v_60574;
wire v_60575;
wire v_60576;
wire v_60577;
wire v_60578;
wire v_60579;
wire v_60580;
wire v_60581;
wire v_60582;
wire v_60583;
wire v_60584;
wire v_60585;
wire v_60586;
wire v_60587;
wire v_60588;
wire v_60589;
wire v_60590;
wire v_60591;
wire v_60592;
wire v_60593;
wire v_60594;
wire v_60595;
wire v_60596;
wire v_60597;
wire v_60598;
wire v_60599;
wire v_60600;
wire v_60601;
wire v_60602;
wire v_60603;
wire v_60604;
wire v_60605;
wire v_60606;
wire v_60607;
wire v_60608;
wire v_60609;
wire v_60610;
wire v_60611;
wire v_60612;
wire v_60613;
wire v_60614;
wire v_60615;
wire v_60616;
wire v_60617;
wire v_60618;
wire v_60619;
wire v_60620;
wire v_60621;
wire v_60622;
wire v_60623;
wire v_60624;
wire v_60625;
wire v_60626;
wire v_60627;
wire v_60628;
wire v_60629;
wire v_60630;
wire v_60631;
wire v_60632;
wire v_60633;
wire v_60634;
wire v_60635;
wire v_60636;
wire v_60637;
wire v_60638;
wire v_60639;
wire v_60640;
wire v_60641;
wire v_60642;
wire v_60643;
wire v_60644;
wire v_60645;
wire v_60646;
wire v_60647;
wire v_60648;
wire v_60649;
wire v_60650;
wire v_60651;
wire v_60652;
wire v_60653;
wire v_60654;
wire v_60655;
wire v_60656;
wire v_60657;
wire v_60658;
wire v_60659;
wire v_60660;
wire v_60661;
wire v_60662;
wire v_60663;
wire v_60664;
wire v_60665;
wire v_60666;
wire v_60667;
wire v_60668;
wire v_60669;
wire v_60670;
wire v_60671;
wire v_60672;
wire v_60673;
wire v_60674;
wire v_60675;
wire v_60676;
wire v_60677;
wire v_60678;
wire v_60679;
wire v_60680;
wire v_60681;
wire v_60682;
wire v_60683;
wire v_60684;
wire v_60685;
wire v_60686;
wire v_60687;
wire v_60688;
wire v_60689;
wire v_60690;
wire v_60691;
wire v_60692;
wire v_60693;
wire v_60694;
wire v_60695;
wire v_60696;
wire v_60697;
wire v_60698;
wire v_60699;
wire v_60700;
wire v_60701;
wire v_60702;
wire v_60703;
wire v_60704;
wire v_60705;
wire v_60706;
wire v_60707;
wire v_60708;
wire v_60709;
wire v_60710;
wire v_60711;
wire v_60712;
wire v_60713;
wire v_60714;
wire v_60715;
wire v_60716;
wire v_60717;
wire v_60718;
wire v_60719;
wire v_60720;
wire v_60721;
wire v_60722;
wire v_60723;
wire v_60724;
wire v_60725;
wire v_60726;
wire v_60727;
wire v_60728;
wire v_60729;
wire v_60730;
wire v_60731;
wire v_60732;
wire v_60733;
wire v_60734;
wire v_60735;
wire v_60736;
wire v_60737;
wire v_60738;
wire v_60739;
wire v_60740;
wire v_60741;
wire v_60742;
wire v_60743;
wire v_60744;
wire v_60745;
wire v_60746;
wire v_60747;
wire v_60748;
wire v_60749;
wire v_60750;
wire v_60751;
wire v_60752;
wire v_60753;
wire v_60754;
wire v_60755;
wire v_60756;
wire v_60757;
wire v_60758;
wire v_60759;
wire v_60760;
wire v_60761;
wire v_60762;
wire v_60763;
wire v_60764;
wire v_60765;
wire v_60766;
wire v_60767;
wire v_60768;
wire v_60769;
wire v_60770;
wire v_60771;
wire v_60772;
wire v_60773;
wire v_60774;
wire v_60775;
wire v_60776;
wire v_60777;
wire v_60778;
wire v_60779;
wire v_60780;
wire v_60781;
wire v_60782;
wire v_60783;
wire v_60784;
wire v_60785;
wire v_60786;
wire v_60787;
wire v_60788;
wire v_60789;
wire v_60790;
wire v_60791;
wire v_60792;
wire v_60793;
wire v_60794;
wire v_60795;
wire v_60796;
wire v_60797;
wire v_60798;
wire v_60799;
wire v_60800;
wire v_60801;
wire v_60802;
wire v_60803;
wire v_60804;
wire v_60805;
wire v_60806;
wire v_60807;
wire v_60808;
wire v_60809;
wire v_60810;
wire v_60811;
wire v_60812;
wire v_60814;
wire v_60815;
wire v_60816;
wire v_60817;
wire v_60818;
wire v_60819;
wire v_60820;
wire v_60821;
wire v_60822;
wire v_60823;
wire v_60824;
wire v_60825;
wire v_60826;
wire v_60827;
wire v_60828;
wire v_60829;
wire v_60830;
wire v_60831;
wire v_60832;
wire v_60833;
wire v_60834;
wire v_60835;
wire v_60836;
wire v_60837;
wire v_60838;
wire v_60839;
wire v_60840;
wire v_60841;
wire v_60842;
wire v_60843;
wire v_60844;
wire v_60845;
wire v_60846;
wire v_60847;
wire v_60848;
wire v_60849;
wire v_60850;
wire v_60851;
wire v_60852;
wire v_60853;
wire v_60854;
wire v_60855;
wire v_60856;
wire v_60857;
wire v_60858;
wire v_60859;
wire v_60860;
wire v_60861;
wire v_60862;
wire v_60863;
wire v_60864;
wire v_60865;
wire v_60866;
wire v_60867;
wire v_60868;
wire v_60869;
wire v_60870;
wire v_60871;
wire v_60872;
wire v_60873;
wire v_60874;
wire v_60875;
wire v_60876;
wire v_60877;
wire v_60878;
wire v_60879;
wire v_60880;
wire v_60881;
wire v_60882;
wire v_60883;
wire v_60884;
wire v_60885;
wire v_60886;
wire v_60887;
wire v_60888;
wire v_60889;
wire v_60890;
wire v_60891;
wire v_60892;
wire v_60893;
wire v_60894;
wire v_60895;
wire v_60896;
wire v_60897;
wire v_60898;
wire v_60899;
wire v_60900;
wire v_60901;
wire v_60902;
wire v_60903;
wire v_60904;
wire v_60905;
wire v_60906;
wire v_60907;
wire v_60908;
wire v_60909;
wire v_60910;
wire v_60911;
wire v_60912;
wire v_60913;
wire v_60914;
wire v_60915;
wire v_60916;
wire v_60917;
wire v_60918;
wire v_60919;
wire v_60920;
wire v_60921;
wire v_60922;
wire v_60923;
wire v_60924;
wire v_60925;
wire v_60926;
wire v_60927;
wire v_60928;
wire v_60929;
wire v_60930;
wire v_60931;
wire v_60932;
wire v_60933;
wire v_60934;
wire v_60935;
wire v_60936;
wire v_60937;
wire v_60938;
wire v_60939;
wire v_60940;
wire v_60941;
wire v_60942;
wire v_60943;
wire v_60944;
wire v_60945;
wire v_60946;
wire v_60947;
wire v_60948;
wire v_60949;
wire v_60950;
wire v_60951;
wire v_60952;
wire v_60953;
wire v_60954;
wire v_60955;
wire v_60956;
wire v_60957;
wire v_60958;
wire v_60959;
wire v_60960;
wire v_60961;
wire v_60962;
wire v_60963;
wire v_60964;
wire v_60965;
wire v_60966;
wire v_60967;
wire v_60968;
wire v_60969;
wire v_60970;
wire v_60971;
wire v_60972;
wire v_60973;
wire v_60974;
wire v_60975;
wire v_60976;
wire v_60977;
wire v_60978;
wire v_60979;
wire v_60980;
wire v_60981;
wire v_60982;
wire v_60983;
wire v_60984;
wire v_60985;
wire v_60986;
wire v_60987;
wire v_60988;
wire v_60989;
wire v_60990;
wire v_60991;
wire v_60992;
wire v_60993;
wire v_60994;
wire v_60995;
wire v_60996;
wire v_60997;
wire v_60998;
wire v_60999;
wire v_61000;
wire v_61001;
wire v_61002;
wire v_61003;
wire v_61004;
wire v_61005;
wire v_61006;
wire v_61007;
wire v_61008;
wire v_61009;
wire v_61010;
wire v_61011;
wire v_61012;
wire v_61013;
wire v_61014;
wire v_61015;
wire v_61016;
wire v_61017;
wire v_61018;
wire v_61019;
wire v_61020;
wire v_61021;
wire v_61022;
wire v_61023;
wire v_61024;
wire v_61025;
wire v_61026;
wire v_61027;
wire v_61028;
wire v_61029;
wire v_61030;
wire v_61031;
wire v_61032;
wire v_61033;
wire v_61034;
wire v_61035;
wire v_61036;
wire v_61037;
wire v_61038;
wire v_61039;
wire v_61040;
wire v_61041;
wire v_61042;
wire v_61043;
wire v_61044;
wire v_61045;
wire v_61046;
wire v_61047;
wire v_61048;
wire v_61049;
wire v_61050;
wire v_61051;
wire v_61052;
wire v_61053;
wire v_61054;
wire v_61055;
wire v_61057;
wire v_61058;
wire v_61059;
wire v_61060;
wire v_61061;
wire v_61062;
wire v_61063;
wire v_61064;
wire v_61065;
wire v_61066;
wire v_61067;
wire v_61068;
wire v_61069;
wire v_61070;
wire v_61071;
wire v_61072;
wire v_61073;
wire v_61074;
wire v_61075;
wire v_61076;
wire v_61077;
wire v_61078;
wire v_61079;
wire v_61080;
wire v_61081;
wire v_61082;
wire v_61083;
wire v_61084;
wire v_61085;
wire v_61086;
wire v_61087;
wire v_61088;
wire v_61089;
wire v_61090;
wire v_61091;
wire v_61092;
wire v_61093;
wire v_61094;
wire v_61095;
wire v_61096;
wire v_61097;
wire v_61098;
wire v_61099;
wire v_61100;
wire v_61101;
wire v_61102;
wire v_61103;
wire v_61104;
wire v_61105;
wire v_61106;
wire v_61107;
wire v_61108;
wire v_61109;
wire v_61110;
wire v_61111;
wire v_61112;
wire v_61113;
wire v_61114;
wire v_61115;
wire v_61116;
wire v_61117;
wire v_61118;
wire v_61119;
wire v_61120;
wire v_61121;
wire v_61122;
wire v_61123;
wire v_61124;
wire v_61125;
wire v_61126;
wire v_61127;
wire v_61128;
wire v_61129;
wire v_61130;
wire v_61131;
wire v_61132;
wire v_61133;
wire v_61134;
wire v_61135;
wire v_61136;
wire v_61137;
wire v_61138;
wire v_61139;
wire v_61140;
wire v_61141;
wire v_61142;
wire v_61143;
wire v_61144;
wire v_61145;
wire v_61146;
wire v_61147;
wire v_61148;
wire v_61149;
wire v_61150;
wire v_61151;
wire v_61152;
wire v_61153;
wire v_61154;
wire v_61155;
wire v_61156;
wire v_61157;
wire v_61158;
wire v_61159;
wire v_61160;
wire v_61161;
wire v_61162;
wire v_61163;
wire v_61164;
wire v_61165;
wire v_61166;
wire v_61167;
wire v_61168;
wire v_61169;
wire v_61170;
wire v_61171;
wire v_61172;
wire v_61173;
wire v_61174;
wire v_61175;
wire v_61176;
wire v_61177;
wire v_61178;
wire v_61179;
wire v_61180;
wire v_61181;
wire v_61182;
wire v_61183;
wire v_61184;
wire v_61185;
wire v_61186;
wire v_61187;
wire v_61188;
wire v_61189;
wire v_61190;
wire v_61191;
wire v_61192;
wire v_61193;
wire v_61194;
wire v_61195;
wire v_61196;
wire v_61197;
wire v_61198;
wire v_61199;
wire v_61200;
wire v_61201;
wire v_61202;
wire v_61203;
wire v_61204;
wire v_61205;
wire v_61206;
wire v_61207;
wire v_61208;
wire v_61209;
wire v_61210;
wire v_61211;
wire v_61212;
wire v_61213;
wire v_61214;
wire v_61215;
wire v_61216;
wire v_61217;
wire v_61218;
wire v_61219;
wire v_61220;
wire v_61221;
wire v_61222;
wire v_61223;
wire v_61224;
wire v_61225;
wire v_61226;
wire v_61227;
wire v_61228;
wire v_61229;
wire v_61230;
wire v_61231;
wire v_61232;
wire v_61233;
wire v_61234;
wire v_61235;
wire v_61236;
wire v_61237;
wire v_61238;
wire v_61239;
wire v_61240;
wire v_61241;
wire v_61242;
wire v_61243;
wire v_61244;
wire v_61245;
wire v_61246;
wire v_61247;
wire v_61248;
wire v_61249;
wire v_61250;
wire v_61251;
wire v_61252;
wire v_61253;
wire v_61254;
wire v_61255;
wire v_61256;
wire v_61257;
wire v_61258;
wire v_61259;
wire v_61260;
wire v_61261;
wire v_61262;
wire v_61263;
wire v_61264;
wire v_61265;
wire v_61266;
wire v_61267;
wire v_61268;
wire v_61269;
wire v_61270;
wire v_61271;
wire v_61272;
wire v_61273;
wire v_61274;
wire v_61275;
wire v_61276;
wire v_61277;
wire v_61278;
wire v_61279;
wire v_61280;
wire v_61281;
wire v_61282;
wire v_61283;
wire v_61284;
wire v_61285;
wire v_61286;
wire v_61287;
wire v_61288;
wire v_61289;
wire v_61290;
wire v_61291;
wire v_61292;
wire v_61293;
wire v_61294;
wire v_61295;
wire v_61296;
wire v_61297;
wire v_61298;
wire v_61300;
wire v_61301;
wire v_61302;
wire v_61303;
wire v_61304;
wire v_61305;
wire v_61306;
wire v_61307;
wire v_61308;
wire v_61309;
wire v_61310;
wire v_61311;
wire v_61312;
wire v_61313;
wire v_61314;
wire v_61315;
wire v_61316;
wire v_61317;
wire v_61318;
wire v_61319;
wire v_61320;
wire v_61321;
wire v_61322;
wire v_61323;
wire v_61324;
wire v_61325;
wire v_61326;
wire v_61327;
wire v_61328;
wire v_61329;
wire v_61330;
wire v_61331;
wire v_61332;
wire v_61333;
wire v_61334;
wire v_61335;
wire v_61336;
wire v_61337;
wire v_61338;
wire v_61339;
wire v_61340;
wire v_61341;
wire v_61342;
wire v_61343;
wire v_61344;
wire v_61345;
wire v_61346;
wire v_61347;
wire v_61348;
wire v_61349;
wire v_61350;
wire v_61351;
wire v_61352;
wire v_61353;
wire v_61354;
wire v_61355;
wire v_61356;
wire v_61357;
wire v_61358;
wire v_61359;
wire v_61360;
wire v_61361;
wire v_61362;
wire v_61363;
wire v_61364;
wire v_61365;
wire v_61366;
wire v_61367;
wire v_61368;
wire v_61369;
wire v_61370;
wire v_61371;
wire v_61372;
wire v_61373;
wire v_61374;
wire v_61375;
wire v_61376;
wire v_61377;
wire v_61378;
wire v_61379;
wire v_61380;
wire v_61381;
wire v_61382;
wire v_61383;
wire v_61384;
wire v_61385;
wire v_61386;
wire v_61387;
wire v_61388;
wire v_61389;
wire v_61390;
wire v_61391;
wire v_61392;
wire v_61393;
wire v_61394;
wire v_61395;
wire v_61396;
wire v_61397;
wire v_61398;
wire v_61399;
wire v_61400;
wire v_61401;
wire v_61402;
wire v_61403;
wire v_61404;
wire v_61405;
wire v_61406;
wire v_61407;
wire v_61408;
wire v_61409;
wire v_61410;
wire v_61411;
wire v_61412;
wire v_61413;
wire v_61414;
wire v_61415;
wire v_61416;
wire v_61417;
wire v_61418;
wire v_61419;
wire v_61420;
wire v_61421;
wire v_61422;
wire v_61423;
wire v_61424;
wire v_61425;
wire v_61426;
wire v_61427;
wire v_61428;
wire v_61429;
wire v_61430;
wire v_61431;
wire v_61432;
wire v_61433;
wire v_61434;
wire v_61435;
wire v_61436;
wire v_61437;
wire v_61438;
wire v_61439;
wire v_61440;
wire v_61441;
wire v_61442;
wire v_61443;
wire v_61444;
wire v_61445;
wire v_61446;
wire v_61447;
wire v_61448;
wire v_61449;
wire v_61450;
wire v_61451;
wire v_61452;
wire v_61453;
wire v_61454;
wire v_61455;
wire v_61456;
wire v_61457;
wire v_61458;
wire v_61459;
wire v_61460;
wire v_61461;
wire v_61462;
wire v_61463;
wire v_61464;
wire v_61465;
wire v_61466;
wire v_61467;
wire v_61468;
wire v_61469;
wire v_61470;
wire v_61471;
wire v_61472;
wire v_61473;
wire v_61474;
wire v_61475;
wire v_61476;
wire v_61477;
wire v_61478;
wire v_61479;
wire v_61480;
wire v_61481;
wire v_61482;
wire v_61483;
wire v_61484;
wire v_61485;
wire v_61486;
wire v_61487;
wire v_61488;
wire v_61489;
wire v_61490;
wire v_61491;
wire v_61492;
wire v_61493;
wire v_61494;
wire v_61495;
wire v_61496;
wire v_61497;
wire v_61498;
wire v_61499;
wire v_61500;
wire v_61501;
wire v_61502;
wire v_61503;
wire v_61504;
wire v_61505;
wire v_61506;
wire v_61507;
wire v_61508;
wire v_61509;
wire v_61510;
wire v_61511;
wire v_61512;
wire v_61513;
wire v_61514;
wire v_61515;
wire v_61516;
wire v_61517;
wire v_61518;
wire v_61519;
wire v_61520;
wire v_61521;
wire v_61522;
wire v_61523;
wire v_61524;
wire v_61525;
wire v_61526;
wire v_61527;
wire v_61528;
wire v_61529;
wire v_61530;
wire v_61531;
wire v_61532;
wire v_61533;
wire v_61534;
wire v_61535;
wire v_61536;
wire v_61537;
wire v_61538;
wire v_61539;
wire v_61540;
wire v_61541;
wire v_61543;
wire v_61544;
wire v_61545;
wire v_61546;
wire v_61547;
wire v_61548;
wire v_61549;
wire v_61550;
wire v_61551;
wire v_61552;
wire v_61553;
wire v_61554;
wire v_61555;
wire v_61556;
wire v_61557;
wire v_61558;
wire v_61559;
wire v_61560;
wire v_61561;
wire v_61562;
wire v_61563;
wire v_61564;
wire v_61565;
wire v_61566;
wire v_61567;
wire v_61568;
wire v_61569;
wire v_61570;
wire v_61571;
wire v_61572;
wire v_61573;
wire v_61574;
wire v_61575;
wire v_61576;
wire v_61577;
wire v_61578;
wire v_61579;
wire v_61580;
wire v_61581;
wire v_61582;
wire v_61583;
wire v_61584;
wire v_61585;
wire v_61586;
wire v_61587;
wire v_61588;
wire v_61589;
wire v_61590;
wire v_61591;
wire v_61592;
wire v_61593;
wire v_61594;
wire v_61595;
wire v_61596;
wire v_61597;
wire v_61598;
wire v_61599;
wire v_61600;
wire v_61601;
wire v_61602;
wire v_61603;
wire v_61604;
wire v_61605;
wire v_61606;
wire v_61607;
wire v_61608;
wire v_61609;
wire v_61610;
wire v_61611;
wire v_61612;
wire v_61613;
wire v_61614;
wire v_61615;
wire v_61616;
wire v_61617;
wire v_61618;
wire v_61619;
wire v_61620;
wire v_61621;
wire v_61622;
wire v_61623;
wire v_61624;
wire v_61625;
wire v_61626;
wire v_61627;
wire v_61628;
wire v_61629;
wire v_61630;
wire v_61631;
wire v_61632;
wire v_61633;
wire v_61634;
wire v_61635;
wire v_61636;
wire v_61637;
wire v_61638;
wire v_61639;
wire v_61640;
wire v_61641;
wire v_61642;
wire v_61643;
wire v_61644;
wire v_61645;
wire v_61646;
wire v_61647;
wire v_61648;
wire v_61649;
wire v_61650;
wire v_61651;
wire v_61652;
wire v_61653;
wire v_61654;
wire v_61655;
wire v_61656;
wire v_61657;
wire v_61658;
wire v_61659;
wire v_61660;
wire v_61661;
wire v_61662;
wire v_61663;
wire v_61664;
wire v_61665;
wire v_61666;
wire v_61667;
wire v_61668;
wire v_61669;
wire v_61670;
wire v_61671;
wire v_61672;
wire v_61673;
wire v_61674;
wire v_61675;
wire v_61676;
wire v_61677;
wire v_61678;
wire v_61679;
wire v_61680;
wire v_61681;
wire v_61682;
wire v_61683;
wire v_61684;
wire v_61685;
wire v_61686;
wire v_61687;
wire v_61688;
wire v_61689;
wire v_61690;
wire v_61691;
wire v_61692;
wire v_61693;
wire v_61694;
wire v_61695;
wire v_61696;
wire v_61697;
wire v_61698;
wire v_61699;
wire v_61700;
wire v_61701;
wire v_61702;
wire v_61703;
wire v_61704;
wire v_61705;
wire v_61706;
wire v_61707;
wire v_61708;
wire v_61709;
wire v_61710;
wire v_61711;
wire v_61712;
wire v_61713;
wire v_61714;
wire v_61715;
wire v_61716;
wire v_61717;
wire v_61718;
wire v_61719;
wire v_61720;
wire v_61721;
wire v_61722;
wire v_61723;
wire v_61724;
wire v_61725;
wire v_61726;
wire v_61727;
wire v_61728;
wire v_61729;
wire v_61730;
wire v_61731;
wire v_61732;
wire v_61733;
wire v_61734;
wire v_61735;
wire v_61736;
wire v_61737;
wire v_61738;
wire v_61739;
wire v_61740;
wire v_61741;
wire v_61742;
wire v_61743;
wire v_61744;
wire v_61745;
wire v_61746;
wire v_61747;
wire v_61748;
wire v_61749;
wire v_61750;
wire v_61751;
wire v_61752;
wire v_61753;
wire v_61754;
wire v_61755;
wire v_61756;
wire v_61757;
wire v_61758;
wire v_61759;
wire v_61760;
wire v_61761;
wire v_61762;
wire v_61763;
wire v_61764;
wire v_61765;
wire v_61766;
wire v_61767;
wire v_61768;
wire v_61769;
wire v_61770;
wire v_61771;
wire v_61772;
wire v_61773;
wire v_61774;
wire v_61775;
wire v_61776;
wire v_61777;
wire v_61778;
wire v_61779;
wire v_61780;
wire v_61781;
wire v_61782;
wire v_61783;
wire v_61784;
wire v_61786;
wire v_61787;
wire v_61788;
wire v_61789;
wire v_61790;
wire v_61791;
wire v_61792;
wire v_61793;
wire v_61794;
wire v_61795;
wire v_61796;
wire v_61797;
wire v_61798;
wire v_61799;
wire v_61800;
wire v_61801;
wire v_61802;
wire v_61803;
wire v_61804;
wire v_61805;
wire v_61806;
wire v_61807;
wire v_61808;
wire v_61809;
wire v_61810;
wire v_61811;
wire v_61812;
wire v_61813;
wire v_61814;
wire v_61815;
wire v_61816;
wire v_61817;
wire v_61818;
wire v_61819;
wire v_61820;
wire v_61821;
wire v_61822;
wire v_61823;
wire v_61824;
wire v_61825;
wire v_61826;
wire v_61827;
wire v_61828;
wire v_61829;
wire v_61830;
wire v_61831;
wire v_61832;
wire v_61833;
wire v_61834;
wire v_61835;
wire v_61836;
wire v_61837;
wire v_61838;
wire v_61839;
wire v_61840;
wire v_61841;
wire v_61842;
wire v_61843;
wire v_61844;
wire v_61845;
wire v_61846;
wire v_61847;
wire v_61848;
wire v_61849;
wire v_61850;
wire v_61851;
wire v_61852;
wire v_61853;
wire v_61854;
wire v_61855;
wire v_61856;
wire v_61857;
wire v_61858;
wire v_61859;
wire v_61860;
wire v_61861;
wire v_61862;
wire v_61863;
wire v_61864;
wire v_61865;
wire v_61866;
wire v_61867;
wire v_61868;
wire v_61869;
wire v_61870;
wire v_61871;
wire v_61872;
wire v_61873;
wire v_61874;
wire v_61875;
wire v_61876;
wire v_61877;
wire v_61878;
wire v_61879;
wire v_61880;
wire v_61881;
wire v_61882;
wire v_61883;
wire v_61884;
wire v_61885;
wire v_61886;
wire v_61887;
wire v_61888;
wire v_61889;
wire v_61890;
wire v_61891;
wire v_61892;
wire v_61893;
wire v_61894;
wire v_61895;
wire v_61896;
wire v_61897;
wire v_61898;
wire v_61899;
wire v_61900;
wire v_61901;
wire v_61902;
wire v_61903;
wire v_61904;
wire v_61905;
wire v_61906;
wire v_61907;
wire v_61908;
wire v_61909;
wire v_61910;
wire v_61911;
wire v_61912;
wire v_61913;
wire v_61914;
wire v_61915;
wire v_61916;
wire v_61917;
wire v_61918;
wire v_61919;
wire v_61920;
wire v_61921;
wire v_61922;
wire v_61923;
wire v_61924;
wire v_61925;
wire v_61926;
wire v_61927;
wire v_61928;
wire v_61929;
wire v_61930;
wire v_61931;
wire v_61932;
wire v_61933;
wire v_61934;
wire v_61935;
wire v_61936;
wire v_61937;
wire v_61938;
wire v_61939;
wire v_61940;
wire v_61941;
wire v_61942;
wire v_61943;
wire v_61944;
wire v_61945;
wire v_61946;
wire v_61947;
wire v_61948;
wire v_61949;
wire v_61950;
wire v_61951;
wire v_61952;
wire v_61953;
wire v_61954;
wire v_61955;
wire v_61956;
wire v_61957;
wire v_61958;
wire v_61959;
wire v_61960;
wire v_61961;
wire v_61962;
wire v_61963;
wire v_61964;
wire v_61965;
wire v_61966;
wire v_61967;
wire v_61968;
wire v_61969;
wire v_61970;
wire v_61971;
wire v_61972;
wire v_61973;
wire v_61974;
wire v_61975;
wire v_61976;
wire v_61977;
wire v_61978;
wire v_61979;
wire v_61980;
wire v_61981;
wire v_61982;
wire v_61983;
wire v_61984;
wire v_61985;
wire v_61986;
wire v_61987;
wire v_61988;
wire v_61989;
wire v_61990;
wire v_61991;
wire v_61992;
wire v_61993;
wire v_61994;
wire v_61995;
wire v_61996;
wire v_61997;
wire v_61998;
wire v_61999;
wire v_62000;
wire v_62001;
wire v_62002;
wire v_62003;
wire v_62004;
wire v_62005;
wire v_62006;
wire v_62007;
wire v_62008;
wire v_62009;
wire v_62010;
wire v_62011;
wire v_62012;
wire v_62013;
wire v_62014;
wire v_62015;
wire v_62016;
wire v_62017;
wire v_62018;
wire v_62019;
wire v_62020;
wire v_62021;
wire v_62022;
wire v_62023;
wire v_62024;
wire v_62025;
wire v_62026;
wire v_62027;
wire v_62029;
wire v_62030;
wire v_62031;
wire v_62032;
wire v_62033;
wire v_62034;
wire v_62035;
wire v_62036;
wire v_62037;
wire v_62038;
wire v_62039;
wire v_62040;
wire v_62041;
wire v_62042;
wire v_62043;
wire v_62044;
wire v_62045;
wire v_62046;
wire v_62047;
wire v_62048;
wire v_62049;
wire v_62050;
wire v_62051;
wire v_62052;
wire v_62053;
wire v_62054;
wire v_62055;
wire v_62056;
wire v_62057;
wire v_62058;
wire v_62059;
wire v_62060;
wire v_62061;
wire v_62062;
wire v_62063;
wire v_62064;
wire v_62065;
wire v_62066;
wire v_62067;
wire v_62068;
wire v_62069;
wire v_62070;
wire v_62071;
wire v_62072;
wire v_62073;
wire v_62074;
wire v_62075;
wire v_62076;
wire v_62077;
wire v_62078;
wire v_62079;
wire v_62080;
wire v_62081;
wire v_62082;
wire v_62083;
wire v_62084;
wire v_62085;
wire v_62086;
wire v_62087;
wire v_62088;
wire v_62089;
wire v_62090;
wire v_62091;
wire v_62092;
wire v_62093;
wire v_62094;
wire v_62095;
wire v_62096;
wire v_62097;
wire v_62098;
wire v_62099;
wire v_62100;
wire v_62101;
wire v_62102;
wire v_62103;
wire v_62104;
wire v_62105;
wire v_62106;
wire v_62107;
wire v_62108;
wire v_62109;
wire v_62110;
wire v_62111;
wire v_62112;
wire v_62113;
wire v_62114;
wire v_62115;
wire v_62116;
wire v_62117;
wire v_62118;
wire v_62119;
wire v_62120;
wire v_62121;
wire v_62122;
wire v_62123;
wire v_62124;
wire v_62125;
wire v_62126;
wire v_62127;
wire v_62128;
wire v_62129;
wire v_62130;
wire v_62131;
wire v_62132;
wire v_62133;
wire v_62134;
wire v_62135;
wire v_62136;
wire v_62137;
wire v_62138;
wire v_62139;
wire v_62140;
wire v_62141;
wire v_62142;
wire v_62143;
wire v_62144;
wire v_62145;
wire v_62146;
wire v_62147;
wire v_62148;
wire v_62149;
wire v_62150;
wire v_62151;
wire v_62152;
wire v_62153;
wire v_62154;
wire v_62155;
wire v_62156;
wire v_62157;
wire v_62158;
wire v_62159;
wire v_62160;
wire v_62161;
wire v_62162;
wire v_62163;
wire v_62164;
wire v_62165;
wire v_62166;
wire v_62167;
wire v_62168;
wire v_62169;
wire v_62170;
wire v_62171;
wire v_62172;
wire v_62173;
wire v_62174;
wire v_62175;
wire v_62176;
wire v_62177;
wire v_62178;
wire v_62179;
wire v_62180;
wire v_62181;
wire v_62182;
wire v_62183;
wire v_62184;
wire v_62185;
wire v_62186;
wire v_62187;
wire v_62188;
wire v_62189;
wire v_62190;
wire v_62191;
wire v_62192;
wire v_62193;
wire v_62194;
wire v_62195;
wire v_62196;
wire v_62197;
wire v_62198;
wire v_62199;
wire v_62200;
wire v_62201;
wire v_62202;
wire v_62203;
wire v_62204;
wire v_62205;
wire v_62206;
wire v_62207;
wire v_62208;
wire v_62209;
wire v_62210;
wire v_62211;
wire v_62212;
wire v_62213;
wire v_62214;
wire v_62215;
wire v_62216;
wire v_62217;
wire v_62218;
wire v_62219;
wire v_62220;
wire v_62221;
wire v_62222;
wire v_62223;
wire v_62224;
wire v_62225;
wire v_62226;
wire v_62227;
wire v_62228;
wire v_62229;
wire v_62230;
wire v_62231;
wire v_62232;
wire v_62233;
wire v_62234;
wire v_62235;
wire v_62236;
wire v_62237;
wire v_62238;
wire v_62239;
wire v_62240;
wire v_62241;
wire v_62242;
wire v_62243;
wire v_62244;
wire v_62245;
wire v_62246;
wire v_62247;
wire v_62248;
wire v_62249;
wire v_62250;
wire v_62251;
wire v_62252;
wire v_62253;
wire v_62254;
wire v_62255;
wire v_62256;
wire v_62257;
wire v_62258;
wire v_62259;
wire v_62260;
wire v_62261;
wire v_62262;
wire v_62263;
wire v_62264;
wire v_62265;
wire v_62266;
wire v_62267;
wire v_62268;
wire v_62269;
wire v_62270;
wire v_62271;
wire v_62272;
wire v_62273;
wire v_62274;
wire v_62275;
wire v_62276;
wire v_62277;
wire v_62278;
wire v_62279;
wire v_62280;
wire v_62281;
wire v_62282;
wire v_62283;
wire v_62284;
wire v_62285;
wire v_62286;
wire v_62287;
wire v_62288;
wire v_62289;
wire v_62290;
wire v_62291;
wire v_62292;
wire v_62293;
wire v_62294;
wire v_62295;
wire v_62296;
wire v_62297;
wire v_62298;
wire v_62299;
wire v_62300;
wire v_62301;
wire v_62302;
wire v_62303;
wire v_62304;
wire v_62305;
wire v_62306;
wire v_62307;
wire v_62308;
wire v_62309;
wire v_62310;
wire v_62311;
wire v_62312;
wire v_62313;
wire v_62314;
wire v_62315;
wire v_62316;
wire v_62317;
wire v_62318;
wire v_62319;
wire v_62320;
wire v_62321;
wire v_62322;
wire v_62323;
wire v_62324;
wire v_62325;
wire v_62326;
wire v_62327;
wire v_62328;
wire v_62329;
wire v_62330;
wire v_62331;
wire v_62332;
wire v_62333;
wire v_62334;
wire v_62335;
wire v_62336;
wire v_62337;
wire v_62338;
wire v_62339;
wire v_62340;
wire v_62341;
wire v_62342;
wire v_62343;
wire v_62344;
wire v_62345;
wire v_62346;
wire v_62347;
wire v_62348;
wire v_62349;
wire v_62350;
wire v_62351;
wire v_62352;
wire v_62353;
wire v_62354;
wire v_62355;
wire v_62356;
wire v_62357;
wire v_62358;
wire v_62359;
wire v_62360;
wire v_62361;
wire v_62362;
wire v_62363;
wire v_62364;
wire v_62365;
wire v_62366;
wire v_62367;
wire v_62368;
wire v_62369;
wire v_62370;
wire v_62371;
wire v_62372;
wire v_62373;
wire v_62374;
wire v_62375;
wire v_62376;
wire v_62377;
wire v_62378;
wire v_62379;
wire v_62380;
wire v_62381;
wire v_62382;
wire v_62383;
wire v_62384;
wire v_62385;
wire v_62386;
wire v_62387;
wire v_62388;
wire v_62389;
wire v_62390;
wire v_62391;
wire v_62392;
wire v_62393;
wire v_62394;
wire v_62395;
wire v_62396;
wire v_62397;
wire v_62398;
wire v_62399;
wire v_62400;
wire v_62401;
wire v_62402;
wire v_62403;
wire v_62404;
wire v_62405;
wire v_62406;
wire v_62407;
wire v_62408;
wire v_62409;
wire v_62410;
wire v_62411;
wire v_62412;
wire v_62413;
wire v_62414;
wire v_62415;
wire v_62416;
wire v_62417;
wire v_62418;
wire v_62419;
wire v_62421;
wire v_62422;
wire v_62423;
wire v_62424;
wire v_62425;
wire v_62426;
wire v_62427;
wire v_62428;
wire v_62429;
wire v_62430;
wire v_62431;
wire v_62432;
wire v_62433;
wire v_62434;
wire v_62435;
wire v_62436;
wire v_62437;
wire v_62438;
wire v_62439;
wire v_62440;
wire v_62441;
wire v_62442;
wire v_62443;
wire v_62444;
wire v_62445;
wire v_62446;
wire v_62447;
wire v_62448;
wire v_62449;
wire v_62450;
wire v_62451;
wire v_62452;
wire v_62453;
wire v_62454;
wire v_62455;
wire v_62456;
wire v_62457;
wire v_62458;
wire v_62459;
wire v_62460;
wire v_62461;
wire v_62462;
wire v_62463;
wire v_62464;
wire v_62465;
wire v_62466;
wire v_62467;
wire v_62468;
wire v_62469;
wire v_62470;
wire v_62471;
wire v_62472;
wire v_62473;
wire v_62474;
wire v_62475;
wire v_62476;
wire v_62477;
wire v_62478;
wire v_62479;
wire v_62480;
wire v_62481;
wire v_62482;
wire v_62483;
wire v_62484;
wire v_62485;
wire v_62486;
wire v_62487;
wire v_62488;
wire v_62489;
wire v_62490;
wire v_62491;
wire v_62492;
wire v_62493;
wire v_62494;
wire v_62495;
wire v_62496;
wire v_62497;
wire v_62498;
wire v_62499;
wire v_62500;
wire v_62501;
wire v_62502;
wire v_62503;
wire v_62504;
wire v_62505;
wire v_62506;
wire v_62507;
wire v_62508;
wire v_62509;
wire v_62510;
wire v_62511;
wire v_62512;
wire v_62513;
wire v_62515;
wire v_62517;
wire v_62518;
wire v_62519;
wire v_62521;
wire v_62522;
wire v_62523;
wire v_62525;
wire v_62526;
wire v_62527;
wire v_62529;
wire v_62530;
wire v_62532;
wire v_62533;
wire v_62534;
wire v_62536;
wire v_62537;
wire v_62538;
wire v_62540;
wire v_62541;
wire v_62542;
wire v_62544;
wire v_62545;
wire v_62546;
wire v_62548;
wire v_62549;
wire v_62550;
wire v_62552;
wire v_62553;
wire v_62554;
wire v_62556;
wire v_62557;
wire v_62558;
wire v_62560;
wire v_62561;
wire v_62562;
wire v_62564;
wire v_62565;
wire v_62566;
wire v_62568;
wire v_62569;
wire v_62570;
wire v_62572;
wire v_62573;
wire v_62574;
wire v_62576;
wire v_62577;
wire v_62578;
wire v_62580;
wire v_62581;
wire v_62582;
wire v_62583;
wire v_62584;
wire v_62585;
wire v_62586;
wire v_62587;
wire v_62588;
wire v_62589;
wire v_62590;
wire v_62591;
wire v_62592;
wire v_62593;
wire v_62594;
wire v_62595;
wire v_62596;
wire v_62597;
wire v_62598;
wire v_62599;
wire v_62600;
wire v_62601;
wire v_62602;
wire v_62603;
wire v_62604;
wire v_62605;
wire v_62606;
wire v_62607;
wire v_62608;
wire v_62609;
wire v_62610;
wire v_62611;
wire v_62612;
wire v_62613;
wire v_62614;
wire v_62615;
wire v_62616;
wire v_62617;
wire v_62618;
wire v_62619;
wire v_62620;
wire v_62621;
wire v_62622;
wire v_62623;
wire v_62624;
wire v_62625;
wire v_62626;
wire v_62627;
wire v_62628;
wire v_62629;
wire v_62630;
wire v_62631;
wire v_62632;
wire v_62633;
wire v_62634;
wire v_62635;
wire v_62636;
wire v_62637;
wire v_62638;
wire v_62639;
wire v_62640;
wire v_62641;
wire v_62642;
wire v_62643;
wire v_62644;
wire v_62645;
wire v_62646;
wire v_62647;
wire v_62648;
wire v_62649;
wire v_62650;
wire v_62651;
wire v_62652;
wire v_62653;
wire v_62654;
wire v_62655;
wire v_62656;
wire v_62657;
wire v_62658;
wire v_62659;
wire v_62660;
wire v_62661;
wire v_62662;
wire v_62663;
wire v_62664;
wire v_62665;
wire v_62666;
wire v_62667;
wire v_62668;
wire v_62669;
wire v_62670;
wire v_62671;
wire v_62672;
wire v_62673;
wire v_62674;
wire v_62675;
wire v_62676;
wire v_62677;
wire v_62678;
wire v_62679;
wire v_62680;
wire v_62681;
wire v_62682;
wire v_62683;
wire v_62684;
wire v_62685;
wire v_62686;
wire v_62687;
wire v_62688;
wire v_62689;
wire v_62690;
wire v_62691;
wire v_62692;
wire v_62693;
wire v_62694;
wire v_62695;
wire v_62696;
wire v_62697;
wire v_62698;
wire v_62699;
wire v_62700;
wire v_62701;
wire v_62702;
wire v_62703;
wire v_62704;
wire v_62705;
wire v_62706;
wire v_62707;
wire v_62708;
wire v_62709;
wire v_62710;
wire v_62711;
wire v_62712;
wire v_62713;
wire v_62714;
wire v_62715;
wire v_62716;
wire v_62717;
wire v_62718;
wire v_62719;
wire v_62720;
wire v_62721;
wire v_62722;
wire v_62723;
wire v_62724;
wire v_62725;
wire v_62726;
wire v_62727;
wire v_62728;
wire v_62729;
wire v_62730;
wire v_62731;
wire v_62732;
wire v_62733;
wire v_62734;
wire v_62735;
wire v_62736;
wire v_62737;
wire v_62738;
wire v_62739;
wire v_62740;
wire v_62741;
wire v_62742;
wire v_62743;
wire v_62744;
wire v_62745;
wire v_62746;
wire v_62747;
wire v_62748;
wire v_62749;
wire v_62750;
wire v_62751;
wire v_62752;
wire v_62753;
wire v_62754;
wire v_62755;
wire v_62756;
wire v_62757;
wire v_62758;
wire v_62759;
wire v_62760;
wire v_62761;
wire v_62762;
wire v_62763;
wire v_62764;
wire v_62765;
wire v_62766;
wire v_62767;
wire v_62768;
wire v_62769;
wire v_62770;
wire v_62771;
wire v_62772;
wire v_62773;
wire v_62775;
wire v_62776;
wire v_62777;
wire v_62778;
wire v_62779;
wire v_62780;
wire v_62781;
wire v_62782;
wire v_62783;
wire v_62784;
wire v_62785;
wire v_62786;
wire v_62787;
wire v_62788;
wire v_62789;
wire v_62790;
wire v_62791;
wire v_62792;
wire v_62793;
wire v_62794;
wire v_62795;
wire v_62796;
wire v_62797;
wire v_62798;
wire v_62799;
wire v_62800;
wire v_62801;
wire v_62802;
wire v_62803;
wire v_62804;
wire v_62805;
wire v_62806;
wire v_62807;
wire v_62808;
wire v_62809;
wire v_62810;
wire v_62811;
wire v_62812;
wire v_62813;
wire v_62814;
wire v_62815;
wire v_62816;
wire v_62817;
wire v_62818;
wire v_62819;
wire v_62820;
wire v_62821;
wire v_62822;
wire v_62823;
wire v_62824;
wire v_62825;
wire v_62826;
wire v_62827;
wire v_62828;
wire v_62829;
wire v_62830;
wire v_62831;
wire v_62832;
wire v_62833;
wire v_62834;
wire v_62835;
wire v_62836;
wire v_62837;
wire v_62838;
wire v_62839;
wire v_62840;
wire v_62841;
wire v_62842;
wire v_62843;
wire v_62844;
wire v_62845;
wire v_62846;
wire v_62847;
wire v_62848;
wire v_62849;
wire v_62850;
wire v_62851;
wire v_62852;
wire v_62853;
wire v_62854;
wire v_62855;
wire v_62856;
wire v_62857;
wire v_62858;
wire v_62859;
wire v_62860;
wire v_62861;
wire v_62862;
wire v_62863;
wire v_62864;
wire v_62865;
wire v_62866;
wire v_62867;
wire v_62868;
wire v_62869;
wire v_62870;
wire v_62871;
wire v_62872;
wire v_62873;
wire v_62874;
wire v_62875;
wire v_62876;
wire v_62877;
wire v_62878;
wire v_62879;
wire v_62880;
wire v_62881;
wire v_62882;
wire v_62883;
wire v_62884;
wire v_62885;
wire v_62886;
wire v_62887;
wire v_62888;
wire v_62889;
wire v_62890;
wire v_62891;
wire v_62892;
wire v_62893;
wire v_62894;
wire v_62895;
wire v_62896;
wire v_62897;
wire v_62898;
wire v_62899;
wire v_62900;
wire v_62901;
wire v_62902;
wire v_62903;
wire v_62904;
wire v_62905;
wire v_62906;
wire v_62907;
wire v_62908;
wire v_62909;
wire v_62910;
wire v_62911;
wire v_62912;
wire v_62913;
wire v_62914;
wire v_62915;
wire v_62916;
wire v_62917;
wire v_62918;
wire v_62919;
wire v_62920;
wire v_62921;
wire v_62922;
wire v_62923;
wire v_62924;
wire v_62925;
wire v_62926;
wire v_62927;
wire v_62928;
wire v_62929;
wire v_62930;
wire v_62931;
wire v_62932;
wire v_62933;
wire v_62934;
wire v_62935;
wire v_62936;
wire v_62937;
wire v_62938;
wire v_62939;
wire v_62940;
wire v_62941;
wire v_62942;
wire v_62943;
wire v_62944;
wire v_62945;
wire v_62946;
wire v_62947;
wire v_62948;
wire v_62949;
wire v_62950;
wire v_62951;
wire v_62952;
wire v_62953;
wire v_62954;
wire v_62955;
wire v_62956;
wire v_62957;
wire v_62958;
wire v_62959;
wire v_62960;
wire v_62961;
wire v_62962;
wire v_62963;
wire v_62964;
wire v_62965;
wire v_62966;
wire v_62967;
wire v_62968;
wire v_62969;
wire v_62970;
wire v_62971;
wire v_62972;
wire v_62973;
wire v_62974;
wire v_62975;
wire v_62976;
wire v_62977;
wire v_62978;
wire v_62979;
wire v_62980;
wire v_62981;
wire v_62982;
wire v_62983;
wire v_62984;
wire v_62985;
wire v_62986;
wire v_62987;
wire v_62988;
wire v_62989;
wire v_62990;
wire v_62991;
wire v_62992;
wire v_62993;
wire v_62994;
wire v_62995;
wire v_62996;
wire v_62997;
wire v_62998;
wire v_62999;
wire v_63000;
wire v_63001;
wire v_63002;
wire v_63003;
wire v_63004;
wire v_63005;
wire v_63006;
wire v_63007;
wire v_63008;
wire v_63009;
wire v_63010;
wire v_63011;
wire v_63012;
wire v_63013;
wire v_63014;
wire v_63015;
wire v_63016;
wire v_63018;
wire v_63019;
wire v_63020;
wire v_63021;
wire v_63022;
wire v_63023;
wire v_63024;
wire v_63025;
wire v_63026;
wire v_63027;
wire v_63028;
wire v_63029;
wire v_63030;
wire v_63031;
wire v_63032;
wire v_63033;
wire v_63034;
wire v_63035;
wire v_63036;
wire v_63037;
wire v_63038;
wire v_63039;
wire v_63040;
wire v_63041;
wire v_63042;
wire v_63043;
wire v_63044;
wire v_63045;
wire v_63046;
wire v_63047;
wire v_63048;
wire v_63049;
wire v_63050;
wire v_63051;
wire v_63052;
wire v_63053;
wire v_63054;
wire v_63055;
wire v_63056;
wire v_63057;
wire v_63058;
wire v_63059;
wire v_63060;
wire v_63061;
wire v_63062;
wire v_63063;
wire v_63064;
wire v_63065;
wire v_63066;
wire v_63067;
wire v_63068;
wire v_63069;
wire v_63070;
wire v_63071;
wire v_63072;
wire v_63073;
wire v_63074;
wire v_63075;
wire v_63076;
wire v_63077;
wire v_63078;
wire v_63079;
wire v_63080;
wire v_63081;
wire v_63082;
wire v_63083;
wire v_63084;
wire v_63085;
wire v_63086;
wire v_63087;
wire v_63088;
wire v_63089;
wire v_63090;
wire v_63091;
wire v_63092;
wire v_63093;
wire v_63094;
wire v_63095;
wire v_63096;
wire v_63097;
wire v_63098;
wire v_63099;
wire v_63100;
wire v_63101;
wire v_63102;
wire v_63103;
wire v_63104;
wire v_63105;
wire v_63106;
wire v_63107;
wire v_63108;
wire v_63109;
wire v_63110;
wire v_63111;
wire v_63112;
wire v_63113;
wire v_63114;
wire v_63115;
wire v_63116;
wire v_63117;
wire v_63118;
wire v_63119;
wire v_63120;
wire v_63121;
wire v_63122;
wire v_63123;
wire v_63124;
wire v_63125;
wire v_63126;
wire v_63127;
wire v_63128;
wire v_63129;
wire v_63130;
wire v_63131;
wire v_63132;
wire v_63133;
wire v_63134;
wire v_63135;
wire v_63136;
wire v_63137;
wire v_63138;
wire v_63139;
wire v_63140;
wire v_63141;
wire v_63142;
wire v_63143;
wire v_63144;
wire v_63145;
wire v_63146;
wire v_63147;
wire v_63148;
wire v_63149;
wire v_63150;
wire v_63151;
wire v_63152;
wire v_63153;
wire v_63154;
wire v_63155;
wire v_63156;
wire v_63157;
wire v_63158;
wire v_63159;
wire v_63160;
wire v_63161;
wire v_63162;
wire v_63163;
wire v_63164;
wire v_63165;
wire v_63166;
wire v_63167;
wire v_63168;
wire v_63169;
wire v_63170;
wire v_63171;
wire v_63172;
wire v_63173;
wire v_63174;
wire v_63175;
wire v_63176;
wire v_63177;
wire v_63178;
wire v_63179;
wire v_63180;
wire v_63181;
wire v_63182;
wire v_63183;
wire v_63184;
wire v_63185;
wire v_63186;
wire v_63187;
wire v_63188;
wire v_63189;
wire v_63190;
wire v_63191;
wire v_63192;
wire v_63193;
wire v_63194;
wire v_63195;
wire v_63196;
wire v_63197;
wire v_63198;
wire v_63199;
wire v_63200;
wire v_63201;
wire v_63202;
wire v_63203;
wire v_63204;
wire v_63205;
wire v_63206;
wire v_63207;
wire v_63208;
wire v_63209;
wire v_63210;
wire v_63211;
wire v_63212;
wire v_63213;
wire v_63214;
wire v_63215;
wire v_63216;
wire v_63217;
wire v_63218;
wire v_63219;
wire v_63220;
wire v_63221;
wire v_63222;
wire v_63223;
wire v_63224;
wire v_63225;
wire v_63226;
wire v_63227;
wire v_63228;
wire v_63229;
wire v_63230;
wire v_63231;
wire v_63232;
wire v_63233;
wire v_63234;
wire v_63235;
wire v_63236;
wire v_63237;
wire v_63238;
wire v_63239;
wire v_63240;
wire v_63241;
wire v_63242;
wire v_63243;
wire v_63244;
wire v_63245;
wire v_63246;
wire v_63247;
wire v_63248;
wire v_63249;
wire v_63250;
wire v_63251;
wire v_63252;
wire v_63253;
wire v_63254;
wire v_63255;
wire v_63256;
wire v_63257;
wire v_63258;
wire v_63259;
wire v_63261;
wire v_63262;
wire v_63263;
wire v_63264;
wire v_63265;
wire v_63266;
wire v_63267;
wire v_63268;
wire v_63269;
wire v_63270;
wire v_63271;
wire v_63272;
wire v_63273;
wire v_63274;
wire v_63275;
wire v_63276;
wire v_63277;
wire v_63278;
wire v_63279;
wire v_63280;
wire v_63281;
wire v_63282;
wire v_63283;
wire v_63284;
wire v_63285;
wire v_63286;
wire v_63287;
wire v_63288;
wire v_63289;
wire v_63290;
wire v_63291;
wire v_63292;
wire v_63293;
wire v_63294;
wire v_63295;
wire v_63296;
wire v_63297;
wire v_63298;
wire v_63299;
wire v_63300;
wire v_63301;
wire v_63302;
wire v_63303;
wire v_63304;
wire v_63305;
wire v_63306;
wire v_63307;
wire v_63308;
wire v_63309;
wire v_63310;
wire v_63311;
wire v_63312;
wire v_63313;
wire v_63314;
wire v_63315;
wire v_63316;
wire v_63317;
wire v_63318;
wire v_63319;
wire v_63320;
wire v_63321;
wire v_63322;
wire v_63323;
wire v_63324;
wire v_63325;
wire v_63326;
wire v_63327;
wire v_63328;
wire v_63329;
wire v_63330;
wire v_63331;
wire v_63332;
wire v_63333;
wire v_63334;
wire v_63335;
wire v_63336;
wire v_63337;
wire v_63338;
wire v_63339;
wire v_63340;
wire v_63341;
wire v_63342;
wire v_63343;
wire v_63344;
wire v_63345;
wire v_63346;
wire v_63347;
wire v_63348;
wire v_63349;
wire v_63350;
wire v_63351;
wire v_63352;
wire v_63353;
wire v_63354;
wire v_63355;
wire v_63356;
wire v_63357;
wire v_63358;
wire v_63359;
wire v_63360;
wire v_63361;
wire v_63362;
wire v_63363;
wire v_63364;
wire v_63365;
wire v_63366;
wire v_63367;
wire v_63368;
wire v_63369;
wire v_63370;
wire v_63371;
wire v_63372;
wire v_63373;
wire v_63374;
wire v_63375;
wire v_63376;
wire v_63377;
wire v_63378;
wire v_63379;
wire v_63380;
wire v_63381;
wire v_63382;
wire v_63383;
wire v_63384;
wire v_63385;
wire v_63386;
wire v_63387;
wire v_63388;
wire v_63389;
wire v_63390;
wire v_63391;
wire v_63392;
wire v_63393;
wire v_63394;
wire v_63395;
wire v_63396;
wire v_63397;
wire v_63398;
wire v_63399;
wire v_63400;
wire v_63401;
wire v_63402;
wire v_63403;
wire v_63404;
wire v_63405;
wire v_63406;
wire v_63407;
wire v_63408;
wire v_63409;
wire v_63410;
wire v_63411;
wire v_63412;
wire v_63413;
wire v_63414;
wire v_63415;
wire v_63416;
wire v_63417;
wire v_63418;
wire v_63419;
wire v_63420;
wire v_63421;
wire v_63422;
wire v_63423;
wire v_63424;
wire v_63425;
wire v_63426;
wire v_63427;
wire v_63428;
wire v_63429;
wire v_63430;
wire v_63431;
wire v_63432;
wire v_63433;
wire v_63434;
wire v_63435;
wire v_63436;
wire v_63437;
wire v_63438;
wire v_63439;
wire v_63440;
wire v_63441;
wire v_63442;
wire v_63443;
wire v_63444;
wire v_63445;
wire v_63446;
wire v_63447;
wire v_63448;
wire v_63449;
wire v_63450;
wire v_63451;
wire v_63452;
wire v_63453;
wire v_63454;
wire v_63455;
wire v_63456;
wire v_63457;
wire v_63458;
wire v_63459;
wire v_63460;
wire v_63461;
wire v_63462;
wire v_63463;
wire v_63464;
wire v_63465;
wire v_63466;
wire v_63467;
wire v_63468;
wire v_63469;
wire v_63470;
wire v_63471;
wire v_63472;
wire v_63473;
wire v_63474;
wire v_63475;
wire v_63476;
wire v_63477;
wire v_63478;
wire v_63479;
wire v_63480;
wire v_63481;
wire v_63482;
wire v_63483;
wire v_63484;
wire v_63485;
wire v_63486;
wire v_63487;
wire v_63488;
wire v_63489;
wire v_63490;
wire v_63491;
wire v_63492;
wire v_63493;
wire v_63494;
wire v_63495;
wire v_63496;
wire v_63497;
wire v_63498;
wire v_63499;
wire v_63500;
wire v_63501;
wire v_63502;
wire v_63504;
wire v_63505;
wire v_63506;
wire v_63507;
wire v_63508;
wire v_63509;
wire v_63510;
wire v_63511;
wire v_63512;
wire v_63513;
wire v_63514;
wire v_63515;
wire v_63516;
wire v_63517;
wire v_63518;
wire v_63519;
wire v_63520;
wire v_63521;
wire v_63522;
wire v_63523;
wire v_63524;
wire v_63525;
wire v_63526;
wire v_63527;
wire v_63528;
wire v_63529;
wire v_63530;
wire v_63531;
wire v_63532;
wire v_63533;
wire v_63534;
wire v_63535;
wire v_63536;
wire v_63537;
wire v_63538;
wire v_63539;
wire v_63540;
wire v_63541;
wire v_63542;
wire v_63543;
wire v_63544;
wire v_63545;
wire v_63546;
wire v_63547;
wire v_63548;
wire v_63549;
wire v_63550;
wire v_63551;
wire v_63552;
wire v_63553;
wire v_63554;
wire v_63555;
wire v_63556;
wire v_63557;
wire v_63558;
wire v_63559;
wire v_63560;
wire v_63561;
wire v_63562;
wire v_63563;
wire v_63564;
wire v_63565;
wire v_63566;
wire v_63567;
wire v_63568;
wire v_63569;
wire v_63570;
wire v_63571;
wire v_63572;
wire v_63573;
wire v_63574;
wire v_63575;
wire v_63576;
wire v_63577;
wire v_63578;
wire v_63579;
wire v_63580;
wire v_63581;
wire v_63582;
wire v_63583;
wire v_63584;
wire v_63585;
wire v_63586;
wire v_63587;
wire v_63588;
wire v_63589;
wire v_63590;
wire v_63591;
wire v_63592;
wire v_63593;
wire v_63594;
wire v_63595;
wire v_63596;
wire v_63597;
wire v_63598;
wire v_63599;
wire v_63600;
wire v_63601;
wire v_63602;
wire v_63603;
wire v_63604;
wire v_63605;
wire v_63606;
wire v_63607;
wire v_63608;
wire v_63609;
wire v_63610;
wire v_63611;
wire v_63612;
wire v_63613;
wire v_63614;
wire v_63615;
wire v_63616;
wire v_63617;
wire v_63618;
wire v_63619;
wire v_63620;
wire v_63621;
wire v_63622;
wire v_63623;
wire v_63624;
wire v_63625;
wire v_63626;
wire v_63627;
wire v_63628;
wire v_63629;
wire v_63630;
wire v_63631;
wire v_63632;
wire v_63633;
wire v_63634;
wire v_63635;
wire v_63636;
wire v_63637;
wire v_63638;
wire v_63639;
wire v_63640;
wire v_63641;
wire v_63642;
wire v_63643;
wire v_63644;
wire v_63645;
wire v_63646;
wire v_63647;
wire v_63648;
wire v_63649;
wire v_63650;
wire v_63651;
wire v_63652;
wire v_63653;
wire v_63654;
wire v_63655;
wire v_63656;
wire v_63657;
wire v_63658;
wire v_63659;
wire v_63660;
wire v_63661;
wire v_63662;
wire v_63663;
wire v_63664;
wire v_63665;
wire v_63666;
wire v_63667;
wire v_63668;
wire v_63669;
wire v_63670;
wire v_63671;
wire v_63672;
wire v_63673;
wire v_63674;
wire v_63675;
wire v_63676;
wire v_63677;
wire v_63678;
wire v_63679;
wire v_63680;
wire v_63681;
wire v_63682;
wire v_63683;
wire v_63684;
wire v_63685;
wire v_63686;
wire v_63687;
wire v_63688;
wire v_63689;
wire v_63690;
wire v_63691;
wire v_63692;
wire v_63693;
wire v_63694;
wire v_63695;
wire v_63696;
wire v_63697;
wire v_63698;
wire v_63699;
wire v_63700;
wire v_63701;
wire v_63702;
wire v_63703;
wire v_63704;
wire v_63705;
wire v_63706;
wire v_63707;
wire v_63708;
wire v_63709;
wire v_63710;
wire v_63711;
wire v_63712;
wire v_63713;
wire v_63714;
wire v_63715;
wire v_63716;
wire v_63717;
wire v_63718;
wire v_63719;
wire v_63720;
wire v_63721;
wire v_63722;
wire v_63723;
wire v_63724;
wire v_63725;
wire v_63726;
wire v_63727;
wire v_63728;
wire v_63729;
wire v_63730;
wire v_63731;
wire v_63732;
wire v_63733;
wire v_63734;
wire v_63735;
wire v_63736;
wire v_63737;
wire v_63738;
wire v_63739;
wire v_63740;
wire v_63741;
wire v_63742;
wire v_63743;
wire v_63744;
wire v_63745;
wire v_63747;
wire v_63748;
wire v_63749;
wire v_63750;
wire v_63751;
wire v_63752;
wire v_63753;
wire v_63754;
wire v_63755;
wire v_63756;
wire v_63757;
wire v_63758;
wire v_63759;
wire v_63760;
wire v_63761;
wire v_63762;
wire v_63763;
wire v_63764;
wire v_63765;
wire v_63766;
wire v_63767;
wire v_63768;
wire v_63769;
wire v_63770;
wire v_63771;
wire v_63772;
wire v_63773;
wire v_63774;
wire v_63775;
wire v_63776;
wire v_63777;
wire v_63778;
wire v_63779;
wire v_63780;
wire v_63781;
wire v_63782;
wire v_63783;
wire v_63784;
wire v_63785;
wire v_63786;
wire v_63787;
wire v_63788;
wire v_63789;
wire v_63790;
wire v_63791;
wire v_63792;
wire v_63793;
wire v_63794;
wire v_63795;
wire v_63796;
wire v_63797;
wire v_63798;
wire v_63799;
wire v_63800;
wire v_63801;
wire v_63802;
wire v_63803;
wire v_63804;
wire v_63805;
wire v_63806;
wire v_63807;
wire v_63808;
wire v_63809;
wire v_63810;
wire v_63811;
wire v_63812;
wire v_63813;
wire v_63814;
wire v_63815;
wire v_63816;
wire v_63817;
wire v_63818;
wire v_63819;
wire v_63820;
wire v_63821;
wire v_63822;
wire v_63823;
wire v_63824;
wire v_63825;
wire v_63826;
wire v_63827;
wire v_63828;
wire v_63829;
wire v_63830;
wire v_63831;
wire v_63832;
wire v_63833;
wire v_63834;
wire v_63835;
wire v_63836;
wire v_63837;
wire v_63838;
wire v_63839;
wire v_63840;
wire v_63841;
wire v_63842;
wire v_63843;
wire v_63844;
wire v_63845;
wire v_63846;
wire v_63847;
wire v_63848;
wire v_63849;
wire v_63850;
wire v_63851;
wire v_63852;
wire v_63853;
wire v_63854;
wire v_63855;
wire v_63856;
wire v_63857;
wire v_63858;
wire v_63859;
wire v_63860;
wire v_63861;
wire v_63862;
wire v_63863;
wire v_63864;
wire v_63865;
wire v_63866;
wire v_63867;
wire v_63868;
wire v_63869;
wire v_63870;
wire v_63871;
wire v_63872;
wire v_63873;
wire v_63874;
wire v_63875;
wire v_63876;
wire v_63877;
wire v_63878;
wire v_63879;
wire v_63880;
wire v_63881;
wire v_63882;
wire v_63883;
wire v_63884;
wire v_63885;
wire v_63886;
wire v_63887;
wire v_63888;
wire v_63889;
wire v_63890;
wire v_63891;
wire v_63892;
wire v_63893;
wire v_63894;
wire v_63895;
wire v_63896;
wire v_63897;
wire v_63898;
wire v_63899;
wire v_63900;
wire v_63901;
wire v_63902;
wire v_63903;
wire v_63904;
wire v_63905;
wire v_63906;
wire v_63907;
wire v_63908;
wire v_63909;
wire v_63910;
wire v_63911;
wire v_63912;
wire v_63913;
wire v_63914;
wire v_63915;
wire v_63916;
wire v_63917;
wire v_63918;
wire v_63919;
wire v_63920;
wire v_63921;
wire v_63922;
wire v_63923;
wire v_63924;
wire v_63925;
wire v_63926;
wire v_63927;
wire v_63928;
wire v_63929;
wire v_63930;
wire v_63931;
wire v_63932;
wire v_63933;
wire v_63934;
wire v_63935;
wire v_63936;
wire v_63937;
wire v_63938;
wire v_63939;
wire v_63940;
wire v_63941;
wire v_63942;
wire v_63943;
wire v_63944;
wire v_63945;
wire v_63946;
wire v_63947;
wire v_63948;
wire v_63949;
wire v_63950;
wire v_63951;
wire v_63952;
wire v_63953;
wire v_63954;
wire v_63955;
wire v_63956;
wire v_63957;
wire v_63958;
wire v_63959;
wire v_63960;
wire v_63961;
wire v_63962;
wire v_63963;
wire v_63964;
wire v_63965;
wire v_63966;
wire v_63967;
wire v_63968;
wire v_63969;
wire v_63970;
wire v_63971;
wire v_63972;
wire v_63973;
wire v_63974;
wire v_63975;
wire v_63976;
wire v_63977;
wire v_63978;
wire v_63979;
wire v_63980;
wire v_63981;
wire v_63982;
wire v_63983;
wire v_63984;
wire v_63985;
wire v_63986;
wire v_63987;
wire v_63988;
wire v_63990;
wire v_63991;
wire v_63992;
wire v_63993;
wire v_63994;
wire v_63995;
wire v_63996;
wire v_63997;
wire v_63998;
wire v_63999;
wire v_64000;
wire v_64001;
wire v_64002;
wire v_64003;
wire v_64004;
wire v_64005;
wire v_64006;
wire v_64007;
wire v_64008;
wire v_64009;
wire v_64010;
wire v_64011;
wire v_64012;
wire v_64013;
wire v_64014;
wire v_64015;
wire v_64016;
wire v_64017;
wire v_64018;
wire v_64019;
wire v_64020;
wire v_64021;
wire v_64022;
wire v_64023;
wire v_64024;
wire v_64025;
wire v_64026;
wire v_64027;
wire v_64028;
wire v_64029;
wire v_64030;
wire v_64031;
wire v_64032;
wire v_64033;
wire v_64034;
wire v_64035;
wire v_64036;
wire v_64037;
wire v_64038;
wire v_64039;
wire v_64040;
wire v_64041;
wire v_64042;
wire v_64043;
wire v_64044;
wire v_64045;
wire v_64046;
wire v_64047;
wire v_64048;
wire v_64049;
wire v_64050;
wire v_64051;
wire v_64052;
wire v_64053;
wire v_64054;
wire v_64055;
wire v_64056;
wire v_64057;
wire v_64058;
wire v_64059;
wire v_64060;
wire v_64061;
wire v_64062;
wire v_64063;
wire v_64064;
wire v_64065;
wire v_64066;
wire v_64067;
wire v_64068;
wire v_64069;
wire v_64070;
wire v_64071;
wire v_64072;
wire v_64073;
wire v_64074;
wire v_64075;
wire v_64076;
wire v_64077;
wire v_64078;
wire v_64079;
wire v_64080;
wire v_64081;
wire v_64082;
wire v_64083;
wire v_64084;
wire v_64085;
wire v_64086;
wire v_64087;
wire v_64088;
wire v_64089;
wire v_64090;
wire v_64091;
wire v_64092;
wire v_64093;
wire v_64094;
wire v_64095;
wire v_64096;
wire v_64097;
wire v_64098;
wire v_64099;
wire v_64100;
wire v_64101;
wire v_64102;
wire v_64103;
wire v_64104;
wire v_64105;
wire v_64106;
wire v_64107;
wire v_64108;
wire v_64109;
wire v_64110;
wire v_64111;
wire v_64112;
wire v_64113;
wire v_64114;
wire v_64115;
wire v_64116;
wire v_64117;
wire v_64118;
wire v_64119;
wire v_64120;
wire v_64121;
wire v_64122;
wire v_64123;
wire v_64124;
wire v_64125;
wire v_64126;
wire v_64127;
wire v_64128;
wire v_64129;
wire v_64130;
wire v_64131;
wire v_64132;
wire v_64133;
wire v_64134;
wire v_64135;
wire v_64136;
wire v_64137;
wire v_64138;
wire v_64139;
wire v_64140;
wire v_64141;
wire v_64142;
wire v_64143;
wire v_64144;
wire v_64145;
wire v_64146;
wire v_64147;
wire v_64148;
wire v_64149;
wire v_64150;
wire v_64151;
wire v_64152;
wire v_64153;
wire v_64154;
wire v_64155;
wire v_64156;
wire v_64157;
wire v_64158;
wire v_64159;
wire v_64160;
wire v_64161;
wire v_64162;
wire v_64163;
wire v_64164;
wire v_64165;
wire v_64166;
wire v_64167;
wire v_64168;
wire v_64169;
wire v_64170;
wire v_64171;
wire v_64172;
wire v_64173;
wire v_64174;
wire v_64175;
wire v_64176;
wire v_64177;
wire v_64178;
wire v_64179;
wire v_64180;
wire v_64181;
wire v_64182;
wire v_64183;
wire v_64184;
wire v_64185;
wire v_64186;
wire v_64187;
wire v_64188;
wire v_64189;
wire v_64190;
wire v_64191;
wire v_64192;
wire v_64193;
wire v_64194;
wire v_64195;
wire v_64196;
wire v_64197;
wire v_64198;
wire v_64199;
wire v_64200;
wire v_64201;
wire v_64202;
wire v_64203;
wire v_64204;
wire v_64205;
wire v_64206;
wire v_64207;
wire v_64208;
wire v_64209;
wire v_64210;
wire v_64211;
wire v_64212;
wire v_64213;
wire v_64214;
wire v_64215;
wire v_64216;
wire v_64217;
wire v_64218;
wire v_64219;
wire v_64220;
wire v_64221;
wire v_64222;
wire v_64223;
wire v_64224;
wire v_64225;
wire v_64226;
wire v_64227;
wire v_64228;
wire v_64229;
wire v_64230;
wire v_64231;
wire v_64233;
wire v_64234;
wire v_64235;
wire v_64236;
wire v_64237;
wire v_64238;
wire v_64239;
wire v_64240;
wire v_64241;
wire v_64242;
wire v_64243;
wire v_64244;
wire v_64245;
wire v_64246;
wire v_64247;
wire v_64248;
wire v_64249;
wire v_64250;
wire v_64251;
wire v_64252;
wire v_64253;
wire v_64254;
wire v_64255;
wire v_64256;
wire v_64257;
wire v_64258;
wire v_64259;
wire v_64260;
wire v_64261;
wire v_64262;
wire v_64263;
wire v_64264;
wire v_64265;
wire v_64266;
wire v_64267;
wire v_64268;
wire v_64269;
wire v_64270;
wire v_64271;
wire v_64272;
wire v_64273;
wire v_64274;
wire v_64275;
wire v_64276;
wire v_64277;
wire v_64278;
wire v_64279;
wire v_64280;
wire v_64281;
wire v_64282;
wire v_64283;
wire v_64284;
wire v_64285;
wire v_64286;
wire v_64287;
wire v_64288;
wire v_64289;
wire v_64290;
wire v_64291;
wire v_64292;
wire v_64293;
wire v_64294;
wire v_64295;
wire v_64296;
wire v_64297;
wire v_64298;
wire v_64299;
wire v_64300;
wire v_64301;
wire v_64302;
wire v_64303;
wire v_64304;
wire v_64305;
wire v_64306;
wire v_64307;
wire v_64308;
wire v_64309;
wire v_64310;
wire v_64311;
wire v_64312;
wire v_64313;
wire v_64314;
wire v_64315;
wire v_64316;
wire v_64317;
wire v_64318;
wire v_64319;
wire v_64320;
wire v_64321;
wire v_64322;
wire v_64323;
wire v_64324;
wire v_64325;
wire v_64326;
wire v_64327;
wire v_64328;
wire v_64329;
wire v_64330;
wire v_64331;
wire v_64332;
wire v_64333;
wire v_64334;
wire v_64335;
wire v_64336;
wire v_64337;
wire v_64338;
wire v_64339;
wire v_64340;
wire v_64341;
wire v_64342;
wire v_64343;
wire v_64344;
wire v_64345;
wire v_64346;
wire v_64347;
wire v_64348;
wire v_64349;
wire v_64350;
wire v_64351;
wire v_64352;
wire v_64353;
wire v_64354;
wire v_64355;
wire v_64356;
wire v_64357;
wire v_64358;
wire v_64359;
wire v_64360;
wire v_64361;
wire v_64362;
wire v_64363;
wire v_64364;
wire v_64365;
wire v_64366;
wire v_64367;
wire v_64368;
wire v_64369;
wire v_64370;
wire v_64371;
wire v_64372;
wire v_64373;
wire v_64374;
wire v_64375;
wire v_64376;
wire v_64377;
wire v_64378;
wire v_64379;
wire v_64380;
wire v_64381;
wire v_64382;
wire v_64383;
wire v_64384;
wire v_64385;
wire v_64386;
wire v_64387;
wire v_64388;
wire v_64389;
wire v_64390;
wire v_64391;
wire v_64392;
wire v_64393;
wire v_64394;
wire v_64395;
wire v_64396;
wire v_64397;
wire v_64398;
wire v_64399;
wire v_64400;
wire v_64401;
wire v_64402;
wire v_64403;
wire v_64404;
wire v_64405;
wire v_64406;
wire v_64407;
wire v_64408;
wire v_64409;
wire v_64410;
wire v_64411;
wire v_64412;
wire v_64413;
wire v_64414;
wire v_64415;
wire v_64416;
wire v_64417;
wire v_64418;
wire v_64419;
wire v_64420;
wire v_64421;
wire v_64422;
wire v_64423;
wire v_64424;
wire v_64425;
wire v_64426;
wire v_64427;
wire v_64428;
wire v_64429;
wire v_64430;
wire v_64431;
wire v_64432;
wire v_64433;
wire v_64434;
wire v_64435;
wire v_64436;
wire v_64437;
wire v_64438;
wire v_64439;
wire v_64440;
wire v_64441;
wire v_64442;
wire v_64443;
wire v_64444;
wire v_64445;
wire v_64446;
wire v_64447;
wire v_64448;
wire v_64449;
wire v_64450;
wire v_64451;
wire v_64452;
wire v_64453;
wire v_64454;
wire v_64455;
wire v_64456;
wire v_64457;
wire v_64458;
wire v_64459;
wire v_64460;
wire v_64461;
wire v_64462;
wire v_64463;
wire v_64464;
wire v_64465;
wire v_64466;
wire v_64467;
wire v_64468;
wire v_64469;
wire v_64470;
wire v_64471;
wire v_64472;
wire v_64473;
wire v_64474;
wire v_64476;
wire v_64477;
wire v_64478;
wire v_64479;
wire v_64480;
wire v_64481;
wire v_64482;
wire v_64483;
wire v_64484;
wire v_64485;
wire v_64486;
wire v_64487;
wire v_64488;
wire v_64489;
wire v_64490;
wire v_64491;
wire v_64492;
wire v_64493;
wire v_64494;
wire v_64495;
wire v_64496;
wire v_64497;
wire v_64498;
wire v_64499;
wire v_64500;
wire v_64501;
wire v_64502;
wire v_64503;
wire v_64504;
wire v_64505;
wire v_64506;
wire v_64507;
wire v_64508;
wire v_64509;
wire v_64510;
wire v_64511;
wire v_64512;
wire v_64513;
wire v_64514;
wire v_64515;
wire v_64516;
wire v_64517;
wire v_64518;
wire v_64519;
wire v_64520;
wire v_64521;
wire v_64522;
wire v_64523;
wire v_64524;
wire v_64525;
wire v_64526;
wire v_64527;
wire v_64528;
wire v_64529;
wire v_64530;
wire v_64531;
wire v_64532;
wire v_64533;
wire v_64534;
wire v_64535;
wire v_64536;
wire v_64537;
wire v_64538;
wire v_64539;
wire v_64540;
wire v_64541;
wire v_64542;
wire v_64543;
wire v_64544;
wire v_64545;
wire v_64546;
wire v_64547;
wire v_64548;
wire v_64549;
wire v_64550;
wire v_64551;
wire v_64552;
wire v_64553;
wire v_64554;
wire v_64555;
wire v_64556;
wire v_64557;
wire v_64558;
wire v_64559;
wire v_64560;
wire v_64561;
wire v_64562;
wire v_64563;
wire v_64564;
wire v_64565;
wire v_64566;
wire v_64567;
wire v_64568;
wire v_64569;
wire v_64570;
wire v_64571;
wire v_64572;
wire v_64573;
wire v_64574;
wire v_64575;
wire v_64576;
wire v_64577;
wire v_64578;
wire v_64579;
wire v_64580;
wire v_64581;
wire v_64582;
wire v_64583;
wire v_64584;
wire v_64585;
wire v_64586;
wire v_64587;
wire v_64588;
wire v_64589;
wire v_64590;
wire v_64591;
wire v_64592;
wire v_64593;
wire v_64594;
wire v_64595;
wire v_64596;
wire v_64597;
wire v_64598;
wire v_64599;
wire v_64600;
wire v_64601;
wire v_64602;
wire v_64603;
wire v_64604;
wire v_64605;
wire v_64606;
wire v_64607;
wire v_64608;
wire v_64609;
wire v_64610;
wire v_64611;
wire v_64612;
wire v_64613;
wire v_64614;
wire v_64615;
wire v_64616;
wire v_64617;
wire v_64618;
wire v_64619;
wire v_64620;
wire v_64621;
wire v_64622;
wire v_64623;
wire v_64624;
wire v_64625;
wire v_64626;
wire v_64627;
wire v_64628;
wire v_64629;
wire v_64630;
wire v_64631;
wire v_64632;
wire v_64633;
wire v_64634;
wire v_64635;
wire v_64636;
wire v_64637;
wire v_64638;
wire v_64639;
wire v_64640;
wire v_64641;
wire v_64642;
wire v_64643;
wire v_64644;
wire v_64645;
wire v_64646;
wire v_64647;
wire v_64648;
wire v_64649;
wire v_64650;
wire v_64651;
wire v_64652;
wire v_64653;
wire v_64654;
wire v_64655;
wire v_64656;
wire v_64657;
wire v_64658;
wire v_64659;
wire v_64660;
wire v_64661;
wire v_64662;
wire v_64663;
wire v_64664;
wire v_64665;
wire v_64666;
wire v_64667;
wire v_64668;
wire v_64669;
wire v_64670;
wire v_64671;
wire v_64672;
wire v_64673;
wire v_64674;
wire v_64675;
wire v_64676;
wire v_64677;
wire v_64678;
wire v_64679;
wire v_64680;
wire v_64681;
wire v_64682;
wire v_64683;
wire v_64684;
wire v_64685;
wire v_64686;
wire v_64687;
wire v_64688;
wire v_64689;
wire v_64690;
wire v_64691;
wire v_64692;
wire v_64693;
wire v_64694;
wire v_64695;
wire v_64696;
wire v_64697;
wire v_64698;
wire v_64699;
wire v_64700;
wire v_64701;
wire v_64702;
wire v_64703;
wire v_64704;
wire v_64705;
wire v_64706;
wire v_64707;
wire v_64708;
wire v_64709;
wire v_64710;
wire v_64711;
wire v_64712;
wire v_64713;
wire v_64714;
wire v_64715;
wire v_64716;
wire v_64717;
wire v_64719;
wire v_64720;
wire v_64721;
wire v_64722;
wire v_64723;
wire v_64724;
wire v_64725;
wire v_64726;
wire v_64727;
wire v_64728;
wire v_64729;
wire v_64730;
wire v_64731;
wire v_64732;
wire v_64733;
wire v_64734;
wire v_64735;
wire v_64736;
wire v_64737;
wire v_64738;
wire v_64739;
wire v_64740;
wire v_64741;
wire v_64742;
wire v_64743;
wire v_64744;
wire v_64745;
wire v_64746;
wire v_64747;
wire v_64748;
wire v_64749;
wire v_64750;
wire v_64751;
wire v_64752;
wire v_64753;
wire v_64754;
wire v_64755;
wire v_64756;
wire v_64757;
wire v_64758;
wire v_64759;
wire v_64760;
wire v_64761;
wire v_64762;
wire v_64763;
wire v_64764;
wire v_64765;
wire v_64766;
wire v_64767;
wire v_64768;
wire v_64769;
wire v_64770;
wire v_64771;
wire v_64772;
wire v_64773;
wire v_64774;
wire v_64775;
wire v_64776;
wire v_64777;
wire v_64778;
wire v_64779;
wire v_64780;
wire v_64781;
wire v_64782;
wire v_64783;
wire v_64784;
wire v_64785;
wire v_64786;
wire v_64787;
wire v_64788;
wire v_64789;
wire v_64790;
wire v_64791;
wire v_64792;
wire v_64793;
wire v_64794;
wire v_64795;
wire v_64796;
wire v_64797;
wire v_64798;
wire v_64799;
wire v_64800;
wire v_64801;
wire v_64802;
wire v_64803;
wire v_64804;
wire v_64805;
wire v_64806;
wire v_64807;
wire v_64808;
wire v_64809;
wire v_64810;
wire v_64811;
wire v_64812;
wire v_64813;
wire v_64814;
wire v_64815;
wire v_64816;
wire v_64817;
wire v_64818;
wire v_64819;
wire v_64820;
wire v_64821;
wire v_64822;
wire v_64823;
wire v_64824;
wire v_64825;
wire v_64826;
wire v_64827;
wire v_64828;
wire v_64829;
wire v_64830;
wire v_64831;
wire v_64832;
wire v_64833;
wire v_64834;
wire v_64835;
wire v_64836;
wire v_64837;
wire v_64838;
wire v_64839;
wire v_64840;
wire v_64841;
wire v_64842;
wire v_64843;
wire v_64844;
wire v_64845;
wire v_64846;
wire v_64847;
wire v_64848;
wire v_64849;
wire v_64850;
wire v_64851;
wire v_64852;
wire v_64853;
wire v_64854;
wire v_64855;
wire v_64856;
wire v_64857;
wire v_64858;
wire v_64859;
wire v_64860;
wire v_64861;
wire v_64862;
wire v_64863;
wire v_64864;
wire v_64865;
wire v_64866;
wire v_64867;
wire v_64868;
wire v_64869;
wire v_64870;
wire v_64871;
wire v_64872;
wire v_64873;
wire v_64874;
wire v_64875;
wire v_64876;
wire v_64877;
wire v_64878;
wire v_64879;
wire v_64880;
wire v_64881;
wire v_64882;
wire v_64883;
wire v_64884;
wire v_64885;
wire v_64886;
wire v_64887;
wire v_64888;
wire v_64889;
wire v_64890;
wire v_64891;
wire v_64892;
wire v_64893;
wire v_64894;
wire v_64895;
wire v_64896;
wire v_64897;
wire v_64898;
wire v_64899;
wire v_64900;
wire v_64901;
wire v_64902;
wire v_64903;
wire v_64904;
wire v_64905;
wire v_64906;
wire v_64907;
wire v_64908;
wire v_64909;
wire v_64910;
wire v_64911;
wire v_64912;
wire v_64913;
wire v_64914;
wire v_64915;
wire v_64916;
wire v_64917;
wire v_64918;
wire v_64919;
wire v_64920;
wire v_64921;
wire v_64922;
wire v_64923;
wire v_64924;
wire v_64925;
wire v_64926;
wire v_64927;
wire v_64928;
wire v_64929;
wire v_64930;
wire v_64931;
wire v_64932;
wire v_64933;
wire v_64934;
wire v_64935;
wire v_64936;
wire v_64937;
wire v_64938;
wire v_64939;
wire v_64940;
wire v_64941;
wire v_64942;
wire v_64943;
wire v_64944;
wire v_64945;
wire v_64946;
wire v_64947;
wire v_64948;
wire v_64949;
wire v_64950;
wire v_64951;
wire v_64952;
wire v_64953;
wire v_64954;
wire v_64955;
wire v_64956;
wire v_64957;
wire v_64958;
wire v_64959;
wire v_64960;
wire v_64962;
wire v_64963;
wire v_64964;
wire v_64965;
wire v_64966;
wire v_64967;
wire v_64968;
wire v_64969;
wire v_64970;
wire v_64971;
wire v_64972;
wire v_64973;
wire v_64974;
wire v_64975;
wire v_64976;
wire v_64977;
wire v_64978;
wire v_64979;
wire v_64980;
wire v_64981;
wire v_64982;
wire v_64983;
wire v_64984;
wire v_64985;
wire v_64986;
wire v_64987;
wire v_64988;
wire v_64989;
wire v_64990;
wire v_64991;
wire v_64992;
wire v_64993;
wire v_64994;
wire v_64995;
wire v_64996;
wire v_64997;
wire v_64998;
wire v_64999;
wire v_65000;
wire v_65001;
wire v_65002;
wire v_65003;
wire v_65004;
wire v_65005;
wire v_65006;
wire v_65007;
wire v_65008;
wire v_65009;
wire v_65010;
wire v_65011;
wire v_65012;
wire v_65013;
wire v_65014;
wire v_65015;
wire v_65016;
wire v_65017;
wire v_65018;
wire v_65019;
wire v_65020;
wire v_65021;
wire v_65022;
wire v_65023;
wire v_65024;
wire v_65025;
wire v_65026;
wire v_65027;
wire v_65028;
wire v_65029;
wire v_65030;
wire v_65031;
wire v_65032;
wire v_65033;
wire v_65034;
wire v_65035;
wire v_65036;
wire v_65037;
wire v_65038;
wire v_65039;
wire v_65040;
wire v_65041;
wire v_65042;
wire v_65043;
wire v_65044;
wire v_65045;
wire v_65046;
wire v_65047;
wire v_65048;
wire v_65049;
wire v_65050;
wire v_65051;
wire v_65052;
wire v_65053;
wire v_65054;
wire v_65055;
wire v_65056;
wire v_65057;
wire v_65058;
wire v_65059;
wire v_65060;
wire v_65061;
wire v_65062;
wire v_65063;
wire v_65064;
wire v_65065;
wire v_65066;
wire v_65067;
wire v_65068;
wire v_65069;
wire v_65070;
wire v_65071;
wire v_65072;
wire v_65073;
wire v_65074;
wire v_65075;
wire v_65076;
wire v_65077;
wire v_65078;
wire v_65079;
wire v_65080;
wire v_65081;
wire v_65082;
wire v_65083;
wire v_65084;
wire v_65085;
wire v_65086;
wire v_65087;
wire v_65088;
wire v_65089;
wire v_65090;
wire v_65091;
wire v_65092;
wire v_65093;
wire v_65094;
wire v_65095;
wire v_65096;
wire v_65097;
wire v_65098;
wire v_65099;
wire v_65100;
wire v_65101;
wire v_65102;
wire v_65103;
wire v_65104;
wire v_65105;
wire v_65106;
wire v_65107;
wire v_65108;
wire v_65109;
wire v_65110;
wire v_65111;
wire v_65112;
wire v_65113;
wire v_65114;
wire v_65115;
wire v_65116;
wire v_65117;
wire v_65118;
wire v_65119;
wire v_65120;
wire v_65121;
wire v_65122;
wire v_65123;
wire v_65124;
wire v_65125;
wire v_65126;
wire v_65127;
wire v_65128;
wire v_65129;
wire v_65130;
wire v_65131;
wire v_65132;
wire v_65133;
wire v_65134;
wire v_65135;
wire v_65136;
wire v_65137;
wire v_65138;
wire v_65139;
wire v_65140;
wire v_65141;
wire v_65142;
wire v_65143;
wire v_65144;
wire v_65145;
wire v_65146;
wire v_65147;
wire v_65148;
wire v_65149;
wire v_65150;
wire v_65151;
wire v_65152;
wire v_65153;
wire v_65154;
wire v_65155;
wire v_65156;
wire v_65157;
wire v_65158;
wire v_65159;
wire v_65160;
wire v_65161;
wire v_65162;
wire v_65163;
wire v_65164;
wire v_65165;
wire v_65166;
wire v_65167;
wire v_65168;
wire v_65169;
wire v_65170;
wire v_65171;
wire v_65172;
wire v_65173;
wire v_65174;
wire v_65175;
wire v_65176;
wire v_65177;
wire v_65178;
wire v_65179;
wire v_65180;
wire v_65181;
wire v_65182;
wire v_65183;
wire v_65184;
wire v_65185;
wire v_65186;
wire v_65187;
wire v_65188;
wire v_65189;
wire v_65190;
wire v_65191;
wire v_65192;
wire v_65193;
wire v_65194;
wire v_65195;
wire v_65196;
wire v_65197;
wire v_65198;
wire v_65199;
wire v_65200;
wire v_65201;
wire v_65202;
wire v_65203;
wire v_65205;
wire v_65206;
wire v_65207;
wire v_65208;
wire v_65209;
wire v_65210;
wire v_65211;
wire v_65212;
wire v_65213;
wire v_65214;
wire v_65215;
wire v_65216;
wire v_65217;
wire v_65218;
wire v_65219;
wire v_65220;
wire v_65221;
wire v_65222;
wire v_65223;
wire v_65224;
wire v_65225;
wire v_65226;
wire v_65227;
wire v_65228;
wire v_65229;
wire v_65230;
wire v_65231;
wire v_65232;
wire v_65233;
wire v_65234;
wire v_65235;
wire v_65236;
wire v_65237;
wire v_65238;
wire v_65239;
wire v_65240;
wire v_65241;
wire v_65242;
wire v_65243;
wire v_65244;
wire v_65245;
wire v_65246;
wire v_65247;
wire v_65248;
wire v_65249;
wire v_65250;
wire v_65251;
wire v_65252;
wire v_65253;
wire v_65254;
wire v_65255;
wire v_65256;
wire v_65257;
wire v_65258;
wire v_65259;
wire v_65260;
wire v_65261;
wire v_65262;
wire v_65263;
wire v_65264;
wire v_65265;
wire v_65266;
wire v_65267;
wire v_65268;
wire v_65269;
wire v_65270;
wire v_65271;
wire v_65272;
wire v_65273;
wire v_65274;
wire v_65275;
wire v_65276;
wire v_65277;
wire v_65278;
wire v_65279;
wire v_65280;
wire v_65281;
wire v_65282;
wire v_65283;
wire v_65284;
wire v_65285;
wire v_65286;
wire v_65287;
wire v_65288;
wire v_65289;
wire v_65290;
wire v_65291;
wire v_65292;
wire v_65293;
wire v_65294;
wire v_65295;
wire v_65296;
wire v_65297;
wire v_65298;
wire v_65299;
wire v_65300;
wire v_65301;
wire v_65302;
wire v_65303;
wire v_65304;
wire v_65305;
wire v_65306;
wire v_65307;
wire v_65308;
wire v_65309;
wire v_65310;
wire v_65311;
wire v_65312;
wire v_65313;
wire v_65314;
wire v_65315;
wire v_65316;
wire v_65317;
wire v_65318;
wire v_65319;
wire v_65320;
wire v_65321;
wire v_65322;
wire v_65323;
wire v_65324;
wire v_65325;
wire v_65326;
wire v_65327;
wire v_65328;
wire v_65329;
wire v_65330;
wire v_65331;
wire v_65332;
wire v_65333;
wire v_65334;
wire v_65335;
wire v_65336;
wire v_65337;
wire v_65338;
wire v_65339;
wire v_65340;
wire v_65341;
wire v_65342;
wire v_65343;
wire v_65344;
wire v_65345;
wire v_65346;
wire v_65347;
wire v_65348;
wire v_65349;
wire v_65350;
wire v_65351;
wire v_65352;
wire v_65353;
wire v_65354;
wire v_65355;
wire v_65356;
wire v_65357;
wire v_65358;
wire v_65359;
wire v_65360;
wire v_65361;
wire v_65362;
wire v_65363;
wire v_65364;
wire v_65365;
wire v_65366;
wire v_65367;
wire v_65368;
wire v_65369;
wire v_65370;
wire v_65371;
wire v_65372;
wire v_65373;
wire v_65374;
wire v_65375;
wire v_65376;
wire v_65377;
wire v_65378;
wire v_65379;
wire v_65380;
wire v_65381;
wire v_65382;
wire v_65383;
wire v_65384;
wire v_65385;
wire v_65386;
wire v_65387;
wire v_65388;
wire v_65389;
wire v_65390;
wire v_65391;
wire v_65392;
wire v_65393;
wire v_65394;
wire v_65395;
wire v_65396;
wire v_65397;
wire v_65398;
wire v_65399;
wire v_65400;
wire v_65401;
wire v_65402;
wire v_65403;
wire v_65404;
wire v_65405;
wire v_65406;
wire v_65407;
wire v_65408;
wire v_65409;
wire v_65410;
wire v_65411;
wire v_65412;
wire v_65413;
wire v_65414;
wire v_65415;
wire v_65416;
wire v_65417;
wire v_65418;
wire v_65419;
wire v_65420;
wire v_65421;
wire v_65422;
wire v_65423;
wire v_65424;
wire v_65425;
wire v_65426;
wire v_65427;
wire v_65428;
wire v_65429;
wire v_65430;
wire v_65431;
wire v_65432;
wire v_65433;
wire v_65434;
wire v_65435;
wire v_65436;
wire v_65437;
wire v_65438;
wire v_65439;
wire v_65440;
wire v_65441;
wire v_65442;
wire v_65443;
wire v_65444;
wire v_65445;
wire v_65446;
wire v_65448;
wire v_65449;
wire v_65450;
wire v_65451;
wire v_65452;
wire v_65453;
wire v_65454;
wire v_65455;
wire v_65456;
wire v_65457;
wire v_65458;
wire v_65459;
wire v_65460;
wire v_65461;
wire v_65462;
wire v_65463;
wire v_65464;
wire v_65465;
wire v_65466;
wire v_65467;
wire v_65468;
wire v_65469;
wire v_65470;
wire v_65471;
wire v_65472;
wire v_65473;
wire v_65474;
wire v_65475;
wire v_65476;
wire v_65477;
wire v_65478;
wire v_65479;
wire v_65480;
wire v_65481;
wire v_65482;
wire v_65483;
wire v_65484;
wire v_65485;
wire v_65486;
wire v_65487;
wire v_65488;
wire v_65489;
wire v_65490;
wire v_65491;
wire v_65492;
wire v_65493;
wire v_65494;
wire v_65495;
wire v_65496;
wire v_65497;
wire v_65498;
wire v_65499;
wire v_65500;
wire v_65501;
wire v_65502;
wire v_65503;
wire v_65504;
wire v_65505;
wire v_65506;
wire v_65507;
wire v_65508;
wire v_65509;
wire v_65510;
wire v_65511;
wire v_65512;
wire v_65513;
wire v_65514;
wire v_65515;
wire v_65516;
wire v_65517;
wire v_65518;
wire v_65519;
wire v_65520;
wire v_65521;
wire v_65522;
wire v_65523;
wire v_65524;
wire v_65525;
wire v_65526;
wire v_65527;
wire v_65528;
wire v_65529;
wire v_65530;
wire v_65531;
wire v_65532;
wire v_65533;
wire v_65534;
wire v_65535;
wire v_65536;
wire v_65537;
wire v_65538;
wire v_65539;
wire v_65540;
wire v_65541;
wire v_65542;
wire v_65543;
wire v_65544;
wire v_65545;
wire v_65546;
wire v_65547;
wire v_65548;
wire v_65549;
wire v_65550;
wire v_65551;
wire v_65552;
wire v_65553;
wire v_65554;
wire v_65555;
wire v_65556;
wire v_65557;
wire v_65558;
wire v_65559;
wire v_65560;
wire v_65561;
wire v_65562;
wire v_65563;
wire v_65564;
wire v_65565;
wire v_65566;
wire v_65567;
wire v_65568;
wire v_65569;
wire v_65570;
wire v_65571;
wire v_65572;
wire v_65573;
wire v_65574;
wire v_65575;
wire v_65576;
wire v_65577;
wire v_65578;
wire v_65579;
wire v_65580;
wire v_65581;
wire v_65582;
wire v_65583;
wire v_65584;
wire v_65585;
wire v_65586;
wire v_65587;
wire v_65588;
wire v_65589;
wire v_65590;
wire v_65591;
wire v_65592;
wire v_65593;
wire v_65594;
wire v_65595;
wire v_65596;
wire v_65597;
wire v_65598;
wire v_65599;
wire v_65600;
wire v_65601;
wire v_65602;
wire v_65603;
wire v_65604;
wire v_65605;
wire v_65606;
wire v_65607;
wire v_65608;
wire v_65609;
wire v_65610;
wire v_65611;
wire v_65612;
wire v_65613;
wire v_65614;
wire v_65615;
wire v_65616;
wire v_65617;
wire v_65618;
wire v_65619;
wire v_65620;
wire v_65621;
wire v_65622;
wire v_65623;
wire v_65624;
wire v_65625;
wire v_65626;
wire v_65627;
wire v_65628;
wire v_65629;
wire v_65630;
wire v_65631;
wire v_65632;
wire v_65633;
wire v_65634;
wire v_65635;
wire v_65636;
wire v_65637;
wire v_65638;
wire v_65639;
wire v_65640;
wire v_65641;
wire v_65642;
wire v_65643;
wire v_65644;
wire v_65645;
wire v_65646;
wire v_65647;
wire v_65648;
wire v_65649;
wire v_65650;
wire v_65651;
wire v_65652;
wire v_65653;
wire v_65654;
wire v_65655;
wire v_65656;
wire v_65657;
wire v_65658;
wire v_65659;
wire v_65660;
wire v_65661;
wire v_65662;
wire v_65663;
wire v_65664;
wire v_65665;
wire v_65666;
wire v_65667;
wire v_65668;
wire v_65669;
wire v_65670;
wire v_65671;
wire v_65672;
wire v_65673;
wire v_65674;
wire v_65675;
wire v_65676;
wire v_65677;
wire v_65678;
wire v_65679;
wire v_65680;
wire v_65681;
wire v_65682;
wire v_65683;
wire v_65684;
wire v_65685;
wire v_65686;
wire v_65687;
wire v_65688;
wire v_65689;
wire v_65691;
wire v_65692;
wire v_65693;
wire v_65694;
wire v_65695;
wire v_65696;
wire v_65697;
wire v_65698;
wire v_65699;
wire v_65700;
wire v_65701;
wire v_65702;
wire v_65703;
wire v_65704;
wire v_65705;
wire v_65706;
wire v_65707;
wire v_65708;
wire v_65709;
wire v_65710;
wire v_65711;
wire v_65712;
wire v_65713;
wire v_65714;
wire v_65715;
wire v_65716;
wire v_65717;
wire v_65718;
wire v_65719;
wire v_65720;
wire v_65721;
wire v_65722;
wire v_65723;
wire v_65724;
wire v_65725;
wire v_65726;
wire v_65727;
wire v_65728;
wire v_65729;
wire v_65730;
wire v_65731;
wire v_65732;
wire v_65733;
wire v_65734;
wire v_65735;
wire v_65736;
wire v_65737;
wire v_65738;
wire v_65739;
wire v_65740;
wire v_65741;
wire v_65742;
wire v_65743;
wire v_65744;
wire v_65745;
wire v_65746;
wire v_65747;
wire v_65748;
wire v_65749;
wire v_65750;
wire v_65751;
wire v_65752;
wire v_65753;
wire v_65754;
wire v_65755;
wire v_65756;
wire v_65757;
wire v_65758;
wire v_65759;
wire v_65760;
wire v_65761;
wire v_65762;
wire v_65763;
wire v_65764;
wire v_65765;
wire v_65766;
wire v_65767;
wire v_65768;
wire v_65769;
wire v_65770;
wire v_65771;
wire v_65772;
wire v_65773;
wire v_65774;
wire v_65775;
wire v_65776;
wire v_65777;
wire v_65778;
wire v_65779;
wire v_65780;
wire v_65781;
wire v_65782;
wire v_65783;
wire v_65784;
wire v_65785;
wire v_65786;
wire v_65787;
wire v_65788;
wire v_65789;
wire v_65790;
wire v_65791;
wire v_65792;
wire v_65793;
wire v_65794;
wire v_65795;
wire v_65796;
wire v_65797;
wire v_65798;
wire v_65799;
wire v_65800;
wire v_65801;
wire v_65802;
wire v_65803;
wire v_65804;
wire v_65805;
wire v_65806;
wire v_65807;
wire v_65808;
wire v_65809;
wire v_65810;
wire v_65811;
wire v_65812;
wire v_65813;
wire v_65814;
wire v_65815;
wire v_65816;
wire v_65817;
wire v_65818;
wire v_65819;
wire v_65820;
wire v_65821;
wire v_65822;
wire v_65823;
wire v_65824;
wire v_65825;
wire v_65826;
wire v_65827;
wire v_65828;
wire v_65829;
wire v_65830;
wire v_65831;
wire v_65832;
wire v_65833;
wire v_65834;
wire v_65835;
wire v_65836;
wire v_65837;
wire v_65838;
wire v_65839;
wire v_65840;
wire v_65841;
wire v_65842;
wire v_65843;
wire v_65844;
wire v_65845;
wire v_65846;
wire v_65847;
wire v_65848;
wire v_65849;
wire v_65850;
wire v_65851;
wire v_65852;
wire v_65853;
wire v_65854;
wire v_65855;
wire v_65856;
wire v_65857;
wire v_65858;
wire v_65859;
wire v_65860;
wire v_65861;
wire v_65862;
wire v_65863;
wire v_65864;
wire v_65865;
wire v_65866;
wire v_65867;
wire v_65868;
wire v_65869;
wire v_65870;
wire v_65871;
wire v_65872;
wire v_65873;
wire v_65874;
wire v_65875;
wire v_65876;
wire v_65877;
wire v_65878;
wire v_65879;
wire v_65880;
wire v_65881;
wire v_65882;
wire v_65883;
wire v_65884;
wire v_65885;
wire v_65886;
wire v_65887;
wire v_65888;
wire v_65889;
wire v_65890;
wire v_65891;
wire v_65892;
wire v_65893;
wire v_65894;
wire v_65895;
wire v_65896;
wire v_65897;
wire v_65898;
wire v_65899;
wire v_65900;
wire v_65901;
wire v_65902;
wire v_65903;
wire v_65904;
wire v_65905;
wire v_65906;
wire v_65907;
wire v_65908;
wire v_65909;
wire v_65910;
wire v_65911;
wire v_65912;
wire v_65913;
wire v_65914;
wire v_65915;
wire v_65916;
wire v_65917;
wire v_65918;
wire v_65919;
wire v_65920;
wire v_65921;
wire v_65922;
wire v_65923;
wire v_65924;
wire v_65925;
wire v_65926;
wire v_65927;
wire v_65928;
wire v_65929;
wire v_65930;
wire v_65931;
wire v_65932;
wire v_65934;
wire v_65935;
wire v_65936;
wire v_65937;
wire v_65938;
wire v_65939;
wire v_65940;
wire v_65941;
wire v_65942;
wire v_65943;
wire v_65944;
wire v_65945;
wire v_65946;
wire v_65947;
wire v_65948;
wire v_65949;
wire v_65950;
wire v_65951;
wire v_65952;
wire v_65953;
wire v_65954;
wire v_65955;
wire v_65956;
wire v_65957;
wire v_65958;
wire v_65959;
wire v_65960;
wire v_65961;
wire v_65962;
wire v_65963;
wire v_65964;
wire v_65965;
wire v_65966;
wire v_65967;
wire v_65968;
wire v_65969;
wire v_65970;
wire v_65971;
wire v_65972;
wire v_65973;
wire v_65974;
wire v_65975;
wire v_65976;
wire v_65977;
wire v_65978;
wire v_65979;
wire v_65980;
wire v_65981;
wire v_65982;
wire v_65983;
wire v_65984;
wire v_65985;
wire v_65986;
wire v_65987;
wire v_65988;
wire v_65989;
wire v_65990;
wire v_65991;
wire v_65992;
wire v_65993;
wire v_65994;
wire v_65995;
wire v_65996;
wire v_65997;
wire v_65998;
wire v_65999;
wire v_66000;
wire v_66001;
wire v_66002;
wire v_66003;
wire v_66004;
wire v_66005;
wire v_66006;
wire v_66007;
wire v_66008;
wire v_66009;
wire v_66010;
wire v_66011;
wire v_66012;
wire v_66013;
wire v_66014;
wire v_66015;
wire v_66016;
wire v_66017;
wire v_66018;
wire v_66019;
wire v_66020;
wire v_66021;
wire v_66022;
wire v_66023;
wire v_66024;
wire v_66025;
wire v_66026;
wire v_66027;
wire v_66028;
wire v_66029;
wire v_66030;
wire v_66031;
wire v_66032;
wire v_66033;
wire v_66034;
wire v_66035;
wire v_66036;
wire v_66037;
wire v_66038;
wire v_66039;
wire v_66040;
wire v_66041;
wire v_66042;
wire v_66043;
wire v_66044;
wire v_66045;
wire v_66046;
wire v_66047;
wire v_66048;
wire v_66049;
wire v_66050;
wire v_66051;
wire v_66052;
wire v_66053;
wire v_66054;
wire v_66055;
wire v_66056;
wire v_66057;
wire v_66058;
wire v_66059;
wire v_66060;
wire v_66061;
wire v_66062;
wire v_66063;
wire v_66064;
wire v_66065;
wire v_66066;
wire v_66067;
wire v_66068;
wire v_66069;
wire v_66070;
wire v_66071;
wire v_66072;
wire v_66073;
wire v_66074;
wire v_66075;
wire v_66076;
wire v_66077;
wire v_66078;
wire v_66079;
wire v_66080;
wire v_66081;
wire v_66082;
wire v_66083;
wire v_66084;
wire v_66085;
wire v_66086;
wire v_66087;
wire v_66088;
wire v_66089;
wire v_66090;
wire v_66091;
wire v_66092;
wire v_66093;
wire v_66094;
wire v_66095;
wire v_66096;
wire v_66097;
wire v_66098;
wire v_66099;
wire v_66100;
wire v_66101;
wire v_66102;
wire v_66103;
wire v_66104;
wire v_66105;
wire v_66106;
wire v_66107;
wire v_66108;
wire v_66109;
wire v_66110;
wire v_66111;
wire v_66112;
wire v_66113;
wire v_66114;
wire v_66115;
wire v_66116;
wire v_66117;
wire v_66118;
wire v_66119;
wire v_66120;
wire v_66121;
wire v_66122;
wire v_66123;
wire v_66124;
wire v_66125;
wire v_66126;
wire v_66127;
wire v_66128;
wire v_66129;
wire v_66130;
wire v_66131;
wire v_66132;
wire v_66133;
wire v_66134;
wire v_66135;
wire v_66136;
wire v_66137;
wire v_66138;
wire v_66139;
wire v_66140;
wire v_66141;
wire v_66142;
wire v_66143;
wire v_66144;
wire v_66145;
wire v_66146;
wire v_66147;
wire v_66148;
wire v_66149;
wire v_66150;
wire v_66151;
wire v_66152;
wire v_66153;
wire v_66154;
wire v_66155;
wire v_66156;
wire v_66157;
wire v_66158;
wire v_66159;
wire v_66160;
wire v_66161;
wire v_66162;
wire v_66163;
wire v_66164;
wire v_66165;
wire v_66166;
wire v_66167;
wire v_66168;
wire v_66169;
wire v_66170;
wire v_66171;
wire v_66172;
wire v_66173;
wire v_66174;
wire v_66175;
wire v_66177;
wire v_66178;
wire v_66179;
wire v_66180;
wire v_66181;
wire v_66182;
wire v_66183;
wire v_66184;
wire v_66185;
wire v_66186;
wire v_66187;
wire v_66188;
wire v_66189;
wire v_66190;
wire v_66191;
wire v_66192;
wire v_66193;
wire v_66194;
wire v_66195;
wire v_66196;
wire v_66197;
wire v_66198;
wire v_66199;
wire v_66200;
wire v_66201;
wire v_66202;
wire v_66203;
wire v_66204;
wire v_66205;
wire v_66206;
wire v_66207;
wire v_66208;
wire v_66209;
wire v_66210;
wire v_66211;
wire v_66212;
wire v_66213;
wire v_66214;
wire v_66215;
wire v_66216;
wire v_66217;
wire v_66218;
wire v_66219;
wire v_66220;
wire v_66221;
wire v_66222;
wire v_66223;
wire v_66224;
wire v_66225;
wire v_66226;
wire v_66227;
wire v_66228;
wire v_66229;
wire v_66230;
wire v_66231;
wire v_66232;
wire v_66233;
wire v_66234;
wire v_66235;
wire v_66236;
wire v_66237;
wire v_66238;
wire v_66239;
wire v_66240;
wire v_66241;
wire v_66242;
wire v_66243;
wire v_66244;
wire v_66245;
wire v_66246;
wire v_66247;
wire v_66248;
wire v_66249;
wire v_66250;
wire v_66251;
wire v_66252;
wire v_66253;
wire v_66254;
wire v_66255;
wire v_66256;
wire v_66257;
wire v_66258;
wire v_66259;
wire v_66260;
wire v_66261;
wire v_66262;
wire v_66263;
wire v_66264;
wire v_66265;
wire v_66266;
wire v_66267;
wire v_66268;
wire v_66269;
wire v_66270;
wire v_66271;
wire v_66272;
wire v_66273;
wire v_66274;
wire v_66275;
wire v_66276;
wire v_66277;
wire v_66278;
wire v_66279;
wire v_66280;
wire v_66281;
wire v_66282;
wire v_66283;
wire v_66284;
wire v_66285;
wire v_66286;
wire v_66287;
wire v_66288;
wire v_66289;
wire v_66290;
wire v_66291;
wire v_66292;
wire v_66293;
wire v_66294;
wire v_66295;
wire v_66296;
wire v_66297;
wire v_66298;
wire v_66299;
wire v_66300;
wire v_66301;
wire v_66302;
wire v_66303;
wire v_66304;
wire v_66305;
wire v_66306;
wire v_66307;
wire v_66308;
wire v_66309;
wire v_66310;
wire v_66311;
wire v_66312;
wire v_66313;
wire v_66314;
wire v_66315;
wire v_66316;
wire v_66317;
wire v_66318;
wire v_66319;
wire v_66320;
wire v_66321;
wire v_66322;
wire v_66323;
wire v_66324;
wire v_66325;
wire v_66326;
wire v_66327;
wire v_66328;
wire v_66329;
wire v_66330;
wire v_66331;
wire v_66332;
wire v_66333;
wire v_66334;
wire v_66335;
wire v_66336;
wire v_66337;
wire v_66338;
wire v_66339;
wire v_66340;
wire v_66341;
wire v_66342;
wire v_66343;
wire v_66344;
wire v_66345;
wire v_66346;
wire v_66347;
wire v_66348;
wire v_66349;
wire v_66350;
wire v_66351;
wire v_66352;
wire v_66353;
wire v_66354;
wire v_66355;
wire v_66356;
wire v_66357;
wire v_66358;
wire v_66359;
wire v_66360;
wire v_66361;
wire v_66362;
wire v_66363;
wire v_66364;
wire v_66365;
wire v_66366;
wire v_66367;
wire v_66368;
wire v_66369;
wire v_66370;
wire v_66371;
wire v_66372;
wire v_66373;
wire v_66374;
wire v_66375;
wire v_66376;
wire v_66377;
wire v_66378;
wire v_66379;
wire v_66380;
wire v_66381;
wire v_66382;
wire v_66383;
wire v_66384;
wire v_66385;
wire v_66386;
wire v_66387;
wire v_66388;
wire v_66389;
wire v_66390;
wire v_66391;
wire v_66392;
wire v_66393;
wire v_66394;
wire v_66395;
wire v_66396;
wire v_66397;
wire v_66398;
wire v_66399;
wire v_66400;
wire v_66401;
wire v_66402;
wire v_66403;
wire v_66404;
wire v_66405;
wire v_66406;
wire v_66407;
wire v_66408;
wire v_66409;
wire v_66410;
wire v_66411;
wire v_66412;
wire v_66413;
wire v_66414;
wire v_66415;
wire v_66416;
wire v_66417;
wire v_66418;
wire v_66419;
wire v_66420;
wire v_66421;
wire v_66422;
wire v_66423;
wire v_66424;
wire v_66425;
wire v_66426;
wire v_66427;
wire v_66428;
wire v_66429;
wire v_66430;
wire v_66431;
wire v_66432;
wire v_66433;
wire v_66434;
wire v_66435;
wire v_66436;
wire v_66437;
wire v_66438;
wire v_66439;
wire v_66440;
wire v_66441;
wire v_66442;
wire v_66443;
wire v_66444;
wire v_66445;
wire v_66446;
wire v_66447;
wire v_66448;
wire v_66449;
wire v_66450;
wire v_66451;
wire v_66452;
wire v_66453;
wire v_66454;
wire v_66455;
wire v_66456;
wire v_66457;
wire v_66458;
wire v_66459;
wire v_66460;
wire v_66461;
wire v_66462;
wire v_66463;
wire v_66464;
wire v_66465;
wire v_66466;
wire v_66467;
wire v_66468;
wire v_66469;
wire v_66470;
wire v_66471;
wire v_66472;
wire v_66473;
wire v_66474;
wire v_66475;
wire v_66476;
wire v_66477;
wire v_66478;
wire v_66479;
wire v_66480;
wire v_66481;
wire v_66482;
wire v_66483;
wire v_66484;
wire v_66485;
wire v_66486;
wire v_66487;
wire v_66488;
wire v_66489;
wire v_66490;
wire v_66491;
wire v_66492;
wire v_66493;
wire v_66494;
wire v_66495;
wire v_66496;
wire v_66497;
wire v_66498;
wire v_66499;
wire v_66500;
wire v_66501;
wire v_66502;
wire v_66503;
wire v_66504;
wire v_66505;
wire v_66506;
wire v_66507;
wire v_66508;
wire v_66509;
wire v_66510;
wire v_66511;
wire v_66512;
wire v_66513;
wire v_66514;
wire v_66515;
wire v_66516;
wire v_66517;
wire v_66518;
wire v_66519;
wire v_66520;
wire v_66521;
wire v_66522;
wire v_66523;
wire v_66524;
wire v_66525;
wire v_66526;
wire v_66527;
wire v_66528;
wire v_66529;
wire v_66530;
wire v_66531;
wire v_66532;
wire v_66533;
wire v_66534;
wire v_66535;
wire v_66536;
wire v_66537;
wire v_66538;
wire v_66539;
wire v_66540;
wire v_66541;
wire v_66542;
wire v_66543;
wire v_66544;
wire v_66545;
wire v_66546;
wire v_66547;
wire v_66548;
wire v_66549;
wire v_66550;
wire v_66551;
wire v_66552;
wire v_66553;
wire v_66554;
wire v_66555;
wire v_66556;
wire v_66557;
wire v_66558;
wire v_66559;
wire v_66560;
wire v_66561;
wire v_66562;
wire v_66563;
wire v_66564;
wire v_66565;
wire v_66566;
wire v_66567;
wire v_66569;
wire v_66570;
wire v_66571;
wire v_66572;
wire v_66573;
wire v_66574;
wire v_66575;
wire v_66576;
wire v_66577;
wire v_66578;
wire v_66579;
wire v_66580;
wire v_66581;
wire v_66582;
wire v_66583;
wire v_66584;
wire v_66585;
wire v_66586;
wire v_66587;
wire v_66588;
wire v_66589;
wire v_66590;
wire v_66591;
wire v_66592;
wire v_66593;
wire v_66594;
wire v_66595;
wire v_66596;
wire v_66597;
wire v_66598;
wire v_66599;
wire v_66600;
wire v_66601;
wire v_66602;
wire v_66603;
wire v_66604;
wire v_66605;
wire v_66606;
wire v_66607;
wire v_66608;
wire v_66609;
wire v_66610;
wire v_66611;
wire v_66612;
wire v_66613;
wire v_66614;
wire v_66615;
wire v_66616;
wire v_66617;
wire v_66618;
wire v_66619;
wire v_66620;
wire v_66621;
wire v_66622;
wire v_66623;
wire v_66624;
wire v_66625;
wire v_66626;
wire v_66627;
wire v_66628;
wire v_66629;
wire v_66630;
wire v_66631;
wire v_66632;
wire v_66633;
wire v_66634;
wire v_66635;
wire v_66636;
wire v_66637;
wire v_66638;
wire v_66639;
wire v_66640;
wire v_66641;
wire v_66642;
wire v_66643;
wire v_66644;
wire v_66645;
wire v_66646;
wire v_66647;
wire v_66648;
wire v_66649;
wire v_66650;
wire v_66651;
wire v_66652;
wire v_66653;
wire v_66654;
wire v_66655;
wire v_66656;
wire v_66657;
wire v_66658;
wire v_66659;
wire v_66660;
wire v_66661;
wire v_66662;
wire v_66664;
wire v_66665;
wire v_66666;
wire v_66668;
wire v_66669;
wire v_66670;
wire v_66672;
wire v_66673;
wire v_66674;
wire v_66676;
wire v_66677;
wire v_66679;
wire v_66680;
wire v_66681;
wire v_66683;
wire v_66684;
wire v_66685;
wire v_66687;
wire v_66688;
wire v_66689;
wire v_66691;
wire v_66692;
wire v_66693;
wire v_66695;
wire v_66696;
wire v_66697;
wire v_66699;
wire v_66700;
wire v_66701;
wire v_66703;
wire v_66704;
wire v_66705;
wire v_66707;
wire v_66708;
wire v_66709;
wire v_66711;
wire v_66712;
wire v_66713;
wire v_66715;
wire v_66716;
wire v_66717;
wire v_66719;
wire v_66720;
wire v_66721;
wire v_66723;
wire v_66724;
wire v_66725;
wire v_66727;
wire v_66728;
wire v_66729;
wire v_66730;
wire v_66731;
wire v_66732;
wire v_66733;
wire v_66734;
wire v_66735;
wire v_66736;
wire v_66737;
wire v_66738;
wire v_66739;
wire v_66740;
wire v_66741;
wire v_66742;
wire v_66743;
wire v_66744;
wire v_66745;
wire v_66746;
wire v_66747;
wire v_66748;
wire v_66749;
wire v_66750;
wire v_66751;
wire v_66752;
wire v_66753;
wire v_66754;
wire v_66755;
wire v_66756;
wire v_66757;
wire v_66758;
wire v_66759;
wire v_66760;
wire v_66761;
wire v_66762;
wire v_66763;
wire v_66764;
wire v_66765;
wire v_66766;
wire v_66767;
wire v_66768;
wire v_66769;
wire v_66770;
wire v_66771;
wire v_66772;
wire v_66773;
wire v_66774;
wire v_66775;
wire v_66776;
wire v_66777;
wire v_66778;
wire v_66779;
wire v_66780;
wire v_66781;
wire v_66782;
wire v_66783;
wire v_66784;
wire v_66785;
wire v_66786;
wire v_66787;
wire v_66788;
wire v_66789;
wire v_66790;
wire v_66791;
wire v_66792;
wire v_66793;
wire v_66794;
wire v_66795;
wire v_66796;
wire v_66797;
wire v_66798;
wire v_66799;
wire v_66800;
wire v_66801;
wire v_66802;
wire v_66803;
wire v_66804;
wire v_66805;
wire v_66806;
wire v_66807;
wire v_66808;
wire v_66809;
wire v_66810;
wire v_66811;
wire v_66812;
wire v_66813;
wire v_66814;
wire v_66815;
wire v_66816;
wire v_66817;
wire v_66818;
wire v_66819;
wire v_66820;
wire v_66821;
wire v_66822;
wire v_66823;
wire v_66824;
wire v_66825;
wire v_66826;
wire v_66827;
wire v_66829;
wire v_66830;
wire v_66831;
wire v_66832;
wire v_66833;
wire v_66834;
wire v_66835;
wire v_66836;
wire v_66837;
wire v_66838;
wire v_66839;
wire v_66840;
wire v_66841;
wire v_66842;
wire v_66843;
wire v_66844;
wire v_66845;
wire v_66846;
wire v_66847;
wire v_66848;
wire v_66849;
wire v_66850;
wire v_66851;
wire v_66852;
wire v_66853;
wire v_66854;
wire v_66855;
wire v_66856;
wire v_66857;
wire v_66858;
wire v_66859;
wire v_66860;
wire v_66861;
wire v_66862;
wire v_66863;
wire v_66864;
wire v_66865;
wire v_66866;
wire v_66867;
wire v_66868;
wire v_66869;
wire v_66870;
wire v_66871;
wire v_66872;
wire v_66873;
wire v_66874;
wire v_66875;
wire v_66876;
wire v_66877;
wire v_66878;
wire v_66879;
wire v_66880;
wire v_66881;
wire v_66882;
wire v_66883;
wire v_66884;
wire v_66885;
wire v_66886;
wire v_66887;
wire v_66888;
wire v_66889;
wire v_66890;
wire v_66891;
wire v_66892;
wire v_66893;
wire v_66894;
wire v_66895;
wire v_66896;
wire v_66897;
wire v_66898;
wire v_66899;
wire v_66900;
wire v_66901;
wire v_66902;
wire v_66903;
wire v_66904;
wire v_66905;
wire v_66906;
wire v_66907;
wire v_66908;
wire v_66909;
wire v_66910;
wire v_66911;
wire v_66912;
wire v_66913;
wire v_66914;
wire v_66915;
wire v_66916;
wire v_66917;
wire v_66918;
wire v_66919;
wire v_66920;
wire v_66921;
wire v_66922;
wire v_66923;
wire v_66924;
wire v_66925;
wire v_66926;
wire v_66927;
wire v_66928;
wire v_66929;
wire v_66930;
wire v_66931;
wire v_66932;
wire v_66933;
wire v_66934;
wire v_66935;
wire v_66936;
wire v_66937;
wire v_66938;
wire v_66939;
wire v_66940;
wire v_66941;
wire v_66942;
wire v_66943;
wire v_66944;
wire v_66945;
wire v_66946;
wire v_66947;
wire v_66948;
wire v_66949;
wire v_66950;
wire v_66951;
wire v_66952;
wire v_66953;
wire v_66954;
wire v_66955;
wire v_66956;
wire v_66957;
wire v_66958;
wire v_66959;
wire v_66960;
wire v_66961;
wire v_66962;
wire v_66963;
wire v_66964;
wire v_66965;
wire v_66966;
wire v_66967;
wire v_66968;
wire v_66969;
wire v_66970;
wire v_66971;
wire v_66972;
wire v_66973;
wire v_66974;
wire v_66975;
wire v_66976;
wire v_66977;
wire v_66978;
wire v_66979;
wire v_66980;
wire v_66981;
wire v_66982;
wire v_66983;
wire v_66984;
wire v_66985;
wire v_66986;
wire v_66987;
wire v_66988;
wire v_66989;
wire v_66990;
wire v_66991;
wire v_66992;
wire v_66993;
wire v_66994;
wire v_66995;
wire v_66996;
wire v_66997;
wire v_66998;
wire v_66999;
wire v_67000;
wire v_67001;
wire v_67002;
wire v_67003;
wire v_67004;
wire v_67005;
wire v_67006;
wire v_67007;
wire v_67008;
wire v_67009;
wire v_67010;
wire v_67011;
wire v_67012;
wire v_67013;
wire v_67014;
wire v_67015;
wire v_67016;
wire v_67017;
wire v_67018;
wire v_67019;
wire v_67020;
wire v_67021;
wire v_67022;
wire v_67023;
wire v_67024;
wire v_67025;
wire v_67026;
wire v_67027;
wire v_67028;
wire v_67029;
wire v_67030;
wire v_67031;
wire v_67032;
wire v_67033;
wire v_67034;
wire v_67035;
wire v_67036;
wire v_67037;
wire v_67038;
wire v_67039;
wire v_67040;
wire v_67041;
wire v_67042;
wire v_67043;
wire v_67044;
wire v_67045;
wire v_67046;
wire v_67047;
wire v_67048;
wire v_67049;
wire v_67050;
wire v_67051;
wire v_67052;
wire v_67053;
wire v_67054;
wire v_67055;
wire v_67056;
wire v_67057;
wire v_67058;
wire v_67059;
wire v_67060;
wire v_67061;
wire v_67062;
wire v_67063;
wire v_67064;
wire v_67065;
wire v_67066;
wire v_67067;
wire v_67068;
wire v_67069;
wire v_67070;
wire v_67072;
wire v_67073;
wire v_67074;
wire v_67075;
wire v_67076;
wire v_67077;
wire v_67078;
wire v_67079;
wire v_67080;
wire v_67081;
wire v_67082;
wire v_67083;
wire v_67084;
wire v_67085;
wire v_67086;
wire v_67087;
wire v_67088;
wire v_67089;
wire v_67090;
wire v_67091;
wire v_67092;
wire v_67093;
wire v_67094;
wire v_67095;
wire v_67096;
wire v_67097;
wire v_67098;
wire v_67099;
wire v_67100;
wire v_67101;
wire v_67102;
wire v_67103;
wire v_67104;
wire v_67105;
wire v_67106;
wire v_67107;
wire v_67108;
wire v_67109;
wire v_67110;
wire v_67111;
wire v_67112;
wire v_67113;
wire v_67114;
wire v_67115;
wire v_67116;
wire v_67117;
wire v_67118;
wire v_67119;
wire v_67120;
wire v_67121;
wire v_67122;
wire v_67123;
wire v_67124;
wire v_67125;
wire v_67126;
wire v_67127;
wire v_67128;
wire v_67129;
wire v_67130;
wire v_67131;
wire v_67132;
wire v_67133;
wire v_67134;
wire v_67135;
wire v_67136;
wire v_67137;
wire v_67138;
wire v_67139;
wire v_67140;
wire v_67141;
wire v_67142;
wire v_67143;
wire v_67144;
wire v_67145;
wire v_67146;
wire v_67147;
wire v_67148;
wire v_67149;
wire v_67150;
wire v_67151;
wire v_67152;
wire v_67153;
wire v_67154;
wire v_67155;
wire v_67156;
wire v_67157;
wire v_67158;
wire v_67159;
wire v_67160;
wire v_67161;
wire v_67162;
wire v_67163;
wire v_67164;
wire v_67165;
wire v_67166;
wire v_67167;
wire v_67168;
wire v_67169;
wire v_67170;
wire v_67171;
wire v_67172;
wire v_67173;
wire v_67174;
wire v_67175;
wire v_67176;
wire v_67177;
wire v_67178;
wire v_67179;
wire v_67180;
wire v_67181;
wire v_67182;
wire v_67183;
wire v_67184;
wire v_67185;
wire v_67186;
wire v_67187;
wire v_67188;
wire v_67189;
wire v_67190;
wire v_67191;
wire v_67192;
wire v_67193;
wire v_67194;
wire v_67195;
wire v_67196;
wire v_67197;
wire v_67198;
wire v_67199;
wire v_67200;
wire v_67201;
wire v_67202;
wire v_67203;
wire v_67204;
wire v_67205;
wire v_67206;
wire v_67207;
wire v_67208;
wire v_67209;
wire v_67210;
wire v_67211;
wire v_67212;
wire v_67213;
wire v_67214;
wire v_67215;
wire v_67216;
wire v_67217;
wire v_67218;
wire v_67219;
wire v_67220;
wire v_67221;
wire v_67222;
wire v_67223;
wire v_67224;
wire v_67225;
wire v_67226;
wire v_67227;
wire v_67228;
wire v_67229;
wire v_67230;
wire v_67231;
wire v_67232;
wire v_67233;
wire v_67234;
wire v_67235;
wire v_67236;
wire v_67237;
wire v_67238;
wire v_67239;
wire v_67240;
wire v_67241;
wire v_67242;
wire v_67243;
wire v_67244;
wire v_67245;
wire v_67246;
wire v_67247;
wire v_67248;
wire v_67249;
wire v_67250;
wire v_67251;
wire v_67252;
wire v_67253;
wire v_67254;
wire v_67255;
wire v_67256;
wire v_67257;
wire v_67258;
wire v_67259;
wire v_67260;
wire v_67261;
wire v_67262;
wire v_67263;
wire v_67264;
wire v_67265;
wire v_67266;
wire v_67267;
wire v_67268;
wire v_67269;
wire v_67270;
wire v_67271;
wire v_67272;
wire v_67273;
wire v_67274;
wire v_67275;
wire v_67276;
wire v_67277;
wire v_67278;
wire v_67279;
wire v_67280;
wire v_67281;
wire v_67282;
wire v_67283;
wire v_67284;
wire v_67285;
wire v_67286;
wire v_67287;
wire v_67288;
wire v_67289;
wire v_67290;
wire v_67291;
wire v_67292;
wire v_67293;
wire v_67294;
wire v_67295;
wire v_67296;
wire v_67297;
wire v_67298;
wire v_67299;
wire v_67300;
wire v_67301;
wire v_67302;
wire v_67303;
wire v_67304;
wire v_67305;
wire v_67306;
wire v_67307;
wire v_67308;
wire v_67309;
wire v_67310;
wire v_67311;
wire v_67312;
wire v_67313;
wire v_67315;
wire v_67316;
wire v_67317;
wire v_67318;
wire v_67319;
wire v_67320;
wire v_67321;
wire v_67322;
wire v_67323;
wire v_67324;
wire v_67325;
wire v_67326;
wire v_67327;
wire v_67328;
wire v_67329;
wire v_67330;
wire v_67331;
wire v_67332;
wire v_67333;
wire v_67334;
wire v_67335;
wire v_67336;
wire v_67337;
wire v_67338;
wire v_67339;
wire v_67340;
wire v_67341;
wire v_67342;
wire v_67343;
wire v_67344;
wire v_67345;
wire v_67346;
wire v_67347;
wire v_67348;
wire v_67349;
wire v_67350;
wire v_67351;
wire v_67352;
wire v_67353;
wire v_67354;
wire v_67355;
wire v_67356;
wire v_67357;
wire v_67358;
wire v_67359;
wire v_67360;
wire v_67361;
wire v_67362;
wire v_67363;
wire v_67364;
wire v_67365;
wire v_67366;
wire v_67367;
wire v_67368;
wire v_67369;
wire v_67370;
wire v_67371;
wire v_67372;
wire v_67373;
wire v_67374;
wire v_67375;
wire v_67376;
wire v_67377;
wire v_67378;
wire v_67379;
wire v_67380;
wire v_67381;
wire v_67382;
wire v_67383;
wire v_67384;
wire v_67385;
wire v_67386;
wire v_67387;
wire v_67388;
wire v_67389;
wire v_67390;
wire v_67391;
wire v_67392;
wire v_67393;
wire v_67394;
wire v_67395;
wire v_67396;
wire v_67397;
wire v_67398;
wire v_67399;
wire v_67400;
wire v_67401;
wire v_67402;
wire v_67403;
wire v_67404;
wire v_67405;
wire v_67406;
wire v_67407;
wire v_67408;
wire v_67409;
wire v_67410;
wire v_67411;
wire v_67412;
wire v_67413;
wire v_67414;
wire v_67415;
wire v_67416;
wire v_67417;
wire v_67418;
wire v_67419;
wire v_67420;
wire v_67421;
wire v_67422;
wire v_67423;
wire v_67424;
wire v_67425;
wire v_67426;
wire v_67427;
wire v_67428;
wire v_67429;
wire v_67430;
wire v_67431;
wire v_67432;
wire v_67433;
wire v_67434;
wire v_67435;
wire v_67436;
wire v_67437;
wire v_67438;
wire v_67439;
wire v_67440;
wire v_67441;
wire v_67442;
wire v_67443;
wire v_67444;
wire v_67445;
wire v_67446;
wire v_67447;
wire v_67448;
wire v_67449;
wire v_67450;
wire v_67451;
wire v_67452;
wire v_67453;
wire v_67454;
wire v_67455;
wire v_67456;
wire v_67457;
wire v_67458;
wire v_67459;
wire v_67460;
wire v_67461;
wire v_67462;
wire v_67463;
wire v_67464;
wire v_67465;
wire v_67466;
wire v_67467;
wire v_67468;
wire v_67469;
wire v_67470;
wire v_67471;
wire v_67472;
wire v_67473;
wire v_67474;
wire v_67475;
wire v_67476;
wire v_67477;
wire v_67478;
wire v_67479;
wire v_67480;
wire v_67481;
wire v_67482;
wire v_67483;
wire v_67484;
wire v_67485;
wire v_67486;
wire v_67487;
wire v_67488;
wire v_67489;
wire v_67490;
wire v_67491;
wire v_67492;
wire v_67493;
wire v_67494;
wire v_67495;
wire v_67496;
wire v_67497;
wire v_67498;
wire v_67499;
wire v_67500;
wire v_67501;
wire v_67502;
wire v_67503;
wire v_67504;
wire v_67505;
wire v_67506;
wire v_67507;
wire v_67508;
wire v_67509;
wire v_67510;
wire v_67511;
wire v_67512;
wire v_67513;
wire v_67514;
wire v_67515;
wire v_67516;
wire v_67517;
wire v_67518;
wire v_67519;
wire v_67520;
wire v_67521;
wire v_67522;
wire v_67523;
wire v_67524;
wire v_67525;
wire v_67526;
wire v_67527;
wire v_67528;
wire v_67529;
wire v_67530;
wire v_67531;
wire v_67532;
wire v_67533;
wire v_67534;
wire v_67535;
wire v_67536;
wire v_67537;
wire v_67538;
wire v_67539;
wire v_67540;
wire v_67541;
wire v_67542;
wire v_67543;
wire v_67544;
wire v_67545;
wire v_67546;
wire v_67547;
wire v_67548;
wire v_67549;
wire v_67550;
wire v_67551;
wire v_67552;
wire v_67553;
wire v_67554;
wire v_67555;
wire v_67556;
wire v_67558;
wire v_67559;
wire v_67560;
wire v_67561;
wire v_67562;
wire v_67563;
wire v_67564;
wire v_67565;
wire v_67566;
wire v_67567;
wire v_67568;
wire v_67569;
wire v_67570;
wire v_67571;
wire v_67572;
wire v_67573;
wire v_67574;
wire v_67575;
wire v_67576;
wire v_67577;
wire v_67578;
wire v_67579;
wire v_67580;
wire v_67581;
wire v_67582;
wire v_67583;
wire v_67584;
wire v_67585;
wire v_67586;
wire v_67587;
wire v_67588;
wire v_67589;
wire v_67590;
wire v_67591;
wire v_67592;
wire v_67593;
wire v_67594;
wire v_67595;
wire v_67596;
wire v_67597;
wire v_67598;
wire v_67599;
wire v_67600;
wire v_67601;
wire v_67602;
wire v_67603;
wire v_67604;
wire v_67605;
wire v_67606;
wire v_67607;
wire v_67608;
wire v_67609;
wire v_67610;
wire v_67611;
wire v_67612;
wire v_67613;
wire v_67614;
wire v_67615;
wire v_67616;
wire v_67617;
wire v_67618;
wire v_67619;
wire v_67620;
wire v_67621;
wire v_67622;
wire v_67623;
wire v_67624;
wire v_67625;
wire v_67626;
wire v_67627;
wire v_67628;
wire v_67629;
wire v_67630;
wire v_67631;
wire v_67632;
wire v_67633;
wire v_67634;
wire v_67635;
wire v_67636;
wire v_67637;
wire v_67638;
wire v_67639;
wire v_67640;
wire v_67641;
wire v_67642;
wire v_67643;
wire v_67644;
wire v_67645;
wire v_67646;
wire v_67647;
wire v_67648;
wire v_67649;
wire v_67650;
wire v_67651;
wire v_67652;
wire v_67653;
wire v_67654;
wire v_67655;
wire v_67656;
wire v_67657;
wire v_67658;
wire v_67659;
wire v_67660;
wire v_67661;
wire v_67662;
wire v_67663;
wire v_67664;
wire v_67665;
wire v_67666;
wire v_67667;
wire v_67668;
wire v_67669;
wire v_67670;
wire v_67671;
wire v_67672;
wire v_67673;
wire v_67674;
wire v_67675;
wire v_67676;
wire v_67677;
wire v_67678;
wire v_67679;
wire v_67680;
wire v_67681;
wire v_67682;
wire v_67683;
wire v_67684;
wire v_67685;
wire v_67686;
wire v_67687;
wire v_67688;
wire v_67689;
wire v_67690;
wire v_67691;
wire v_67692;
wire v_67693;
wire v_67694;
wire v_67695;
wire v_67696;
wire v_67697;
wire v_67698;
wire v_67699;
wire v_67700;
wire v_67701;
wire v_67702;
wire v_67703;
wire v_67704;
wire v_67705;
wire v_67706;
wire v_67707;
wire v_67708;
wire v_67709;
wire v_67710;
wire v_67711;
wire v_67712;
wire v_67713;
wire v_67714;
wire v_67715;
wire v_67716;
wire v_67717;
wire v_67718;
wire v_67719;
wire v_67720;
wire v_67721;
wire v_67722;
wire v_67723;
wire v_67724;
wire v_67725;
wire v_67726;
wire v_67727;
wire v_67728;
wire v_67729;
wire v_67730;
wire v_67731;
wire v_67732;
wire v_67733;
wire v_67734;
wire v_67735;
wire v_67736;
wire v_67737;
wire v_67738;
wire v_67739;
wire v_67740;
wire v_67741;
wire v_67742;
wire v_67743;
wire v_67744;
wire v_67745;
wire v_67746;
wire v_67747;
wire v_67748;
wire v_67749;
wire v_67750;
wire v_67751;
wire v_67752;
wire v_67753;
wire v_67754;
wire v_67755;
wire v_67756;
wire v_67757;
wire v_67758;
wire v_67759;
wire v_67760;
wire v_67761;
wire v_67762;
wire v_67763;
wire v_67764;
wire v_67765;
wire v_67766;
wire v_67767;
wire v_67768;
wire v_67769;
wire v_67770;
wire v_67771;
wire v_67772;
wire v_67773;
wire v_67774;
wire v_67775;
wire v_67776;
wire v_67777;
wire v_67778;
wire v_67779;
wire v_67780;
wire v_67781;
wire v_67782;
wire v_67783;
wire v_67784;
wire v_67785;
wire v_67786;
wire v_67787;
wire v_67788;
wire v_67789;
wire v_67790;
wire v_67791;
wire v_67792;
wire v_67793;
wire v_67794;
wire v_67795;
wire v_67796;
wire v_67797;
wire v_67798;
wire v_67799;
wire v_67801;
wire v_67802;
wire v_67803;
wire v_67804;
wire v_67805;
wire v_67806;
wire v_67807;
wire v_67808;
wire v_67809;
wire v_67810;
wire v_67811;
wire v_67812;
wire v_67813;
wire v_67814;
wire v_67815;
wire v_67816;
wire v_67817;
wire v_67818;
wire v_67819;
wire v_67820;
wire v_67821;
wire v_67822;
wire v_67823;
wire v_67824;
wire v_67825;
wire v_67826;
wire v_67827;
wire v_67828;
wire v_67829;
wire v_67830;
wire v_67831;
wire v_67832;
wire v_67833;
wire v_67834;
wire v_67835;
wire v_67836;
wire v_67837;
wire v_67838;
wire v_67839;
wire v_67840;
wire v_67841;
wire v_67842;
wire v_67843;
wire v_67844;
wire v_67845;
wire v_67846;
wire v_67847;
wire v_67848;
wire v_67849;
wire v_67850;
wire v_67851;
wire v_67852;
wire v_67853;
wire v_67854;
wire v_67855;
wire v_67856;
wire v_67857;
wire v_67858;
wire v_67859;
wire v_67860;
wire v_67861;
wire v_67862;
wire v_67863;
wire v_67864;
wire v_67865;
wire v_67866;
wire v_67867;
wire v_67868;
wire v_67869;
wire v_67870;
wire v_67871;
wire v_67872;
wire v_67873;
wire v_67874;
wire v_67875;
wire v_67876;
wire v_67877;
wire v_67878;
wire v_67879;
wire v_67880;
wire v_67881;
wire v_67882;
wire v_67883;
wire v_67884;
wire v_67885;
wire v_67886;
wire v_67887;
wire v_67888;
wire v_67889;
wire v_67890;
wire v_67891;
wire v_67892;
wire v_67893;
wire v_67894;
wire v_67895;
wire v_67896;
wire v_67897;
wire v_67898;
wire v_67899;
wire v_67900;
wire v_67901;
wire v_67902;
wire v_67903;
wire v_67904;
wire v_67905;
wire v_67906;
wire v_67907;
wire v_67908;
wire v_67909;
wire v_67910;
wire v_67911;
wire v_67912;
wire v_67913;
wire v_67914;
wire v_67915;
wire v_67916;
wire v_67917;
wire v_67918;
wire v_67919;
wire v_67920;
wire v_67921;
wire v_67922;
wire v_67923;
wire v_67924;
wire v_67925;
wire v_67926;
wire v_67927;
wire v_67928;
wire v_67929;
wire v_67930;
wire v_67931;
wire v_67932;
wire v_67933;
wire v_67934;
wire v_67935;
wire v_67936;
wire v_67937;
wire v_67938;
wire v_67939;
wire v_67940;
wire v_67941;
wire v_67942;
wire v_67943;
wire v_67944;
wire v_67945;
wire v_67946;
wire v_67947;
wire v_67948;
wire v_67949;
wire v_67950;
wire v_67951;
wire v_67952;
wire v_67953;
wire v_67954;
wire v_67955;
wire v_67956;
wire v_67957;
wire v_67958;
wire v_67959;
wire v_67960;
wire v_67961;
wire v_67962;
wire v_67963;
wire v_67964;
wire v_67965;
wire v_67966;
wire v_67967;
wire v_67968;
wire v_67969;
wire v_67970;
wire v_67971;
wire v_67972;
wire v_67973;
wire v_67974;
wire v_67975;
wire v_67976;
wire v_67977;
wire v_67978;
wire v_67979;
wire v_67980;
wire v_67981;
wire v_67982;
wire v_67983;
wire v_67984;
wire v_67985;
wire v_67986;
wire v_67987;
wire v_67988;
wire v_67989;
wire v_67990;
wire v_67991;
wire v_67992;
wire v_67993;
wire v_67994;
wire v_67995;
wire v_67996;
wire v_67997;
wire v_67998;
wire v_67999;
wire v_68000;
wire v_68001;
wire v_68002;
wire v_68003;
wire v_68004;
wire v_68005;
wire v_68006;
wire v_68007;
wire v_68008;
wire v_68009;
wire v_68010;
wire v_68011;
wire v_68012;
wire v_68013;
wire v_68014;
wire v_68015;
wire v_68016;
wire v_68017;
wire v_68018;
wire v_68019;
wire v_68020;
wire v_68021;
wire v_68022;
wire v_68023;
wire v_68024;
wire v_68025;
wire v_68026;
wire v_68027;
wire v_68028;
wire v_68029;
wire v_68030;
wire v_68031;
wire v_68032;
wire v_68033;
wire v_68034;
wire v_68035;
wire v_68036;
wire v_68037;
wire v_68038;
wire v_68039;
wire v_68040;
wire v_68041;
wire v_68042;
wire v_68044;
wire v_68045;
wire v_68046;
wire v_68047;
wire v_68048;
wire v_68049;
wire v_68050;
wire v_68051;
wire v_68052;
wire v_68053;
wire v_68054;
wire v_68055;
wire v_68056;
wire v_68057;
wire v_68058;
wire v_68059;
wire v_68060;
wire v_68061;
wire v_68062;
wire v_68063;
wire v_68064;
wire v_68065;
wire v_68066;
wire v_68067;
wire v_68068;
wire v_68069;
wire v_68070;
wire v_68071;
wire v_68072;
wire v_68073;
wire v_68074;
wire v_68075;
wire v_68076;
wire v_68077;
wire v_68078;
wire v_68079;
wire v_68080;
wire v_68081;
wire v_68082;
wire v_68083;
wire v_68084;
wire v_68085;
wire v_68086;
wire v_68087;
wire v_68088;
wire v_68089;
wire v_68090;
wire v_68091;
wire v_68092;
wire v_68093;
wire v_68094;
wire v_68095;
wire v_68096;
wire v_68097;
wire v_68098;
wire v_68099;
wire v_68100;
wire v_68101;
wire v_68102;
wire v_68103;
wire v_68104;
wire v_68105;
wire v_68106;
wire v_68107;
wire v_68108;
wire v_68109;
wire v_68110;
wire v_68111;
wire v_68112;
wire v_68113;
wire v_68114;
wire v_68115;
wire v_68116;
wire v_68117;
wire v_68118;
wire v_68119;
wire v_68120;
wire v_68121;
wire v_68122;
wire v_68123;
wire v_68124;
wire v_68125;
wire v_68126;
wire v_68127;
wire v_68128;
wire v_68129;
wire v_68130;
wire v_68131;
wire v_68132;
wire v_68133;
wire v_68134;
wire v_68135;
wire v_68136;
wire v_68137;
wire v_68138;
wire v_68139;
wire v_68140;
wire v_68141;
wire v_68142;
wire v_68143;
wire v_68144;
wire v_68145;
wire v_68146;
wire v_68147;
wire v_68148;
wire v_68149;
wire v_68150;
wire v_68151;
wire v_68152;
wire v_68153;
wire v_68154;
wire v_68155;
wire v_68156;
wire v_68157;
wire v_68158;
wire v_68159;
wire v_68160;
wire v_68161;
wire v_68162;
wire v_68163;
wire v_68164;
wire v_68165;
wire v_68166;
wire v_68167;
wire v_68168;
wire v_68169;
wire v_68170;
wire v_68171;
wire v_68172;
wire v_68173;
wire v_68174;
wire v_68175;
wire v_68176;
wire v_68177;
wire v_68178;
wire v_68179;
wire v_68180;
wire v_68181;
wire v_68182;
wire v_68183;
wire v_68184;
wire v_68185;
wire v_68186;
wire v_68187;
wire v_68188;
wire v_68189;
wire v_68190;
wire v_68191;
wire v_68192;
wire v_68193;
wire v_68194;
wire v_68195;
wire v_68196;
wire v_68197;
wire v_68198;
wire v_68199;
wire v_68200;
wire v_68201;
wire v_68202;
wire v_68203;
wire v_68204;
wire v_68205;
wire v_68206;
wire v_68207;
wire v_68208;
wire v_68209;
wire v_68210;
wire v_68211;
wire v_68212;
wire v_68213;
wire v_68214;
wire v_68215;
wire v_68216;
wire v_68217;
wire v_68218;
wire v_68219;
wire v_68220;
wire v_68221;
wire v_68222;
wire v_68223;
wire v_68224;
wire v_68225;
wire v_68226;
wire v_68227;
wire v_68228;
wire v_68229;
wire v_68230;
wire v_68231;
wire v_68232;
wire v_68233;
wire v_68234;
wire v_68235;
wire v_68236;
wire v_68237;
wire v_68238;
wire v_68239;
wire v_68240;
wire v_68241;
wire v_68242;
wire v_68243;
wire v_68244;
wire v_68245;
wire v_68246;
wire v_68247;
wire v_68248;
wire v_68249;
wire v_68250;
wire v_68251;
wire v_68252;
wire v_68253;
wire v_68254;
wire v_68255;
wire v_68256;
wire v_68257;
wire v_68258;
wire v_68259;
wire v_68260;
wire v_68261;
wire v_68262;
wire v_68263;
wire v_68264;
wire v_68265;
wire v_68266;
wire v_68267;
wire v_68268;
wire v_68269;
wire v_68270;
wire v_68271;
wire v_68272;
wire v_68273;
wire v_68274;
wire v_68275;
wire v_68276;
wire v_68277;
wire v_68278;
wire v_68279;
wire v_68280;
wire v_68281;
wire v_68282;
wire v_68283;
wire v_68284;
wire v_68285;
wire v_68287;
wire v_68288;
wire v_68289;
wire v_68290;
wire v_68291;
wire v_68292;
wire v_68293;
wire v_68294;
wire v_68295;
wire v_68296;
wire v_68297;
wire v_68298;
wire v_68299;
wire v_68300;
wire v_68301;
wire v_68302;
wire v_68303;
wire v_68304;
wire v_68305;
wire v_68306;
wire v_68307;
wire v_68308;
wire v_68309;
wire v_68310;
wire v_68311;
wire v_68312;
wire v_68313;
wire v_68314;
wire v_68315;
wire v_68316;
wire v_68317;
wire v_68318;
wire v_68319;
wire v_68320;
wire v_68321;
wire v_68322;
wire v_68323;
wire v_68324;
wire v_68325;
wire v_68326;
wire v_68327;
wire v_68328;
wire v_68329;
wire v_68330;
wire v_68331;
wire v_68332;
wire v_68333;
wire v_68334;
wire v_68335;
wire v_68336;
wire v_68337;
wire v_68338;
wire v_68339;
wire v_68340;
wire v_68341;
wire v_68342;
wire v_68343;
wire v_68344;
wire v_68345;
wire v_68346;
wire v_68347;
wire v_68348;
wire v_68349;
wire v_68350;
wire v_68351;
wire v_68352;
wire v_68353;
wire v_68354;
wire v_68355;
wire v_68356;
wire v_68357;
wire v_68358;
wire v_68359;
wire v_68360;
wire v_68361;
wire v_68362;
wire v_68363;
wire v_68364;
wire v_68365;
wire v_68366;
wire v_68367;
wire v_68368;
wire v_68369;
wire v_68370;
wire v_68371;
wire v_68372;
wire v_68373;
wire v_68374;
wire v_68375;
wire v_68376;
wire v_68377;
wire v_68378;
wire v_68379;
wire v_68380;
wire v_68381;
wire v_68382;
wire v_68383;
wire v_68384;
wire v_68385;
wire v_68386;
wire v_68387;
wire v_68388;
wire v_68389;
wire v_68390;
wire v_68391;
wire v_68392;
wire v_68393;
wire v_68394;
wire v_68395;
wire v_68396;
wire v_68397;
wire v_68398;
wire v_68399;
wire v_68400;
wire v_68401;
wire v_68402;
wire v_68403;
wire v_68404;
wire v_68405;
wire v_68406;
wire v_68407;
wire v_68408;
wire v_68409;
wire v_68410;
wire v_68411;
wire v_68412;
wire v_68413;
wire v_68414;
wire v_68415;
wire v_68416;
wire v_68417;
wire v_68418;
wire v_68419;
wire v_68420;
wire v_68421;
wire v_68422;
wire v_68423;
wire v_68424;
wire v_68425;
wire v_68426;
wire v_68427;
wire v_68428;
wire v_68429;
wire v_68430;
wire v_68431;
wire v_68432;
wire v_68433;
wire v_68434;
wire v_68435;
wire v_68436;
wire v_68437;
wire v_68438;
wire v_68439;
wire v_68440;
wire v_68441;
wire v_68442;
wire v_68443;
wire v_68444;
wire v_68445;
wire v_68446;
wire v_68447;
wire v_68448;
wire v_68449;
wire v_68450;
wire v_68451;
wire v_68452;
wire v_68453;
wire v_68454;
wire v_68455;
wire v_68456;
wire v_68457;
wire v_68458;
wire v_68459;
wire v_68460;
wire v_68461;
wire v_68462;
wire v_68463;
wire v_68464;
wire v_68465;
wire v_68466;
wire v_68467;
wire v_68468;
wire v_68469;
wire v_68470;
wire v_68471;
wire v_68472;
wire v_68473;
wire v_68474;
wire v_68475;
wire v_68476;
wire v_68477;
wire v_68478;
wire v_68479;
wire v_68480;
wire v_68481;
wire v_68482;
wire v_68483;
wire v_68484;
wire v_68485;
wire v_68486;
wire v_68487;
wire v_68488;
wire v_68489;
wire v_68490;
wire v_68491;
wire v_68492;
wire v_68493;
wire v_68494;
wire v_68495;
wire v_68496;
wire v_68497;
wire v_68498;
wire v_68499;
wire v_68500;
wire v_68501;
wire v_68502;
wire v_68503;
wire v_68504;
wire v_68505;
wire v_68506;
wire v_68507;
wire v_68508;
wire v_68509;
wire v_68510;
wire v_68511;
wire v_68512;
wire v_68513;
wire v_68514;
wire v_68515;
wire v_68516;
wire v_68517;
wire v_68518;
wire v_68519;
wire v_68520;
wire v_68521;
wire v_68522;
wire v_68523;
wire v_68524;
wire v_68525;
wire v_68526;
wire v_68527;
wire v_68528;
wire v_68530;
wire v_68531;
wire v_68532;
wire v_68533;
wire v_68534;
wire v_68535;
wire v_68536;
wire v_68537;
wire v_68538;
wire v_68539;
wire v_68540;
wire v_68541;
wire v_68542;
wire v_68543;
wire v_68544;
wire v_68545;
wire v_68546;
wire v_68547;
wire v_68548;
wire v_68549;
wire v_68550;
wire v_68551;
wire v_68552;
wire v_68553;
wire v_68554;
wire v_68555;
wire v_68556;
wire v_68557;
wire v_68558;
wire v_68559;
wire v_68560;
wire v_68561;
wire v_68562;
wire v_68563;
wire v_68564;
wire v_68565;
wire v_68566;
wire v_68567;
wire v_68568;
wire v_68569;
wire v_68570;
wire v_68571;
wire v_68572;
wire v_68573;
wire v_68574;
wire v_68575;
wire v_68576;
wire v_68577;
wire v_68578;
wire v_68579;
wire v_68580;
wire v_68581;
wire v_68582;
wire v_68583;
wire v_68584;
wire v_68585;
wire v_68586;
wire v_68587;
wire v_68588;
wire v_68589;
wire v_68590;
wire v_68591;
wire v_68592;
wire v_68593;
wire v_68594;
wire v_68595;
wire v_68596;
wire v_68597;
wire v_68598;
wire v_68599;
wire v_68600;
wire v_68601;
wire v_68602;
wire v_68603;
wire v_68604;
wire v_68605;
wire v_68606;
wire v_68607;
wire v_68608;
wire v_68609;
wire v_68610;
wire v_68611;
wire v_68612;
wire v_68613;
wire v_68614;
wire v_68615;
wire v_68616;
wire v_68617;
wire v_68618;
wire v_68619;
wire v_68620;
wire v_68621;
wire v_68622;
wire v_68623;
wire v_68624;
wire v_68625;
wire v_68626;
wire v_68627;
wire v_68628;
wire v_68629;
wire v_68630;
wire v_68631;
wire v_68632;
wire v_68633;
wire v_68634;
wire v_68635;
wire v_68636;
wire v_68637;
wire v_68638;
wire v_68639;
wire v_68640;
wire v_68641;
wire v_68642;
wire v_68643;
wire v_68644;
wire v_68645;
wire v_68646;
wire v_68647;
wire v_68648;
wire v_68649;
wire v_68650;
wire v_68651;
wire v_68652;
wire v_68653;
wire v_68654;
wire v_68655;
wire v_68656;
wire v_68657;
wire v_68658;
wire v_68659;
wire v_68660;
wire v_68661;
wire v_68662;
wire v_68663;
wire v_68664;
wire v_68665;
wire v_68666;
wire v_68667;
wire v_68668;
wire v_68669;
wire v_68670;
wire v_68671;
wire v_68672;
wire v_68673;
wire v_68674;
wire v_68675;
wire v_68676;
wire v_68677;
wire v_68678;
wire v_68679;
wire v_68680;
wire v_68681;
wire v_68682;
wire v_68683;
wire v_68684;
wire v_68685;
wire v_68686;
wire v_68687;
wire v_68688;
wire v_68689;
wire v_68690;
wire v_68691;
wire v_68692;
wire v_68693;
wire v_68694;
wire v_68695;
wire v_68696;
wire v_68697;
wire v_68698;
wire v_68699;
wire v_68700;
wire v_68701;
wire v_68702;
wire v_68703;
wire v_68704;
wire v_68705;
wire v_68706;
wire v_68707;
wire v_68708;
wire v_68709;
wire v_68710;
wire v_68711;
wire v_68712;
wire v_68713;
wire v_68714;
wire v_68715;
wire v_68716;
wire v_68717;
wire v_68718;
wire v_68719;
wire v_68720;
wire v_68721;
wire v_68722;
wire v_68723;
wire v_68724;
wire v_68725;
wire v_68726;
wire v_68727;
wire v_68728;
wire v_68729;
wire v_68730;
wire v_68731;
wire v_68732;
wire v_68733;
wire v_68734;
wire v_68735;
wire v_68736;
wire v_68737;
wire v_68738;
wire v_68739;
wire v_68740;
wire v_68741;
wire v_68742;
wire v_68743;
wire v_68744;
wire v_68745;
wire v_68746;
wire v_68747;
wire v_68748;
wire v_68749;
wire v_68750;
wire v_68751;
wire v_68752;
wire v_68753;
wire v_68754;
wire v_68755;
wire v_68756;
wire v_68757;
wire v_68758;
wire v_68759;
wire v_68760;
wire v_68761;
wire v_68762;
wire v_68763;
wire v_68764;
wire v_68765;
wire v_68766;
wire v_68767;
wire v_68768;
wire v_68769;
wire v_68770;
wire v_68771;
wire v_68773;
wire v_68774;
wire v_68775;
wire v_68776;
wire v_68777;
wire v_68778;
wire v_68779;
wire v_68780;
wire v_68781;
wire v_68782;
wire v_68783;
wire v_68784;
wire v_68785;
wire v_68786;
wire v_68787;
wire v_68788;
wire v_68789;
wire v_68790;
wire v_68791;
wire v_68792;
wire v_68793;
wire v_68794;
wire v_68795;
wire v_68796;
wire v_68797;
wire v_68798;
wire v_68799;
wire v_68800;
wire v_68801;
wire v_68802;
wire v_68803;
wire v_68804;
wire v_68805;
wire v_68806;
wire v_68807;
wire v_68808;
wire v_68809;
wire v_68810;
wire v_68811;
wire v_68812;
wire v_68813;
wire v_68814;
wire v_68815;
wire v_68816;
wire v_68817;
wire v_68818;
wire v_68819;
wire v_68820;
wire v_68821;
wire v_68822;
wire v_68823;
wire v_68824;
wire v_68825;
wire v_68826;
wire v_68827;
wire v_68828;
wire v_68829;
wire v_68830;
wire v_68831;
wire v_68832;
wire v_68833;
wire v_68834;
wire v_68835;
wire v_68836;
wire v_68837;
wire v_68838;
wire v_68839;
wire v_68840;
wire v_68841;
wire v_68842;
wire v_68843;
wire v_68844;
wire v_68845;
wire v_68846;
wire v_68847;
wire v_68848;
wire v_68849;
wire v_68850;
wire v_68851;
wire v_68852;
wire v_68853;
wire v_68854;
wire v_68855;
wire v_68856;
wire v_68857;
wire v_68858;
wire v_68859;
wire v_68860;
wire v_68861;
wire v_68862;
wire v_68863;
wire v_68864;
wire v_68865;
wire v_68866;
wire v_68867;
wire v_68868;
wire v_68869;
wire v_68870;
wire v_68871;
wire v_68872;
wire v_68873;
wire v_68874;
wire v_68875;
wire v_68876;
wire v_68877;
wire v_68878;
wire v_68879;
wire v_68880;
wire v_68881;
wire v_68882;
wire v_68883;
wire v_68884;
wire v_68885;
wire v_68886;
wire v_68887;
wire v_68888;
wire v_68889;
wire v_68890;
wire v_68891;
wire v_68892;
wire v_68893;
wire v_68894;
wire v_68895;
wire v_68896;
wire v_68897;
wire v_68898;
wire v_68899;
wire v_68900;
wire v_68901;
wire v_68902;
wire v_68903;
wire v_68904;
wire v_68905;
wire v_68906;
wire v_68907;
wire v_68908;
wire v_68909;
wire v_68910;
wire v_68911;
wire v_68912;
wire v_68913;
wire v_68914;
wire v_68915;
wire v_68916;
wire v_68917;
wire v_68918;
wire v_68919;
wire v_68920;
wire v_68921;
wire v_68922;
wire v_68923;
wire v_68924;
wire v_68925;
wire v_68926;
wire v_68927;
wire v_68928;
wire v_68929;
wire v_68930;
wire v_68931;
wire v_68932;
wire v_68933;
wire v_68934;
wire v_68935;
wire v_68936;
wire v_68937;
wire v_68938;
wire v_68939;
wire v_68940;
wire v_68941;
wire v_68942;
wire v_68943;
wire v_68944;
wire v_68945;
wire v_68946;
wire v_68947;
wire v_68948;
wire v_68949;
wire v_68950;
wire v_68951;
wire v_68952;
wire v_68953;
wire v_68954;
wire v_68955;
wire v_68956;
wire v_68957;
wire v_68958;
wire v_68959;
wire v_68960;
wire v_68961;
wire v_68962;
wire v_68963;
wire v_68964;
wire v_68965;
wire v_68966;
wire v_68967;
wire v_68968;
wire v_68969;
wire v_68970;
wire v_68971;
wire v_68972;
wire v_68973;
wire v_68974;
wire v_68975;
wire v_68976;
wire v_68977;
wire v_68978;
wire v_68979;
wire v_68980;
wire v_68981;
wire v_68982;
wire v_68983;
wire v_68984;
wire v_68985;
wire v_68986;
wire v_68987;
wire v_68988;
wire v_68989;
wire v_68990;
wire v_68991;
wire v_68992;
wire v_68993;
wire v_68994;
wire v_68995;
wire v_68996;
wire v_68997;
wire v_68998;
wire v_68999;
wire v_69000;
wire v_69001;
wire v_69002;
wire v_69003;
wire v_69004;
wire v_69005;
wire v_69006;
wire v_69007;
wire v_69008;
wire v_69009;
wire v_69010;
wire v_69011;
wire v_69012;
wire v_69013;
wire v_69014;
wire v_69016;
wire v_69017;
wire v_69018;
wire v_69019;
wire v_69020;
wire v_69021;
wire v_69022;
wire v_69023;
wire v_69024;
wire v_69025;
wire v_69026;
wire v_69027;
wire v_69028;
wire v_69029;
wire v_69030;
wire v_69031;
wire v_69032;
wire v_69033;
wire v_69034;
wire v_69035;
wire v_69036;
wire v_69037;
wire v_69038;
wire v_69039;
wire v_69040;
wire v_69041;
wire v_69042;
wire v_69043;
wire v_69044;
wire v_69045;
wire v_69046;
wire v_69047;
wire v_69048;
wire v_69049;
wire v_69050;
wire v_69051;
wire v_69052;
wire v_69053;
wire v_69054;
wire v_69055;
wire v_69056;
wire v_69057;
wire v_69058;
wire v_69059;
wire v_69060;
wire v_69061;
wire v_69062;
wire v_69063;
wire v_69064;
wire v_69065;
wire v_69066;
wire v_69067;
wire v_69068;
wire v_69069;
wire v_69070;
wire v_69071;
wire v_69072;
wire v_69073;
wire v_69074;
wire v_69075;
wire v_69076;
wire v_69077;
wire v_69078;
wire v_69079;
wire v_69080;
wire v_69081;
wire v_69082;
wire v_69083;
wire v_69084;
wire v_69085;
wire v_69086;
wire v_69087;
wire v_69088;
wire v_69089;
wire v_69090;
wire v_69091;
wire v_69092;
wire v_69093;
wire v_69094;
wire v_69095;
wire v_69096;
wire v_69097;
wire v_69098;
wire v_69099;
wire v_69100;
wire v_69101;
wire v_69102;
wire v_69103;
wire v_69104;
wire v_69105;
wire v_69106;
wire v_69107;
wire v_69108;
wire v_69109;
wire v_69110;
wire v_69111;
wire v_69112;
wire v_69113;
wire v_69114;
wire v_69115;
wire v_69116;
wire v_69117;
wire v_69118;
wire v_69119;
wire v_69120;
wire v_69121;
wire v_69122;
wire v_69123;
wire v_69124;
wire v_69125;
wire v_69126;
wire v_69127;
wire v_69128;
wire v_69129;
wire v_69130;
wire v_69131;
wire v_69132;
wire v_69133;
wire v_69134;
wire v_69135;
wire v_69136;
wire v_69137;
wire v_69138;
wire v_69139;
wire v_69140;
wire v_69141;
wire v_69142;
wire v_69143;
wire v_69144;
wire v_69145;
wire v_69146;
wire v_69147;
wire v_69148;
wire v_69149;
wire v_69150;
wire v_69151;
wire v_69152;
wire v_69153;
wire v_69154;
wire v_69155;
wire v_69156;
wire v_69157;
wire v_69158;
wire v_69159;
wire v_69160;
wire v_69161;
wire v_69162;
wire v_69163;
wire v_69164;
wire v_69165;
wire v_69166;
wire v_69167;
wire v_69168;
wire v_69169;
wire v_69170;
wire v_69171;
wire v_69172;
wire v_69173;
wire v_69174;
wire v_69175;
wire v_69176;
wire v_69177;
wire v_69178;
wire v_69179;
wire v_69180;
wire v_69181;
wire v_69182;
wire v_69183;
wire v_69184;
wire v_69185;
wire v_69186;
wire v_69187;
wire v_69188;
wire v_69189;
wire v_69190;
wire v_69191;
wire v_69192;
wire v_69193;
wire v_69194;
wire v_69195;
wire v_69196;
wire v_69197;
wire v_69198;
wire v_69199;
wire v_69200;
wire v_69201;
wire v_69202;
wire v_69203;
wire v_69204;
wire v_69205;
wire v_69206;
wire v_69207;
wire v_69208;
wire v_69209;
wire v_69210;
wire v_69211;
wire v_69212;
wire v_69213;
wire v_69214;
wire v_69215;
wire v_69216;
wire v_69217;
wire v_69218;
wire v_69219;
wire v_69220;
wire v_69221;
wire v_69222;
wire v_69223;
wire v_69224;
wire v_69225;
wire v_69226;
wire v_69227;
wire v_69228;
wire v_69229;
wire v_69230;
wire v_69231;
wire v_69232;
wire v_69233;
wire v_69234;
wire v_69235;
wire v_69236;
wire v_69237;
wire v_69238;
wire v_69239;
wire v_69240;
wire v_69241;
wire v_69242;
wire v_69243;
wire v_69244;
wire v_69245;
wire v_69246;
wire v_69247;
wire v_69248;
wire v_69249;
wire v_69250;
wire v_69251;
wire v_69252;
wire v_69253;
wire v_69254;
wire v_69255;
wire v_69256;
wire v_69257;
wire v_69259;
wire v_69260;
wire v_69261;
wire v_69262;
wire v_69263;
wire v_69264;
wire v_69265;
wire v_69266;
wire v_69267;
wire v_69268;
wire v_69269;
wire v_69270;
wire v_69271;
wire v_69272;
wire v_69273;
wire v_69274;
wire v_69275;
wire v_69276;
wire v_69277;
wire v_69278;
wire v_69279;
wire v_69280;
wire v_69281;
wire v_69282;
wire v_69283;
wire v_69284;
wire v_69285;
wire v_69286;
wire v_69287;
wire v_69288;
wire v_69289;
wire v_69290;
wire v_69291;
wire v_69292;
wire v_69293;
wire v_69294;
wire v_69295;
wire v_69296;
wire v_69297;
wire v_69298;
wire v_69299;
wire v_69300;
wire v_69301;
wire v_69302;
wire v_69303;
wire v_69304;
wire v_69305;
wire v_69306;
wire v_69307;
wire v_69308;
wire v_69309;
wire v_69310;
wire v_69311;
wire v_69312;
wire v_69313;
wire v_69314;
wire v_69315;
wire v_69316;
wire v_69317;
wire v_69318;
wire v_69319;
wire v_69320;
wire v_69321;
wire v_69322;
wire v_69323;
wire v_69324;
wire v_69325;
wire v_69326;
wire v_69327;
wire v_69328;
wire v_69329;
wire v_69330;
wire v_69331;
wire v_69332;
wire v_69333;
wire v_69334;
wire v_69335;
wire v_69336;
wire v_69337;
wire v_69338;
wire v_69339;
wire v_69340;
wire v_69341;
wire v_69342;
wire v_69343;
wire v_69344;
wire v_69345;
wire v_69346;
wire v_69347;
wire v_69348;
wire v_69349;
wire v_69350;
wire v_69351;
wire v_69352;
wire v_69353;
wire v_69354;
wire v_69355;
wire v_69356;
wire v_69357;
wire v_69358;
wire v_69359;
wire v_69360;
wire v_69361;
wire v_69362;
wire v_69363;
wire v_69364;
wire v_69365;
wire v_69366;
wire v_69367;
wire v_69368;
wire v_69369;
wire v_69370;
wire v_69371;
wire v_69372;
wire v_69373;
wire v_69374;
wire v_69375;
wire v_69376;
wire v_69377;
wire v_69378;
wire v_69379;
wire v_69380;
wire v_69381;
wire v_69382;
wire v_69383;
wire v_69384;
wire v_69385;
wire v_69386;
wire v_69387;
wire v_69388;
wire v_69389;
wire v_69390;
wire v_69391;
wire v_69392;
wire v_69393;
wire v_69394;
wire v_69395;
wire v_69396;
wire v_69397;
wire v_69398;
wire v_69399;
wire v_69400;
wire v_69401;
wire v_69402;
wire v_69403;
wire v_69404;
wire v_69405;
wire v_69406;
wire v_69407;
wire v_69408;
wire v_69409;
wire v_69410;
wire v_69411;
wire v_69412;
wire v_69413;
wire v_69414;
wire v_69415;
wire v_69416;
wire v_69417;
wire v_69418;
wire v_69419;
wire v_69420;
wire v_69421;
wire v_69422;
wire v_69423;
wire v_69424;
wire v_69425;
wire v_69426;
wire v_69427;
wire v_69428;
wire v_69429;
wire v_69430;
wire v_69431;
wire v_69432;
wire v_69433;
wire v_69434;
wire v_69435;
wire v_69436;
wire v_69437;
wire v_69438;
wire v_69439;
wire v_69440;
wire v_69441;
wire v_69442;
wire v_69443;
wire v_69444;
wire v_69445;
wire v_69446;
wire v_69447;
wire v_69448;
wire v_69449;
wire v_69450;
wire v_69451;
wire v_69452;
wire v_69453;
wire v_69454;
wire v_69455;
wire v_69456;
wire v_69457;
wire v_69458;
wire v_69459;
wire v_69460;
wire v_69461;
wire v_69462;
wire v_69463;
wire v_69464;
wire v_69465;
wire v_69466;
wire v_69467;
wire v_69468;
wire v_69469;
wire v_69470;
wire v_69471;
wire v_69472;
wire v_69473;
wire v_69474;
wire v_69475;
wire v_69476;
wire v_69477;
wire v_69478;
wire v_69479;
wire v_69480;
wire v_69481;
wire v_69482;
wire v_69483;
wire v_69484;
wire v_69485;
wire v_69486;
wire v_69487;
wire v_69488;
wire v_69489;
wire v_69490;
wire v_69491;
wire v_69492;
wire v_69493;
wire v_69494;
wire v_69495;
wire v_69496;
wire v_69497;
wire v_69498;
wire v_69499;
wire v_69500;
wire v_69502;
wire v_69503;
wire v_69504;
wire v_69505;
wire v_69506;
wire v_69507;
wire v_69508;
wire v_69509;
wire v_69510;
wire v_69511;
wire v_69512;
wire v_69513;
wire v_69514;
wire v_69515;
wire v_69516;
wire v_69517;
wire v_69518;
wire v_69519;
wire v_69520;
wire v_69521;
wire v_69522;
wire v_69523;
wire v_69524;
wire v_69525;
wire v_69526;
wire v_69527;
wire v_69528;
wire v_69529;
wire v_69530;
wire v_69531;
wire v_69532;
wire v_69533;
wire v_69534;
wire v_69535;
wire v_69536;
wire v_69537;
wire v_69538;
wire v_69539;
wire v_69540;
wire v_69541;
wire v_69542;
wire v_69543;
wire v_69544;
wire v_69545;
wire v_69546;
wire v_69547;
wire v_69548;
wire v_69549;
wire v_69550;
wire v_69551;
wire v_69552;
wire v_69553;
wire v_69554;
wire v_69555;
wire v_69556;
wire v_69557;
wire v_69558;
wire v_69559;
wire v_69560;
wire v_69561;
wire v_69562;
wire v_69563;
wire v_69564;
wire v_69565;
wire v_69566;
wire v_69567;
wire v_69568;
wire v_69569;
wire v_69570;
wire v_69571;
wire v_69572;
wire v_69573;
wire v_69574;
wire v_69575;
wire v_69576;
wire v_69577;
wire v_69578;
wire v_69579;
wire v_69580;
wire v_69581;
wire v_69582;
wire v_69583;
wire v_69584;
wire v_69585;
wire v_69586;
wire v_69587;
wire v_69588;
wire v_69589;
wire v_69590;
wire v_69591;
wire v_69592;
wire v_69593;
wire v_69594;
wire v_69595;
wire v_69596;
wire v_69597;
wire v_69598;
wire v_69599;
wire v_69600;
wire v_69601;
wire v_69602;
wire v_69603;
wire v_69604;
wire v_69605;
wire v_69606;
wire v_69607;
wire v_69608;
wire v_69609;
wire v_69610;
wire v_69611;
wire v_69612;
wire v_69613;
wire v_69614;
wire v_69615;
wire v_69616;
wire v_69617;
wire v_69618;
wire v_69619;
wire v_69620;
wire v_69621;
wire v_69622;
wire v_69623;
wire v_69624;
wire v_69625;
wire v_69626;
wire v_69627;
wire v_69628;
wire v_69629;
wire v_69630;
wire v_69631;
wire v_69632;
wire v_69633;
wire v_69634;
wire v_69635;
wire v_69636;
wire v_69637;
wire v_69638;
wire v_69639;
wire v_69640;
wire v_69641;
wire v_69642;
wire v_69643;
wire v_69644;
wire v_69645;
wire v_69646;
wire v_69647;
wire v_69648;
wire v_69649;
wire v_69650;
wire v_69651;
wire v_69652;
wire v_69653;
wire v_69654;
wire v_69655;
wire v_69656;
wire v_69657;
wire v_69658;
wire v_69659;
wire v_69660;
wire v_69661;
wire v_69662;
wire v_69663;
wire v_69664;
wire v_69665;
wire v_69666;
wire v_69667;
wire v_69668;
wire v_69669;
wire v_69670;
wire v_69671;
wire v_69672;
wire v_69673;
wire v_69674;
wire v_69675;
wire v_69676;
wire v_69677;
wire v_69678;
wire v_69679;
wire v_69680;
wire v_69681;
wire v_69682;
wire v_69683;
wire v_69684;
wire v_69685;
wire v_69686;
wire v_69687;
wire v_69688;
wire v_69689;
wire v_69690;
wire v_69691;
wire v_69692;
wire v_69693;
wire v_69694;
wire v_69695;
wire v_69696;
wire v_69697;
wire v_69698;
wire v_69699;
wire v_69700;
wire v_69701;
wire v_69702;
wire v_69703;
wire v_69704;
wire v_69705;
wire v_69706;
wire v_69707;
wire v_69708;
wire v_69709;
wire v_69710;
wire v_69711;
wire v_69712;
wire v_69713;
wire v_69714;
wire v_69715;
wire v_69716;
wire v_69717;
wire v_69718;
wire v_69719;
wire v_69720;
wire v_69721;
wire v_69722;
wire v_69723;
wire v_69724;
wire v_69725;
wire v_69726;
wire v_69727;
wire v_69728;
wire v_69729;
wire v_69730;
wire v_69731;
wire v_69732;
wire v_69733;
wire v_69734;
wire v_69735;
wire v_69736;
wire v_69737;
wire v_69738;
wire v_69739;
wire v_69740;
wire v_69741;
wire v_69742;
wire v_69743;
wire v_69745;
wire v_69746;
wire v_69747;
wire v_69748;
wire v_69749;
wire v_69750;
wire v_69751;
wire v_69752;
wire v_69753;
wire v_69754;
wire v_69755;
wire v_69756;
wire v_69757;
wire v_69758;
wire v_69759;
wire v_69760;
wire v_69761;
wire v_69762;
wire v_69763;
wire v_69764;
wire v_69765;
wire v_69766;
wire v_69767;
wire v_69768;
wire v_69769;
wire v_69770;
wire v_69771;
wire v_69772;
wire v_69773;
wire v_69774;
wire v_69775;
wire v_69776;
wire v_69777;
wire v_69778;
wire v_69779;
wire v_69780;
wire v_69781;
wire v_69782;
wire v_69783;
wire v_69784;
wire v_69785;
wire v_69786;
wire v_69787;
wire v_69788;
wire v_69789;
wire v_69790;
wire v_69791;
wire v_69792;
wire v_69793;
wire v_69794;
wire v_69795;
wire v_69796;
wire v_69797;
wire v_69798;
wire v_69799;
wire v_69800;
wire v_69801;
wire v_69802;
wire v_69803;
wire v_69804;
wire v_69805;
wire v_69806;
wire v_69807;
wire v_69808;
wire v_69809;
wire v_69810;
wire v_69811;
wire v_69812;
wire v_69813;
wire v_69814;
wire v_69815;
wire v_69816;
wire v_69817;
wire v_69818;
wire v_69819;
wire v_69820;
wire v_69821;
wire v_69822;
wire v_69823;
wire v_69824;
wire v_69825;
wire v_69826;
wire v_69827;
wire v_69828;
wire v_69829;
wire v_69830;
wire v_69831;
wire v_69832;
wire v_69833;
wire v_69834;
wire v_69835;
wire v_69836;
wire v_69837;
wire v_69838;
wire v_69839;
wire v_69840;
wire v_69841;
wire v_69842;
wire v_69843;
wire v_69844;
wire v_69845;
wire v_69846;
wire v_69847;
wire v_69848;
wire v_69849;
wire v_69850;
wire v_69851;
wire v_69852;
wire v_69853;
wire v_69854;
wire v_69855;
wire v_69856;
wire v_69857;
wire v_69858;
wire v_69859;
wire v_69860;
wire v_69861;
wire v_69862;
wire v_69863;
wire v_69864;
wire v_69865;
wire v_69866;
wire v_69867;
wire v_69868;
wire v_69869;
wire v_69870;
wire v_69871;
wire v_69872;
wire v_69873;
wire v_69874;
wire v_69875;
wire v_69876;
wire v_69877;
wire v_69878;
wire v_69879;
wire v_69880;
wire v_69881;
wire v_69882;
wire v_69883;
wire v_69884;
wire v_69885;
wire v_69886;
wire v_69887;
wire v_69888;
wire v_69889;
wire v_69890;
wire v_69891;
wire v_69892;
wire v_69893;
wire v_69894;
wire v_69895;
wire v_69896;
wire v_69897;
wire v_69898;
wire v_69899;
wire v_69900;
wire v_69901;
wire v_69902;
wire v_69903;
wire v_69904;
wire v_69905;
wire v_69906;
wire v_69907;
wire v_69908;
wire v_69909;
wire v_69910;
wire v_69911;
wire v_69912;
wire v_69913;
wire v_69914;
wire v_69915;
wire v_69916;
wire v_69917;
wire v_69918;
wire v_69919;
wire v_69920;
wire v_69921;
wire v_69922;
wire v_69923;
wire v_69924;
wire v_69925;
wire v_69926;
wire v_69927;
wire v_69928;
wire v_69929;
wire v_69930;
wire v_69931;
wire v_69932;
wire v_69933;
wire v_69934;
wire v_69935;
wire v_69936;
wire v_69937;
wire v_69938;
wire v_69939;
wire v_69940;
wire v_69941;
wire v_69942;
wire v_69943;
wire v_69944;
wire v_69945;
wire v_69946;
wire v_69947;
wire v_69948;
wire v_69949;
wire v_69950;
wire v_69951;
wire v_69952;
wire v_69953;
wire v_69954;
wire v_69955;
wire v_69956;
wire v_69957;
wire v_69958;
wire v_69959;
wire v_69960;
wire v_69961;
wire v_69962;
wire v_69963;
wire v_69964;
wire v_69965;
wire v_69966;
wire v_69967;
wire v_69968;
wire v_69969;
wire v_69970;
wire v_69971;
wire v_69972;
wire v_69973;
wire v_69974;
wire v_69975;
wire v_69976;
wire v_69977;
wire v_69978;
wire v_69979;
wire v_69980;
wire v_69981;
wire v_69982;
wire v_69983;
wire v_69984;
wire v_69985;
wire v_69986;
wire v_69988;
wire v_69989;
wire v_69990;
wire v_69991;
wire v_69992;
wire v_69993;
wire v_69994;
wire v_69995;
wire v_69996;
wire v_69997;
wire v_69998;
wire v_69999;
wire v_70000;
wire v_70001;
wire v_70002;
wire v_70003;
wire v_70004;
wire v_70005;
wire v_70006;
wire v_70007;
wire v_70008;
wire v_70009;
wire v_70010;
wire v_70011;
wire v_70012;
wire v_70013;
wire v_70014;
wire v_70015;
wire v_70016;
wire v_70017;
wire v_70018;
wire v_70019;
wire v_70020;
wire v_70021;
wire v_70022;
wire v_70023;
wire v_70024;
wire v_70025;
wire v_70026;
wire v_70027;
wire v_70028;
wire v_70029;
wire v_70030;
wire v_70031;
wire v_70032;
wire v_70033;
wire v_70034;
wire v_70035;
wire v_70036;
wire v_70037;
wire v_70038;
wire v_70039;
wire v_70040;
wire v_70041;
wire v_70042;
wire v_70043;
wire v_70044;
wire v_70045;
wire v_70046;
wire v_70047;
wire v_70048;
wire v_70049;
wire v_70050;
wire v_70051;
wire v_70052;
wire v_70053;
wire v_70054;
wire v_70055;
wire v_70056;
wire v_70057;
wire v_70058;
wire v_70059;
wire v_70060;
wire v_70061;
wire v_70062;
wire v_70063;
wire v_70064;
wire v_70065;
wire v_70066;
wire v_70067;
wire v_70068;
wire v_70069;
wire v_70070;
wire v_70071;
wire v_70072;
wire v_70073;
wire v_70074;
wire v_70075;
wire v_70076;
wire v_70077;
wire v_70078;
wire v_70079;
wire v_70080;
wire v_70081;
wire v_70082;
wire v_70083;
wire v_70084;
wire v_70085;
wire v_70086;
wire v_70087;
wire v_70088;
wire v_70089;
wire v_70090;
wire v_70091;
wire v_70092;
wire v_70093;
wire v_70094;
wire v_70095;
wire v_70096;
wire v_70097;
wire v_70098;
wire v_70099;
wire v_70100;
wire v_70101;
wire v_70102;
wire v_70103;
wire v_70104;
wire v_70105;
wire v_70106;
wire v_70107;
wire v_70108;
wire v_70109;
wire v_70110;
wire v_70111;
wire v_70112;
wire v_70113;
wire v_70114;
wire v_70115;
wire v_70116;
wire v_70117;
wire v_70118;
wire v_70119;
wire v_70120;
wire v_70121;
wire v_70122;
wire v_70123;
wire v_70124;
wire v_70125;
wire v_70126;
wire v_70127;
wire v_70128;
wire v_70129;
wire v_70130;
wire v_70131;
wire v_70132;
wire v_70133;
wire v_70134;
wire v_70135;
wire v_70136;
wire v_70137;
wire v_70138;
wire v_70139;
wire v_70140;
wire v_70141;
wire v_70142;
wire v_70143;
wire v_70144;
wire v_70145;
wire v_70146;
wire v_70147;
wire v_70148;
wire v_70149;
wire v_70150;
wire v_70151;
wire v_70152;
wire v_70153;
wire v_70154;
wire v_70155;
wire v_70156;
wire v_70157;
wire v_70158;
wire v_70159;
wire v_70160;
wire v_70161;
wire v_70162;
wire v_70163;
wire v_70164;
wire v_70165;
wire v_70166;
wire v_70167;
wire v_70168;
wire v_70169;
wire v_70170;
wire v_70171;
wire v_70172;
wire v_70173;
wire v_70174;
wire v_70175;
wire v_70176;
wire v_70177;
wire v_70178;
wire v_70179;
wire v_70180;
wire v_70181;
wire v_70182;
wire v_70183;
wire v_70184;
wire v_70185;
wire v_70186;
wire v_70187;
wire v_70188;
wire v_70189;
wire v_70190;
wire v_70191;
wire v_70192;
wire v_70193;
wire v_70194;
wire v_70195;
wire v_70196;
wire v_70197;
wire v_70198;
wire v_70199;
wire v_70200;
wire v_70201;
wire v_70202;
wire v_70203;
wire v_70204;
wire v_70205;
wire v_70206;
wire v_70207;
wire v_70208;
wire v_70209;
wire v_70210;
wire v_70211;
wire v_70212;
wire v_70213;
wire v_70214;
wire v_70215;
wire v_70216;
wire v_70217;
wire v_70218;
wire v_70219;
wire v_70220;
wire v_70221;
wire v_70222;
wire v_70223;
wire v_70224;
wire v_70225;
wire v_70226;
wire v_70227;
wire v_70228;
wire v_70229;
wire v_70231;
wire v_70232;
wire v_70233;
wire v_70234;
wire v_70235;
wire v_70236;
wire v_70237;
wire v_70238;
wire v_70239;
wire v_70240;
wire v_70241;
wire v_70242;
wire v_70243;
wire v_70244;
wire v_70245;
wire v_70246;
wire v_70247;
wire v_70248;
wire v_70249;
wire v_70250;
wire v_70251;
wire v_70252;
wire v_70253;
wire v_70254;
wire v_70255;
wire v_70256;
wire v_70257;
wire v_70258;
wire v_70259;
wire v_70260;
wire v_70261;
wire v_70262;
wire v_70263;
wire v_70264;
wire v_70265;
wire v_70266;
wire v_70267;
wire v_70268;
wire v_70269;
wire v_70270;
wire v_70271;
wire v_70272;
wire v_70273;
wire v_70274;
wire v_70275;
wire v_70276;
wire v_70277;
wire v_70278;
wire v_70279;
wire v_70280;
wire v_70281;
wire v_70282;
wire v_70283;
wire v_70284;
wire v_70285;
wire v_70286;
wire v_70287;
wire v_70288;
wire v_70289;
wire v_70290;
wire v_70291;
wire v_70292;
wire v_70293;
wire v_70294;
wire v_70295;
wire v_70296;
wire v_70297;
wire v_70298;
wire v_70299;
wire v_70300;
wire v_70301;
wire v_70302;
wire v_70303;
wire v_70304;
wire v_70305;
wire v_70306;
wire v_70307;
wire v_70308;
wire v_70309;
wire v_70310;
wire v_70311;
wire v_70312;
wire v_70313;
wire v_70314;
wire v_70315;
wire v_70316;
wire v_70317;
wire v_70318;
wire v_70319;
wire v_70320;
wire v_70321;
wire v_70322;
wire v_70323;
wire v_70324;
wire v_70325;
wire v_70326;
wire v_70327;
wire v_70328;
wire v_70329;
wire v_70330;
wire v_70331;
wire v_70332;
wire v_70333;
wire v_70334;
wire v_70335;
wire v_70336;
wire v_70337;
wire v_70338;
wire v_70339;
wire v_70340;
wire v_70341;
wire v_70342;
wire v_70343;
wire v_70344;
wire v_70345;
wire v_70346;
wire v_70347;
wire v_70348;
wire v_70349;
wire v_70350;
wire v_70351;
wire v_70352;
wire v_70353;
wire v_70354;
wire v_70355;
wire v_70356;
wire v_70357;
wire v_70358;
wire v_70359;
wire v_70360;
wire v_70361;
wire v_70362;
wire v_70363;
wire v_70364;
wire v_70365;
wire v_70366;
wire v_70367;
wire v_70368;
wire v_70369;
wire v_70370;
wire v_70371;
wire v_70372;
wire v_70373;
wire v_70374;
wire v_70375;
wire v_70376;
wire v_70377;
wire v_70378;
wire v_70379;
wire v_70380;
wire v_70381;
wire v_70382;
wire v_70383;
wire v_70384;
wire v_70385;
wire v_70386;
wire v_70387;
wire v_70388;
wire v_70389;
wire v_70390;
wire v_70391;
wire v_70392;
wire v_70393;
wire v_70394;
wire v_70395;
wire v_70396;
wire v_70397;
wire v_70398;
wire v_70399;
wire v_70400;
wire v_70401;
wire v_70402;
wire v_70403;
wire v_70404;
wire v_70405;
wire v_70406;
wire v_70407;
wire v_70408;
wire v_70409;
wire v_70410;
wire v_70411;
wire v_70412;
wire v_70413;
wire v_70414;
wire v_70415;
wire v_70416;
wire v_70417;
wire v_70418;
wire v_70419;
wire v_70420;
wire v_70421;
wire v_70422;
wire v_70423;
wire v_70424;
wire v_70425;
wire v_70426;
wire v_70427;
wire v_70428;
wire v_70429;
wire v_70430;
wire v_70431;
wire v_70432;
wire v_70433;
wire v_70434;
wire v_70435;
wire v_70436;
wire v_70437;
wire v_70438;
wire v_70439;
wire v_70440;
wire v_70441;
wire v_70442;
wire v_70443;
wire v_70444;
wire v_70445;
wire v_70446;
wire v_70447;
wire v_70448;
wire v_70449;
wire v_70450;
wire v_70451;
wire v_70452;
wire v_70453;
wire v_70454;
wire v_70455;
wire v_70456;
wire v_70457;
wire v_70458;
wire v_70459;
wire v_70460;
wire v_70461;
wire v_70462;
wire v_70463;
wire v_70464;
wire v_70465;
wire v_70466;
wire v_70467;
wire v_70468;
wire v_70469;
wire v_70470;
wire v_70471;
wire v_70472;
wire v_70474;
wire v_70475;
wire v_70476;
wire v_70477;
wire v_70478;
wire v_70479;
wire v_70480;
wire v_70481;
wire v_70482;
wire v_70483;
wire v_70484;
wire v_70485;
wire v_70486;
wire v_70487;
wire v_70488;
wire v_70489;
wire v_70490;
wire v_70491;
wire v_70492;
wire v_70493;
wire v_70494;
wire v_70495;
wire v_70496;
wire v_70497;
wire v_70498;
wire v_70499;
wire v_70500;
wire v_70501;
wire v_70502;
wire v_70503;
wire v_70504;
wire v_70505;
wire v_70506;
wire v_70507;
wire v_70508;
wire v_70509;
wire v_70510;
wire v_70511;
wire v_70512;
wire v_70513;
wire v_70514;
wire v_70515;
wire v_70516;
wire v_70517;
wire v_70518;
wire v_70519;
wire v_70520;
wire v_70521;
wire v_70522;
wire v_70523;
wire v_70524;
wire v_70525;
wire v_70526;
wire v_70527;
wire v_70528;
wire v_70529;
wire v_70530;
wire v_70531;
wire v_70532;
wire v_70533;
wire v_70534;
wire v_70535;
wire v_70536;
wire v_70537;
wire v_70538;
wire v_70539;
wire v_70540;
wire v_70541;
wire v_70542;
wire v_70543;
wire v_70544;
wire v_70545;
wire v_70546;
wire v_70547;
wire v_70548;
wire v_70549;
wire v_70550;
wire v_70551;
wire v_70552;
wire v_70553;
wire v_70554;
wire v_70555;
wire v_70556;
wire v_70557;
wire v_70558;
wire v_70559;
wire v_70560;
wire v_70561;
wire v_70562;
wire v_70563;
wire v_70564;
wire v_70565;
wire v_70566;
wire v_70567;
wire v_70568;
wire v_70569;
wire v_70570;
wire v_70571;
wire v_70572;
wire v_70573;
wire v_70574;
wire v_70575;
wire v_70576;
wire v_70577;
wire v_70578;
wire v_70579;
wire v_70580;
wire v_70581;
wire v_70582;
wire v_70583;
wire v_70584;
wire v_70585;
wire v_70586;
wire v_70587;
wire v_70588;
wire v_70589;
wire v_70590;
wire v_70591;
wire v_70592;
wire v_70593;
wire v_70594;
wire v_70595;
wire v_70596;
wire v_70597;
wire v_70598;
wire v_70599;
wire v_70600;
wire v_70601;
wire v_70602;
wire v_70603;
wire v_70604;
wire v_70605;
wire v_70606;
wire v_70607;
wire v_70608;
wire v_70609;
wire v_70610;
wire v_70611;
wire v_70612;
wire v_70613;
wire v_70614;
wire v_70615;
wire v_70616;
wire v_70617;
wire v_70618;
wire v_70619;
wire v_70620;
wire v_70621;
wire v_70622;
wire v_70623;
wire v_70624;
wire v_70625;
wire v_70626;
wire v_70627;
wire v_70628;
wire v_70629;
wire v_70630;
wire v_70631;
wire v_70632;
wire v_70633;
wire v_70634;
wire v_70635;
wire v_70636;
wire v_70637;
wire v_70638;
wire v_70639;
wire v_70640;
wire v_70641;
wire v_70642;
wire v_70643;
wire v_70644;
wire v_70645;
wire v_70646;
wire v_70647;
wire v_70648;
wire v_70649;
wire v_70650;
wire v_70651;
wire v_70652;
wire v_70653;
wire v_70654;
wire v_70655;
wire v_70656;
wire v_70657;
wire v_70658;
wire v_70659;
wire v_70660;
wire v_70661;
wire v_70662;
wire v_70663;
wire v_70664;
wire v_70665;
wire v_70666;
wire v_70667;
wire v_70668;
wire v_70669;
wire v_70670;
wire v_70671;
wire v_70672;
wire v_70673;
wire v_70674;
wire v_70675;
wire v_70676;
wire v_70677;
wire v_70678;
wire v_70679;
wire v_70680;
wire v_70681;
wire v_70682;
wire v_70683;
wire v_70684;
wire v_70685;
wire v_70686;
wire v_70687;
wire v_70688;
wire v_70689;
wire v_70690;
wire v_70691;
wire v_70692;
wire v_70693;
wire v_70694;
wire v_70695;
wire v_70696;
wire v_70697;
wire v_70698;
wire v_70699;
wire v_70700;
wire v_70701;
wire v_70702;
wire v_70703;
wire v_70704;
wire v_70705;
wire v_70706;
wire v_70707;
wire v_70708;
wire v_70709;
wire v_70710;
wire v_70711;
wire v_70712;
wire v_70713;
wire v_70714;
wire v_70715;
wire v_70717;
wire v_70718;
wire v_70719;
wire v_70720;
wire v_70721;
wire v_70722;
wire v_70723;
wire v_70724;
wire v_70725;
wire v_70726;
wire v_70727;
wire v_70728;
wire v_70729;
wire v_70730;
wire v_70731;
wire v_70732;
wire v_70733;
wire v_70734;
wire v_70735;
wire v_70736;
wire v_70737;
wire v_70738;
wire v_70739;
wire v_70740;
wire v_70741;
wire v_70742;
wire v_70743;
wire v_70744;
wire v_70745;
wire v_70746;
wire v_70747;
wire v_70748;
wire v_70749;
wire v_70750;
wire v_70751;
wire v_70752;
wire v_70753;
wire v_70754;
wire v_70755;
wire v_70756;
wire v_70757;
wire v_70758;
wire v_70759;
wire v_70760;
wire v_70761;
wire v_70762;
wire v_70763;
wire v_70764;
wire v_70765;
wire v_70766;
wire v_70767;
wire v_70768;
wire v_70769;
wire v_70770;
wire v_70771;
wire v_70772;
wire v_70773;
wire v_70774;
wire v_70775;
wire v_70776;
wire v_70777;
wire v_70778;
wire v_70779;
wire v_70780;
wire v_70781;
wire v_70782;
wire v_70783;
wire v_70784;
wire v_70785;
wire v_70786;
wire v_70787;
wire v_70788;
wire v_70789;
wire v_70790;
wire v_70791;
wire v_70792;
wire v_70793;
wire v_70794;
wire v_70795;
wire v_70796;
wire v_70797;
wire v_70798;
wire v_70799;
wire v_70800;
wire v_70801;
wire v_70802;
wire v_70803;
wire v_70804;
wire v_70805;
wire v_70806;
wire v_70807;
wire v_70808;
wire v_70809;
wire v_70810;
wire v_70811;
wire v_70812;
wire v_70813;
wire v_70814;
wire v_70815;
wire v_70816;
wire v_70817;
wire v_70818;
wire v_70819;
wire v_70820;
wire v_70821;
wire v_70822;
wire v_70823;
wire v_70824;
wire v_70825;
wire v_70826;
wire v_70827;
wire v_70828;
wire v_70829;
wire v_70830;
wire v_70831;
wire v_70832;
wire v_70833;
wire v_70834;
wire v_70835;
wire v_70836;
wire v_70837;
wire v_70838;
wire v_70839;
wire v_70840;
wire v_70841;
wire v_70842;
wire v_70843;
wire v_70844;
wire v_70845;
wire v_70846;
wire v_70847;
wire v_70848;
wire v_70849;
wire v_70850;
wire v_70851;
wire v_70852;
wire v_70853;
wire v_70854;
wire v_70855;
wire v_70856;
wire v_70857;
wire v_70858;
wire v_70859;
wire v_70860;
wire v_70861;
wire v_70862;
wire v_70863;
wire v_70864;
wire v_70865;
wire v_70866;
wire v_70867;
wire v_70868;
wire v_70869;
wire v_70870;
wire v_70871;
wire v_70872;
wire v_70873;
wire v_70874;
wire v_70875;
wire v_70876;
wire v_70877;
wire v_70878;
wire v_70879;
wire v_70880;
wire v_70881;
wire v_70882;
wire v_70883;
wire v_70884;
wire v_70885;
wire v_70886;
wire v_70887;
wire v_70888;
wire v_70889;
wire v_70890;
wire v_70891;
wire v_70892;
wire v_70893;
wire v_70894;
wire v_70895;
wire v_70896;
wire v_70897;
wire v_70898;
wire v_70899;
wire v_70900;
wire v_70901;
wire v_70902;
wire v_70903;
wire v_70904;
wire v_70905;
wire v_70906;
wire v_70907;
wire v_70908;
wire v_70909;
wire v_70910;
wire v_70911;
wire v_70912;
wire v_70913;
wire v_70914;
wire v_70915;
wire v_70916;
wire v_70917;
wire v_70918;
wire v_70919;
wire v_70920;
wire v_70921;
wire v_70922;
wire v_70923;
wire v_70924;
wire v_70925;
wire v_70926;
wire v_70927;
wire v_70928;
wire v_70929;
wire v_70930;
wire v_70931;
wire v_70932;
wire v_70933;
wire v_70934;
wire v_70935;
wire v_70936;
wire v_70937;
wire v_70938;
wire v_70939;
wire v_70940;
wire v_70941;
wire v_70942;
wire v_70943;
wire v_70944;
wire v_70945;
wire v_70946;
wire v_70947;
wire v_70948;
wire v_70949;
wire v_70950;
wire v_70951;
wire v_70952;
wire v_70953;
wire v_70954;
wire v_70955;
wire v_70956;
wire v_70957;
wire v_70958;
wire v_70959;
wire v_70960;
wire v_70961;
wire v_70962;
wire v_70963;
wire v_70964;
wire v_70965;
wire v_70966;
wire v_70967;
wire v_70968;
wire v_70969;
wire v_70970;
wire v_70971;
wire v_70972;
wire v_70973;
wire v_70974;
wire v_70975;
wire v_70976;
wire v_70977;
wire v_70978;
wire v_70979;
wire v_70980;
wire v_70981;
wire v_70982;
wire v_70983;
wire v_70984;
wire v_70985;
wire v_70986;
wire v_70987;
wire v_70988;
wire v_70989;
wire v_70990;
wire v_70991;
wire v_70992;
wire v_70993;
wire v_70994;
wire v_70995;
wire v_70996;
wire v_70997;
wire v_70998;
wire v_70999;
wire v_71000;
wire v_71001;
wire v_71002;
wire v_71003;
wire v_71004;
wire v_71005;
wire v_71006;
wire v_71007;
wire v_71008;
wire v_71009;
wire v_71010;
wire v_71011;
wire v_71012;
wire v_71013;
wire v_71014;
wire v_71015;
wire v_71016;
wire v_71017;
wire v_71018;
wire v_71019;
wire v_71020;
wire v_71021;
wire v_71022;
wire v_71023;
wire v_71024;
wire v_71025;
wire v_71026;
wire v_71027;
wire v_71028;
wire v_71029;
wire v_71030;
wire v_71031;
wire v_71032;
wire v_71033;
wire v_71034;
wire v_71035;
wire v_71036;
wire v_71037;
wire v_71038;
wire v_71039;
wire v_71040;
wire v_71041;
wire v_71042;
wire v_71043;
wire v_71044;
wire v_71045;
wire v_71046;
wire v_71047;
wire v_71048;
wire v_71049;
wire v_71050;
wire v_71051;
wire v_71052;
wire v_71053;
wire v_71054;
wire v_71055;
wire v_71056;
wire v_71057;
wire v_71058;
wire v_71059;
wire v_71060;
wire v_71061;
wire v_71062;
wire v_71063;
wire v_71064;
wire v_71065;
wire v_71066;
wire v_71067;
wire v_71068;
wire v_71069;
wire v_71070;
wire v_71071;
wire v_71072;
wire v_71073;
wire v_71074;
wire v_71075;
wire v_71076;
wire v_71077;
wire v_71078;
wire v_71079;
wire v_71080;
wire v_71081;
wire v_71082;
wire v_71083;
wire v_71084;
wire v_71085;
wire v_71086;
wire v_71087;
wire v_71088;
wire v_71089;
wire v_71090;
wire v_71091;
wire v_71092;
wire v_71093;
wire v_71094;
wire v_71095;
wire v_71096;
wire v_71097;
wire v_71098;
wire v_71099;
wire v_71100;
wire v_71101;
wire v_71102;
wire v_71103;
wire v_71104;
wire v_71105;
wire v_71106;
wire v_71107;
wire v_71108;
wire v_71109;
wire v_71110;
wire v_71111;
wire v_71112;
wire v_71113;
wire v_71114;
wire v_71115;
wire v_71116;
wire v_71117;
wire v_71118;
wire v_71119;
wire v_71120;
wire v_71121;
wire v_71122;
wire v_71123;
wire v_71124;
wire v_71125;
wire v_71126;
wire v_71127;
wire v_71128;
wire v_71129;
wire v_71130;
wire v_71131;
wire v_71132;
wire v_71133;
wire v_71134;
wire v_71135;
wire v_71136;
wire v_71137;
wire v_71138;
wire v_71139;
wire v_71140;
wire v_71141;
wire v_71142;
wire v_71143;
wire v_71144;
wire v_71145;
wire v_71146;
wire v_71147;
wire v_71148;
wire v_71149;
wire v_71150;
wire v_71151;
wire v_71152;
wire v_71153;
wire v_71154;
wire v_71155;
wire v_71156;
wire v_71157;
wire v_71158;
wire v_71159;
wire v_71160;
wire v_71161;
wire v_71162;
wire v_71163;
wire v_71164;
wire v_71165;
wire v_71166;
wire v_71167;
wire v_71168;
wire v_71169;
wire v_71170;
wire v_71171;
wire v_71172;
wire v_71173;
wire v_71174;
wire v_71175;
wire v_71176;
wire v_71177;
wire v_71178;
wire v_71179;
wire v_71180;
wire v_71181;
wire v_71182;
wire v_71183;
wire v_71184;
wire v_71185;
wire v_71186;
wire v_71187;
wire v_71188;
wire v_71189;
wire v_71190;
wire v_71191;
wire v_71192;
wire v_71193;
wire v_71194;
wire v_71195;
wire v_71196;
wire v_71197;
wire v_71198;
wire v_71199;
wire v_71200;
wire v_71201;
wire v_71202;
wire v_71203;
wire v_71204;
wire v_71205;
wire v_71206;
wire v_71207;
wire v_71208;
wire v_71209;
wire v_71210;
wire v_71211;
wire v_71212;
wire v_71213;
wire v_71214;
wire v_71215;
wire v_71216;
wire v_71217;
wire v_71218;
wire v_71219;
wire v_71220;
wire v_71221;
wire v_71222;
wire v_71223;
wire v_71224;
wire v_71225;
wire v_71226;
wire v_71227;
wire v_71228;
wire v_71229;
wire v_71230;
wire v_71231;
wire v_71232;
wire v_71233;
wire v_71234;
wire v_71235;
wire v_71236;
wire v_71237;
wire v_71238;
wire v_71239;
wire v_71240;
wire v_71241;
wire v_71242;
wire v_71243;
wire v_71244;
wire v_71245;
wire v_71246;
wire v_71247;
wire v_71248;
wire v_71249;
wire v_71250;
wire v_71251;
wire v_71252;
wire v_71253;
wire v_71254;
wire v_71255;
wire v_71256;
wire v_71257;
wire v_71258;
wire v_71259;
wire v_71260;
wire v_71261;
wire v_71262;
wire v_71263;
wire v_71264;
wire v_71265;
wire v_71266;
wire v_71267;
wire v_71268;
wire v_71269;
wire v_71270;
wire v_71271;
wire v_71272;
wire v_71273;
wire v_71274;
wire v_71275;
wire v_71276;
wire v_71277;
wire v_71278;
wire v_71279;
wire v_71280;
wire v_71281;
wire v_71282;
wire v_71283;
wire v_71284;
wire v_71285;
wire v_71286;
wire v_71287;
wire v_71288;
wire v_71289;
wire v_71290;
wire v_71291;
wire v_71292;
wire v_71293;
wire v_71294;
wire v_71295;
wire v_71296;
wire v_71297;
wire v_71298;
wire v_71299;
wire v_71300;
wire v_71301;
wire v_71302;
wire v_71303;
wire v_71304;
wire v_71305;
wire v_71306;
wire v_71307;
wire v_71308;
wire v_71309;
wire v_71310;
wire v_71311;
wire v_71312;
wire v_71313;
wire v_71314;
wire v_71315;
wire v_71316;
wire v_71317;
wire v_71318;
wire v_71319;
wire v_71320;
wire v_71321;
wire v_71322;
wire v_71323;
wire v_71324;
wire v_71325;
wire v_71326;
wire v_71327;
wire v_71328;
wire v_71329;
wire v_71330;
wire v_71331;
wire v_71332;
wire v_71333;
wire v_71334;
wire v_71335;
wire v_71336;
wire v_71337;
wire v_71338;
wire v_71339;
wire v_71340;
wire v_71341;
wire v_71342;
wire v_71343;
wire v_71344;
wire v_71345;
wire v_71346;
wire v_71347;
wire v_71348;
wire v_71349;
wire v_71350;
wire v_71351;
wire v_71352;
wire v_71353;
wire v_71354;
wire v_71355;
wire v_71356;
wire v_71357;
wire v_71358;
wire v_71359;
wire v_71360;
wire v_71361;
wire v_71362;
wire v_71363;
wire v_71364;
wire v_71365;
wire v_71366;
wire v_71367;
wire v_71368;
wire v_71369;
wire v_71370;
wire v_71371;
wire v_71372;
wire v_71373;
wire v_71374;
wire v_71375;
wire v_71376;
wire v_71377;
wire v_71378;
wire v_71379;
wire v_71380;
wire v_71381;
wire v_71382;
wire v_71383;
wire v_71384;
wire v_71385;
wire v_71386;
wire v_71387;
wire v_71388;
wire v_71389;
wire v_71390;
wire v_71391;
wire v_71392;
wire v_71393;
wire v_71394;
wire v_71395;
wire v_71396;
wire v_71397;
wire v_71398;
wire v_71399;
wire v_71400;
wire v_71401;
wire v_71402;
wire v_71403;
wire v_71404;
wire v_71405;
wire v_71406;
wire v_71407;
wire v_71408;
wire v_71409;
wire v_71410;
wire v_71411;
wire v_71412;
wire v_71413;
wire v_71414;
wire v_71415;
wire v_71416;
wire v_71417;
wire v_71418;
wire v_71419;
wire v_71420;
wire v_71421;
wire v_71422;
wire v_71423;
wire v_71424;
wire v_71425;
wire v_71426;
wire v_71427;
wire v_71428;
wire v_71429;
wire v_71430;
wire v_71431;
wire v_71432;
wire v_71433;
wire v_71434;
wire v_71435;
wire v_71436;
wire v_71437;
wire v_71438;
wire v_71439;
wire v_71440;
wire v_71441;
wire v_71442;
wire v_71443;
wire v_71444;
wire v_71445;
wire v_71446;
wire v_71447;
wire v_71448;
wire v_71449;
wire v_71450;
wire v_71451;
wire v_71452;
wire v_71453;
wire v_71454;
wire v_71455;
wire v_71456;
wire v_71457;
wire v_71458;
wire v_71459;
wire v_71460;
wire v_71461;
wire v_71462;
wire v_71463;
wire v_71464;
wire v_71465;
wire v_71466;
wire v_71467;
wire v_71468;
wire v_71469;
wire v_71470;
wire v_71471;
wire v_71472;
wire v_71473;
wire v_71474;
wire v_71475;
wire v_71476;
wire v_71477;
wire v_71478;
wire v_71479;
wire v_71480;
wire v_71481;
wire v_71482;
wire v_71483;
wire v_71484;
wire v_71485;
wire v_71486;
wire v_71487;
wire v_71488;
wire v_71489;
wire v_71490;
wire v_71491;
wire v_71492;
wire v_71493;
wire v_71494;
wire v_71495;
wire v_71496;
wire v_71497;
wire v_71498;
wire v_71499;
wire v_71500;
wire v_71501;
wire v_71502;
wire v_71503;
wire v_71504;
wire v_71505;
wire v_71506;
wire v_71507;
wire v_71508;
wire v_71509;
wire v_71510;
wire v_71511;
wire v_71512;
wire v_71513;
wire v_71514;
wire v_71515;
wire v_71516;
wire v_71517;
wire v_71518;
wire v_71519;
wire v_71520;
wire v_71521;
wire v_71522;
wire v_71523;
wire v_71524;
wire v_71525;
wire v_71526;
wire v_71527;
wire v_71528;
wire v_71529;
wire v_71530;
wire v_71531;
wire v_71532;
wire v_71533;
wire v_71534;
wire v_71535;
wire v_71536;
wire v_71537;
wire v_71538;
wire v_71539;
wire v_71540;
wire v_71541;
wire v_71542;
wire v_71543;
wire v_71544;
wire v_71545;
wire v_71546;
wire v_71547;
wire v_71548;
wire v_71549;
wire v_71550;
wire v_71551;
wire v_71552;
wire v_71553;
wire v_71554;
wire v_71555;
wire v_71556;
wire v_71557;
wire v_71558;
wire v_71559;
wire v_71560;
wire v_71561;
wire v_71562;
wire v_71563;
wire v_71564;
wire v_71565;
wire v_71566;
wire v_71567;
wire v_71568;
wire v_71569;
wire v_71570;
wire v_71571;
wire v_71572;
wire v_71573;
wire v_71574;
wire v_71575;
wire v_71576;
wire v_71577;
wire v_71578;
wire v_71579;
wire v_71580;
wire v_71581;
wire v_71582;
wire v_71583;
wire v_71584;
wire v_71585;
wire v_71586;
wire v_71587;
wire v_71588;
wire v_71589;
wire v_71590;
wire v_71591;
wire v_71592;
wire v_71593;
wire v_71594;
wire v_71595;
wire v_71596;
wire v_71597;
wire v_71598;
wire v_71599;
wire v_71600;
wire v_71601;
wire v_71602;
wire v_71603;
wire v_71604;
wire v_71605;
wire v_71606;
wire v_71607;
wire v_71608;
wire v_71609;
wire v_71610;
wire v_71611;
wire v_71612;
wire v_71613;
wire v_71614;
wire v_71615;
wire v_71616;
wire v_71617;
wire v_71618;
wire v_71619;
wire v_71620;
wire v_71621;
wire v_71622;
wire v_71623;
wire v_71624;
wire v_71625;
wire v_71626;
wire v_71627;
wire v_71628;
wire v_71629;
wire v_71630;
wire v_71631;
wire v_71632;
wire v_71633;
wire v_71634;
wire v_71635;
wire v_71636;
wire v_71637;
wire v_71638;
wire v_71639;
wire v_71640;
wire v_71641;
wire v_71642;
wire v_71643;
wire v_71644;
wire v_71645;
wire v_71646;
wire v_71647;
wire v_71648;
wire v_71649;
wire v_71650;
wire v_71651;
wire v_71652;
wire v_71653;
wire v_71654;
wire v_71655;
wire v_71656;
wire v_71657;
wire v_71658;
wire v_71659;
wire v_71660;
wire v_71661;
wire v_71662;
wire v_71663;
wire v_71664;
wire v_71665;
wire v_71666;
wire v_71667;
wire v_71668;
wire v_71669;
wire v_71670;
wire v_71671;
wire v_71672;
wire v_71673;
wire v_71674;
wire v_71675;
wire v_71676;
wire v_71677;
wire v_71678;
wire v_71679;
wire v_71680;
wire v_71681;
wire v_71682;
wire v_71683;
wire v_71684;
wire v_71685;
wire v_71686;
wire v_71687;
wire v_71688;
wire v_71689;
wire v_71690;
wire v_71691;
wire v_71692;
wire v_71693;
wire v_71694;
wire v_71695;
wire v_71696;
wire v_71697;
wire v_71698;
wire v_71699;
wire v_71700;
wire v_71701;
wire v_71702;
wire v_71703;
wire v_71704;
wire v_71705;
wire v_71706;
wire v_71707;
wire v_71708;
wire v_71709;
wire v_71710;
wire v_71711;
wire v_71712;
wire v_71713;
wire v_71714;
wire v_71715;
wire v_71716;
wire v_71717;
wire v_71718;
wire v_71719;
wire v_71720;
wire v_71721;
wire v_71722;
wire v_71723;
wire v_71724;
wire v_71725;
wire v_71726;
wire v_71727;
wire v_71728;
wire v_71729;
wire v_71730;
wire v_71731;
wire v_71732;
wire v_71733;
wire v_71734;
wire v_71735;
wire v_71736;
wire v_71737;
wire v_71738;
wire v_71739;
wire v_71740;
wire v_71741;
wire v_71742;
wire v_71743;
wire v_71744;
wire v_71745;
wire v_71746;
wire v_71747;
wire v_71748;
wire v_71749;
wire v_71750;
wire v_71751;
wire v_71752;
wire v_71753;
wire v_71754;
wire v_71755;
wire v_71756;
wire v_71757;
wire v_71758;
wire v_71759;
wire v_71760;
wire v_71761;
wire v_71762;
wire v_71763;
wire v_71764;
wire v_71765;
wire v_71766;
wire v_71767;
wire v_71768;
wire v_71769;
wire v_71770;
wire v_71771;
wire v_71772;
wire v_71773;
wire v_71774;
wire v_71775;
wire v_71776;
wire v_71777;
wire v_71778;
wire v_71779;
wire v_71780;
wire v_71781;
wire v_71782;
wire v_71783;
wire v_71784;
wire v_71785;
wire v_71786;
wire v_71787;
wire v_71788;
wire v_71789;
wire v_71790;
wire v_71791;
wire v_71792;
wire v_71793;
wire v_71794;
wire v_71795;
wire v_71796;
wire v_71797;
wire v_71798;
wire v_71799;
wire v_71800;
wire v_71801;
wire v_71802;
wire v_71803;
wire v_71804;
wire v_71805;
wire v_71806;
wire v_71807;
wire v_71808;
wire v_71809;
wire v_71810;
wire v_71811;
wire v_71812;
wire v_71813;
wire v_71814;
wire v_71815;
wire v_71816;
wire v_71817;
wire v_71818;
wire v_71819;
wire v_71820;
wire v_71821;
wire v_71822;
wire v_71823;
wire v_71824;
wire v_71825;
wire v_71826;
wire v_71827;
wire v_71828;
wire v_71829;
wire v_71830;
wire v_71831;
wire v_71832;
wire v_71833;
wire v_71834;
wire v_71835;
wire v_71836;
wire v_71837;
wire v_71838;
wire v_71839;
wire v_71840;
wire v_71841;
wire v_71842;
wire v_71843;
wire v_71844;
wire v_71845;
wire v_71846;
wire v_71847;
wire v_71848;
wire v_71849;
wire v_71850;
wire v_71851;
wire v_71852;
wire v_71853;
wire v_71854;
wire v_71855;
wire v_71856;
wire v_71857;
wire v_71858;
wire v_71859;
wire v_71860;
wire v_71861;
wire v_71862;
wire v_71863;
wire v_71864;
wire v_71865;
wire v_71866;
wire v_71867;
wire v_71868;
wire v_71869;
wire v_71870;
wire v_71871;
wire v_71872;
wire v_71873;
wire v_71874;
wire v_71875;
wire v_71876;
wire v_71877;
wire v_71878;
wire v_71879;
wire v_71880;
wire v_71881;
wire v_71882;
wire v_71883;
wire v_71884;
wire v_71885;
wire v_71886;
wire v_71887;
wire v_71888;
wire v_71889;
wire v_71890;
wire v_71891;
wire v_71892;
wire v_71893;
wire v_71894;
wire v_71895;
wire v_71896;
wire v_71897;
wire v_71898;
wire v_71899;
wire v_71900;
wire v_71901;
wire v_71902;
wire v_71903;
wire v_71904;
wire v_71905;
wire v_71906;
wire v_71907;
wire v_71908;
wire v_71909;
wire v_71910;
wire v_71911;
wire v_71912;
wire v_71913;
wire v_71914;
wire v_71915;
wire v_71916;
wire v_71917;
wire v_71918;
wire v_71919;
wire v_71920;
wire v_71921;
wire v_71922;
wire v_71923;
wire v_71924;
wire v_71925;
wire v_71926;
wire v_71927;
wire v_71928;
wire v_71929;
wire v_71930;
wire v_71931;
wire v_71932;
wire v_71933;
wire v_71934;
wire v_71935;
wire v_71936;
wire v_71937;
wire v_71938;
wire v_71939;
wire v_71940;
wire v_71941;
wire v_71942;
wire v_71943;
wire v_71944;
wire v_71945;
wire v_71946;
wire v_71947;
wire v_71948;
wire v_71949;
wire v_71950;
wire v_71951;
wire v_71952;
wire v_71953;
wire v_71954;
wire v_71955;
wire v_71956;
wire v_71957;
wire v_71958;
wire v_71959;
wire v_71960;
wire v_71961;
wire v_71962;
wire v_71963;
wire v_71964;
wire v_71965;
wire v_71966;
wire v_71967;
wire v_71968;
wire v_71969;
wire v_71970;
wire v_71971;
wire v_71972;
wire v_71973;
wire v_71974;
wire v_71975;
wire v_71976;
wire v_71977;
wire v_71978;
wire v_71979;
wire v_71980;
wire v_71981;
wire v_71982;
wire v_71983;
wire v_71984;
wire v_71985;
wire v_71986;
wire v_71987;
wire v_71988;
wire v_71989;
wire v_71990;
wire v_71991;
wire v_71992;
wire v_71993;
wire v_71994;
wire v_71995;
wire v_71996;
wire v_71997;
wire v_71998;
wire v_71999;
wire v_72000;
wire v_72001;
wire v_72002;
wire v_72003;
wire v_72004;
wire v_72005;
wire v_72006;
wire v_72007;
wire v_72008;
wire v_72009;
wire v_72010;
wire v_72011;
wire v_72012;
wire v_72013;
wire v_72014;
wire v_72015;
wire v_72016;
wire v_72017;
wire v_72018;
wire v_72019;
wire v_72020;
wire v_72021;
wire v_72022;
wire v_72023;
wire v_72024;
wire v_72025;
wire v_72026;
wire v_72027;
wire v_72028;
wire v_72029;
wire v_72030;
wire v_72031;
wire v_72032;
wire v_72033;
wire v_72034;
wire v_72035;
wire v_72036;
wire v_72037;
wire v_72038;
wire v_72039;
wire v_72040;
wire v_72041;
wire v_72042;
wire v_72043;
wire v_72044;
wire v_72045;
wire v_72046;
wire v_72047;
wire v_72048;
wire v_72049;
wire v_72050;
wire v_72051;
wire v_72052;
wire v_72053;
wire v_72054;
wire v_72055;
wire v_72056;
wire v_72057;
wire v_72058;
wire v_72059;
wire v_72060;
wire v_72061;
wire v_72062;
wire v_72063;
wire v_72064;
wire v_72065;
wire v_72066;
wire v_72067;
wire v_72068;
wire v_72069;
wire v_72070;
wire v_72071;
wire v_72072;
wire v_72073;
wire v_72074;
wire v_72075;
wire v_72076;
wire v_72077;
wire v_72078;
wire v_72079;
wire v_72080;
wire v_72081;
wire v_72082;
wire v_72083;
wire v_72084;
wire v_72085;
wire v_72086;
wire v_72087;
wire v_72088;
wire v_72089;
wire v_72090;
wire v_72091;
wire v_72092;
wire v_72093;
wire v_72094;
wire v_72095;
wire v_72096;
wire v_72097;
wire v_72098;
wire v_72099;
wire v_72100;
wire v_72101;
wire v_72102;
wire v_72103;
wire v_72104;
wire v_72105;
wire v_72106;
wire v_72107;
wire v_72108;
wire v_72109;
wire v_72110;
wire v_72111;
wire v_72112;
wire v_72113;
wire v_72114;
wire v_72115;
wire v_72116;
wire v_72117;
wire v_72118;
wire v_72119;
wire v_72120;
wire v_72121;
wire v_72122;
wire v_72123;
wire v_72124;
wire v_72125;
wire v_72126;
wire v_72127;
wire v_72128;
wire v_72129;
wire v_72130;
wire v_72131;
wire v_72132;
wire v_72133;
wire v_72134;
wire v_72135;
wire v_72136;
wire v_72137;
wire v_72138;
wire v_72139;
wire v_72140;
wire v_72141;
wire v_72142;
wire v_72143;
wire v_72144;
wire v_72145;
wire v_72146;
wire v_72147;
wire v_72148;
wire v_72149;
wire v_72150;
wire v_72151;
wire v_72152;
wire v_72153;
wire v_72154;
wire v_72155;
wire v_72156;
wire v_72157;
wire v_72158;
wire v_72159;
wire v_72160;
wire v_72161;
wire v_72162;
wire v_72163;
wire v_72164;
wire v_72165;
wire v_72166;
wire v_72167;
wire v_72168;
wire v_72169;
wire v_72170;
wire v_72171;
wire v_72172;
wire v_72173;
wire v_72174;
wire v_72175;
wire v_72176;
wire v_72177;
wire v_72178;
wire v_72179;
wire v_72180;
wire v_72181;
wire v_72182;
wire v_72183;
wire v_72184;
wire v_72185;
wire v_72186;
wire v_72187;
wire v_72188;
wire v_72189;
wire v_72190;
wire v_72191;
wire v_72192;
wire v_72193;
wire v_72194;
wire v_72195;
wire v_72196;
wire v_72197;
wire v_72198;
wire v_72199;
wire v_72200;
wire v_72201;
wire v_72202;
wire v_72203;
wire v_72204;
wire v_72205;
wire v_72206;
wire v_72207;
wire v_72208;
wire v_72209;
wire v_72210;
wire v_72211;
wire v_72212;
wire v_72213;
wire v_72214;
wire v_72215;
wire v_72216;
wire v_72217;
wire v_72218;
wire v_72219;
wire v_72220;
wire v_72221;
wire v_72222;
wire v_72223;
wire v_72224;
wire v_72225;
wire v_72226;
wire v_72227;
wire v_72228;
wire v_72229;
wire v_72230;
wire v_72231;
wire v_72232;
wire v_72233;
wire v_72234;
wire v_72235;
wire v_72236;
wire v_72237;
wire v_72238;
wire v_72239;
wire v_72240;
wire v_72241;
wire v_72242;
wire v_72243;
wire v_72244;
wire v_72245;
wire v_72246;
wire v_72247;
wire v_72248;
wire v_72249;
wire v_72250;
wire v_72251;
wire v_72252;
wire v_72253;
wire v_72254;
wire v_72255;
wire v_72256;
wire v_72257;
wire v_72258;
wire v_72259;
wire v_72260;
wire v_72261;
wire v_72262;
wire v_72263;
wire v_72264;
wire v_72265;
wire v_72266;
wire v_72267;
wire v_72268;
wire v_72269;
wire v_72270;
wire v_72271;
wire v_72272;
wire v_72273;
wire v_72274;
wire v_72275;
wire v_72276;
wire v_72277;
wire v_72278;
wire v_72279;
wire v_72280;
wire v_72281;
wire v_72282;
wire v_72283;
wire v_72284;
wire v_72285;
wire v_72286;
wire v_72287;
wire v_72288;
wire v_72289;
wire v_72290;
wire v_72291;
wire v_72292;
wire v_72293;
wire v_72294;
wire v_72295;
wire v_72296;
wire v_72297;
wire v_72298;
wire v_72299;
wire v_72300;
wire v_72301;
wire v_72302;
wire v_72303;
wire v_72304;
wire v_72305;
wire v_72306;
wire v_72307;
wire v_72308;
wire v_72309;
wire v_72310;
wire v_72311;
wire v_72312;
wire v_72313;
wire v_72314;
wire v_72315;
wire v_72316;
wire v_72317;
wire v_72318;
wire v_72319;
wire v_72320;
wire v_72321;
wire v_72322;
wire v_72323;
wire v_72324;
wire v_72325;
wire v_72326;
wire v_72327;
wire v_72328;
wire v_72329;
wire v_72330;
wire v_72331;
wire v_72332;
wire v_72333;
wire v_72334;
wire v_72335;
wire v_72336;
wire v_72337;
wire v_72338;
wire v_72339;
wire v_72340;
wire v_72341;
wire v_72342;
wire v_72343;
wire v_72344;
wire v_72345;
wire v_72346;
wire v_72347;
wire v_72348;
wire v_72349;
wire v_72350;
wire v_72351;
wire v_72352;
wire v_72353;
wire v_72354;
wire v_72355;
wire v_72356;
wire v_72357;
wire v_72358;
wire v_72359;
wire v_72360;
wire v_72361;
wire v_72362;
wire v_72363;
wire v_72364;
wire v_72365;
wire v_72366;
wire v_72367;
wire v_72368;
wire v_72369;
wire v_72370;
wire v_72371;
wire v_72372;
wire v_72373;
wire v_72374;
wire v_72375;
wire v_72376;
wire v_72377;
wire v_72378;
wire v_72379;
wire v_72380;
wire v_72381;
wire v_72382;
wire v_72383;
wire v_72384;
wire v_72385;
wire v_72386;
wire v_72387;
wire v_72388;
wire v_72389;
wire v_72390;
wire v_72391;
wire v_72392;
wire v_72393;
wire v_72394;
wire v_72395;
wire v_72396;
wire v_72397;
wire v_72398;
wire v_72399;
wire v_72400;
wire v_72401;
wire v_72402;
wire v_72403;
wire v_72404;
wire v_72405;
wire v_72406;
wire v_72407;
wire v_72408;
wire v_72409;
wire v_72410;
wire v_72411;
wire v_72412;
wire v_72413;
wire v_72414;
wire v_72415;
wire v_72416;
wire v_72417;
wire v_72418;
wire v_72419;
wire v_72420;
wire v_72421;
wire v_72422;
wire v_72423;
wire v_72424;
wire v_72425;
wire v_72426;
wire v_72427;
wire v_72428;
wire v_72429;
wire v_72430;
wire v_72431;
wire v_72432;
wire v_72433;
wire v_72434;
wire v_72435;
wire v_72436;
wire v_72437;
wire v_72438;
wire v_72439;
wire v_72440;
wire v_72441;
wire v_72442;
wire v_72443;
wire v_72444;
wire v_72445;
wire v_72446;
wire v_72447;
wire v_72448;
wire v_72449;
wire v_72450;
wire v_72451;
wire v_72452;
wire v_72453;
wire v_72454;
wire v_72455;
wire v_72456;
wire v_72457;
wire v_72458;
wire v_72459;
wire v_72460;
wire v_72461;
wire v_72462;
wire v_72463;
wire v_72464;
wire v_72465;
wire v_72466;
wire v_72467;
wire v_72468;
wire v_72469;
wire v_72470;
wire v_72471;
wire v_72472;
wire v_72473;
wire v_72474;
wire v_72475;
wire v_72476;
wire v_72477;
wire v_72478;
wire v_72479;
wire v_72480;
wire v_72481;
wire v_72482;
wire v_72483;
wire v_72484;
wire v_72485;
wire v_72486;
wire v_72487;
wire v_72488;
wire v_72489;
wire v_72490;
wire v_72491;
wire v_72492;
wire v_72493;
wire v_72494;
wire v_72495;
wire v_72496;
wire v_72497;
wire v_72498;
wire v_72499;
wire v_72500;
wire v_72501;
wire v_72502;
wire v_72503;
wire v_72504;
wire v_72505;
wire v_72506;
wire v_72507;
wire v_72508;
wire v_72509;
wire v_72510;
wire v_72511;
wire v_72512;
wire v_72513;
wire v_72514;
wire v_72515;
wire v_72516;
wire v_72517;
wire v_72518;
wire v_72519;
wire v_72520;
wire v_72521;
wire v_72522;
wire v_72523;
wire v_72524;
wire v_72525;
wire v_72526;
wire v_72527;
wire v_72528;
wire v_72529;
wire v_72530;
wire v_72531;
wire v_72532;
wire v_72533;
wire v_72534;
wire v_72535;
wire v_72536;
wire v_72537;
wire v_72538;
wire v_72539;
wire v_72540;
wire v_72541;
wire v_72542;
wire v_72543;
wire v_72544;
wire v_72545;
wire v_72546;
wire v_72547;
wire v_72548;
wire v_72549;
wire v_72550;
wire v_72551;
wire v_72552;
wire v_72553;
wire v_72554;
wire v_72555;
wire v_72556;
wire v_72557;
wire v_72558;
wire v_72559;
wire v_72560;
wire v_72561;
wire v_72562;
wire v_72563;
wire v_72564;
wire v_72565;
wire v_72566;
wire v_72567;
wire v_72568;
wire v_72569;
wire v_72570;
wire v_72571;
wire v_72572;
wire v_72573;
wire v_72574;
wire v_72575;
wire v_72576;
wire v_72577;
wire v_72578;
wire v_72579;
wire v_72580;
wire v_72581;
wire v_72582;
wire v_72583;
wire v_72584;
wire v_72585;
wire v_72586;
wire v_72587;
wire v_72588;
wire v_72589;
wire v_72590;
wire v_72591;
wire v_72592;
wire v_72593;
wire v_72594;
wire v_72595;
wire v_72596;
wire v_72597;
wire v_72598;
wire v_72599;
wire v_72600;
wire v_72601;
wire v_72602;
wire v_72603;
wire v_72604;
wire v_72605;
wire v_72606;
wire v_72607;
wire v_72608;
wire v_72609;
wire v_72610;
wire v_72611;
wire v_72612;
wire v_72613;
wire v_72614;
wire v_72615;
wire v_72616;
wire v_72617;
wire v_72618;
wire v_72619;
wire v_72620;
wire v_72621;
wire v_72622;
wire v_72623;
wire v_72624;
wire v_72625;
wire v_72626;
wire v_72627;
wire v_72628;
wire v_72629;
wire v_72630;
wire v_72631;
wire v_72632;
wire v_72633;
wire v_72634;
wire v_72635;
wire v_72636;
wire v_72637;
wire v_72638;
wire v_72639;
wire v_72640;
wire v_72641;
wire v_72642;
wire v_72643;
wire v_72644;
wire v_72645;
wire v_72646;
wire v_72647;
wire v_72648;
wire v_72649;
wire v_72650;
wire v_72651;
wire v_72652;
wire v_72653;
wire v_72654;
wire v_72655;
wire v_72656;
wire v_72657;
wire v_72658;
wire v_72659;
wire v_72660;
wire v_72661;
wire v_72662;
wire v_72663;
wire v_72664;
wire v_72665;
wire v_72666;
wire v_72667;
wire v_72668;
wire v_72669;
wire v_72670;
wire v_72671;
wire v_72672;
wire v_72673;
wire v_72674;
wire v_72675;
wire v_72676;
wire v_72677;
wire v_72678;
wire v_72679;
wire v_72680;
wire v_72681;
wire v_72682;
wire v_72683;
wire v_72684;
wire v_72685;
wire v_72686;
wire v_72687;
wire v_72688;
wire v_72689;
wire v_72690;
wire v_72691;
wire v_72692;
wire v_72693;
wire v_72694;
wire v_72695;
wire v_72696;
wire v_72697;
wire v_72698;
wire v_72699;
wire v_72700;
wire v_72701;
wire v_72702;
wire v_72703;
wire v_72704;
wire v_72705;
wire v_72706;
wire v_72707;
wire v_72708;
wire v_72709;
wire v_72710;
wire v_72711;
wire v_72712;
wire v_72713;
wire v_72714;
wire v_72715;
wire v_72716;
wire v_72717;
wire v_72718;
wire v_72719;
wire v_72720;
wire v_72721;
wire v_72722;
wire v_72723;
wire v_72724;
wire v_72725;
wire v_72726;
wire v_72727;
wire v_72728;
wire v_72729;
wire v_72730;
wire v_72731;
wire v_72732;
wire v_72733;
wire v_72734;
wire v_72735;
wire v_72736;
wire v_72737;
wire v_72738;
wire v_72739;
wire v_72740;
wire v_72741;
wire v_72742;
wire v_72743;
wire v_72744;
wire v_72745;
wire v_72746;
wire v_72747;
wire v_72748;
wire v_72749;
wire v_72750;
wire v_72751;
wire v_72752;
wire v_72753;
wire v_72754;
wire v_72755;
wire v_72756;
wire v_72757;
wire v_72758;
wire v_72759;
wire v_72760;
wire v_72761;
wire v_72762;
wire v_72763;
wire v_72764;
wire v_72765;
wire v_72766;
wire v_72767;
wire v_72768;
wire v_72769;
wire v_72770;
wire v_72771;
wire v_72772;
wire v_72773;
wire v_72774;
wire v_72775;
wire v_72776;
wire v_72777;
wire v_72778;
wire v_72779;
wire v_72780;
wire v_72781;
wire v_72782;
wire v_72783;
wire v_72784;
wire v_72785;
wire v_72786;
wire v_72787;
wire v_72788;
wire v_72789;
wire v_72790;
wire v_72791;
wire v_72792;
wire v_72793;
wire v_72794;
wire v_72795;
wire v_72796;
wire v_72797;
wire v_72798;
wire v_72799;
wire v_72800;
wire v_72801;
wire v_72802;
wire v_72803;
wire v_72804;
wire v_72805;
wire v_72806;
wire v_72807;
wire v_72808;
wire v_72809;
wire v_72810;
wire v_72811;
wire v_72812;
wire v_72813;
wire v_72814;
wire v_72815;
wire v_72816;
wire v_72817;
wire v_72818;
wire v_72819;
wire v_72820;
wire v_72821;
wire v_72822;
wire v_72823;
wire v_72824;
wire v_72825;
wire v_72826;
wire v_72827;
wire v_72828;
wire v_72829;
wire v_72830;
wire v_72831;
wire v_72832;
wire v_72833;
wire v_72834;
wire v_72835;
wire v_72836;
wire v_72837;
wire v_72838;
wire v_72839;
wire v_72840;
wire v_72841;
wire v_72842;
wire v_72843;
wire v_72844;
wire v_72845;
wire v_72846;
wire v_72847;
wire v_72848;
wire v_72849;
wire v_72850;
wire v_72851;
wire v_72852;
wire v_72853;
wire v_72854;
wire v_72855;
wire v_72856;
wire v_72857;
wire v_72858;
wire v_72859;
wire v_72860;
wire v_72861;
wire v_72862;
wire v_72863;
wire v_72864;
wire v_72865;
wire v_72866;
wire v_72867;
wire v_72868;
wire v_72869;
wire v_72870;
wire v_72871;
wire v_72872;
wire v_72873;
wire v_72874;
wire v_72875;
wire v_72876;
wire v_72877;
wire v_72878;
wire v_72879;
wire v_72880;
wire v_72881;
wire v_72882;
wire v_72883;
wire v_72884;
wire v_72885;
wire v_72886;
wire v_72887;
wire v_72888;
wire v_72889;
wire v_72890;
wire v_72891;
wire v_72892;
wire v_72893;
wire v_72894;
wire v_72895;
wire v_72896;
wire v_72897;
wire v_72898;
wire v_72899;
wire v_72900;
wire v_72901;
wire v_72902;
wire v_72903;
wire v_72904;
wire v_72905;
wire v_72906;
wire v_72907;
wire v_72908;
wire v_72909;
wire v_72910;
wire v_72911;
wire v_72912;
wire v_72913;
wire v_72914;
wire v_72915;
wire v_72916;
wire v_72917;
wire v_72918;
wire v_72919;
wire v_72920;
wire v_72921;
wire v_72922;
wire v_72923;
wire v_72924;
wire v_72925;
wire v_72926;
wire v_72927;
wire v_72928;
wire v_72929;
wire v_72930;
wire v_72931;
wire v_72932;
wire v_72933;
wire v_72934;
wire v_72935;
wire v_72936;
wire v_72937;
wire v_72938;
wire v_72939;
wire v_72940;
wire v_72941;
wire v_72942;
wire v_72943;
wire v_72944;
wire v_72945;
wire v_72946;
wire v_72947;
wire v_72948;
wire v_72949;
wire v_72950;
wire v_72951;
wire v_72952;
wire v_72953;
wire v_72954;
wire v_72955;
wire v_72956;
wire v_72957;
wire v_72958;
wire v_72959;
wire v_72960;
wire v_72961;
wire v_72962;
wire v_72963;
wire v_72964;
wire v_72965;
wire v_72966;
wire v_72967;
wire v_72968;
wire v_72969;
wire v_72970;
wire v_72971;
wire v_72972;
wire v_72973;
wire v_72974;
wire v_72975;
wire v_72976;
wire v_72977;
wire v_72978;
wire v_72979;
wire v_72980;
wire v_72981;
wire v_72982;
wire v_72983;
wire v_72984;
wire v_72985;
wire v_72986;
wire v_72987;
wire v_72988;
wire v_72989;
wire v_72990;
wire v_72991;
wire v_72992;
wire v_72993;
wire v_72994;
wire v_72995;
wire v_72996;
wire v_72997;
wire v_72998;
wire v_72999;
wire v_73000;
wire v_73001;
wire v_73002;
wire v_73003;
wire v_73004;
wire v_73005;
wire v_73006;
wire v_73007;
wire v_73008;
wire v_73009;
wire v_73010;
wire v_73011;
wire v_73012;
wire v_73013;
wire v_73014;
wire v_73015;
wire v_73016;
wire v_73017;
wire v_73018;
wire v_73019;
wire v_73020;
wire v_73021;
wire v_73022;
wire v_73023;
wire v_73024;
wire v_73025;
wire v_73026;
wire v_73027;
wire v_73028;
wire v_73029;
wire v_73030;
wire v_73031;
wire v_73032;
wire v_73033;
wire v_73034;
wire v_73035;
wire v_73036;
wire v_73037;
wire v_73038;
wire v_73039;
wire v_73040;
wire v_73041;
wire v_73042;
wire v_73043;
wire v_73044;
wire v_73045;
wire v_73046;
wire v_73047;
wire v_73048;
wire v_73049;
wire v_73050;
wire v_73051;
wire v_73052;
wire v_73053;
wire v_73054;
wire v_73055;
wire v_73056;
wire v_73057;
wire v_73058;
wire v_73059;
wire v_73060;
wire v_73061;
wire v_73062;
wire v_73063;
wire v_73064;
wire v_73065;
wire v_73066;
wire v_73067;
wire v_73068;
wire v_73069;
wire v_73070;
wire v_73071;
wire v_73072;
wire v_73073;
wire v_73074;
wire v_73075;
wire v_73076;
wire v_73077;
wire v_73078;
wire v_73079;
wire v_73080;
wire v_73081;
wire v_73082;
wire v_73083;
wire v_73084;
wire v_73085;
wire v_73086;
wire v_73087;
wire v_73088;
wire v_73089;
wire v_73090;
wire v_73091;
wire v_73092;
wire v_73093;
wire v_73094;
wire v_73095;
wire v_73096;
wire v_73097;
wire v_73098;
wire v_73099;
wire v_73100;
wire v_73101;
wire v_73102;
wire v_73103;
wire v_73104;
wire v_73105;
wire v_73106;
wire v_73107;
wire v_73108;
wire v_73109;
wire v_73110;
wire v_73111;
wire v_73112;
wire v_73113;
wire v_73114;
wire v_73115;
wire v_73116;
wire v_73117;
wire v_73118;
wire v_73119;
wire v_73120;
wire v_73121;
wire v_73122;
wire v_73123;
wire x_1;
assign v_11 = 0;
assign v_7 = 1;
assign v_73123 = 1;
assign v_2 = v_1;
assign v_3 = v_2;
assign v_8 = ~v_6;
assign v_10 = ~v_9;
assign v_12 = v_9;
assign v_14 = ~v_13;
assign v_16 = ~v_15;
assign v_17 = v_15;
assign v_19 = ~v_18;
assign v_21 = ~v_20;
assign v_22 = v_20;
assign v_24 = ~v_23;
assign v_26 = ~v_25;
assign v_27 = v_25;
assign v_29 = ~v_28;
assign v_31 = ~v_30;
assign v_32 = v_30;
assign v_34 = ~v_33;
assign v_36 = ~v_35;
assign v_37 = v_35;
assign v_39 = ~v_38;
assign v_41 = ~v_40;
assign v_42 = v_40;
assign v_44 = ~v_43;
assign v_46 = ~v_45;
assign v_47 = v_45;
assign v_49 = ~v_48;
assign v_51 = ~v_50;
assign v_52 = v_50;
assign v_54 = ~v_53;
assign v_56 = ~v_55;
assign v_57 = v_55;
assign v_59 = ~v_58;
assign v_61 = ~v_60;
assign v_62 = v_60;
assign v_64 = ~v_63;
assign v_66 = ~v_65;
assign v_67 = v_65;
assign v_69 = ~v_68;
assign v_71 = ~v_70;
assign v_72 = v_70;
assign v_74 = ~v_73;
assign v_76 = ~v_75;
assign v_77 = v_75;
assign v_79 = ~v_78;
assign v_81 = ~v_80;
assign v_82 = v_80;
assign v_84 = ~v_83;
assign v_86 = ~v_85;
assign v_87 = v_85;
assign v_89 = ~v_88;
assign v_91 = ~v_90;
assign v_92 = v_91;
assign v_94 = v_93;
assign v_96 = v_86 & v_95;
assign v_98 = v_83;
assign v_100 = v_97 & v_99;
assign v_102 = v_81 & v_101;
assign v_104 = v_78;
assign v_106 = v_103 & v_105;
assign v_108 = v_76 & v_107;
assign v_110 = v_73;
assign v_112 = v_109 & v_111;
assign v_114 = v_71 & v_113;
assign v_116 = v_68;
assign v_118 = v_115 & v_117;
assign v_120 = v_66 & v_119;
assign v_122 = v_63;
assign v_124 = v_121 & v_123;
assign v_126 = v_61 & v_125;
assign v_128 = v_58;
assign v_130 = v_127 & v_129;
assign v_132 = v_56 & v_131;
assign v_134 = v_53;
assign v_136 = v_133 & v_135;
assign v_138 = v_51 & v_137;
assign v_140 = v_48;
assign v_142 = v_139 & v_141;
assign v_144 = v_46 & v_143;
assign v_146 = v_43;
assign v_148 = v_145 & v_147;
assign v_150 = v_41 & v_149;
assign v_152 = v_38;
assign v_154 = v_151 & v_153;
assign v_156 = v_36 & v_155;
assign v_158 = v_33;
assign v_160 = v_157 & v_159;
assign v_162 = v_31 & v_161;
assign v_164 = v_28;
assign v_166 = v_163 & v_165;
assign v_168 = v_26 & v_167;
assign v_170 = v_23;
assign v_172 = v_169 & v_171;
assign v_174 = v_21 & v_173;
assign v_176 = v_18;
assign v_178 = v_175 & v_177;
assign v_180 = v_16 & v_179;
assign v_182 = v_13;
assign v_184 = v_181 & v_183;
assign v_186 = v_10 & v_185;
assign v_188 = v_6;
assign v_190 = v_187 & v_189;
assign v_191 = v_190;
assign v_193 = v_88;
assign v_194 = v_90;
assign v_195 = v_194;
assign v_196 = v_193 & v_195;
assign v_197 = v_196;
assign v_198 = v_86 & v_197;
assign v_200 = v_98 & v_199;
assign v_201 = v_84 & v_197;
assign v_203 = v_81 & v_202;
assign v_205 = v_104 & v_204;
assign v_206 = v_79 & v_202;
assign v_208 = v_76 & v_207;
assign v_210 = v_110 & v_209;
assign v_211 = v_74 & v_207;
assign v_213 = v_71 & v_212;
assign v_215 = v_116 & v_214;
assign v_216 = v_69 & v_212;
assign v_218 = v_66 & v_217;
assign v_220 = v_122 & v_219;
assign v_221 = v_64 & v_217;
assign v_223 = v_61 & v_222;
assign v_225 = v_128 & v_224;
assign v_226 = v_59 & v_222;
assign v_228 = v_56 & v_227;
assign v_230 = v_134 & v_229;
assign v_231 = v_54 & v_227;
assign v_233 = v_51 & v_232;
assign v_235 = v_140 & v_234;
assign v_236 = v_49 & v_232;
assign v_238 = v_46 & v_237;
assign v_240 = v_146 & v_239;
assign v_241 = v_44 & v_237;
assign v_243 = v_41 & v_242;
assign v_245 = v_152 & v_244;
assign v_246 = v_39 & v_242;
assign v_248 = v_36 & v_247;
assign v_250 = v_158 & v_249;
assign v_251 = v_34 & v_247;
assign v_253 = v_31 & v_252;
assign v_255 = v_164 & v_254;
assign v_256 = v_29 & v_252;
assign v_258 = v_26 & v_257;
assign v_260 = v_170 & v_259;
assign v_261 = v_24 & v_257;
assign v_263 = v_21 & v_262;
assign v_265 = v_176 & v_264;
assign v_266 = v_19 & v_262;
assign v_268 = v_16 & v_267;
assign v_270 = v_182 & v_269;
assign v_271 = v_14 & v_267;
assign v_273 = v_10 & v_272;
assign v_275 = v_188 & v_274;
assign v_276 = v_8 & v_272;
assign v_278 = v_277;
assign v_280 = v_192 & v_279;
assign v_281 = v_280;
assign v_284 = ~v_283;
assign v_285 = ~v_9;
assign v_286 = v_9;
assign v_288 = ~v_287;
assign v_289 = ~v_15;
assign v_290 = v_15;
assign v_292 = ~v_291;
assign v_293 = ~v_20;
assign v_294 = v_20;
assign v_296 = ~v_295;
assign v_297 = ~v_25;
assign v_298 = v_25;
assign v_299 = ~v_28;
assign v_301 = ~v_300;
assign v_302 = v_300;
assign v_303 = ~v_33;
assign v_305 = ~v_304;
assign v_306 = v_304;
assign v_307 = ~v_38;
assign v_309 = ~v_308;
assign v_310 = v_308;
assign v_311 = ~v_43;
assign v_313 = ~v_312;
assign v_314 = v_312;
assign v_315 = ~v_48;
assign v_317 = ~v_316;
assign v_318 = v_316;
assign v_319 = ~v_53;
assign v_321 = ~v_320;
assign v_322 = v_320;
assign v_323 = ~v_58;
assign v_325 = ~v_324;
assign v_326 = v_324;
assign v_327 = ~v_63;
assign v_329 = ~v_328;
assign v_330 = v_328;
assign v_331 = ~v_68;
assign v_333 = ~v_332;
assign v_334 = v_332;
assign v_335 = ~v_73;
assign v_337 = ~v_336;
assign v_338 = v_336;
assign v_339 = ~v_78;
assign v_341 = ~v_340;
assign v_342 = v_340;
assign v_343 = ~v_83;
assign v_345 = ~v_344;
assign v_346 = v_344;
assign v_347 = ~v_88;
assign v_349 = ~v_348;
assign v_350 = v_349;
assign v_352 = v_351;
assign v_354 = v_345 & v_353;
assign v_356 = v_83;
assign v_358 = v_355 & v_357;
assign v_360 = v_341 & v_359;
assign v_362 = v_78;
assign v_364 = v_361 & v_363;
assign v_366 = v_337 & v_365;
assign v_368 = v_73;
assign v_370 = v_367 & v_369;
assign v_372 = v_333 & v_371;
assign v_374 = v_68;
assign v_376 = v_373 & v_375;
assign v_378 = v_329 & v_377;
assign v_380 = v_63;
assign v_382 = v_379 & v_381;
assign v_384 = v_325 & v_383;
assign v_386 = v_58;
assign v_388 = v_385 & v_387;
assign v_390 = v_321 & v_389;
assign v_392 = v_53;
assign v_394 = v_391 & v_393;
assign v_396 = v_317 & v_395;
assign v_398 = v_48;
assign v_400 = v_397 & v_399;
assign v_402 = v_313 & v_401;
assign v_404 = v_43;
assign v_406 = v_403 & v_405;
assign v_408 = v_309 & v_407;
assign v_410 = v_38;
assign v_412 = v_409 & v_411;
assign v_414 = v_305 & v_413;
assign v_416 = v_33;
assign v_418 = v_415 & v_417;
assign v_420 = v_301 & v_419;
assign v_422 = v_28;
assign v_424 = v_421 & v_423;
assign v_426 = v_297 & v_425;
assign v_428 = v_295;
assign v_430 = v_427 & v_429;
assign v_432 = v_293 & v_431;
assign v_434 = v_291;
assign v_436 = v_433 & v_435;
assign v_438 = v_289 & v_437;
assign v_440 = v_287;
assign v_442 = v_439 & v_441;
assign v_444 = v_285 & v_443;
assign v_446 = v_283;
assign v_448 = v_445 & v_447;
assign v_449 = v_448;
assign v_451 = v_88;
assign v_452 = v_348;
assign v_453 = v_452;
assign v_454 = v_451 & v_453;
assign v_455 = v_454;
assign v_456 = v_345 & v_455;
assign v_458 = v_356 & v_457;
assign v_459 = v_343 & v_455;
assign v_461 = v_341 & v_460;
assign v_463 = v_362 & v_462;
assign v_464 = v_339 & v_460;
assign v_466 = v_337 & v_465;
assign v_468 = v_368 & v_467;
assign v_469 = v_335 & v_465;
assign v_471 = v_333 & v_470;
assign v_473 = v_374 & v_472;
assign v_474 = v_331 & v_470;
assign v_476 = v_329 & v_475;
assign v_478 = v_380 & v_477;
assign v_479 = v_327 & v_475;
assign v_481 = v_325 & v_480;
assign v_483 = v_386 & v_482;
assign v_484 = v_323 & v_480;
assign v_486 = v_321 & v_485;
assign v_488 = v_392 & v_487;
assign v_489 = v_319 & v_485;
assign v_491 = v_317 & v_490;
assign v_493 = v_398 & v_492;
assign v_494 = v_315 & v_490;
assign v_496 = v_313 & v_495;
assign v_498 = v_404 & v_497;
assign v_499 = v_311 & v_495;
assign v_501 = v_309 & v_500;
assign v_503 = v_410 & v_502;
assign v_504 = v_307 & v_500;
assign v_506 = v_305 & v_505;
assign v_508 = v_416 & v_507;
assign v_509 = v_303 & v_505;
assign v_511 = v_301 & v_510;
assign v_513 = v_422 & v_512;
assign v_514 = v_299 & v_510;
assign v_516 = v_297 & v_515;
assign v_518 = v_428 & v_517;
assign v_519 = v_296 & v_515;
assign v_521 = v_293 & v_520;
assign v_523 = v_434 & v_522;
assign v_524 = v_292 & v_520;
assign v_526 = v_289 & v_525;
assign v_528 = v_440 & v_527;
assign v_529 = v_288 & v_525;
assign v_531 = v_285 & v_530;
assign v_533 = v_446 & v_532;
assign v_534 = v_284 & v_530;
assign v_536 = v_535;
assign v_538 = v_450 & v_537;
assign v_539 = v_538;
assign v_541 = v_540;
assign v_544 = ~v_543;
assign v_545 = ~v_9;
assign v_546 = v_9;
assign v_548 = ~v_547;
assign v_549 = ~v_15;
assign v_550 = v_15;
assign v_552 = ~v_551;
assign v_553 = ~v_20;
assign v_554 = v_20;
assign v_556 = ~v_555;
assign v_557 = ~v_25;
assign v_558 = v_25;
assign v_559 = ~v_28;
assign v_561 = ~v_560;
assign v_562 = v_560;
assign v_563 = ~v_33;
assign v_565 = ~v_564;
assign v_566 = v_564;
assign v_567 = ~v_38;
assign v_569 = ~v_568;
assign v_570 = v_568;
assign v_571 = ~v_43;
assign v_573 = ~v_572;
assign v_574 = v_572;
assign v_575 = ~v_48;
assign v_577 = ~v_576;
assign v_578 = v_576;
assign v_579 = ~v_53;
assign v_581 = ~v_580;
assign v_582 = v_580;
assign v_583 = ~v_58;
assign v_585 = ~v_584;
assign v_586 = v_584;
assign v_587 = ~v_63;
assign v_589 = ~v_588;
assign v_590 = v_588;
assign v_591 = ~v_68;
assign v_593 = ~v_592;
assign v_594 = v_592;
assign v_595 = ~v_73;
assign v_597 = ~v_596;
assign v_598 = v_596;
assign v_599 = ~v_78;
assign v_601 = ~v_600;
assign v_602 = v_600;
assign v_603 = ~v_83;
assign v_605 = ~v_604;
assign v_606 = v_604;
assign v_607 = ~v_88;
assign v_609 = ~v_608;
assign v_610 = v_609;
assign v_612 = v_611;
assign v_614 = v_605 & v_613;
assign v_616 = v_83;
assign v_618 = v_615 & v_617;
assign v_620 = v_601 & v_619;
assign v_622 = v_78;
assign v_624 = v_621 & v_623;
assign v_626 = v_597 & v_625;
assign v_628 = v_73;
assign v_630 = v_627 & v_629;
assign v_632 = v_593 & v_631;
assign v_634 = v_68;
assign v_636 = v_633 & v_635;
assign v_638 = v_589 & v_637;
assign v_640 = v_63;
assign v_642 = v_639 & v_641;
assign v_644 = v_585 & v_643;
assign v_646 = v_58;
assign v_648 = v_645 & v_647;
assign v_650 = v_581 & v_649;
assign v_652 = v_53;
assign v_654 = v_651 & v_653;
assign v_656 = v_577 & v_655;
assign v_658 = v_48;
assign v_660 = v_657 & v_659;
assign v_662 = v_573 & v_661;
assign v_664 = v_43;
assign v_666 = v_663 & v_665;
assign v_668 = v_569 & v_667;
assign v_670 = v_38;
assign v_672 = v_669 & v_671;
assign v_674 = v_565 & v_673;
assign v_676 = v_33;
assign v_678 = v_675 & v_677;
assign v_680 = v_561 & v_679;
assign v_682 = v_28;
assign v_684 = v_681 & v_683;
assign v_686 = v_557 & v_685;
assign v_688 = v_555;
assign v_690 = v_687 & v_689;
assign v_692 = v_553 & v_691;
assign v_694 = v_551;
assign v_696 = v_693 & v_695;
assign v_698 = v_549 & v_697;
assign v_700 = v_547;
assign v_702 = v_699 & v_701;
assign v_704 = v_545 & v_703;
assign v_706 = v_543;
assign v_708 = v_705 & v_707;
assign v_709 = v_708;
assign v_711 = v_88;
assign v_712 = v_608;
assign v_713 = v_712;
assign v_714 = v_711 & v_713;
assign v_715 = v_714;
assign v_716 = v_605 & v_715;
assign v_718 = v_616 & v_717;
assign v_719 = v_603 & v_715;
assign v_721 = v_601 & v_720;
assign v_723 = v_622 & v_722;
assign v_724 = v_599 & v_720;
assign v_726 = v_597 & v_725;
assign v_728 = v_628 & v_727;
assign v_729 = v_595 & v_725;
assign v_731 = v_593 & v_730;
assign v_733 = v_634 & v_732;
assign v_734 = v_591 & v_730;
assign v_736 = v_589 & v_735;
assign v_738 = v_640 & v_737;
assign v_739 = v_587 & v_735;
assign v_741 = v_585 & v_740;
assign v_743 = v_646 & v_742;
assign v_744 = v_583 & v_740;
assign v_746 = v_581 & v_745;
assign v_748 = v_652 & v_747;
assign v_749 = v_579 & v_745;
assign v_751 = v_577 & v_750;
assign v_753 = v_658 & v_752;
assign v_754 = v_575 & v_750;
assign v_756 = v_573 & v_755;
assign v_758 = v_664 & v_757;
assign v_759 = v_571 & v_755;
assign v_761 = v_569 & v_760;
assign v_763 = v_670 & v_762;
assign v_764 = v_567 & v_760;
assign v_766 = v_565 & v_765;
assign v_768 = v_676 & v_767;
assign v_769 = v_563 & v_765;
assign v_771 = v_561 & v_770;
assign v_773 = v_682 & v_772;
assign v_774 = v_559 & v_770;
assign v_776 = v_557 & v_775;
assign v_778 = v_688 & v_777;
assign v_779 = v_556 & v_775;
assign v_781 = v_553 & v_780;
assign v_783 = v_694 & v_782;
assign v_784 = v_552 & v_780;
assign v_786 = v_549 & v_785;
assign v_788 = v_700 & v_787;
assign v_789 = v_548 & v_785;
assign v_791 = v_545 & v_790;
assign v_793 = v_706 & v_792;
assign v_794 = v_544 & v_790;
assign v_796 = v_795;
assign v_798 = v_710 & v_797;
assign v_799 = v_798;
assign v_801 = v_800;
assign v_804 = ~v_803;
assign v_805 = ~v_9;
assign v_806 = v_9;
assign v_808 = ~v_807;
assign v_809 = ~v_15;
assign v_810 = v_15;
assign v_812 = ~v_811;
assign v_813 = ~v_20;
assign v_814 = v_20;
assign v_816 = ~v_815;
assign v_817 = ~v_25;
assign v_818 = v_25;
assign v_819 = ~v_28;
assign v_821 = ~v_820;
assign v_822 = v_820;
assign v_823 = ~v_33;
assign v_825 = ~v_824;
assign v_826 = v_824;
assign v_827 = ~v_38;
assign v_829 = ~v_828;
assign v_830 = v_828;
assign v_831 = ~v_43;
assign v_833 = ~v_832;
assign v_834 = v_832;
assign v_835 = ~v_48;
assign v_837 = ~v_836;
assign v_838 = v_836;
assign v_839 = ~v_53;
assign v_841 = ~v_840;
assign v_842 = v_840;
assign v_843 = ~v_58;
assign v_845 = ~v_844;
assign v_846 = v_844;
assign v_847 = ~v_63;
assign v_849 = ~v_848;
assign v_850 = v_848;
assign v_851 = ~v_68;
assign v_853 = ~v_852;
assign v_854 = v_852;
assign v_855 = ~v_73;
assign v_857 = ~v_856;
assign v_858 = v_856;
assign v_859 = ~v_78;
assign v_861 = ~v_860;
assign v_862 = v_860;
assign v_863 = ~v_83;
assign v_865 = ~v_864;
assign v_866 = v_864;
assign v_867 = ~v_88;
assign v_869 = ~v_868;
assign v_870 = v_869;
assign v_872 = v_871;
assign v_874 = v_865 & v_873;
assign v_876 = v_83;
assign v_878 = v_875 & v_877;
assign v_880 = v_861 & v_879;
assign v_882 = v_78;
assign v_884 = v_881 & v_883;
assign v_886 = v_857 & v_885;
assign v_888 = v_73;
assign v_890 = v_887 & v_889;
assign v_892 = v_853 & v_891;
assign v_894 = v_68;
assign v_896 = v_893 & v_895;
assign v_898 = v_849 & v_897;
assign v_900 = v_63;
assign v_902 = v_899 & v_901;
assign v_904 = v_845 & v_903;
assign v_906 = v_58;
assign v_908 = v_905 & v_907;
assign v_910 = v_841 & v_909;
assign v_912 = v_53;
assign v_914 = v_911 & v_913;
assign v_916 = v_837 & v_915;
assign v_918 = v_48;
assign v_920 = v_917 & v_919;
assign v_922 = v_833 & v_921;
assign v_924 = v_43;
assign v_926 = v_923 & v_925;
assign v_928 = v_829 & v_927;
assign v_930 = v_38;
assign v_932 = v_929 & v_931;
assign v_934 = v_825 & v_933;
assign v_936 = v_33;
assign v_938 = v_935 & v_937;
assign v_940 = v_821 & v_939;
assign v_942 = v_28;
assign v_944 = v_941 & v_943;
assign v_946 = v_817 & v_945;
assign v_948 = v_815;
assign v_950 = v_947 & v_949;
assign v_952 = v_813 & v_951;
assign v_954 = v_811;
assign v_956 = v_953 & v_955;
assign v_958 = v_809 & v_957;
assign v_960 = v_807;
assign v_962 = v_959 & v_961;
assign v_964 = v_805 & v_963;
assign v_966 = v_803;
assign v_968 = v_965 & v_967;
assign v_969 = v_968;
assign v_971 = v_88;
assign v_972 = v_868;
assign v_973 = v_972;
assign v_974 = v_971 & v_973;
assign v_975 = v_974;
assign v_976 = v_865 & v_975;
assign v_978 = v_876 & v_977;
assign v_979 = v_863 & v_975;
assign v_981 = v_861 & v_980;
assign v_983 = v_882 & v_982;
assign v_984 = v_859 & v_980;
assign v_986 = v_857 & v_985;
assign v_988 = v_888 & v_987;
assign v_989 = v_855 & v_985;
assign v_991 = v_853 & v_990;
assign v_993 = v_894 & v_992;
assign v_994 = v_851 & v_990;
assign v_996 = v_849 & v_995;
assign v_998 = v_900 & v_997;
assign v_999 = v_847 & v_995;
assign v_1001 = v_845 & v_1000;
assign v_1003 = v_906 & v_1002;
assign v_1004 = v_843 & v_1000;
assign v_1006 = v_841 & v_1005;
assign v_1008 = v_912 & v_1007;
assign v_1009 = v_839 & v_1005;
assign v_1011 = v_837 & v_1010;
assign v_1013 = v_918 & v_1012;
assign v_1014 = v_835 & v_1010;
assign v_1016 = v_833 & v_1015;
assign v_1018 = v_924 & v_1017;
assign v_1019 = v_831 & v_1015;
assign v_1021 = v_829 & v_1020;
assign v_1023 = v_930 & v_1022;
assign v_1024 = v_827 & v_1020;
assign v_1026 = v_825 & v_1025;
assign v_1028 = v_936 & v_1027;
assign v_1029 = v_823 & v_1025;
assign v_1031 = v_821 & v_1030;
assign v_1033 = v_942 & v_1032;
assign v_1034 = v_819 & v_1030;
assign v_1036 = v_817 & v_1035;
assign v_1038 = v_948 & v_1037;
assign v_1039 = v_816 & v_1035;
assign v_1041 = v_813 & v_1040;
assign v_1043 = v_954 & v_1042;
assign v_1044 = v_812 & v_1040;
assign v_1046 = v_809 & v_1045;
assign v_1048 = v_960 & v_1047;
assign v_1049 = v_808 & v_1045;
assign v_1051 = v_805 & v_1050;
assign v_1053 = v_966 & v_1052;
assign v_1054 = v_804 & v_1050;
assign v_1056 = v_1055;
assign v_1058 = v_970 & v_1057;
assign v_1059 = v_1058;
assign v_1061 = v_1060;
assign v_1064 = ~v_1063;
assign v_1065 = ~v_9;
assign v_1066 = v_9;
assign v_1068 = ~v_1067;
assign v_1069 = ~v_15;
assign v_1070 = v_15;
assign v_1072 = ~v_1071;
assign v_1073 = ~v_20;
assign v_1074 = v_20;
assign v_1076 = ~v_1075;
assign v_1077 = ~v_25;
assign v_1078 = v_25;
assign v_1079 = ~v_28;
assign v_1081 = ~v_1080;
assign v_1082 = v_1080;
assign v_1083 = ~v_33;
assign v_1085 = ~v_1084;
assign v_1086 = v_1084;
assign v_1087 = ~v_38;
assign v_1089 = ~v_1088;
assign v_1090 = v_1088;
assign v_1091 = ~v_43;
assign v_1093 = ~v_1092;
assign v_1094 = v_1092;
assign v_1095 = ~v_48;
assign v_1097 = ~v_1096;
assign v_1098 = v_1096;
assign v_1099 = ~v_53;
assign v_1101 = ~v_1100;
assign v_1102 = v_1100;
assign v_1103 = ~v_58;
assign v_1105 = ~v_1104;
assign v_1106 = v_1104;
assign v_1107 = ~v_63;
assign v_1109 = ~v_1108;
assign v_1110 = v_1108;
assign v_1111 = ~v_68;
assign v_1113 = ~v_1112;
assign v_1114 = v_1112;
assign v_1115 = ~v_73;
assign v_1117 = ~v_1116;
assign v_1118 = v_1116;
assign v_1119 = ~v_78;
assign v_1121 = ~v_1120;
assign v_1122 = v_1120;
assign v_1123 = ~v_83;
assign v_1125 = ~v_1124;
assign v_1126 = v_1124;
assign v_1127 = ~v_88;
assign v_1129 = ~v_1128;
assign v_1130 = v_1129;
assign v_1132 = v_1131;
assign v_1134 = v_1125 & v_1133;
assign v_1136 = v_83;
assign v_1138 = v_1135 & v_1137;
assign v_1140 = v_1121 & v_1139;
assign v_1142 = v_78;
assign v_1144 = v_1141 & v_1143;
assign v_1146 = v_1117 & v_1145;
assign v_1148 = v_73;
assign v_1150 = v_1147 & v_1149;
assign v_1152 = v_1113 & v_1151;
assign v_1154 = v_68;
assign v_1156 = v_1153 & v_1155;
assign v_1158 = v_1109 & v_1157;
assign v_1160 = v_63;
assign v_1162 = v_1159 & v_1161;
assign v_1164 = v_1105 & v_1163;
assign v_1166 = v_58;
assign v_1168 = v_1165 & v_1167;
assign v_1170 = v_1101 & v_1169;
assign v_1172 = v_53;
assign v_1174 = v_1171 & v_1173;
assign v_1176 = v_1097 & v_1175;
assign v_1178 = v_48;
assign v_1180 = v_1177 & v_1179;
assign v_1182 = v_1093 & v_1181;
assign v_1184 = v_43;
assign v_1186 = v_1183 & v_1185;
assign v_1188 = v_1089 & v_1187;
assign v_1190 = v_38;
assign v_1192 = v_1189 & v_1191;
assign v_1194 = v_1085 & v_1193;
assign v_1196 = v_33;
assign v_1198 = v_1195 & v_1197;
assign v_1200 = v_1081 & v_1199;
assign v_1202 = v_28;
assign v_1204 = v_1201 & v_1203;
assign v_1206 = v_1077 & v_1205;
assign v_1208 = v_1075;
assign v_1210 = v_1207 & v_1209;
assign v_1212 = v_1073 & v_1211;
assign v_1214 = v_1071;
assign v_1216 = v_1213 & v_1215;
assign v_1218 = v_1069 & v_1217;
assign v_1220 = v_1067;
assign v_1222 = v_1219 & v_1221;
assign v_1224 = v_1065 & v_1223;
assign v_1226 = v_1063;
assign v_1228 = v_1225 & v_1227;
assign v_1229 = v_1228;
assign v_1231 = v_88;
assign v_1232 = v_1128;
assign v_1233 = v_1232;
assign v_1234 = v_1231 & v_1233;
assign v_1235 = v_1234;
assign v_1236 = v_1125 & v_1235;
assign v_1238 = v_1136 & v_1237;
assign v_1239 = v_1123 & v_1235;
assign v_1241 = v_1121 & v_1240;
assign v_1243 = v_1142 & v_1242;
assign v_1244 = v_1119 & v_1240;
assign v_1246 = v_1117 & v_1245;
assign v_1248 = v_1148 & v_1247;
assign v_1249 = v_1115 & v_1245;
assign v_1251 = v_1113 & v_1250;
assign v_1253 = v_1154 & v_1252;
assign v_1254 = v_1111 & v_1250;
assign v_1256 = v_1109 & v_1255;
assign v_1258 = v_1160 & v_1257;
assign v_1259 = v_1107 & v_1255;
assign v_1261 = v_1105 & v_1260;
assign v_1263 = v_1166 & v_1262;
assign v_1264 = v_1103 & v_1260;
assign v_1266 = v_1101 & v_1265;
assign v_1268 = v_1172 & v_1267;
assign v_1269 = v_1099 & v_1265;
assign v_1271 = v_1097 & v_1270;
assign v_1273 = v_1178 & v_1272;
assign v_1274 = v_1095 & v_1270;
assign v_1276 = v_1093 & v_1275;
assign v_1278 = v_1184 & v_1277;
assign v_1279 = v_1091 & v_1275;
assign v_1281 = v_1089 & v_1280;
assign v_1283 = v_1190 & v_1282;
assign v_1284 = v_1087 & v_1280;
assign v_1286 = v_1085 & v_1285;
assign v_1288 = v_1196 & v_1287;
assign v_1289 = v_1083 & v_1285;
assign v_1291 = v_1081 & v_1290;
assign v_1293 = v_1202 & v_1292;
assign v_1294 = v_1079 & v_1290;
assign v_1296 = v_1077 & v_1295;
assign v_1298 = v_1208 & v_1297;
assign v_1299 = v_1076 & v_1295;
assign v_1301 = v_1073 & v_1300;
assign v_1303 = v_1214 & v_1302;
assign v_1304 = v_1072 & v_1300;
assign v_1306 = v_1069 & v_1305;
assign v_1308 = v_1220 & v_1307;
assign v_1309 = v_1068 & v_1305;
assign v_1311 = v_1065 & v_1310;
assign v_1313 = v_1226 & v_1312;
assign v_1314 = v_1064 & v_1310;
assign v_1316 = v_1315;
assign v_1318 = v_1230 & v_1317;
assign v_1319 = v_1318;
assign v_1321 = v_1320;
assign v_1324 = ~v_1323;
assign v_1325 = ~v_9;
assign v_1326 = v_9;
assign v_1328 = ~v_1327;
assign v_1329 = ~v_15;
assign v_1330 = v_15;
assign v_1332 = ~v_1331;
assign v_1333 = ~v_20;
assign v_1334 = v_20;
assign v_1336 = ~v_1335;
assign v_1337 = ~v_25;
assign v_1338 = v_25;
assign v_1339 = ~v_28;
assign v_1341 = ~v_1340;
assign v_1342 = v_1340;
assign v_1343 = ~v_33;
assign v_1345 = ~v_1344;
assign v_1346 = v_1344;
assign v_1347 = ~v_38;
assign v_1349 = ~v_1348;
assign v_1350 = v_1348;
assign v_1351 = ~v_43;
assign v_1353 = ~v_1352;
assign v_1354 = v_1352;
assign v_1355 = ~v_48;
assign v_1357 = ~v_1356;
assign v_1358 = v_1356;
assign v_1359 = ~v_53;
assign v_1361 = ~v_1360;
assign v_1362 = v_1360;
assign v_1363 = ~v_58;
assign v_1365 = ~v_1364;
assign v_1366 = v_1364;
assign v_1367 = ~v_63;
assign v_1369 = ~v_1368;
assign v_1370 = v_1368;
assign v_1371 = ~v_68;
assign v_1373 = ~v_1372;
assign v_1374 = v_1372;
assign v_1375 = ~v_73;
assign v_1377 = ~v_1376;
assign v_1378 = v_1376;
assign v_1379 = ~v_78;
assign v_1381 = ~v_1380;
assign v_1382 = v_1380;
assign v_1383 = ~v_83;
assign v_1385 = ~v_1384;
assign v_1386 = v_1384;
assign v_1387 = ~v_88;
assign v_1389 = ~v_1388;
assign v_1390 = v_1389;
assign v_1392 = v_1391;
assign v_1394 = v_1385 & v_1393;
assign v_1396 = v_83;
assign v_1398 = v_1395 & v_1397;
assign v_1400 = v_1381 & v_1399;
assign v_1402 = v_78;
assign v_1404 = v_1401 & v_1403;
assign v_1406 = v_1377 & v_1405;
assign v_1408 = v_73;
assign v_1410 = v_1407 & v_1409;
assign v_1412 = v_1373 & v_1411;
assign v_1414 = v_68;
assign v_1416 = v_1413 & v_1415;
assign v_1418 = v_1369 & v_1417;
assign v_1420 = v_63;
assign v_1422 = v_1419 & v_1421;
assign v_1424 = v_1365 & v_1423;
assign v_1426 = v_58;
assign v_1428 = v_1425 & v_1427;
assign v_1430 = v_1361 & v_1429;
assign v_1432 = v_53;
assign v_1434 = v_1431 & v_1433;
assign v_1436 = v_1357 & v_1435;
assign v_1438 = v_48;
assign v_1440 = v_1437 & v_1439;
assign v_1442 = v_1353 & v_1441;
assign v_1444 = v_43;
assign v_1446 = v_1443 & v_1445;
assign v_1448 = v_1349 & v_1447;
assign v_1450 = v_38;
assign v_1452 = v_1449 & v_1451;
assign v_1454 = v_1345 & v_1453;
assign v_1456 = v_33;
assign v_1458 = v_1455 & v_1457;
assign v_1460 = v_1341 & v_1459;
assign v_1462 = v_28;
assign v_1464 = v_1461 & v_1463;
assign v_1466 = v_1337 & v_1465;
assign v_1468 = v_1335;
assign v_1470 = v_1467 & v_1469;
assign v_1472 = v_1333 & v_1471;
assign v_1474 = v_1331;
assign v_1476 = v_1473 & v_1475;
assign v_1478 = v_1329 & v_1477;
assign v_1480 = v_1327;
assign v_1482 = v_1479 & v_1481;
assign v_1484 = v_1325 & v_1483;
assign v_1486 = v_1323;
assign v_1488 = v_1485 & v_1487;
assign v_1489 = v_1488;
assign v_1491 = v_88;
assign v_1492 = v_1388;
assign v_1493 = v_1492;
assign v_1494 = v_1491 & v_1493;
assign v_1495 = v_1494;
assign v_1496 = v_1385 & v_1495;
assign v_1498 = v_1396 & v_1497;
assign v_1499 = v_1383 & v_1495;
assign v_1501 = v_1381 & v_1500;
assign v_1503 = v_1402 & v_1502;
assign v_1504 = v_1379 & v_1500;
assign v_1506 = v_1377 & v_1505;
assign v_1508 = v_1408 & v_1507;
assign v_1509 = v_1375 & v_1505;
assign v_1511 = v_1373 & v_1510;
assign v_1513 = v_1414 & v_1512;
assign v_1514 = v_1371 & v_1510;
assign v_1516 = v_1369 & v_1515;
assign v_1518 = v_1420 & v_1517;
assign v_1519 = v_1367 & v_1515;
assign v_1521 = v_1365 & v_1520;
assign v_1523 = v_1426 & v_1522;
assign v_1524 = v_1363 & v_1520;
assign v_1526 = v_1361 & v_1525;
assign v_1528 = v_1432 & v_1527;
assign v_1529 = v_1359 & v_1525;
assign v_1531 = v_1357 & v_1530;
assign v_1533 = v_1438 & v_1532;
assign v_1534 = v_1355 & v_1530;
assign v_1536 = v_1353 & v_1535;
assign v_1538 = v_1444 & v_1537;
assign v_1539 = v_1351 & v_1535;
assign v_1541 = v_1349 & v_1540;
assign v_1543 = v_1450 & v_1542;
assign v_1544 = v_1347 & v_1540;
assign v_1546 = v_1345 & v_1545;
assign v_1548 = v_1456 & v_1547;
assign v_1549 = v_1343 & v_1545;
assign v_1551 = v_1341 & v_1550;
assign v_1553 = v_1462 & v_1552;
assign v_1554 = v_1339 & v_1550;
assign v_1556 = v_1337 & v_1555;
assign v_1558 = v_1468 & v_1557;
assign v_1559 = v_1336 & v_1555;
assign v_1561 = v_1333 & v_1560;
assign v_1563 = v_1474 & v_1562;
assign v_1564 = v_1332 & v_1560;
assign v_1566 = v_1329 & v_1565;
assign v_1568 = v_1480 & v_1567;
assign v_1569 = v_1328 & v_1565;
assign v_1571 = v_1325 & v_1570;
assign v_1573 = v_1486 & v_1572;
assign v_1574 = v_1324 & v_1570;
assign v_1576 = v_1575;
assign v_1578 = v_1490 & v_1577;
assign v_1579 = v_1578;
assign v_1581 = v_1580;
assign v_1584 = ~v_1583;
assign v_1585 = ~v_9;
assign v_1586 = v_9;
assign v_1588 = ~v_1587;
assign v_1589 = ~v_15;
assign v_1590 = v_15;
assign v_1592 = ~v_1591;
assign v_1593 = ~v_20;
assign v_1594 = v_20;
assign v_1596 = ~v_1595;
assign v_1597 = ~v_25;
assign v_1598 = v_25;
assign v_1599 = ~v_28;
assign v_1601 = ~v_1600;
assign v_1602 = v_1600;
assign v_1603 = ~v_33;
assign v_1605 = ~v_1604;
assign v_1606 = v_1604;
assign v_1607 = ~v_38;
assign v_1609 = ~v_1608;
assign v_1610 = v_1608;
assign v_1611 = ~v_43;
assign v_1613 = ~v_1612;
assign v_1614 = v_1612;
assign v_1615 = ~v_48;
assign v_1617 = ~v_1616;
assign v_1618 = v_1616;
assign v_1619 = ~v_53;
assign v_1621 = ~v_1620;
assign v_1622 = v_1620;
assign v_1623 = ~v_58;
assign v_1625 = ~v_1624;
assign v_1626 = v_1624;
assign v_1627 = ~v_63;
assign v_1629 = ~v_1628;
assign v_1630 = v_1628;
assign v_1631 = ~v_68;
assign v_1633 = ~v_1632;
assign v_1634 = v_1632;
assign v_1635 = ~v_73;
assign v_1637 = ~v_1636;
assign v_1638 = v_1636;
assign v_1639 = ~v_78;
assign v_1641 = ~v_1640;
assign v_1642 = v_1640;
assign v_1643 = ~v_83;
assign v_1645 = ~v_1644;
assign v_1646 = v_1644;
assign v_1647 = ~v_88;
assign v_1649 = ~v_1648;
assign v_1650 = v_1649;
assign v_1652 = v_1651;
assign v_1654 = v_1645 & v_1653;
assign v_1656 = v_83;
assign v_1658 = v_1655 & v_1657;
assign v_1660 = v_1641 & v_1659;
assign v_1662 = v_78;
assign v_1664 = v_1661 & v_1663;
assign v_1666 = v_1637 & v_1665;
assign v_1668 = v_73;
assign v_1670 = v_1667 & v_1669;
assign v_1672 = v_1633 & v_1671;
assign v_1674 = v_68;
assign v_1676 = v_1673 & v_1675;
assign v_1678 = v_1629 & v_1677;
assign v_1680 = v_63;
assign v_1682 = v_1679 & v_1681;
assign v_1684 = v_1625 & v_1683;
assign v_1686 = v_58;
assign v_1688 = v_1685 & v_1687;
assign v_1690 = v_1621 & v_1689;
assign v_1692 = v_53;
assign v_1694 = v_1691 & v_1693;
assign v_1696 = v_1617 & v_1695;
assign v_1698 = v_48;
assign v_1700 = v_1697 & v_1699;
assign v_1702 = v_1613 & v_1701;
assign v_1704 = v_43;
assign v_1706 = v_1703 & v_1705;
assign v_1708 = v_1609 & v_1707;
assign v_1710 = v_38;
assign v_1712 = v_1709 & v_1711;
assign v_1714 = v_1605 & v_1713;
assign v_1716 = v_33;
assign v_1718 = v_1715 & v_1717;
assign v_1720 = v_1601 & v_1719;
assign v_1722 = v_28;
assign v_1724 = v_1721 & v_1723;
assign v_1726 = v_1597 & v_1725;
assign v_1728 = v_1595;
assign v_1730 = v_1727 & v_1729;
assign v_1732 = v_1593 & v_1731;
assign v_1734 = v_1591;
assign v_1736 = v_1733 & v_1735;
assign v_1738 = v_1589 & v_1737;
assign v_1740 = v_1587;
assign v_1742 = v_1739 & v_1741;
assign v_1744 = v_1585 & v_1743;
assign v_1746 = v_1583;
assign v_1748 = v_1745 & v_1747;
assign v_1749 = v_1748;
assign v_1751 = v_88;
assign v_1752 = v_1648;
assign v_1753 = v_1752;
assign v_1754 = v_1751 & v_1753;
assign v_1755 = v_1754;
assign v_1756 = v_1645 & v_1755;
assign v_1758 = v_1656 & v_1757;
assign v_1759 = v_1643 & v_1755;
assign v_1761 = v_1641 & v_1760;
assign v_1763 = v_1662 & v_1762;
assign v_1764 = v_1639 & v_1760;
assign v_1766 = v_1637 & v_1765;
assign v_1768 = v_1668 & v_1767;
assign v_1769 = v_1635 & v_1765;
assign v_1771 = v_1633 & v_1770;
assign v_1773 = v_1674 & v_1772;
assign v_1774 = v_1631 & v_1770;
assign v_1776 = v_1629 & v_1775;
assign v_1778 = v_1680 & v_1777;
assign v_1779 = v_1627 & v_1775;
assign v_1781 = v_1625 & v_1780;
assign v_1783 = v_1686 & v_1782;
assign v_1784 = v_1623 & v_1780;
assign v_1786 = v_1621 & v_1785;
assign v_1788 = v_1692 & v_1787;
assign v_1789 = v_1619 & v_1785;
assign v_1791 = v_1617 & v_1790;
assign v_1793 = v_1698 & v_1792;
assign v_1794 = v_1615 & v_1790;
assign v_1796 = v_1613 & v_1795;
assign v_1798 = v_1704 & v_1797;
assign v_1799 = v_1611 & v_1795;
assign v_1801 = v_1609 & v_1800;
assign v_1803 = v_1710 & v_1802;
assign v_1804 = v_1607 & v_1800;
assign v_1806 = v_1605 & v_1805;
assign v_1808 = v_1716 & v_1807;
assign v_1809 = v_1603 & v_1805;
assign v_1811 = v_1601 & v_1810;
assign v_1813 = v_1722 & v_1812;
assign v_1814 = v_1599 & v_1810;
assign v_1816 = v_1597 & v_1815;
assign v_1818 = v_1728 & v_1817;
assign v_1819 = v_1596 & v_1815;
assign v_1821 = v_1593 & v_1820;
assign v_1823 = v_1734 & v_1822;
assign v_1824 = v_1592 & v_1820;
assign v_1826 = v_1589 & v_1825;
assign v_1828 = v_1740 & v_1827;
assign v_1829 = v_1588 & v_1825;
assign v_1831 = v_1585 & v_1830;
assign v_1833 = v_1746 & v_1832;
assign v_1834 = v_1584 & v_1830;
assign v_1836 = v_1835;
assign v_1838 = v_1750 & v_1837;
assign v_1839 = v_1838;
assign v_1841 = v_1840;
assign v_1844 = ~v_1843;
assign v_1845 = ~v_9;
assign v_1846 = v_9;
assign v_1848 = ~v_1847;
assign v_1849 = ~v_15;
assign v_1850 = v_15;
assign v_1852 = ~v_1851;
assign v_1853 = ~v_20;
assign v_1854 = v_20;
assign v_1856 = ~v_1855;
assign v_1857 = ~v_25;
assign v_1858 = v_25;
assign v_1859 = ~v_28;
assign v_1861 = ~v_1860;
assign v_1862 = v_1860;
assign v_1863 = ~v_33;
assign v_1865 = ~v_1864;
assign v_1866 = v_1864;
assign v_1867 = ~v_38;
assign v_1869 = ~v_1868;
assign v_1870 = v_1868;
assign v_1871 = ~v_43;
assign v_1873 = ~v_1872;
assign v_1874 = v_1872;
assign v_1875 = ~v_48;
assign v_1877 = ~v_1876;
assign v_1878 = v_1876;
assign v_1879 = ~v_53;
assign v_1881 = ~v_1880;
assign v_1882 = v_1880;
assign v_1883 = ~v_58;
assign v_1885 = ~v_1884;
assign v_1886 = v_1884;
assign v_1887 = ~v_63;
assign v_1889 = ~v_1888;
assign v_1890 = v_1888;
assign v_1891 = ~v_68;
assign v_1893 = ~v_1892;
assign v_1894 = v_1892;
assign v_1895 = ~v_73;
assign v_1897 = ~v_1896;
assign v_1898 = v_1896;
assign v_1899 = ~v_78;
assign v_1901 = ~v_1900;
assign v_1902 = v_1900;
assign v_1903 = ~v_83;
assign v_1905 = ~v_1904;
assign v_1906 = v_1904;
assign v_1907 = ~v_88;
assign v_1909 = ~v_1908;
assign v_1910 = v_1909;
assign v_1912 = v_1911;
assign v_1914 = v_1905 & v_1913;
assign v_1916 = v_83;
assign v_1918 = v_1915 & v_1917;
assign v_1920 = v_1901 & v_1919;
assign v_1922 = v_78;
assign v_1924 = v_1921 & v_1923;
assign v_1926 = v_1897 & v_1925;
assign v_1928 = v_73;
assign v_1930 = v_1927 & v_1929;
assign v_1932 = v_1893 & v_1931;
assign v_1934 = v_68;
assign v_1936 = v_1933 & v_1935;
assign v_1938 = v_1889 & v_1937;
assign v_1940 = v_63;
assign v_1942 = v_1939 & v_1941;
assign v_1944 = v_1885 & v_1943;
assign v_1946 = v_58;
assign v_1948 = v_1945 & v_1947;
assign v_1950 = v_1881 & v_1949;
assign v_1952 = v_53;
assign v_1954 = v_1951 & v_1953;
assign v_1956 = v_1877 & v_1955;
assign v_1958 = v_48;
assign v_1960 = v_1957 & v_1959;
assign v_1962 = v_1873 & v_1961;
assign v_1964 = v_43;
assign v_1966 = v_1963 & v_1965;
assign v_1968 = v_1869 & v_1967;
assign v_1970 = v_38;
assign v_1972 = v_1969 & v_1971;
assign v_1974 = v_1865 & v_1973;
assign v_1976 = v_33;
assign v_1978 = v_1975 & v_1977;
assign v_1980 = v_1861 & v_1979;
assign v_1982 = v_28;
assign v_1984 = v_1981 & v_1983;
assign v_1986 = v_1857 & v_1985;
assign v_1988 = v_1855;
assign v_1990 = v_1987 & v_1989;
assign v_1992 = v_1853 & v_1991;
assign v_1994 = v_1851;
assign v_1996 = v_1993 & v_1995;
assign v_1998 = v_1849 & v_1997;
assign v_2000 = v_1847;
assign v_2002 = v_1999 & v_2001;
assign v_2004 = v_1845 & v_2003;
assign v_2006 = v_1843;
assign v_2008 = v_2005 & v_2007;
assign v_2009 = v_2008;
assign v_2011 = v_88;
assign v_2012 = v_1908;
assign v_2013 = v_2012;
assign v_2014 = v_2011 & v_2013;
assign v_2015 = v_2014;
assign v_2016 = v_1905 & v_2015;
assign v_2018 = v_1916 & v_2017;
assign v_2019 = v_1903 & v_2015;
assign v_2021 = v_1901 & v_2020;
assign v_2023 = v_1922 & v_2022;
assign v_2024 = v_1899 & v_2020;
assign v_2026 = v_1897 & v_2025;
assign v_2028 = v_1928 & v_2027;
assign v_2029 = v_1895 & v_2025;
assign v_2031 = v_1893 & v_2030;
assign v_2033 = v_1934 & v_2032;
assign v_2034 = v_1891 & v_2030;
assign v_2036 = v_1889 & v_2035;
assign v_2038 = v_1940 & v_2037;
assign v_2039 = v_1887 & v_2035;
assign v_2041 = v_1885 & v_2040;
assign v_2043 = v_1946 & v_2042;
assign v_2044 = v_1883 & v_2040;
assign v_2046 = v_1881 & v_2045;
assign v_2048 = v_1952 & v_2047;
assign v_2049 = v_1879 & v_2045;
assign v_2051 = v_1877 & v_2050;
assign v_2053 = v_1958 & v_2052;
assign v_2054 = v_1875 & v_2050;
assign v_2056 = v_1873 & v_2055;
assign v_2058 = v_1964 & v_2057;
assign v_2059 = v_1871 & v_2055;
assign v_2061 = v_1869 & v_2060;
assign v_2063 = v_1970 & v_2062;
assign v_2064 = v_1867 & v_2060;
assign v_2066 = v_1865 & v_2065;
assign v_2068 = v_1976 & v_2067;
assign v_2069 = v_1863 & v_2065;
assign v_2071 = v_1861 & v_2070;
assign v_2073 = v_1982 & v_2072;
assign v_2074 = v_1859 & v_2070;
assign v_2076 = v_1857 & v_2075;
assign v_2078 = v_1988 & v_2077;
assign v_2079 = v_1856 & v_2075;
assign v_2081 = v_1853 & v_2080;
assign v_2083 = v_1994 & v_2082;
assign v_2084 = v_1852 & v_2080;
assign v_2086 = v_1849 & v_2085;
assign v_2088 = v_2000 & v_2087;
assign v_2089 = v_1848 & v_2085;
assign v_2091 = v_1845 & v_2090;
assign v_2093 = v_2006 & v_2092;
assign v_2094 = v_1844 & v_2090;
assign v_2096 = v_2095;
assign v_2098 = v_2010 & v_2097;
assign v_2099 = v_2098;
assign v_2101 = v_2100;
assign v_2104 = ~v_2103;
assign v_2105 = ~v_9;
assign v_2106 = v_9;
assign v_2108 = ~v_2107;
assign v_2109 = ~v_15;
assign v_2110 = v_15;
assign v_2112 = ~v_2111;
assign v_2113 = ~v_20;
assign v_2114 = v_20;
assign v_2116 = ~v_2115;
assign v_2117 = ~v_25;
assign v_2118 = v_25;
assign v_2119 = ~v_28;
assign v_2121 = ~v_2120;
assign v_2122 = v_2120;
assign v_2123 = ~v_33;
assign v_2125 = ~v_2124;
assign v_2126 = v_2124;
assign v_2127 = ~v_38;
assign v_2129 = ~v_2128;
assign v_2130 = v_2128;
assign v_2131 = ~v_43;
assign v_2133 = ~v_2132;
assign v_2134 = v_2132;
assign v_2135 = ~v_48;
assign v_2137 = ~v_2136;
assign v_2138 = v_2136;
assign v_2139 = ~v_53;
assign v_2141 = ~v_2140;
assign v_2142 = v_2140;
assign v_2143 = ~v_58;
assign v_2145 = ~v_2144;
assign v_2146 = v_2144;
assign v_2147 = ~v_63;
assign v_2149 = ~v_2148;
assign v_2150 = v_2148;
assign v_2151 = ~v_68;
assign v_2153 = ~v_2152;
assign v_2154 = v_2152;
assign v_2155 = ~v_73;
assign v_2157 = ~v_2156;
assign v_2158 = v_2156;
assign v_2159 = ~v_78;
assign v_2161 = ~v_2160;
assign v_2162 = v_2160;
assign v_2163 = ~v_83;
assign v_2165 = ~v_2164;
assign v_2166 = v_2164;
assign v_2167 = ~v_88;
assign v_2169 = ~v_2168;
assign v_2170 = v_2169;
assign v_2172 = v_2171;
assign v_2174 = v_2165 & v_2173;
assign v_2176 = v_83;
assign v_2178 = v_2175 & v_2177;
assign v_2180 = v_2161 & v_2179;
assign v_2182 = v_78;
assign v_2184 = v_2181 & v_2183;
assign v_2186 = v_2157 & v_2185;
assign v_2188 = v_73;
assign v_2190 = v_2187 & v_2189;
assign v_2192 = v_2153 & v_2191;
assign v_2194 = v_68;
assign v_2196 = v_2193 & v_2195;
assign v_2198 = v_2149 & v_2197;
assign v_2200 = v_63;
assign v_2202 = v_2199 & v_2201;
assign v_2204 = v_2145 & v_2203;
assign v_2206 = v_58;
assign v_2208 = v_2205 & v_2207;
assign v_2210 = v_2141 & v_2209;
assign v_2212 = v_53;
assign v_2214 = v_2211 & v_2213;
assign v_2216 = v_2137 & v_2215;
assign v_2218 = v_48;
assign v_2220 = v_2217 & v_2219;
assign v_2222 = v_2133 & v_2221;
assign v_2224 = v_43;
assign v_2226 = v_2223 & v_2225;
assign v_2228 = v_2129 & v_2227;
assign v_2230 = v_38;
assign v_2232 = v_2229 & v_2231;
assign v_2234 = v_2125 & v_2233;
assign v_2236 = v_33;
assign v_2238 = v_2235 & v_2237;
assign v_2240 = v_2121 & v_2239;
assign v_2242 = v_28;
assign v_2244 = v_2241 & v_2243;
assign v_2246 = v_2117 & v_2245;
assign v_2248 = v_2115;
assign v_2250 = v_2247 & v_2249;
assign v_2252 = v_2113 & v_2251;
assign v_2254 = v_2111;
assign v_2256 = v_2253 & v_2255;
assign v_2258 = v_2109 & v_2257;
assign v_2260 = v_2107;
assign v_2262 = v_2259 & v_2261;
assign v_2264 = v_2105 & v_2263;
assign v_2266 = v_2103;
assign v_2268 = v_2265 & v_2267;
assign v_2269 = v_2268;
assign v_2271 = v_88;
assign v_2272 = v_2168;
assign v_2273 = v_2272;
assign v_2274 = v_2271 & v_2273;
assign v_2275 = v_2274;
assign v_2276 = v_2165 & v_2275;
assign v_2278 = v_2176 & v_2277;
assign v_2279 = v_2163 & v_2275;
assign v_2281 = v_2161 & v_2280;
assign v_2283 = v_2182 & v_2282;
assign v_2284 = v_2159 & v_2280;
assign v_2286 = v_2157 & v_2285;
assign v_2288 = v_2188 & v_2287;
assign v_2289 = v_2155 & v_2285;
assign v_2291 = v_2153 & v_2290;
assign v_2293 = v_2194 & v_2292;
assign v_2294 = v_2151 & v_2290;
assign v_2296 = v_2149 & v_2295;
assign v_2298 = v_2200 & v_2297;
assign v_2299 = v_2147 & v_2295;
assign v_2301 = v_2145 & v_2300;
assign v_2303 = v_2206 & v_2302;
assign v_2304 = v_2143 & v_2300;
assign v_2306 = v_2141 & v_2305;
assign v_2308 = v_2212 & v_2307;
assign v_2309 = v_2139 & v_2305;
assign v_2311 = v_2137 & v_2310;
assign v_2313 = v_2218 & v_2312;
assign v_2314 = v_2135 & v_2310;
assign v_2316 = v_2133 & v_2315;
assign v_2318 = v_2224 & v_2317;
assign v_2319 = v_2131 & v_2315;
assign v_2321 = v_2129 & v_2320;
assign v_2323 = v_2230 & v_2322;
assign v_2324 = v_2127 & v_2320;
assign v_2326 = v_2125 & v_2325;
assign v_2328 = v_2236 & v_2327;
assign v_2329 = v_2123 & v_2325;
assign v_2331 = v_2121 & v_2330;
assign v_2333 = v_2242 & v_2332;
assign v_2334 = v_2119 & v_2330;
assign v_2336 = v_2117 & v_2335;
assign v_2338 = v_2248 & v_2337;
assign v_2339 = v_2116 & v_2335;
assign v_2341 = v_2113 & v_2340;
assign v_2343 = v_2254 & v_2342;
assign v_2344 = v_2112 & v_2340;
assign v_2346 = v_2109 & v_2345;
assign v_2348 = v_2260 & v_2347;
assign v_2349 = v_2108 & v_2345;
assign v_2351 = v_2105 & v_2350;
assign v_2353 = v_2266 & v_2352;
assign v_2354 = v_2104 & v_2350;
assign v_2356 = v_2355;
assign v_2358 = v_2270 & v_2357;
assign v_2359 = v_2358;
assign v_2361 = v_2360;
assign v_2364 = ~v_2363;
assign v_2365 = ~v_9;
assign v_2366 = v_9;
assign v_2368 = ~v_2367;
assign v_2369 = ~v_15;
assign v_2370 = v_15;
assign v_2372 = ~v_2371;
assign v_2373 = ~v_20;
assign v_2374 = v_20;
assign v_2376 = ~v_2375;
assign v_2377 = ~v_25;
assign v_2378 = v_25;
assign v_2379 = ~v_28;
assign v_2381 = ~v_2380;
assign v_2382 = v_2380;
assign v_2383 = ~v_33;
assign v_2385 = ~v_2384;
assign v_2386 = v_2384;
assign v_2387 = ~v_38;
assign v_2389 = ~v_2388;
assign v_2390 = v_2388;
assign v_2391 = ~v_43;
assign v_2393 = ~v_2392;
assign v_2394 = v_2392;
assign v_2395 = ~v_48;
assign v_2397 = ~v_2396;
assign v_2398 = v_2396;
assign v_2399 = ~v_53;
assign v_2401 = ~v_2400;
assign v_2402 = v_2400;
assign v_2403 = ~v_58;
assign v_2405 = ~v_2404;
assign v_2406 = v_2404;
assign v_2407 = ~v_63;
assign v_2409 = ~v_2408;
assign v_2410 = v_2408;
assign v_2411 = ~v_68;
assign v_2413 = ~v_2412;
assign v_2414 = v_2412;
assign v_2415 = ~v_73;
assign v_2417 = ~v_2416;
assign v_2418 = v_2416;
assign v_2419 = ~v_78;
assign v_2421 = ~v_2420;
assign v_2422 = v_2420;
assign v_2423 = ~v_83;
assign v_2425 = ~v_2424;
assign v_2426 = v_2424;
assign v_2427 = ~v_88;
assign v_2429 = ~v_2428;
assign v_2430 = v_2429;
assign v_2432 = v_2431;
assign v_2434 = v_2425 & v_2433;
assign v_2436 = v_83;
assign v_2438 = v_2435 & v_2437;
assign v_2440 = v_2421 & v_2439;
assign v_2442 = v_78;
assign v_2444 = v_2441 & v_2443;
assign v_2446 = v_2417 & v_2445;
assign v_2448 = v_73;
assign v_2450 = v_2447 & v_2449;
assign v_2452 = v_2413 & v_2451;
assign v_2454 = v_68;
assign v_2456 = v_2453 & v_2455;
assign v_2458 = v_2409 & v_2457;
assign v_2460 = v_63;
assign v_2462 = v_2459 & v_2461;
assign v_2464 = v_2405 & v_2463;
assign v_2466 = v_58;
assign v_2468 = v_2465 & v_2467;
assign v_2470 = v_2401 & v_2469;
assign v_2472 = v_53;
assign v_2474 = v_2471 & v_2473;
assign v_2476 = v_2397 & v_2475;
assign v_2478 = v_48;
assign v_2480 = v_2477 & v_2479;
assign v_2482 = v_2393 & v_2481;
assign v_2484 = v_43;
assign v_2486 = v_2483 & v_2485;
assign v_2488 = v_2389 & v_2487;
assign v_2490 = v_38;
assign v_2492 = v_2489 & v_2491;
assign v_2494 = v_2385 & v_2493;
assign v_2496 = v_33;
assign v_2498 = v_2495 & v_2497;
assign v_2500 = v_2381 & v_2499;
assign v_2502 = v_28;
assign v_2504 = v_2501 & v_2503;
assign v_2506 = v_2377 & v_2505;
assign v_2508 = v_2375;
assign v_2510 = v_2507 & v_2509;
assign v_2512 = v_2373 & v_2511;
assign v_2514 = v_2371;
assign v_2516 = v_2513 & v_2515;
assign v_2518 = v_2369 & v_2517;
assign v_2520 = v_2367;
assign v_2522 = v_2519 & v_2521;
assign v_2524 = v_2365 & v_2523;
assign v_2526 = v_2363;
assign v_2528 = v_2525 & v_2527;
assign v_2529 = v_2528;
assign v_2531 = v_88;
assign v_2532 = v_2428;
assign v_2533 = v_2532;
assign v_2534 = v_2531 & v_2533;
assign v_2535 = v_2534;
assign v_2536 = v_2425 & v_2535;
assign v_2538 = v_2436 & v_2537;
assign v_2539 = v_2423 & v_2535;
assign v_2541 = v_2421 & v_2540;
assign v_2543 = v_2442 & v_2542;
assign v_2544 = v_2419 & v_2540;
assign v_2546 = v_2417 & v_2545;
assign v_2548 = v_2448 & v_2547;
assign v_2549 = v_2415 & v_2545;
assign v_2551 = v_2413 & v_2550;
assign v_2553 = v_2454 & v_2552;
assign v_2554 = v_2411 & v_2550;
assign v_2556 = v_2409 & v_2555;
assign v_2558 = v_2460 & v_2557;
assign v_2559 = v_2407 & v_2555;
assign v_2561 = v_2405 & v_2560;
assign v_2563 = v_2466 & v_2562;
assign v_2564 = v_2403 & v_2560;
assign v_2566 = v_2401 & v_2565;
assign v_2568 = v_2472 & v_2567;
assign v_2569 = v_2399 & v_2565;
assign v_2571 = v_2397 & v_2570;
assign v_2573 = v_2478 & v_2572;
assign v_2574 = v_2395 & v_2570;
assign v_2576 = v_2393 & v_2575;
assign v_2578 = v_2484 & v_2577;
assign v_2579 = v_2391 & v_2575;
assign v_2581 = v_2389 & v_2580;
assign v_2583 = v_2490 & v_2582;
assign v_2584 = v_2387 & v_2580;
assign v_2586 = v_2385 & v_2585;
assign v_2588 = v_2496 & v_2587;
assign v_2589 = v_2383 & v_2585;
assign v_2591 = v_2381 & v_2590;
assign v_2593 = v_2502 & v_2592;
assign v_2594 = v_2379 & v_2590;
assign v_2596 = v_2377 & v_2595;
assign v_2598 = v_2508 & v_2597;
assign v_2599 = v_2376 & v_2595;
assign v_2601 = v_2373 & v_2600;
assign v_2603 = v_2514 & v_2602;
assign v_2604 = v_2372 & v_2600;
assign v_2606 = v_2369 & v_2605;
assign v_2608 = v_2520 & v_2607;
assign v_2609 = v_2368 & v_2605;
assign v_2611 = v_2365 & v_2610;
assign v_2613 = v_2526 & v_2612;
assign v_2614 = v_2364 & v_2610;
assign v_2616 = v_2615;
assign v_2618 = v_2530 & v_2617;
assign v_2619 = v_2618;
assign v_2621 = v_2620;
assign v_2624 = ~v_2623;
assign v_2625 = ~v_9;
assign v_2626 = v_9;
assign v_2628 = ~v_2627;
assign v_2629 = ~v_15;
assign v_2630 = v_15;
assign v_2632 = ~v_2631;
assign v_2633 = ~v_20;
assign v_2634 = v_20;
assign v_2636 = ~v_2635;
assign v_2637 = ~v_25;
assign v_2638 = v_25;
assign v_2639 = ~v_28;
assign v_2641 = ~v_2640;
assign v_2642 = v_2640;
assign v_2643 = ~v_33;
assign v_2645 = ~v_2644;
assign v_2646 = v_2644;
assign v_2647 = ~v_38;
assign v_2649 = ~v_2648;
assign v_2650 = v_2648;
assign v_2651 = ~v_43;
assign v_2653 = ~v_2652;
assign v_2654 = v_2652;
assign v_2655 = ~v_48;
assign v_2657 = ~v_2656;
assign v_2658 = v_2656;
assign v_2659 = ~v_53;
assign v_2661 = ~v_2660;
assign v_2662 = v_2660;
assign v_2663 = ~v_58;
assign v_2665 = ~v_2664;
assign v_2666 = v_2664;
assign v_2667 = ~v_63;
assign v_2669 = ~v_2668;
assign v_2670 = v_2668;
assign v_2671 = ~v_68;
assign v_2673 = ~v_2672;
assign v_2674 = v_2672;
assign v_2675 = ~v_73;
assign v_2677 = ~v_2676;
assign v_2678 = v_2676;
assign v_2679 = ~v_78;
assign v_2681 = ~v_2680;
assign v_2682 = v_2680;
assign v_2683 = ~v_83;
assign v_2685 = ~v_2684;
assign v_2686 = v_2684;
assign v_2687 = ~v_88;
assign v_2689 = ~v_2688;
assign v_2690 = v_2689;
assign v_2692 = v_2691;
assign v_2694 = v_2685 & v_2693;
assign v_2696 = v_83;
assign v_2698 = v_2695 & v_2697;
assign v_2700 = v_2681 & v_2699;
assign v_2702 = v_78;
assign v_2704 = v_2701 & v_2703;
assign v_2706 = v_2677 & v_2705;
assign v_2708 = v_73;
assign v_2710 = v_2707 & v_2709;
assign v_2712 = v_2673 & v_2711;
assign v_2714 = v_68;
assign v_2716 = v_2713 & v_2715;
assign v_2718 = v_2669 & v_2717;
assign v_2720 = v_63;
assign v_2722 = v_2719 & v_2721;
assign v_2724 = v_2665 & v_2723;
assign v_2726 = v_58;
assign v_2728 = v_2725 & v_2727;
assign v_2730 = v_2661 & v_2729;
assign v_2732 = v_53;
assign v_2734 = v_2731 & v_2733;
assign v_2736 = v_2657 & v_2735;
assign v_2738 = v_48;
assign v_2740 = v_2737 & v_2739;
assign v_2742 = v_2653 & v_2741;
assign v_2744 = v_43;
assign v_2746 = v_2743 & v_2745;
assign v_2748 = v_2649 & v_2747;
assign v_2750 = v_38;
assign v_2752 = v_2749 & v_2751;
assign v_2754 = v_2645 & v_2753;
assign v_2756 = v_33;
assign v_2758 = v_2755 & v_2757;
assign v_2760 = v_2641 & v_2759;
assign v_2762 = v_28;
assign v_2764 = v_2761 & v_2763;
assign v_2766 = v_2637 & v_2765;
assign v_2768 = v_2635;
assign v_2770 = v_2767 & v_2769;
assign v_2772 = v_2633 & v_2771;
assign v_2774 = v_2631;
assign v_2776 = v_2773 & v_2775;
assign v_2778 = v_2629 & v_2777;
assign v_2780 = v_2627;
assign v_2782 = v_2779 & v_2781;
assign v_2784 = v_2625 & v_2783;
assign v_2786 = v_2623;
assign v_2788 = v_2785 & v_2787;
assign v_2789 = v_2788;
assign v_2791 = v_88;
assign v_2792 = v_2688;
assign v_2793 = v_2792;
assign v_2794 = v_2791 & v_2793;
assign v_2795 = v_2794;
assign v_2796 = v_2685 & v_2795;
assign v_2798 = v_2696 & v_2797;
assign v_2799 = v_2683 & v_2795;
assign v_2801 = v_2681 & v_2800;
assign v_2803 = v_2702 & v_2802;
assign v_2804 = v_2679 & v_2800;
assign v_2806 = v_2677 & v_2805;
assign v_2808 = v_2708 & v_2807;
assign v_2809 = v_2675 & v_2805;
assign v_2811 = v_2673 & v_2810;
assign v_2813 = v_2714 & v_2812;
assign v_2814 = v_2671 & v_2810;
assign v_2816 = v_2669 & v_2815;
assign v_2818 = v_2720 & v_2817;
assign v_2819 = v_2667 & v_2815;
assign v_2821 = v_2665 & v_2820;
assign v_2823 = v_2726 & v_2822;
assign v_2824 = v_2663 & v_2820;
assign v_2826 = v_2661 & v_2825;
assign v_2828 = v_2732 & v_2827;
assign v_2829 = v_2659 & v_2825;
assign v_2831 = v_2657 & v_2830;
assign v_2833 = v_2738 & v_2832;
assign v_2834 = v_2655 & v_2830;
assign v_2836 = v_2653 & v_2835;
assign v_2838 = v_2744 & v_2837;
assign v_2839 = v_2651 & v_2835;
assign v_2841 = v_2649 & v_2840;
assign v_2843 = v_2750 & v_2842;
assign v_2844 = v_2647 & v_2840;
assign v_2846 = v_2645 & v_2845;
assign v_2848 = v_2756 & v_2847;
assign v_2849 = v_2643 & v_2845;
assign v_2851 = v_2641 & v_2850;
assign v_2853 = v_2762 & v_2852;
assign v_2854 = v_2639 & v_2850;
assign v_2856 = v_2637 & v_2855;
assign v_2858 = v_2768 & v_2857;
assign v_2859 = v_2636 & v_2855;
assign v_2861 = v_2633 & v_2860;
assign v_2863 = v_2774 & v_2862;
assign v_2864 = v_2632 & v_2860;
assign v_2866 = v_2629 & v_2865;
assign v_2868 = v_2780 & v_2867;
assign v_2869 = v_2628 & v_2865;
assign v_2871 = v_2625 & v_2870;
assign v_2873 = v_2786 & v_2872;
assign v_2874 = v_2624 & v_2870;
assign v_2876 = v_2875;
assign v_2878 = v_2790 & v_2877;
assign v_2879 = v_2878;
assign v_2881 = v_2880;
assign v_2884 = ~v_2883;
assign v_2885 = ~v_9;
assign v_2886 = v_9;
assign v_2888 = ~v_2887;
assign v_2889 = ~v_15;
assign v_2890 = v_15;
assign v_2892 = ~v_2891;
assign v_2893 = ~v_20;
assign v_2894 = v_20;
assign v_2896 = ~v_2895;
assign v_2897 = ~v_25;
assign v_2898 = v_25;
assign v_2899 = ~v_28;
assign v_2901 = ~v_2900;
assign v_2902 = v_2900;
assign v_2903 = ~v_33;
assign v_2905 = ~v_2904;
assign v_2906 = v_2904;
assign v_2907 = ~v_38;
assign v_2909 = ~v_2908;
assign v_2910 = v_2908;
assign v_2911 = ~v_43;
assign v_2913 = ~v_2912;
assign v_2914 = v_2912;
assign v_2915 = ~v_48;
assign v_2917 = ~v_2916;
assign v_2918 = v_2916;
assign v_2919 = ~v_53;
assign v_2921 = ~v_2920;
assign v_2922 = v_2920;
assign v_2923 = ~v_58;
assign v_2925 = ~v_2924;
assign v_2926 = v_2924;
assign v_2927 = ~v_63;
assign v_2929 = ~v_2928;
assign v_2930 = v_2928;
assign v_2931 = ~v_68;
assign v_2933 = ~v_2932;
assign v_2934 = v_2932;
assign v_2935 = ~v_73;
assign v_2937 = ~v_2936;
assign v_2938 = v_2936;
assign v_2939 = ~v_78;
assign v_2941 = ~v_2940;
assign v_2942 = v_2940;
assign v_2943 = ~v_83;
assign v_2945 = ~v_2944;
assign v_2946 = v_2944;
assign v_2947 = ~v_88;
assign v_2949 = ~v_2948;
assign v_2950 = v_2949;
assign v_2952 = v_2951;
assign v_2954 = v_2945 & v_2953;
assign v_2956 = v_83;
assign v_2958 = v_2955 & v_2957;
assign v_2960 = v_2941 & v_2959;
assign v_2962 = v_78;
assign v_2964 = v_2961 & v_2963;
assign v_2966 = v_2937 & v_2965;
assign v_2968 = v_73;
assign v_2970 = v_2967 & v_2969;
assign v_2972 = v_2933 & v_2971;
assign v_2974 = v_68;
assign v_2976 = v_2973 & v_2975;
assign v_2978 = v_2929 & v_2977;
assign v_2980 = v_63;
assign v_2982 = v_2979 & v_2981;
assign v_2984 = v_2925 & v_2983;
assign v_2986 = v_58;
assign v_2988 = v_2985 & v_2987;
assign v_2990 = v_2921 & v_2989;
assign v_2992 = v_53;
assign v_2994 = v_2991 & v_2993;
assign v_2996 = v_2917 & v_2995;
assign v_2998 = v_48;
assign v_3000 = v_2997 & v_2999;
assign v_3002 = v_2913 & v_3001;
assign v_3004 = v_43;
assign v_3006 = v_3003 & v_3005;
assign v_3008 = v_2909 & v_3007;
assign v_3010 = v_38;
assign v_3012 = v_3009 & v_3011;
assign v_3014 = v_2905 & v_3013;
assign v_3016 = v_33;
assign v_3018 = v_3015 & v_3017;
assign v_3020 = v_2901 & v_3019;
assign v_3022 = v_28;
assign v_3024 = v_3021 & v_3023;
assign v_3026 = v_2897 & v_3025;
assign v_3028 = v_2895;
assign v_3030 = v_3027 & v_3029;
assign v_3032 = v_2893 & v_3031;
assign v_3034 = v_2891;
assign v_3036 = v_3033 & v_3035;
assign v_3038 = v_2889 & v_3037;
assign v_3040 = v_2887;
assign v_3042 = v_3039 & v_3041;
assign v_3044 = v_2885 & v_3043;
assign v_3046 = v_2883;
assign v_3048 = v_3045 & v_3047;
assign v_3049 = v_3048;
assign v_3051 = v_88;
assign v_3052 = v_2948;
assign v_3053 = v_3052;
assign v_3054 = v_3051 & v_3053;
assign v_3055 = v_3054;
assign v_3056 = v_2945 & v_3055;
assign v_3058 = v_2956 & v_3057;
assign v_3059 = v_2943 & v_3055;
assign v_3061 = v_2941 & v_3060;
assign v_3063 = v_2962 & v_3062;
assign v_3064 = v_2939 & v_3060;
assign v_3066 = v_2937 & v_3065;
assign v_3068 = v_2968 & v_3067;
assign v_3069 = v_2935 & v_3065;
assign v_3071 = v_2933 & v_3070;
assign v_3073 = v_2974 & v_3072;
assign v_3074 = v_2931 & v_3070;
assign v_3076 = v_2929 & v_3075;
assign v_3078 = v_2980 & v_3077;
assign v_3079 = v_2927 & v_3075;
assign v_3081 = v_2925 & v_3080;
assign v_3083 = v_2986 & v_3082;
assign v_3084 = v_2923 & v_3080;
assign v_3086 = v_2921 & v_3085;
assign v_3088 = v_2992 & v_3087;
assign v_3089 = v_2919 & v_3085;
assign v_3091 = v_2917 & v_3090;
assign v_3093 = v_2998 & v_3092;
assign v_3094 = v_2915 & v_3090;
assign v_3096 = v_2913 & v_3095;
assign v_3098 = v_3004 & v_3097;
assign v_3099 = v_2911 & v_3095;
assign v_3101 = v_2909 & v_3100;
assign v_3103 = v_3010 & v_3102;
assign v_3104 = v_2907 & v_3100;
assign v_3106 = v_2905 & v_3105;
assign v_3108 = v_3016 & v_3107;
assign v_3109 = v_2903 & v_3105;
assign v_3111 = v_2901 & v_3110;
assign v_3113 = v_3022 & v_3112;
assign v_3114 = v_2899 & v_3110;
assign v_3116 = v_2897 & v_3115;
assign v_3118 = v_3028 & v_3117;
assign v_3119 = v_2896 & v_3115;
assign v_3121 = v_2893 & v_3120;
assign v_3123 = v_3034 & v_3122;
assign v_3124 = v_2892 & v_3120;
assign v_3126 = v_2889 & v_3125;
assign v_3128 = v_3040 & v_3127;
assign v_3129 = v_2888 & v_3125;
assign v_3131 = v_2885 & v_3130;
assign v_3133 = v_3046 & v_3132;
assign v_3134 = v_2884 & v_3130;
assign v_3136 = v_3135;
assign v_3138 = v_3050 & v_3137;
assign v_3139 = v_3138;
assign v_3141 = v_3140;
assign v_3144 = ~v_3143;
assign v_3145 = ~v_9;
assign v_3146 = v_9;
assign v_3148 = ~v_3147;
assign v_3149 = ~v_15;
assign v_3150 = v_15;
assign v_3152 = ~v_3151;
assign v_3153 = ~v_20;
assign v_3154 = v_20;
assign v_3156 = ~v_3155;
assign v_3157 = ~v_25;
assign v_3158 = v_25;
assign v_3159 = ~v_28;
assign v_3161 = ~v_3160;
assign v_3162 = v_3160;
assign v_3163 = ~v_33;
assign v_3165 = ~v_3164;
assign v_3166 = v_3164;
assign v_3167 = ~v_38;
assign v_3169 = ~v_3168;
assign v_3170 = v_3168;
assign v_3171 = ~v_43;
assign v_3173 = ~v_3172;
assign v_3174 = v_3172;
assign v_3175 = ~v_48;
assign v_3177 = ~v_3176;
assign v_3178 = v_3176;
assign v_3179 = ~v_53;
assign v_3181 = ~v_3180;
assign v_3182 = v_3180;
assign v_3183 = ~v_58;
assign v_3185 = ~v_3184;
assign v_3186 = v_3184;
assign v_3187 = ~v_63;
assign v_3189 = ~v_3188;
assign v_3190 = v_3188;
assign v_3191 = ~v_68;
assign v_3193 = ~v_3192;
assign v_3194 = v_3192;
assign v_3195 = ~v_73;
assign v_3197 = ~v_3196;
assign v_3198 = v_3196;
assign v_3199 = ~v_78;
assign v_3201 = ~v_3200;
assign v_3202 = v_3200;
assign v_3203 = ~v_83;
assign v_3205 = ~v_3204;
assign v_3206 = v_3204;
assign v_3207 = ~v_88;
assign v_3209 = ~v_3208;
assign v_3210 = v_3209;
assign v_3212 = v_3211;
assign v_3214 = v_3205 & v_3213;
assign v_3216 = v_83;
assign v_3218 = v_3215 & v_3217;
assign v_3220 = v_3201 & v_3219;
assign v_3222 = v_78;
assign v_3224 = v_3221 & v_3223;
assign v_3226 = v_3197 & v_3225;
assign v_3228 = v_73;
assign v_3230 = v_3227 & v_3229;
assign v_3232 = v_3193 & v_3231;
assign v_3234 = v_68;
assign v_3236 = v_3233 & v_3235;
assign v_3238 = v_3189 & v_3237;
assign v_3240 = v_63;
assign v_3242 = v_3239 & v_3241;
assign v_3244 = v_3185 & v_3243;
assign v_3246 = v_58;
assign v_3248 = v_3245 & v_3247;
assign v_3250 = v_3181 & v_3249;
assign v_3252 = v_53;
assign v_3254 = v_3251 & v_3253;
assign v_3256 = v_3177 & v_3255;
assign v_3258 = v_48;
assign v_3260 = v_3257 & v_3259;
assign v_3262 = v_3173 & v_3261;
assign v_3264 = v_43;
assign v_3266 = v_3263 & v_3265;
assign v_3268 = v_3169 & v_3267;
assign v_3270 = v_38;
assign v_3272 = v_3269 & v_3271;
assign v_3274 = v_3165 & v_3273;
assign v_3276 = v_33;
assign v_3278 = v_3275 & v_3277;
assign v_3280 = v_3161 & v_3279;
assign v_3282 = v_28;
assign v_3284 = v_3281 & v_3283;
assign v_3286 = v_3157 & v_3285;
assign v_3288 = v_3155;
assign v_3290 = v_3287 & v_3289;
assign v_3292 = v_3153 & v_3291;
assign v_3294 = v_3151;
assign v_3296 = v_3293 & v_3295;
assign v_3298 = v_3149 & v_3297;
assign v_3300 = v_3147;
assign v_3302 = v_3299 & v_3301;
assign v_3304 = v_3145 & v_3303;
assign v_3306 = v_3143;
assign v_3308 = v_3305 & v_3307;
assign v_3309 = v_3308;
assign v_3311 = v_88;
assign v_3312 = v_3208;
assign v_3313 = v_3312;
assign v_3314 = v_3311 & v_3313;
assign v_3315 = v_3314;
assign v_3316 = v_3205 & v_3315;
assign v_3318 = v_3216 & v_3317;
assign v_3319 = v_3203 & v_3315;
assign v_3321 = v_3201 & v_3320;
assign v_3323 = v_3222 & v_3322;
assign v_3324 = v_3199 & v_3320;
assign v_3326 = v_3197 & v_3325;
assign v_3328 = v_3228 & v_3327;
assign v_3329 = v_3195 & v_3325;
assign v_3331 = v_3193 & v_3330;
assign v_3333 = v_3234 & v_3332;
assign v_3334 = v_3191 & v_3330;
assign v_3336 = v_3189 & v_3335;
assign v_3338 = v_3240 & v_3337;
assign v_3339 = v_3187 & v_3335;
assign v_3341 = v_3185 & v_3340;
assign v_3343 = v_3246 & v_3342;
assign v_3344 = v_3183 & v_3340;
assign v_3346 = v_3181 & v_3345;
assign v_3348 = v_3252 & v_3347;
assign v_3349 = v_3179 & v_3345;
assign v_3351 = v_3177 & v_3350;
assign v_3353 = v_3258 & v_3352;
assign v_3354 = v_3175 & v_3350;
assign v_3356 = v_3173 & v_3355;
assign v_3358 = v_3264 & v_3357;
assign v_3359 = v_3171 & v_3355;
assign v_3361 = v_3169 & v_3360;
assign v_3363 = v_3270 & v_3362;
assign v_3364 = v_3167 & v_3360;
assign v_3366 = v_3165 & v_3365;
assign v_3368 = v_3276 & v_3367;
assign v_3369 = v_3163 & v_3365;
assign v_3371 = v_3161 & v_3370;
assign v_3373 = v_3282 & v_3372;
assign v_3374 = v_3159 & v_3370;
assign v_3376 = v_3157 & v_3375;
assign v_3378 = v_3288 & v_3377;
assign v_3379 = v_3156 & v_3375;
assign v_3381 = v_3153 & v_3380;
assign v_3383 = v_3294 & v_3382;
assign v_3384 = v_3152 & v_3380;
assign v_3386 = v_3149 & v_3385;
assign v_3388 = v_3300 & v_3387;
assign v_3389 = v_3148 & v_3385;
assign v_3391 = v_3145 & v_3390;
assign v_3393 = v_3306 & v_3392;
assign v_3394 = v_3144 & v_3390;
assign v_3396 = v_3395;
assign v_3398 = v_3310 & v_3397;
assign v_3399 = v_3398;
assign v_3401 = v_3400;
assign v_3404 = ~v_3403;
assign v_3405 = ~v_9;
assign v_3406 = v_9;
assign v_3408 = ~v_3407;
assign v_3409 = ~v_15;
assign v_3410 = v_15;
assign v_3412 = ~v_3411;
assign v_3413 = ~v_20;
assign v_3414 = v_20;
assign v_3416 = ~v_3415;
assign v_3417 = ~v_25;
assign v_3418 = v_25;
assign v_3419 = ~v_28;
assign v_3421 = ~v_3420;
assign v_3422 = v_3420;
assign v_3423 = ~v_33;
assign v_3425 = ~v_3424;
assign v_3426 = v_3424;
assign v_3427 = ~v_38;
assign v_3429 = ~v_3428;
assign v_3430 = v_3428;
assign v_3431 = ~v_43;
assign v_3433 = ~v_3432;
assign v_3434 = v_3432;
assign v_3435 = ~v_48;
assign v_3437 = ~v_3436;
assign v_3438 = v_3436;
assign v_3439 = ~v_53;
assign v_3441 = ~v_3440;
assign v_3442 = v_3440;
assign v_3443 = ~v_58;
assign v_3445 = ~v_3444;
assign v_3446 = v_3444;
assign v_3447 = ~v_63;
assign v_3449 = ~v_3448;
assign v_3450 = v_3448;
assign v_3451 = ~v_68;
assign v_3453 = ~v_3452;
assign v_3454 = v_3452;
assign v_3455 = ~v_73;
assign v_3457 = ~v_3456;
assign v_3458 = v_3456;
assign v_3459 = ~v_78;
assign v_3461 = ~v_3460;
assign v_3462 = v_3460;
assign v_3463 = ~v_83;
assign v_3465 = ~v_3464;
assign v_3466 = v_3464;
assign v_3467 = ~v_88;
assign v_3469 = ~v_3468;
assign v_3470 = v_3469;
assign v_3472 = v_3471;
assign v_3474 = v_3465 & v_3473;
assign v_3476 = v_83;
assign v_3478 = v_3475 & v_3477;
assign v_3480 = v_3461 & v_3479;
assign v_3482 = v_78;
assign v_3484 = v_3481 & v_3483;
assign v_3486 = v_3457 & v_3485;
assign v_3488 = v_73;
assign v_3490 = v_3487 & v_3489;
assign v_3492 = v_3453 & v_3491;
assign v_3494 = v_68;
assign v_3496 = v_3493 & v_3495;
assign v_3498 = v_3449 & v_3497;
assign v_3500 = v_63;
assign v_3502 = v_3499 & v_3501;
assign v_3504 = v_3445 & v_3503;
assign v_3506 = v_58;
assign v_3508 = v_3505 & v_3507;
assign v_3510 = v_3441 & v_3509;
assign v_3512 = v_53;
assign v_3514 = v_3511 & v_3513;
assign v_3516 = v_3437 & v_3515;
assign v_3518 = v_48;
assign v_3520 = v_3517 & v_3519;
assign v_3522 = v_3433 & v_3521;
assign v_3524 = v_43;
assign v_3526 = v_3523 & v_3525;
assign v_3528 = v_3429 & v_3527;
assign v_3530 = v_38;
assign v_3532 = v_3529 & v_3531;
assign v_3534 = v_3425 & v_3533;
assign v_3536 = v_33;
assign v_3538 = v_3535 & v_3537;
assign v_3540 = v_3421 & v_3539;
assign v_3542 = v_28;
assign v_3544 = v_3541 & v_3543;
assign v_3546 = v_3417 & v_3545;
assign v_3548 = v_3415;
assign v_3550 = v_3547 & v_3549;
assign v_3552 = v_3413 & v_3551;
assign v_3554 = v_3411;
assign v_3556 = v_3553 & v_3555;
assign v_3558 = v_3409 & v_3557;
assign v_3560 = v_3407;
assign v_3562 = v_3559 & v_3561;
assign v_3564 = v_3405 & v_3563;
assign v_3566 = v_3403;
assign v_3568 = v_3565 & v_3567;
assign v_3569 = v_3568;
assign v_3571 = v_88;
assign v_3572 = v_3468;
assign v_3573 = v_3572;
assign v_3574 = v_3571 & v_3573;
assign v_3575 = v_3574;
assign v_3576 = v_3465 & v_3575;
assign v_3578 = v_3476 & v_3577;
assign v_3579 = v_3463 & v_3575;
assign v_3581 = v_3461 & v_3580;
assign v_3583 = v_3482 & v_3582;
assign v_3584 = v_3459 & v_3580;
assign v_3586 = v_3457 & v_3585;
assign v_3588 = v_3488 & v_3587;
assign v_3589 = v_3455 & v_3585;
assign v_3591 = v_3453 & v_3590;
assign v_3593 = v_3494 & v_3592;
assign v_3594 = v_3451 & v_3590;
assign v_3596 = v_3449 & v_3595;
assign v_3598 = v_3500 & v_3597;
assign v_3599 = v_3447 & v_3595;
assign v_3601 = v_3445 & v_3600;
assign v_3603 = v_3506 & v_3602;
assign v_3604 = v_3443 & v_3600;
assign v_3606 = v_3441 & v_3605;
assign v_3608 = v_3512 & v_3607;
assign v_3609 = v_3439 & v_3605;
assign v_3611 = v_3437 & v_3610;
assign v_3613 = v_3518 & v_3612;
assign v_3614 = v_3435 & v_3610;
assign v_3616 = v_3433 & v_3615;
assign v_3618 = v_3524 & v_3617;
assign v_3619 = v_3431 & v_3615;
assign v_3621 = v_3429 & v_3620;
assign v_3623 = v_3530 & v_3622;
assign v_3624 = v_3427 & v_3620;
assign v_3626 = v_3425 & v_3625;
assign v_3628 = v_3536 & v_3627;
assign v_3629 = v_3423 & v_3625;
assign v_3631 = v_3421 & v_3630;
assign v_3633 = v_3542 & v_3632;
assign v_3634 = v_3419 & v_3630;
assign v_3636 = v_3417 & v_3635;
assign v_3638 = v_3548 & v_3637;
assign v_3639 = v_3416 & v_3635;
assign v_3641 = v_3413 & v_3640;
assign v_3643 = v_3554 & v_3642;
assign v_3644 = v_3412 & v_3640;
assign v_3646 = v_3409 & v_3645;
assign v_3648 = v_3560 & v_3647;
assign v_3649 = v_3408 & v_3645;
assign v_3651 = v_3405 & v_3650;
assign v_3653 = v_3566 & v_3652;
assign v_3654 = v_3404 & v_3650;
assign v_3656 = v_3655;
assign v_3658 = v_3570 & v_3657;
assign v_3659 = v_3658;
assign v_3661 = v_3660;
assign v_3664 = ~v_3663;
assign v_3665 = ~v_9;
assign v_3666 = v_9;
assign v_3668 = ~v_3667;
assign v_3669 = ~v_15;
assign v_3670 = v_15;
assign v_3672 = ~v_3671;
assign v_3673 = ~v_20;
assign v_3674 = v_20;
assign v_3676 = ~v_3675;
assign v_3677 = ~v_25;
assign v_3678 = v_25;
assign v_3679 = ~v_28;
assign v_3681 = ~v_3680;
assign v_3682 = v_3680;
assign v_3683 = ~v_33;
assign v_3685 = ~v_3684;
assign v_3686 = v_3684;
assign v_3687 = ~v_38;
assign v_3689 = ~v_3688;
assign v_3690 = v_3688;
assign v_3691 = ~v_43;
assign v_3693 = ~v_3692;
assign v_3694 = v_3692;
assign v_3695 = ~v_48;
assign v_3697 = ~v_3696;
assign v_3698 = v_3696;
assign v_3699 = ~v_53;
assign v_3701 = ~v_3700;
assign v_3702 = v_3700;
assign v_3703 = ~v_58;
assign v_3705 = ~v_3704;
assign v_3706 = v_3704;
assign v_3707 = ~v_63;
assign v_3709 = ~v_3708;
assign v_3710 = v_3708;
assign v_3711 = ~v_68;
assign v_3713 = ~v_3712;
assign v_3714 = v_3712;
assign v_3715 = ~v_73;
assign v_3717 = ~v_3716;
assign v_3718 = v_3716;
assign v_3719 = ~v_78;
assign v_3721 = ~v_3720;
assign v_3722 = v_3720;
assign v_3723 = ~v_83;
assign v_3725 = ~v_3724;
assign v_3726 = v_3724;
assign v_3727 = ~v_88;
assign v_3729 = ~v_3728;
assign v_3730 = v_3729;
assign v_3732 = v_3731;
assign v_3734 = v_3725 & v_3733;
assign v_3736 = v_83;
assign v_3738 = v_3735 & v_3737;
assign v_3740 = v_3721 & v_3739;
assign v_3742 = v_78;
assign v_3744 = v_3741 & v_3743;
assign v_3746 = v_3717 & v_3745;
assign v_3748 = v_73;
assign v_3750 = v_3747 & v_3749;
assign v_3752 = v_3713 & v_3751;
assign v_3754 = v_68;
assign v_3756 = v_3753 & v_3755;
assign v_3758 = v_3709 & v_3757;
assign v_3760 = v_63;
assign v_3762 = v_3759 & v_3761;
assign v_3764 = v_3705 & v_3763;
assign v_3766 = v_58;
assign v_3768 = v_3765 & v_3767;
assign v_3770 = v_3701 & v_3769;
assign v_3772 = v_53;
assign v_3774 = v_3771 & v_3773;
assign v_3776 = v_3697 & v_3775;
assign v_3778 = v_48;
assign v_3780 = v_3777 & v_3779;
assign v_3782 = v_3693 & v_3781;
assign v_3784 = v_43;
assign v_3786 = v_3783 & v_3785;
assign v_3788 = v_3689 & v_3787;
assign v_3790 = v_38;
assign v_3792 = v_3789 & v_3791;
assign v_3794 = v_3685 & v_3793;
assign v_3796 = v_33;
assign v_3798 = v_3795 & v_3797;
assign v_3800 = v_3681 & v_3799;
assign v_3802 = v_28;
assign v_3804 = v_3801 & v_3803;
assign v_3806 = v_3677 & v_3805;
assign v_3808 = v_3675;
assign v_3810 = v_3807 & v_3809;
assign v_3812 = v_3673 & v_3811;
assign v_3814 = v_3671;
assign v_3816 = v_3813 & v_3815;
assign v_3818 = v_3669 & v_3817;
assign v_3820 = v_3667;
assign v_3822 = v_3819 & v_3821;
assign v_3824 = v_3665 & v_3823;
assign v_3826 = v_3663;
assign v_3828 = v_3825 & v_3827;
assign v_3829 = v_3828;
assign v_3831 = v_88;
assign v_3832 = v_3728;
assign v_3833 = v_3832;
assign v_3834 = v_3831 & v_3833;
assign v_3835 = v_3834;
assign v_3836 = v_3725 & v_3835;
assign v_3838 = v_3736 & v_3837;
assign v_3839 = v_3723 & v_3835;
assign v_3841 = v_3721 & v_3840;
assign v_3843 = v_3742 & v_3842;
assign v_3844 = v_3719 & v_3840;
assign v_3846 = v_3717 & v_3845;
assign v_3848 = v_3748 & v_3847;
assign v_3849 = v_3715 & v_3845;
assign v_3851 = v_3713 & v_3850;
assign v_3853 = v_3754 & v_3852;
assign v_3854 = v_3711 & v_3850;
assign v_3856 = v_3709 & v_3855;
assign v_3858 = v_3760 & v_3857;
assign v_3859 = v_3707 & v_3855;
assign v_3861 = v_3705 & v_3860;
assign v_3863 = v_3766 & v_3862;
assign v_3864 = v_3703 & v_3860;
assign v_3866 = v_3701 & v_3865;
assign v_3868 = v_3772 & v_3867;
assign v_3869 = v_3699 & v_3865;
assign v_3871 = v_3697 & v_3870;
assign v_3873 = v_3778 & v_3872;
assign v_3874 = v_3695 & v_3870;
assign v_3876 = v_3693 & v_3875;
assign v_3878 = v_3784 & v_3877;
assign v_3879 = v_3691 & v_3875;
assign v_3881 = v_3689 & v_3880;
assign v_3883 = v_3790 & v_3882;
assign v_3884 = v_3687 & v_3880;
assign v_3886 = v_3685 & v_3885;
assign v_3888 = v_3796 & v_3887;
assign v_3889 = v_3683 & v_3885;
assign v_3891 = v_3681 & v_3890;
assign v_3893 = v_3802 & v_3892;
assign v_3894 = v_3679 & v_3890;
assign v_3896 = v_3677 & v_3895;
assign v_3898 = v_3808 & v_3897;
assign v_3899 = v_3676 & v_3895;
assign v_3901 = v_3673 & v_3900;
assign v_3903 = v_3814 & v_3902;
assign v_3904 = v_3672 & v_3900;
assign v_3906 = v_3669 & v_3905;
assign v_3908 = v_3820 & v_3907;
assign v_3909 = v_3668 & v_3905;
assign v_3911 = v_3665 & v_3910;
assign v_3913 = v_3826 & v_3912;
assign v_3914 = v_3664 & v_3910;
assign v_3916 = v_3915;
assign v_3918 = v_3830 & v_3917;
assign v_3919 = v_3918;
assign v_3921 = v_3920;
assign v_3924 = ~v_3923;
assign v_3925 = ~v_9;
assign v_3926 = v_9;
assign v_3928 = ~v_3927;
assign v_3929 = ~v_15;
assign v_3930 = v_15;
assign v_3932 = ~v_3931;
assign v_3933 = ~v_20;
assign v_3934 = v_20;
assign v_3936 = ~v_3935;
assign v_3937 = ~v_25;
assign v_3938 = v_25;
assign v_3939 = ~v_28;
assign v_3941 = ~v_3940;
assign v_3942 = v_3940;
assign v_3943 = ~v_33;
assign v_3945 = ~v_3944;
assign v_3946 = v_3944;
assign v_3947 = ~v_38;
assign v_3949 = ~v_3948;
assign v_3950 = v_3948;
assign v_3951 = ~v_43;
assign v_3953 = ~v_3952;
assign v_3954 = v_3952;
assign v_3955 = ~v_48;
assign v_3957 = ~v_3956;
assign v_3958 = v_3956;
assign v_3959 = ~v_53;
assign v_3961 = ~v_3960;
assign v_3962 = v_3960;
assign v_3963 = ~v_58;
assign v_3965 = ~v_3964;
assign v_3966 = v_3964;
assign v_3967 = ~v_63;
assign v_3969 = ~v_3968;
assign v_3970 = v_3968;
assign v_3971 = ~v_68;
assign v_3973 = ~v_3972;
assign v_3974 = v_3972;
assign v_3975 = ~v_73;
assign v_3977 = ~v_3976;
assign v_3978 = v_3976;
assign v_3979 = ~v_78;
assign v_3981 = ~v_3980;
assign v_3982 = v_3980;
assign v_3983 = ~v_83;
assign v_3985 = ~v_3984;
assign v_3986 = v_3984;
assign v_3987 = ~v_88;
assign v_3989 = ~v_3988;
assign v_3990 = v_3989;
assign v_3992 = v_3991;
assign v_3994 = v_3985 & v_3993;
assign v_3996 = v_83;
assign v_3998 = v_3995 & v_3997;
assign v_4000 = v_3981 & v_3999;
assign v_4002 = v_78;
assign v_4004 = v_4001 & v_4003;
assign v_4006 = v_3977 & v_4005;
assign v_4008 = v_73;
assign v_4010 = v_4007 & v_4009;
assign v_4012 = v_3973 & v_4011;
assign v_4014 = v_68;
assign v_4016 = v_4013 & v_4015;
assign v_4018 = v_3969 & v_4017;
assign v_4020 = v_63;
assign v_4022 = v_4019 & v_4021;
assign v_4024 = v_3965 & v_4023;
assign v_4026 = v_58;
assign v_4028 = v_4025 & v_4027;
assign v_4030 = v_3961 & v_4029;
assign v_4032 = v_53;
assign v_4034 = v_4031 & v_4033;
assign v_4036 = v_3957 & v_4035;
assign v_4038 = v_48;
assign v_4040 = v_4037 & v_4039;
assign v_4042 = v_3953 & v_4041;
assign v_4044 = v_43;
assign v_4046 = v_4043 & v_4045;
assign v_4048 = v_3949 & v_4047;
assign v_4050 = v_38;
assign v_4052 = v_4049 & v_4051;
assign v_4054 = v_3945 & v_4053;
assign v_4056 = v_33;
assign v_4058 = v_4055 & v_4057;
assign v_4060 = v_3941 & v_4059;
assign v_4062 = v_28;
assign v_4064 = v_4061 & v_4063;
assign v_4066 = v_3937 & v_4065;
assign v_4068 = v_3935;
assign v_4070 = v_4067 & v_4069;
assign v_4072 = v_3933 & v_4071;
assign v_4074 = v_3931;
assign v_4076 = v_4073 & v_4075;
assign v_4078 = v_3929 & v_4077;
assign v_4080 = v_3927;
assign v_4082 = v_4079 & v_4081;
assign v_4084 = v_3925 & v_4083;
assign v_4086 = v_3923;
assign v_4088 = v_4085 & v_4087;
assign v_4089 = v_4088;
assign v_4091 = v_88;
assign v_4092 = v_3988;
assign v_4093 = v_4092;
assign v_4094 = v_4091 & v_4093;
assign v_4095 = v_4094;
assign v_4096 = v_3985 & v_4095;
assign v_4098 = v_3996 & v_4097;
assign v_4099 = v_3983 & v_4095;
assign v_4101 = v_3981 & v_4100;
assign v_4103 = v_4002 & v_4102;
assign v_4104 = v_3979 & v_4100;
assign v_4106 = v_3977 & v_4105;
assign v_4108 = v_4008 & v_4107;
assign v_4109 = v_3975 & v_4105;
assign v_4111 = v_3973 & v_4110;
assign v_4113 = v_4014 & v_4112;
assign v_4114 = v_3971 & v_4110;
assign v_4116 = v_3969 & v_4115;
assign v_4118 = v_4020 & v_4117;
assign v_4119 = v_3967 & v_4115;
assign v_4121 = v_3965 & v_4120;
assign v_4123 = v_4026 & v_4122;
assign v_4124 = v_3963 & v_4120;
assign v_4126 = v_3961 & v_4125;
assign v_4128 = v_4032 & v_4127;
assign v_4129 = v_3959 & v_4125;
assign v_4131 = v_3957 & v_4130;
assign v_4133 = v_4038 & v_4132;
assign v_4134 = v_3955 & v_4130;
assign v_4136 = v_3953 & v_4135;
assign v_4138 = v_4044 & v_4137;
assign v_4139 = v_3951 & v_4135;
assign v_4141 = v_3949 & v_4140;
assign v_4143 = v_4050 & v_4142;
assign v_4144 = v_3947 & v_4140;
assign v_4146 = v_3945 & v_4145;
assign v_4148 = v_4056 & v_4147;
assign v_4149 = v_3943 & v_4145;
assign v_4151 = v_3941 & v_4150;
assign v_4153 = v_4062 & v_4152;
assign v_4154 = v_3939 & v_4150;
assign v_4156 = v_3937 & v_4155;
assign v_4158 = v_4068 & v_4157;
assign v_4159 = v_3936 & v_4155;
assign v_4161 = v_3933 & v_4160;
assign v_4163 = v_4074 & v_4162;
assign v_4164 = v_3932 & v_4160;
assign v_4166 = v_3929 & v_4165;
assign v_4168 = v_4080 & v_4167;
assign v_4169 = v_3928 & v_4165;
assign v_4171 = v_3925 & v_4170;
assign v_4173 = v_4086 & v_4172;
assign v_4174 = v_3924 & v_4170;
assign v_4176 = v_4175;
assign v_4178 = v_4090 & v_4177;
assign v_4179 = v_4178;
assign v_4181 = v_4180;
assign v_4183 = ~v_4182;
assign v_4184 = ~v_9;
assign v_4185 = v_9;
assign v_4187 = ~v_4186;
assign v_4188 = ~v_15;
assign v_4189 = v_15;
assign v_4191 = ~v_4190;
assign v_4192 = ~v_20;
assign v_4193 = v_20;
assign v_4195 = ~v_4194;
assign v_4196 = ~v_25;
assign v_4197 = v_25;
assign v_4198 = ~v_28;
assign v_4200 = ~v_4199;
assign v_4201 = v_4199;
assign v_4202 = ~v_33;
assign v_4204 = ~v_4203;
assign v_4205 = v_4203;
assign v_4206 = ~v_38;
assign v_4208 = ~v_4207;
assign v_4209 = v_4207;
assign v_4210 = ~v_43;
assign v_4212 = ~v_4211;
assign v_4213 = v_4211;
assign v_4214 = ~v_48;
assign v_4216 = ~v_4215;
assign v_4217 = v_4215;
assign v_4218 = ~v_53;
assign v_4220 = ~v_4219;
assign v_4221 = v_4219;
assign v_4222 = ~v_58;
assign v_4224 = ~v_4223;
assign v_4225 = v_4223;
assign v_4226 = ~v_63;
assign v_4228 = ~v_4227;
assign v_4229 = v_4227;
assign v_4230 = ~v_68;
assign v_4232 = ~v_4231;
assign v_4233 = v_4231;
assign v_4234 = ~v_73;
assign v_4236 = ~v_4235;
assign v_4237 = v_4235;
assign v_4238 = ~v_78;
assign v_4240 = ~v_4239;
assign v_4241 = v_4239;
assign v_4242 = ~v_83;
assign v_4244 = ~v_4243;
assign v_4245 = v_4243;
assign v_4246 = ~v_88;
assign v_4248 = ~v_4247;
assign v_4249 = v_4248;
assign v_4251 = v_4250;
assign v_4253 = v_4244 & v_4252;
assign v_4255 = v_83;
assign v_4257 = v_4254 & v_4256;
assign v_4259 = v_4240 & v_4258;
assign v_4261 = v_78;
assign v_4263 = v_4260 & v_4262;
assign v_4265 = v_4236 & v_4264;
assign v_4267 = v_73;
assign v_4269 = v_4266 & v_4268;
assign v_4271 = v_4232 & v_4270;
assign v_4273 = v_68;
assign v_4275 = v_4272 & v_4274;
assign v_4277 = v_4228 & v_4276;
assign v_4279 = v_63;
assign v_4281 = v_4278 & v_4280;
assign v_4283 = v_4224 & v_4282;
assign v_4285 = v_58;
assign v_4287 = v_4284 & v_4286;
assign v_4289 = v_4220 & v_4288;
assign v_4291 = v_53;
assign v_4293 = v_4290 & v_4292;
assign v_4295 = v_4216 & v_4294;
assign v_4297 = v_48;
assign v_4299 = v_4296 & v_4298;
assign v_4301 = v_4212 & v_4300;
assign v_4303 = v_43;
assign v_4305 = v_4302 & v_4304;
assign v_4307 = v_4208 & v_4306;
assign v_4309 = v_38;
assign v_4311 = v_4308 & v_4310;
assign v_4313 = v_4204 & v_4312;
assign v_4315 = v_33;
assign v_4317 = v_4314 & v_4316;
assign v_4319 = v_4200 & v_4318;
assign v_4321 = v_28;
assign v_4323 = v_4320 & v_4322;
assign v_4325 = v_4196 & v_4324;
assign v_4327 = v_4194;
assign v_4329 = v_4326 & v_4328;
assign v_4331 = v_4192 & v_4330;
assign v_4333 = v_4190;
assign v_4335 = v_4332 & v_4334;
assign v_4337 = v_4188 & v_4336;
assign v_4339 = v_4186;
assign v_4341 = v_4338 & v_4340;
assign v_4343 = v_4184 & v_4342;
assign v_4345 = v_4182;
assign v_4347 = v_4344 & v_4346;
assign v_4349 = ~v_4348;
assign v_4351 = v_88;
assign v_4352 = v_4247;
assign v_4353 = v_4352;
assign v_4354 = v_4351 & v_4353;
assign v_4355 = v_4354;
assign v_4356 = v_4244 & v_4355;
assign v_4358 = v_4255 & v_4357;
assign v_4359 = v_4242 & v_4355;
assign v_4361 = v_4240 & v_4360;
assign v_4363 = v_4261 & v_4362;
assign v_4364 = v_4238 & v_4360;
assign v_4366 = v_4236 & v_4365;
assign v_4368 = v_4267 & v_4367;
assign v_4369 = v_4234 & v_4365;
assign v_4371 = v_4232 & v_4370;
assign v_4373 = v_4273 & v_4372;
assign v_4374 = v_4230 & v_4370;
assign v_4376 = v_4228 & v_4375;
assign v_4378 = v_4279 & v_4377;
assign v_4379 = v_4226 & v_4375;
assign v_4381 = v_4224 & v_4380;
assign v_4383 = v_4285 & v_4382;
assign v_4384 = v_4222 & v_4380;
assign v_4386 = v_4220 & v_4385;
assign v_4388 = v_4291 & v_4387;
assign v_4389 = v_4218 & v_4385;
assign v_4391 = v_4216 & v_4390;
assign v_4393 = v_4297 & v_4392;
assign v_4394 = v_4214 & v_4390;
assign v_4396 = v_4212 & v_4395;
assign v_4398 = v_4303 & v_4397;
assign v_4399 = v_4210 & v_4395;
assign v_4401 = v_4208 & v_4400;
assign v_4403 = v_4309 & v_4402;
assign v_4404 = v_4206 & v_4400;
assign v_4406 = v_4204 & v_4405;
assign v_4408 = v_4315 & v_4407;
assign v_4409 = v_4202 & v_4405;
assign v_4411 = v_4200 & v_4410;
assign v_4413 = v_4321 & v_4412;
assign v_4414 = v_4198 & v_4410;
assign v_4416 = v_4196 & v_4415;
assign v_4418 = v_4327 & v_4417;
assign v_4419 = v_4195 & v_4415;
assign v_4421 = v_4192 & v_4420;
assign v_4423 = v_4333 & v_4422;
assign v_4424 = v_4191 & v_4420;
assign v_4426 = v_4188 & v_4425;
assign v_4428 = v_4339 & v_4427;
assign v_4429 = v_4187 & v_4425;
assign v_4431 = v_4184 & v_4430;
assign v_4433 = v_4345 & v_4432;
assign v_4434 = v_4183 & v_4430;
assign v_4436 = v_4348;
assign v_4438 = v_4350 & v_4437;
assign v_4439 = v_4438;
assign v_4441 = v_4440;
assign v_4443 = ~v_6;
assign v_4445 = ~v_4444;
assign v_4446 = v_4444;
assign v_4447 = ~v_13;
assign v_4449 = ~v_4448;
assign v_4450 = v_4448;
assign v_4451 = ~v_18;
assign v_4453 = ~v_4452;
assign v_4454 = v_4452;
assign v_4455 = ~v_23;
assign v_4457 = ~v_4456;
assign v_4458 = v_4456;
assign v_4460 = ~v_4459;
assign v_4461 = ~v_30;
assign v_4462 = v_30;
assign v_4464 = ~v_4463;
assign v_4465 = ~v_35;
assign v_4466 = v_35;
assign v_4468 = ~v_4467;
assign v_4469 = ~v_40;
assign v_4470 = v_40;
assign v_4472 = ~v_4471;
assign v_4473 = ~v_45;
assign v_4474 = v_45;
assign v_4476 = ~v_4475;
assign v_4477 = ~v_50;
assign v_4478 = v_50;
assign v_4480 = ~v_4479;
assign v_4481 = ~v_55;
assign v_4482 = v_55;
assign v_4484 = ~v_4483;
assign v_4485 = ~v_60;
assign v_4486 = v_60;
assign v_4488 = ~v_4487;
assign v_4489 = ~v_65;
assign v_4490 = v_65;
assign v_4492 = ~v_4491;
assign v_4493 = ~v_70;
assign v_4494 = v_70;
assign v_4496 = ~v_4495;
assign v_4497 = ~v_75;
assign v_4498 = v_75;
assign v_4500 = ~v_4499;
assign v_4501 = ~v_80;
assign v_4502 = v_80;
assign v_4504 = ~v_4503;
assign v_4505 = ~v_85;
assign v_4506 = v_85;
assign v_4508 = ~v_4507;
assign v_4509 = ~v_90;
assign v_4510 = v_4509;
assign v_4512 = v_4511;
assign v_4514 = v_4505 & v_4513;
assign v_4516 = v_4503;
assign v_4518 = v_4515 & v_4517;
assign v_4520 = v_4501 & v_4519;
assign v_4522 = v_4499;
assign v_4524 = v_4521 & v_4523;
assign v_4526 = v_4497 & v_4525;
assign v_4528 = v_4495;
assign v_4530 = v_4527 & v_4529;
assign v_4532 = v_4493 & v_4531;
assign v_4534 = v_4491;
assign v_4536 = v_4533 & v_4535;
assign v_4538 = v_4489 & v_4537;
assign v_4540 = v_4487;
assign v_4542 = v_4539 & v_4541;
assign v_4544 = v_4485 & v_4543;
assign v_4546 = v_4483;
assign v_4548 = v_4545 & v_4547;
assign v_4550 = v_4481 & v_4549;
assign v_4552 = v_4479;
assign v_4554 = v_4551 & v_4553;
assign v_4556 = v_4477 & v_4555;
assign v_4558 = v_4475;
assign v_4560 = v_4557 & v_4559;
assign v_4562 = v_4473 & v_4561;
assign v_4564 = v_4471;
assign v_4566 = v_4563 & v_4565;
assign v_4568 = v_4469 & v_4567;
assign v_4570 = v_4467;
assign v_4572 = v_4569 & v_4571;
assign v_4574 = v_4465 & v_4573;
assign v_4576 = v_4463;
assign v_4578 = v_4575 & v_4577;
assign v_4580 = v_4461 & v_4579;
assign v_4582 = v_4459;
assign v_4584 = v_4581 & v_4583;
assign v_4586 = v_4457 & v_4585;
assign v_4588 = v_23;
assign v_4590 = v_4587 & v_4589;
assign v_4592 = v_4453 & v_4591;
assign v_4594 = v_18;
assign v_4596 = v_4593 & v_4595;
assign v_4598 = v_4449 & v_4597;
assign v_4600 = v_13;
assign v_4602 = v_4599 & v_4601;
assign v_4604 = v_4445 & v_4603;
assign v_4606 = v_6;
assign v_4608 = v_4605 & v_4607;
assign v_4609 = v_4608;
assign v_4611 = v_4507;
assign v_4612 = v_90;
assign v_4613 = v_4612;
assign v_4614 = v_4611 & v_4613;
assign v_4615 = v_4614;
assign v_4616 = v_4505 & v_4615;
assign v_4618 = v_4516 & v_4617;
assign v_4619 = v_4504 & v_4615;
assign v_4621 = v_4501 & v_4620;
assign v_4623 = v_4522 & v_4622;
assign v_4624 = v_4500 & v_4620;
assign v_4626 = v_4497 & v_4625;
assign v_4628 = v_4528 & v_4627;
assign v_4629 = v_4496 & v_4625;
assign v_4631 = v_4493 & v_4630;
assign v_4633 = v_4534 & v_4632;
assign v_4634 = v_4492 & v_4630;
assign v_4636 = v_4489 & v_4635;
assign v_4638 = v_4540 & v_4637;
assign v_4639 = v_4488 & v_4635;
assign v_4641 = v_4485 & v_4640;
assign v_4643 = v_4546 & v_4642;
assign v_4644 = v_4484 & v_4640;
assign v_4646 = v_4481 & v_4645;
assign v_4648 = v_4552 & v_4647;
assign v_4649 = v_4480 & v_4645;
assign v_4651 = v_4477 & v_4650;
assign v_4653 = v_4558 & v_4652;
assign v_4654 = v_4476 & v_4650;
assign v_4656 = v_4473 & v_4655;
assign v_4658 = v_4564 & v_4657;
assign v_4659 = v_4472 & v_4655;
assign v_4661 = v_4469 & v_4660;
assign v_4663 = v_4570 & v_4662;
assign v_4664 = v_4468 & v_4660;
assign v_4666 = v_4465 & v_4665;
assign v_4668 = v_4576 & v_4667;
assign v_4669 = v_4464 & v_4665;
assign v_4671 = v_4461 & v_4670;
assign v_4673 = v_4582 & v_4672;
assign v_4674 = v_4460 & v_4670;
assign v_4676 = v_4457 & v_4675;
assign v_4678 = v_4588 & v_4677;
assign v_4679 = v_4455 & v_4675;
assign v_4681 = v_4453 & v_4680;
assign v_4683 = v_4594 & v_4682;
assign v_4684 = v_4451 & v_4680;
assign v_4686 = v_4449 & v_4685;
assign v_4688 = v_4600 & v_4687;
assign v_4689 = v_4447 & v_4685;
assign v_4691 = v_4445 & v_4690;
assign v_4693 = v_4606 & v_4692;
assign v_4694 = v_4443 & v_4690;
assign v_4696 = v_4695;
assign v_4698 = v_4610 & v_4697;
assign v_4699 = v_4698;
assign v_4701 = v_4700;
assign v_4703 = ~v_283;
assign v_4704 = ~v_4444;
assign v_4705 = v_4444;
assign v_4706 = ~v_287;
assign v_4707 = ~v_4448;
assign v_4708 = v_4448;
assign v_4709 = ~v_291;
assign v_4710 = ~v_4452;
assign v_4711 = v_4452;
assign v_4712 = ~v_295;
assign v_4713 = ~v_4456;
assign v_4714 = v_4456;
assign v_4715 = ~v_4459;
assign v_4716 = ~v_300;
assign v_4717 = v_300;
assign v_4718 = ~v_4463;
assign v_4719 = ~v_304;
assign v_4720 = v_304;
assign v_4721 = ~v_4467;
assign v_4722 = ~v_308;
assign v_4723 = v_308;
assign v_4724 = ~v_4471;
assign v_4725 = ~v_312;
assign v_4726 = v_312;
assign v_4727 = ~v_4475;
assign v_4728 = ~v_316;
assign v_4729 = v_316;
assign v_4730 = ~v_4479;
assign v_4731 = ~v_320;
assign v_4732 = v_320;
assign v_4733 = ~v_4483;
assign v_4734 = ~v_324;
assign v_4735 = v_324;
assign v_4736 = ~v_4487;
assign v_4737 = ~v_328;
assign v_4738 = v_328;
assign v_4739 = ~v_4491;
assign v_4740 = ~v_332;
assign v_4741 = v_332;
assign v_4742 = ~v_4495;
assign v_4743 = ~v_336;
assign v_4744 = v_336;
assign v_4745 = ~v_4499;
assign v_4746 = ~v_340;
assign v_4747 = v_340;
assign v_4748 = ~v_4503;
assign v_4749 = ~v_344;
assign v_4750 = v_344;
assign v_4751 = ~v_4507;
assign v_4752 = ~v_348;
assign v_4753 = v_4752;
assign v_4755 = v_4754;
assign v_4757 = v_4749 & v_4756;
assign v_4759 = v_4503;
assign v_4761 = v_4758 & v_4760;
assign v_4763 = v_4746 & v_4762;
assign v_4765 = v_4499;
assign v_4767 = v_4764 & v_4766;
assign v_4769 = v_4743 & v_4768;
assign v_4771 = v_4495;
assign v_4773 = v_4770 & v_4772;
assign v_4775 = v_4740 & v_4774;
assign v_4777 = v_4491;
assign v_4779 = v_4776 & v_4778;
assign v_4781 = v_4737 & v_4780;
assign v_4783 = v_4487;
assign v_4785 = v_4782 & v_4784;
assign v_4787 = v_4734 & v_4786;
assign v_4789 = v_4483;
assign v_4791 = v_4788 & v_4790;
assign v_4793 = v_4731 & v_4792;
assign v_4795 = v_4479;
assign v_4797 = v_4794 & v_4796;
assign v_4799 = v_4728 & v_4798;
assign v_4801 = v_4475;
assign v_4803 = v_4800 & v_4802;
assign v_4805 = v_4725 & v_4804;
assign v_4807 = v_4471;
assign v_4809 = v_4806 & v_4808;
assign v_4811 = v_4722 & v_4810;
assign v_4813 = v_4467;
assign v_4815 = v_4812 & v_4814;
assign v_4817 = v_4719 & v_4816;
assign v_4819 = v_4463;
assign v_4821 = v_4818 & v_4820;
assign v_4823 = v_4716 & v_4822;
assign v_4825 = v_4459;
assign v_4827 = v_4824 & v_4826;
assign v_4829 = v_4713 & v_4828;
assign v_4831 = v_295;
assign v_4833 = v_4830 & v_4832;
assign v_4835 = v_4710 & v_4834;
assign v_4837 = v_291;
assign v_4839 = v_4836 & v_4838;
assign v_4841 = v_4707 & v_4840;
assign v_4843 = v_287;
assign v_4845 = v_4842 & v_4844;
assign v_4847 = v_4704 & v_4846;
assign v_4849 = v_283;
assign v_4851 = v_4848 & v_4850;
assign v_4852 = v_4851;
assign v_4854 = v_4507;
assign v_4855 = v_348;
assign v_4856 = v_4855;
assign v_4857 = v_4854 & v_4856;
assign v_4858 = v_4857;
assign v_4859 = v_4749 & v_4858;
assign v_4861 = v_4759 & v_4860;
assign v_4862 = v_4748 & v_4858;
assign v_4864 = v_4746 & v_4863;
assign v_4866 = v_4765 & v_4865;
assign v_4867 = v_4745 & v_4863;
assign v_4869 = v_4743 & v_4868;
assign v_4871 = v_4771 & v_4870;
assign v_4872 = v_4742 & v_4868;
assign v_4874 = v_4740 & v_4873;
assign v_4876 = v_4777 & v_4875;
assign v_4877 = v_4739 & v_4873;
assign v_4879 = v_4737 & v_4878;
assign v_4881 = v_4783 & v_4880;
assign v_4882 = v_4736 & v_4878;
assign v_4884 = v_4734 & v_4883;
assign v_4886 = v_4789 & v_4885;
assign v_4887 = v_4733 & v_4883;
assign v_4889 = v_4731 & v_4888;
assign v_4891 = v_4795 & v_4890;
assign v_4892 = v_4730 & v_4888;
assign v_4894 = v_4728 & v_4893;
assign v_4896 = v_4801 & v_4895;
assign v_4897 = v_4727 & v_4893;
assign v_4899 = v_4725 & v_4898;
assign v_4901 = v_4807 & v_4900;
assign v_4902 = v_4724 & v_4898;
assign v_4904 = v_4722 & v_4903;
assign v_4906 = v_4813 & v_4905;
assign v_4907 = v_4721 & v_4903;
assign v_4909 = v_4719 & v_4908;
assign v_4911 = v_4819 & v_4910;
assign v_4912 = v_4718 & v_4908;
assign v_4914 = v_4716 & v_4913;
assign v_4916 = v_4825 & v_4915;
assign v_4917 = v_4715 & v_4913;
assign v_4919 = v_4713 & v_4918;
assign v_4921 = v_4831 & v_4920;
assign v_4922 = v_4712 & v_4918;
assign v_4924 = v_4710 & v_4923;
assign v_4926 = v_4837 & v_4925;
assign v_4927 = v_4709 & v_4923;
assign v_4929 = v_4707 & v_4928;
assign v_4931 = v_4843 & v_4930;
assign v_4932 = v_4706 & v_4928;
assign v_4934 = v_4704 & v_4933;
assign v_4936 = v_4849 & v_4935;
assign v_4937 = v_4703 & v_4933;
assign v_4939 = v_4938;
assign v_4941 = v_4853 & v_4940;
assign v_4942 = v_4941;
assign v_4944 = v_4943;
assign v_4946 = ~v_543;
assign v_4947 = ~v_4444;
assign v_4948 = v_4444;
assign v_4949 = ~v_547;
assign v_4950 = ~v_4448;
assign v_4951 = v_4448;
assign v_4952 = ~v_551;
assign v_4953 = ~v_4452;
assign v_4954 = v_4452;
assign v_4955 = ~v_555;
assign v_4956 = ~v_4456;
assign v_4957 = v_4456;
assign v_4958 = ~v_4459;
assign v_4959 = ~v_560;
assign v_4960 = v_560;
assign v_4961 = ~v_4463;
assign v_4962 = ~v_564;
assign v_4963 = v_564;
assign v_4964 = ~v_4467;
assign v_4965 = ~v_568;
assign v_4966 = v_568;
assign v_4967 = ~v_4471;
assign v_4968 = ~v_572;
assign v_4969 = v_572;
assign v_4970 = ~v_4475;
assign v_4971 = ~v_576;
assign v_4972 = v_576;
assign v_4973 = ~v_4479;
assign v_4974 = ~v_580;
assign v_4975 = v_580;
assign v_4976 = ~v_4483;
assign v_4977 = ~v_584;
assign v_4978 = v_584;
assign v_4979 = ~v_4487;
assign v_4980 = ~v_588;
assign v_4981 = v_588;
assign v_4982 = ~v_4491;
assign v_4983 = ~v_592;
assign v_4984 = v_592;
assign v_4985 = ~v_4495;
assign v_4986 = ~v_596;
assign v_4987 = v_596;
assign v_4988 = ~v_4499;
assign v_4989 = ~v_600;
assign v_4990 = v_600;
assign v_4991 = ~v_4503;
assign v_4992 = ~v_604;
assign v_4993 = v_604;
assign v_4994 = ~v_4507;
assign v_4995 = ~v_608;
assign v_4996 = v_4995;
assign v_4998 = v_4997;
assign v_5000 = v_4992 & v_4999;
assign v_5002 = v_4503;
assign v_5004 = v_5001 & v_5003;
assign v_5006 = v_4989 & v_5005;
assign v_5008 = v_4499;
assign v_5010 = v_5007 & v_5009;
assign v_5012 = v_4986 & v_5011;
assign v_5014 = v_4495;
assign v_5016 = v_5013 & v_5015;
assign v_5018 = v_4983 & v_5017;
assign v_5020 = v_4491;
assign v_5022 = v_5019 & v_5021;
assign v_5024 = v_4980 & v_5023;
assign v_5026 = v_4487;
assign v_5028 = v_5025 & v_5027;
assign v_5030 = v_4977 & v_5029;
assign v_5032 = v_4483;
assign v_5034 = v_5031 & v_5033;
assign v_5036 = v_4974 & v_5035;
assign v_5038 = v_4479;
assign v_5040 = v_5037 & v_5039;
assign v_5042 = v_4971 & v_5041;
assign v_5044 = v_4475;
assign v_5046 = v_5043 & v_5045;
assign v_5048 = v_4968 & v_5047;
assign v_5050 = v_4471;
assign v_5052 = v_5049 & v_5051;
assign v_5054 = v_4965 & v_5053;
assign v_5056 = v_4467;
assign v_5058 = v_5055 & v_5057;
assign v_5060 = v_4962 & v_5059;
assign v_5062 = v_4463;
assign v_5064 = v_5061 & v_5063;
assign v_5066 = v_4959 & v_5065;
assign v_5068 = v_4459;
assign v_5070 = v_5067 & v_5069;
assign v_5072 = v_4956 & v_5071;
assign v_5074 = v_555;
assign v_5076 = v_5073 & v_5075;
assign v_5078 = v_4953 & v_5077;
assign v_5080 = v_551;
assign v_5082 = v_5079 & v_5081;
assign v_5084 = v_4950 & v_5083;
assign v_5086 = v_547;
assign v_5088 = v_5085 & v_5087;
assign v_5090 = v_4947 & v_5089;
assign v_5092 = v_543;
assign v_5094 = v_5091 & v_5093;
assign v_5095 = v_5094;
assign v_5097 = v_4507;
assign v_5098 = v_608;
assign v_5099 = v_5098;
assign v_5100 = v_5097 & v_5099;
assign v_5101 = v_5100;
assign v_5102 = v_4992 & v_5101;
assign v_5104 = v_5002 & v_5103;
assign v_5105 = v_4991 & v_5101;
assign v_5107 = v_4989 & v_5106;
assign v_5109 = v_5008 & v_5108;
assign v_5110 = v_4988 & v_5106;
assign v_5112 = v_4986 & v_5111;
assign v_5114 = v_5014 & v_5113;
assign v_5115 = v_4985 & v_5111;
assign v_5117 = v_4983 & v_5116;
assign v_5119 = v_5020 & v_5118;
assign v_5120 = v_4982 & v_5116;
assign v_5122 = v_4980 & v_5121;
assign v_5124 = v_5026 & v_5123;
assign v_5125 = v_4979 & v_5121;
assign v_5127 = v_4977 & v_5126;
assign v_5129 = v_5032 & v_5128;
assign v_5130 = v_4976 & v_5126;
assign v_5132 = v_4974 & v_5131;
assign v_5134 = v_5038 & v_5133;
assign v_5135 = v_4973 & v_5131;
assign v_5137 = v_4971 & v_5136;
assign v_5139 = v_5044 & v_5138;
assign v_5140 = v_4970 & v_5136;
assign v_5142 = v_4968 & v_5141;
assign v_5144 = v_5050 & v_5143;
assign v_5145 = v_4967 & v_5141;
assign v_5147 = v_4965 & v_5146;
assign v_5149 = v_5056 & v_5148;
assign v_5150 = v_4964 & v_5146;
assign v_5152 = v_4962 & v_5151;
assign v_5154 = v_5062 & v_5153;
assign v_5155 = v_4961 & v_5151;
assign v_5157 = v_4959 & v_5156;
assign v_5159 = v_5068 & v_5158;
assign v_5160 = v_4958 & v_5156;
assign v_5162 = v_4956 & v_5161;
assign v_5164 = v_5074 & v_5163;
assign v_5165 = v_4955 & v_5161;
assign v_5167 = v_4953 & v_5166;
assign v_5169 = v_5080 & v_5168;
assign v_5170 = v_4952 & v_5166;
assign v_5172 = v_4950 & v_5171;
assign v_5174 = v_5086 & v_5173;
assign v_5175 = v_4949 & v_5171;
assign v_5177 = v_4947 & v_5176;
assign v_5179 = v_5092 & v_5178;
assign v_5180 = v_4946 & v_5176;
assign v_5182 = v_5181;
assign v_5184 = v_5096 & v_5183;
assign v_5185 = v_5184;
assign v_5187 = v_5186;
assign v_5189 = ~v_803;
assign v_5190 = ~v_4444;
assign v_5191 = v_4444;
assign v_5192 = ~v_807;
assign v_5193 = ~v_4448;
assign v_5194 = v_4448;
assign v_5195 = ~v_811;
assign v_5196 = ~v_4452;
assign v_5197 = v_4452;
assign v_5198 = ~v_815;
assign v_5199 = ~v_4456;
assign v_5200 = v_4456;
assign v_5201 = ~v_4459;
assign v_5202 = ~v_820;
assign v_5203 = v_820;
assign v_5204 = ~v_4463;
assign v_5205 = ~v_824;
assign v_5206 = v_824;
assign v_5207 = ~v_4467;
assign v_5208 = ~v_828;
assign v_5209 = v_828;
assign v_5210 = ~v_4471;
assign v_5211 = ~v_832;
assign v_5212 = v_832;
assign v_5213 = ~v_4475;
assign v_5214 = ~v_836;
assign v_5215 = v_836;
assign v_5216 = ~v_4479;
assign v_5217 = ~v_840;
assign v_5218 = v_840;
assign v_5219 = ~v_4483;
assign v_5220 = ~v_844;
assign v_5221 = v_844;
assign v_5222 = ~v_4487;
assign v_5223 = ~v_848;
assign v_5224 = v_848;
assign v_5225 = ~v_4491;
assign v_5226 = ~v_852;
assign v_5227 = v_852;
assign v_5228 = ~v_4495;
assign v_5229 = ~v_856;
assign v_5230 = v_856;
assign v_5231 = ~v_4499;
assign v_5232 = ~v_860;
assign v_5233 = v_860;
assign v_5234 = ~v_4503;
assign v_5235 = ~v_864;
assign v_5236 = v_864;
assign v_5237 = ~v_4507;
assign v_5238 = ~v_868;
assign v_5239 = v_5238;
assign v_5241 = v_5240;
assign v_5243 = v_5235 & v_5242;
assign v_5245 = v_4503;
assign v_5247 = v_5244 & v_5246;
assign v_5249 = v_5232 & v_5248;
assign v_5251 = v_4499;
assign v_5253 = v_5250 & v_5252;
assign v_5255 = v_5229 & v_5254;
assign v_5257 = v_4495;
assign v_5259 = v_5256 & v_5258;
assign v_5261 = v_5226 & v_5260;
assign v_5263 = v_4491;
assign v_5265 = v_5262 & v_5264;
assign v_5267 = v_5223 & v_5266;
assign v_5269 = v_4487;
assign v_5271 = v_5268 & v_5270;
assign v_5273 = v_5220 & v_5272;
assign v_5275 = v_4483;
assign v_5277 = v_5274 & v_5276;
assign v_5279 = v_5217 & v_5278;
assign v_5281 = v_4479;
assign v_5283 = v_5280 & v_5282;
assign v_5285 = v_5214 & v_5284;
assign v_5287 = v_4475;
assign v_5289 = v_5286 & v_5288;
assign v_5291 = v_5211 & v_5290;
assign v_5293 = v_4471;
assign v_5295 = v_5292 & v_5294;
assign v_5297 = v_5208 & v_5296;
assign v_5299 = v_4467;
assign v_5301 = v_5298 & v_5300;
assign v_5303 = v_5205 & v_5302;
assign v_5305 = v_4463;
assign v_5307 = v_5304 & v_5306;
assign v_5309 = v_5202 & v_5308;
assign v_5311 = v_4459;
assign v_5313 = v_5310 & v_5312;
assign v_5315 = v_5199 & v_5314;
assign v_5317 = v_815;
assign v_5319 = v_5316 & v_5318;
assign v_5321 = v_5196 & v_5320;
assign v_5323 = v_811;
assign v_5325 = v_5322 & v_5324;
assign v_5327 = v_5193 & v_5326;
assign v_5329 = v_807;
assign v_5331 = v_5328 & v_5330;
assign v_5333 = v_5190 & v_5332;
assign v_5335 = v_803;
assign v_5337 = v_5334 & v_5336;
assign v_5338 = v_5337;
assign v_5340 = v_4507;
assign v_5341 = v_868;
assign v_5342 = v_5341;
assign v_5343 = v_5340 & v_5342;
assign v_5344 = v_5343;
assign v_5345 = v_5235 & v_5344;
assign v_5347 = v_5245 & v_5346;
assign v_5348 = v_5234 & v_5344;
assign v_5350 = v_5232 & v_5349;
assign v_5352 = v_5251 & v_5351;
assign v_5353 = v_5231 & v_5349;
assign v_5355 = v_5229 & v_5354;
assign v_5357 = v_5257 & v_5356;
assign v_5358 = v_5228 & v_5354;
assign v_5360 = v_5226 & v_5359;
assign v_5362 = v_5263 & v_5361;
assign v_5363 = v_5225 & v_5359;
assign v_5365 = v_5223 & v_5364;
assign v_5367 = v_5269 & v_5366;
assign v_5368 = v_5222 & v_5364;
assign v_5370 = v_5220 & v_5369;
assign v_5372 = v_5275 & v_5371;
assign v_5373 = v_5219 & v_5369;
assign v_5375 = v_5217 & v_5374;
assign v_5377 = v_5281 & v_5376;
assign v_5378 = v_5216 & v_5374;
assign v_5380 = v_5214 & v_5379;
assign v_5382 = v_5287 & v_5381;
assign v_5383 = v_5213 & v_5379;
assign v_5385 = v_5211 & v_5384;
assign v_5387 = v_5293 & v_5386;
assign v_5388 = v_5210 & v_5384;
assign v_5390 = v_5208 & v_5389;
assign v_5392 = v_5299 & v_5391;
assign v_5393 = v_5207 & v_5389;
assign v_5395 = v_5205 & v_5394;
assign v_5397 = v_5305 & v_5396;
assign v_5398 = v_5204 & v_5394;
assign v_5400 = v_5202 & v_5399;
assign v_5402 = v_5311 & v_5401;
assign v_5403 = v_5201 & v_5399;
assign v_5405 = v_5199 & v_5404;
assign v_5407 = v_5317 & v_5406;
assign v_5408 = v_5198 & v_5404;
assign v_5410 = v_5196 & v_5409;
assign v_5412 = v_5323 & v_5411;
assign v_5413 = v_5195 & v_5409;
assign v_5415 = v_5193 & v_5414;
assign v_5417 = v_5329 & v_5416;
assign v_5418 = v_5192 & v_5414;
assign v_5420 = v_5190 & v_5419;
assign v_5422 = v_5335 & v_5421;
assign v_5423 = v_5189 & v_5419;
assign v_5425 = v_5424;
assign v_5427 = v_5339 & v_5426;
assign v_5428 = v_5427;
assign v_5430 = v_5429;
assign v_5432 = ~v_1063;
assign v_5433 = ~v_4444;
assign v_5434 = v_4444;
assign v_5435 = ~v_1067;
assign v_5436 = ~v_4448;
assign v_5437 = v_4448;
assign v_5438 = ~v_1071;
assign v_5439 = ~v_4452;
assign v_5440 = v_4452;
assign v_5441 = ~v_1075;
assign v_5442 = ~v_4456;
assign v_5443 = v_4456;
assign v_5444 = ~v_4459;
assign v_5445 = ~v_1080;
assign v_5446 = v_1080;
assign v_5447 = ~v_4463;
assign v_5448 = ~v_1084;
assign v_5449 = v_1084;
assign v_5450 = ~v_4467;
assign v_5451 = ~v_1088;
assign v_5452 = v_1088;
assign v_5453 = ~v_4471;
assign v_5454 = ~v_1092;
assign v_5455 = v_1092;
assign v_5456 = ~v_4475;
assign v_5457 = ~v_1096;
assign v_5458 = v_1096;
assign v_5459 = ~v_4479;
assign v_5460 = ~v_1100;
assign v_5461 = v_1100;
assign v_5462 = ~v_4483;
assign v_5463 = ~v_1104;
assign v_5464 = v_1104;
assign v_5465 = ~v_4487;
assign v_5466 = ~v_1108;
assign v_5467 = v_1108;
assign v_5468 = ~v_4491;
assign v_5469 = ~v_1112;
assign v_5470 = v_1112;
assign v_5471 = ~v_4495;
assign v_5472 = ~v_1116;
assign v_5473 = v_1116;
assign v_5474 = ~v_4499;
assign v_5475 = ~v_1120;
assign v_5476 = v_1120;
assign v_5477 = ~v_4503;
assign v_5478 = ~v_1124;
assign v_5479 = v_1124;
assign v_5480 = ~v_4507;
assign v_5481 = ~v_1128;
assign v_5482 = v_5481;
assign v_5484 = v_5483;
assign v_5486 = v_5478 & v_5485;
assign v_5488 = v_4503;
assign v_5490 = v_5487 & v_5489;
assign v_5492 = v_5475 & v_5491;
assign v_5494 = v_4499;
assign v_5496 = v_5493 & v_5495;
assign v_5498 = v_5472 & v_5497;
assign v_5500 = v_4495;
assign v_5502 = v_5499 & v_5501;
assign v_5504 = v_5469 & v_5503;
assign v_5506 = v_4491;
assign v_5508 = v_5505 & v_5507;
assign v_5510 = v_5466 & v_5509;
assign v_5512 = v_4487;
assign v_5514 = v_5511 & v_5513;
assign v_5516 = v_5463 & v_5515;
assign v_5518 = v_4483;
assign v_5520 = v_5517 & v_5519;
assign v_5522 = v_5460 & v_5521;
assign v_5524 = v_4479;
assign v_5526 = v_5523 & v_5525;
assign v_5528 = v_5457 & v_5527;
assign v_5530 = v_4475;
assign v_5532 = v_5529 & v_5531;
assign v_5534 = v_5454 & v_5533;
assign v_5536 = v_4471;
assign v_5538 = v_5535 & v_5537;
assign v_5540 = v_5451 & v_5539;
assign v_5542 = v_4467;
assign v_5544 = v_5541 & v_5543;
assign v_5546 = v_5448 & v_5545;
assign v_5548 = v_4463;
assign v_5550 = v_5547 & v_5549;
assign v_5552 = v_5445 & v_5551;
assign v_5554 = v_4459;
assign v_5556 = v_5553 & v_5555;
assign v_5558 = v_5442 & v_5557;
assign v_5560 = v_1075;
assign v_5562 = v_5559 & v_5561;
assign v_5564 = v_5439 & v_5563;
assign v_5566 = v_1071;
assign v_5568 = v_5565 & v_5567;
assign v_5570 = v_5436 & v_5569;
assign v_5572 = v_1067;
assign v_5574 = v_5571 & v_5573;
assign v_5576 = v_5433 & v_5575;
assign v_5578 = v_1063;
assign v_5580 = v_5577 & v_5579;
assign v_5581 = v_5580;
assign v_5583 = v_4507;
assign v_5584 = v_1128;
assign v_5585 = v_5584;
assign v_5586 = v_5583 & v_5585;
assign v_5587 = v_5586;
assign v_5588 = v_5478 & v_5587;
assign v_5590 = v_5488 & v_5589;
assign v_5591 = v_5477 & v_5587;
assign v_5593 = v_5475 & v_5592;
assign v_5595 = v_5494 & v_5594;
assign v_5596 = v_5474 & v_5592;
assign v_5598 = v_5472 & v_5597;
assign v_5600 = v_5500 & v_5599;
assign v_5601 = v_5471 & v_5597;
assign v_5603 = v_5469 & v_5602;
assign v_5605 = v_5506 & v_5604;
assign v_5606 = v_5468 & v_5602;
assign v_5608 = v_5466 & v_5607;
assign v_5610 = v_5512 & v_5609;
assign v_5611 = v_5465 & v_5607;
assign v_5613 = v_5463 & v_5612;
assign v_5615 = v_5518 & v_5614;
assign v_5616 = v_5462 & v_5612;
assign v_5618 = v_5460 & v_5617;
assign v_5620 = v_5524 & v_5619;
assign v_5621 = v_5459 & v_5617;
assign v_5623 = v_5457 & v_5622;
assign v_5625 = v_5530 & v_5624;
assign v_5626 = v_5456 & v_5622;
assign v_5628 = v_5454 & v_5627;
assign v_5630 = v_5536 & v_5629;
assign v_5631 = v_5453 & v_5627;
assign v_5633 = v_5451 & v_5632;
assign v_5635 = v_5542 & v_5634;
assign v_5636 = v_5450 & v_5632;
assign v_5638 = v_5448 & v_5637;
assign v_5640 = v_5548 & v_5639;
assign v_5641 = v_5447 & v_5637;
assign v_5643 = v_5445 & v_5642;
assign v_5645 = v_5554 & v_5644;
assign v_5646 = v_5444 & v_5642;
assign v_5648 = v_5442 & v_5647;
assign v_5650 = v_5560 & v_5649;
assign v_5651 = v_5441 & v_5647;
assign v_5653 = v_5439 & v_5652;
assign v_5655 = v_5566 & v_5654;
assign v_5656 = v_5438 & v_5652;
assign v_5658 = v_5436 & v_5657;
assign v_5660 = v_5572 & v_5659;
assign v_5661 = v_5435 & v_5657;
assign v_5663 = v_5433 & v_5662;
assign v_5665 = v_5578 & v_5664;
assign v_5666 = v_5432 & v_5662;
assign v_5668 = v_5667;
assign v_5670 = v_5582 & v_5669;
assign v_5671 = v_5670;
assign v_5673 = v_5672;
assign v_5675 = ~v_1323;
assign v_5676 = ~v_4444;
assign v_5677 = v_4444;
assign v_5678 = ~v_1327;
assign v_5679 = ~v_4448;
assign v_5680 = v_4448;
assign v_5681 = ~v_1331;
assign v_5682 = ~v_4452;
assign v_5683 = v_4452;
assign v_5684 = ~v_1335;
assign v_5685 = ~v_4456;
assign v_5686 = v_4456;
assign v_5687 = ~v_4459;
assign v_5688 = ~v_1340;
assign v_5689 = v_1340;
assign v_5690 = ~v_4463;
assign v_5691 = ~v_1344;
assign v_5692 = v_1344;
assign v_5693 = ~v_4467;
assign v_5694 = ~v_1348;
assign v_5695 = v_1348;
assign v_5696 = ~v_4471;
assign v_5697 = ~v_1352;
assign v_5698 = v_1352;
assign v_5699 = ~v_4475;
assign v_5700 = ~v_1356;
assign v_5701 = v_1356;
assign v_5702 = ~v_4479;
assign v_5703 = ~v_1360;
assign v_5704 = v_1360;
assign v_5705 = ~v_4483;
assign v_5706 = ~v_1364;
assign v_5707 = v_1364;
assign v_5708 = ~v_4487;
assign v_5709 = ~v_1368;
assign v_5710 = v_1368;
assign v_5711 = ~v_4491;
assign v_5712 = ~v_1372;
assign v_5713 = v_1372;
assign v_5714 = ~v_4495;
assign v_5715 = ~v_1376;
assign v_5716 = v_1376;
assign v_5717 = ~v_4499;
assign v_5718 = ~v_1380;
assign v_5719 = v_1380;
assign v_5720 = ~v_4503;
assign v_5721 = ~v_1384;
assign v_5722 = v_1384;
assign v_5723 = ~v_4507;
assign v_5724 = ~v_1388;
assign v_5725 = v_5724;
assign v_5727 = v_5726;
assign v_5729 = v_5721 & v_5728;
assign v_5731 = v_4503;
assign v_5733 = v_5730 & v_5732;
assign v_5735 = v_5718 & v_5734;
assign v_5737 = v_4499;
assign v_5739 = v_5736 & v_5738;
assign v_5741 = v_5715 & v_5740;
assign v_5743 = v_4495;
assign v_5745 = v_5742 & v_5744;
assign v_5747 = v_5712 & v_5746;
assign v_5749 = v_4491;
assign v_5751 = v_5748 & v_5750;
assign v_5753 = v_5709 & v_5752;
assign v_5755 = v_4487;
assign v_5757 = v_5754 & v_5756;
assign v_5759 = v_5706 & v_5758;
assign v_5761 = v_4483;
assign v_5763 = v_5760 & v_5762;
assign v_5765 = v_5703 & v_5764;
assign v_5767 = v_4479;
assign v_5769 = v_5766 & v_5768;
assign v_5771 = v_5700 & v_5770;
assign v_5773 = v_4475;
assign v_5775 = v_5772 & v_5774;
assign v_5777 = v_5697 & v_5776;
assign v_5779 = v_4471;
assign v_5781 = v_5778 & v_5780;
assign v_5783 = v_5694 & v_5782;
assign v_5785 = v_4467;
assign v_5787 = v_5784 & v_5786;
assign v_5789 = v_5691 & v_5788;
assign v_5791 = v_4463;
assign v_5793 = v_5790 & v_5792;
assign v_5795 = v_5688 & v_5794;
assign v_5797 = v_4459;
assign v_5799 = v_5796 & v_5798;
assign v_5801 = v_5685 & v_5800;
assign v_5803 = v_1335;
assign v_5805 = v_5802 & v_5804;
assign v_5807 = v_5682 & v_5806;
assign v_5809 = v_1331;
assign v_5811 = v_5808 & v_5810;
assign v_5813 = v_5679 & v_5812;
assign v_5815 = v_1327;
assign v_5817 = v_5814 & v_5816;
assign v_5819 = v_5676 & v_5818;
assign v_5821 = v_1323;
assign v_5823 = v_5820 & v_5822;
assign v_5824 = v_5823;
assign v_5826 = v_4507;
assign v_5827 = v_1388;
assign v_5828 = v_5827;
assign v_5829 = v_5826 & v_5828;
assign v_5830 = v_5829;
assign v_5831 = v_5721 & v_5830;
assign v_5833 = v_5731 & v_5832;
assign v_5834 = v_5720 & v_5830;
assign v_5836 = v_5718 & v_5835;
assign v_5838 = v_5737 & v_5837;
assign v_5839 = v_5717 & v_5835;
assign v_5841 = v_5715 & v_5840;
assign v_5843 = v_5743 & v_5842;
assign v_5844 = v_5714 & v_5840;
assign v_5846 = v_5712 & v_5845;
assign v_5848 = v_5749 & v_5847;
assign v_5849 = v_5711 & v_5845;
assign v_5851 = v_5709 & v_5850;
assign v_5853 = v_5755 & v_5852;
assign v_5854 = v_5708 & v_5850;
assign v_5856 = v_5706 & v_5855;
assign v_5858 = v_5761 & v_5857;
assign v_5859 = v_5705 & v_5855;
assign v_5861 = v_5703 & v_5860;
assign v_5863 = v_5767 & v_5862;
assign v_5864 = v_5702 & v_5860;
assign v_5866 = v_5700 & v_5865;
assign v_5868 = v_5773 & v_5867;
assign v_5869 = v_5699 & v_5865;
assign v_5871 = v_5697 & v_5870;
assign v_5873 = v_5779 & v_5872;
assign v_5874 = v_5696 & v_5870;
assign v_5876 = v_5694 & v_5875;
assign v_5878 = v_5785 & v_5877;
assign v_5879 = v_5693 & v_5875;
assign v_5881 = v_5691 & v_5880;
assign v_5883 = v_5791 & v_5882;
assign v_5884 = v_5690 & v_5880;
assign v_5886 = v_5688 & v_5885;
assign v_5888 = v_5797 & v_5887;
assign v_5889 = v_5687 & v_5885;
assign v_5891 = v_5685 & v_5890;
assign v_5893 = v_5803 & v_5892;
assign v_5894 = v_5684 & v_5890;
assign v_5896 = v_5682 & v_5895;
assign v_5898 = v_5809 & v_5897;
assign v_5899 = v_5681 & v_5895;
assign v_5901 = v_5679 & v_5900;
assign v_5903 = v_5815 & v_5902;
assign v_5904 = v_5678 & v_5900;
assign v_5906 = v_5676 & v_5905;
assign v_5908 = v_5821 & v_5907;
assign v_5909 = v_5675 & v_5905;
assign v_5911 = v_5910;
assign v_5913 = v_5825 & v_5912;
assign v_5914 = v_5913;
assign v_5916 = v_5915;
assign v_5918 = ~v_1583;
assign v_5919 = ~v_4444;
assign v_5920 = v_4444;
assign v_5921 = ~v_1587;
assign v_5922 = ~v_4448;
assign v_5923 = v_4448;
assign v_5924 = ~v_1591;
assign v_5925 = ~v_4452;
assign v_5926 = v_4452;
assign v_5927 = ~v_1595;
assign v_5928 = ~v_4456;
assign v_5929 = v_4456;
assign v_5930 = ~v_4459;
assign v_5931 = ~v_1600;
assign v_5932 = v_1600;
assign v_5933 = ~v_4463;
assign v_5934 = ~v_1604;
assign v_5935 = v_1604;
assign v_5936 = ~v_4467;
assign v_5937 = ~v_1608;
assign v_5938 = v_1608;
assign v_5939 = ~v_4471;
assign v_5940 = ~v_1612;
assign v_5941 = v_1612;
assign v_5942 = ~v_4475;
assign v_5943 = ~v_1616;
assign v_5944 = v_1616;
assign v_5945 = ~v_4479;
assign v_5946 = ~v_1620;
assign v_5947 = v_1620;
assign v_5948 = ~v_4483;
assign v_5949 = ~v_1624;
assign v_5950 = v_1624;
assign v_5951 = ~v_4487;
assign v_5952 = ~v_1628;
assign v_5953 = v_1628;
assign v_5954 = ~v_4491;
assign v_5955 = ~v_1632;
assign v_5956 = v_1632;
assign v_5957 = ~v_4495;
assign v_5958 = ~v_1636;
assign v_5959 = v_1636;
assign v_5960 = ~v_4499;
assign v_5961 = ~v_1640;
assign v_5962 = v_1640;
assign v_5963 = ~v_4503;
assign v_5964 = ~v_1644;
assign v_5965 = v_1644;
assign v_5966 = ~v_4507;
assign v_5967 = ~v_1648;
assign v_5968 = v_5967;
assign v_5970 = v_5969;
assign v_5972 = v_5964 & v_5971;
assign v_5974 = v_4503;
assign v_5976 = v_5973 & v_5975;
assign v_5978 = v_5961 & v_5977;
assign v_5980 = v_4499;
assign v_5982 = v_5979 & v_5981;
assign v_5984 = v_5958 & v_5983;
assign v_5986 = v_4495;
assign v_5988 = v_5985 & v_5987;
assign v_5990 = v_5955 & v_5989;
assign v_5992 = v_4491;
assign v_5994 = v_5991 & v_5993;
assign v_5996 = v_5952 & v_5995;
assign v_5998 = v_4487;
assign v_6000 = v_5997 & v_5999;
assign v_6002 = v_5949 & v_6001;
assign v_6004 = v_4483;
assign v_6006 = v_6003 & v_6005;
assign v_6008 = v_5946 & v_6007;
assign v_6010 = v_4479;
assign v_6012 = v_6009 & v_6011;
assign v_6014 = v_5943 & v_6013;
assign v_6016 = v_4475;
assign v_6018 = v_6015 & v_6017;
assign v_6020 = v_5940 & v_6019;
assign v_6022 = v_4471;
assign v_6024 = v_6021 & v_6023;
assign v_6026 = v_5937 & v_6025;
assign v_6028 = v_4467;
assign v_6030 = v_6027 & v_6029;
assign v_6032 = v_5934 & v_6031;
assign v_6034 = v_4463;
assign v_6036 = v_6033 & v_6035;
assign v_6038 = v_5931 & v_6037;
assign v_6040 = v_4459;
assign v_6042 = v_6039 & v_6041;
assign v_6044 = v_5928 & v_6043;
assign v_6046 = v_1595;
assign v_6048 = v_6045 & v_6047;
assign v_6050 = v_5925 & v_6049;
assign v_6052 = v_1591;
assign v_6054 = v_6051 & v_6053;
assign v_6056 = v_5922 & v_6055;
assign v_6058 = v_1587;
assign v_6060 = v_6057 & v_6059;
assign v_6062 = v_5919 & v_6061;
assign v_6064 = v_1583;
assign v_6066 = v_6063 & v_6065;
assign v_6067 = v_6066;
assign v_6069 = v_4507;
assign v_6070 = v_1648;
assign v_6071 = v_6070;
assign v_6072 = v_6069 & v_6071;
assign v_6073 = v_6072;
assign v_6074 = v_5964 & v_6073;
assign v_6076 = v_5974 & v_6075;
assign v_6077 = v_5963 & v_6073;
assign v_6079 = v_5961 & v_6078;
assign v_6081 = v_5980 & v_6080;
assign v_6082 = v_5960 & v_6078;
assign v_6084 = v_5958 & v_6083;
assign v_6086 = v_5986 & v_6085;
assign v_6087 = v_5957 & v_6083;
assign v_6089 = v_5955 & v_6088;
assign v_6091 = v_5992 & v_6090;
assign v_6092 = v_5954 & v_6088;
assign v_6094 = v_5952 & v_6093;
assign v_6096 = v_5998 & v_6095;
assign v_6097 = v_5951 & v_6093;
assign v_6099 = v_5949 & v_6098;
assign v_6101 = v_6004 & v_6100;
assign v_6102 = v_5948 & v_6098;
assign v_6104 = v_5946 & v_6103;
assign v_6106 = v_6010 & v_6105;
assign v_6107 = v_5945 & v_6103;
assign v_6109 = v_5943 & v_6108;
assign v_6111 = v_6016 & v_6110;
assign v_6112 = v_5942 & v_6108;
assign v_6114 = v_5940 & v_6113;
assign v_6116 = v_6022 & v_6115;
assign v_6117 = v_5939 & v_6113;
assign v_6119 = v_5937 & v_6118;
assign v_6121 = v_6028 & v_6120;
assign v_6122 = v_5936 & v_6118;
assign v_6124 = v_5934 & v_6123;
assign v_6126 = v_6034 & v_6125;
assign v_6127 = v_5933 & v_6123;
assign v_6129 = v_5931 & v_6128;
assign v_6131 = v_6040 & v_6130;
assign v_6132 = v_5930 & v_6128;
assign v_6134 = v_5928 & v_6133;
assign v_6136 = v_6046 & v_6135;
assign v_6137 = v_5927 & v_6133;
assign v_6139 = v_5925 & v_6138;
assign v_6141 = v_6052 & v_6140;
assign v_6142 = v_5924 & v_6138;
assign v_6144 = v_5922 & v_6143;
assign v_6146 = v_6058 & v_6145;
assign v_6147 = v_5921 & v_6143;
assign v_6149 = v_5919 & v_6148;
assign v_6151 = v_6064 & v_6150;
assign v_6152 = v_5918 & v_6148;
assign v_6154 = v_6153;
assign v_6156 = v_6068 & v_6155;
assign v_6157 = v_6156;
assign v_6159 = v_6158;
assign v_6161 = ~v_1843;
assign v_6162 = ~v_4444;
assign v_6163 = v_4444;
assign v_6164 = ~v_1847;
assign v_6165 = ~v_4448;
assign v_6166 = v_4448;
assign v_6167 = ~v_1851;
assign v_6168 = ~v_4452;
assign v_6169 = v_4452;
assign v_6170 = ~v_1855;
assign v_6171 = ~v_4456;
assign v_6172 = v_4456;
assign v_6173 = ~v_4459;
assign v_6174 = ~v_1860;
assign v_6175 = v_1860;
assign v_6176 = ~v_4463;
assign v_6177 = ~v_1864;
assign v_6178 = v_1864;
assign v_6179 = ~v_4467;
assign v_6180 = ~v_1868;
assign v_6181 = v_1868;
assign v_6182 = ~v_4471;
assign v_6183 = ~v_1872;
assign v_6184 = v_1872;
assign v_6185 = ~v_4475;
assign v_6186 = ~v_1876;
assign v_6187 = v_1876;
assign v_6188 = ~v_4479;
assign v_6189 = ~v_1880;
assign v_6190 = v_1880;
assign v_6191 = ~v_4483;
assign v_6192 = ~v_1884;
assign v_6193 = v_1884;
assign v_6194 = ~v_4487;
assign v_6195 = ~v_1888;
assign v_6196 = v_1888;
assign v_6197 = ~v_4491;
assign v_6198 = ~v_1892;
assign v_6199 = v_1892;
assign v_6200 = ~v_4495;
assign v_6201 = ~v_1896;
assign v_6202 = v_1896;
assign v_6203 = ~v_4499;
assign v_6204 = ~v_1900;
assign v_6205 = v_1900;
assign v_6206 = ~v_4503;
assign v_6207 = ~v_1904;
assign v_6208 = v_1904;
assign v_6209 = ~v_4507;
assign v_6210 = ~v_1908;
assign v_6211 = v_6210;
assign v_6213 = v_6212;
assign v_6215 = v_6207 & v_6214;
assign v_6217 = v_4503;
assign v_6219 = v_6216 & v_6218;
assign v_6221 = v_6204 & v_6220;
assign v_6223 = v_4499;
assign v_6225 = v_6222 & v_6224;
assign v_6227 = v_6201 & v_6226;
assign v_6229 = v_4495;
assign v_6231 = v_6228 & v_6230;
assign v_6233 = v_6198 & v_6232;
assign v_6235 = v_4491;
assign v_6237 = v_6234 & v_6236;
assign v_6239 = v_6195 & v_6238;
assign v_6241 = v_4487;
assign v_6243 = v_6240 & v_6242;
assign v_6245 = v_6192 & v_6244;
assign v_6247 = v_4483;
assign v_6249 = v_6246 & v_6248;
assign v_6251 = v_6189 & v_6250;
assign v_6253 = v_4479;
assign v_6255 = v_6252 & v_6254;
assign v_6257 = v_6186 & v_6256;
assign v_6259 = v_4475;
assign v_6261 = v_6258 & v_6260;
assign v_6263 = v_6183 & v_6262;
assign v_6265 = v_4471;
assign v_6267 = v_6264 & v_6266;
assign v_6269 = v_6180 & v_6268;
assign v_6271 = v_4467;
assign v_6273 = v_6270 & v_6272;
assign v_6275 = v_6177 & v_6274;
assign v_6277 = v_4463;
assign v_6279 = v_6276 & v_6278;
assign v_6281 = v_6174 & v_6280;
assign v_6283 = v_4459;
assign v_6285 = v_6282 & v_6284;
assign v_6287 = v_6171 & v_6286;
assign v_6289 = v_1855;
assign v_6291 = v_6288 & v_6290;
assign v_6293 = v_6168 & v_6292;
assign v_6295 = v_1851;
assign v_6297 = v_6294 & v_6296;
assign v_6299 = v_6165 & v_6298;
assign v_6301 = v_1847;
assign v_6303 = v_6300 & v_6302;
assign v_6305 = v_6162 & v_6304;
assign v_6307 = v_1843;
assign v_6309 = v_6306 & v_6308;
assign v_6310 = v_6309;
assign v_6312 = v_4507;
assign v_6313 = v_1908;
assign v_6314 = v_6313;
assign v_6315 = v_6312 & v_6314;
assign v_6316 = v_6315;
assign v_6317 = v_6207 & v_6316;
assign v_6319 = v_6217 & v_6318;
assign v_6320 = v_6206 & v_6316;
assign v_6322 = v_6204 & v_6321;
assign v_6324 = v_6223 & v_6323;
assign v_6325 = v_6203 & v_6321;
assign v_6327 = v_6201 & v_6326;
assign v_6329 = v_6229 & v_6328;
assign v_6330 = v_6200 & v_6326;
assign v_6332 = v_6198 & v_6331;
assign v_6334 = v_6235 & v_6333;
assign v_6335 = v_6197 & v_6331;
assign v_6337 = v_6195 & v_6336;
assign v_6339 = v_6241 & v_6338;
assign v_6340 = v_6194 & v_6336;
assign v_6342 = v_6192 & v_6341;
assign v_6344 = v_6247 & v_6343;
assign v_6345 = v_6191 & v_6341;
assign v_6347 = v_6189 & v_6346;
assign v_6349 = v_6253 & v_6348;
assign v_6350 = v_6188 & v_6346;
assign v_6352 = v_6186 & v_6351;
assign v_6354 = v_6259 & v_6353;
assign v_6355 = v_6185 & v_6351;
assign v_6357 = v_6183 & v_6356;
assign v_6359 = v_6265 & v_6358;
assign v_6360 = v_6182 & v_6356;
assign v_6362 = v_6180 & v_6361;
assign v_6364 = v_6271 & v_6363;
assign v_6365 = v_6179 & v_6361;
assign v_6367 = v_6177 & v_6366;
assign v_6369 = v_6277 & v_6368;
assign v_6370 = v_6176 & v_6366;
assign v_6372 = v_6174 & v_6371;
assign v_6374 = v_6283 & v_6373;
assign v_6375 = v_6173 & v_6371;
assign v_6377 = v_6171 & v_6376;
assign v_6379 = v_6289 & v_6378;
assign v_6380 = v_6170 & v_6376;
assign v_6382 = v_6168 & v_6381;
assign v_6384 = v_6295 & v_6383;
assign v_6385 = v_6167 & v_6381;
assign v_6387 = v_6165 & v_6386;
assign v_6389 = v_6301 & v_6388;
assign v_6390 = v_6164 & v_6386;
assign v_6392 = v_6162 & v_6391;
assign v_6394 = v_6307 & v_6393;
assign v_6395 = v_6161 & v_6391;
assign v_6397 = v_6396;
assign v_6399 = v_6311 & v_6398;
assign v_6400 = v_6399;
assign v_6402 = v_6401;
assign v_6404 = ~v_2103;
assign v_6405 = ~v_4444;
assign v_6406 = v_4444;
assign v_6407 = ~v_2107;
assign v_6408 = ~v_4448;
assign v_6409 = v_4448;
assign v_6410 = ~v_2111;
assign v_6411 = ~v_4452;
assign v_6412 = v_4452;
assign v_6413 = ~v_2115;
assign v_6414 = ~v_4456;
assign v_6415 = v_4456;
assign v_6416 = ~v_4459;
assign v_6417 = ~v_2120;
assign v_6418 = v_2120;
assign v_6419 = ~v_4463;
assign v_6420 = ~v_2124;
assign v_6421 = v_2124;
assign v_6422 = ~v_4467;
assign v_6423 = ~v_2128;
assign v_6424 = v_2128;
assign v_6425 = ~v_4471;
assign v_6426 = ~v_2132;
assign v_6427 = v_2132;
assign v_6428 = ~v_4475;
assign v_6429 = ~v_2136;
assign v_6430 = v_2136;
assign v_6431 = ~v_4479;
assign v_6432 = ~v_2140;
assign v_6433 = v_2140;
assign v_6434 = ~v_4483;
assign v_6435 = ~v_2144;
assign v_6436 = v_2144;
assign v_6437 = ~v_4487;
assign v_6438 = ~v_2148;
assign v_6439 = v_2148;
assign v_6440 = ~v_4491;
assign v_6441 = ~v_2152;
assign v_6442 = v_2152;
assign v_6443 = ~v_4495;
assign v_6444 = ~v_2156;
assign v_6445 = v_2156;
assign v_6446 = ~v_4499;
assign v_6447 = ~v_2160;
assign v_6448 = v_2160;
assign v_6449 = ~v_4503;
assign v_6450 = ~v_2164;
assign v_6451 = v_2164;
assign v_6452 = ~v_4507;
assign v_6453 = ~v_2168;
assign v_6454 = v_6453;
assign v_6456 = v_6455;
assign v_6458 = v_6450 & v_6457;
assign v_6460 = v_4503;
assign v_6462 = v_6459 & v_6461;
assign v_6464 = v_6447 & v_6463;
assign v_6466 = v_4499;
assign v_6468 = v_6465 & v_6467;
assign v_6470 = v_6444 & v_6469;
assign v_6472 = v_4495;
assign v_6474 = v_6471 & v_6473;
assign v_6476 = v_6441 & v_6475;
assign v_6478 = v_4491;
assign v_6480 = v_6477 & v_6479;
assign v_6482 = v_6438 & v_6481;
assign v_6484 = v_4487;
assign v_6486 = v_6483 & v_6485;
assign v_6488 = v_6435 & v_6487;
assign v_6490 = v_4483;
assign v_6492 = v_6489 & v_6491;
assign v_6494 = v_6432 & v_6493;
assign v_6496 = v_4479;
assign v_6498 = v_6495 & v_6497;
assign v_6500 = v_6429 & v_6499;
assign v_6502 = v_4475;
assign v_6504 = v_6501 & v_6503;
assign v_6506 = v_6426 & v_6505;
assign v_6508 = v_4471;
assign v_6510 = v_6507 & v_6509;
assign v_6512 = v_6423 & v_6511;
assign v_6514 = v_4467;
assign v_6516 = v_6513 & v_6515;
assign v_6518 = v_6420 & v_6517;
assign v_6520 = v_4463;
assign v_6522 = v_6519 & v_6521;
assign v_6524 = v_6417 & v_6523;
assign v_6526 = v_4459;
assign v_6528 = v_6525 & v_6527;
assign v_6530 = v_6414 & v_6529;
assign v_6532 = v_2115;
assign v_6534 = v_6531 & v_6533;
assign v_6536 = v_6411 & v_6535;
assign v_6538 = v_2111;
assign v_6540 = v_6537 & v_6539;
assign v_6542 = v_6408 & v_6541;
assign v_6544 = v_2107;
assign v_6546 = v_6543 & v_6545;
assign v_6548 = v_6405 & v_6547;
assign v_6550 = v_2103;
assign v_6552 = v_6549 & v_6551;
assign v_6553 = v_6552;
assign v_6555 = v_4507;
assign v_6556 = v_2168;
assign v_6557 = v_6556;
assign v_6558 = v_6555 & v_6557;
assign v_6559 = v_6558;
assign v_6560 = v_6450 & v_6559;
assign v_6562 = v_6460 & v_6561;
assign v_6563 = v_6449 & v_6559;
assign v_6565 = v_6447 & v_6564;
assign v_6567 = v_6466 & v_6566;
assign v_6568 = v_6446 & v_6564;
assign v_6570 = v_6444 & v_6569;
assign v_6572 = v_6472 & v_6571;
assign v_6573 = v_6443 & v_6569;
assign v_6575 = v_6441 & v_6574;
assign v_6577 = v_6478 & v_6576;
assign v_6578 = v_6440 & v_6574;
assign v_6580 = v_6438 & v_6579;
assign v_6582 = v_6484 & v_6581;
assign v_6583 = v_6437 & v_6579;
assign v_6585 = v_6435 & v_6584;
assign v_6587 = v_6490 & v_6586;
assign v_6588 = v_6434 & v_6584;
assign v_6590 = v_6432 & v_6589;
assign v_6592 = v_6496 & v_6591;
assign v_6593 = v_6431 & v_6589;
assign v_6595 = v_6429 & v_6594;
assign v_6597 = v_6502 & v_6596;
assign v_6598 = v_6428 & v_6594;
assign v_6600 = v_6426 & v_6599;
assign v_6602 = v_6508 & v_6601;
assign v_6603 = v_6425 & v_6599;
assign v_6605 = v_6423 & v_6604;
assign v_6607 = v_6514 & v_6606;
assign v_6608 = v_6422 & v_6604;
assign v_6610 = v_6420 & v_6609;
assign v_6612 = v_6520 & v_6611;
assign v_6613 = v_6419 & v_6609;
assign v_6615 = v_6417 & v_6614;
assign v_6617 = v_6526 & v_6616;
assign v_6618 = v_6416 & v_6614;
assign v_6620 = v_6414 & v_6619;
assign v_6622 = v_6532 & v_6621;
assign v_6623 = v_6413 & v_6619;
assign v_6625 = v_6411 & v_6624;
assign v_6627 = v_6538 & v_6626;
assign v_6628 = v_6410 & v_6624;
assign v_6630 = v_6408 & v_6629;
assign v_6632 = v_6544 & v_6631;
assign v_6633 = v_6407 & v_6629;
assign v_6635 = v_6405 & v_6634;
assign v_6637 = v_6550 & v_6636;
assign v_6638 = v_6404 & v_6634;
assign v_6640 = v_6639;
assign v_6642 = v_6554 & v_6641;
assign v_6643 = v_6642;
assign v_6645 = v_6644;
assign v_6647 = ~v_2363;
assign v_6648 = ~v_4444;
assign v_6649 = v_4444;
assign v_6650 = ~v_2367;
assign v_6651 = ~v_4448;
assign v_6652 = v_4448;
assign v_6653 = ~v_2371;
assign v_6654 = ~v_4452;
assign v_6655 = v_4452;
assign v_6656 = ~v_2375;
assign v_6657 = ~v_4456;
assign v_6658 = v_4456;
assign v_6659 = ~v_4459;
assign v_6660 = ~v_2380;
assign v_6661 = v_2380;
assign v_6662 = ~v_4463;
assign v_6663 = ~v_2384;
assign v_6664 = v_2384;
assign v_6665 = ~v_4467;
assign v_6666 = ~v_2388;
assign v_6667 = v_2388;
assign v_6668 = ~v_4471;
assign v_6669 = ~v_2392;
assign v_6670 = v_2392;
assign v_6671 = ~v_4475;
assign v_6672 = ~v_2396;
assign v_6673 = v_2396;
assign v_6674 = ~v_4479;
assign v_6675 = ~v_2400;
assign v_6676 = v_2400;
assign v_6677 = ~v_4483;
assign v_6678 = ~v_2404;
assign v_6679 = v_2404;
assign v_6680 = ~v_4487;
assign v_6681 = ~v_2408;
assign v_6682 = v_2408;
assign v_6683 = ~v_4491;
assign v_6684 = ~v_2412;
assign v_6685 = v_2412;
assign v_6686 = ~v_4495;
assign v_6687 = ~v_2416;
assign v_6688 = v_2416;
assign v_6689 = ~v_4499;
assign v_6690 = ~v_2420;
assign v_6691 = v_2420;
assign v_6692 = ~v_4503;
assign v_6693 = ~v_2424;
assign v_6694 = v_2424;
assign v_6695 = ~v_4507;
assign v_6696 = ~v_2428;
assign v_6697 = v_6696;
assign v_6699 = v_6698;
assign v_6701 = v_6693 & v_6700;
assign v_6703 = v_4503;
assign v_6705 = v_6702 & v_6704;
assign v_6707 = v_6690 & v_6706;
assign v_6709 = v_4499;
assign v_6711 = v_6708 & v_6710;
assign v_6713 = v_6687 & v_6712;
assign v_6715 = v_4495;
assign v_6717 = v_6714 & v_6716;
assign v_6719 = v_6684 & v_6718;
assign v_6721 = v_4491;
assign v_6723 = v_6720 & v_6722;
assign v_6725 = v_6681 & v_6724;
assign v_6727 = v_4487;
assign v_6729 = v_6726 & v_6728;
assign v_6731 = v_6678 & v_6730;
assign v_6733 = v_4483;
assign v_6735 = v_6732 & v_6734;
assign v_6737 = v_6675 & v_6736;
assign v_6739 = v_4479;
assign v_6741 = v_6738 & v_6740;
assign v_6743 = v_6672 & v_6742;
assign v_6745 = v_4475;
assign v_6747 = v_6744 & v_6746;
assign v_6749 = v_6669 & v_6748;
assign v_6751 = v_4471;
assign v_6753 = v_6750 & v_6752;
assign v_6755 = v_6666 & v_6754;
assign v_6757 = v_4467;
assign v_6759 = v_6756 & v_6758;
assign v_6761 = v_6663 & v_6760;
assign v_6763 = v_4463;
assign v_6765 = v_6762 & v_6764;
assign v_6767 = v_6660 & v_6766;
assign v_6769 = v_4459;
assign v_6771 = v_6768 & v_6770;
assign v_6773 = v_6657 & v_6772;
assign v_6775 = v_2375;
assign v_6777 = v_6774 & v_6776;
assign v_6779 = v_6654 & v_6778;
assign v_6781 = v_2371;
assign v_6783 = v_6780 & v_6782;
assign v_6785 = v_6651 & v_6784;
assign v_6787 = v_2367;
assign v_6789 = v_6786 & v_6788;
assign v_6791 = v_6648 & v_6790;
assign v_6793 = v_2363;
assign v_6795 = v_6792 & v_6794;
assign v_6796 = v_6795;
assign v_6798 = v_4507;
assign v_6799 = v_2428;
assign v_6800 = v_6799;
assign v_6801 = v_6798 & v_6800;
assign v_6802 = v_6801;
assign v_6803 = v_6693 & v_6802;
assign v_6805 = v_6703 & v_6804;
assign v_6806 = v_6692 & v_6802;
assign v_6808 = v_6690 & v_6807;
assign v_6810 = v_6709 & v_6809;
assign v_6811 = v_6689 & v_6807;
assign v_6813 = v_6687 & v_6812;
assign v_6815 = v_6715 & v_6814;
assign v_6816 = v_6686 & v_6812;
assign v_6818 = v_6684 & v_6817;
assign v_6820 = v_6721 & v_6819;
assign v_6821 = v_6683 & v_6817;
assign v_6823 = v_6681 & v_6822;
assign v_6825 = v_6727 & v_6824;
assign v_6826 = v_6680 & v_6822;
assign v_6828 = v_6678 & v_6827;
assign v_6830 = v_6733 & v_6829;
assign v_6831 = v_6677 & v_6827;
assign v_6833 = v_6675 & v_6832;
assign v_6835 = v_6739 & v_6834;
assign v_6836 = v_6674 & v_6832;
assign v_6838 = v_6672 & v_6837;
assign v_6840 = v_6745 & v_6839;
assign v_6841 = v_6671 & v_6837;
assign v_6843 = v_6669 & v_6842;
assign v_6845 = v_6751 & v_6844;
assign v_6846 = v_6668 & v_6842;
assign v_6848 = v_6666 & v_6847;
assign v_6850 = v_6757 & v_6849;
assign v_6851 = v_6665 & v_6847;
assign v_6853 = v_6663 & v_6852;
assign v_6855 = v_6763 & v_6854;
assign v_6856 = v_6662 & v_6852;
assign v_6858 = v_6660 & v_6857;
assign v_6860 = v_6769 & v_6859;
assign v_6861 = v_6659 & v_6857;
assign v_6863 = v_6657 & v_6862;
assign v_6865 = v_6775 & v_6864;
assign v_6866 = v_6656 & v_6862;
assign v_6868 = v_6654 & v_6867;
assign v_6870 = v_6781 & v_6869;
assign v_6871 = v_6653 & v_6867;
assign v_6873 = v_6651 & v_6872;
assign v_6875 = v_6787 & v_6874;
assign v_6876 = v_6650 & v_6872;
assign v_6878 = v_6648 & v_6877;
assign v_6880 = v_6793 & v_6879;
assign v_6881 = v_6647 & v_6877;
assign v_6883 = v_6882;
assign v_6885 = v_6797 & v_6884;
assign v_6886 = v_6885;
assign v_6888 = v_6887;
assign v_6890 = ~v_2623;
assign v_6891 = ~v_4444;
assign v_6892 = v_4444;
assign v_6893 = ~v_2627;
assign v_6894 = ~v_4448;
assign v_6895 = v_4448;
assign v_6896 = ~v_2631;
assign v_6897 = ~v_4452;
assign v_6898 = v_4452;
assign v_6899 = ~v_2635;
assign v_6900 = ~v_4456;
assign v_6901 = v_4456;
assign v_6902 = ~v_4459;
assign v_6903 = ~v_2640;
assign v_6904 = v_2640;
assign v_6905 = ~v_4463;
assign v_6906 = ~v_2644;
assign v_6907 = v_2644;
assign v_6908 = ~v_4467;
assign v_6909 = ~v_2648;
assign v_6910 = v_2648;
assign v_6911 = ~v_4471;
assign v_6912 = ~v_2652;
assign v_6913 = v_2652;
assign v_6914 = ~v_4475;
assign v_6915 = ~v_2656;
assign v_6916 = v_2656;
assign v_6917 = ~v_4479;
assign v_6918 = ~v_2660;
assign v_6919 = v_2660;
assign v_6920 = ~v_4483;
assign v_6921 = ~v_2664;
assign v_6922 = v_2664;
assign v_6923 = ~v_4487;
assign v_6924 = ~v_2668;
assign v_6925 = v_2668;
assign v_6926 = ~v_4491;
assign v_6927 = ~v_2672;
assign v_6928 = v_2672;
assign v_6929 = ~v_4495;
assign v_6930 = ~v_2676;
assign v_6931 = v_2676;
assign v_6932 = ~v_4499;
assign v_6933 = ~v_2680;
assign v_6934 = v_2680;
assign v_6935 = ~v_4503;
assign v_6936 = ~v_2684;
assign v_6937 = v_2684;
assign v_6938 = ~v_4507;
assign v_6939 = ~v_2688;
assign v_6940 = v_6939;
assign v_6942 = v_6941;
assign v_6944 = v_6936 & v_6943;
assign v_6946 = v_4503;
assign v_6948 = v_6945 & v_6947;
assign v_6950 = v_6933 & v_6949;
assign v_6952 = v_4499;
assign v_6954 = v_6951 & v_6953;
assign v_6956 = v_6930 & v_6955;
assign v_6958 = v_4495;
assign v_6960 = v_6957 & v_6959;
assign v_6962 = v_6927 & v_6961;
assign v_6964 = v_4491;
assign v_6966 = v_6963 & v_6965;
assign v_6968 = v_6924 & v_6967;
assign v_6970 = v_4487;
assign v_6972 = v_6969 & v_6971;
assign v_6974 = v_6921 & v_6973;
assign v_6976 = v_4483;
assign v_6978 = v_6975 & v_6977;
assign v_6980 = v_6918 & v_6979;
assign v_6982 = v_4479;
assign v_6984 = v_6981 & v_6983;
assign v_6986 = v_6915 & v_6985;
assign v_6988 = v_4475;
assign v_6990 = v_6987 & v_6989;
assign v_6992 = v_6912 & v_6991;
assign v_6994 = v_4471;
assign v_6996 = v_6993 & v_6995;
assign v_6998 = v_6909 & v_6997;
assign v_7000 = v_4467;
assign v_7002 = v_6999 & v_7001;
assign v_7004 = v_6906 & v_7003;
assign v_7006 = v_4463;
assign v_7008 = v_7005 & v_7007;
assign v_7010 = v_6903 & v_7009;
assign v_7012 = v_4459;
assign v_7014 = v_7011 & v_7013;
assign v_7016 = v_6900 & v_7015;
assign v_7018 = v_2635;
assign v_7020 = v_7017 & v_7019;
assign v_7022 = v_6897 & v_7021;
assign v_7024 = v_2631;
assign v_7026 = v_7023 & v_7025;
assign v_7028 = v_6894 & v_7027;
assign v_7030 = v_2627;
assign v_7032 = v_7029 & v_7031;
assign v_7034 = v_6891 & v_7033;
assign v_7036 = v_2623;
assign v_7038 = v_7035 & v_7037;
assign v_7039 = v_7038;
assign v_7041 = v_4507;
assign v_7042 = v_2688;
assign v_7043 = v_7042;
assign v_7044 = v_7041 & v_7043;
assign v_7045 = v_7044;
assign v_7046 = v_6936 & v_7045;
assign v_7048 = v_6946 & v_7047;
assign v_7049 = v_6935 & v_7045;
assign v_7051 = v_6933 & v_7050;
assign v_7053 = v_6952 & v_7052;
assign v_7054 = v_6932 & v_7050;
assign v_7056 = v_6930 & v_7055;
assign v_7058 = v_6958 & v_7057;
assign v_7059 = v_6929 & v_7055;
assign v_7061 = v_6927 & v_7060;
assign v_7063 = v_6964 & v_7062;
assign v_7064 = v_6926 & v_7060;
assign v_7066 = v_6924 & v_7065;
assign v_7068 = v_6970 & v_7067;
assign v_7069 = v_6923 & v_7065;
assign v_7071 = v_6921 & v_7070;
assign v_7073 = v_6976 & v_7072;
assign v_7074 = v_6920 & v_7070;
assign v_7076 = v_6918 & v_7075;
assign v_7078 = v_6982 & v_7077;
assign v_7079 = v_6917 & v_7075;
assign v_7081 = v_6915 & v_7080;
assign v_7083 = v_6988 & v_7082;
assign v_7084 = v_6914 & v_7080;
assign v_7086 = v_6912 & v_7085;
assign v_7088 = v_6994 & v_7087;
assign v_7089 = v_6911 & v_7085;
assign v_7091 = v_6909 & v_7090;
assign v_7093 = v_7000 & v_7092;
assign v_7094 = v_6908 & v_7090;
assign v_7096 = v_6906 & v_7095;
assign v_7098 = v_7006 & v_7097;
assign v_7099 = v_6905 & v_7095;
assign v_7101 = v_6903 & v_7100;
assign v_7103 = v_7012 & v_7102;
assign v_7104 = v_6902 & v_7100;
assign v_7106 = v_6900 & v_7105;
assign v_7108 = v_7018 & v_7107;
assign v_7109 = v_6899 & v_7105;
assign v_7111 = v_6897 & v_7110;
assign v_7113 = v_7024 & v_7112;
assign v_7114 = v_6896 & v_7110;
assign v_7116 = v_6894 & v_7115;
assign v_7118 = v_7030 & v_7117;
assign v_7119 = v_6893 & v_7115;
assign v_7121 = v_6891 & v_7120;
assign v_7123 = v_7036 & v_7122;
assign v_7124 = v_6890 & v_7120;
assign v_7126 = v_7125;
assign v_7128 = v_7040 & v_7127;
assign v_7129 = v_7128;
assign v_7131 = v_7130;
assign v_7133 = ~v_2883;
assign v_7134 = ~v_4444;
assign v_7135 = v_4444;
assign v_7136 = ~v_2887;
assign v_7137 = ~v_4448;
assign v_7138 = v_4448;
assign v_7139 = ~v_2891;
assign v_7140 = ~v_4452;
assign v_7141 = v_4452;
assign v_7142 = ~v_2895;
assign v_7143 = ~v_4456;
assign v_7144 = v_4456;
assign v_7145 = ~v_4459;
assign v_7146 = ~v_2900;
assign v_7147 = v_2900;
assign v_7148 = ~v_4463;
assign v_7149 = ~v_2904;
assign v_7150 = v_2904;
assign v_7151 = ~v_4467;
assign v_7152 = ~v_2908;
assign v_7153 = v_2908;
assign v_7154 = ~v_4471;
assign v_7155 = ~v_2912;
assign v_7156 = v_2912;
assign v_7157 = ~v_4475;
assign v_7158 = ~v_2916;
assign v_7159 = v_2916;
assign v_7160 = ~v_4479;
assign v_7161 = ~v_2920;
assign v_7162 = v_2920;
assign v_7163 = ~v_4483;
assign v_7164 = ~v_2924;
assign v_7165 = v_2924;
assign v_7166 = ~v_4487;
assign v_7167 = ~v_2928;
assign v_7168 = v_2928;
assign v_7169 = ~v_4491;
assign v_7170 = ~v_2932;
assign v_7171 = v_2932;
assign v_7172 = ~v_4495;
assign v_7173 = ~v_2936;
assign v_7174 = v_2936;
assign v_7175 = ~v_4499;
assign v_7176 = ~v_2940;
assign v_7177 = v_2940;
assign v_7178 = ~v_4503;
assign v_7179 = ~v_2944;
assign v_7180 = v_2944;
assign v_7181 = ~v_4507;
assign v_7182 = ~v_2948;
assign v_7183 = v_7182;
assign v_7185 = v_7184;
assign v_7187 = v_7179 & v_7186;
assign v_7189 = v_4503;
assign v_7191 = v_7188 & v_7190;
assign v_7193 = v_7176 & v_7192;
assign v_7195 = v_4499;
assign v_7197 = v_7194 & v_7196;
assign v_7199 = v_7173 & v_7198;
assign v_7201 = v_4495;
assign v_7203 = v_7200 & v_7202;
assign v_7205 = v_7170 & v_7204;
assign v_7207 = v_4491;
assign v_7209 = v_7206 & v_7208;
assign v_7211 = v_7167 & v_7210;
assign v_7213 = v_4487;
assign v_7215 = v_7212 & v_7214;
assign v_7217 = v_7164 & v_7216;
assign v_7219 = v_4483;
assign v_7221 = v_7218 & v_7220;
assign v_7223 = v_7161 & v_7222;
assign v_7225 = v_4479;
assign v_7227 = v_7224 & v_7226;
assign v_7229 = v_7158 & v_7228;
assign v_7231 = v_4475;
assign v_7233 = v_7230 & v_7232;
assign v_7235 = v_7155 & v_7234;
assign v_7237 = v_4471;
assign v_7239 = v_7236 & v_7238;
assign v_7241 = v_7152 & v_7240;
assign v_7243 = v_4467;
assign v_7245 = v_7242 & v_7244;
assign v_7247 = v_7149 & v_7246;
assign v_7249 = v_4463;
assign v_7251 = v_7248 & v_7250;
assign v_7253 = v_7146 & v_7252;
assign v_7255 = v_4459;
assign v_7257 = v_7254 & v_7256;
assign v_7259 = v_7143 & v_7258;
assign v_7261 = v_2895;
assign v_7263 = v_7260 & v_7262;
assign v_7265 = v_7140 & v_7264;
assign v_7267 = v_2891;
assign v_7269 = v_7266 & v_7268;
assign v_7271 = v_7137 & v_7270;
assign v_7273 = v_2887;
assign v_7275 = v_7272 & v_7274;
assign v_7277 = v_7134 & v_7276;
assign v_7279 = v_2883;
assign v_7281 = v_7278 & v_7280;
assign v_7282 = v_7281;
assign v_7284 = v_4507;
assign v_7285 = v_2948;
assign v_7286 = v_7285;
assign v_7287 = v_7284 & v_7286;
assign v_7288 = v_7287;
assign v_7289 = v_7179 & v_7288;
assign v_7291 = v_7189 & v_7290;
assign v_7292 = v_7178 & v_7288;
assign v_7294 = v_7176 & v_7293;
assign v_7296 = v_7195 & v_7295;
assign v_7297 = v_7175 & v_7293;
assign v_7299 = v_7173 & v_7298;
assign v_7301 = v_7201 & v_7300;
assign v_7302 = v_7172 & v_7298;
assign v_7304 = v_7170 & v_7303;
assign v_7306 = v_7207 & v_7305;
assign v_7307 = v_7169 & v_7303;
assign v_7309 = v_7167 & v_7308;
assign v_7311 = v_7213 & v_7310;
assign v_7312 = v_7166 & v_7308;
assign v_7314 = v_7164 & v_7313;
assign v_7316 = v_7219 & v_7315;
assign v_7317 = v_7163 & v_7313;
assign v_7319 = v_7161 & v_7318;
assign v_7321 = v_7225 & v_7320;
assign v_7322 = v_7160 & v_7318;
assign v_7324 = v_7158 & v_7323;
assign v_7326 = v_7231 & v_7325;
assign v_7327 = v_7157 & v_7323;
assign v_7329 = v_7155 & v_7328;
assign v_7331 = v_7237 & v_7330;
assign v_7332 = v_7154 & v_7328;
assign v_7334 = v_7152 & v_7333;
assign v_7336 = v_7243 & v_7335;
assign v_7337 = v_7151 & v_7333;
assign v_7339 = v_7149 & v_7338;
assign v_7341 = v_7249 & v_7340;
assign v_7342 = v_7148 & v_7338;
assign v_7344 = v_7146 & v_7343;
assign v_7346 = v_7255 & v_7345;
assign v_7347 = v_7145 & v_7343;
assign v_7349 = v_7143 & v_7348;
assign v_7351 = v_7261 & v_7350;
assign v_7352 = v_7142 & v_7348;
assign v_7354 = v_7140 & v_7353;
assign v_7356 = v_7267 & v_7355;
assign v_7357 = v_7139 & v_7353;
assign v_7359 = v_7137 & v_7358;
assign v_7361 = v_7273 & v_7360;
assign v_7362 = v_7136 & v_7358;
assign v_7364 = v_7134 & v_7363;
assign v_7366 = v_7279 & v_7365;
assign v_7367 = v_7133 & v_7363;
assign v_7369 = v_7368;
assign v_7371 = v_7283 & v_7370;
assign v_7372 = v_7371;
assign v_7374 = v_7373;
assign v_7376 = ~v_3143;
assign v_7377 = ~v_4444;
assign v_7378 = v_4444;
assign v_7379 = ~v_3147;
assign v_7380 = ~v_4448;
assign v_7381 = v_4448;
assign v_7382 = ~v_3151;
assign v_7383 = ~v_4452;
assign v_7384 = v_4452;
assign v_7385 = ~v_3155;
assign v_7386 = ~v_4456;
assign v_7387 = v_4456;
assign v_7388 = ~v_4459;
assign v_7389 = ~v_3160;
assign v_7390 = v_3160;
assign v_7391 = ~v_4463;
assign v_7392 = ~v_3164;
assign v_7393 = v_3164;
assign v_7394 = ~v_4467;
assign v_7395 = ~v_3168;
assign v_7396 = v_3168;
assign v_7397 = ~v_4471;
assign v_7398 = ~v_3172;
assign v_7399 = v_3172;
assign v_7400 = ~v_4475;
assign v_7401 = ~v_3176;
assign v_7402 = v_3176;
assign v_7403 = ~v_4479;
assign v_7404 = ~v_3180;
assign v_7405 = v_3180;
assign v_7406 = ~v_4483;
assign v_7407 = ~v_3184;
assign v_7408 = v_3184;
assign v_7409 = ~v_4487;
assign v_7410 = ~v_3188;
assign v_7411 = v_3188;
assign v_7412 = ~v_4491;
assign v_7413 = ~v_3192;
assign v_7414 = v_3192;
assign v_7415 = ~v_4495;
assign v_7416 = ~v_3196;
assign v_7417 = v_3196;
assign v_7418 = ~v_4499;
assign v_7419 = ~v_3200;
assign v_7420 = v_3200;
assign v_7421 = ~v_4503;
assign v_7422 = ~v_3204;
assign v_7423 = v_3204;
assign v_7424 = ~v_4507;
assign v_7425 = ~v_3208;
assign v_7426 = v_7425;
assign v_7428 = v_7427;
assign v_7430 = v_7422 & v_7429;
assign v_7432 = v_4503;
assign v_7434 = v_7431 & v_7433;
assign v_7436 = v_7419 & v_7435;
assign v_7438 = v_4499;
assign v_7440 = v_7437 & v_7439;
assign v_7442 = v_7416 & v_7441;
assign v_7444 = v_4495;
assign v_7446 = v_7443 & v_7445;
assign v_7448 = v_7413 & v_7447;
assign v_7450 = v_4491;
assign v_7452 = v_7449 & v_7451;
assign v_7454 = v_7410 & v_7453;
assign v_7456 = v_4487;
assign v_7458 = v_7455 & v_7457;
assign v_7460 = v_7407 & v_7459;
assign v_7462 = v_4483;
assign v_7464 = v_7461 & v_7463;
assign v_7466 = v_7404 & v_7465;
assign v_7468 = v_4479;
assign v_7470 = v_7467 & v_7469;
assign v_7472 = v_7401 & v_7471;
assign v_7474 = v_4475;
assign v_7476 = v_7473 & v_7475;
assign v_7478 = v_7398 & v_7477;
assign v_7480 = v_4471;
assign v_7482 = v_7479 & v_7481;
assign v_7484 = v_7395 & v_7483;
assign v_7486 = v_4467;
assign v_7488 = v_7485 & v_7487;
assign v_7490 = v_7392 & v_7489;
assign v_7492 = v_4463;
assign v_7494 = v_7491 & v_7493;
assign v_7496 = v_7389 & v_7495;
assign v_7498 = v_4459;
assign v_7500 = v_7497 & v_7499;
assign v_7502 = v_7386 & v_7501;
assign v_7504 = v_3155;
assign v_7506 = v_7503 & v_7505;
assign v_7508 = v_7383 & v_7507;
assign v_7510 = v_3151;
assign v_7512 = v_7509 & v_7511;
assign v_7514 = v_7380 & v_7513;
assign v_7516 = v_3147;
assign v_7518 = v_7515 & v_7517;
assign v_7520 = v_7377 & v_7519;
assign v_7522 = v_3143;
assign v_7524 = v_7521 & v_7523;
assign v_7525 = v_7524;
assign v_7527 = v_4507;
assign v_7528 = v_3208;
assign v_7529 = v_7528;
assign v_7530 = v_7527 & v_7529;
assign v_7531 = v_7530;
assign v_7532 = v_7422 & v_7531;
assign v_7534 = v_7432 & v_7533;
assign v_7535 = v_7421 & v_7531;
assign v_7537 = v_7419 & v_7536;
assign v_7539 = v_7438 & v_7538;
assign v_7540 = v_7418 & v_7536;
assign v_7542 = v_7416 & v_7541;
assign v_7544 = v_7444 & v_7543;
assign v_7545 = v_7415 & v_7541;
assign v_7547 = v_7413 & v_7546;
assign v_7549 = v_7450 & v_7548;
assign v_7550 = v_7412 & v_7546;
assign v_7552 = v_7410 & v_7551;
assign v_7554 = v_7456 & v_7553;
assign v_7555 = v_7409 & v_7551;
assign v_7557 = v_7407 & v_7556;
assign v_7559 = v_7462 & v_7558;
assign v_7560 = v_7406 & v_7556;
assign v_7562 = v_7404 & v_7561;
assign v_7564 = v_7468 & v_7563;
assign v_7565 = v_7403 & v_7561;
assign v_7567 = v_7401 & v_7566;
assign v_7569 = v_7474 & v_7568;
assign v_7570 = v_7400 & v_7566;
assign v_7572 = v_7398 & v_7571;
assign v_7574 = v_7480 & v_7573;
assign v_7575 = v_7397 & v_7571;
assign v_7577 = v_7395 & v_7576;
assign v_7579 = v_7486 & v_7578;
assign v_7580 = v_7394 & v_7576;
assign v_7582 = v_7392 & v_7581;
assign v_7584 = v_7492 & v_7583;
assign v_7585 = v_7391 & v_7581;
assign v_7587 = v_7389 & v_7586;
assign v_7589 = v_7498 & v_7588;
assign v_7590 = v_7388 & v_7586;
assign v_7592 = v_7386 & v_7591;
assign v_7594 = v_7504 & v_7593;
assign v_7595 = v_7385 & v_7591;
assign v_7597 = v_7383 & v_7596;
assign v_7599 = v_7510 & v_7598;
assign v_7600 = v_7382 & v_7596;
assign v_7602 = v_7380 & v_7601;
assign v_7604 = v_7516 & v_7603;
assign v_7605 = v_7379 & v_7601;
assign v_7607 = v_7377 & v_7606;
assign v_7609 = v_7522 & v_7608;
assign v_7610 = v_7376 & v_7606;
assign v_7612 = v_7611;
assign v_7614 = v_7526 & v_7613;
assign v_7615 = v_7614;
assign v_7617 = v_7616;
assign v_7619 = ~v_3403;
assign v_7620 = ~v_4444;
assign v_7621 = v_4444;
assign v_7622 = ~v_3407;
assign v_7623 = ~v_4448;
assign v_7624 = v_4448;
assign v_7625 = ~v_3411;
assign v_7626 = ~v_4452;
assign v_7627 = v_4452;
assign v_7628 = ~v_3415;
assign v_7629 = ~v_4456;
assign v_7630 = v_4456;
assign v_7631 = ~v_4459;
assign v_7632 = ~v_3420;
assign v_7633 = v_3420;
assign v_7634 = ~v_4463;
assign v_7635 = ~v_3424;
assign v_7636 = v_3424;
assign v_7637 = ~v_4467;
assign v_7638 = ~v_3428;
assign v_7639 = v_3428;
assign v_7640 = ~v_4471;
assign v_7641 = ~v_3432;
assign v_7642 = v_3432;
assign v_7643 = ~v_4475;
assign v_7644 = ~v_3436;
assign v_7645 = v_3436;
assign v_7646 = ~v_4479;
assign v_7647 = ~v_3440;
assign v_7648 = v_3440;
assign v_7649 = ~v_4483;
assign v_7650 = ~v_3444;
assign v_7651 = v_3444;
assign v_7652 = ~v_4487;
assign v_7653 = ~v_3448;
assign v_7654 = v_3448;
assign v_7655 = ~v_4491;
assign v_7656 = ~v_3452;
assign v_7657 = v_3452;
assign v_7658 = ~v_4495;
assign v_7659 = ~v_3456;
assign v_7660 = v_3456;
assign v_7661 = ~v_4499;
assign v_7662 = ~v_3460;
assign v_7663 = v_3460;
assign v_7664 = ~v_4503;
assign v_7665 = ~v_3464;
assign v_7666 = v_3464;
assign v_7667 = ~v_4507;
assign v_7668 = ~v_3468;
assign v_7669 = v_7668;
assign v_7671 = v_7670;
assign v_7673 = v_7665 & v_7672;
assign v_7675 = v_4503;
assign v_7677 = v_7674 & v_7676;
assign v_7679 = v_7662 & v_7678;
assign v_7681 = v_4499;
assign v_7683 = v_7680 & v_7682;
assign v_7685 = v_7659 & v_7684;
assign v_7687 = v_4495;
assign v_7689 = v_7686 & v_7688;
assign v_7691 = v_7656 & v_7690;
assign v_7693 = v_4491;
assign v_7695 = v_7692 & v_7694;
assign v_7697 = v_7653 & v_7696;
assign v_7699 = v_4487;
assign v_7701 = v_7698 & v_7700;
assign v_7703 = v_7650 & v_7702;
assign v_7705 = v_4483;
assign v_7707 = v_7704 & v_7706;
assign v_7709 = v_7647 & v_7708;
assign v_7711 = v_4479;
assign v_7713 = v_7710 & v_7712;
assign v_7715 = v_7644 & v_7714;
assign v_7717 = v_4475;
assign v_7719 = v_7716 & v_7718;
assign v_7721 = v_7641 & v_7720;
assign v_7723 = v_4471;
assign v_7725 = v_7722 & v_7724;
assign v_7727 = v_7638 & v_7726;
assign v_7729 = v_4467;
assign v_7731 = v_7728 & v_7730;
assign v_7733 = v_7635 & v_7732;
assign v_7735 = v_4463;
assign v_7737 = v_7734 & v_7736;
assign v_7739 = v_7632 & v_7738;
assign v_7741 = v_4459;
assign v_7743 = v_7740 & v_7742;
assign v_7745 = v_7629 & v_7744;
assign v_7747 = v_3415;
assign v_7749 = v_7746 & v_7748;
assign v_7751 = v_7626 & v_7750;
assign v_7753 = v_3411;
assign v_7755 = v_7752 & v_7754;
assign v_7757 = v_7623 & v_7756;
assign v_7759 = v_3407;
assign v_7761 = v_7758 & v_7760;
assign v_7763 = v_7620 & v_7762;
assign v_7765 = v_3403;
assign v_7767 = v_7764 & v_7766;
assign v_7768 = v_7767;
assign v_7770 = v_4507;
assign v_7771 = v_3468;
assign v_7772 = v_7771;
assign v_7773 = v_7770 & v_7772;
assign v_7774 = v_7773;
assign v_7775 = v_7665 & v_7774;
assign v_7777 = v_7675 & v_7776;
assign v_7778 = v_7664 & v_7774;
assign v_7780 = v_7662 & v_7779;
assign v_7782 = v_7681 & v_7781;
assign v_7783 = v_7661 & v_7779;
assign v_7785 = v_7659 & v_7784;
assign v_7787 = v_7687 & v_7786;
assign v_7788 = v_7658 & v_7784;
assign v_7790 = v_7656 & v_7789;
assign v_7792 = v_7693 & v_7791;
assign v_7793 = v_7655 & v_7789;
assign v_7795 = v_7653 & v_7794;
assign v_7797 = v_7699 & v_7796;
assign v_7798 = v_7652 & v_7794;
assign v_7800 = v_7650 & v_7799;
assign v_7802 = v_7705 & v_7801;
assign v_7803 = v_7649 & v_7799;
assign v_7805 = v_7647 & v_7804;
assign v_7807 = v_7711 & v_7806;
assign v_7808 = v_7646 & v_7804;
assign v_7810 = v_7644 & v_7809;
assign v_7812 = v_7717 & v_7811;
assign v_7813 = v_7643 & v_7809;
assign v_7815 = v_7641 & v_7814;
assign v_7817 = v_7723 & v_7816;
assign v_7818 = v_7640 & v_7814;
assign v_7820 = v_7638 & v_7819;
assign v_7822 = v_7729 & v_7821;
assign v_7823 = v_7637 & v_7819;
assign v_7825 = v_7635 & v_7824;
assign v_7827 = v_7735 & v_7826;
assign v_7828 = v_7634 & v_7824;
assign v_7830 = v_7632 & v_7829;
assign v_7832 = v_7741 & v_7831;
assign v_7833 = v_7631 & v_7829;
assign v_7835 = v_7629 & v_7834;
assign v_7837 = v_7747 & v_7836;
assign v_7838 = v_7628 & v_7834;
assign v_7840 = v_7626 & v_7839;
assign v_7842 = v_7753 & v_7841;
assign v_7843 = v_7625 & v_7839;
assign v_7845 = v_7623 & v_7844;
assign v_7847 = v_7759 & v_7846;
assign v_7848 = v_7622 & v_7844;
assign v_7850 = v_7620 & v_7849;
assign v_7852 = v_7765 & v_7851;
assign v_7853 = v_7619 & v_7849;
assign v_7855 = v_7854;
assign v_7857 = v_7769 & v_7856;
assign v_7858 = v_7857;
assign v_7860 = v_7859;
assign v_7862 = ~v_3663;
assign v_7863 = ~v_4444;
assign v_7864 = v_4444;
assign v_7865 = ~v_3667;
assign v_7866 = ~v_4448;
assign v_7867 = v_4448;
assign v_7868 = ~v_3671;
assign v_7869 = ~v_4452;
assign v_7870 = v_4452;
assign v_7871 = ~v_3675;
assign v_7872 = ~v_4456;
assign v_7873 = v_4456;
assign v_7874 = ~v_4459;
assign v_7875 = ~v_3680;
assign v_7876 = v_3680;
assign v_7877 = ~v_4463;
assign v_7878 = ~v_3684;
assign v_7879 = v_3684;
assign v_7880 = ~v_4467;
assign v_7881 = ~v_3688;
assign v_7882 = v_3688;
assign v_7883 = ~v_4471;
assign v_7884 = ~v_3692;
assign v_7885 = v_3692;
assign v_7886 = ~v_4475;
assign v_7887 = ~v_3696;
assign v_7888 = v_3696;
assign v_7889 = ~v_4479;
assign v_7890 = ~v_3700;
assign v_7891 = v_3700;
assign v_7892 = ~v_4483;
assign v_7893 = ~v_3704;
assign v_7894 = v_3704;
assign v_7895 = ~v_4487;
assign v_7896 = ~v_3708;
assign v_7897 = v_3708;
assign v_7898 = ~v_4491;
assign v_7899 = ~v_3712;
assign v_7900 = v_3712;
assign v_7901 = ~v_4495;
assign v_7902 = ~v_3716;
assign v_7903 = v_3716;
assign v_7904 = ~v_4499;
assign v_7905 = ~v_3720;
assign v_7906 = v_3720;
assign v_7907 = ~v_4503;
assign v_7908 = ~v_3724;
assign v_7909 = v_3724;
assign v_7910 = ~v_4507;
assign v_7911 = ~v_3728;
assign v_7912 = v_7911;
assign v_7914 = v_7913;
assign v_7916 = v_7908 & v_7915;
assign v_7918 = v_4503;
assign v_7920 = v_7917 & v_7919;
assign v_7922 = v_7905 & v_7921;
assign v_7924 = v_4499;
assign v_7926 = v_7923 & v_7925;
assign v_7928 = v_7902 & v_7927;
assign v_7930 = v_4495;
assign v_7932 = v_7929 & v_7931;
assign v_7934 = v_7899 & v_7933;
assign v_7936 = v_4491;
assign v_7938 = v_7935 & v_7937;
assign v_7940 = v_7896 & v_7939;
assign v_7942 = v_4487;
assign v_7944 = v_7941 & v_7943;
assign v_7946 = v_7893 & v_7945;
assign v_7948 = v_4483;
assign v_7950 = v_7947 & v_7949;
assign v_7952 = v_7890 & v_7951;
assign v_7954 = v_4479;
assign v_7956 = v_7953 & v_7955;
assign v_7958 = v_7887 & v_7957;
assign v_7960 = v_4475;
assign v_7962 = v_7959 & v_7961;
assign v_7964 = v_7884 & v_7963;
assign v_7966 = v_4471;
assign v_7968 = v_7965 & v_7967;
assign v_7970 = v_7881 & v_7969;
assign v_7972 = v_4467;
assign v_7974 = v_7971 & v_7973;
assign v_7976 = v_7878 & v_7975;
assign v_7978 = v_4463;
assign v_7980 = v_7977 & v_7979;
assign v_7982 = v_7875 & v_7981;
assign v_7984 = v_4459;
assign v_7986 = v_7983 & v_7985;
assign v_7988 = v_7872 & v_7987;
assign v_7990 = v_3675;
assign v_7992 = v_7989 & v_7991;
assign v_7994 = v_7869 & v_7993;
assign v_7996 = v_3671;
assign v_7998 = v_7995 & v_7997;
assign v_8000 = v_7866 & v_7999;
assign v_8002 = v_3667;
assign v_8004 = v_8001 & v_8003;
assign v_8006 = v_7863 & v_8005;
assign v_8008 = v_3663;
assign v_8010 = v_8007 & v_8009;
assign v_8011 = v_8010;
assign v_8013 = v_4507;
assign v_8014 = v_3728;
assign v_8015 = v_8014;
assign v_8016 = v_8013 & v_8015;
assign v_8017 = v_8016;
assign v_8018 = v_7908 & v_8017;
assign v_8020 = v_7918 & v_8019;
assign v_8021 = v_7907 & v_8017;
assign v_8023 = v_7905 & v_8022;
assign v_8025 = v_7924 & v_8024;
assign v_8026 = v_7904 & v_8022;
assign v_8028 = v_7902 & v_8027;
assign v_8030 = v_7930 & v_8029;
assign v_8031 = v_7901 & v_8027;
assign v_8033 = v_7899 & v_8032;
assign v_8035 = v_7936 & v_8034;
assign v_8036 = v_7898 & v_8032;
assign v_8038 = v_7896 & v_8037;
assign v_8040 = v_7942 & v_8039;
assign v_8041 = v_7895 & v_8037;
assign v_8043 = v_7893 & v_8042;
assign v_8045 = v_7948 & v_8044;
assign v_8046 = v_7892 & v_8042;
assign v_8048 = v_7890 & v_8047;
assign v_8050 = v_7954 & v_8049;
assign v_8051 = v_7889 & v_8047;
assign v_8053 = v_7887 & v_8052;
assign v_8055 = v_7960 & v_8054;
assign v_8056 = v_7886 & v_8052;
assign v_8058 = v_7884 & v_8057;
assign v_8060 = v_7966 & v_8059;
assign v_8061 = v_7883 & v_8057;
assign v_8063 = v_7881 & v_8062;
assign v_8065 = v_7972 & v_8064;
assign v_8066 = v_7880 & v_8062;
assign v_8068 = v_7878 & v_8067;
assign v_8070 = v_7978 & v_8069;
assign v_8071 = v_7877 & v_8067;
assign v_8073 = v_7875 & v_8072;
assign v_8075 = v_7984 & v_8074;
assign v_8076 = v_7874 & v_8072;
assign v_8078 = v_7872 & v_8077;
assign v_8080 = v_7990 & v_8079;
assign v_8081 = v_7871 & v_8077;
assign v_8083 = v_7869 & v_8082;
assign v_8085 = v_7996 & v_8084;
assign v_8086 = v_7868 & v_8082;
assign v_8088 = v_7866 & v_8087;
assign v_8090 = v_8002 & v_8089;
assign v_8091 = v_7865 & v_8087;
assign v_8093 = v_7863 & v_8092;
assign v_8095 = v_8008 & v_8094;
assign v_8096 = v_7862 & v_8092;
assign v_8098 = v_8097;
assign v_8100 = v_8012 & v_8099;
assign v_8101 = v_8100;
assign v_8103 = v_8102;
assign v_8105 = ~v_3923;
assign v_8106 = ~v_4444;
assign v_8107 = v_4444;
assign v_8108 = ~v_3927;
assign v_8109 = ~v_4448;
assign v_8110 = v_4448;
assign v_8111 = ~v_3931;
assign v_8112 = ~v_4452;
assign v_8113 = v_4452;
assign v_8114 = ~v_3935;
assign v_8115 = ~v_4456;
assign v_8116 = v_4456;
assign v_8117 = ~v_4459;
assign v_8118 = ~v_3940;
assign v_8119 = v_3940;
assign v_8120 = ~v_4463;
assign v_8121 = ~v_3944;
assign v_8122 = v_3944;
assign v_8123 = ~v_4467;
assign v_8124 = ~v_3948;
assign v_8125 = v_3948;
assign v_8126 = ~v_4471;
assign v_8127 = ~v_3952;
assign v_8128 = v_3952;
assign v_8129 = ~v_4475;
assign v_8130 = ~v_3956;
assign v_8131 = v_3956;
assign v_8132 = ~v_4479;
assign v_8133 = ~v_3960;
assign v_8134 = v_3960;
assign v_8135 = ~v_4483;
assign v_8136 = ~v_3964;
assign v_8137 = v_3964;
assign v_8138 = ~v_4487;
assign v_8139 = ~v_3968;
assign v_8140 = v_3968;
assign v_8141 = ~v_4491;
assign v_8142 = ~v_3972;
assign v_8143 = v_3972;
assign v_8144 = ~v_4495;
assign v_8145 = ~v_3976;
assign v_8146 = v_3976;
assign v_8147 = ~v_4499;
assign v_8148 = ~v_3980;
assign v_8149 = v_3980;
assign v_8150 = ~v_4503;
assign v_8151 = ~v_3984;
assign v_8152 = v_3984;
assign v_8153 = ~v_4507;
assign v_8154 = ~v_3988;
assign v_8155 = v_8154;
assign v_8157 = v_8156;
assign v_8159 = v_8151 & v_8158;
assign v_8161 = v_4503;
assign v_8163 = v_8160 & v_8162;
assign v_8165 = v_8148 & v_8164;
assign v_8167 = v_4499;
assign v_8169 = v_8166 & v_8168;
assign v_8171 = v_8145 & v_8170;
assign v_8173 = v_4495;
assign v_8175 = v_8172 & v_8174;
assign v_8177 = v_8142 & v_8176;
assign v_8179 = v_4491;
assign v_8181 = v_8178 & v_8180;
assign v_8183 = v_8139 & v_8182;
assign v_8185 = v_4487;
assign v_8187 = v_8184 & v_8186;
assign v_8189 = v_8136 & v_8188;
assign v_8191 = v_4483;
assign v_8193 = v_8190 & v_8192;
assign v_8195 = v_8133 & v_8194;
assign v_8197 = v_4479;
assign v_8199 = v_8196 & v_8198;
assign v_8201 = v_8130 & v_8200;
assign v_8203 = v_4475;
assign v_8205 = v_8202 & v_8204;
assign v_8207 = v_8127 & v_8206;
assign v_8209 = v_4471;
assign v_8211 = v_8208 & v_8210;
assign v_8213 = v_8124 & v_8212;
assign v_8215 = v_4467;
assign v_8217 = v_8214 & v_8216;
assign v_8219 = v_8121 & v_8218;
assign v_8221 = v_4463;
assign v_8223 = v_8220 & v_8222;
assign v_8225 = v_8118 & v_8224;
assign v_8227 = v_4459;
assign v_8229 = v_8226 & v_8228;
assign v_8231 = v_8115 & v_8230;
assign v_8233 = v_3935;
assign v_8235 = v_8232 & v_8234;
assign v_8237 = v_8112 & v_8236;
assign v_8239 = v_3931;
assign v_8241 = v_8238 & v_8240;
assign v_8243 = v_8109 & v_8242;
assign v_8245 = v_3927;
assign v_8247 = v_8244 & v_8246;
assign v_8249 = v_8106 & v_8248;
assign v_8251 = v_3923;
assign v_8253 = v_8250 & v_8252;
assign v_8254 = v_8253;
assign v_8256 = v_4507;
assign v_8257 = v_3988;
assign v_8258 = v_8257;
assign v_8259 = v_8256 & v_8258;
assign v_8260 = v_8259;
assign v_8261 = v_8151 & v_8260;
assign v_8263 = v_8161 & v_8262;
assign v_8264 = v_8150 & v_8260;
assign v_8266 = v_8148 & v_8265;
assign v_8268 = v_8167 & v_8267;
assign v_8269 = v_8147 & v_8265;
assign v_8271 = v_8145 & v_8270;
assign v_8273 = v_8173 & v_8272;
assign v_8274 = v_8144 & v_8270;
assign v_8276 = v_8142 & v_8275;
assign v_8278 = v_8179 & v_8277;
assign v_8279 = v_8141 & v_8275;
assign v_8281 = v_8139 & v_8280;
assign v_8283 = v_8185 & v_8282;
assign v_8284 = v_8138 & v_8280;
assign v_8286 = v_8136 & v_8285;
assign v_8288 = v_8191 & v_8287;
assign v_8289 = v_8135 & v_8285;
assign v_8291 = v_8133 & v_8290;
assign v_8293 = v_8197 & v_8292;
assign v_8294 = v_8132 & v_8290;
assign v_8296 = v_8130 & v_8295;
assign v_8298 = v_8203 & v_8297;
assign v_8299 = v_8129 & v_8295;
assign v_8301 = v_8127 & v_8300;
assign v_8303 = v_8209 & v_8302;
assign v_8304 = v_8126 & v_8300;
assign v_8306 = v_8124 & v_8305;
assign v_8308 = v_8215 & v_8307;
assign v_8309 = v_8123 & v_8305;
assign v_8311 = v_8121 & v_8310;
assign v_8313 = v_8221 & v_8312;
assign v_8314 = v_8120 & v_8310;
assign v_8316 = v_8118 & v_8315;
assign v_8318 = v_8227 & v_8317;
assign v_8319 = v_8117 & v_8315;
assign v_8321 = v_8115 & v_8320;
assign v_8323 = v_8233 & v_8322;
assign v_8324 = v_8114 & v_8320;
assign v_8326 = v_8112 & v_8325;
assign v_8328 = v_8239 & v_8327;
assign v_8329 = v_8111 & v_8325;
assign v_8331 = v_8109 & v_8330;
assign v_8333 = v_8245 & v_8332;
assign v_8334 = v_8108 & v_8330;
assign v_8336 = v_8106 & v_8335;
assign v_8338 = v_8251 & v_8337;
assign v_8339 = v_8105 & v_8335;
assign v_8341 = v_8340;
assign v_8343 = v_8255 & v_8342;
assign v_8344 = v_8343;
assign v_8346 = v_8345;
assign v_8347 = ~v_4182;
assign v_8348 = ~v_4444;
assign v_8349 = v_4444;
assign v_8350 = ~v_4186;
assign v_8351 = ~v_4448;
assign v_8352 = v_4448;
assign v_8353 = ~v_4190;
assign v_8354 = ~v_4452;
assign v_8355 = v_4452;
assign v_8356 = ~v_4194;
assign v_8357 = ~v_4456;
assign v_8358 = v_4456;
assign v_8359 = ~v_4459;
assign v_8360 = ~v_4199;
assign v_8361 = v_4199;
assign v_8362 = ~v_4463;
assign v_8363 = ~v_4203;
assign v_8364 = v_4203;
assign v_8365 = ~v_4467;
assign v_8366 = ~v_4207;
assign v_8367 = v_4207;
assign v_8368 = ~v_4471;
assign v_8369 = ~v_4211;
assign v_8370 = v_4211;
assign v_8371 = ~v_4475;
assign v_8372 = ~v_4215;
assign v_8373 = v_4215;
assign v_8374 = ~v_4479;
assign v_8375 = ~v_4219;
assign v_8376 = v_4219;
assign v_8377 = ~v_4483;
assign v_8378 = ~v_4223;
assign v_8379 = v_4223;
assign v_8380 = ~v_4487;
assign v_8381 = ~v_4227;
assign v_8382 = v_4227;
assign v_8383 = ~v_4491;
assign v_8384 = ~v_4231;
assign v_8385 = v_4231;
assign v_8386 = ~v_4495;
assign v_8387 = ~v_4235;
assign v_8388 = v_4235;
assign v_8389 = ~v_4499;
assign v_8390 = ~v_4239;
assign v_8391 = v_4239;
assign v_8392 = ~v_4503;
assign v_8393 = ~v_4243;
assign v_8394 = v_4243;
assign v_8395 = ~v_4507;
assign v_8396 = ~v_4247;
assign v_8397 = v_8396;
assign v_8399 = v_8398;
assign v_8401 = v_8393 & v_8400;
assign v_8403 = v_4503;
assign v_8405 = v_8402 & v_8404;
assign v_8407 = v_8390 & v_8406;
assign v_8409 = v_4499;
assign v_8411 = v_8408 & v_8410;
assign v_8413 = v_8387 & v_8412;
assign v_8415 = v_4495;
assign v_8417 = v_8414 & v_8416;
assign v_8419 = v_8384 & v_8418;
assign v_8421 = v_4491;
assign v_8423 = v_8420 & v_8422;
assign v_8425 = v_8381 & v_8424;
assign v_8427 = v_4487;
assign v_8429 = v_8426 & v_8428;
assign v_8431 = v_8378 & v_8430;
assign v_8433 = v_4483;
assign v_8435 = v_8432 & v_8434;
assign v_8437 = v_8375 & v_8436;
assign v_8439 = v_4479;
assign v_8441 = v_8438 & v_8440;
assign v_8443 = v_8372 & v_8442;
assign v_8445 = v_4475;
assign v_8447 = v_8444 & v_8446;
assign v_8449 = v_8369 & v_8448;
assign v_8451 = v_4471;
assign v_8453 = v_8450 & v_8452;
assign v_8455 = v_8366 & v_8454;
assign v_8457 = v_4467;
assign v_8459 = v_8456 & v_8458;
assign v_8461 = v_8363 & v_8460;
assign v_8463 = v_4463;
assign v_8465 = v_8462 & v_8464;
assign v_8467 = v_8360 & v_8466;
assign v_8469 = v_4459;
assign v_8471 = v_8468 & v_8470;
assign v_8473 = v_8357 & v_8472;
assign v_8475 = v_4194;
assign v_8477 = v_8474 & v_8476;
assign v_8479 = v_8354 & v_8478;
assign v_8481 = v_4190;
assign v_8483 = v_8480 & v_8482;
assign v_8485 = v_8351 & v_8484;
assign v_8487 = v_4186;
assign v_8489 = v_8486 & v_8488;
assign v_8491 = v_8348 & v_8490;
assign v_8493 = v_4182;
assign v_8495 = v_8492 & v_8494;
assign v_8497 = ~v_8496;
assign v_8499 = v_4507;
assign v_8500 = v_4247;
assign v_8501 = v_8500;
assign v_8502 = v_8499 & v_8501;
assign v_8503 = v_8502;
assign v_8504 = v_8393 & v_8503;
assign v_8506 = v_8403 & v_8505;
assign v_8507 = v_8392 & v_8503;
assign v_8509 = v_8390 & v_8508;
assign v_8511 = v_8409 & v_8510;
assign v_8512 = v_8389 & v_8508;
assign v_8514 = v_8387 & v_8513;
assign v_8516 = v_8415 & v_8515;
assign v_8517 = v_8386 & v_8513;
assign v_8519 = v_8384 & v_8518;
assign v_8521 = v_8421 & v_8520;
assign v_8522 = v_8383 & v_8518;
assign v_8524 = v_8381 & v_8523;
assign v_8526 = v_8427 & v_8525;
assign v_8527 = v_8380 & v_8523;
assign v_8529 = v_8378 & v_8528;
assign v_8531 = v_8433 & v_8530;
assign v_8532 = v_8377 & v_8528;
assign v_8534 = v_8375 & v_8533;
assign v_8536 = v_8439 & v_8535;
assign v_8537 = v_8374 & v_8533;
assign v_8539 = v_8372 & v_8538;
assign v_8541 = v_8445 & v_8540;
assign v_8542 = v_8371 & v_8538;
assign v_8544 = v_8369 & v_8543;
assign v_8546 = v_8451 & v_8545;
assign v_8547 = v_8368 & v_8543;
assign v_8549 = v_8366 & v_8548;
assign v_8551 = v_8457 & v_8550;
assign v_8552 = v_8365 & v_8548;
assign v_8554 = v_8363 & v_8553;
assign v_8556 = v_8463 & v_8555;
assign v_8557 = v_8362 & v_8553;
assign v_8559 = v_8360 & v_8558;
assign v_8561 = v_8469 & v_8560;
assign v_8562 = v_8359 & v_8558;
assign v_8564 = v_8357 & v_8563;
assign v_8566 = v_8475 & v_8565;
assign v_8567 = v_8356 & v_8563;
assign v_8569 = v_8354 & v_8568;
assign v_8571 = v_8481 & v_8570;
assign v_8572 = v_8353 & v_8568;
assign v_8574 = v_8351 & v_8573;
assign v_8576 = v_8487 & v_8575;
assign v_8577 = v_8350 & v_8573;
assign v_8579 = v_8348 & v_8578;
assign v_8581 = v_8493 & v_8580;
assign v_8582 = v_8347 & v_8578;
assign v_8584 = v_8496;
assign v_8586 = v_8498 & v_8585;
assign v_8587 = v_8586;
assign v_8589 = v_8588;
assign v_8591 = ~v_6;
assign v_8593 = ~v_8592;
assign v_8594 = v_8592;
assign v_8595 = ~v_13;
assign v_8597 = ~v_8596;
assign v_8598 = v_8596;
assign v_8599 = ~v_18;
assign v_8601 = ~v_8600;
assign v_8602 = v_8600;
assign v_8603 = ~v_23;
assign v_8605 = ~v_8604;
assign v_8606 = v_8604;
assign v_8608 = ~v_8607;
assign v_8609 = ~v_30;
assign v_8610 = v_30;
assign v_8612 = ~v_8611;
assign v_8613 = ~v_35;
assign v_8614 = v_35;
assign v_8616 = ~v_8615;
assign v_8617 = ~v_40;
assign v_8618 = v_40;
assign v_8620 = ~v_8619;
assign v_8621 = ~v_45;
assign v_8622 = v_45;
assign v_8624 = ~v_8623;
assign v_8625 = ~v_50;
assign v_8626 = v_50;
assign v_8628 = ~v_8627;
assign v_8629 = ~v_55;
assign v_8630 = v_55;
assign v_8632 = ~v_8631;
assign v_8633 = ~v_60;
assign v_8634 = v_60;
assign v_8636 = ~v_8635;
assign v_8637 = ~v_65;
assign v_8638 = v_65;
assign v_8640 = ~v_8639;
assign v_8641 = ~v_70;
assign v_8642 = v_70;
assign v_8644 = ~v_8643;
assign v_8645 = ~v_75;
assign v_8646 = v_75;
assign v_8648 = ~v_8647;
assign v_8649 = ~v_80;
assign v_8650 = v_80;
assign v_8652 = ~v_8651;
assign v_8653 = ~v_85;
assign v_8654 = v_85;
assign v_8656 = ~v_8655;
assign v_8657 = ~v_90;
assign v_8658 = v_8657;
assign v_8660 = v_8659;
assign v_8662 = v_8653 & v_8661;
assign v_8664 = v_8651;
assign v_8666 = v_8663 & v_8665;
assign v_8668 = v_8649 & v_8667;
assign v_8670 = v_8647;
assign v_8672 = v_8669 & v_8671;
assign v_8674 = v_8645 & v_8673;
assign v_8676 = v_8643;
assign v_8678 = v_8675 & v_8677;
assign v_8680 = v_8641 & v_8679;
assign v_8682 = v_8639;
assign v_8684 = v_8681 & v_8683;
assign v_8686 = v_8637 & v_8685;
assign v_8688 = v_8635;
assign v_8690 = v_8687 & v_8689;
assign v_8692 = v_8633 & v_8691;
assign v_8694 = v_8631;
assign v_8696 = v_8693 & v_8695;
assign v_8698 = v_8629 & v_8697;
assign v_8700 = v_8627;
assign v_8702 = v_8699 & v_8701;
assign v_8704 = v_8625 & v_8703;
assign v_8706 = v_8623;
assign v_8708 = v_8705 & v_8707;
assign v_8710 = v_8621 & v_8709;
assign v_8712 = v_8619;
assign v_8714 = v_8711 & v_8713;
assign v_8716 = v_8617 & v_8715;
assign v_8718 = v_8615;
assign v_8720 = v_8717 & v_8719;
assign v_8722 = v_8613 & v_8721;
assign v_8724 = v_8611;
assign v_8726 = v_8723 & v_8725;
assign v_8728 = v_8609 & v_8727;
assign v_8730 = v_8607;
assign v_8732 = v_8729 & v_8731;
assign v_8734 = v_8605 & v_8733;
assign v_8736 = v_23;
assign v_8738 = v_8735 & v_8737;
assign v_8740 = v_8601 & v_8739;
assign v_8742 = v_18;
assign v_8744 = v_8741 & v_8743;
assign v_8746 = v_8597 & v_8745;
assign v_8748 = v_13;
assign v_8750 = v_8747 & v_8749;
assign v_8752 = v_8593 & v_8751;
assign v_8754 = v_6;
assign v_8756 = v_8753 & v_8755;
assign v_8757 = v_8756;
assign v_8759 = v_8655;
assign v_8760 = v_90;
assign v_8761 = v_8760;
assign v_8762 = v_8759 & v_8761;
assign v_8763 = v_8762;
assign v_8764 = v_8653 & v_8763;
assign v_8766 = v_8664 & v_8765;
assign v_8767 = v_8652 & v_8763;
assign v_8769 = v_8649 & v_8768;
assign v_8771 = v_8670 & v_8770;
assign v_8772 = v_8648 & v_8768;
assign v_8774 = v_8645 & v_8773;
assign v_8776 = v_8676 & v_8775;
assign v_8777 = v_8644 & v_8773;
assign v_8779 = v_8641 & v_8778;
assign v_8781 = v_8682 & v_8780;
assign v_8782 = v_8640 & v_8778;
assign v_8784 = v_8637 & v_8783;
assign v_8786 = v_8688 & v_8785;
assign v_8787 = v_8636 & v_8783;
assign v_8789 = v_8633 & v_8788;
assign v_8791 = v_8694 & v_8790;
assign v_8792 = v_8632 & v_8788;
assign v_8794 = v_8629 & v_8793;
assign v_8796 = v_8700 & v_8795;
assign v_8797 = v_8628 & v_8793;
assign v_8799 = v_8625 & v_8798;
assign v_8801 = v_8706 & v_8800;
assign v_8802 = v_8624 & v_8798;
assign v_8804 = v_8621 & v_8803;
assign v_8806 = v_8712 & v_8805;
assign v_8807 = v_8620 & v_8803;
assign v_8809 = v_8617 & v_8808;
assign v_8811 = v_8718 & v_8810;
assign v_8812 = v_8616 & v_8808;
assign v_8814 = v_8613 & v_8813;
assign v_8816 = v_8724 & v_8815;
assign v_8817 = v_8612 & v_8813;
assign v_8819 = v_8609 & v_8818;
assign v_8821 = v_8730 & v_8820;
assign v_8822 = v_8608 & v_8818;
assign v_8824 = v_8605 & v_8823;
assign v_8826 = v_8736 & v_8825;
assign v_8827 = v_8603 & v_8823;
assign v_8829 = v_8601 & v_8828;
assign v_8831 = v_8742 & v_8830;
assign v_8832 = v_8599 & v_8828;
assign v_8834 = v_8597 & v_8833;
assign v_8836 = v_8748 & v_8835;
assign v_8837 = v_8595 & v_8833;
assign v_8839 = v_8593 & v_8838;
assign v_8841 = v_8754 & v_8840;
assign v_8842 = v_8591 & v_8838;
assign v_8844 = v_8843;
assign v_8846 = v_8758 & v_8845;
assign v_8847 = v_8846;
assign v_8849 = v_8848;
assign v_8851 = ~v_283;
assign v_8852 = ~v_8592;
assign v_8853 = v_8592;
assign v_8854 = ~v_287;
assign v_8855 = ~v_8596;
assign v_8856 = v_8596;
assign v_8857 = ~v_291;
assign v_8858 = ~v_8600;
assign v_8859 = v_8600;
assign v_8860 = ~v_295;
assign v_8861 = ~v_8604;
assign v_8862 = v_8604;
assign v_8863 = ~v_8607;
assign v_8864 = ~v_300;
assign v_8865 = v_300;
assign v_8866 = ~v_8611;
assign v_8867 = ~v_304;
assign v_8868 = v_304;
assign v_8869 = ~v_8615;
assign v_8870 = ~v_308;
assign v_8871 = v_308;
assign v_8872 = ~v_8619;
assign v_8873 = ~v_312;
assign v_8874 = v_312;
assign v_8875 = ~v_8623;
assign v_8876 = ~v_316;
assign v_8877 = v_316;
assign v_8878 = ~v_8627;
assign v_8879 = ~v_320;
assign v_8880 = v_320;
assign v_8881 = ~v_8631;
assign v_8882 = ~v_324;
assign v_8883 = v_324;
assign v_8884 = ~v_8635;
assign v_8885 = ~v_328;
assign v_8886 = v_328;
assign v_8887 = ~v_8639;
assign v_8888 = ~v_332;
assign v_8889 = v_332;
assign v_8890 = ~v_8643;
assign v_8891 = ~v_336;
assign v_8892 = v_336;
assign v_8893 = ~v_8647;
assign v_8894 = ~v_340;
assign v_8895 = v_340;
assign v_8896 = ~v_8651;
assign v_8897 = ~v_344;
assign v_8898 = v_344;
assign v_8899 = ~v_8655;
assign v_8900 = ~v_348;
assign v_8901 = v_8900;
assign v_8903 = v_8902;
assign v_8905 = v_8897 & v_8904;
assign v_8907 = v_8651;
assign v_8909 = v_8906 & v_8908;
assign v_8911 = v_8894 & v_8910;
assign v_8913 = v_8647;
assign v_8915 = v_8912 & v_8914;
assign v_8917 = v_8891 & v_8916;
assign v_8919 = v_8643;
assign v_8921 = v_8918 & v_8920;
assign v_8923 = v_8888 & v_8922;
assign v_8925 = v_8639;
assign v_8927 = v_8924 & v_8926;
assign v_8929 = v_8885 & v_8928;
assign v_8931 = v_8635;
assign v_8933 = v_8930 & v_8932;
assign v_8935 = v_8882 & v_8934;
assign v_8937 = v_8631;
assign v_8939 = v_8936 & v_8938;
assign v_8941 = v_8879 & v_8940;
assign v_8943 = v_8627;
assign v_8945 = v_8942 & v_8944;
assign v_8947 = v_8876 & v_8946;
assign v_8949 = v_8623;
assign v_8951 = v_8948 & v_8950;
assign v_8953 = v_8873 & v_8952;
assign v_8955 = v_8619;
assign v_8957 = v_8954 & v_8956;
assign v_8959 = v_8870 & v_8958;
assign v_8961 = v_8615;
assign v_8963 = v_8960 & v_8962;
assign v_8965 = v_8867 & v_8964;
assign v_8967 = v_8611;
assign v_8969 = v_8966 & v_8968;
assign v_8971 = v_8864 & v_8970;
assign v_8973 = v_8607;
assign v_8975 = v_8972 & v_8974;
assign v_8977 = v_8861 & v_8976;
assign v_8979 = v_295;
assign v_8981 = v_8978 & v_8980;
assign v_8983 = v_8858 & v_8982;
assign v_8985 = v_291;
assign v_8987 = v_8984 & v_8986;
assign v_8989 = v_8855 & v_8988;
assign v_8991 = v_287;
assign v_8993 = v_8990 & v_8992;
assign v_8995 = v_8852 & v_8994;
assign v_8997 = v_283;
assign v_8999 = v_8996 & v_8998;
assign v_9000 = v_8999;
assign v_9002 = v_8655;
assign v_9003 = v_348;
assign v_9004 = v_9003;
assign v_9005 = v_9002 & v_9004;
assign v_9006 = v_9005;
assign v_9007 = v_8897 & v_9006;
assign v_9009 = v_8907 & v_9008;
assign v_9010 = v_8896 & v_9006;
assign v_9012 = v_8894 & v_9011;
assign v_9014 = v_8913 & v_9013;
assign v_9015 = v_8893 & v_9011;
assign v_9017 = v_8891 & v_9016;
assign v_9019 = v_8919 & v_9018;
assign v_9020 = v_8890 & v_9016;
assign v_9022 = v_8888 & v_9021;
assign v_9024 = v_8925 & v_9023;
assign v_9025 = v_8887 & v_9021;
assign v_9027 = v_8885 & v_9026;
assign v_9029 = v_8931 & v_9028;
assign v_9030 = v_8884 & v_9026;
assign v_9032 = v_8882 & v_9031;
assign v_9034 = v_8937 & v_9033;
assign v_9035 = v_8881 & v_9031;
assign v_9037 = v_8879 & v_9036;
assign v_9039 = v_8943 & v_9038;
assign v_9040 = v_8878 & v_9036;
assign v_9042 = v_8876 & v_9041;
assign v_9044 = v_8949 & v_9043;
assign v_9045 = v_8875 & v_9041;
assign v_9047 = v_8873 & v_9046;
assign v_9049 = v_8955 & v_9048;
assign v_9050 = v_8872 & v_9046;
assign v_9052 = v_8870 & v_9051;
assign v_9054 = v_8961 & v_9053;
assign v_9055 = v_8869 & v_9051;
assign v_9057 = v_8867 & v_9056;
assign v_9059 = v_8967 & v_9058;
assign v_9060 = v_8866 & v_9056;
assign v_9062 = v_8864 & v_9061;
assign v_9064 = v_8973 & v_9063;
assign v_9065 = v_8863 & v_9061;
assign v_9067 = v_8861 & v_9066;
assign v_9069 = v_8979 & v_9068;
assign v_9070 = v_8860 & v_9066;
assign v_9072 = v_8858 & v_9071;
assign v_9074 = v_8985 & v_9073;
assign v_9075 = v_8857 & v_9071;
assign v_9077 = v_8855 & v_9076;
assign v_9079 = v_8991 & v_9078;
assign v_9080 = v_8854 & v_9076;
assign v_9082 = v_8852 & v_9081;
assign v_9084 = v_8997 & v_9083;
assign v_9085 = v_8851 & v_9081;
assign v_9087 = v_9086;
assign v_9089 = v_9001 & v_9088;
assign v_9090 = v_9089;
assign v_9092 = v_9091;
assign v_9094 = ~v_543;
assign v_9095 = ~v_8592;
assign v_9096 = v_8592;
assign v_9097 = ~v_547;
assign v_9098 = ~v_8596;
assign v_9099 = v_8596;
assign v_9100 = ~v_551;
assign v_9101 = ~v_8600;
assign v_9102 = v_8600;
assign v_9103 = ~v_555;
assign v_9104 = ~v_8604;
assign v_9105 = v_8604;
assign v_9106 = ~v_8607;
assign v_9107 = ~v_560;
assign v_9108 = v_560;
assign v_9109 = ~v_8611;
assign v_9110 = ~v_564;
assign v_9111 = v_564;
assign v_9112 = ~v_8615;
assign v_9113 = ~v_568;
assign v_9114 = v_568;
assign v_9115 = ~v_8619;
assign v_9116 = ~v_572;
assign v_9117 = v_572;
assign v_9118 = ~v_8623;
assign v_9119 = ~v_576;
assign v_9120 = v_576;
assign v_9121 = ~v_8627;
assign v_9122 = ~v_580;
assign v_9123 = v_580;
assign v_9124 = ~v_8631;
assign v_9125 = ~v_584;
assign v_9126 = v_584;
assign v_9127 = ~v_8635;
assign v_9128 = ~v_588;
assign v_9129 = v_588;
assign v_9130 = ~v_8639;
assign v_9131 = ~v_592;
assign v_9132 = v_592;
assign v_9133 = ~v_8643;
assign v_9134 = ~v_596;
assign v_9135 = v_596;
assign v_9136 = ~v_8647;
assign v_9137 = ~v_600;
assign v_9138 = v_600;
assign v_9139 = ~v_8651;
assign v_9140 = ~v_604;
assign v_9141 = v_604;
assign v_9142 = ~v_8655;
assign v_9143 = ~v_608;
assign v_9144 = v_9143;
assign v_9146 = v_9145;
assign v_9148 = v_9140 & v_9147;
assign v_9150 = v_8651;
assign v_9152 = v_9149 & v_9151;
assign v_9154 = v_9137 & v_9153;
assign v_9156 = v_8647;
assign v_9158 = v_9155 & v_9157;
assign v_9160 = v_9134 & v_9159;
assign v_9162 = v_8643;
assign v_9164 = v_9161 & v_9163;
assign v_9166 = v_9131 & v_9165;
assign v_9168 = v_8639;
assign v_9170 = v_9167 & v_9169;
assign v_9172 = v_9128 & v_9171;
assign v_9174 = v_8635;
assign v_9176 = v_9173 & v_9175;
assign v_9178 = v_9125 & v_9177;
assign v_9180 = v_8631;
assign v_9182 = v_9179 & v_9181;
assign v_9184 = v_9122 & v_9183;
assign v_9186 = v_8627;
assign v_9188 = v_9185 & v_9187;
assign v_9190 = v_9119 & v_9189;
assign v_9192 = v_8623;
assign v_9194 = v_9191 & v_9193;
assign v_9196 = v_9116 & v_9195;
assign v_9198 = v_8619;
assign v_9200 = v_9197 & v_9199;
assign v_9202 = v_9113 & v_9201;
assign v_9204 = v_8615;
assign v_9206 = v_9203 & v_9205;
assign v_9208 = v_9110 & v_9207;
assign v_9210 = v_8611;
assign v_9212 = v_9209 & v_9211;
assign v_9214 = v_9107 & v_9213;
assign v_9216 = v_8607;
assign v_9218 = v_9215 & v_9217;
assign v_9220 = v_9104 & v_9219;
assign v_9222 = v_555;
assign v_9224 = v_9221 & v_9223;
assign v_9226 = v_9101 & v_9225;
assign v_9228 = v_551;
assign v_9230 = v_9227 & v_9229;
assign v_9232 = v_9098 & v_9231;
assign v_9234 = v_547;
assign v_9236 = v_9233 & v_9235;
assign v_9238 = v_9095 & v_9237;
assign v_9240 = v_543;
assign v_9242 = v_9239 & v_9241;
assign v_9243 = v_9242;
assign v_9245 = v_8655;
assign v_9246 = v_608;
assign v_9247 = v_9246;
assign v_9248 = v_9245 & v_9247;
assign v_9249 = v_9248;
assign v_9250 = v_9140 & v_9249;
assign v_9252 = v_9150 & v_9251;
assign v_9253 = v_9139 & v_9249;
assign v_9255 = v_9137 & v_9254;
assign v_9257 = v_9156 & v_9256;
assign v_9258 = v_9136 & v_9254;
assign v_9260 = v_9134 & v_9259;
assign v_9262 = v_9162 & v_9261;
assign v_9263 = v_9133 & v_9259;
assign v_9265 = v_9131 & v_9264;
assign v_9267 = v_9168 & v_9266;
assign v_9268 = v_9130 & v_9264;
assign v_9270 = v_9128 & v_9269;
assign v_9272 = v_9174 & v_9271;
assign v_9273 = v_9127 & v_9269;
assign v_9275 = v_9125 & v_9274;
assign v_9277 = v_9180 & v_9276;
assign v_9278 = v_9124 & v_9274;
assign v_9280 = v_9122 & v_9279;
assign v_9282 = v_9186 & v_9281;
assign v_9283 = v_9121 & v_9279;
assign v_9285 = v_9119 & v_9284;
assign v_9287 = v_9192 & v_9286;
assign v_9288 = v_9118 & v_9284;
assign v_9290 = v_9116 & v_9289;
assign v_9292 = v_9198 & v_9291;
assign v_9293 = v_9115 & v_9289;
assign v_9295 = v_9113 & v_9294;
assign v_9297 = v_9204 & v_9296;
assign v_9298 = v_9112 & v_9294;
assign v_9300 = v_9110 & v_9299;
assign v_9302 = v_9210 & v_9301;
assign v_9303 = v_9109 & v_9299;
assign v_9305 = v_9107 & v_9304;
assign v_9307 = v_9216 & v_9306;
assign v_9308 = v_9106 & v_9304;
assign v_9310 = v_9104 & v_9309;
assign v_9312 = v_9222 & v_9311;
assign v_9313 = v_9103 & v_9309;
assign v_9315 = v_9101 & v_9314;
assign v_9317 = v_9228 & v_9316;
assign v_9318 = v_9100 & v_9314;
assign v_9320 = v_9098 & v_9319;
assign v_9322 = v_9234 & v_9321;
assign v_9323 = v_9097 & v_9319;
assign v_9325 = v_9095 & v_9324;
assign v_9327 = v_9240 & v_9326;
assign v_9328 = v_9094 & v_9324;
assign v_9330 = v_9329;
assign v_9332 = v_9244 & v_9331;
assign v_9333 = v_9332;
assign v_9335 = v_9334;
assign v_9337 = ~v_803;
assign v_9338 = ~v_8592;
assign v_9339 = v_8592;
assign v_9340 = ~v_807;
assign v_9341 = ~v_8596;
assign v_9342 = v_8596;
assign v_9343 = ~v_811;
assign v_9344 = ~v_8600;
assign v_9345 = v_8600;
assign v_9346 = ~v_815;
assign v_9347 = ~v_8604;
assign v_9348 = v_8604;
assign v_9349 = ~v_8607;
assign v_9350 = ~v_820;
assign v_9351 = v_820;
assign v_9352 = ~v_8611;
assign v_9353 = ~v_824;
assign v_9354 = v_824;
assign v_9355 = ~v_8615;
assign v_9356 = ~v_828;
assign v_9357 = v_828;
assign v_9358 = ~v_8619;
assign v_9359 = ~v_832;
assign v_9360 = v_832;
assign v_9361 = ~v_8623;
assign v_9362 = ~v_836;
assign v_9363 = v_836;
assign v_9364 = ~v_8627;
assign v_9365 = ~v_840;
assign v_9366 = v_840;
assign v_9367 = ~v_8631;
assign v_9368 = ~v_844;
assign v_9369 = v_844;
assign v_9370 = ~v_8635;
assign v_9371 = ~v_848;
assign v_9372 = v_848;
assign v_9373 = ~v_8639;
assign v_9374 = ~v_852;
assign v_9375 = v_852;
assign v_9376 = ~v_8643;
assign v_9377 = ~v_856;
assign v_9378 = v_856;
assign v_9379 = ~v_8647;
assign v_9380 = ~v_860;
assign v_9381 = v_860;
assign v_9382 = ~v_8651;
assign v_9383 = ~v_864;
assign v_9384 = v_864;
assign v_9385 = ~v_8655;
assign v_9386 = ~v_868;
assign v_9387 = v_9386;
assign v_9389 = v_9388;
assign v_9391 = v_9383 & v_9390;
assign v_9393 = v_8651;
assign v_9395 = v_9392 & v_9394;
assign v_9397 = v_9380 & v_9396;
assign v_9399 = v_8647;
assign v_9401 = v_9398 & v_9400;
assign v_9403 = v_9377 & v_9402;
assign v_9405 = v_8643;
assign v_9407 = v_9404 & v_9406;
assign v_9409 = v_9374 & v_9408;
assign v_9411 = v_8639;
assign v_9413 = v_9410 & v_9412;
assign v_9415 = v_9371 & v_9414;
assign v_9417 = v_8635;
assign v_9419 = v_9416 & v_9418;
assign v_9421 = v_9368 & v_9420;
assign v_9423 = v_8631;
assign v_9425 = v_9422 & v_9424;
assign v_9427 = v_9365 & v_9426;
assign v_9429 = v_8627;
assign v_9431 = v_9428 & v_9430;
assign v_9433 = v_9362 & v_9432;
assign v_9435 = v_8623;
assign v_9437 = v_9434 & v_9436;
assign v_9439 = v_9359 & v_9438;
assign v_9441 = v_8619;
assign v_9443 = v_9440 & v_9442;
assign v_9445 = v_9356 & v_9444;
assign v_9447 = v_8615;
assign v_9449 = v_9446 & v_9448;
assign v_9451 = v_9353 & v_9450;
assign v_9453 = v_8611;
assign v_9455 = v_9452 & v_9454;
assign v_9457 = v_9350 & v_9456;
assign v_9459 = v_8607;
assign v_9461 = v_9458 & v_9460;
assign v_9463 = v_9347 & v_9462;
assign v_9465 = v_815;
assign v_9467 = v_9464 & v_9466;
assign v_9469 = v_9344 & v_9468;
assign v_9471 = v_811;
assign v_9473 = v_9470 & v_9472;
assign v_9475 = v_9341 & v_9474;
assign v_9477 = v_807;
assign v_9479 = v_9476 & v_9478;
assign v_9481 = v_9338 & v_9480;
assign v_9483 = v_803;
assign v_9485 = v_9482 & v_9484;
assign v_9486 = v_9485;
assign v_9488 = v_8655;
assign v_9489 = v_868;
assign v_9490 = v_9489;
assign v_9491 = v_9488 & v_9490;
assign v_9492 = v_9491;
assign v_9493 = v_9383 & v_9492;
assign v_9495 = v_9393 & v_9494;
assign v_9496 = v_9382 & v_9492;
assign v_9498 = v_9380 & v_9497;
assign v_9500 = v_9399 & v_9499;
assign v_9501 = v_9379 & v_9497;
assign v_9503 = v_9377 & v_9502;
assign v_9505 = v_9405 & v_9504;
assign v_9506 = v_9376 & v_9502;
assign v_9508 = v_9374 & v_9507;
assign v_9510 = v_9411 & v_9509;
assign v_9511 = v_9373 & v_9507;
assign v_9513 = v_9371 & v_9512;
assign v_9515 = v_9417 & v_9514;
assign v_9516 = v_9370 & v_9512;
assign v_9518 = v_9368 & v_9517;
assign v_9520 = v_9423 & v_9519;
assign v_9521 = v_9367 & v_9517;
assign v_9523 = v_9365 & v_9522;
assign v_9525 = v_9429 & v_9524;
assign v_9526 = v_9364 & v_9522;
assign v_9528 = v_9362 & v_9527;
assign v_9530 = v_9435 & v_9529;
assign v_9531 = v_9361 & v_9527;
assign v_9533 = v_9359 & v_9532;
assign v_9535 = v_9441 & v_9534;
assign v_9536 = v_9358 & v_9532;
assign v_9538 = v_9356 & v_9537;
assign v_9540 = v_9447 & v_9539;
assign v_9541 = v_9355 & v_9537;
assign v_9543 = v_9353 & v_9542;
assign v_9545 = v_9453 & v_9544;
assign v_9546 = v_9352 & v_9542;
assign v_9548 = v_9350 & v_9547;
assign v_9550 = v_9459 & v_9549;
assign v_9551 = v_9349 & v_9547;
assign v_9553 = v_9347 & v_9552;
assign v_9555 = v_9465 & v_9554;
assign v_9556 = v_9346 & v_9552;
assign v_9558 = v_9344 & v_9557;
assign v_9560 = v_9471 & v_9559;
assign v_9561 = v_9343 & v_9557;
assign v_9563 = v_9341 & v_9562;
assign v_9565 = v_9477 & v_9564;
assign v_9566 = v_9340 & v_9562;
assign v_9568 = v_9338 & v_9567;
assign v_9570 = v_9483 & v_9569;
assign v_9571 = v_9337 & v_9567;
assign v_9573 = v_9572;
assign v_9575 = v_9487 & v_9574;
assign v_9576 = v_9575;
assign v_9578 = v_9577;
assign v_9580 = ~v_1063;
assign v_9581 = ~v_8592;
assign v_9582 = v_8592;
assign v_9583 = ~v_1067;
assign v_9584 = ~v_8596;
assign v_9585 = v_8596;
assign v_9586 = ~v_1071;
assign v_9587 = ~v_8600;
assign v_9588 = v_8600;
assign v_9589 = ~v_1075;
assign v_9590 = ~v_8604;
assign v_9591 = v_8604;
assign v_9592 = ~v_8607;
assign v_9593 = ~v_1080;
assign v_9594 = v_1080;
assign v_9595 = ~v_8611;
assign v_9596 = ~v_1084;
assign v_9597 = v_1084;
assign v_9598 = ~v_8615;
assign v_9599 = ~v_1088;
assign v_9600 = v_1088;
assign v_9601 = ~v_8619;
assign v_9602 = ~v_1092;
assign v_9603 = v_1092;
assign v_9604 = ~v_8623;
assign v_9605 = ~v_1096;
assign v_9606 = v_1096;
assign v_9607 = ~v_8627;
assign v_9608 = ~v_1100;
assign v_9609 = v_1100;
assign v_9610 = ~v_8631;
assign v_9611 = ~v_1104;
assign v_9612 = v_1104;
assign v_9613 = ~v_8635;
assign v_9614 = ~v_1108;
assign v_9615 = v_1108;
assign v_9616 = ~v_8639;
assign v_9617 = ~v_1112;
assign v_9618 = v_1112;
assign v_9619 = ~v_8643;
assign v_9620 = ~v_1116;
assign v_9621 = v_1116;
assign v_9622 = ~v_8647;
assign v_9623 = ~v_1120;
assign v_9624 = v_1120;
assign v_9625 = ~v_8651;
assign v_9626 = ~v_1124;
assign v_9627 = v_1124;
assign v_9628 = ~v_8655;
assign v_9629 = ~v_1128;
assign v_9630 = v_9629;
assign v_9632 = v_9631;
assign v_9634 = v_9626 & v_9633;
assign v_9636 = v_8651;
assign v_9638 = v_9635 & v_9637;
assign v_9640 = v_9623 & v_9639;
assign v_9642 = v_8647;
assign v_9644 = v_9641 & v_9643;
assign v_9646 = v_9620 & v_9645;
assign v_9648 = v_8643;
assign v_9650 = v_9647 & v_9649;
assign v_9652 = v_9617 & v_9651;
assign v_9654 = v_8639;
assign v_9656 = v_9653 & v_9655;
assign v_9658 = v_9614 & v_9657;
assign v_9660 = v_8635;
assign v_9662 = v_9659 & v_9661;
assign v_9664 = v_9611 & v_9663;
assign v_9666 = v_8631;
assign v_9668 = v_9665 & v_9667;
assign v_9670 = v_9608 & v_9669;
assign v_9672 = v_8627;
assign v_9674 = v_9671 & v_9673;
assign v_9676 = v_9605 & v_9675;
assign v_9678 = v_8623;
assign v_9680 = v_9677 & v_9679;
assign v_9682 = v_9602 & v_9681;
assign v_9684 = v_8619;
assign v_9686 = v_9683 & v_9685;
assign v_9688 = v_9599 & v_9687;
assign v_9690 = v_8615;
assign v_9692 = v_9689 & v_9691;
assign v_9694 = v_9596 & v_9693;
assign v_9696 = v_8611;
assign v_9698 = v_9695 & v_9697;
assign v_9700 = v_9593 & v_9699;
assign v_9702 = v_8607;
assign v_9704 = v_9701 & v_9703;
assign v_9706 = v_9590 & v_9705;
assign v_9708 = v_1075;
assign v_9710 = v_9707 & v_9709;
assign v_9712 = v_9587 & v_9711;
assign v_9714 = v_1071;
assign v_9716 = v_9713 & v_9715;
assign v_9718 = v_9584 & v_9717;
assign v_9720 = v_1067;
assign v_9722 = v_9719 & v_9721;
assign v_9724 = v_9581 & v_9723;
assign v_9726 = v_1063;
assign v_9728 = v_9725 & v_9727;
assign v_9729 = v_9728;
assign v_9731 = v_8655;
assign v_9732 = v_1128;
assign v_9733 = v_9732;
assign v_9734 = v_9731 & v_9733;
assign v_9735 = v_9734;
assign v_9736 = v_9626 & v_9735;
assign v_9738 = v_9636 & v_9737;
assign v_9739 = v_9625 & v_9735;
assign v_9741 = v_9623 & v_9740;
assign v_9743 = v_9642 & v_9742;
assign v_9744 = v_9622 & v_9740;
assign v_9746 = v_9620 & v_9745;
assign v_9748 = v_9648 & v_9747;
assign v_9749 = v_9619 & v_9745;
assign v_9751 = v_9617 & v_9750;
assign v_9753 = v_9654 & v_9752;
assign v_9754 = v_9616 & v_9750;
assign v_9756 = v_9614 & v_9755;
assign v_9758 = v_9660 & v_9757;
assign v_9759 = v_9613 & v_9755;
assign v_9761 = v_9611 & v_9760;
assign v_9763 = v_9666 & v_9762;
assign v_9764 = v_9610 & v_9760;
assign v_9766 = v_9608 & v_9765;
assign v_9768 = v_9672 & v_9767;
assign v_9769 = v_9607 & v_9765;
assign v_9771 = v_9605 & v_9770;
assign v_9773 = v_9678 & v_9772;
assign v_9774 = v_9604 & v_9770;
assign v_9776 = v_9602 & v_9775;
assign v_9778 = v_9684 & v_9777;
assign v_9779 = v_9601 & v_9775;
assign v_9781 = v_9599 & v_9780;
assign v_9783 = v_9690 & v_9782;
assign v_9784 = v_9598 & v_9780;
assign v_9786 = v_9596 & v_9785;
assign v_9788 = v_9696 & v_9787;
assign v_9789 = v_9595 & v_9785;
assign v_9791 = v_9593 & v_9790;
assign v_9793 = v_9702 & v_9792;
assign v_9794 = v_9592 & v_9790;
assign v_9796 = v_9590 & v_9795;
assign v_9798 = v_9708 & v_9797;
assign v_9799 = v_9589 & v_9795;
assign v_9801 = v_9587 & v_9800;
assign v_9803 = v_9714 & v_9802;
assign v_9804 = v_9586 & v_9800;
assign v_9806 = v_9584 & v_9805;
assign v_9808 = v_9720 & v_9807;
assign v_9809 = v_9583 & v_9805;
assign v_9811 = v_9581 & v_9810;
assign v_9813 = v_9726 & v_9812;
assign v_9814 = v_9580 & v_9810;
assign v_9816 = v_9815;
assign v_9818 = v_9730 & v_9817;
assign v_9819 = v_9818;
assign v_9821 = v_9820;
assign v_9823 = ~v_1323;
assign v_9824 = ~v_8592;
assign v_9825 = v_8592;
assign v_9826 = ~v_1327;
assign v_9827 = ~v_8596;
assign v_9828 = v_8596;
assign v_9829 = ~v_1331;
assign v_9830 = ~v_8600;
assign v_9831 = v_8600;
assign v_9832 = ~v_1335;
assign v_9833 = ~v_8604;
assign v_9834 = v_8604;
assign v_9835 = ~v_8607;
assign v_9836 = ~v_1340;
assign v_9837 = v_1340;
assign v_9838 = ~v_8611;
assign v_9839 = ~v_1344;
assign v_9840 = v_1344;
assign v_9841 = ~v_8615;
assign v_9842 = ~v_1348;
assign v_9843 = v_1348;
assign v_9844 = ~v_8619;
assign v_9845 = ~v_1352;
assign v_9846 = v_1352;
assign v_9847 = ~v_8623;
assign v_9848 = ~v_1356;
assign v_9849 = v_1356;
assign v_9850 = ~v_8627;
assign v_9851 = ~v_1360;
assign v_9852 = v_1360;
assign v_9853 = ~v_8631;
assign v_9854 = ~v_1364;
assign v_9855 = v_1364;
assign v_9856 = ~v_8635;
assign v_9857 = ~v_1368;
assign v_9858 = v_1368;
assign v_9859 = ~v_8639;
assign v_9860 = ~v_1372;
assign v_9861 = v_1372;
assign v_9862 = ~v_8643;
assign v_9863 = ~v_1376;
assign v_9864 = v_1376;
assign v_9865 = ~v_8647;
assign v_9866 = ~v_1380;
assign v_9867 = v_1380;
assign v_9868 = ~v_8651;
assign v_9869 = ~v_1384;
assign v_9870 = v_1384;
assign v_9871 = ~v_8655;
assign v_9872 = ~v_1388;
assign v_9873 = v_9872;
assign v_9875 = v_9874;
assign v_9877 = v_9869 & v_9876;
assign v_9879 = v_8651;
assign v_9881 = v_9878 & v_9880;
assign v_9883 = v_9866 & v_9882;
assign v_9885 = v_8647;
assign v_9887 = v_9884 & v_9886;
assign v_9889 = v_9863 & v_9888;
assign v_9891 = v_8643;
assign v_9893 = v_9890 & v_9892;
assign v_9895 = v_9860 & v_9894;
assign v_9897 = v_8639;
assign v_9899 = v_9896 & v_9898;
assign v_9901 = v_9857 & v_9900;
assign v_9903 = v_8635;
assign v_9905 = v_9902 & v_9904;
assign v_9907 = v_9854 & v_9906;
assign v_9909 = v_8631;
assign v_9911 = v_9908 & v_9910;
assign v_9913 = v_9851 & v_9912;
assign v_9915 = v_8627;
assign v_9917 = v_9914 & v_9916;
assign v_9919 = v_9848 & v_9918;
assign v_9921 = v_8623;
assign v_9923 = v_9920 & v_9922;
assign v_9925 = v_9845 & v_9924;
assign v_9927 = v_8619;
assign v_9929 = v_9926 & v_9928;
assign v_9931 = v_9842 & v_9930;
assign v_9933 = v_8615;
assign v_9935 = v_9932 & v_9934;
assign v_9937 = v_9839 & v_9936;
assign v_9939 = v_8611;
assign v_9941 = v_9938 & v_9940;
assign v_9943 = v_9836 & v_9942;
assign v_9945 = v_8607;
assign v_9947 = v_9944 & v_9946;
assign v_9949 = v_9833 & v_9948;
assign v_9951 = v_1335;
assign v_9953 = v_9950 & v_9952;
assign v_9955 = v_9830 & v_9954;
assign v_9957 = v_1331;
assign v_9959 = v_9956 & v_9958;
assign v_9961 = v_9827 & v_9960;
assign v_9963 = v_1327;
assign v_9965 = v_9962 & v_9964;
assign v_9967 = v_9824 & v_9966;
assign v_9969 = v_1323;
assign v_9971 = v_9968 & v_9970;
assign v_9972 = v_9971;
assign v_9974 = v_8655;
assign v_9975 = v_1388;
assign v_9976 = v_9975;
assign v_9977 = v_9974 & v_9976;
assign v_9978 = v_9977;
assign v_9979 = v_9869 & v_9978;
assign v_9981 = v_9879 & v_9980;
assign v_9982 = v_9868 & v_9978;
assign v_9984 = v_9866 & v_9983;
assign v_9986 = v_9885 & v_9985;
assign v_9987 = v_9865 & v_9983;
assign v_9989 = v_9863 & v_9988;
assign v_9991 = v_9891 & v_9990;
assign v_9992 = v_9862 & v_9988;
assign v_9994 = v_9860 & v_9993;
assign v_9996 = v_9897 & v_9995;
assign v_9997 = v_9859 & v_9993;
assign v_9999 = v_9857 & v_9998;
assign v_10001 = v_9903 & v_10000;
assign v_10002 = v_9856 & v_9998;
assign v_10004 = v_9854 & v_10003;
assign v_10006 = v_9909 & v_10005;
assign v_10007 = v_9853 & v_10003;
assign v_10009 = v_9851 & v_10008;
assign v_10011 = v_9915 & v_10010;
assign v_10012 = v_9850 & v_10008;
assign v_10014 = v_9848 & v_10013;
assign v_10016 = v_9921 & v_10015;
assign v_10017 = v_9847 & v_10013;
assign v_10019 = v_9845 & v_10018;
assign v_10021 = v_9927 & v_10020;
assign v_10022 = v_9844 & v_10018;
assign v_10024 = v_9842 & v_10023;
assign v_10026 = v_9933 & v_10025;
assign v_10027 = v_9841 & v_10023;
assign v_10029 = v_9839 & v_10028;
assign v_10031 = v_9939 & v_10030;
assign v_10032 = v_9838 & v_10028;
assign v_10034 = v_9836 & v_10033;
assign v_10036 = v_9945 & v_10035;
assign v_10037 = v_9835 & v_10033;
assign v_10039 = v_9833 & v_10038;
assign v_10041 = v_9951 & v_10040;
assign v_10042 = v_9832 & v_10038;
assign v_10044 = v_9830 & v_10043;
assign v_10046 = v_9957 & v_10045;
assign v_10047 = v_9829 & v_10043;
assign v_10049 = v_9827 & v_10048;
assign v_10051 = v_9963 & v_10050;
assign v_10052 = v_9826 & v_10048;
assign v_10054 = v_9824 & v_10053;
assign v_10056 = v_9969 & v_10055;
assign v_10057 = v_9823 & v_10053;
assign v_10059 = v_10058;
assign v_10061 = v_9973 & v_10060;
assign v_10062 = v_10061;
assign v_10064 = v_10063;
assign v_10066 = ~v_1583;
assign v_10067 = ~v_8592;
assign v_10068 = v_8592;
assign v_10069 = ~v_1587;
assign v_10070 = ~v_8596;
assign v_10071 = v_8596;
assign v_10072 = ~v_1591;
assign v_10073 = ~v_8600;
assign v_10074 = v_8600;
assign v_10075 = ~v_1595;
assign v_10076 = ~v_8604;
assign v_10077 = v_8604;
assign v_10078 = ~v_8607;
assign v_10079 = ~v_1600;
assign v_10080 = v_1600;
assign v_10081 = ~v_8611;
assign v_10082 = ~v_1604;
assign v_10083 = v_1604;
assign v_10084 = ~v_8615;
assign v_10085 = ~v_1608;
assign v_10086 = v_1608;
assign v_10087 = ~v_8619;
assign v_10088 = ~v_1612;
assign v_10089 = v_1612;
assign v_10090 = ~v_8623;
assign v_10091 = ~v_1616;
assign v_10092 = v_1616;
assign v_10093 = ~v_8627;
assign v_10094 = ~v_1620;
assign v_10095 = v_1620;
assign v_10096 = ~v_8631;
assign v_10097 = ~v_1624;
assign v_10098 = v_1624;
assign v_10099 = ~v_8635;
assign v_10100 = ~v_1628;
assign v_10101 = v_1628;
assign v_10102 = ~v_8639;
assign v_10103 = ~v_1632;
assign v_10104 = v_1632;
assign v_10105 = ~v_8643;
assign v_10106 = ~v_1636;
assign v_10107 = v_1636;
assign v_10108 = ~v_8647;
assign v_10109 = ~v_1640;
assign v_10110 = v_1640;
assign v_10111 = ~v_8651;
assign v_10112 = ~v_1644;
assign v_10113 = v_1644;
assign v_10114 = ~v_8655;
assign v_10115 = ~v_1648;
assign v_10116 = v_10115;
assign v_10118 = v_10117;
assign v_10120 = v_10112 & v_10119;
assign v_10122 = v_8651;
assign v_10124 = v_10121 & v_10123;
assign v_10126 = v_10109 & v_10125;
assign v_10128 = v_8647;
assign v_10130 = v_10127 & v_10129;
assign v_10132 = v_10106 & v_10131;
assign v_10134 = v_8643;
assign v_10136 = v_10133 & v_10135;
assign v_10138 = v_10103 & v_10137;
assign v_10140 = v_8639;
assign v_10142 = v_10139 & v_10141;
assign v_10144 = v_10100 & v_10143;
assign v_10146 = v_8635;
assign v_10148 = v_10145 & v_10147;
assign v_10150 = v_10097 & v_10149;
assign v_10152 = v_8631;
assign v_10154 = v_10151 & v_10153;
assign v_10156 = v_10094 & v_10155;
assign v_10158 = v_8627;
assign v_10160 = v_10157 & v_10159;
assign v_10162 = v_10091 & v_10161;
assign v_10164 = v_8623;
assign v_10166 = v_10163 & v_10165;
assign v_10168 = v_10088 & v_10167;
assign v_10170 = v_8619;
assign v_10172 = v_10169 & v_10171;
assign v_10174 = v_10085 & v_10173;
assign v_10176 = v_8615;
assign v_10178 = v_10175 & v_10177;
assign v_10180 = v_10082 & v_10179;
assign v_10182 = v_8611;
assign v_10184 = v_10181 & v_10183;
assign v_10186 = v_10079 & v_10185;
assign v_10188 = v_8607;
assign v_10190 = v_10187 & v_10189;
assign v_10192 = v_10076 & v_10191;
assign v_10194 = v_1595;
assign v_10196 = v_10193 & v_10195;
assign v_10198 = v_10073 & v_10197;
assign v_10200 = v_1591;
assign v_10202 = v_10199 & v_10201;
assign v_10204 = v_10070 & v_10203;
assign v_10206 = v_1587;
assign v_10208 = v_10205 & v_10207;
assign v_10210 = v_10067 & v_10209;
assign v_10212 = v_1583;
assign v_10214 = v_10211 & v_10213;
assign v_10215 = v_10214;
assign v_10217 = v_8655;
assign v_10218 = v_1648;
assign v_10219 = v_10218;
assign v_10220 = v_10217 & v_10219;
assign v_10221 = v_10220;
assign v_10222 = v_10112 & v_10221;
assign v_10224 = v_10122 & v_10223;
assign v_10225 = v_10111 & v_10221;
assign v_10227 = v_10109 & v_10226;
assign v_10229 = v_10128 & v_10228;
assign v_10230 = v_10108 & v_10226;
assign v_10232 = v_10106 & v_10231;
assign v_10234 = v_10134 & v_10233;
assign v_10235 = v_10105 & v_10231;
assign v_10237 = v_10103 & v_10236;
assign v_10239 = v_10140 & v_10238;
assign v_10240 = v_10102 & v_10236;
assign v_10242 = v_10100 & v_10241;
assign v_10244 = v_10146 & v_10243;
assign v_10245 = v_10099 & v_10241;
assign v_10247 = v_10097 & v_10246;
assign v_10249 = v_10152 & v_10248;
assign v_10250 = v_10096 & v_10246;
assign v_10252 = v_10094 & v_10251;
assign v_10254 = v_10158 & v_10253;
assign v_10255 = v_10093 & v_10251;
assign v_10257 = v_10091 & v_10256;
assign v_10259 = v_10164 & v_10258;
assign v_10260 = v_10090 & v_10256;
assign v_10262 = v_10088 & v_10261;
assign v_10264 = v_10170 & v_10263;
assign v_10265 = v_10087 & v_10261;
assign v_10267 = v_10085 & v_10266;
assign v_10269 = v_10176 & v_10268;
assign v_10270 = v_10084 & v_10266;
assign v_10272 = v_10082 & v_10271;
assign v_10274 = v_10182 & v_10273;
assign v_10275 = v_10081 & v_10271;
assign v_10277 = v_10079 & v_10276;
assign v_10279 = v_10188 & v_10278;
assign v_10280 = v_10078 & v_10276;
assign v_10282 = v_10076 & v_10281;
assign v_10284 = v_10194 & v_10283;
assign v_10285 = v_10075 & v_10281;
assign v_10287 = v_10073 & v_10286;
assign v_10289 = v_10200 & v_10288;
assign v_10290 = v_10072 & v_10286;
assign v_10292 = v_10070 & v_10291;
assign v_10294 = v_10206 & v_10293;
assign v_10295 = v_10069 & v_10291;
assign v_10297 = v_10067 & v_10296;
assign v_10299 = v_10212 & v_10298;
assign v_10300 = v_10066 & v_10296;
assign v_10302 = v_10301;
assign v_10304 = v_10216 & v_10303;
assign v_10305 = v_10304;
assign v_10307 = v_10306;
assign v_10309 = ~v_1843;
assign v_10310 = ~v_8592;
assign v_10311 = v_8592;
assign v_10312 = ~v_1847;
assign v_10313 = ~v_8596;
assign v_10314 = v_8596;
assign v_10315 = ~v_1851;
assign v_10316 = ~v_8600;
assign v_10317 = v_8600;
assign v_10318 = ~v_1855;
assign v_10319 = ~v_8604;
assign v_10320 = v_8604;
assign v_10321 = ~v_8607;
assign v_10322 = ~v_1860;
assign v_10323 = v_1860;
assign v_10324 = ~v_8611;
assign v_10325 = ~v_1864;
assign v_10326 = v_1864;
assign v_10327 = ~v_8615;
assign v_10328 = ~v_1868;
assign v_10329 = v_1868;
assign v_10330 = ~v_8619;
assign v_10331 = ~v_1872;
assign v_10332 = v_1872;
assign v_10333 = ~v_8623;
assign v_10334 = ~v_1876;
assign v_10335 = v_1876;
assign v_10336 = ~v_8627;
assign v_10337 = ~v_1880;
assign v_10338 = v_1880;
assign v_10339 = ~v_8631;
assign v_10340 = ~v_1884;
assign v_10341 = v_1884;
assign v_10342 = ~v_8635;
assign v_10343 = ~v_1888;
assign v_10344 = v_1888;
assign v_10345 = ~v_8639;
assign v_10346 = ~v_1892;
assign v_10347 = v_1892;
assign v_10348 = ~v_8643;
assign v_10349 = ~v_1896;
assign v_10350 = v_1896;
assign v_10351 = ~v_8647;
assign v_10352 = ~v_1900;
assign v_10353 = v_1900;
assign v_10354 = ~v_8651;
assign v_10355 = ~v_1904;
assign v_10356 = v_1904;
assign v_10357 = ~v_8655;
assign v_10358 = ~v_1908;
assign v_10359 = v_10358;
assign v_10361 = v_10360;
assign v_10363 = v_10355 & v_10362;
assign v_10365 = v_8651;
assign v_10367 = v_10364 & v_10366;
assign v_10369 = v_10352 & v_10368;
assign v_10371 = v_8647;
assign v_10373 = v_10370 & v_10372;
assign v_10375 = v_10349 & v_10374;
assign v_10377 = v_8643;
assign v_10379 = v_10376 & v_10378;
assign v_10381 = v_10346 & v_10380;
assign v_10383 = v_8639;
assign v_10385 = v_10382 & v_10384;
assign v_10387 = v_10343 & v_10386;
assign v_10389 = v_8635;
assign v_10391 = v_10388 & v_10390;
assign v_10393 = v_10340 & v_10392;
assign v_10395 = v_8631;
assign v_10397 = v_10394 & v_10396;
assign v_10399 = v_10337 & v_10398;
assign v_10401 = v_8627;
assign v_10403 = v_10400 & v_10402;
assign v_10405 = v_10334 & v_10404;
assign v_10407 = v_8623;
assign v_10409 = v_10406 & v_10408;
assign v_10411 = v_10331 & v_10410;
assign v_10413 = v_8619;
assign v_10415 = v_10412 & v_10414;
assign v_10417 = v_10328 & v_10416;
assign v_10419 = v_8615;
assign v_10421 = v_10418 & v_10420;
assign v_10423 = v_10325 & v_10422;
assign v_10425 = v_8611;
assign v_10427 = v_10424 & v_10426;
assign v_10429 = v_10322 & v_10428;
assign v_10431 = v_8607;
assign v_10433 = v_10430 & v_10432;
assign v_10435 = v_10319 & v_10434;
assign v_10437 = v_1855;
assign v_10439 = v_10436 & v_10438;
assign v_10441 = v_10316 & v_10440;
assign v_10443 = v_1851;
assign v_10445 = v_10442 & v_10444;
assign v_10447 = v_10313 & v_10446;
assign v_10449 = v_1847;
assign v_10451 = v_10448 & v_10450;
assign v_10453 = v_10310 & v_10452;
assign v_10455 = v_1843;
assign v_10457 = v_10454 & v_10456;
assign v_10458 = v_10457;
assign v_10460 = v_8655;
assign v_10461 = v_1908;
assign v_10462 = v_10461;
assign v_10463 = v_10460 & v_10462;
assign v_10464 = v_10463;
assign v_10465 = v_10355 & v_10464;
assign v_10467 = v_10365 & v_10466;
assign v_10468 = v_10354 & v_10464;
assign v_10470 = v_10352 & v_10469;
assign v_10472 = v_10371 & v_10471;
assign v_10473 = v_10351 & v_10469;
assign v_10475 = v_10349 & v_10474;
assign v_10477 = v_10377 & v_10476;
assign v_10478 = v_10348 & v_10474;
assign v_10480 = v_10346 & v_10479;
assign v_10482 = v_10383 & v_10481;
assign v_10483 = v_10345 & v_10479;
assign v_10485 = v_10343 & v_10484;
assign v_10487 = v_10389 & v_10486;
assign v_10488 = v_10342 & v_10484;
assign v_10490 = v_10340 & v_10489;
assign v_10492 = v_10395 & v_10491;
assign v_10493 = v_10339 & v_10489;
assign v_10495 = v_10337 & v_10494;
assign v_10497 = v_10401 & v_10496;
assign v_10498 = v_10336 & v_10494;
assign v_10500 = v_10334 & v_10499;
assign v_10502 = v_10407 & v_10501;
assign v_10503 = v_10333 & v_10499;
assign v_10505 = v_10331 & v_10504;
assign v_10507 = v_10413 & v_10506;
assign v_10508 = v_10330 & v_10504;
assign v_10510 = v_10328 & v_10509;
assign v_10512 = v_10419 & v_10511;
assign v_10513 = v_10327 & v_10509;
assign v_10515 = v_10325 & v_10514;
assign v_10517 = v_10425 & v_10516;
assign v_10518 = v_10324 & v_10514;
assign v_10520 = v_10322 & v_10519;
assign v_10522 = v_10431 & v_10521;
assign v_10523 = v_10321 & v_10519;
assign v_10525 = v_10319 & v_10524;
assign v_10527 = v_10437 & v_10526;
assign v_10528 = v_10318 & v_10524;
assign v_10530 = v_10316 & v_10529;
assign v_10532 = v_10443 & v_10531;
assign v_10533 = v_10315 & v_10529;
assign v_10535 = v_10313 & v_10534;
assign v_10537 = v_10449 & v_10536;
assign v_10538 = v_10312 & v_10534;
assign v_10540 = v_10310 & v_10539;
assign v_10542 = v_10455 & v_10541;
assign v_10543 = v_10309 & v_10539;
assign v_10545 = v_10544;
assign v_10547 = v_10459 & v_10546;
assign v_10548 = v_10547;
assign v_10550 = v_10549;
assign v_10552 = ~v_2103;
assign v_10553 = ~v_8592;
assign v_10554 = v_8592;
assign v_10555 = ~v_2107;
assign v_10556 = ~v_8596;
assign v_10557 = v_8596;
assign v_10558 = ~v_2111;
assign v_10559 = ~v_8600;
assign v_10560 = v_8600;
assign v_10561 = ~v_2115;
assign v_10562 = ~v_8604;
assign v_10563 = v_8604;
assign v_10564 = ~v_8607;
assign v_10565 = ~v_2120;
assign v_10566 = v_2120;
assign v_10567 = ~v_8611;
assign v_10568 = ~v_2124;
assign v_10569 = v_2124;
assign v_10570 = ~v_8615;
assign v_10571 = ~v_2128;
assign v_10572 = v_2128;
assign v_10573 = ~v_8619;
assign v_10574 = ~v_2132;
assign v_10575 = v_2132;
assign v_10576 = ~v_8623;
assign v_10577 = ~v_2136;
assign v_10578 = v_2136;
assign v_10579 = ~v_8627;
assign v_10580 = ~v_2140;
assign v_10581 = v_2140;
assign v_10582 = ~v_8631;
assign v_10583 = ~v_2144;
assign v_10584 = v_2144;
assign v_10585 = ~v_8635;
assign v_10586 = ~v_2148;
assign v_10587 = v_2148;
assign v_10588 = ~v_8639;
assign v_10589 = ~v_2152;
assign v_10590 = v_2152;
assign v_10591 = ~v_8643;
assign v_10592 = ~v_2156;
assign v_10593 = v_2156;
assign v_10594 = ~v_8647;
assign v_10595 = ~v_2160;
assign v_10596 = v_2160;
assign v_10597 = ~v_8651;
assign v_10598 = ~v_2164;
assign v_10599 = v_2164;
assign v_10600 = ~v_8655;
assign v_10601 = ~v_2168;
assign v_10602 = v_10601;
assign v_10604 = v_10603;
assign v_10606 = v_10598 & v_10605;
assign v_10608 = v_8651;
assign v_10610 = v_10607 & v_10609;
assign v_10612 = v_10595 & v_10611;
assign v_10614 = v_8647;
assign v_10616 = v_10613 & v_10615;
assign v_10618 = v_10592 & v_10617;
assign v_10620 = v_8643;
assign v_10622 = v_10619 & v_10621;
assign v_10624 = v_10589 & v_10623;
assign v_10626 = v_8639;
assign v_10628 = v_10625 & v_10627;
assign v_10630 = v_10586 & v_10629;
assign v_10632 = v_8635;
assign v_10634 = v_10631 & v_10633;
assign v_10636 = v_10583 & v_10635;
assign v_10638 = v_8631;
assign v_10640 = v_10637 & v_10639;
assign v_10642 = v_10580 & v_10641;
assign v_10644 = v_8627;
assign v_10646 = v_10643 & v_10645;
assign v_10648 = v_10577 & v_10647;
assign v_10650 = v_8623;
assign v_10652 = v_10649 & v_10651;
assign v_10654 = v_10574 & v_10653;
assign v_10656 = v_8619;
assign v_10658 = v_10655 & v_10657;
assign v_10660 = v_10571 & v_10659;
assign v_10662 = v_8615;
assign v_10664 = v_10661 & v_10663;
assign v_10666 = v_10568 & v_10665;
assign v_10668 = v_8611;
assign v_10670 = v_10667 & v_10669;
assign v_10672 = v_10565 & v_10671;
assign v_10674 = v_8607;
assign v_10676 = v_10673 & v_10675;
assign v_10678 = v_10562 & v_10677;
assign v_10680 = v_2115;
assign v_10682 = v_10679 & v_10681;
assign v_10684 = v_10559 & v_10683;
assign v_10686 = v_2111;
assign v_10688 = v_10685 & v_10687;
assign v_10690 = v_10556 & v_10689;
assign v_10692 = v_2107;
assign v_10694 = v_10691 & v_10693;
assign v_10696 = v_10553 & v_10695;
assign v_10698 = v_2103;
assign v_10700 = v_10697 & v_10699;
assign v_10701 = v_10700;
assign v_10703 = v_8655;
assign v_10704 = v_2168;
assign v_10705 = v_10704;
assign v_10706 = v_10703 & v_10705;
assign v_10707 = v_10706;
assign v_10708 = v_10598 & v_10707;
assign v_10710 = v_10608 & v_10709;
assign v_10711 = v_10597 & v_10707;
assign v_10713 = v_10595 & v_10712;
assign v_10715 = v_10614 & v_10714;
assign v_10716 = v_10594 & v_10712;
assign v_10718 = v_10592 & v_10717;
assign v_10720 = v_10620 & v_10719;
assign v_10721 = v_10591 & v_10717;
assign v_10723 = v_10589 & v_10722;
assign v_10725 = v_10626 & v_10724;
assign v_10726 = v_10588 & v_10722;
assign v_10728 = v_10586 & v_10727;
assign v_10730 = v_10632 & v_10729;
assign v_10731 = v_10585 & v_10727;
assign v_10733 = v_10583 & v_10732;
assign v_10735 = v_10638 & v_10734;
assign v_10736 = v_10582 & v_10732;
assign v_10738 = v_10580 & v_10737;
assign v_10740 = v_10644 & v_10739;
assign v_10741 = v_10579 & v_10737;
assign v_10743 = v_10577 & v_10742;
assign v_10745 = v_10650 & v_10744;
assign v_10746 = v_10576 & v_10742;
assign v_10748 = v_10574 & v_10747;
assign v_10750 = v_10656 & v_10749;
assign v_10751 = v_10573 & v_10747;
assign v_10753 = v_10571 & v_10752;
assign v_10755 = v_10662 & v_10754;
assign v_10756 = v_10570 & v_10752;
assign v_10758 = v_10568 & v_10757;
assign v_10760 = v_10668 & v_10759;
assign v_10761 = v_10567 & v_10757;
assign v_10763 = v_10565 & v_10762;
assign v_10765 = v_10674 & v_10764;
assign v_10766 = v_10564 & v_10762;
assign v_10768 = v_10562 & v_10767;
assign v_10770 = v_10680 & v_10769;
assign v_10771 = v_10561 & v_10767;
assign v_10773 = v_10559 & v_10772;
assign v_10775 = v_10686 & v_10774;
assign v_10776 = v_10558 & v_10772;
assign v_10778 = v_10556 & v_10777;
assign v_10780 = v_10692 & v_10779;
assign v_10781 = v_10555 & v_10777;
assign v_10783 = v_10553 & v_10782;
assign v_10785 = v_10698 & v_10784;
assign v_10786 = v_10552 & v_10782;
assign v_10788 = v_10787;
assign v_10790 = v_10702 & v_10789;
assign v_10791 = v_10790;
assign v_10793 = v_10792;
assign v_10795 = ~v_2363;
assign v_10796 = ~v_8592;
assign v_10797 = v_8592;
assign v_10798 = ~v_2367;
assign v_10799 = ~v_8596;
assign v_10800 = v_8596;
assign v_10801 = ~v_2371;
assign v_10802 = ~v_8600;
assign v_10803 = v_8600;
assign v_10804 = ~v_2375;
assign v_10805 = ~v_8604;
assign v_10806 = v_8604;
assign v_10807 = ~v_8607;
assign v_10808 = ~v_2380;
assign v_10809 = v_2380;
assign v_10810 = ~v_8611;
assign v_10811 = ~v_2384;
assign v_10812 = v_2384;
assign v_10813 = ~v_8615;
assign v_10814 = ~v_2388;
assign v_10815 = v_2388;
assign v_10816 = ~v_8619;
assign v_10817 = ~v_2392;
assign v_10818 = v_2392;
assign v_10819 = ~v_8623;
assign v_10820 = ~v_2396;
assign v_10821 = v_2396;
assign v_10822 = ~v_8627;
assign v_10823 = ~v_2400;
assign v_10824 = v_2400;
assign v_10825 = ~v_8631;
assign v_10826 = ~v_2404;
assign v_10827 = v_2404;
assign v_10828 = ~v_8635;
assign v_10829 = ~v_2408;
assign v_10830 = v_2408;
assign v_10831 = ~v_8639;
assign v_10832 = ~v_2412;
assign v_10833 = v_2412;
assign v_10834 = ~v_8643;
assign v_10835 = ~v_2416;
assign v_10836 = v_2416;
assign v_10837 = ~v_8647;
assign v_10838 = ~v_2420;
assign v_10839 = v_2420;
assign v_10840 = ~v_8651;
assign v_10841 = ~v_2424;
assign v_10842 = v_2424;
assign v_10843 = ~v_8655;
assign v_10844 = ~v_2428;
assign v_10845 = v_10844;
assign v_10847 = v_10846;
assign v_10849 = v_10841 & v_10848;
assign v_10851 = v_8651;
assign v_10853 = v_10850 & v_10852;
assign v_10855 = v_10838 & v_10854;
assign v_10857 = v_8647;
assign v_10859 = v_10856 & v_10858;
assign v_10861 = v_10835 & v_10860;
assign v_10863 = v_8643;
assign v_10865 = v_10862 & v_10864;
assign v_10867 = v_10832 & v_10866;
assign v_10869 = v_8639;
assign v_10871 = v_10868 & v_10870;
assign v_10873 = v_10829 & v_10872;
assign v_10875 = v_8635;
assign v_10877 = v_10874 & v_10876;
assign v_10879 = v_10826 & v_10878;
assign v_10881 = v_8631;
assign v_10883 = v_10880 & v_10882;
assign v_10885 = v_10823 & v_10884;
assign v_10887 = v_8627;
assign v_10889 = v_10886 & v_10888;
assign v_10891 = v_10820 & v_10890;
assign v_10893 = v_8623;
assign v_10895 = v_10892 & v_10894;
assign v_10897 = v_10817 & v_10896;
assign v_10899 = v_8619;
assign v_10901 = v_10898 & v_10900;
assign v_10903 = v_10814 & v_10902;
assign v_10905 = v_8615;
assign v_10907 = v_10904 & v_10906;
assign v_10909 = v_10811 & v_10908;
assign v_10911 = v_8611;
assign v_10913 = v_10910 & v_10912;
assign v_10915 = v_10808 & v_10914;
assign v_10917 = v_8607;
assign v_10919 = v_10916 & v_10918;
assign v_10921 = v_10805 & v_10920;
assign v_10923 = v_2375;
assign v_10925 = v_10922 & v_10924;
assign v_10927 = v_10802 & v_10926;
assign v_10929 = v_2371;
assign v_10931 = v_10928 & v_10930;
assign v_10933 = v_10799 & v_10932;
assign v_10935 = v_2367;
assign v_10937 = v_10934 & v_10936;
assign v_10939 = v_10796 & v_10938;
assign v_10941 = v_2363;
assign v_10943 = v_10940 & v_10942;
assign v_10944 = v_10943;
assign v_10946 = v_8655;
assign v_10947 = v_2428;
assign v_10948 = v_10947;
assign v_10949 = v_10946 & v_10948;
assign v_10950 = v_10949;
assign v_10951 = v_10841 & v_10950;
assign v_10953 = v_10851 & v_10952;
assign v_10954 = v_10840 & v_10950;
assign v_10956 = v_10838 & v_10955;
assign v_10958 = v_10857 & v_10957;
assign v_10959 = v_10837 & v_10955;
assign v_10961 = v_10835 & v_10960;
assign v_10963 = v_10863 & v_10962;
assign v_10964 = v_10834 & v_10960;
assign v_10966 = v_10832 & v_10965;
assign v_10968 = v_10869 & v_10967;
assign v_10969 = v_10831 & v_10965;
assign v_10971 = v_10829 & v_10970;
assign v_10973 = v_10875 & v_10972;
assign v_10974 = v_10828 & v_10970;
assign v_10976 = v_10826 & v_10975;
assign v_10978 = v_10881 & v_10977;
assign v_10979 = v_10825 & v_10975;
assign v_10981 = v_10823 & v_10980;
assign v_10983 = v_10887 & v_10982;
assign v_10984 = v_10822 & v_10980;
assign v_10986 = v_10820 & v_10985;
assign v_10988 = v_10893 & v_10987;
assign v_10989 = v_10819 & v_10985;
assign v_10991 = v_10817 & v_10990;
assign v_10993 = v_10899 & v_10992;
assign v_10994 = v_10816 & v_10990;
assign v_10996 = v_10814 & v_10995;
assign v_10998 = v_10905 & v_10997;
assign v_10999 = v_10813 & v_10995;
assign v_11001 = v_10811 & v_11000;
assign v_11003 = v_10911 & v_11002;
assign v_11004 = v_10810 & v_11000;
assign v_11006 = v_10808 & v_11005;
assign v_11008 = v_10917 & v_11007;
assign v_11009 = v_10807 & v_11005;
assign v_11011 = v_10805 & v_11010;
assign v_11013 = v_10923 & v_11012;
assign v_11014 = v_10804 & v_11010;
assign v_11016 = v_10802 & v_11015;
assign v_11018 = v_10929 & v_11017;
assign v_11019 = v_10801 & v_11015;
assign v_11021 = v_10799 & v_11020;
assign v_11023 = v_10935 & v_11022;
assign v_11024 = v_10798 & v_11020;
assign v_11026 = v_10796 & v_11025;
assign v_11028 = v_10941 & v_11027;
assign v_11029 = v_10795 & v_11025;
assign v_11031 = v_11030;
assign v_11033 = v_10945 & v_11032;
assign v_11034 = v_11033;
assign v_11036 = v_11035;
assign v_11038 = ~v_2623;
assign v_11039 = ~v_8592;
assign v_11040 = v_8592;
assign v_11041 = ~v_2627;
assign v_11042 = ~v_8596;
assign v_11043 = v_8596;
assign v_11044 = ~v_2631;
assign v_11045 = ~v_8600;
assign v_11046 = v_8600;
assign v_11047 = ~v_2635;
assign v_11048 = ~v_8604;
assign v_11049 = v_8604;
assign v_11050 = ~v_8607;
assign v_11051 = ~v_2640;
assign v_11052 = v_2640;
assign v_11053 = ~v_8611;
assign v_11054 = ~v_2644;
assign v_11055 = v_2644;
assign v_11056 = ~v_8615;
assign v_11057 = ~v_2648;
assign v_11058 = v_2648;
assign v_11059 = ~v_8619;
assign v_11060 = ~v_2652;
assign v_11061 = v_2652;
assign v_11062 = ~v_8623;
assign v_11063 = ~v_2656;
assign v_11064 = v_2656;
assign v_11065 = ~v_8627;
assign v_11066 = ~v_2660;
assign v_11067 = v_2660;
assign v_11068 = ~v_8631;
assign v_11069 = ~v_2664;
assign v_11070 = v_2664;
assign v_11071 = ~v_8635;
assign v_11072 = ~v_2668;
assign v_11073 = v_2668;
assign v_11074 = ~v_8639;
assign v_11075 = ~v_2672;
assign v_11076 = v_2672;
assign v_11077 = ~v_8643;
assign v_11078 = ~v_2676;
assign v_11079 = v_2676;
assign v_11080 = ~v_8647;
assign v_11081 = ~v_2680;
assign v_11082 = v_2680;
assign v_11083 = ~v_8651;
assign v_11084 = ~v_2684;
assign v_11085 = v_2684;
assign v_11086 = ~v_8655;
assign v_11087 = ~v_2688;
assign v_11088 = v_11087;
assign v_11090 = v_11089;
assign v_11092 = v_11084 & v_11091;
assign v_11094 = v_8651;
assign v_11096 = v_11093 & v_11095;
assign v_11098 = v_11081 & v_11097;
assign v_11100 = v_8647;
assign v_11102 = v_11099 & v_11101;
assign v_11104 = v_11078 & v_11103;
assign v_11106 = v_8643;
assign v_11108 = v_11105 & v_11107;
assign v_11110 = v_11075 & v_11109;
assign v_11112 = v_8639;
assign v_11114 = v_11111 & v_11113;
assign v_11116 = v_11072 & v_11115;
assign v_11118 = v_8635;
assign v_11120 = v_11117 & v_11119;
assign v_11122 = v_11069 & v_11121;
assign v_11124 = v_8631;
assign v_11126 = v_11123 & v_11125;
assign v_11128 = v_11066 & v_11127;
assign v_11130 = v_8627;
assign v_11132 = v_11129 & v_11131;
assign v_11134 = v_11063 & v_11133;
assign v_11136 = v_8623;
assign v_11138 = v_11135 & v_11137;
assign v_11140 = v_11060 & v_11139;
assign v_11142 = v_8619;
assign v_11144 = v_11141 & v_11143;
assign v_11146 = v_11057 & v_11145;
assign v_11148 = v_8615;
assign v_11150 = v_11147 & v_11149;
assign v_11152 = v_11054 & v_11151;
assign v_11154 = v_8611;
assign v_11156 = v_11153 & v_11155;
assign v_11158 = v_11051 & v_11157;
assign v_11160 = v_8607;
assign v_11162 = v_11159 & v_11161;
assign v_11164 = v_11048 & v_11163;
assign v_11166 = v_2635;
assign v_11168 = v_11165 & v_11167;
assign v_11170 = v_11045 & v_11169;
assign v_11172 = v_2631;
assign v_11174 = v_11171 & v_11173;
assign v_11176 = v_11042 & v_11175;
assign v_11178 = v_2627;
assign v_11180 = v_11177 & v_11179;
assign v_11182 = v_11039 & v_11181;
assign v_11184 = v_2623;
assign v_11186 = v_11183 & v_11185;
assign v_11187 = v_11186;
assign v_11189 = v_8655;
assign v_11190 = v_2688;
assign v_11191 = v_11190;
assign v_11192 = v_11189 & v_11191;
assign v_11193 = v_11192;
assign v_11194 = v_11084 & v_11193;
assign v_11196 = v_11094 & v_11195;
assign v_11197 = v_11083 & v_11193;
assign v_11199 = v_11081 & v_11198;
assign v_11201 = v_11100 & v_11200;
assign v_11202 = v_11080 & v_11198;
assign v_11204 = v_11078 & v_11203;
assign v_11206 = v_11106 & v_11205;
assign v_11207 = v_11077 & v_11203;
assign v_11209 = v_11075 & v_11208;
assign v_11211 = v_11112 & v_11210;
assign v_11212 = v_11074 & v_11208;
assign v_11214 = v_11072 & v_11213;
assign v_11216 = v_11118 & v_11215;
assign v_11217 = v_11071 & v_11213;
assign v_11219 = v_11069 & v_11218;
assign v_11221 = v_11124 & v_11220;
assign v_11222 = v_11068 & v_11218;
assign v_11224 = v_11066 & v_11223;
assign v_11226 = v_11130 & v_11225;
assign v_11227 = v_11065 & v_11223;
assign v_11229 = v_11063 & v_11228;
assign v_11231 = v_11136 & v_11230;
assign v_11232 = v_11062 & v_11228;
assign v_11234 = v_11060 & v_11233;
assign v_11236 = v_11142 & v_11235;
assign v_11237 = v_11059 & v_11233;
assign v_11239 = v_11057 & v_11238;
assign v_11241 = v_11148 & v_11240;
assign v_11242 = v_11056 & v_11238;
assign v_11244 = v_11054 & v_11243;
assign v_11246 = v_11154 & v_11245;
assign v_11247 = v_11053 & v_11243;
assign v_11249 = v_11051 & v_11248;
assign v_11251 = v_11160 & v_11250;
assign v_11252 = v_11050 & v_11248;
assign v_11254 = v_11048 & v_11253;
assign v_11256 = v_11166 & v_11255;
assign v_11257 = v_11047 & v_11253;
assign v_11259 = v_11045 & v_11258;
assign v_11261 = v_11172 & v_11260;
assign v_11262 = v_11044 & v_11258;
assign v_11264 = v_11042 & v_11263;
assign v_11266 = v_11178 & v_11265;
assign v_11267 = v_11041 & v_11263;
assign v_11269 = v_11039 & v_11268;
assign v_11271 = v_11184 & v_11270;
assign v_11272 = v_11038 & v_11268;
assign v_11274 = v_11273;
assign v_11276 = v_11188 & v_11275;
assign v_11277 = v_11276;
assign v_11279 = v_11278;
assign v_11281 = ~v_2883;
assign v_11282 = ~v_8592;
assign v_11283 = v_8592;
assign v_11284 = ~v_2887;
assign v_11285 = ~v_8596;
assign v_11286 = v_8596;
assign v_11287 = ~v_2891;
assign v_11288 = ~v_8600;
assign v_11289 = v_8600;
assign v_11290 = ~v_2895;
assign v_11291 = ~v_8604;
assign v_11292 = v_8604;
assign v_11293 = ~v_8607;
assign v_11294 = ~v_2900;
assign v_11295 = v_2900;
assign v_11296 = ~v_8611;
assign v_11297 = ~v_2904;
assign v_11298 = v_2904;
assign v_11299 = ~v_8615;
assign v_11300 = ~v_2908;
assign v_11301 = v_2908;
assign v_11302 = ~v_8619;
assign v_11303 = ~v_2912;
assign v_11304 = v_2912;
assign v_11305 = ~v_8623;
assign v_11306 = ~v_2916;
assign v_11307 = v_2916;
assign v_11308 = ~v_8627;
assign v_11309 = ~v_2920;
assign v_11310 = v_2920;
assign v_11311 = ~v_8631;
assign v_11312 = ~v_2924;
assign v_11313 = v_2924;
assign v_11314 = ~v_8635;
assign v_11315 = ~v_2928;
assign v_11316 = v_2928;
assign v_11317 = ~v_8639;
assign v_11318 = ~v_2932;
assign v_11319 = v_2932;
assign v_11320 = ~v_8643;
assign v_11321 = ~v_2936;
assign v_11322 = v_2936;
assign v_11323 = ~v_8647;
assign v_11324 = ~v_2940;
assign v_11325 = v_2940;
assign v_11326 = ~v_8651;
assign v_11327 = ~v_2944;
assign v_11328 = v_2944;
assign v_11329 = ~v_8655;
assign v_11330 = ~v_2948;
assign v_11331 = v_11330;
assign v_11333 = v_11332;
assign v_11335 = v_11327 & v_11334;
assign v_11337 = v_8651;
assign v_11339 = v_11336 & v_11338;
assign v_11341 = v_11324 & v_11340;
assign v_11343 = v_8647;
assign v_11345 = v_11342 & v_11344;
assign v_11347 = v_11321 & v_11346;
assign v_11349 = v_8643;
assign v_11351 = v_11348 & v_11350;
assign v_11353 = v_11318 & v_11352;
assign v_11355 = v_8639;
assign v_11357 = v_11354 & v_11356;
assign v_11359 = v_11315 & v_11358;
assign v_11361 = v_8635;
assign v_11363 = v_11360 & v_11362;
assign v_11365 = v_11312 & v_11364;
assign v_11367 = v_8631;
assign v_11369 = v_11366 & v_11368;
assign v_11371 = v_11309 & v_11370;
assign v_11373 = v_8627;
assign v_11375 = v_11372 & v_11374;
assign v_11377 = v_11306 & v_11376;
assign v_11379 = v_8623;
assign v_11381 = v_11378 & v_11380;
assign v_11383 = v_11303 & v_11382;
assign v_11385 = v_8619;
assign v_11387 = v_11384 & v_11386;
assign v_11389 = v_11300 & v_11388;
assign v_11391 = v_8615;
assign v_11393 = v_11390 & v_11392;
assign v_11395 = v_11297 & v_11394;
assign v_11397 = v_8611;
assign v_11399 = v_11396 & v_11398;
assign v_11401 = v_11294 & v_11400;
assign v_11403 = v_8607;
assign v_11405 = v_11402 & v_11404;
assign v_11407 = v_11291 & v_11406;
assign v_11409 = v_2895;
assign v_11411 = v_11408 & v_11410;
assign v_11413 = v_11288 & v_11412;
assign v_11415 = v_2891;
assign v_11417 = v_11414 & v_11416;
assign v_11419 = v_11285 & v_11418;
assign v_11421 = v_2887;
assign v_11423 = v_11420 & v_11422;
assign v_11425 = v_11282 & v_11424;
assign v_11427 = v_2883;
assign v_11429 = v_11426 & v_11428;
assign v_11430 = v_11429;
assign v_11432 = v_8655;
assign v_11433 = v_2948;
assign v_11434 = v_11433;
assign v_11435 = v_11432 & v_11434;
assign v_11436 = v_11435;
assign v_11437 = v_11327 & v_11436;
assign v_11439 = v_11337 & v_11438;
assign v_11440 = v_11326 & v_11436;
assign v_11442 = v_11324 & v_11441;
assign v_11444 = v_11343 & v_11443;
assign v_11445 = v_11323 & v_11441;
assign v_11447 = v_11321 & v_11446;
assign v_11449 = v_11349 & v_11448;
assign v_11450 = v_11320 & v_11446;
assign v_11452 = v_11318 & v_11451;
assign v_11454 = v_11355 & v_11453;
assign v_11455 = v_11317 & v_11451;
assign v_11457 = v_11315 & v_11456;
assign v_11459 = v_11361 & v_11458;
assign v_11460 = v_11314 & v_11456;
assign v_11462 = v_11312 & v_11461;
assign v_11464 = v_11367 & v_11463;
assign v_11465 = v_11311 & v_11461;
assign v_11467 = v_11309 & v_11466;
assign v_11469 = v_11373 & v_11468;
assign v_11470 = v_11308 & v_11466;
assign v_11472 = v_11306 & v_11471;
assign v_11474 = v_11379 & v_11473;
assign v_11475 = v_11305 & v_11471;
assign v_11477 = v_11303 & v_11476;
assign v_11479 = v_11385 & v_11478;
assign v_11480 = v_11302 & v_11476;
assign v_11482 = v_11300 & v_11481;
assign v_11484 = v_11391 & v_11483;
assign v_11485 = v_11299 & v_11481;
assign v_11487 = v_11297 & v_11486;
assign v_11489 = v_11397 & v_11488;
assign v_11490 = v_11296 & v_11486;
assign v_11492 = v_11294 & v_11491;
assign v_11494 = v_11403 & v_11493;
assign v_11495 = v_11293 & v_11491;
assign v_11497 = v_11291 & v_11496;
assign v_11499 = v_11409 & v_11498;
assign v_11500 = v_11290 & v_11496;
assign v_11502 = v_11288 & v_11501;
assign v_11504 = v_11415 & v_11503;
assign v_11505 = v_11287 & v_11501;
assign v_11507 = v_11285 & v_11506;
assign v_11509 = v_11421 & v_11508;
assign v_11510 = v_11284 & v_11506;
assign v_11512 = v_11282 & v_11511;
assign v_11514 = v_11427 & v_11513;
assign v_11515 = v_11281 & v_11511;
assign v_11517 = v_11516;
assign v_11519 = v_11431 & v_11518;
assign v_11520 = v_11519;
assign v_11522 = v_11521;
assign v_11524 = ~v_3143;
assign v_11525 = ~v_8592;
assign v_11526 = v_8592;
assign v_11527 = ~v_3147;
assign v_11528 = ~v_8596;
assign v_11529 = v_8596;
assign v_11530 = ~v_3151;
assign v_11531 = ~v_8600;
assign v_11532 = v_8600;
assign v_11533 = ~v_3155;
assign v_11534 = ~v_8604;
assign v_11535 = v_8604;
assign v_11536 = ~v_8607;
assign v_11537 = ~v_3160;
assign v_11538 = v_3160;
assign v_11539 = ~v_8611;
assign v_11540 = ~v_3164;
assign v_11541 = v_3164;
assign v_11542 = ~v_8615;
assign v_11543 = ~v_3168;
assign v_11544 = v_3168;
assign v_11545 = ~v_8619;
assign v_11546 = ~v_3172;
assign v_11547 = v_3172;
assign v_11548 = ~v_8623;
assign v_11549 = ~v_3176;
assign v_11550 = v_3176;
assign v_11551 = ~v_8627;
assign v_11552 = ~v_3180;
assign v_11553 = v_3180;
assign v_11554 = ~v_8631;
assign v_11555 = ~v_3184;
assign v_11556 = v_3184;
assign v_11557 = ~v_8635;
assign v_11558 = ~v_3188;
assign v_11559 = v_3188;
assign v_11560 = ~v_8639;
assign v_11561 = ~v_3192;
assign v_11562 = v_3192;
assign v_11563 = ~v_8643;
assign v_11564 = ~v_3196;
assign v_11565 = v_3196;
assign v_11566 = ~v_8647;
assign v_11567 = ~v_3200;
assign v_11568 = v_3200;
assign v_11569 = ~v_8651;
assign v_11570 = ~v_3204;
assign v_11571 = v_3204;
assign v_11572 = ~v_8655;
assign v_11573 = ~v_3208;
assign v_11574 = v_11573;
assign v_11576 = v_11575;
assign v_11578 = v_11570 & v_11577;
assign v_11580 = v_8651;
assign v_11582 = v_11579 & v_11581;
assign v_11584 = v_11567 & v_11583;
assign v_11586 = v_8647;
assign v_11588 = v_11585 & v_11587;
assign v_11590 = v_11564 & v_11589;
assign v_11592 = v_8643;
assign v_11594 = v_11591 & v_11593;
assign v_11596 = v_11561 & v_11595;
assign v_11598 = v_8639;
assign v_11600 = v_11597 & v_11599;
assign v_11602 = v_11558 & v_11601;
assign v_11604 = v_8635;
assign v_11606 = v_11603 & v_11605;
assign v_11608 = v_11555 & v_11607;
assign v_11610 = v_8631;
assign v_11612 = v_11609 & v_11611;
assign v_11614 = v_11552 & v_11613;
assign v_11616 = v_8627;
assign v_11618 = v_11615 & v_11617;
assign v_11620 = v_11549 & v_11619;
assign v_11622 = v_8623;
assign v_11624 = v_11621 & v_11623;
assign v_11626 = v_11546 & v_11625;
assign v_11628 = v_8619;
assign v_11630 = v_11627 & v_11629;
assign v_11632 = v_11543 & v_11631;
assign v_11634 = v_8615;
assign v_11636 = v_11633 & v_11635;
assign v_11638 = v_11540 & v_11637;
assign v_11640 = v_8611;
assign v_11642 = v_11639 & v_11641;
assign v_11644 = v_11537 & v_11643;
assign v_11646 = v_8607;
assign v_11648 = v_11645 & v_11647;
assign v_11650 = v_11534 & v_11649;
assign v_11652 = v_3155;
assign v_11654 = v_11651 & v_11653;
assign v_11656 = v_11531 & v_11655;
assign v_11658 = v_3151;
assign v_11660 = v_11657 & v_11659;
assign v_11662 = v_11528 & v_11661;
assign v_11664 = v_3147;
assign v_11666 = v_11663 & v_11665;
assign v_11668 = v_11525 & v_11667;
assign v_11670 = v_3143;
assign v_11672 = v_11669 & v_11671;
assign v_11673 = v_11672;
assign v_11675 = v_8655;
assign v_11676 = v_3208;
assign v_11677 = v_11676;
assign v_11678 = v_11675 & v_11677;
assign v_11679 = v_11678;
assign v_11680 = v_11570 & v_11679;
assign v_11682 = v_11580 & v_11681;
assign v_11683 = v_11569 & v_11679;
assign v_11685 = v_11567 & v_11684;
assign v_11687 = v_11586 & v_11686;
assign v_11688 = v_11566 & v_11684;
assign v_11690 = v_11564 & v_11689;
assign v_11692 = v_11592 & v_11691;
assign v_11693 = v_11563 & v_11689;
assign v_11695 = v_11561 & v_11694;
assign v_11697 = v_11598 & v_11696;
assign v_11698 = v_11560 & v_11694;
assign v_11700 = v_11558 & v_11699;
assign v_11702 = v_11604 & v_11701;
assign v_11703 = v_11557 & v_11699;
assign v_11705 = v_11555 & v_11704;
assign v_11707 = v_11610 & v_11706;
assign v_11708 = v_11554 & v_11704;
assign v_11710 = v_11552 & v_11709;
assign v_11712 = v_11616 & v_11711;
assign v_11713 = v_11551 & v_11709;
assign v_11715 = v_11549 & v_11714;
assign v_11717 = v_11622 & v_11716;
assign v_11718 = v_11548 & v_11714;
assign v_11720 = v_11546 & v_11719;
assign v_11722 = v_11628 & v_11721;
assign v_11723 = v_11545 & v_11719;
assign v_11725 = v_11543 & v_11724;
assign v_11727 = v_11634 & v_11726;
assign v_11728 = v_11542 & v_11724;
assign v_11730 = v_11540 & v_11729;
assign v_11732 = v_11640 & v_11731;
assign v_11733 = v_11539 & v_11729;
assign v_11735 = v_11537 & v_11734;
assign v_11737 = v_11646 & v_11736;
assign v_11738 = v_11536 & v_11734;
assign v_11740 = v_11534 & v_11739;
assign v_11742 = v_11652 & v_11741;
assign v_11743 = v_11533 & v_11739;
assign v_11745 = v_11531 & v_11744;
assign v_11747 = v_11658 & v_11746;
assign v_11748 = v_11530 & v_11744;
assign v_11750 = v_11528 & v_11749;
assign v_11752 = v_11664 & v_11751;
assign v_11753 = v_11527 & v_11749;
assign v_11755 = v_11525 & v_11754;
assign v_11757 = v_11670 & v_11756;
assign v_11758 = v_11524 & v_11754;
assign v_11760 = v_11759;
assign v_11762 = v_11674 & v_11761;
assign v_11763 = v_11762;
assign v_11765 = v_11764;
assign v_11767 = ~v_3403;
assign v_11768 = ~v_8592;
assign v_11769 = v_8592;
assign v_11770 = ~v_3407;
assign v_11771 = ~v_8596;
assign v_11772 = v_8596;
assign v_11773 = ~v_3411;
assign v_11774 = ~v_8600;
assign v_11775 = v_8600;
assign v_11776 = ~v_3415;
assign v_11777 = ~v_8604;
assign v_11778 = v_8604;
assign v_11779 = ~v_8607;
assign v_11780 = ~v_3420;
assign v_11781 = v_3420;
assign v_11782 = ~v_8611;
assign v_11783 = ~v_3424;
assign v_11784 = v_3424;
assign v_11785 = ~v_8615;
assign v_11786 = ~v_3428;
assign v_11787 = v_3428;
assign v_11788 = ~v_8619;
assign v_11789 = ~v_3432;
assign v_11790 = v_3432;
assign v_11791 = ~v_8623;
assign v_11792 = ~v_3436;
assign v_11793 = v_3436;
assign v_11794 = ~v_8627;
assign v_11795 = ~v_3440;
assign v_11796 = v_3440;
assign v_11797 = ~v_8631;
assign v_11798 = ~v_3444;
assign v_11799 = v_3444;
assign v_11800 = ~v_8635;
assign v_11801 = ~v_3448;
assign v_11802 = v_3448;
assign v_11803 = ~v_8639;
assign v_11804 = ~v_3452;
assign v_11805 = v_3452;
assign v_11806 = ~v_8643;
assign v_11807 = ~v_3456;
assign v_11808 = v_3456;
assign v_11809 = ~v_8647;
assign v_11810 = ~v_3460;
assign v_11811 = v_3460;
assign v_11812 = ~v_8651;
assign v_11813 = ~v_3464;
assign v_11814 = v_3464;
assign v_11815 = ~v_8655;
assign v_11816 = ~v_3468;
assign v_11817 = v_11816;
assign v_11819 = v_11818;
assign v_11821 = v_11813 & v_11820;
assign v_11823 = v_8651;
assign v_11825 = v_11822 & v_11824;
assign v_11827 = v_11810 & v_11826;
assign v_11829 = v_8647;
assign v_11831 = v_11828 & v_11830;
assign v_11833 = v_11807 & v_11832;
assign v_11835 = v_8643;
assign v_11837 = v_11834 & v_11836;
assign v_11839 = v_11804 & v_11838;
assign v_11841 = v_8639;
assign v_11843 = v_11840 & v_11842;
assign v_11845 = v_11801 & v_11844;
assign v_11847 = v_8635;
assign v_11849 = v_11846 & v_11848;
assign v_11851 = v_11798 & v_11850;
assign v_11853 = v_8631;
assign v_11855 = v_11852 & v_11854;
assign v_11857 = v_11795 & v_11856;
assign v_11859 = v_8627;
assign v_11861 = v_11858 & v_11860;
assign v_11863 = v_11792 & v_11862;
assign v_11865 = v_8623;
assign v_11867 = v_11864 & v_11866;
assign v_11869 = v_11789 & v_11868;
assign v_11871 = v_8619;
assign v_11873 = v_11870 & v_11872;
assign v_11875 = v_11786 & v_11874;
assign v_11877 = v_8615;
assign v_11879 = v_11876 & v_11878;
assign v_11881 = v_11783 & v_11880;
assign v_11883 = v_8611;
assign v_11885 = v_11882 & v_11884;
assign v_11887 = v_11780 & v_11886;
assign v_11889 = v_8607;
assign v_11891 = v_11888 & v_11890;
assign v_11893 = v_11777 & v_11892;
assign v_11895 = v_3415;
assign v_11897 = v_11894 & v_11896;
assign v_11899 = v_11774 & v_11898;
assign v_11901 = v_3411;
assign v_11903 = v_11900 & v_11902;
assign v_11905 = v_11771 & v_11904;
assign v_11907 = v_3407;
assign v_11909 = v_11906 & v_11908;
assign v_11911 = v_11768 & v_11910;
assign v_11913 = v_3403;
assign v_11915 = v_11912 & v_11914;
assign v_11916 = v_11915;
assign v_11918 = v_8655;
assign v_11919 = v_3468;
assign v_11920 = v_11919;
assign v_11921 = v_11918 & v_11920;
assign v_11922 = v_11921;
assign v_11923 = v_11813 & v_11922;
assign v_11925 = v_11823 & v_11924;
assign v_11926 = v_11812 & v_11922;
assign v_11928 = v_11810 & v_11927;
assign v_11930 = v_11829 & v_11929;
assign v_11931 = v_11809 & v_11927;
assign v_11933 = v_11807 & v_11932;
assign v_11935 = v_11835 & v_11934;
assign v_11936 = v_11806 & v_11932;
assign v_11938 = v_11804 & v_11937;
assign v_11940 = v_11841 & v_11939;
assign v_11941 = v_11803 & v_11937;
assign v_11943 = v_11801 & v_11942;
assign v_11945 = v_11847 & v_11944;
assign v_11946 = v_11800 & v_11942;
assign v_11948 = v_11798 & v_11947;
assign v_11950 = v_11853 & v_11949;
assign v_11951 = v_11797 & v_11947;
assign v_11953 = v_11795 & v_11952;
assign v_11955 = v_11859 & v_11954;
assign v_11956 = v_11794 & v_11952;
assign v_11958 = v_11792 & v_11957;
assign v_11960 = v_11865 & v_11959;
assign v_11961 = v_11791 & v_11957;
assign v_11963 = v_11789 & v_11962;
assign v_11965 = v_11871 & v_11964;
assign v_11966 = v_11788 & v_11962;
assign v_11968 = v_11786 & v_11967;
assign v_11970 = v_11877 & v_11969;
assign v_11971 = v_11785 & v_11967;
assign v_11973 = v_11783 & v_11972;
assign v_11975 = v_11883 & v_11974;
assign v_11976 = v_11782 & v_11972;
assign v_11978 = v_11780 & v_11977;
assign v_11980 = v_11889 & v_11979;
assign v_11981 = v_11779 & v_11977;
assign v_11983 = v_11777 & v_11982;
assign v_11985 = v_11895 & v_11984;
assign v_11986 = v_11776 & v_11982;
assign v_11988 = v_11774 & v_11987;
assign v_11990 = v_11901 & v_11989;
assign v_11991 = v_11773 & v_11987;
assign v_11993 = v_11771 & v_11992;
assign v_11995 = v_11907 & v_11994;
assign v_11996 = v_11770 & v_11992;
assign v_11998 = v_11768 & v_11997;
assign v_12000 = v_11913 & v_11999;
assign v_12001 = v_11767 & v_11997;
assign v_12003 = v_12002;
assign v_12005 = v_11917 & v_12004;
assign v_12006 = v_12005;
assign v_12008 = v_12007;
assign v_12010 = ~v_3663;
assign v_12011 = ~v_8592;
assign v_12012 = v_8592;
assign v_12013 = ~v_3667;
assign v_12014 = ~v_8596;
assign v_12015 = v_8596;
assign v_12016 = ~v_3671;
assign v_12017 = ~v_8600;
assign v_12018 = v_8600;
assign v_12019 = ~v_3675;
assign v_12020 = ~v_8604;
assign v_12021 = v_8604;
assign v_12022 = ~v_8607;
assign v_12023 = ~v_3680;
assign v_12024 = v_3680;
assign v_12025 = ~v_8611;
assign v_12026 = ~v_3684;
assign v_12027 = v_3684;
assign v_12028 = ~v_8615;
assign v_12029 = ~v_3688;
assign v_12030 = v_3688;
assign v_12031 = ~v_8619;
assign v_12032 = ~v_3692;
assign v_12033 = v_3692;
assign v_12034 = ~v_8623;
assign v_12035 = ~v_3696;
assign v_12036 = v_3696;
assign v_12037 = ~v_8627;
assign v_12038 = ~v_3700;
assign v_12039 = v_3700;
assign v_12040 = ~v_8631;
assign v_12041 = ~v_3704;
assign v_12042 = v_3704;
assign v_12043 = ~v_8635;
assign v_12044 = ~v_3708;
assign v_12045 = v_3708;
assign v_12046 = ~v_8639;
assign v_12047 = ~v_3712;
assign v_12048 = v_3712;
assign v_12049 = ~v_8643;
assign v_12050 = ~v_3716;
assign v_12051 = v_3716;
assign v_12052 = ~v_8647;
assign v_12053 = ~v_3720;
assign v_12054 = v_3720;
assign v_12055 = ~v_8651;
assign v_12056 = ~v_3724;
assign v_12057 = v_3724;
assign v_12058 = ~v_8655;
assign v_12059 = ~v_3728;
assign v_12060 = v_12059;
assign v_12062 = v_12061;
assign v_12064 = v_12056 & v_12063;
assign v_12066 = v_8651;
assign v_12068 = v_12065 & v_12067;
assign v_12070 = v_12053 & v_12069;
assign v_12072 = v_8647;
assign v_12074 = v_12071 & v_12073;
assign v_12076 = v_12050 & v_12075;
assign v_12078 = v_8643;
assign v_12080 = v_12077 & v_12079;
assign v_12082 = v_12047 & v_12081;
assign v_12084 = v_8639;
assign v_12086 = v_12083 & v_12085;
assign v_12088 = v_12044 & v_12087;
assign v_12090 = v_8635;
assign v_12092 = v_12089 & v_12091;
assign v_12094 = v_12041 & v_12093;
assign v_12096 = v_8631;
assign v_12098 = v_12095 & v_12097;
assign v_12100 = v_12038 & v_12099;
assign v_12102 = v_8627;
assign v_12104 = v_12101 & v_12103;
assign v_12106 = v_12035 & v_12105;
assign v_12108 = v_8623;
assign v_12110 = v_12107 & v_12109;
assign v_12112 = v_12032 & v_12111;
assign v_12114 = v_8619;
assign v_12116 = v_12113 & v_12115;
assign v_12118 = v_12029 & v_12117;
assign v_12120 = v_8615;
assign v_12122 = v_12119 & v_12121;
assign v_12124 = v_12026 & v_12123;
assign v_12126 = v_8611;
assign v_12128 = v_12125 & v_12127;
assign v_12130 = v_12023 & v_12129;
assign v_12132 = v_8607;
assign v_12134 = v_12131 & v_12133;
assign v_12136 = v_12020 & v_12135;
assign v_12138 = v_3675;
assign v_12140 = v_12137 & v_12139;
assign v_12142 = v_12017 & v_12141;
assign v_12144 = v_3671;
assign v_12146 = v_12143 & v_12145;
assign v_12148 = v_12014 & v_12147;
assign v_12150 = v_3667;
assign v_12152 = v_12149 & v_12151;
assign v_12154 = v_12011 & v_12153;
assign v_12156 = v_3663;
assign v_12158 = v_12155 & v_12157;
assign v_12159 = v_12158;
assign v_12161 = v_8655;
assign v_12162 = v_3728;
assign v_12163 = v_12162;
assign v_12164 = v_12161 & v_12163;
assign v_12165 = v_12164;
assign v_12166 = v_12056 & v_12165;
assign v_12168 = v_12066 & v_12167;
assign v_12169 = v_12055 & v_12165;
assign v_12171 = v_12053 & v_12170;
assign v_12173 = v_12072 & v_12172;
assign v_12174 = v_12052 & v_12170;
assign v_12176 = v_12050 & v_12175;
assign v_12178 = v_12078 & v_12177;
assign v_12179 = v_12049 & v_12175;
assign v_12181 = v_12047 & v_12180;
assign v_12183 = v_12084 & v_12182;
assign v_12184 = v_12046 & v_12180;
assign v_12186 = v_12044 & v_12185;
assign v_12188 = v_12090 & v_12187;
assign v_12189 = v_12043 & v_12185;
assign v_12191 = v_12041 & v_12190;
assign v_12193 = v_12096 & v_12192;
assign v_12194 = v_12040 & v_12190;
assign v_12196 = v_12038 & v_12195;
assign v_12198 = v_12102 & v_12197;
assign v_12199 = v_12037 & v_12195;
assign v_12201 = v_12035 & v_12200;
assign v_12203 = v_12108 & v_12202;
assign v_12204 = v_12034 & v_12200;
assign v_12206 = v_12032 & v_12205;
assign v_12208 = v_12114 & v_12207;
assign v_12209 = v_12031 & v_12205;
assign v_12211 = v_12029 & v_12210;
assign v_12213 = v_12120 & v_12212;
assign v_12214 = v_12028 & v_12210;
assign v_12216 = v_12026 & v_12215;
assign v_12218 = v_12126 & v_12217;
assign v_12219 = v_12025 & v_12215;
assign v_12221 = v_12023 & v_12220;
assign v_12223 = v_12132 & v_12222;
assign v_12224 = v_12022 & v_12220;
assign v_12226 = v_12020 & v_12225;
assign v_12228 = v_12138 & v_12227;
assign v_12229 = v_12019 & v_12225;
assign v_12231 = v_12017 & v_12230;
assign v_12233 = v_12144 & v_12232;
assign v_12234 = v_12016 & v_12230;
assign v_12236 = v_12014 & v_12235;
assign v_12238 = v_12150 & v_12237;
assign v_12239 = v_12013 & v_12235;
assign v_12241 = v_12011 & v_12240;
assign v_12243 = v_12156 & v_12242;
assign v_12244 = v_12010 & v_12240;
assign v_12246 = v_12245;
assign v_12248 = v_12160 & v_12247;
assign v_12249 = v_12248;
assign v_12251 = v_12250;
assign v_12253 = ~v_3923;
assign v_12254 = ~v_8592;
assign v_12255 = v_8592;
assign v_12256 = ~v_3927;
assign v_12257 = ~v_8596;
assign v_12258 = v_8596;
assign v_12259 = ~v_3931;
assign v_12260 = ~v_8600;
assign v_12261 = v_8600;
assign v_12262 = ~v_3935;
assign v_12263 = ~v_8604;
assign v_12264 = v_8604;
assign v_12265 = ~v_8607;
assign v_12266 = ~v_3940;
assign v_12267 = v_3940;
assign v_12268 = ~v_8611;
assign v_12269 = ~v_3944;
assign v_12270 = v_3944;
assign v_12271 = ~v_8615;
assign v_12272 = ~v_3948;
assign v_12273 = v_3948;
assign v_12274 = ~v_8619;
assign v_12275 = ~v_3952;
assign v_12276 = v_3952;
assign v_12277 = ~v_8623;
assign v_12278 = ~v_3956;
assign v_12279 = v_3956;
assign v_12280 = ~v_8627;
assign v_12281 = ~v_3960;
assign v_12282 = v_3960;
assign v_12283 = ~v_8631;
assign v_12284 = ~v_3964;
assign v_12285 = v_3964;
assign v_12286 = ~v_8635;
assign v_12287 = ~v_3968;
assign v_12288 = v_3968;
assign v_12289 = ~v_8639;
assign v_12290 = ~v_3972;
assign v_12291 = v_3972;
assign v_12292 = ~v_8643;
assign v_12293 = ~v_3976;
assign v_12294 = v_3976;
assign v_12295 = ~v_8647;
assign v_12296 = ~v_3980;
assign v_12297 = v_3980;
assign v_12298 = ~v_8651;
assign v_12299 = ~v_3984;
assign v_12300 = v_3984;
assign v_12301 = ~v_8655;
assign v_12302 = ~v_3988;
assign v_12303 = v_12302;
assign v_12305 = v_12304;
assign v_12307 = v_12299 & v_12306;
assign v_12309 = v_8651;
assign v_12311 = v_12308 & v_12310;
assign v_12313 = v_12296 & v_12312;
assign v_12315 = v_8647;
assign v_12317 = v_12314 & v_12316;
assign v_12319 = v_12293 & v_12318;
assign v_12321 = v_8643;
assign v_12323 = v_12320 & v_12322;
assign v_12325 = v_12290 & v_12324;
assign v_12327 = v_8639;
assign v_12329 = v_12326 & v_12328;
assign v_12331 = v_12287 & v_12330;
assign v_12333 = v_8635;
assign v_12335 = v_12332 & v_12334;
assign v_12337 = v_12284 & v_12336;
assign v_12339 = v_8631;
assign v_12341 = v_12338 & v_12340;
assign v_12343 = v_12281 & v_12342;
assign v_12345 = v_8627;
assign v_12347 = v_12344 & v_12346;
assign v_12349 = v_12278 & v_12348;
assign v_12351 = v_8623;
assign v_12353 = v_12350 & v_12352;
assign v_12355 = v_12275 & v_12354;
assign v_12357 = v_8619;
assign v_12359 = v_12356 & v_12358;
assign v_12361 = v_12272 & v_12360;
assign v_12363 = v_8615;
assign v_12365 = v_12362 & v_12364;
assign v_12367 = v_12269 & v_12366;
assign v_12369 = v_8611;
assign v_12371 = v_12368 & v_12370;
assign v_12373 = v_12266 & v_12372;
assign v_12375 = v_8607;
assign v_12377 = v_12374 & v_12376;
assign v_12379 = v_12263 & v_12378;
assign v_12381 = v_3935;
assign v_12383 = v_12380 & v_12382;
assign v_12385 = v_12260 & v_12384;
assign v_12387 = v_3931;
assign v_12389 = v_12386 & v_12388;
assign v_12391 = v_12257 & v_12390;
assign v_12393 = v_3927;
assign v_12395 = v_12392 & v_12394;
assign v_12397 = v_12254 & v_12396;
assign v_12399 = v_3923;
assign v_12401 = v_12398 & v_12400;
assign v_12402 = v_12401;
assign v_12404 = v_8655;
assign v_12405 = v_3988;
assign v_12406 = v_12405;
assign v_12407 = v_12404 & v_12406;
assign v_12408 = v_12407;
assign v_12409 = v_12299 & v_12408;
assign v_12411 = v_12309 & v_12410;
assign v_12412 = v_12298 & v_12408;
assign v_12414 = v_12296 & v_12413;
assign v_12416 = v_12315 & v_12415;
assign v_12417 = v_12295 & v_12413;
assign v_12419 = v_12293 & v_12418;
assign v_12421 = v_12321 & v_12420;
assign v_12422 = v_12292 & v_12418;
assign v_12424 = v_12290 & v_12423;
assign v_12426 = v_12327 & v_12425;
assign v_12427 = v_12289 & v_12423;
assign v_12429 = v_12287 & v_12428;
assign v_12431 = v_12333 & v_12430;
assign v_12432 = v_12286 & v_12428;
assign v_12434 = v_12284 & v_12433;
assign v_12436 = v_12339 & v_12435;
assign v_12437 = v_12283 & v_12433;
assign v_12439 = v_12281 & v_12438;
assign v_12441 = v_12345 & v_12440;
assign v_12442 = v_12280 & v_12438;
assign v_12444 = v_12278 & v_12443;
assign v_12446 = v_12351 & v_12445;
assign v_12447 = v_12277 & v_12443;
assign v_12449 = v_12275 & v_12448;
assign v_12451 = v_12357 & v_12450;
assign v_12452 = v_12274 & v_12448;
assign v_12454 = v_12272 & v_12453;
assign v_12456 = v_12363 & v_12455;
assign v_12457 = v_12271 & v_12453;
assign v_12459 = v_12269 & v_12458;
assign v_12461 = v_12369 & v_12460;
assign v_12462 = v_12268 & v_12458;
assign v_12464 = v_12266 & v_12463;
assign v_12466 = v_12375 & v_12465;
assign v_12467 = v_12265 & v_12463;
assign v_12469 = v_12263 & v_12468;
assign v_12471 = v_12381 & v_12470;
assign v_12472 = v_12262 & v_12468;
assign v_12474 = v_12260 & v_12473;
assign v_12476 = v_12387 & v_12475;
assign v_12477 = v_12259 & v_12473;
assign v_12479 = v_12257 & v_12478;
assign v_12481 = v_12393 & v_12480;
assign v_12482 = v_12256 & v_12478;
assign v_12484 = v_12254 & v_12483;
assign v_12486 = v_12399 & v_12485;
assign v_12487 = v_12253 & v_12483;
assign v_12489 = v_12488;
assign v_12491 = v_12403 & v_12490;
assign v_12492 = v_12491;
assign v_12494 = v_12493;
assign v_12495 = ~v_4182;
assign v_12496 = ~v_8592;
assign v_12497 = v_8592;
assign v_12498 = ~v_4186;
assign v_12499 = ~v_8596;
assign v_12500 = v_8596;
assign v_12501 = ~v_4190;
assign v_12502 = ~v_8600;
assign v_12503 = v_8600;
assign v_12504 = ~v_4194;
assign v_12505 = ~v_8604;
assign v_12506 = v_8604;
assign v_12507 = ~v_8607;
assign v_12508 = ~v_4199;
assign v_12509 = v_4199;
assign v_12510 = ~v_8611;
assign v_12511 = ~v_4203;
assign v_12512 = v_4203;
assign v_12513 = ~v_8615;
assign v_12514 = ~v_4207;
assign v_12515 = v_4207;
assign v_12516 = ~v_8619;
assign v_12517 = ~v_4211;
assign v_12518 = v_4211;
assign v_12519 = ~v_8623;
assign v_12520 = ~v_4215;
assign v_12521 = v_4215;
assign v_12522 = ~v_8627;
assign v_12523 = ~v_4219;
assign v_12524 = v_4219;
assign v_12525 = ~v_8631;
assign v_12526 = ~v_4223;
assign v_12527 = v_4223;
assign v_12528 = ~v_8635;
assign v_12529 = ~v_4227;
assign v_12530 = v_4227;
assign v_12531 = ~v_8639;
assign v_12532 = ~v_4231;
assign v_12533 = v_4231;
assign v_12534 = ~v_8643;
assign v_12535 = ~v_4235;
assign v_12536 = v_4235;
assign v_12537 = ~v_8647;
assign v_12538 = ~v_4239;
assign v_12539 = v_4239;
assign v_12540 = ~v_8651;
assign v_12541 = ~v_4243;
assign v_12542 = v_4243;
assign v_12543 = ~v_8655;
assign v_12544 = ~v_4247;
assign v_12545 = v_12544;
assign v_12547 = v_12546;
assign v_12549 = v_12541 & v_12548;
assign v_12551 = v_8651;
assign v_12553 = v_12550 & v_12552;
assign v_12555 = v_12538 & v_12554;
assign v_12557 = v_8647;
assign v_12559 = v_12556 & v_12558;
assign v_12561 = v_12535 & v_12560;
assign v_12563 = v_8643;
assign v_12565 = v_12562 & v_12564;
assign v_12567 = v_12532 & v_12566;
assign v_12569 = v_8639;
assign v_12571 = v_12568 & v_12570;
assign v_12573 = v_12529 & v_12572;
assign v_12575 = v_8635;
assign v_12577 = v_12574 & v_12576;
assign v_12579 = v_12526 & v_12578;
assign v_12581 = v_8631;
assign v_12583 = v_12580 & v_12582;
assign v_12585 = v_12523 & v_12584;
assign v_12587 = v_8627;
assign v_12589 = v_12586 & v_12588;
assign v_12591 = v_12520 & v_12590;
assign v_12593 = v_8623;
assign v_12595 = v_12592 & v_12594;
assign v_12597 = v_12517 & v_12596;
assign v_12599 = v_8619;
assign v_12601 = v_12598 & v_12600;
assign v_12603 = v_12514 & v_12602;
assign v_12605 = v_8615;
assign v_12607 = v_12604 & v_12606;
assign v_12609 = v_12511 & v_12608;
assign v_12611 = v_8611;
assign v_12613 = v_12610 & v_12612;
assign v_12615 = v_12508 & v_12614;
assign v_12617 = v_8607;
assign v_12619 = v_12616 & v_12618;
assign v_12621 = v_12505 & v_12620;
assign v_12623 = v_4194;
assign v_12625 = v_12622 & v_12624;
assign v_12627 = v_12502 & v_12626;
assign v_12629 = v_4190;
assign v_12631 = v_12628 & v_12630;
assign v_12633 = v_12499 & v_12632;
assign v_12635 = v_4186;
assign v_12637 = v_12634 & v_12636;
assign v_12639 = v_12496 & v_12638;
assign v_12641 = v_4182;
assign v_12643 = v_12640 & v_12642;
assign v_12645 = ~v_12644;
assign v_12647 = v_8655;
assign v_12648 = v_4247;
assign v_12649 = v_12648;
assign v_12650 = v_12647 & v_12649;
assign v_12651 = v_12650;
assign v_12652 = v_12541 & v_12651;
assign v_12654 = v_12551 & v_12653;
assign v_12655 = v_12540 & v_12651;
assign v_12657 = v_12538 & v_12656;
assign v_12659 = v_12557 & v_12658;
assign v_12660 = v_12537 & v_12656;
assign v_12662 = v_12535 & v_12661;
assign v_12664 = v_12563 & v_12663;
assign v_12665 = v_12534 & v_12661;
assign v_12667 = v_12532 & v_12666;
assign v_12669 = v_12569 & v_12668;
assign v_12670 = v_12531 & v_12666;
assign v_12672 = v_12529 & v_12671;
assign v_12674 = v_12575 & v_12673;
assign v_12675 = v_12528 & v_12671;
assign v_12677 = v_12526 & v_12676;
assign v_12679 = v_12581 & v_12678;
assign v_12680 = v_12525 & v_12676;
assign v_12682 = v_12523 & v_12681;
assign v_12684 = v_12587 & v_12683;
assign v_12685 = v_12522 & v_12681;
assign v_12687 = v_12520 & v_12686;
assign v_12689 = v_12593 & v_12688;
assign v_12690 = v_12519 & v_12686;
assign v_12692 = v_12517 & v_12691;
assign v_12694 = v_12599 & v_12693;
assign v_12695 = v_12516 & v_12691;
assign v_12697 = v_12514 & v_12696;
assign v_12699 = v_12605 & v_12698;
assign v_12700 = v_12513 & v_12696;
assign v_12702 = v_12511 & v_12701;
assign v_12704 = v_12611 & v_12703;
assign v_12705 = v_12510 & v_12701;
assign v_12707 = v_12508 & v_12706;
assign v_12709 = v_12617 & v_12708;
assign v_12710 = v_12507 & v_12706;
assign v_12712 = v_12505 & v_12711;
assign v_12714 = v_12623 & v_12713;
assign v_12715 = v_12504 & v_12711;
assign v_12717 = v_12502 & v_12716;
assign v_12719 = v_12629 & v_12718;
assign v_12720 = v_12501 & v_12716;
assign v_12722 = v_12499 & v_12721;
assign v_12724 = v_12635 & v_12723;
assign v_12725 = v_12498 & v_12721;
assign v_12727 = v_12496 & v_12726;
assign v_12729 = v_12641 & v_12728;
assign v_12730 = v_12495 & v_12726;
assign v_12732 = v_12644;
assign v_12734 = v_12646 & v_12733;
assign v_12735 = v_12734;
assign v_12737 = v_12736;
assign v_12739 = ~v_6;
assign v_12741 = ~v_12740;
assign v_12742 = v_12740;
assign v_12743 = ~v_13;
assign v_12745 = ~v_12744;
assign v_12746 = v_12744;
assign v_12747 = ~v_18;
assign v_12749 = ~v_12748;
assign v_12750 = v_12748;
assign v_12751 = ~v_23;
assign v_12753 = ~v_12752;
assign v_12754 = v_12752;
assign v_12756 = ~v_12755;
assign v_12757 = ~v_30;
assign v_12758 = v_30;
assign v_12760 = ~v_12759;
assign v_12761 = ~v_35;
assign v_12762 = v_35;
assign v_12764 = ~v_12763;
assign v_12765 = ~v_40;
assign v_12766 = v_40;
assign v_12768 = ~v_12767;
assign v_12769 = ~v_45;
assign v_12770 = v_45;
assign v_12772 = ~v_12771;
assign v_12773 = ~v_50;
assign v_12774 = v_50;
assign v_12776 = ~v_12775;
assign v_12777 = ~v_55;
assign v_12778 = v_55;
assign v_12780 = ~v_12779;
assign v_12781 = ~v_60;
assign v_12782 = v_60;
assign v_12784 = ~v_12783;
assign v_12785 = ~v_65;
assign v_12786 = v_65;
assign v_12788 = ~v_12787;
assign v_12789 = ~v_70;
assign v_12790 = v_70;
assign v_12792 = ~v_12791;
assign v_12793 = ~v_75;
assign v_12794 = v_75;
assign v_12796 = ~v_12795;
assign v_12797 = ~v_80;
assign v_12798 = v_80;
assign v_12800 = ~v_12799;
assign v_12801 = ~v_85;
assign v_12802 = v_85;
assign v_12804 = ~v_12803;
assign v_12805 = ~v_90;
assign v_12806 = v_12805;
assign v_12808 = v_12807;
assign v_12810 = v_12801 & v_12809;
assign v_12812 = v_12799;
assign v_12814 = v_12811 & v_12813;
assign v_12816 = v_12797 & v_12815;
assign v_12818 = v_12795;
assign v_12820 = v_12817 & v_12819;
assign v_12822 = v_12793 & v_12821;
assign v_12824 = v_12791;
assign v_12826 = v_12823 & v_12825;
assign v_12828 = v_12789 & v_12827;
assign v_12830 = v_12787;
assign v_12832 = v_12829 & v_12831;
assign v_12834 = v_12785 & v_12833;
assign v_12836 = v_12783;
assign v_12838 = v_12835 & v_12837;
assign v_12840 = v_12781 & v_12839;
assign v_12842 = v_12779;
assign v_12844 = v_12841 & v_12843;
assign v_12846 = v_12777 & v_12845;
assign v_12848 = v_12775;
assign v_12850 = v_12847 & v_12849;
assign v_12852 = v_12773 & v_12851;
assign v_12854 = v_12771;
assign v_12856 = v_12853 & v_12855;
assign v_12858 = v_12769 & v_12857;
assign v_12860 = v_12767;
assign v_12862 = v_12859 & v_12861;
assign v_12864 = v_12765 & v_12863;
assign v_12866 = v_12763;
assign v_12868 = v_12865 & v_12867;
assign v_12870 = v_12761 & v_12869;
assign v_12872 = v_12759;
assign v_12874 = v_12871 & v_12873;
assign v_12876 = v_12757 & v_12875;
assign v_12878 = v_12755;
assign v_12880 = v_12877 & v_12879;
assign v_12882 = v_12753 & v_12881;
assign v_12884 = v_23;
assign v_12886 = v_12883 & v_12885;
assign v_12888 = v_12749 & v_12887;
assign v_12890 = v_18;
assign v_12892 = v_12889 & v_12891;
assign v_12894 = v_12745 & v_12893;
assign v_12896 = v_13;
assign v_12898 = v_12895 & v_12897;
assign v_12900 = v_12741 & v_12899;
assign v_12902 = v_6;
assign v_12904 = v_12901 & v_12903;
assign v_12905 = v_12904;
assign v_12907 = v_12803;
assign v_12908 = v_90;
assign v_12909 = v_12908;
assign v_12910 = v_12907 & v_12909;
assign v_12911 = v_12910;
assign v_12912 = v_12801 & v_12911;
assign v_12914 = v_12812 & v_12913;
assign v_12915 = v_12800 & v_12911;
assign v_12917 = v_12797 & v_12916;
assign v_12919 = v_12818 & v_12918;
assign v_12920 = v_12796 & v_12916;
assign v_12922 = v_12793 & v_12921;
assign v_12924 = v_12824 & v_12923;
assign v_12925 = v_12792 & v_12921;
assign v_12927 = v_12789 & v_12926;
assign v_12929 = v_12830 & v_12928;
assign v_12930 = v_12788 & v_12926;
assign v_12932 = v_12785 & v_12931;
assign v_12934 = v_12836 & v_12933;
assign v_12935 = v_12784 & v_12931;
assign v_12937 = v_12781 & v_12936;
assign v_12939 = v_12842 & v_12938;
assign v_12940 = v_12780 & v_12936;
assign v_12942 = v_12777 & v_12941;
assign v_12944 = v_12848 & v_12943;
assign v_12945 = v_12776 & v_12941;
assign v_12947 = v_12773 & v_12946;
assign v_12949 = v_12854 & v_12948;
assign v_12950 = v_12772 & v_12946;
assign v_12952 = v_12769 & v_12951;
assign v_12954 = v_12860 & v_12953;
assign v_12955 = v_12768 & v_12951;
assign v_12957 = v_12765 & v_12956;
assign v_12959 = v_12866 & v_12958;
assign v_12960 = v_12764 & v_12956;
assign v_12962 = v_12761 & v_12961;
assign v_12964 = v_12872 & v_12963;
assign v_12965 = v_12760 & v_12961;
assign v_12967 = v_12757 & v_12966;
assign v_12969 = v_12878 & v_12968;
assign v_12970 = v_12756 & v_12966;
assign v_12972 = v_12753 & v_12971;
assign v_12974 = v_12884 & v_12973;
assign v_12975 = v_12751 & v_12971;
assign v_12977 = v_12749 & v_12976;
assign v_12979 = v_12890 & v_12978;
assign v_12980 = v_12747 & v_12976;
assign v_12982 = v_12745 & v_12981;
assign v_12984 = v_12896 & v_12983;
assign v_12985 = v_12743 & v_12981;
assign v_12987 = v_12741 & v_12986;
assign v_12989 = v_12902 & v_12988;
assign v_12990 = v_12739 & v_12986;
assign v_12992 = v_12991;
assign v_12994 = v_12906 & v_12993;
assign v_12995 = v_12994;
assign v_12997 = v_12996;
assign v_12999 = ~v_283;
assign v_13000 = ~v_12740;
assign v_13001 = v_12740;
assign v_13002 = ~v_287;
assign v_13003 = ~v_12744;
assign v_13004 = v_12744;
assign v_13005 = ~v_291;
assign v_13006 = ~v_12748;
assign v_13007 = v_12748;
assign v_13008 = ~v_295;
assign v_13009 = ~v_12752;
assign v_13010 = v_12752;
assign v_13011 = ~v_12755;
assign v_13012 = ~v_300;
assign v_13013 = v_300;
assign v_13014 = ~v_12759;
assign v_13015 = ~v_304;
assign v_13016 = v_304;
assign v_13017 = ~v_12763;
assign v_13018 = ~v_308;
assign v_13019 = v_308;
assign v_13020 = ~v_12767;
assign v_13021 = ~v_312;
assign v_13022 = v_312;
assign v_13023 = ~v_12771;
assign v_13024 = ~v_316;
assign v_13025 = v_316;
assign v_13026 = ~v_12775;
assign v_13027 = ~v_320;
assign v_13028 = v_320;
assign v_13029 = ~v_12779;
assign v_13030 = ~v_324;
assign v_13031 = v_324;
assign v_13032 = ~v_12783;
assign v_13033 = ~v_328;
assign v_13034 = v_328;
assign v_13035 = ~v_12787;
assign v_13036 = ~v_332;
assign v_13037 = v_332;
assign v_13038 = ~v_12791;
assign v_13039 = ~v_336;
assign v_13040 = v_336;
assign v_13041 = ~v_12795;
assign v_13042 = ~v_340;
assign v_13043 = v_340;
assign v_13044 = ~v_12799;
assign v_13045 = ~v_344;
assign v_13046 = v_344;
assign v_13047 = ~v_12803;
assign v_13048 = ~v_348;
assign v_13049 = v_13048;
assign v_13051 = v_13050;
assign v_13053 = v_13045 & v_13052;
assign v_13055 = v_12799;
assign v_13057 = v_13054 & v_13056;
assign v_13059 = v_13042 & v_13058;
assign v_13061 = v_12795;
assign v_13063 = v_13060 & v_13062;
assign v_13065 = v_13039 & v_13064;
assign v_13067 = v_12791;
assign v_13069 = v_13066 & v_13068;
assign v_13071 = v_13036 & v_13070;
assign v_13073 = v_12787;
assign v_13075 = v_13072 & v_13074;
assign v_13077 = v_13033 & v_13076;
assign v_13079 = v_12783;
assign v_13081 = v_13078 & v_13080;
assign v_13083 = v_13030 & v_13082;
assign v_13085 = v_12779;
assign v_13087 = v_13084 & v_13086;
assign v_13089 = v_13027 & v_13088;
assign v_13091 = v_12775;
assign v_13093 = v_13090 & v_13092;
assign v_13095 = v_13024 & v_13094;
assign v_13097 = v_12771;
assign v_13099 = v_13096 & v_13098;
assign v_13101 = v_13021 & v_13100;
assign v_13103 = v_12767;
assign v_13105 = v_13102 & v_13104;
assign v_13107 = v_13018 & v_13106;
assign v_13109 = v_12763;
assign v_13111 = v_13108 & v_13110;
assign v_13113 = v_13015 & v_13112;
assign v_13115 = v_12759;
assign v_13117 = v_13114 & v_13116;
assign v_13119 = v_13012 & v_13118;
assign v_13121 = v_12755;
assign v_13123 = v_13120 & v_13122;
assign v_13125 = v_13009 & v_13124;
assign v_13127 = v_295;
assign v_13129 = v_13126 & v_13128;
assign v_13131 = v_13006 & v_13130;
assign v_13133 = v_291;
assign v_13135 = v_13132 & v_13134;
assign v_13137 = v_13003 & v_13136;
assign v_13139 = v_287;
assign v_13141 = v_13138 & v_13140;
assign v_13143 = v_13000 & v_13142;
assign v_13145 = v_283;
assign v_13147 = v_13144 & v_13146;
assign v_13148 = v_13147;
assign v_13150 = v_12803;
assign v_13151 = v_348;
assign v_13152 = v_13151;
assign v_13153 = v_13150 & v_13152;
assign v_13154 = v_13153;
assign v_13155 = v_13045 & v_13154;
assign v_13157 = v_13055 & v_13156;
assign v_13158 = v_13044 & v_13154;
assign v_13160 = v_13042 & v_13159;
assign v_13162 = v_13061 & v_13161;
assign v_13163 = v_13041 & v_13159;
assign v_13165 = v_13039 & v_13164;
assign v_13167 = v_13067 & v_13166;
assign v_13168 = v_13038 & v_13164;
assign v_13170 = v_13036 & v_13169;
assign v_13172 = v_13073 & v_13171;
assign v_13173 = v_13035 & v_13169;
assign v_13175 = v_13033 & v_13174;
assign v_13177 = v_13079 & v_13176;
assign v_13178 = v_13032 & v_13174;
assign v_13180 = v_13030 & v_13179;
assign v_13182 = v_13085 & v_13181;
assign v_13183 = v_13029 & v_13179;
assign v_13185 = v_13027 & v_13184;
assign v_13187 = v_13091 & v_13186;
assign v_13188 = v_13026 & v_13184;
assign v_13190 = v_13024 & v_13189;
assign v_13192 = v_13097 & v_13191;
assign v_13193 = v_13023 & v_13189;
assign v_13195 = v_13021 & v_13194;
assign v_13197 = v_13103 & v_13196;
assign v_13198 = v_13020 & v_13194;
assign v_13200 = v_13018 & v_13199;
assign v_13202 = v_13109 & v_13201;
assign v_13203 = v_13017 & v_13199;
assign v_13205 = v_13015 & v_13204;
assign v_13207 = v_13115 & v_13206;
assign v_13208 = v_13014 & v_13204;
assign v_13210 = v_13012 & v_13209;
assign v_13212 = v_13121 & v_13211;
assign v_13213 = v_13011 & v_13209;
assign v_13215 = v_13009 & v_13214;
assign v_13217 = v_13127 & v_13216;
assign v_13218 = v_13008 & v_13214;
assign v_13220 = v_13006 & v_13219;
assign v_13222 = v_13133 & v_13221;
assign v_13223 = v_13005 & v_13219;
assign v_13225 = v_13003 & v_13224;
assign v_13227 = v_13139 & v_13226;
assign v_13228 = v_13002 & v_13224;
assign v_13230 = v_13000 & v_13229;
assign v_13232 = v_13145 & v_13231;
assign v_13233 = v_12999 & v_13229;
assign v_13235 = v_13234;
assign v_13237 = v_13149 & v_13236;
assign v_13238 = v_13237;
assign v_13240 = v_13239;
assign v_13242 = ~v_543;
assign v_13243 = ~v_12740;
assign v_13244 = v_12740;
assign v_13245 = ~v_547;
assign v_13246 = ~v_12744;
assign v_13247 = v_12744;
assign v_13248 = ~v_551;
assign v_13249 = ~v_12748;
assign v_13250 = v_12748;
assign v_13251 = ~v_555;
assign v_13252 = ~v_12752;
assign v_13253 = v_12752;
assign v_13254 = ~v_12755;
assign v_13255 = ~v_560;
assign v_13256 = v_560;
assign v_13257 = ~v_12759;
assign v_13258 = ~v_564;
assign v_13259 = v_564;
assign v_13260 = ~v_12763;
assign v_13261 = ~v_568;
assign v_13262 = v_568;
assign v_13263 = ~v_12767;
assign v_13264 = ~v_572;
assign v_13265 = v_572;
assign v_13266 = ~v_12771;
assign v_13267 = ~v_576;
assign v_13268 = v_576;
assign v_13269 = ~v_12775;
assign v_13270 = ~v_580;
assign v_13271 = v_580;
assign v_13272 = ~v_12779;
assign v_13273 = ~v_584;
assign v_13274 = v_584;
assign v_13275 = ~v_12783;
assign v_13276 = ~v_588;
assign v_13277 = v_588;
assign v_13278 = ~v_12787;
assign v_13279 = ~v_592;
assign v_13280 = v_592;
assign v_13281 = ~v_12791;
assign v_13282 = ~v_596;
assign v_13283 = v_596;
assign v_13284 = ~v_12795;
assign v_13285 = ~v_600;
assign v_13286 = v_600;
assign v_13287 = ~v_12799;
assign v_13288 = ~v_604;
assign v_13289 = v_604;
assign v_13290 = ~v_12803;
assign v_13291 = ~v_608;
assign v_13292 = v_13291;
assign v_13294 = v_13293;
assign v_13296 = v_13288 & v_13295;
assign v_13298 = v_12799;
assign v_13300 = v_13297 & v_13299;
assign v_13302 = v_13285 & v_13301;
assign v_13304 = v_12795;
assign v_13306 = v_13303 & v_13305;
assign v_13308 = v_13282 & v_13307;
assign v_13310 = v_12791;
assign v_13312 = v_13309 & v_13311;
assign v_13314 = v_13279 & v_13313;
assign v_13316 = v_12787;
assign v_13318 = v_13315 & v_13317;
assign v_13320 = v_13276 & v_13319;
assign v_13322 = v_12783;
assign v_13324 = v_13321 & v_13323;
assign v_13326 = v_13273 & v_13325;
assign v_13328 = v_12779;
assign v_13330 = v_13327 & v_13329;
assign v_13332 = v_13270 & v_13331;
assign v_13334 = v_12775;
assign v_13336 = v_13333 & v_13335;
assign v_13338 = v_13267 & v_13337;
assign v_13340 = v_12771;
assign v_13342 = v_13339 & v_13341;
assign v_13344 = v_13264 & v_13343;
assign v_13346 = v_12767;
assign v_13348 = v_13345 & v_13347;
assign v_13350 = v_13261 & v_13349;
assign v_13352 = v_12763;
assign v_13354 = v_13351 & v_13353;
assign v_13356 = v_13258 & v_13355;
assign v_13358 = v_12759;
assign v_13360 = v_13357 & v_13359;
assign v_13362 = v_13255 & v_13361;
assign v_13364 = v_12755;
assign v_13366 = v_13363 & v_13365;
assign v_13368 = v_13252 & v_13367;
assign v_13370 = v_555;
assign v_13372 = v_13369 & v_13371;
assign v_13374 = v_13249 & v_13373;
assign v_13376 = v_551;
assign v_13378 = v_13375 & v_13377;
assign v_13380 = v_13246 & v_13379;
assign v_13382 = v_547;
assign v_13384 = v_13381 & v_13383;
assign v_13386 = v_13243 & v_13385;
assign v_13388 = v_543;
assign v_13390 = v_13387 & v_13389;
assign v_13391 = v_13390;
assign v_13393 = v_12803;
assign v_13394 = v_608;
assign v_13395 = v_13394;
assign v_13396 = v_13393 & v_13395;
assign v_13397 = v_13396;
assign v_13398 = v_13288 & v_13397;
assign v_13400 = v_13298 & v_13399;
assign v_13401 = v_13287 & v_13397;
assign v_13403 = v_13285 & v_13402;
assign v_13405 = v_13304 & v_13404;
assign v_13406 = v_13284 & v_13402;
assign v_13408 = v_13282 & v_13407;
assign v_13410 = v_13310 & v_13409;
assign v_13411 = v_13281 & v_13407;
assign v_13413 = v_13279 & v_13412;
assign v_13415 = v_13316 & v_13414;
assign v_13416 = v_13278 & v_13412;
assign v_13418 = v_13276 & v_13417;
assign v_13420 = v_13322 & v_13419;
assign v_13421 = v_13275 & v_13417;
assign v_13423 = v_13273 & v_13422;
assign v_13425 = v_13328 & v_13424;
assign v_13426 = v_13272 & v_13422;
assign v_13428 = v_13270 & v_13427;
assign v_13430 = v_13334 & v_13429;
assign v_13431 = v_13269 & v_13427;
assign v_13433 = v_13267 & v_13432;
assign v_13435 = v_13340 & v_13434;
assign v_13436 = v_13266 & v_13432;
assign v_13438 = v_13264 & v_13437;
assign v_13440 = v_13346 & v_13439;
assign v_13441 = v_13263 & v_13437;
assign v_13443 = v_13261 & v_13442;
assign v_13445 = v_13352 & v_13444;
assign v_13446 = v_13260 & v_13442;
assign v_13448 = v_13258 & v_13447;
assign v_13450 = v_13358 & v_13449;
assign v_13451 = v_13257 & v_13447;
assign v_13453 = v_13255 & v_13452;
assign v_13455 = v_13364 & v_13454;
assign v_13456 = v_13254 & v_13452;
assign v_13458 = v_13252 & v_13457;
assign v_13460 = v_13370 & v_13459;
assign v_13461 = v_13251 & v_13457;
assign v_13463 = v_13249 & v_13462;
assign v_13465 = v_13376 & v_13464;
assign v_13466 = v_13248 & v_13462;
assign v_13468 = v_13246 & v_13467;
assign v_13470 = v_13382 & v_13469;
assign v_13471 = v_13245 & v_13467;
assign v_13473 = v_13243 & v_13472;
assign v_13475 = v_13388 & v_13474;
assign v_13476 = v_13242 & v_13472;
assign v_13478 = v_13477;
assign v_13480 = v_13392 & v_13479;
assign v_13481 = v_13480;
assign v_13483 = v_13482;
assign v_13485 = ~v_803;
assign v_13486 = ~v_12740;
assign v_13487 = v_12740;
assign v_13488 = ~v_807;
assign v_13489 = ~v_12744;
assign v_13490 = v_12744;
assign v_13491 = ~v_811;
assign v_13492 = ~v_12748;
assign v_13493 = v_12748;
assign v_13494 = ~v_815;
assign v_13495 = ~v_12752;
assign v_13496 = v_12752;
assign v_13497 = ~v_12755;
assign v_13498 = ~v_820;
assign v_13499 = v_820;
assign v_13500 = ~v_12759;
assign v_13501 = ~v_824;
assign v_13502 = v_824;
assign v_13503 = ~v_12763;
assign v_13504 = ~v_828;
assign v_13505 = v_828;
assign v_13506 = ~v_12767;
assign v_13507 = ~v_832;
assign v_13508 = v_832;
assign v_13509 = ~v_12771;
assign v_13510 = ~v_836;
assign v_13511 = v_836;
assign v_13512 = ~v_12775;
assign v_13513 = ~v_840;
assign v_13514 = v_840;
assign v_13515 = ~v_12779;
assign v_13516 = ~v_844;
assign v_13517 = v_844;
assign v_13518 = ~v_12783;
assign v_13519 = ~v_848;
assign v_13520 = v_848;
assign v_13521 = ~v_12787;
assign v_13522 = ~v_852;
assign v_13523 = v_852;
assign v_13524 = ~v_12791;
assign v_13525 = ~v_856;
assign v_13526 = v_856;
assign v_13527 = ~v_12795;
assign v_13528 = ~v_860;
assign v_13529 = v_860;
assign v_13530 = ~v_12799;
assign v_13531 = ~v_864;
assign v_13532 = v_864;
assign v_13533 = ~v_12803;
assign v_13534 = ~v_868;
assign v_13535 = v_13534;
assign v_13537 = v_13536;
assign v_13539 = v_13531 & v_13538;
assign v_13541 = v_12799;
assign v_13543 = v_13540 & v_13542;
assign v_13545 = v_13528 & v_13544;
assign v_13547 = v_12795;
assign v_13549 = v_13546 & v_13548;
assign v_13551 = v_13525 & v_13550;
assign v_13553 = v_12791;
assign v_13555 = v_13552 & v_13554;
assign v_13557 = v_13522 & v_13556;
assign v_13559 = v_12787;
assign v_13561 = v_13558 & v_13560;
assign v_13563 = v_13519 & v_13562;
assign v_13565 = v_12783;
assign v_13567 = v_13564 & v_13566;
assign v_13569 = v_13516 & v_13568;
assign v_13571 = v_12779;
assign v_13573 = v_13570 & v_13572;
assign v_13575 = v_13513 & v_13574;
assign v_13577 = v_12775;
assign v_13579 = v_13576 & v_13578;
assign v_13581 = v_13510 & v_13580;
assign v_13583 = v_12771;
assign v_13585 = v_13582 & v_13584;
assign v_13587 = v_13507 & v_13586;
assign v_13589 = v_12767;
assign v_13591 = v_13588 & v_13590;
assign v_13593 = v_13504 & v_13592;
assign v_13595 = v_12763;
assign v_13597 = v_13594 & v_13596;
assign v_13599 = v_13501 & v_13598;
assign v_13601 = v_12759;
assign v_13603 = v_13600 & v_13602;
assign v_13605 = v_13498 & v_13604;
assign v_13607 = v_12755;
assign v_13609 = v_13606 & v_13608;
assign v_13611 = v_13495 & v_13610;
assign v_13613 = v_815;
assign v_13615 = v_13612 & v_13614;
assign v_13617 = v_13492 & v_13616;
assign v_13619 = v_811;
assign v_13621 = v_13618 & v_13620;
assign v_13623 = v_13489 & v_13622;
assign v_13625 = v_807;
assign v_13627 = v_13624 & v_13626;
assign v_13629 = v_13486 & v_13628;
assign v_13631 = v_803;
assign v_13633 = v_13630 & v_13632;
assign v_13634 = v_13633;
assign v_13636 = v_12803;
assign v_13637 = v_868;
assign v_13638 = v_13637;
assign v_13639 = v_13636 & v_13638;
assign v_13640 = v_13639;
assign v_13641 = v_13531 & v_13640;
assign v_13643 = v_13541 & v_13642;
assign v_13644 = v_13530 & v_13640;
assign v_13646 = v_13528 & v_13645;
assign v_13648 = v_13547 & v_13647;
assign v_13649 = v_13527 & v_13645;
assign v_13651 = v_13525 & v_13650;
assign v_13653 = v_13553 & v_13652;
assign v_13654 = v_13524 & v_13650;
assign v_13656 = v_13522 & v_13655;
assign v_13658 = v_13559 & v_13657;
assign v_13659 = v_13521 & v_13655;
assign v_13661 = v_13519 & v_13660;
assign v_13663 = v_13565 & v_13662;
assign v_13664 = v_13518 & v_13660;
assign v_13666 = v_13516 & v_13665;
assign v_13668 = v_13571 & v_13667;
assign v_13669 = v_13515 & v_13665;
assign v_13671 = v_13513 & v_13670;
assign v_13673 = v_13577 & v_13672;
assign v_13674 = v_13512 & v_13670;
assign v_13676 = v_13510 & v_13675;
assign v_13678 = v_13583 & v_13677;
assign v_13679 = v_13509 & v_13675;
assign v_13681 = v_13507 & v_13680;
assign v_13683 = v_13589 & v_13682;
assign v_13684 = v_13506 & v_13680;
assign v_13686 = v_13504 & v_13685;
assign v_13688 = v_13595 & v_13687;
assign v_13689 = v_13503 & v_13685;
assign v_13691 = v_13501 & v_13690;
assign v_13693 = v_13601 & v_13692;
assign v_13694 = v_13500 & v_13690;
assign v_13696 = v_13498 & v_13695;
assign v_13698 = v_13607 & v_13697;
assign v_13699 = v_13497 & v_13695;
assign v_13701 = v_13495 & v_13700;
assign v_13703 = v_13613 & v_13702;
assign v_13704 = v_13494 & v_13700;
assign v_13706 = v_13492 & v_13705;
assign v_13708 = v_13619 & v_13707;
assign v_13709 = v_13491 & v_13705;
assign v_13711 = v_13489 & v_13710;
assign v_13713 = v_13625 & v_13712;
assign v_13714 = v_13488 & v_13710;
assign v_13716 = v_13486 & v_13715;
assign v_13718 = v_13631 & v_13717;
assign v_13719 = v_13485 & v_13715;
assign v_13721 = v_13720;
assign v_13723 = v_13635 & v_13722;
assign v_13724 = v_13723;
assign v_13726 = v_13725;
assign v_13728 = ~v_1063;
assign v_13729 = ~v_12740;
assign v_13730 = v_12740;
assign v_13731 = ~v_1067;
assign v_13732 = ~v_12744;
assign v_13733 = v_12744;
assign v_13734 = ~v_1071;
assign v_13735 = ~v_12748;
assign v_13736 = v_12748;
assign v_13737 = ~v_1075;
assign v_13738 = ~v_12752;
assign v_13739 = v_12752;
assign v_13740 = ~v_12755;
assign v_13741 = ~v_1080;
assign v_13742 = v_1080;
assign v_13743 = ~v_12759;
assign v_13744 = ~v_1084;
assign v_13745 = v_1084;
assign v_13746 = ~v_12763;
assign v_13747 = ~v_1088;
assign v_13748 = v_1088;
assign v_13749 = ~v_12767;
assign v_13750 = ~v_1092;
assign v_13751 = v_1092;
assign v_13752 = ~v_12771;
assign v_13753 = ~v_1096;
assign v_13754 = v_1096;
assign v_13755 = ~v_12775;
assign v_13756 = ~v_1100;
assign v_13757 = v_1100;
assign v_13758 = ~v_12779;
assign v_13759 = ~v_1104;
assign v_13760 = v_1104;
assign v_13761 = ~v_12783;
assign v_13762 = ~v_1108;
assign v_13763 = v_1108;
assign v_13764 = ~v_12787;
assign v_13765 = ~v_1112;
assign v_13766 = v_1112;
assign v_13767 = ~v_12791;
assign v_13768 = ~v_1116;
assign v_13769 = v_1116;
assign v_13770 = ~v_12795;
assign v_13771 = ~v_1120;
assign v_13772 = v_1120;
assign v_13773 = ~v_12799;
assign v_13774 = ~v_1124;
assign v_13775 = v_1124;
assign v_13776 = ~v_12803;
assign v_13777 = ~v_1128;
assign v_13778 = v_13777;
assign v_13780 = v_13779;
assign v_13782 = v_13774 & v_13781;
assign v_13784 = v_12799;
assign v_13786 = v_13783 & v_13785;
assign v_13788 = v_13771 & v_13787;
assign v_13790 = v_12795;
assign v_13792 = v_13789 & v_13791;
assign v_13794 = v_13768 & v_13793;
assign v_13796 = v_12791;
assign v_13798 = v_13795 & v_13797;
assign v_13800 = v_13765 & v_13799;
assign v_13802 = v_12787;
assign v_13804 = v_13801 & v_13803;
assign v_13806 = v_13762 & v_13805;
assign v_13808 = v_12783;
assign v_13810 = v_13807 & v_13809;
assign v_13812 = v_13759 & v_13811;
assign v_13814 = v_12779;
assign v_13816 = v_13813 & v_13815;
assign v_13818 = v_13756 & v_13817;
assign v_13820 = v_12775;
assign v_13822 = v_13819 & v_13821;
assign v_13824 = v_13753 & v_13823;
assign v_13826 = v_12771;
assign v_13828 = v_13825 & v_13827;
assign v_13830 = v_13750 & v_13829;
assign v_13832 = v_12767;
assign v_13834 = v_13831 & v_13833;
assign v_13836 = v_13747 & v_13835;
assign v_13838 = v_12763;
assign v_13840 = v_13837 & v_13839;
assign v_13842 = v_13744 & v_13841;
assign v_13844 = v_12759;
assign v_13846 = v_13843 & v_13845;
assign v_13848 = v_13741 & v_13847;
assign v_13850 = v_12755;
assign v_13852 = v_13849 & v_13851;
assign v_13854 = v_13738 & v_13853;
assign v_13856 = v_1075;
assign v_13858 = v_13855 & v_13857;
assign v_13860 = v_13735 & v_13859;
assign v_13862 = v_1071;
assign v_13864 = v_13861 & v_13863;
assign v_13866 = v_13732 & v_13865;
assign v_13868 = v_1067;
assign v_13870 = v_13867 & v_13869;
assign v_13872 = v_13729 & v_13871;
assign v_13874 = v_1063;
assign v_13876 = v_13873 & v_13875;
assign v_13877 = v_13876;
assign v_13879 = v_12803;
assign v_13880 = v_1128;
assign v_13881 = v_13880;
assign v_13882 = v_13879 & v_13881;
assign v_13883 = v_13882;
assign v_13884 = v_13774 & v_13883;
assign v_13886 = v_13784 & v_13885;
assign v_13887 = v_13773 & v_13883;
assign v_13889 = v_13771 & v_13888;
assign v_13891 = v_13790 & v_13890;
assign v_13892 = v_13770 & v_13888;
assign v_13894 = v_13768 & v_13893;
assign v_13896 = v_13796 & v_13895;
assign v_13897 = v_13767 & v_13893;
assign v_13899 = v_13765 & v_13898;
assign v_13901 = v_13802 & v_13900;
assign v_13902 = v_13764 & v_13898;
assign v_13904 = v_13762 & v_13903;
assign v_13906 = v_13808 & v_13905;
assign v_13907 = v_13761 & v_13903;
assign v_13909 = v_13759 & v_13908;
assign v_13911 = v_13814 & v_13910;
assign v_13912 = v_13758 & v_13908;
assign v_13914 = v_13756 & v_13913;
assign v_13916 = v_13820 & v_13915;
assign v_13917 = v_13755 & v_13913;
assign v_13919 = v_13753 & v_13918;
assign v_13921 = v_13826 & v_13920;
assign v_13922 = v_13752 & v_13918;
assign v_13924 = v_13750 & v_13923;
assign v_13926 = v_13832 & v_13925;
assign v_13927 = v_13749 & v_13923;
assign v_13929 = v_13747 & v_13928;
assign v_13931 = v_13838 & v_13930;
assign v_13932 = v_13746 & v_13928;
assign v_13934 = v_13744 & v_13933;
assign v_13936 = v_13844 & v_13935;
assign v_13937 = v_13743 & v_13933;
assign v_13939 = v_13741 & v_13938;
assign v_13941 = v_13850 & v_13940;
assign v_13942 = v_13740 & v_13938;
assign v_13944 = v_13738 & v_13943;
assign v_13946 = v_13856 & v_13945;
assign v_13947 = v_13737 & v_13943;
assign v_13949 = v_13735 & v_13948;
assign v_13951 = v_13862 & v_13950;
assign v_13952 = v_13734 & v_13948;
assign v_13954 = v_13732 & v_13953;
assign v_13956 = v_13868 & v_13955;
assign v_13957 = v_13731 & v_13953;
assign v_13959 = v_13729 & v_13958;
assign v_13961 = v_13874 & v_13960;
assign v_13962 = v_13728 & v_13958;
assign v_13964 = v_13963;
assign v_13966 = v_13878 & v_13965;
assign v_13967 = v_13966;
assign v_13969 = v_13968;
assign v_13971 = ~v_1323;
assign v_13972 = ~v_12740;
assign v_13973 = v_12740;
assign v_13974 = ~v_1327;
assign v_13975 = ~v_12744;
assign v_13976 = v_12744;
assign v_13977 = ~v_1331;
assign v_13978 = ~v_12748;
assign v_13979 = v_12748;
assign v_13980 = ~v_1335;
assign v_13981 = ~v_12752;
assign v_13982 = v_12752;
assign v_13983 = ~v_12755;
assign v_13984 = ~v_1340;
assign v_13985 = v_1340;
assign v_13986 = ~v_12759;
assign v_13987 = ~v_1344;
assign v_13988 = v_1344;
assign v_13989 = ~v_12763;
assign v_13990 = ~v_1348;
assign v_13991 = v_1348;
assign v_13992 = ~v_12767;
assign v_13993 = ~v_1352;
assign v_13994 = v_1352;
assign v_13995 = ~v_12771;
assign v_13996 = ~v_1356;
assign v_13997 = v_1356;
assign v_13998 = ~v_12775;
assign v_13999 = ~v_1360;
assign v_14000 = v_1360;
assign v_14001 = ~v_12779;
assign v_14002 = ~v_1364;
assign v_14003 = v_1364;
assign v_14004 = ~v_12783;
assign v_14005 = ~v_1368;
assign v_14006 = v_1368;
assign v_14007 = ~v_12787;
assign v_14008 = ~v_1372;
assign v_14009 = v_1372;
assign v_14010 = ~v_12791;
assign v_14011 = ~v_1376;
assign v_14012 = v_1376;
assign v_14013 = ~v_12795;
assign v_14014 = ~v_1380;
assign v_14015 = v_1380;
assign v_14016 = ~v_12799;
assign v_14017 = ~v_1384;
assign v_14018 = v_1384;
assign v_14019 = ~v_12803;
assign v_14020 = ~v_1388;
assign v_14021 = v_14020;
assign v_14023 = v_14022;
assign v_14025 = v_14017 & v_14024;
assign v_14027 = v_12799;
assign v_14029 = v_14026 & v_14028;
assign v_14031 = v_14014 & v_14030;
assign v_14033 = v_12795;
assign v_14035 = v_14032 & v_14034;
assign v_14037 = v_14011 & v_14036;
assign v_14039 = v_12791;
assign v_14041 = v_14038 & v_14040;
assign v_14043 = v_14008 & v_14042;
assign v_14045 = v_12787;
assign v_14047 = v_14044 & v_14046;
assign v_14049 = v_14005 & v_14048;
assign v_14051 = v_12783;
assign v_14053 = v_14050 & v_14052;
assign v_14055 = v_14002 & v_14054;
assign v_14057 = v_12779;
assign v_14059 = v_14056 & v_14058;
assign v_14061 = v_13999 & v_14060;
assign v_14063 = v_12775;
assign v_14065 = v_14062 & v_14064;
assign v_14067 = v_13996 & v_14066;
assign v_14069 = v_12771;
assign v_14071 = v_14068 & v_14070;
assign v_14073 = v_13993 & v_14072;
assign v_14075 = v_12767;
assign v_14077 = v_14074 & v_14076;
assign v_14079 = v_13990 & v_14078;
assign v_14081 = v_12763;
assign v_14083 = v_14080 & v_14082;
assign v_14085 = v_13987 & v_14084;
assign v_14087 = v_12759;
assign v_14089 = v_14086 & v_14088;
assign v_14091 = v_13984 & v_14090;
assign v_14093 = v_12755;
assign v_14095 = v_14092 & v_14094;
assign v_14097 = v_13981 & v_14096;
assign v_14099 = v_1335;
assign v_14101 = v_14098 & v_14100;
assign v_14103 = v_13978 & v_14102;
assign v_14105 = v_1331;
assign v_14107 = v_14104 & v_14106;
assign v_14109 = v_13975 & v_14108;
assign v_14111 = v_1327;
assign v_14113 = v_14110 & v_14112;
assign v_14115 = v_13972 & v_14114;
assign v_14117 = v_1323;
assign v_14119 = v_14116 & v_14118;
assign v_14120 = v_14119;
assign v_14122 = v_12803;
assign v_14123 = v_1388;
assign v_14124 = v_14123;
assign v_14125 = v_14122 & v_14124;
assign v_14126 = v_14125;
assign v_14127 = v_14017 & v_14126;
assign v_14129 = v_14027 & v_14128;
assign v_14130 = v_14016 & v_14126;
assign v_14132 = v_14014 & v_14131;
assign v_14134 = v_14033 & v_14133;
assign v_14135 = v_14013 & v_14131;
assign v_14137 = v_14011 & v_14136;
assign v_14139 = v_14039 & v_14138;
assign v_14140 = v_14010 & v_14136;
assign v_14142 = v_14008 & v_14141;
assign v_14144 = v_14045 & v_14143;
assign v_14145 = v_14007 & v_14141;
assign v_14147 = v_14005 & v_14146;
assign v_14149 = v_14051 & v_14148;
assign v_14150 = v_14004 & v_14146;
assign v_14152 = v_14002 & v_14151;
assign v_14154 = v_14057 & v_14153;
assign v_14155 = v_14001 & v_14151;
assign v_14157 = v_13999 & v_14156;
assign v_14159 = v_14063 & v_14158;
assign v_14160 = v_13998 & v_14156;
assign v_14162 = v_13996 & v_14161;
assign v_14164 = v_14069 & v_14163;
assign v_14165 = v_13995 & v_14161;
assign v_14167 = v_13993 & v_14166;
assign v_14169 = v_14075 & v_14168;
assign v_14170 = v_13992 & v_14166;
assign v_14172 = v_13990 & v_14171;
assign v_14174 = v_14081 & v_14173;
assign v_14175 = v_13989 & v_14171;
assign v_14177 = v_13987 & v_14176;
assign v_14179 = v_14087 & v_14178;
assign v_14180 = v_13986 & v_14176;
assign v_14182 = v_13984 & v_14181;
assign v_14184 = v_14093 & v_14183;
assign v_14185 = v_13983 & v_14181;
assign v_14187 = v_13981 & v_14186;
assign v_14189 = v_14099 & v_14188;
assign v_14190 = v_13980 & v_14186;
assign v_14192 = v_13978 & v_14191;
assign v_14194 = v_14105 & v_14193;
assign v_14195 = v_13977 & v_14191;
assign v_14197 = v_13975 & v_14196;
assign v_14199 = v_14111 & v_14198;
assign v_14200 = v_13974 & v_14196;
assign v_14202 = v_13972 & v_14201;
assign v_14204 = v_14117 & v_14203;
assign v_14205 = v_13971 & v_14201;
assign v_14207 = v_14206;
assign v_14209 = v_14121 & v_14208;
assign v_14210 = v_14209;
assign v_14212 = v_14211;
assign v_14214 = ~v_1583;
assign v_14215 = ~v_12740;
assign v_14216 = v_12740;
assign v_14217 = ~v_1587;
assign v_14218 = ~v_12744;
assign v_14219 = v_12744;
assign v_14220 = ~v_1591;
assign v_14221 = ~v_12748;
assign v_14222 = v_12748;
assign v_14223 = ~v_1595;
assign v_14224 = ~v_12752;
assign v_14225 = v_12752;
assign v_14226 = ~v_12755;
assign v_14227 = ~v_1600;
assign v_14228 = v_1600;
assign v_14229 = ~v_12759;
assign v_14230 = ~v_1604;
assign v_14231 = v_1604;
assign v_14232 = ~v_12763;
assign v_14233 = ~v_1608;
assign v_14234 = v_1608;
assign v_14235 = ~v_12767;
assign v_14236 = ~v_1612;
assign v_14237 = v_1612;
assign v_14238 = ~v_12771;
assign v_14239 = ~v_1616;
assign v_14240 = v_1616;
assign v_14241 = ~v_12775;
assign v_14242 = ~v_1620;
assign v_14243 = v_1620;
assign v_14244 = ~v_12779;
assign v_14245 = ~v_1624;
assign v_14246 = v_1624;
assign v_14247 = ~v_12783;
assign v_14248 = ~v_1628;
assign v_14249 = v_1628;
assign v_14250 = ~v_12787;
assign v_14251 = ~v_1632;
assign v_14252 = v_1632;
assign v_14253 = ~v_12791;
assign v_14254 = ~v_1636;
assign v_14255 = v_1636;
assign v_14256 = ~v_12795;
assign v_14257 = ~v_1640;
assign v_14258 = v_1640;
assign v_14259 = ~v_12799;
assign v_14260 = ~v_1644;
assign v_14261 = v_1644;
assign v_14262 = ~v_12803;
assign v_14263 = ~v_1648;
assign v_14264 = v_14263;
assign v_14266 = v_14265;
assign v_14268 = v_14260 & v_14267;
assign v_14270 = v_12799;
assign v_14272 = v_14269 & v_14271;
assign v_14274 = v_14257 & v_14273;
assign v_14276 = v_12795;
assign v_14278 = v_14275 & v_14277;
assign v_14280 = v_14254 & v_14279;
assign v_14282 = v_12791;
assign v_14284 = v_14281 & v_14283;
assign v_14286 = v_14251 & v_14285;
assign v_14288 = v_12787;
assign v_14290 = v_14287 & v_14289;
assign v_14292 = v_14248 & v_14291;
assign v_14294 = v_12783;
assign v_14296 = v_14293 & v_14295;
assign v_14298 = v_14245 & v_14297;
assign v_14300 = v_12779;
assign v_14302 = v_14299 & v_14301;
assign v_14304 = v_14242 & v_14303;
assign v_14306 = v_12775;
assign v_14308 = v_14305 & v_14307;
assign v_14310 = v_14239 & v_14309;
assign v_14312 = v_12771;
assign v_14314 = v_14311 & v_14313;
assign v_14316 = v_14236 & v_14315;
assign v_14318 = v_12767;
assign v_14320 = v_14317 & v_14319;
assign v_14322 = v_14233 & v_14321;
assign v_14324 = v_12763;
assign v_14326 = v_14323 & v_14325;
assign v_14328 = v_14230 & v_14327;
assign v_14330 = v_12759;
assign v_14332 = v_14329 & v_14331;
assign v_14334 = v_14227 & v_14333;
assign v_14336 = v_12755;
assign v_14338 = v_14335 & v_14337;
assign v_14340 = v_14224 & v_14339;
assign v_14342 = v_1595;
assign v_14344 = v_14341 & v_14343;
assign v_14346 = v_14221 & v_14345;
assign v_14348 = v_1591;
assign v_14350 = v_14347 & v_14349;
assign v_14352 = v_14218 & v_14351;
assign v_14354 = v_1587;
assign v_14356 = v_14353 & v_14355;
assign v_14358 = v_14215 & v_14357;
assign v_14360 = v_1583;
assign v_14362 = v_14359 & v_14361;
assign v_14363 = v_14362;
assign v_14365 = v_12803;
assign v_14366 = v_1648;
assign v_14367 = v_14366;
assign v_14368 = v_14365 & v_14367;
assign v_14369 = v_14368;
assign v_14370 = v_14260 & v_14369;
assign v_14372 = v_14270 & v_14371;
assign v_14373 = v_14259 & v_14369;
assign v_14375 = v_14257 & v_14374;
assign v_14377 = v_14276 & v_14376;
assign v_14378 = v_14256 & v_14374;
assign v_14380 = v_14254 & v_14379;
assign v_14382 = v_14282 & v_14381;
assign v_14383 = v_14253 & v_14379;
assign v_14385 = v_14251 & v_14384;
assign v_14387 = v_14288 & v_14386;
assign v_14388 = v_14250 & v_14384;
assign v_14390 = v_14248 & v_14389;
assign v_14392 = v_14294 & v_14391;
assign v_14393 = v_14247 & v_14389;
assign v_14395 = v_14245 & v_14394;
assign v_14397 = v_14300 & v_14396;
assign v_14398 = v_14244 & v_14394;
assign v_14400 = v_14242 & v_14399;
assign v_14402 = v_14306 & v_14401;
assign v_14403 = v_14241 & v_14399;
assign v_14405 = v_14239 & v_14404;
assign v_14407 = v_14312 & v_14406;
assign v_14408 = v_14238 & v_14404;
assign v_14410 = v_14236 & v_14409;
assign v_14412 = v_14318 & v_14411;
assign v_14413 = v_14235 & v_14409;
assign v_14415 = v_14233 & v_14414;
assign v_14417 = v_14324 & v_14416;
assign v_14418 = v_14232 & v_14414;
assign v_14420 = v_14230 & v_14419;
assign v_14422 = v_14330 & v_14421;
assign v_14423 = v_14229 & v_14419;
assign v_14425 = v_14227 & v_14424;
assign v_14427 = v_14336 & v_14426;
assign v_14428 = v_14226 & v_14424;
assign v_14430 = v_14224 & v_14429;
assign v_14432 = v_14342 & v_14431;
assign v_14433 = v_14223 & v_14429;
assign v_14435 = v_14221 & v_14434;
assign v_14437 = v_14348 & v_14436;
assign v_14438 = v_14220 & v_14434;
assign v_14440 = v_14218 & v_14439;
assign v_14442 = v_14354 & v_14441;
assign v_14443 = v_14217 & v_14439;
assign v_14445 = v_14215 & v_14444;
assign v_14447 = v_14360 & v_14446;
assign v_14448 = v_14214 & v_14444;
assign v_14450 = v_14449;
assign v_14452 = v_14364 & v_14451;
assign v_14453 = v_14452;
assign v_14455 = v_14454;
assign v_14457 = ~v_1843;
assign v_14458 = ~v_12740;
assign v_14459 = v_12740;
assign v_14460 = ~v_1847;
assign v_14461 = ~v_12744;
assign v_14462 = v_12744;
assign v_14463 = ~v_1851;
assign v_14464 = ~v_12748;
assign v_14465 = v_12748;
assign v_14466 = ~v_1855;
assign v_14467 = ~v_12752;
assign v_14468 = v_12752;
assign v_14469 = ~v_12755;
assign v_14470 = ~v_1860;
assign v_14471 = v_1860;
assign v_14472 = ~v_12759;
assign v_14473 = ~v_1864;
assign v_14474 = v_1864;
assign v_14475 = ~v_12763;
assign v_14476 = ~v_1868;
assign v_14477 = v_1868;
assign v_14478 = ~v_12767;
assign v_14479 = ~v_1872;
assign v_14480 = v_1872;
assign v_14481 = ~v_12771;
assign v_14482 = ~v_1876;
assign v_14483 = v_1876;
assign v_14484 = ~v_12775;
assign v_14485 = ~v_1880;
assign v_14486 = v_1880;
assign v_14487 = ~v_12779;
assign v_14488 = ~v_1884;
assign v_14489 = v_1884;
assign v_14490 = ~v_12783;
assign v_14491 = ~v_1888;
assign v_14492 = v_1888;
assign v_14493 = ~v_12787;
assign v_14494 = ~v_1892;
assign v_14495 = v_1892;
assign v_14496 = ~v_12791;
assign v_14497 = ~v_1896;
assign v_14498 = v_1896;
assign v_14499 = ~v_12795;
assign v_14500 = ~v_1900;
assign v_14501 = v_1900;
assign v_14502 = ~v_12799;
assign v_14503 = ~v_1904;
assign v_14504 = v_1904;
assign v_14505 = ~v_12803;
assign v_14506 = ~v_1908;
assign v_14507 = v_14506;
assign v_14509 = v_14508;
assign v_14511 = v_14503 & v_14510;
assign v_14513 = v_12799;
assign v_14515 = v_14512 & v_14514;
assign v_14517 = v_14500 & v_14516;
assign v_14519 = v_12795;
assign v_14521 = v_14518 & v_14520;
assign v_14523 = v_14497 & v_14522;
assign v_14525 = v_12791;
assign v_14527 = v_14524 & v_14526;
assign v_14529 = v_14494 & v_14528;
assign v_14531 = v_12787;
assign v_14533 = v_14530 & v_14532;
assign v_14535 = v_14491 & v_14534;
assign v_14537 = v_12783;
assign v_14539 = v_14536 & v_14538;
assign v_14541 = v_14488 & v_14540;
assign v_14543 = v_12779;
assign v_14545 = v_14542 & v_14544;
assign v_14547 = v_14485 & v_14546;
assign v_14549 = v_12775;
assign v_14551 = v_14548 & v_14550;
assign v_14553 = v_14482 & v_14552;
assign v_14555 = v_12771;
assign v_14557 = v_14554 & v_14556;
assign v_14559 = v_14479 & v_14558;
assign v_14561 = v_12767;
assign v_14563 = v_14560 & v_14562;
assign v_14565 = v_14476 & v_14564;
assign v_14567 = v_12763;
assign v_14569 = v_14566 & v_14568;
assign v_14571 = v_14473 & v_14570;
assign v_14573 = v_12759;
assign v_14575 = v_14572 & v_14574;
assign v_14577 = v_14470 & v_14576;
assign v_14579 = v_12755;
assign v_14581 = v_14578 & v_14580;
assign v_14583 = v_14467 & v_14582;
assign v_14585 = v_1855;
assign v_14587 = v_14584 & v_14586;
assign v_14589 = v_14464 & v_14588;
assign v_14591 = v_1851;
assign v_14593 = v_14590 & v_14592;
assign v_14595 = v_14461 & v_14594;
assign v_14597 = v_1847;
assign v_14599 = v_14596 & v_14598;
assign v_14601 = v_14458 & v_14600;
assign v_14603 = v_1843;
assign v_14605 = v_14602 & v_14604;
assign v_14606 = v_14605;
assign v_14608 = v_12803;
assign v_14609 = v_1908;
assign v_14610 = v_14609;
assign v_14611 = v_14608 & v_14610;
assign v_14612 = v_14611;
assign v_14613 = v_14503 & v_14612;
assign v_14615 = v_14513 & v_14614;
assign v_14616 = v_14502 & v_14612;
assign v_14618 = v_14500 & v_14617;
assign v_14620 = v_14519 & v_14619;
assign v_14621 = v_14499 & v_14617;
assign v_14623 = v_14497 & v_14622;
assign v_14625 = v_14525 & v_14624;
assign v_14626 = v_14496 & v_14622;
assign v_14628 = v_14494 & v_14627;
assign v_14630 = v_14531 & v_14629;
assign v_14631 = v_14493 & v_14627;
assign v_14633 = v_14491 & v_14632;
assign v_14635 = v_14537 & v_14634;
assign v_14636 = v_14490 & v_14632;
assign v_14638 = v_14488 & v_14637;
assign v_14640 = v_14543 & v_14639;
assign v_14641 = v_14487 & v_14637;
assign v_14643 = v_14485 & v_14642;
assign v_14645 = v_14549 & v_14644;
assign v_14646 = v_14484 & v_14642;
assign v_14648 = v_14482 & v_14647;
assign v_14650 = v_14555 & v_14649;
assign v_14651 = v_14481 & v_14647;
assign v_14653 = v_14479 & v_14652;
assign v_14655 = v_14561 & v_14654;
assign v_14656 = v_14478 & v_14652;
assign v_14658 = v_14476 & v_14657;
assign v_14660 = v_14567 & v_14659;
assign v_14661 = v_14475 & v_14657;
assign v_14663 = v_14473 & v_14662;
assign v_14665 = v_14573 & v_14664;
assign v_14666 = v_14472 & v_14662;
assign v_14668 = v_14470 & v_14667;
assign v_14670 = v_14579 & v_14669;
assign v_14671 = v_14469 & v_14667;
assign v_14673 = v_14467 & v_14672;
assign v_14675 = v_14585 & v_14674;
assign v_14676 = v_14466 & v_14672;
assign v_14678 = v_14464 & v_14677;
assign v_14680 = v_14591 & v_14679;
assign v_14681 = v_14463 & v_14677;
assign v_14683 = v_14461 & v_14682;
assign v_14685 = v_14597 & v_14684;
assign v_14686 = v_14460 & v_14682;
assign v_14688 = v_14458 & v_14687;
assign v_14690 = v_14603 & v_14689;
assign v_14691 = v_14457 & v_14687;
assign v_14693 = v_14692;
assign v_14695 = v_14607 & v_14694;
assign v_14696 = v_14695;
assign v_14698 = v_14697;
assign v_14700 = ~v_2103;
assign v_14701 = ~v_12740;
assign v_14702 = v_12740;
assign v_14703 = ~v_2107;
assign v_14704 = ~v_12744;
assign v_14705 = v_12744;
assign v_14706 = ~v_2111;
assign v_14707 = ~v_12748;
assign v_14708 = v_12748;
assign v_14709 = ~v_2115;
assign v_14710 = ~v_12752;
assign v_14711 = v_12752;
assign v_14712 = ~v_12755;
assign v_14713 = ~v_2120;
assign v_14714 = v_2120;
assign v_14715 = ~v_12759;
assign v_14716 = ~v_2124;
assign v_14717 = v_2124;
assign v_14718 = ~v_12763;
assign v_14719 = ~v_2128;
assign v_14720 = v_2128;
assign v_14721 = ~v_12767;
assign v_14722 = ~v_2132;
assign v_14723 = v_2132;
assign v_14724 = ~v_12771;
assign v_14725 = ~v_2136;
assign v_14726 = v_2136;
assign v_14727 = ~v_12775;
assign v_14728 = ~v_2140;
assign v_14729 = v_2140;
assign v_14730 = ~v_12779;
assign v_14731 = ~v_2144;
assign v_14732 = v_2144;
assign v_14733 = ~v_12783;
assign v_14734 = ~v_2148;
assign v_14735 = v_2148;
assign v_14736 = ~v_12787;
assign v_14737 = ~v_2152;
assign v_14738 = v_2152;
assign v_14739 = ~v_12791;
assign v_14740 = ~v_2156;
assign v_14741 = v_2156;
assign v_14742 = ~v_12795;
assign v_14743 = ~v_2160;
assign v_14744 = v_2160;
assign v_14745 = ~v_12799;
assign v_14746 = ~v_2164;
assign v_14747 = v_2164;
assign v_14748 = ~v_12803;
assign v_14749 = ~v_2168;
assign v_14750 = v_14749;
assign v_14752 = v_14751;
assign v_14754 = v_14746 & v_14753;
assign v_14756 = v_12799;
assign v_14758 = v_14755 & v_14757;
assign v_14760 = v_14743 & v_14759;
assign v_14762 = v_12795;
assign v_14764 = v_14761 & v_14763;
assign v_14766 = v_14740 & v_14765;
assign v_14768 = v_12791;
assign v_14770 = v_14767 & v_14769;
assign v_14772 = v_14737 & v_14771;
assign v_14774 = v_12787;
assign v_14776 = v_14773 & v_14775;
assign v_14778 = v_14734 & v_14777;
assign v_14780 = v_12783;
assign v_14782 = v_14779 & v_14781;
assign v_14784 = v_14731 & v_14783;
assign v_14786 = v_12779;
assign v_14788 = v_14785 & v_14787;
assign v_14790 = v_14728 & v_14789;
assign v_14792 = v_12775;
assign v_14794 = v_14791 & v_14793;
assign v_14796 = v_14725 & v_14795;
assign v_14798 = v_12771;
assign v_14800 = v_14797 & v_14799;
assign v_14802 = v_14722 & v_14801;
assign v_14804 = v_12767;
assign v_14806 = v_14803 & v_14805;
assign v_14808 = v_14719 & v_14807;
assign v_14810 = v_12763;
assign v_14812 = v_14809 & v_14811;
assign v_14814 = v_14716 & v_14813;
assign v_14816 = v_12759;
assign v_14818 = v_14815 & v_14817;
assign v_14820 = v_14713 & v_14819;
assign v_14822 = v_12755;
assign v_14824 = v_14821 & v_14823;
assign v_14826 = v_14710 & v_14825;
assign v_14828 = v_2115;
assign v_14830 = v_14827 & v_14829;
assign v_14832 = v_14707 & v_14831;
assign v_14834 = v_2111;
assign v_14836 = v_14833 & v_14835;
assign v_14838 = v_14704 & v_14837;
assign v_14840 = v_2107;
assign v_14842 = v_14839 & v_14841;
assign v_14844 = v_14701 & v_14843;
assign v_14846 = v_2103;
assign v_14848 = v_14845 & v_14847;
assign v_14849 = v_14848;
assign v_14851 = v_12803;
assign v_14852 = v_2168;
assign v_14853 = v_14852;
assign v_14854 = v_14851 & v_14853;
assign v_14855 = v_14854;
assign v_14856 = v_14746 & v_14855;
assign v_14858 = v_14756 & v_14857;
assign v_14859 = v_14745 & v_14855;
assign v_14861 = v_14743 & v_14860;
assign v_14863 = v_14762 & v_14862;
assign v_14864 = v_14742 & v_14860;
assign v_14866 = v_14740 & v_14865;
assign v_14868 = v_14768 & v_14867;
assign v_14869 = v_14739 & v_14865;
assign v_14871 = v_14737 & v_14870;
assign v_14873 = v_14774 & v_14872;
assign v_14874 = v_14736 & v_14870;
assign v_14876 = v_14734 & v_14875;
assign v_14878 = v_14780 & v_14877;
assign v_14879 = v_14733 & v_14875;
assign v_14881 = v_14731 & v_14880;
assign v_14883 = v_14786 & v_14882;
assign v_14884 = v_14730 & v_14880;
assign v_14886 = v_14728 & v_14885;
assign v_14888 = v_14792 & v_14887;
assign v_14889 = v_14727 & v_14885;
assign v_14891 = v_14725 & v_14890;
assign v_14893 = v_14798 & v_14892;
assign v_14894 = v_14724 & v_14890;
assign v_14896 = v_14722 & v_14895;
assign v_14898 = v_14804 & v_14897;
assign v_14899 = v_14721 & v_14895;
assign v_14901 = v_14719 & v_14900;
assign v_14903 = v_14810 & v_14902;
assign v_14904 = v_14718 & v_14900;
assign v_14906 = v_14716 & v_14905;
assign v_14908 = v_14816 & v_14907;
assign v_14909 = v_14715 & v_14905;
assign v_14911 = v_14713 & v_14910;
assign v_14913 = v_14822 & v_14912;
assign v_14914 = v_14712 & v_14910;
assign v_14916 = v_14710 & v_14915;
assign v_14918 = v_14828 & v_14917;
assign v_14919 = v_14709 & v_14915;
assign v_14921 = v_14707 & v_14920;
assign v_14923 = v_14834 & v_14922;
assign v_14924 = v_14706 & v_14920;
assign v_14926 = v_14704 & v_14925;
assign v_14928 = v_14840 & v_14927;
assign v_14929 = v_14703 & v_14925;
assign v_14931 = v_14701 & v_14930;
assign v_14933 = v_14846 & v_14932;
assign v_14934 = v_14700 & v_14930;
assign v_14936 = v_14935;
assign v_14938 = v_14850 & v_14937;
assign v_14939 = v_14938;
assign v_14941 = v_14940;
assign v_14943 = ~v_2363;
assign v_14944 = ~v_12740;
assign v_14945 = v_12740;
assign v_14946 = ~v_2367;
assign v_14947 = ~v_12744;
assign v_14948 = v_12744;
assign v_14949 = ~v_2371;
assign v_14950 = ~v_12748;
assign v_14951 = v_12748;
assign v_14952 = ~v_2375;
assign v_14953 = ~v_12752;
assign v_14954 = v_12752;
assign v_14955 = ~v_12755;
assign v_14956 = ~v_2380;
assign v_14957 = v_2380;
assign v_14958 = ~v_12759;
assign v_14959 = ~v_2384;
assign v_14960 = v_2384;
assign v_14961 = ~v_12763;
assign v_14962 = ~v_2388;
assign v_14963 = v_2388;
assign v_14964 = ~v_12767;
assign v_14965 = ~v_2392;
assign v_14966 = v_2392;
assign v_14967 = ~v_12771;
assign v_14968 = ~v_2396;
assign v_14969 = v_2396;
assign v_14970 = ~v_12775;
assign v_14971 = ~v_2400;
assign v_14972 = v_2400;
assign v_14973 = ~v_12779;
assign v_14974 = ~v_2404;
assign v_14975 = v_2404;
assign v_14976 = ~v_12783;
assign v_14977 = ~v_2408;
assign v_14978 = v_2408;
assign v_14979 = ~v_12787;
assign v_14980 = ~v_2412;
assign v_14981 = v_2412;
assign v_14982 = ~v_12791;
assign v_14983 = ~v_2416;
assign v_14984 = v_2416;
assign v_14985 = ~v_12795;
assign v_14986 = ~v_2420;
assign v_14987 = v_2420;
assign v_14988 = ~v_12799;
assign v_14989 = ~v_2424;
assign v_14990 = v_2424;
assign v_14991 = ~v_12803;
assign v_14992 = ~v_2428;
assign v_14993 = v_14992;
assign v_14995 = v_14994;
assign v_14997 = v_14989 & v_14996;
assign v_14999 = v_12799;
assign v_15001 = v_14998 & v_15000;
assign v_15003 = v_14986 & v_15002;
assign v_15005 = v_12795;
assign v_15007 = v_15004 & v_15006;
assign v_15009 = v_14983 & v_15008;
assign v_15011 = v_12791;
assign v_15013 = v_15010 & v_15012;
assign v_15015 = v_14980 & v_15014;
assign v_15017 = v_12787;
assign v_15019 = v_15016 & v_15018;
assign v_15021 = v_14977 & v_15020;
assign v_15023 = v_12783;
assign v_15025 = v_15022 & v_15024;
assign v_15027 = v_14974 & v_15026;
assign v_15029 = v_12779;
assign v_15031 = v_15028 & v_15030;
assign v_15033 = v_14971 & v_15032;
assign v_15035 = v_12775;
assign v_15037 = v_15034 & v_15036;
assign v_15039 = v_14968 & v_15038;
assign v_15041 = v_12771;
assign v_15043 = v_15040 & v_15042;
assign v_15045 = v_14965 & v_15044;
assign v_15047 = v_12767;
assign v_15049 = v_15046 & v_15048;
assign v_15051 = v_14962 & v_15050;
assign v_15053 = v_12763;
assign v_15055 = v_15052 & v_15054;
assign v_15057 = v_14959 & v_15056;
assign v_15059 = v_12759;
assign v_15061 = v_15058 & v_15060;
assign v_15063 = v_14956 & v_15062;
assign v_15065 = v_12755;
assign v_15067 = v_15064 & v_15066;
assign v_15069 = v_14953 & v_15068;
assign v_15071 = v_2375;
assign v_15073 = v_15070 & v_15072;
assign v_15075 = v_14950 & v_15074;
assign v_15077 = v_2371;
assign v_15079 = v_15076 & v_15078;
assign v_15081 = v_14947 & v_15080;
assign v_15083 = v_2367;
assign v_15085 = v_15082 & v_15084;
assign v_15087 = v_14944 & v_15086;
assign v_15089 = v_2363;
assign v_15091 = v_15088 & v_15090;
assign v_15092 = v_15091;
assign v_15094 = v_12803;
assign v_15095 = v_2428;
assign v_15096 = v_15095;
assign v_15097 = v_15094 & v_15096;
assign v_15098 = v_15097;
assign v_15099 = v_14989 & v_15098;
assign v_15101 = v_14999 & v_15100;
assign v_15102 = v_14988 & v_15098;
assign v_15104 = v_14986 & v_15103;
assign v_15106 = v_15005 & v_15105;
assign v_15107 = v_14985 & v_15103;
assign v_15109 = v_14983 & v_15108;
assign v_15111 = v_15011 & v_15110;
assign v_15112 = v_14982 & v_15108;
assign v_15114 = v_14980 & v_15113;
assign v_15116 = v_15017 & v_15115;
assign v_15117 = v_14979 & v_15113;
assign v_15119 = v_14977 & v_15118;
assign v_15121 = v_15023 & v_15120;
assign v_15122 = v_14976 & v_15118;
assign v_15124 = v_14974 & v_15123;
assign v_15126 = v_15029 & v_15125;
assign v_15127 = v_14973 & v_15123;
assign v_15129 = v_14971 & v_15128;
assign v_15131 = v_15035 & v_15130;
assign v_15132 = v_14970 & v_15128;
assign v_15134 = v_14968 & v_15133;
assign v_15136 = v_15041 & v_15135;
assign v_15137 = v_14967 & v_15133;
assign v_15139 = v_14965 & v_15138;
assign v_15141 = v_15047 & v_15140;
assign v_15142 = v_14964 & v_15138;
assign v_15144 = v_14962 & v_15143;
assign v_15146 = v_15053 & v_15145;
assign v_15147 = v_14961 & v_15143;
assign v_15149 = v_14959 & v_15148;
assign v_15151 = v_15059 & v_15150;
assign v_15152 = v_14958 & v_15148;
assign v_15154 = v_14956 & v_15153;
assign v_15156 = v_15065 & v_15155;
assign v_15157 = v_14955 & v_15153;
assign v_15159 = v_14953 & v_15158;
assign v_15161 = v_15071 & v_15160;
assign v_15162 = v_14952 & v_15158;
assign v_15164 = v_14950 & v_15163;
assign v_15166 = v_15077 & v_15165;
assign v_15167 = v_14949 & v_15163;
assign v_15169 = v_14947 & v_15168;
assign v_15171 = v_15083 & v_15170;
assign v_15172 = v_14946 & v_15168;
assign v_15174 = v_14944 & v_15173;
assign v_15176 = v_15089 & v_15175;
assign v_15177 = v_14943 & v_15173;
assign v_15179 = v_15178;
assign v_15181 = v_15093 & v_15180;
assign v_15182 = v_15181;
assign v_15184 = v_15183;
assign v_15186 = ~v_2623;
assign v_15187 = ~v_12740;
assign v_15188 = v_12740;
assign v_15189 = ~v_2627;
assign v_15190 = ~v_12744;
assign v_15191 = v_12744;
assign v_15192 = ~v_2631;
assign v_15193 = ~v_12748;
assign v_15194 = v_12748;
assign v_15195 = ~v_2635;
assign v_15196 = ~v_12752;
assign v_15197 = v_12752;
assign v_15198 = ~v_12755;
assign v_15199 = ~v_2640;
assign v_15200 = v_2640;
assign v_15201 = ~v_12759;
assign v_15202 = ~v_2644;
assign v_15203 = v_2644;
assign v_15204 = ~v_12763;
assign v_15205 = ~v_2648;
assign v_15206 = v_2648;
assign v_15207 = ~v_12767;
assign v_15208 = ~v_2652;
assign v_15209 = v_2652;
assign v_15210 = ~v_12771;
assign v_15211 = ~v_2656;
assign v_15212 = v_2656;
assign v_15213 = ~v_12775;
assign v_15214 = ~v_2660;
assign v_15215 = v_2660;
assign v_15216 = ~v_12779;
assign v_15217 = ~v_2664;
assign v_15218 = v_2664;
assign v_15219 = ~v_12783;
assign v_15220 = ~v_2668;
assign v_15221 = v_2668;
assign v_15222 = ~v_12787;
assign v_15223 = ~v_2672;
assign v_15224 = v_2672;
assign v_15225 = ~v_12791;
assign v_15226 = ~v_2676;
assign v_15227 = v_2676;
assign v_15228 = ~v_12795;
assign v_15229 = ~v_2680;
assign v_15230 = v_2680;
assign v_15231 = ~v_12799;
assign v_15232 = ~v_2684;
assign v_15233 = v_2684;
assign v_15234 = ~v_12803;
assign v_15235 = ~v_2688;
assign v_15236 = v_15235;
assign v_15238 = v_15237;
assign v_15240 = v_15232 & v_15239;
assign v_15242 = v_12799;
assign v_15244 = v_15241 & v_15243;
assign v_15246 = v_15229 & v_15245;
assign v_15248 = v_12795;
assign v_15250 = v_15247 & v_15249;
assign v_15252 = v_15226 & v_15251;
assign v_15254 = v_12791;
assign v_15256 = v_15253 & v_15255;
assign v_15258 = v_15223 & v_15257;
assign v_15260 = v_12787;
assign v_15262 = v_15259 & v_15261;
assign v_15264 = v_15220 & v_15263;
assign v_15266 = v_12783;
assign v_15268 = v_15265 & v_15267;
assign v_15270 = v_15217 & v_15269;
assign v_15272 = v_12779;
assign v_15274 = v_15271 & v_15273;
assign v_15276 = v_15214 & v_15275;
assign v_15278 = v_12775;
assign v_15280 = v_15277 & v_15279;
assign v_15282 = v_15211 & v_15281;
assign v_15284 = v_12771;
assign v_15286 = v_15283 & v_15285;
assign v_15288 = v_15208 & v_15287;
assign v_15290 = v_12767;
assign v_15292 = v_15289 & v_15291;
assign v_15294 = v_15205 & v_15293;
assign v_15296 = v_12763;
assign v_15298 = v_15295 & v_15297;
assign v_15300 = v_15202 & v_15299;
assign v_15302 = v_12759;
assign v_15304 = v_15301 & v_15303;
assign v_15306 = v_15199 & v_15305;
assign v_15308 = v_12755;
assign v_15310 = v_15307 & v_15309;
assign v_15312 = v_15196 & v_15311;
assign v_15314 = v_2635;
assign v_15316 = v_15313 & v_15315;
assign v_15318 = v_15193 & v_15317;
assign v_15320 = v_2631;
assign v_15322 = v_15319 & v_15321;
assign v_15324 = v_15190 & v_15323;
assign v_15326 = v_2627;
assign v_15328 = v_15325 & v_15327;
assign v_15330 = v_15187 & v_15329;
assign v_15332 = v_2623;
assign v_15334 = v_15331 & v_15333;
assign v_15335 = v_15334;
assign v_15337 = v_12803;
assign v_15338 = v_2688;
assign v_15339 = v_15338;
assign v_15340 = v_15337 & v_15339;
assign v_15341 = v_15340;
assign v_15342 = v_15232 & v_15341;
assign v_15344 = v_15242 & v_15343;
assign v_15345 = v_15231 & v_15341;
assign v_15347 = v_15229 & v_15346;
assign v_15349 = v_15248 & v_15348;
assign v_15350 = v_15228 & v_15346;
assign v_15352 = v_15226 & v_15351;
assign v_15354 = v_15254 & v_15353;
assign v_15355 = v_15225 & v_15351;
assign v_15357 = v_15223 & v_15356;
assign v_15359 = v_15260 & v_15358;
assign v_15360 = v_15222 & v_15356;
assign v_15362 = v_15220 & v_15361;
assign v_15364 = v_15266 & v_15363;
assign v_15365 = v_15219 & v_15361;
assign v_15367 = v_15217 & v_15366;
assign v_15369 = v_15272 & v_15368;
assign v_15370 = v_15216 & v_15366;
assign v_15372 = v_15214 & v_15371;
assign v_15374 = v_15278 & v_15373;
assign v_15375 = v_15213 & v_15371;
assign v_15377 = v_15211 & v_15376;
assign v_15379 = v_15284 & v_15378;
assign v_15380 = v_15210 & v_15376;
assign v_15382 = v_15208 & v_15381;
assign v_15384 = v_15290 & v_15383;
assign v_15385 = v_15207 & v_15381;
assign v_15387 = v_15205 & v_15386;
assign v_15389 = v_15296 & v_15388;
assign v_15390 = v_15204 & v_15386;
assign v_15392 = v_15202 & v_15391;
assign v_15394 = v_15302 & v_15393;
assign v_15395 = v_15201 & v_15391;
assign v_15397 = v_15199 & v_15396;
assign v_15399 = v_15308 & v_15398;
assign v_15400 = v_15198 & v_15396;
assign v_15402 = v_15196 & v_15401;
assign v_15404 = v_15314 & v_15403;
assign v_15405 = v_15195 & v_15401;
assign v_15407 = v_15193 & v_15406;
assign v_15409 = v_15320 & v_15408;
assign v_15410 = v_15192 & v_15406;
assign v_15412 = v_15190 & v_15411;
assign v_15414 = v_15326 & v_15413;
assign v_15415 = v_15189 & v_15411;
assign v_15417 = v_15187 & v_15416;
assign v_15419 = v_15332 & v_15418;
assign v_15420 = v_15186 & v_15416;
assign v_15422 = v_15421;
assign v_15424 = v_15336 & v_15423;
assign v_15425 = v_15424;
assign v_15427 = v_15426;
assign v_15429 = ~v_2883;
assign v_15430 = ~v_12740;
assign v_15431 = v_12740;
assign v_15432 = ~v_2887;
assign v_15433 = ~v_12744;
assign v_15434 = v_12744;
assign v_15435 = ~v_2891;
assign v_15436 = ~v_12748;
assign v_15437 = v_12748;
assign v_15438 = ~v_2895;
assign v_15439 = ~v_12752;
assign v_15440 = v_12752;
assign v_15441 = ~v_12755;
assign v_15442 = ~v_2900;
assign v_15443 = v_2900;
assign v_15444 = ~v_12759;
assign v_15445 = ~v_2904;
assign v_15446 = v_2904;
assign v_15447 = ~v_12763;
assign v_15448 = ~v_2908;
assign v_15449 = v_2908;
assign v_15450 = ~v_12767;
assign v_15451 = ~v_2912;
assign v_15452 = v_2912;
assign v_15453 = ~v_12771;
assign v_15454 = ~v_2916;
assign v_15455 = v_2916;
assign v_15456 = ~v_12775;
assign v_15457 = ~v_2920;
assign v_15458 = v_2920;
assign v_15459 = ~v_12779;
assign v_15460 = ~v_2924;
assign v_15461 = v_2924;
assign v_15462 = ~v_12783;
assign v_15463 = ~v_2928;
assign v_15464 = v_2928;
assign v_15465 = ~v_12787;
assign v_15466 = ~v_2932;
assign v_15467 = v_2932;
assign v_15468 = ~v_12791;
assign v_15469 = ~v_2936;
assign v_15470 = v_2936;
assign v_15471 = ~v_12795;
assign v_15472 = ~v_2940;
assign v_15473 = v_2940;
assign v_15474 = ~v_12799;
assign v_15475 = ~v_2944;
assign v_15476 = v_2944;
assign v_15477 = ~v_12803;
assign v_15478 = ~v_2948;
assign v_15479 = v_15478;
assign v_15481 = v_15480;
assign v_15483 = v_15475 & v_15482;
assign v_15485 = v_12799;
assign v_15487 = v_15484 & v_15486;
assign v_15489 = v_15472 & v_15488;
assign v_15491 = v_12795;
assign v_15493 = v_15490 & v_15492;
assign v_15495 = v_15469 & v_15494;
assign v_15497 = v_12791;
assign v_15499 = v_15496 & v_15498;
assign v_15501 = v_15466 & v_15500;
assign v_15503 = v_12787;
assign v_15505 = v_15502 & v_15504;
assign v_15507 = v_15463 & v_15506;
assign v_15509 = v_12783;
assign v_15511 = v_15508 & v_15510;
assign v_15513 = v_15460 & v_15512;
assign v_15515 = v_12779;
assign v_15517 = v_15514 & v_15516;
assign v_15519 = v_15457 & v_15518;
assign v_15521 = v_12775;
assign v_15523 = v_15520 & v_15522;
assign v_15525 = v_15454 & v_15524;
assign v_15527 = v_12771;
assign v_15529 = v_15526 & v_15528;
assign v_15531 = v_15451 & v_15530;
assign v_15533 = v_12767;
assign v_15535 = v_15532 & v_15534;
assign v_15537 = v_15448 & v_15536;
assign v_15539 = v_12763;
assign v_15541 = v_15538 & v_15540;
assign v_15543 = v_15445 & v_15542;
assign v_15545 = v_12759;
assign v_15547 = v_15544 & v_15546;
assign v_15549 = v_15442 & v_15548;
assign v_15551 = v_12755;
assign v_15553 = v_15550 & v_15552;
assign v_15555 = v_15439 & v_15554;
assign v_15557 = v_2895;
assign v_15559 = v_15556 & v_15558;
assign v_15561 = v_15436 & v_15560;
assign v_15563 = v_2891;
assign v_15565 = v_15562 & v_15564;
assign v_15567 = v_15433 & v_15566;
assign v_15569 = v_2887;
assign v_15571 = v_15568 & v_15570;
assign v_15573 = v_15430 & v_15572;
assign v_15575 = v_2883;
assign v_15577 = v_15574 & v_15576;
assign v_15578 = v_15577;
assign v_15580 = v_12803;
assign v_15581 = v_2948;
assign v_15582 = v_15581;
assign v_15583 = v_15580 & v_15582;
assign v_15584 = v_15583;
assign v_15585 = v_15475 & v_15584;
assign v_15587 = v_15485 & v_15586;
assign v_15588 = v_15474 & v_15584;
assign v_15590 = v_15472 & v_15589;
assign v_15592 = v_15491 & v_15591;
assign v_15593 = v_15471 & v_15589;
assign v_15595 = v_15469 & v_15594;
assign v_15597 = v_15497 & v_15596;
assign v_15598 = v_15468 & v_15594;
assign v_15600 = v_15466 & v_15599;
assign v_15602 = v_15503 & v_15601;
assign v_15603 = v_15465 & v_15599;
assign v_15605 = v_15463 & v_15604;
assign v_15607 = v_15509 & v_15606;
assign v_15608 = v_15462 & v_15604;
assign v_15610 = v_15460 & v_15609;
assign v_15612 = v_15515 & v_15611;
assign v_15613 = v_15459 & v_15609;
assign v_15615 = v_15457 & v_15614;
assign v_15617 = v_15521 & v_15616;
assign v_15618 = v_15456 & v_15614;
assign v_15620 = v_15454 & v_15619;
assign v_15622 = v_15527 & v_15621;
assign v_15623 = v_15453 & v_15619;
assign v_15625 = v_15451 & v_15624;
assign v_15627 = v_15533 & v_15626;
assign v_15628 = v_15450 & v_15624;
assign v_15630 = v_15448 & v_15629;
assign v_15632 = v_15539 & v_15631;
assign v_15633 = v_15447 & v_15629;
assign v_15635 = v_15445 & v_15634;
assign v_15637 = v_15545 & v_15636;
assign v_15638 = v_15444 & v_15634;
assign v_15640 = v_15442 & v_15639;
assign v_15642 = v_15551 & v_15641;
assign v_15643 = v_15441 & v_15639;
assign v_15645 = v_15439 & v_15644;
assign v_15647 = v_15557 & v_15646;
assign v_15648 = v_15438 & v_15644;
assign v_15650 = v_15436 & v_15649;
assign v_15652 = v_15563 & v_15651;
assign v_15653 = v_15435 & v_15649;
assign v_15655 = v_15433 & v_15654;
assign v_15657 = v_15569 & v_15656;
assign v_15658 = v_15432 & v_15654;
assign v_15660 = v_15430 & v_15659;
assign v_15662 = v_15575 & v_15661;
assign v_15663 = v_15429 & v_15659;
assign v_15665 = v_15664;
assign v_15667 = v_15579 & v_15666;
assign v_15668 = v_15667;
assign v_15670 = v_15669;
assign v_15672 = ~v_3143;
assign v_15673 = ~v_12740;
assign v_15674 = v_12740;
assign v_15675 = ~v_3147;
assign v_15676 = ~v_12744;
assign v_15677 = v_12744;
assign v_15678 = ~v_3151;
assign v_15679 = ~v_12748;
assign v_15680 = v_12748;
assign v_15681 = ~v_3155;
assign v_15682 = ~v_12752;
assign v_15683 = v_12752;
assign v_15684 = ~v_12755;
assign v_15685 = ~v_3160;
assign v_15686 = v_3160;
assign v_15687 = ~v_12759;
assign v_15688 = ~v_3164;
assign v_15689 = v_3164;
assign v_15690 = ~v_12763;
assign v_15691 = ~v_3168;
assign v_15692 = v_3168;
assign v_15693 = ~v_12767;
assign v_15694 = ~v_3172;
assign v_15695 = v_3172;
assign v_15696 = ~v_12771;
assign v_15697 = ~v_3176;
assign v_15698 = v_3176;
assign v_15699 = ~v_12775;
assign v_15700 = ~v_3180;
assign v_15701 = v_3180;
assign v_15702 = ~v_12779;
assign v_15703 = ~v_3184;
assign v_15704 = v_3184;
assign v_15705 = ~v_12783;
assign v_15706 = ~v_3188;
assign v_15707 = v_3188;
assign v_15708 = ~v_12787;
assign v_15709 = ~v_3192;
assign v_15710 = v_3192;
assign v_15711 = ~v_12791;
assign v_15712 = ~v_3196;
assign v_15713 = v_3196;
assign v_15714 = ~v_12795;
assign v_15715 = ~v_3200;
assign v_15716 = v_3200;
assign v_15717 = ~v_12799;
assign v_15718 = ~v_3204;
assign v_15719 = v_3204;
assign v_15720 = ~v_12803;
assign v_15721 = ~v_3208;
assign v_15722 = v_15721;
assign v_15724 = v_15723;
assign v_15726 = v_15718 & v_15725;
assign v_15728 = v_12799;
assign v_15730 = v_15727 & v_15729;
assign v_15732 = v_15715 & v_15731;
assign v_15734 = v_12795;
assign v_15736 = v_15733 & v_15735;
assign v_15738 = v_15712 & v_15737;
assign v_15740 = v_12791;
assign v_15742 = v_15739 & v_15741;
assign v_15744 = v_15709 & v_15743;
assign v_15746 = v_12787;
assign v_15748 = v_15745 & v_15747;
assign v_15750 = v_15706 & v_15749;
assign v_15752 = v_12783;
assign v_15754 = v_15751 & v_15753;
assign v_15756 = v_15703 & v_15755;
assign v_15758 = v_12779;
assign v_15760 = v_15757 & v_15759;
assign v_15762 = v_15700 & v_15761;
assign v_15764 = v_12775;
assign v_15766 = v_15763 & v_15765;
assign v_15768 = v_15697 & v_15767;
assign v_15770 = v_12771;
assign v_15772 = v_15769 & v_15771;
assign v_15774 = v_15694 & v_15773;
assign v_15776 = v_12767;
assign v_15778 = v_15775 & v_15777;
assign v_15780 = v_15691 & v_15779;
assign v_15782 = v_12763;
assign v_15784 = v_15781 & v_15783;
assign v_15786 = v_15688 & v_15785;
assign v_15788 = v_12759;
assign v_15790 = v_15787 & v_15789;
assign v_15792 = v_15685 & v_15791;
assign v_15794 = v_12755;
assign v_15796 = v_15793 & v_15795;
assign v_15798 = v_15682 & v_15797;
assign v_15800 = v_3155;
assign v_15802 = v_15799 & v_15801;
assign v_15804 = v_15679 & v_15803;
assign v_15806 = v_3151;
assign v_15808 = v_15805 & v_15807;
assign v_15810 = v_15676 & v_15809;
assign v_15812 = v_3147;
assign v_15814 = v_15811 & v_15813;
assign v_15816 = v_15673 & v_15815;
assign v_15818 = v_3143;
assign v_15820 = v_15817 & v_15819;
assign v_15821 = v_15820;
assign v_15823 = v_12803;
assign v_15824 = v_3208;
assign v_15825 = v_15824;
assign v_15826 = v_15823 & v_15825;
assign v_15827 = v_15826;
assign v_15828 = v_15718 & v_15827;
assign v_15830 = v_15728 & v_15829;
assign v_15831 = v_15717 & v_15827;
assign v_15833 = v_15715 & v_15832;
assign v_15835 = v_15734 & v_15834;
assign v_15836 = v_15714 & v_15832;
assign v_15838 = v_15712 & v_15837;
assign v_15840 = v_15740 & v_15839;
assign v_15841 = v_15711 & v_15837;
assign v_15843 = v_15709 & v_15842;
assign v_15845 = v_15746 & v_15844;
assign v_15846 = v_15708 & v_15842;
assign v_15848 = v_15706 & v_15847;
assign v_15850 = v_15752 & v_15849;
assign v_15851 = v_15705 & v_15847;
assign v_15853 = v_15703 & v_15852;
assign v_15855 = v_15758 & v_15854;
assign v_15856 = v_15702 & v_15852;
assign v_15858 = v_15700 & v_15857;
assign v_15860 = v_15764 & v_15859;
assign v_15861 = v_15699 & v_15857;
assign v_15863 = v_15697 & v_15862;
assign v_15865 = v_15770 & v_15864;
assign v_15866 = v_15696 & v_15862;
assign v_15868 = v_15694 & v_15867;
assign v_15870 = v_15776 & v_15869;
assign v_15871 = v_15693 & v_15867;
assign v_15873 = v_15691 & v_15872;
assign v_15875 = v_15782 & v_15874;
assign v_15876 = v_15690 & v_15872;
assign v_15878 = v_15688 & v_15877;
assign v_15880 = v_15788 & v_15879;
assign v_15881 = v_15687 & v_15877;
assign v_15883 = v_15685 & v_15882;
assign v_15885 = v_15794 & v_15884;
assign v_15886 = v_15684 & v_15882;
assign v_15888 = v_15682 & v_15887;
assign v_15890 = v_15800 & v_15889;
assign v_15891 = v_15681 & v_15887;
assign v_15893 = v_15679 & v_15892;
assign v_15895 = v_15806 & v_15894;
assign v_15896 = v_15678 & v_15892;
assign v_15898 = v_15676 & v_15897;
assign v_15900 = v_15812 & v_15899;
assign v_15901 = v_15675 & v_15897;
assign v_15903 = v_15673 & v_15902;
assign v_15905 = v_15818 & v_15904;
assign v_15906 = v_15672 & v_15902;
assign v_15908 = v_15907;
assign v_15910 = v_15822 & v_15909;
assign v_15911 = v_15910;
assign v_15913 = v_15912;
assign v_15915 = ~v_3403;
assign v_15916 = ~v_12740;
assign v_15917 = v_12740;
assign v_15918 = ~v_3407;
assign v_15919 = ~v_12744;
assign v_15920 = v_12744;
assign v_15921 = ~v_3411;
assign v_15922 = ~v_12748;
assign v_15923 = v_12748;
assign v_15924 = ~v_3415;
assign v_15925 = ~v_12752;
assign v_15926 = v_12752;
assign v_15927 = ~v_12755;
assign v_15928 = ~v_3420;
assign v_15929 = v_3420;
assign v_15930 = ~v_12759;
assign v_15931 = ~v_3424;
assign v_15932 = v_3424;
assign v_15933 = ~v_12763;
assign v_15934 = ~v_3428;
assign v_15935 = v_3428;
assign v_15936 = ~v_12767;
assign v_15937 = ~v_3432;
assign v_15938 = v_3432;
assign v_15939 = ~v_12771;
assign v_15940 = ~v_3436;
assign v_15941 = v_3436;
assign v_15942 = ~v_12775;
assign v_15943 = ~v_3440;
assign v_15944 = v_3440;
assign v_15945 = ~v_12779;
assign v_15946 = ~v_3444;
assign v_15947 = v_3444;
assign v_15948 = ~v_12783;
assign v_15949 = ~v_3448;
assign v_15950 = v_3448;
assign v_15951 = ~v_12787;
assign v_15952 = ~v_3452;
assign v_15953 = v_3452;
assign v_15954 = ~v_12791;
assign v_15955 = ~v_3456;
assign v_15956 = v_3456;
assign v_15957 = ~v_12795;
assign v_15958 = ~v_3460;
assign v_15959 = v_3460;
assign v_15960 = ~v_12799;
assign v_15961 = ~v_3464;
assign v_15962 = v_3464;
assign v_15963 = ~v_12803;
assign v_15964 = ~v_3468;
assign v_15965 = v_15964;
assign v_15967 = v_15966;
assign v_15969 = v_15961 & v_15968;
assign v_15971 = v_12799;
assign v_15973 = v_15970 & v_15972;
assign v_15975 = v_15958 & v_15974;
assign v_15977 = v_12795;
assign v_15979 = v_15976 & v_15978;
assign v_15981 = v_15955 & v_15980;
assign v_15983 = v_12791;
assign v_15985 = v_15982 & v_15984;
assign v_15987 = v_15952 & v_15986;
assign v_15989 = v_12787;
assign v_15991 = v_15988 & v_15990;
assign v_15993 = v_15949 & v_15992;
assign v_15995 = v_12783;
assign v_15997 = v_15994 & v_15996;
assign v_15999 = v_15946 & v_15998;
assign v_16001 = v_12779;
assign v_16003 = v_16000 & v_16002;
assign v_16005 = v_15943 & v_16004;
assign v_16007 = v_12775;
assign v_16009 = v_16006 & v_16008;
assign v_16011 = v_15940 & v_16010;
assign v_16013 = v_12771;
assign v_16015 = v_16012 & v_16014;
assign v_16017 = v_15937 & v_16016;
assign v_16019 = v_12767;
assign v_16021 = v_16018 & v_16020;
assign v_16023 = v_15934 & v_16022;
assign v_16025 = v_12763;
assign v_16027 = v_16024 & v_16026;
assign v_16029 = v_15931 & v_16028;
assign v_16031 = v_12759;
assign v_16033 = v_16030 & v_16032;
assign v_16035 = v_15928 & v_16034;
assign v_16037 = v_12755;
assign v_16039 = v_16036 & v_16038;
assign v_16041 = v_15925 & v_16040;
assign v_16043 = v_3415;
assign v_16045 = v_16042 & v_16044;
assign v_16047 = v_15922 & v_16046;
assign v_16049 = v_3411;
assign v_16051 = v_16048 & v_16050;
assign v_16053 = v_15919 & v_16052;
assign v_16055 = v_3407;
assign v_16057 = v_16054 & v_16056;
assign v_16059 = v_15916 & v_16058;
assign v_16061 = v_3403;
assign v_16063 = v_16060 & v_16062;
assign v_16064 = v_16063;
assign v_16066 = v_12803;
assign v_16067 = v_3468;
assign v_16068 = v_16067;
assign v_16069 = v_16066 & v_16068;
assign v_16070 = v_16069;
assign v_16071 = v_15961 & v_16070;
assign v_16073 = v_15971 & v_16072;
assign v_16074 = v_15960 & v_16070;
assign v_16076 = v_15958 & v_16075;
assign v_16078 = v_15977 & v_16077;
assign v_16079 = v_15957 & v_16075;
assign v_16081 = v_15955 & v_16080;
assign v_16083 = v_15983 & v_16082;
assign v_16084 = v_15954 & v_16080;
assign v_16086 = v_15952 & v_16085;
assign v_16088 = v_15989 & v_16087;
assign v_16089 = v_15951 & v_16085;
assign v_16091 = v_15949 & v_16090;
assign v_16093 = v_15995 & v_16092;
assign v_16094 = v_15948 & v_16090;
assign v_16096 = v_15946 & v_16095;
assign v_16098 = v_16001 & v_16097;
assign v_16099 = v_15945 & v_16095;
assign v_16101 = v_15943 & v_16100;
assign v_16103 = v_16007 & v_16102;
assign v_16104 = v_15942 & v_16100;
assign v_16106 = v_15940 & v_16105;
assign v_16108 = v_16013 & v_16107;
assign v_16109 = v_15939 & v_16105;
assign v_16111 = v_15937 & v_16110;
assign v_16113 = v_16019 & v_16112;
assign v_16114 = v_15936 & v_16110;
assign v_16116 = v_15934 & v_16115;
assign v_16118 = v_16025 & v_16117;
assign v_16119 = v_15933 & v_16115;
assign v_16121 = v_15931 & v_16120;
assign v_16123 = v_16031 & v_16122;
assign v_16124 = v_15930 & v_16120;
assign v_16126 = v_15928 & v_16125;
assign v_16128 = v_16037 & v_16127;
assign v_16129 = v_15927 & v_16125;
assign v_16131 = v_15925 & v_16130;
assign v_16133 = v_16043 & v_16132;
assign v_16134 = v_15924 & v_16130;
assign v_16136 = v_15922 & v_16135;
assign v_16138 = v_16049 & v_16137;
assign v_16139 = v_15921 & v_16135;
assign v_16141 = v_15919 & v_16140;
assign v_16143 = v_16055 & v_16142;
assign v_16144 = v_15918 & v_16140;
assign v_16146 = v_15916 & v_16145;
assign v_16148 = v_16061 & v_16147;
assign v_16149 = v_15915 & v_16145;
assign v_16151 = v_16150;
assign v_16153 = v_16065 & v_16152;
assign v_16154 = v_16153;
assign v_16156 = v_16155;
assign v_16158 = ~v_3663;
assign v_16159 = ~v_12740;
assign v_16160 = v_12740;
assign v_16161 = ~v_3667;
assign v_16162 = ~v_12744;
assign v_16163 = v_12744;
assign v_16164 = ~v_3671;
assign v_16165 = ~v_12748;
assign v_16166 = v_12748;
assign v_16167 = ~v_3675;
assign v_16168 = ~v_12752;
assign v_16169 = v_12752;
assign v_16170 = ~v_12755;
assign v_16171 = ~v_3680;
assign v_16172 = v_3680;
assign v_16173 = ~v_12759;
assign v_16174 = ~v_3684;
assign v_16175 = v_3684;
assign v_16176 = ~v_12763;
assign v_16177 = ~v_3688;
assign v_16178 = v_3688;
assign v_16179 = ~v_12767;
assign v_16180 = ~v_3692;
assign v_16181 = v_3692;
assign v_16182 = ~v_12771;
assign v_16183 = ~v_3696;
assign v_16184 = v_3696;
assign v_16185 = ~v_12775;
assign v_16186 = ~v_3700;
assign v_16187 = v_3700;
assign v_16188 = ~v_12779;
assign v_16189 = ~v_3704;
assign v_16190 = v_3704;
assign v_16191 = ~v_12783;
assign v_16192 = ~v_3708;
assign v_16193 = v_3708;
assign v_16194 = ~v_12787;
assign v_16195 = ~v_3712;
assign v_16196 = v_3712;
assign v_16197 = ~v_12791;
assign v_16198 = ~v_3716;
assign v_16199 = v_3716;
assign v_16200 = ~v_12795;
assign v_16201 = ~v_3720;
assign v_16202 = v_3720;
assign v_16203 = ~v_12799;
assign v_16204 = ~v_3724;
assign v_16205 = v_3724;
assign v_16206 = ~v_12803;
assign v_16207 = ~v_3728;
assign v_16208 = v_16207;
assign v_16210 = v_16209;
assign v_16212 = v_16204 & v_16211;
assign v_16214 = v_12799;
assign v_16216 = v_16213 & v_16215;
assign v_16218 = v_16201 & v_16217;
assign v_16220 = v_12795;
assign v_16222 = v_16219 & v_16221;
assign v_16224 = v_16198 & v_16223;
assign v_16226 = v_12791;
assign v_16228 = v_16225 & v_16227;
assign v_16230 = v_16195 & v_16229;
assign v_16232 = v_12787;
assign v_16234 = v_16231 & v_16233;
assign v_16236 = v_16192 & v_16235;
assign v_16238 = v_12783;
assign v_16240 = v_16237 & v_16239;
assign v_16242 = v_16189 & v_16241;
assign v_16244 = v_12779;
assign v_16246 = v_16243 & v_16245;
assign v_16248 = v_16186 & v_16247;
assign v_16250 = v_12775;
assign v_16252 = v_16249 & v_16251;
assign v_16254 = v_16183 & v_16253;
assign v_16256 = v_12771;
assign v_16258 = v_16255 & v_16257;
assign v_16260 = v_16180 & v_16259;
assign v_16262 = v_12767;
assign v_16264 = v_16261 & v_16263;
assign v_16266 = v_16177 & v_16265;
assign v_16268 = v_12763;
assign v_16270 = v_16267 & v_16269;
assign v_16272 = v_16174 & v_16271;
assign v_16274 = v_12759;
assign v_16276 = v_16273 & v_16275;
assign v_16278 = v_16171 & v_16277;
assign v_16280 = v_12755;
assign v_16282 = v_16279 & v_16281;
assign v_16284 = v_16168 & v_16283;
assign v_16286 = v_3675;
assign v_16288 = v_16285 & v_16287;
assign v_16290 = v_16165 & v_16289;
assign v_16292 = v_3671;
assign v_16294 = v_16291 & v_16293;
assign v_16296 = v_16162 & v_16295;
assign v_16298 = v_3667;
assign v_16300 = v_16297 & v_16299;
assign v_16302 = v_16159 & v_16301;
assign v_16304 = v_3663;
assign v_16306 = v_16303 & v_16305;
assign v_16307 = v_16306;
assign v_16309 = v_12803;
assign v_16310 = v_3728;
assign v_16311 = v_16310;
assign v_16312 = v_16309 & v_16311;
assign v_16313 = v_16312;
assign v_16314 = v_16204 & v_16313;
assign v_16316 = v_16214 & v_16315;
assign v_16317 = v_16203 & v_16313;
assign v_16319 = v_16201 & v_16318;
assign v_16321 = v_16220 & v_16320;
assign v_16322 = v_16200 & v_16318;
assign v_16324 = v_16198 & v_16323;
assign v_16326 = v_16226 & v_16325;
assign v_16327 = v_16197 & v_16323;
assign v_16329 = v_16195 & v_16328;
assign v_16331 = v_16232 & v_16330;
assign v_16332 = v_16194 & v_16328;
assign v_16334 = v_16192 & v_16333;
assign v_16336 = v_16238 & v_16335;
assign v_16337 = v_16191 & v_16333;
assign v_16339 = v_16189 & v_16338;
assign v_16341 = v_16244 & v_16340;
assign v_16342 = v_16188 & v_16338;
assign v_16344 = v_16186 & v_16343;
assign v_16346 = v_16250 & v_16345;
assign v_16347 = v_16185 & v_16343;
assign v_16349 = v_16183 & v_16348;
assign v_16351 = v_16256 & v_16350;
assign v_16352 = v_16182 & v_16348;
assign v_16354 = v_16180 & v_16353;
assign v_16356 = v_16262 & v_16355;
assign v_16357 = v_16179 & v_16353;
assign v_16359 = v_16177 & v_16358;
assign v_16361 = v_16268 & v_16360;
assign v_16362 = v_16176 & v_16358;
assign v_16364 = v_16174 & v_16363;
assign v_16366 = v_16274 & v_16365;
assign v_16367 = v_16173 & v_16363;
assign v_16369 = v_16171 & v_16368;
assign v_16371 = v_16280 & v_16370;
assign v_16372 = v_16170 & v_16368;
assign v_16374 = v_16168 & v_16373;
assign v_16376 = v_16286 & v_16375;
assign v_16377 = v_16167 & v_16373;
assign v_16379 = v_16165 & v_16378;
assign v_16381 = v_16292 & v_16380;
assign v_16382 = v_16164 & v_16378;
assign v_16384 = v_16162 & v_16383;
assign v_16386 = v_16298 & v_16385;
assign v_16387 = v_16161 & v_16383;
assign v_16389 = v_16159 & v_16388;
assign v_16391 = v_16304 & v_16390;
assign v_16392 = v_16158 & v_16388;
assign v_16394 = v_16393;
assign v_16396 = v_16308 & v_16395;
assign v_16397 = v_16396;
assign v_16399 = v_16398;
assign v_16401 = ~v_3923;
assign v_16402 = ~v_12740;
assign v_16403 = v_12740;
assign v_16404 = ~v_3927;
assign v_16405 = ~v_12744;
assign v_16406 = v_12744;
assign v_16407 = ~v_3931;
assign v_16408 = ~v_12748;
assign v_16409 = v_12748;
assign v_16410 = ~v_3935;
assign v_16411 = ~v_12752;
assign v_16412 = v_12752;
assign v_16413 = ~v_12755;
assign v_16414 = ~v_3940;
assign v_16415 = v_3940;
assign v_16416 = ~v_12759;
assign v_16417 = ~v_3944;
assign v_16418 = v_3944;
assign v_16419 = ~v_12763;
assign v_16420 = ~v_3948;
assign v_16421 = v_3948;
assign v_16422 = ~v_12767;
assign v_16423 = ~v_3952;
assign v_16424 = v_3952;
assign v_16425 = ~v_12771;
assign v_16426 = ~v_3956;
assign v_16427 = v_3956;
assign v_16428 = ~v_12775;
assign v_16429 = ~v_3960;
assign v_16430 = v_3960;
assign v_16431 = ~v_12779;
assign v_16432 = ~v_3964;
assign v_16433 = v_3964;
assign v_16434 = ~v_12783;
assign v_16435 = ~v_3968;
assign v_16436 = v_3968;
assign v_16437 = ~v_12787;
assign v_16438 = ~v_3972;
assign v_16439 = v_3972;
assign v_16440 = ~v_12791;
assign v_16441 = ~v_3976;
assign v_16442 = v_3976;
assign v_16443 = ~v_12795;
assign v_16444 = ~v_3980;
assign v_16445 = v_3980;
assign v_16446 = ~v_12799;
assign v_16447 = ~v_3984;
assign v_16448 = v_3984;
assign v_16449 = ~v_12803;
assign v_16450 = ~v_3988;
assign v_16451 = v_16450;
assign v_16453 = v_16452;
assign v_16455 = v_16447 & v_16454;
assign v_16457 = v_12799;
assign v_16459 = v_16456 & v_16458;
assign v_16461 = v_16444 & v_16460;
assign v_16463 = v_12795;
assign v_16465 = v_16462 & v_16464;
assign v_16467 = v_16441 & v_16466;
assign v_16469 = v_12791;
assign v_16471 = v_16468 & v_16470;
assign v_16473 = v_16438 & v_16472;
assign v_16475 = v_12787;
assign v_16477 = v_16474 & v_16476;
assign v_16479 = v_16435 & v_16478;
assign v_16481 = v_12783;
assign v_16483 = v_16480 & v_16482;
assign v_16485 = v_16432 & v_16484;
assign v_16487 = v_12779;
assign v_16489 = v_16486 & v_16488;
assign v_16491 = v_16429 & v_16490;
assign v_16493 = v_12775;
assign v_16495 = v_16492 & v_16494;
assign v_16497 = v_16426 & v_16496;
assign v_16499 = v_12771;
assign v_16501 = v_16498 & v_16500;
assign v_16503 = v_16423 & v_16502;
assign v_16505 = v_12767;
assign v_16507 = v_16504 & v_16506;
assign v_16509 = v_16420 & v_16508;
assign v_16511 = v_12763;
assign v_16513 = v_16510 & v_16512;
assign v_16515 = v_16417 & v_16514;
assign v_16517 = v_12759;
assign v_16519 = v_16516 & v_16518;
assign v_16521 = v_16414 & v_16520;
assign v_16523 = v_12755;
assign v_16525 = v_16522 & v_16524;
assign v_16527 = v_16411 & v_16526;
assign v_16529 = v_3935;
assign v_16531 = v_16528 & v_16530;
assign v_16533 = v_16408 & v_16532;
assign v_16535 = v_3931;
assign v_16537 = v_16534 & v_16536;
assign v_16539 = v_16405 & v_16538;
assign v_16541 = v_3927;
assign v_16543 = v_16540 & v_16542;
assign v_16545 = v_16402 & v_16544;
assign v_16547 = v_3923;
assign v_16549 = v_16546 & v_16548;
assign v_16550 = v_16549;
assign v_16552 = v_12803;
assign v_16553 = v_3988;
assign v_16554 = v_16553;
assign v_16555 = v_16552 & v_16554;
assign v_16556 = v_16555;
assign v_16557 = v_16447 & v_16556;
assign v_16559 = v_16457 & v_16558;
assign v_16560 = v_16446 & v_16556;
assign v_16562 = v_16444 & v_16561;
assign v_16564 = v_16463 & v_16563;
assign v_16565 = v_16443 & v_16561;
assign v_16567 = v_16441 & v_16566;
assign v_16569 = v_16469 & v_16568;
assign v_16570 = v_16440 & v_16566;
assign v_16572 = v_16438 & v_16571;
assign v_16574 = v_16475 & v_16573;
assign v_16575 = v_16437 & v_16571;
assign v_16577 = v_16435 & v_16576;
assign v_16579 = v_16481 & v_16578;
assign v_16580 = v_16434 & v_16576;
assign v_16582 = v_16432 & v_16581;
assign v_16584 = v_16487 & v_16583;
assign v_16585 = v_16431 & v_16581;
assign v_16587 = v_16429 & v_16586;
assign v_16589 = v_16493 & v_16588;
assign v_16590 = v_16428 & v_16586;
assign v_16592 = v_16426 & v_16591;
assign v_16594 = v_16499 & v_16593;
assign v_16595 = v_16425 & v_16591;
assign v_16597 = v_16423 & v_16596;
assign v_16599 = v_16505 & v_16598;
assign v_16600 = v_16422 & v_16596;
assign v_16602 = v_16420 & v_16601;
assign v_16604 = v_16511 & v_16603;
assign v_16605 = v_16419 & v_16601;
assign v_16607 = v_16417 & v_16606;
assign v_16609 = v_16517 & v_16608;
assign v_16610 = v_16416 & v_16606;
assign v_16612 = v_16414 & v_16611;
assign v_16614 = v_16523 & v_16613;
assign v_16615 = v_16413 & v_16611;
assign v_16617 = v_16411 & v_16616;
assign v_16619 = v_16529 & v_16618;
assign v_16620 = v_16410 & v_16616;
assign v_16622 = v_16408 & v_16621;
assign v_16624 = v_16535 & v_16623;
assign v_16625 = v_16407 & v_16621;
assign v_16627 = v_16405 & v_16626;
assign v_16629 = v_16541 & v_16628;
assign v_16630 = v_16404 & v_16626;
assign v_16632 = v_16402 & v_16631;
assign v_16634 = v_16547 & v_16633;
assign v_16635 = v_16401 & v_16631;
assign v_16637 = v_16636;
assign v_16639 = v_16551 & v_16638;
assign v_16640 = v_16639;
assign v_16642 = v_16641;
assign v_16643 = ~v_4182;
assign v_16644 = ~v_12740;
assign v_16645 = v_12740;
assign v_16646 = ~v_4186;
assign v_16647 = ~v_12744;
assign v_16648 = v_12744;
assign v_16649 = ~v_4190;
assign v_16650 = ~v_12748;
assign v_16651 = v_12748;
assign v_16652 = ~v_4194;
assign v_16653 = ~v_12752;
assign v_16654 = v_12752;
assign v_16655 = ~v_12755;
assign v_16656 = ~v_4199;
assign v_16657 = v_4199;
assign v_16658 = ~v_12759;
assign v_16659 = ~v_4203;
assign v_16660 = v_4203;
assign v_16661 = ~v_12763;
assign v_16662 = ~v_4207;
assign v_16663 = v_4207;
assign v_16664 = ~v_12767;
assign v_16665 = ~v_4211;
assign v_16666 = v_4211;
assign v_16667 = ~v_12771;
assign v_16668 = ~v_4215;
assign v_16669 = v_4215;
assign v_16670 = ~v_12775;
assign v_16671 = ~v_4219;
assign v_16672 = v_4219;
assign v_16673 = ~v_12779;
assign v_16674 = ~v_4223;
assign v_16675 = v_4223;
assign v_16676 = ~v_12783;
assign v_16677 = ~v_4227;
assign v_16678 = v_4227;
assign v_16679 = ~v_12787;
assign v_16680 = ~v_4231;
assign v_16681 = v_4231;
assign v_16682 = ~v_12791;
assign v_16683 = ~v_4235;
assign v_16684 = v_4235;
assign v_16685 = ~v_12795;
assign v_16686 = ~v_4239;
assign v_16687 = v_4239;
assign v_16688 = ~v_12799;
assign v_16689 = ~v_4243;
assign v_16690 = v_4243;
assign v_16691 = ~v_12803;
assign v_16692 = ~v_4247;
assign v_16693 = v_16692;
assign v_16695 = v_16694;
assign v_16697 = v_16689 & v_16696;
assign v_16699 = v_12799;
assign v_16701 = v_16698 & v_16700;
assign v_16703 = v_16686 & v_16702;
assign v_16705 = v_12795;
assign v_16707 = v_16704 & v_16706;
assign v_16709 = v_16683 & v_16708;
assign v_16711 = v_12791;
assign v_16713 = v_16710 & v_16712;
assign v_16715 = v_16680 & v_16714;
assign v_16717 = v_12787;
assign v_16719 = v_16716 & v_16718;
assign v_16721 = v_16677 & v_16720;
assign v_16723 = v_12783;
assign v_16725 = v_16722 & v_16724;
assign v_16727 = v_16674 & v_16726;
assign v_16729 = v_12779;
assign v_16731 = v_16728 & v_16730;
assign v_16733 = v_16671 & v_16732;
assign v_16735 = v_12775;
assign v_16737 = v_16734 & v_16736;
assign v_16739 = v_16668 & v_16738;
assign v_16741 = v_12771;
assign v_16743 = v_16740 & v_16742;
assign v_16745 = v_16665 & v_16744;
assign v_16747 = v_12767;
assign v_16749 = v_16746 & v_16748;
assign v_16751 = v_16662 & v_16750;
assign v_16753 = v_12763;
assign v_16755 = v_16752 & v_16754;
assign v_16757 = v_16659 & v_16756;
assign v_16759 = v_12759;
assign v_16761 = v_16758 & v_16760;
assign v_16763 = v_16656 & v_16762;
assign v_16765 = v_12755;
assign v_16767 = v_16764 & v_16766;
assign v_16769 = v_16653 & v_16768;
assign v_16771 = v_4194;
assign v_16773 = v_16770 & v_16772;
assign v_16775 = v_16650 & v_16774;
assign v_16777 = v_4190;
assign v_16779 = v_16776 & v_16778;
assign v_16781 = v_16647 & v_16780;
assign v_16783 = v_4186;
assign v_16785 = v_16782 & v_16784;
assign v_16787 = v_16644 & v_16786;
assign v_16789 = v_4182;
assign v_16791 = v_16788 & v_16790;
assign v_16793 = ~v_16792;
assign v_16795 = v_12803;
assign v_16796 = v_4247;
assign v_16797 = v_16796;
assign v_16798 = v_16795 & v_16797;
assign v_16799 = v_16798;
assign v_16800 = v_16689 & v_16799;
assign v_16802 = v_16699 & v_16801;
assign v_16803 = v_16688 & v_16799;
assign v_16805 = v_16686 & v_16804;
assign v_16807 = v_16705 & v_16806;
assign v_16808 = v_16685 & v_16804;
assign v_16810 = v_16683 & v_16809;
assign v_16812 = v_16711 & v_16811;
assign v_16813 = v_16682 & v_16809;
assign v_16815 = v_16680 & v_16814;
assign v_16817 = v_16717 & v_16816;
assign v_16818 = v_16679 & v_16814;
assign v_16820 = v_16677 & v_16819;
assign v_16822 = v_16723 & v_16821;
assign v_16823 = v_16676 & v_16819;
assign v_16825 = v_16674 & v_16824;
assign v_16827 = v_16729 & v_16826;
assign v_16828 = v_16673 & v_16824;
assign v_16830 = v_16671 & v_16829;
assign v_16832 = v_16735 & v_16831;
assign v_16833 = v_16670 & v_16829;
assign v_16835 = v_16668 & v_16834;
assign v_16837 = v_16741 & v_16836;
assign v_16838 = v_16667 & v_16834;
assign v_16840 = v_16665 & v_16839;
assign v_16842 = v_16747 & v_16841;
assign v_16843 = v_16664 & v_16839;
assign v_16845 = v_16662 & v_16844;
assign v_16847 = v_16753 & v_16846;
assign v_16848 = v_16661 & v_16844;
assign v_16850 = v_16659 & v_16849;
assign v_16852 = v_16759 & v_16851;
assign v_16853 = v_16658 & v_16849;
assign v_16855 = v_16656 & v_16854;
assign v_16857 = v_16765 & v_16856;
assign v_16858 = v_16655 & v_16854;
assign v_16860 = v_16653 & v_16859;
assign v_16862 = v_16771 & v_16861;
assign v_16863 = v_16652 & v_16859;
assign v_16865 = v_16650 & v_16864;
assign v_16867 = v_16777 & v_16866;
assign v_16868 = v_16649 & v_16864;
assign v_16870 = v_16647 & v_16869;
assign v_16872 = v_16783 & v_16871;
assign v_16873 = v_16646 & v_16869;
assign v_16875 = v_16644 & v_16874;
assign v_16877 = v_16789 & v_16876;
assign v_16878 = v_16643 & v_16874;
assign v_16880 = v_16792;
assign v_16882 = v_16794 & v_16881;
assign v_16883 = v_16882;
assign v_16885 = v_16884;
assign v_16887 = ~v_6;
assign v_16889 = ~v_16888;
assign v_16890 = v_16888;
assign v_16891 = ~v_13;
assign v_16893 = ~v_16892;
assign v_16894 = v_16892;
assign v_16895 = ~v_18;
assign v_16897 = ~v_16896;
assign v_16898 = v_16896;
assign v_16899 = ~v_23;
assign v_16901 = ~v_16900;
assign v_16902 = v_16900;
assign v_16904 = ~v_16903;
assign v_16905 = ~v_30;
assign v_16906 = v_30;
assign v_16908 = ~v_16907;
assign v_16909 = ~v_35;
assign v_16910 = v_35;
assign v_16912 = ~v_16911;
assign v_16913 = ~v_40;
assign v_16914 = v_40;
assign v_16916 = ~v_16915;
assign v_16917 = ~v_45;
assign v_16918 = v_45;
assign v_16920 = ~v_16919;
assign v_16921 = ~v_50;
assign v_16922 = v_50;
assign v_16924 = ~v_16923;
assign v_16925 = ~v_55;
assign v_16926 = v_55;
assign v_16928 = ~v_16927;
assign v_16929 = ~v_60;
assign v_16930 = v_60;
assign v_16932 = ~v_16931;
assign v_16933 = ~v_65;
assign v_16934 = v_65;
assign v_16936 = ~v_16935;
assign v_16937 = ~v_70;
assign v_16938 = v_70;
assign v_16940 = ~v_16939;
assign v_16941 = ~v_75;
assign v_16942 = v_75;
assign v_16944 = ~v_16943;
assign v_16945 = ~v_80;
assign v_16946 = v_80;
assign v_16948 = ~v_16947;
assign v_16949 = ~v_85;
assign v_16950 = v_85;
assign v_16952 = ~v_16951;
assign v_16953 = ~v_90;
assign v_16954 = v_16953;
assign v_16956 = v_16955;
assign v_16958 = v_16949 & v_16957;
assign v_16960 = v_16947;
assign v_16962 = v_16959 & v_16961;
assign v_16964 = v_16945 & v_16963;
assign v_16966 = v_16943;
assign v_16968 = v_16965 & v_16967;
assign v_16970 = v_16941 & v_16969;
assign v_16972 = v_16939;
assign v_16974 = v_16971 & v_16973;
assign v_16976 = v_16937 & v_16975;
assign v_16978 = v_16935;
assign v_16980 = v_16977 & v_16979;
assign v_16982 = v_16933 & v_16981;
assign v_16984 = v_16931;
assign v_16986 = v_16983 & v_16985;
assign v_16988 = v_16929 & v_16987;
assign v_16990 = v_16927;
assign v_16992 = v_16989 & v_16991;
assign v_16994 = v_16925 & v_16993;
assign v_16996 = v_16923;
assign v_16998 = v_16995 & v_16997;
assign v_17000 = v_16921 & v_16999;
assign v_17002 = v_16919;
assign v_17004 = v_17001 & v_17003;
assign v_17006 = v_16917 & v_17005;
assign v_17008 = v_16915;
assign v_17010 = v_17007 & v_17009;
assign v_17012 = v_16913 & v_17011;
assign v_17014 = v_16911;
assign v_17016 = v_17013 & v_17015;
assign v_17018 = v_16909 & v_17017;
assign v_17020 = v_16907;
assign v_17022 = v_17019 & v_17021;
assign v_17024 = v_16905 & v_17023;
assign v_17026 = v_16903;
assign v_17028 = v_17025 & v_17027;
assign v_17030 = v_16901 & v_17029;
assign v_17032 = v_23;
assign v_17034 = v_17031 & v_17033;
assign v_17036 = v_16897 & v_17035;
assign v_17038 = v_18;
assign v_17040 = v_17037 & v_17039;
assign v_17042 = v_16893 & v_17041;
assign v_17044 = v_13;
assign v_17046 = v_17043 & v_17045;
assign v_17048 = v_16889 & v_17047;
assign v_17050 = v_6;
assign v_17052 = v_17049 & v_17051;
assign v_17053 = v_17052;
assign v_17055 = v_16951;
assign v_17056 = v_90;
assign v_17057 = v_17056;
assign v_17058 = v_17055 & v_17057;
assign v_17059 = v_17058;
assign v_17060 = v_16949 & v_17059;
assign v_17062 = v_16960 & v_17061;
assign v_17063 = v_16948 & v_17059;
assign v_17065 = v_16945 & v_17064;
assign v_17067 = v_16966 & v_17066;
assign v_17068 = v_16944 & v_17064;
assign v_17070 = v_16941 & v_17069;
assign v_17072 = v_16972 & v_17071;
assign v_17073 = v_16940 & v_17069;
assign v_17075 = v_16937 & v_17074;
assign v_17077 = v_16978 & v_17076;
assign v_17078 = v_16936 & v_17074;
assign v_17080 = v_16933 & v_17079;
assign v_17082 = v_16984 & v_17081;
assign v_17083 = v_16932 & v_17079;
assign v_17085 = v_16929 & v_17084;
assign v_17087 = v_16990 & v_17086;
assign v_17088 = v_16928 & v_17084;
assign v_17090 = v_16925 & v_17089;
assign v_17092 = v_16996 & v_17091;
assign v_17093 = v_16924 & v_17089;
assign v_17095 = v_16921 & v_17094;
assign v_17097 = v_17002 & v_17096;
assign v_17098 = v_16920 & v_17094;
assign v_17100 = v_16917 & v_17099;
assign v_17102 = v_17008 & v_17101;
assign v_17103 = v_16916 & v_17099;
assign v_17105 = v_16913 & v_17104;
assign v_17107 = v_17014 & v_17106;
assign v_17108 = v_16912 & v_17104;
assign v_17110 = v_16909 & v_17109;
assign v_17112 = v_17020 & v_17111;
assign v_17113 = v_16908 & v_17109;
assign v_17115 = v_16905 & v_17114;
assign v_17117 = v_17026 & v_17116;
assign v_17118 = v_16904 & v_17114;
assign v_17120 = v_16901 & v_17119;
assign v_17122 = v_17032 & v_17121;
assign v_17123 = v_16899 & v_17119;
assign v_17125 = v_16897 & v_17124;
assign v_17127 = v_17038 & v_17126;
assign v_17128 = v_16895 & v_17124;
assign v_17130 = v_16893 & v_17129;
assign v_17132 = v_17044 & v_17131;
assign v_17133 = v_16891 & v_17129;
assign v_17135 = v_16889 & v_17134;
assign v_17137 = v_17050 & v_17136;
assign v_17138 = v_16887 & v_17134;
assign v_17140 = v_17139;
assign v_17142 = v_17054 & v_17141;
assign v_17143 = v_17142;
assign v_17145 = v_17144;
assign v_17147 = ~v_283;
assign v_17148 = ~v_16888;
assign v_17149 = v_16888;
assign v_17150 = ~v_287;
assign v_17151 = ~v_16892;
assign v_17152 = v_16892;
assign v_17153 = ~v_291;
assign v_17154 = ~v_16896;
assign v_17155 = v_16896;
assign v_17156 = ~v_295;
assign v_17157 = ~v_16900;
assign v_17158 = v_16900;
assign v_17159 = ~v_16903;
assign v_17160 = ~v_300;
assign v_17161 = v_300;
assign v_17162 = ~v_16907;
assign v_17163 = ~v_304;
assign v_17164 = v_304;
assign v_17165 = ~v_16911;
assign v_17166 = ~v_308;
assign v_17167 = v_308;
assign v_17168 = ~v_16915;
assign v_17169 = ~v_312;
assign v_17170 = v_312;
assign v_17171 = ~v_16919;
assign v_17172 = ~v_316;
assign v_17173 = v_316;
assign v_17174 = ~v_16923;
assign v_17175 = ~v_320;
assign v_17176 = v_320;
assign v_17177 = ~v_16927;
assign v_17178 = ~v_324;
assign v_17179 = v_324;
assign v_17180 = ~v_16931;
assign v_17181 = ~v_328;
assign v_17182 = v_328;
assign v_17183 = ~v_16935;
assign v_17184 = ~v_332;
assign v_17185 = v_332;
assign v_17186 = ~v_16939;
assign v_17187 = ~v_336;
assign v_17188 = v_336;
assign v_17189 = ~v_16943;
assign v_17190 = ~v_340;
assign v_17191 = v_340;
assign v_17192 = ~v_16947;
assign v_17193 = ~v_344;
assign v_17194 = v_344;
assign v_17195 = ~v_16951;
assign v_17196 = ~v_348;
assign v_17197 = v_17196;
assign v_17199 = v_17198;
assign v_17201 = v_17193 & v_17200;
assign v_17203 = v_16947;
assign v_17205 = v_17202 & v_17204;
assign v_17207 = v_17190 & v_17206;
assign v_17209 = v_16943;
assign v_17211 = v_17208 & v_17210;
assign v_17213 = v_17187 & v_17212;
assign v_17215 = v_16939;
assign v_17217 = v_17214 & v_17216;
assign v_17219 = v_17184 & v_17218;
assign v_17221 = v_16935;
assign v_17223 = v_17220 & v_17222;
assign v_17225 = v_17181 & v_17224;
assign v_17227 = v_16931;
assign v_17229 = v_17226 & v_17228;
assign v_17231 = v_17178 & v_17230;
assign v_17233 = v_16927;
assign v_17235 = v_17232 & v_17234;
assign v_17237 = v_17175 & v_17236;
assign v_17239 = v_16923;
assign v_17241 = v_17238 & v_17240;
assign v_17243 = v_17172 & v_17242;
assign v_17245 = v_16919;
assign v_17247 = v_17244 & v_17246;
assign v_17249 = v_17169 & v_17248;
assign v_17251 = v_16915;
assign v_17253 = v_17250 & v_17252;
assign v_17255 = v_17166 & v_17254;
assign v_17257 = v_16911;
assign v_17259 = v_17256 & v_17258;
assign v_17261 = v_17163 & v_17260;
assign v_17263 = v_16907;
assign v_17265 = v_17262 & v_17264;
assign v_17267 = v_17160 & v_17266;
assign v_17269 = v_16903;
assign v_17271 = v_17268 & v_17270;
assign v_17273 = v_17157 & v_17272;
assign v_17275 = v_295;
assign v_17277 = v_17274 & v_17276;
assign v_17279 = v_17154 & v_17278;
assign v_17281 = v_291;
assign v_17283 = v_17280 & v_17282;
assign v_17285 = v_17151 & v_17284;
assign v_17287 = v_287;
assign v_17289 = v_17286 & v_17288;
assign v_17291 = v_17148 & v_17290;
assign v_17293 = v_283;
assign v_17295 = v_17292 & v_17294;
assign v_17296 = v_17295;
assign v_17298 = v_16951;
assign v_17299 = v_348;
assign v_17300 = v_17299;
assign v_17301 = v_17298 & v_17300;
assign v_17302 = v_17301;
assign v_17303 = v_17193 & v_17302;
assign v_17305 = v_17203 & v_17304;
assign v_17306 = v_17192 & v_17302;
assign v_17308 = v_17190 & v_17307;
assign v_17310 = v_17209 & v_17309;
assign v_17311 = v_17189 & v_17307;
assign v_17313 = v_17187 & v_17312;
assign v_17315 = v_17215 & v_17314;
assign v_17316 = v_17186 & v_17312;
assign v_17318 = v_17184 & v_17317;
assign v_17320 = v_17221 & v_17319;
assign v_17321 = v_17183 & v_17317;
assign v_17323 = v_17181 & v_17322;
assign v_17325 = v_17227 & v_17324;
assign v_17326 = v_17180 & v_17322;
assign v_17328 = v_17178 & v_17327;
assign v_17330 = v_17233 & v_17329;
assign v_17331 = v_17177 & v_17327;
assign v_17333 = v_17175 & v_17332;
assign v_17335 = v_17239 & v_17334;
assign v_17336 = v_17174 & v_17332;
assign v_17338 = v_17172 & v_17337;
assign v_17340 = v_17245 & v_17339;
assign v_17341 = v_17171 & v_17337;
assign v_17343 = v_17169 & v_17342;
assign v_17345 = v_17251 & v_17344;
assign v_17346 = v_17168 & v_17342;
assign v_17348 = v_17166 & v_17347;
assign v_17350 = v_17257 & v_17349;
assign v_17351 = v_17165 & v_17347;
assign v_17353 = v_17163 & v_17352;
assign v_17355 = v_17263 & v_17354;
assign v_17356 = v_17162 & v_17352;
assign v_17358 = v_17160 & v_17357;
assign v_17360 = v_17269 & v_17359;
assign v_17361 = v_17159 & v_17357;
assign v_17363 = v_17157 & v_17362;
assign v_17365 = v_17275 & v_17364;
assign v_17366 = v_17156 & v_17362;
assign v_17368 = v_17154 & v_17367;
assign v_17370 = v_17281 & v_17369;
assign v_17371 = v_17153 & v_17367;
assign v_17373 = v_17151 & v_17372;
assign v_17375 = v_17287 & v_17374;
assign v_17376 = v_17150 & v_17372;
assign v_17378 = v_17148 & v_17377;
assign v_17380 = v_17293 & v_17379;
assign v_17381 = v_17147 & v_17377;
assign v_17383 = v_17382;
assign v_17385 = v_17297 & v_17384;
assign v_17386 = v_17385;
assign v_17388 = v_17387;
assign v_17390 = ~v_543;
assign v_17391 = ~v_16888;
assign v_17392 = v_16888;
assign v_17393 = ~v_547;
assign v_17394 = ~v_16892;
assign v_17395 = v_16892;
assign v_17396 = ~v_551;
assign v_17397 = ~v_16896;
assign v_17398 = v_16896;
assign v_17399 = ~v_555;
assign v_17400 = ~v_16900;
assign v_17401 = v_16900;
assign v_17402 = ~v_16903;
assign v_17403 = ~v_560;
assign v_17404 = v_560;
assign v_17405 = ~v_16907;
assign v_17406 = ~v_564;
assign v_17407 = v_564;
assign v_17408 = ~v_16911;
assign v_17409 = ~v_568;
assign v_17410 = v_568;
assign v_17411 = ~v_16915;
assign v_17412 = ~v_572;
assign v_17413 = v_572;
assign v_17414 = ~v_16919;
assign v_17415 = ~v_576;
assign v_17416 = v_576;
assign v_17417 = ~v_16923;
assign v_17418 = ~v_580;
assign v_17419 = v_580;
assign v_17420 = ~v_16927;
assign v_17421 = ~v_584;
assign v_17422 = v_584;
assign v_17423 = ~v_16931;
assign v_17424 = ~v_588;
assign v_17425 = v_588;
assign v_17426 = ~v_16935;
assign v_17427 = ~v_592;
assign v_17428 = v_592;
assign v_17429 = ~v_16939;
assign v_17430 = ~v_596;
assign v_17431 = v_596;
assign v_17432 = ~v_16943;
assign v_17433 = ~v_600;
assign v_17434 = v_600;
assign v_17435 = ~v_16947;
assign v_17436 = ~v_604;
assign v_17437 = v_604;
assign v_17438 = ~v_16951;
assign v_17439 = ~v_608;
assign v_17440 = v_17439;
assign v_17442 = v_17441;
assign v_17444 = v_17436 & v_17443;
assign v_17446 = v_16947;
assign v_17448 = v_17445 & v_17447;
assign v_17450 = v_17433 & v_17449;
assign v_17452 = v_16943;
assign v_17454 = v_17451 & v_17453;
assign v_17456 = v_17430 & v_17455;
assign v_17458 = v_16939;
assign v_17460 = v_17457 & v_17459;
assign v_17462 = v_17427 & v_17461;
assign v_17464 = v_16935;
assign v_17466 = v_17463 & v_17465;
assign v_17468 = v_17424 & v_17467;
assign v_17470 = v_16931;
assign v_17472 = v_17469 & v_17471;
assign v_17474 = v_17421 & v_17473;
assign v_17476 = v_16927;
assign v_17478 = v_17475 & v_17477;
assign v_17480 = v_17418 & v_17479;
assign v_17482 = v_16923;
assign v_17484 = v_17481 & v_17483;
assign v_17486 = v_17415 & v_17485;
assign v_17488 = v_16919;
assign v_17490 = v_17487 & v_17489;
assign v_17492 = v_17412 & v_17491;
assign v_17494 = v_16915;
assign v_17496 = v_17493 & v_17495;
assign v_17498 = v_17409 & v_17497;
assign v_17500 = v_16911;
assign v_17502 = v_17499 & v_17501;
assign v_17504 = v_17406 & v_17503;
assign v_17506 = v_16907;
assign v_17508 = v_17505 & v_17507;
assign v_17510 = v_17403 & v_17509;
assign v_17512 = v_16903;
assign v_17514 = v_17511 & v_17513;
assign v_17516 = v_17400 & v_17515;
assign v_17518 = v_555;
assign v_17520 = v_17517 & v_17519;
assign v_17522 = v_17397 & v_17521;
assign v_17524 = v_551;
assign v_17526 = v_17523 & v_17525;
assign v_17528 = v_17394 & v_17527;
assign v_17530 = v_547;
assign v_17532 = v_17529 & v_17531;
assign v_17534 = v_17391 & v_17533;
assign v_17536 = v_543;
assign v_17538 = v_17535 & v_17537;
assign v_17539 = v_17538;
assign v_17541 = v_16951;
assign v_17542 = v_608;
assign v_17543 = v_17542;
assign v_17544 = v_17541 & v_17543;
assign v_17545 = v_17544;
assign v_17546 = v_17436 & v_17545;
assign v_17548 = v_17446 & v_17547;
assign v_17549 = v_17435 & v_17545;
assign v_17551 = v_17433 & v_17550;
assign v_17553 = v_17452 & v_17552;
assign v_17554 = v_17432 & v_17550;
assign v_17556 = v_17430 & v_17555;
assign v_17558 = v_17458 & v_17557;
assign v_17559 = v_17429 & v_17555;
assign v_17561 = v_17427 & v_17560;
assign v_17563 = v_17464 & v_17562;
assign v_17564 = v_17426 & v_17560;
assign v_17566 = v_17424 & v_17565;
assign v_17568 = v_17470 & v_17567;
assign v_17569 = v_17423 & v_17565;
assign v_17571 = v_17421 & v_17570;
assign v_17573 = v_17476 & v_17572;
assign v_17574 = v_17420 & v_17570;
assign v_17576 = v_17418 & v_17575;
assign v_17578 = v_17482 & v_17577;
assign v_17579 = v_17417 & v_17575;
assign v_17581 = v_17415 & v_17580;
assign v_17583 = v_17488 & v_17582;
assign v_17584 = v_17414 & v_17580;
assign v_17586 = v_17412 & v_17585;
assign v_17588 = v_17494 & v_17587;
assign v_17589 = v_17411 & v_17585;
assign v_17591 = v_17409 & v_17590;
assign v_17593 = v_17500 & v_17592;
assign v_17594 = v_17408 & v_17590;
assign v_17596 = v_17406 & v_17595;
assign v_17598 = v_17506 & v_17597;
assign v_17599 = v_17405 & v_17595;
assign v_17601 = v_17403 & v_17600;
assign v_17603 = v_17512 & v_17602;
assign v_17604 = v_17402 & v_17600;
assign v_17606 = v_17400 & v_17605;
assign v_17608 = v_17518 & v_17607;
assign v_17609 = v_17399 & v_17605;
assign v_17611 = v_17397 & v_17610;
assign v_17613 = v_17524 & v_17612;
assign v_17614 = v_17396 & v_17610;
assign v_17616 = v_17394 & v_17615;
assign v_17618 = v_17530 & v_17617;
assign v_17619 = v_17393 & v_17615;
assign v_17621 = v_17391 & v_17620;
assign v_17623 = v_17536 & v_17622;
assign v_17624 = v_17390 & v_17620;
assign v_17626 = v_17625;
assign v_17628 = v_17540 & v_17627;
assign v_17629 = v_17628;
assign v_17631 = v_17630;
assign v_17633 = ~v_803;
assign v_17634 = ~v_16888;
assign v_17635 = v_16888;
assign v_17636 = ~v_807;
assign v_17637 = ~v_16892;
assign v_17638 = v_16892;
assign v_17639 = ~v_811;
assign v_17640 = ~v_16896;
assign v_17641 = v_16896;
assign v_17642 = ~v_815;
assign v_17643 = ~v_16900;
assign v_17644 = v_16900;
assign v_17645 = ~v_16903;
assign v_17646 = ~v_820;
assign v_17647 = v_820;
assign v_17648 = ~v_16907;
assign v_17649 = ~v_824;
assign v_17650 = v_824;
assign v_17651 = ~v_16911;
assign v_17652 = ~v_828;
assign v_17653 = v_828;
assign v_17654 = ~v_16915;
assign v_17655 = ~v_832;
assign v_17656 = v_832;
assign v_17657 = ~v_16919;
assign v_17658 = ~v_836;
assign v_17659 = v_836;
assign v_17660 = ~v_16923;
assign v_17661 = ~v_840;
assign v_17662 = v_840;
assign v_17663 = ~v_16927;
assign v_17664 = ~v_844;
assign v_17665 = v_844;
assign v_17666 = ~v_16931;
assign v_17667 = ~v_848;
assign v_17668 = v_848;
assign v_17669 = ~v_16935;
assign v_17670 = ~v_852;
assign v_17671 = v_852;
assign v_17672 = ~v_16939;
assign v_17673 = ~v_856;
assign v_17674 = v_856;
assign v_17675 = ~v_16943;
assign v_17676 = ~v_860;
assign v_17677 = v_860;
assign v_17678 = ~v_16947;
assign v_17679 = ~v_864;
assign v_17680 = v_864;
assign v_17681 = ~v_16951;
assign v_17682 = ~v_868;
assign v_17683 = v_17682;
assign v_17685 = v_17684;
assign v_17687 = v_17679 & v_17686;
assign v_17689 = v_16947;
assign v_17691 = v_17688 & v_17690;
assign v_17693 = v_17676 & v_17692;
assign v_17695 = v_16943;
assign v_17697 = v_17694 & v_17696;
assign v_17699 = v_17673 & v_17698;
assign v_17701 = v_16939;
assign v_17703 = v_17700 & v_17702;
assign v_17705 = v_17670 & v_17704;
assign v_17707 = v_16935;
assign v_17709 = v_17706 & v_17708;
assign v_17711 = v_17667 & v_17710;
assign v_17713 = v_16931;
assign v_17715 = v_17712 & v_17714;
assign v_17717 = v_17664 & v_17716;
assign v_17719 = v_16927;
assign v_17721 = v_17718 & v_17720;
assign v_17723 = v_17661 & v_17722;
assign v_17725 = v_16923;
assign v_17727 = v_17724 & v_17726;
assign v_17729 = v_17658 & v_17728;
assign v_17731 = v_16919;
assign v_17733 = v_17730 & v_17732;
assign v_17735 = v_17655 & v_17734;
assign v_17737 = v_16915;
assign v_17739 = v_17736 & v_17738;
assign v_17741 = v_17652 & v_17740;
assign v_17743 = v_16911;
assign v_17745 = v_17742 & v_17744;
assign v_17747 = v_17649 & v_17746;
assign v_17749 = v_16907;
assign v_17751 = v_17748 & v_17750;
assign v_17753 = v_17646 & v_17752;
assign v_17755 = v_16903;
assign v_17757 = v_17754 & v_17756;
assign v_17759 = v_17643 & v_17758;
assign v_17761 = v_815;
assign v_17763 = v_17760 & v_17762;
assign v_17765 = v_17640 & v_17764;
assign v_17767 = v_811;
assign v_17769 = v_17766 & v_17768;
assign v_17771 = v_17637 & v_17770;
assign v_17773 = v_807;
assign v_17775 = v_17772 & v_17774;
assign v_17777 = v_17634 & v_17776;
assign v_17779 = v_803;
assign v_17781 = v_17778 & v_17780;
assign v_17782 = v_17781;
assign v_17784 = v_16951;
assign v_17785 = v_868;
assign v_17786 = v_17785;
assign v_17787 = v_17784 & v_17786;
assign v_17788 = v_17787;
assign v_17789 = v_17679 & v_17788;
assign v_17791 = v_17689 & v_17790;
assign v_17792 = v_17678 & v_17788;
assign v_17794 = v_17676 & v_17793;
assign v_17796 = v_17695 & v_17795;
assign v_17797 = v_17675 & v_17793;
assign v_17799 = v_17673 & v_17798;
assign v_17801 = v_17701 & v_17800;
assign v_17802 = v_17672 & v_17798;
assign v_17804 = v_17670 & v_17803;
assign v_17806 = v_17707 & v_17805;
assign v_17807 = v_17669 & v_17803;
assign v_17809 = v_17667 & v_17808;
assign v_17811 = v_17713 & v_17810;
assign v_17812 = v_17666 & v_17808;
assign v_17814 = v_17664 & v_17813;
assign v_17816 = v_17719 & v_17815;
assign v_17817 = v_17663 & v_17813;
assign v_17819 = v_17661 & v_17818;
assign v_17821 = v_17725 & v_17820;
assign v_17822 = v_17660 & v_17818;
assign v_17824 = v_17658 & v_17823;
assign v_17826 = v_17731 & v_17825;
assign v_17827 = v_17657 & v_17823;
assign v_17829 = v_17655 & v_17828;
assign v_17831 = v_17737 & v_17830;
assign v_17832 = v_17654 & v_17828;
assign v_17834 = v_17652 & v_17833;
assign v_17836 = v_17743 & v_17835;
assign v_17837 = v_17651 & v_17833;
assign v_17839 = v_17649 & v_17838;
assign v_17841 = v_17749 & v_17840;
assign v_17842 = v_17648 & v_17838;
assign v_17844 = v_17646 & v_17843;
assign v_17846 = v_17755 & v_17845;
assign v_17847 = v_17645 & v_17843;
assign v_17849 = v_17643 & v_17848;
assign v_17851 = v_17761 & v_17850;
assign v_17852 = v_17642 & v_17848;
assign v_17854 = v_17640 & v_17853;
assign v_17856 = v_17767 & v_17855;
assign v_17857 = v_17639 & v_17853;
assign v_17859 = v_17637 & v_17858;
assign v_17861 = v_17773 & v_17860;
assign v_17862 = v_17636 & v_17858;
assign v_17864 = v_17634 & v_17863;
assign v_17866 = v_17779 & v_17865;
assign v_17867 = v_17633 & v_17863;
assign v_17869 = v_17868;
assign v_17871 = v_17783 & v_17870;
assign v_17872 = v_17871;
assign v_17874 = v_17873;
assign v_17876 = ~v_1063;
assign v_17877 = ~v_16888;
assign v_17878 = v_16888;
assign v_17879 = ~v_1067;
assign v_17880 = ~v_16892;
assign v_17881 = v_16892;
assign v_17882 = ~v_1071;
assign v_17883 = ~v_16896;
assign v_17884 = v_16896;
assign v_17885 = ~v_1075;
assign v_17886 = ~v_16900;
assign v_17887 = v_16900;
assign v_17888 = ~v_16903;
assign v_17889 = ~v_1080;
assign v_17890 = v_1080;
assign v_17891 = ~v_16907;
assign v_17892 = ~v_1084;
assign v_17893 = v_1084;
assign v_17894 = ~v_16911;
assign v_17895 = ~v_1088;
assign v_17896 = v_1088;
assign v_17897 = ~v_16915;
assign v_17898 = ~v_1092;
assign v_17899 = v_1092;
assign v_17900 = ~v_16919;
assign v_17901 = ~v_1096;
assign v_17902 = v_1096;
assign v_17903 = ~v_16923;
assign v_17904 = ~v_1100;
assign v_17905 = v_1100;
assign v_17906 = ~v_16927;
assign v_17907 = ~v_1104;
assign v_17908 = v_1104;
assign v_17909 = ~v_16931;
assign v_17910 = ~v_1108;
assign v_17911 = v_1108;
assign v_17912 = ~v_16935;
assign v_17913 = ~v_1112;
assign v_17914 = v_1112;
assign v_17915 = ~v_16939;
assign v_17916 = ~v_1116;
assign v_17917 = v_1116;
assign v_17918 = ~v_16943;
assign v_17919 = ~v_1120;
assign v_17920 = v_1120;
assign v_17921 = ~v_16947;
assign v_17922 = ~v_1124;
assign v_17923 = v_1124;
assign v_17924 = ~v_16951;
assign v_17925 = ~v_1128;
assign v_17926 = v_17925;
assign v_17928 = v_17927;
assign v_17930 = v_17922 & v_17929;
assign v_17932 = v_16947;
assign v_17934 = v_17931 & v_17933;
assign v_17936 = v_17919 & v_17935;
assign v_17938 = v_16943;
assign v_17940 = v_17937 & v_17939;
assign v_17942 = v_17916 & v_17941;
assign v_17944 = v_16939;
assign v_17946 = v_17943 & v_17945;
assign v_17948 = v_17913 & v_17947;
assign v_17950 = v_16935;
assign v_17952 = v_17949 & v_17951;
assign v_17954 = v_17910 & v_17953;
assign v_17956 = v_16931;
assign v_17958 = v_17955 & v_17957;
assign v_17960 = v_17907 & v_17959;
assign v_17962 = v_16927;
assign v_17964 = v_17961 & v_17963;
assign v_17966 = v_17904 & v_17965;
assign v_17968 = v_16923;
assign v_17970 = v_17967 & v_17969;
assign v_17972 = v_17901 & v_17971;
assign v_17974 = v_16919;
assign v_17976 = v_17973 & v_17975;
assign v_17978 = v_17898 & v_17977;
assign v_17980 = v_16915;
assign v_17982 = v_17979 & v_17981;
assign v_17984 = v_17895 & v_17983;
assign v_17986 = v_16911;
assign v_17988 = v_17985 & v_17987;
assign v_17990 = v_17892 & v_17989;
assign v_17992 = v_16907;
assign v_17994 = v_17991 & v_17993;
assign v_17996 = v_17889 & v_17995;
assign v_17998 = v_16903;
assign v_18000 = v_17997 & v_17999;
assign v_18002 = v_17886 & v_18001;
assign v_18004 = v_1075;
assign v_18006 = v_18003 & v_18005;
assign v_18008 = v_17883 & v_18007;
assign v_18010 = v_1071;
assign v_18012 = v_18009 & v_18011;
assign v_18014 = v_17880 & v_18013;
assign v_18016 = v_1067;
assign v_18018 = v_18015 & v_18017;
assign v_18020 = v_17877 & v_18019;
assign v_18022 = v_1063;
assign v_18024 = v_18021 & v_18023;
assign v_18025 = v_18024;
assign v_18027 = v_16951;
assign v_18028 = v_1128;
assign v_18029 = v_18028;
assign v_18030 = v_18027 & v_18029;
assign v_18031 = v_18030;
assign v_18032 = v_17922 & v_18031;
assign v_18034 = v_17932 & v_18033;
assign v_18035 = v_17921 & v_18031;
assign v_18037 = v_17919 & v_18036;
assign v_18039 = v_17938 & v_18038;
assign v_18040 = v_17918 & v_18036;
assign v_18042 = v_17916 & v_18041;
assign v_18044 = v_17944 & v_18043;
assign v_18045 = v_17915 & v_18041;
assign v_18047 = v_17913 & v_18046;
assign v_18049 = v_17950 & v_18048;
assign v_18050 = v_17912 & v_18046;
assign v_18052 = v_17910 & v_18051;
assign v_18054 = v_17956 & v_18053;
assign v_18055 = v_17909 & v_18051;
assign v_18057 = v_17907 & v_18056;
assign v_18059 = v_17962 & v_18058;
assign v_18060 = v_17906 & v_18056;
assign v_18062 = v_17904 & v_18061;
assign v_18064 = v_17968 & v_18063;
assign v_18065 = v_17903 & v_18061;
assign v_18067 = v_17901 & v_18066;
assign v_18069 = v_17974 & v_18068;
assign v_18070 = v_17900 & v_18066;
assign v_18072 = v_17898 & v_18071;
assign v_18074 = v_17980 & v_18073;
assign v_18075 = v_17897 & v_18071;
assign v_18077 = v_17895 & v_18076;
assign v_18079 = v_17986 & v_18078;
assign v_18080 = v_17894 & v_18076;
assign v_18082 = v_17892 & v_18081;
assign v_18084 = v_17992 & v_18083;
assign v_18085 = v_17891 & v_18081;
assign v_18087 = v_17889 & v_18086;
assign v_18089 = v_17998 & v_18088;
assign v_18090 = v_17888 & v_18086;
assign v_18092 = v_17886 & v_18091;
assign v_18094 = v_18004 & v_18093;
assign v_18095 = v_17885 & v_18091;
assign v_18097 = v_17883 & v_18096;
assign v_18099 = v_18010 & v_18098;
assign v_18100 = v_17882 & v_18096;
assign v_18102 = v_17880 & v_18101;
assign v_18104 = v_18016 & v_18103;
assign v_18105 = v_17879 & v_18101;
assign v_18107 = v_17877 & v_18106;
assign v_18109 = v_18022 & v_18108;
assign v_18110 = v_17876 & v_18106;
assign v_18112 = v_18111;
assign v_18114 = v_18026 & v_18113;
assign v_18115 = v_18114;
assign v_18117 = v_18116;
assign v_18119 = ~v_1323;
assign v_18120 = ~v_16888;
assign v_18121 = v_16888;
assign v_18122 = ~v_1327;
assign v_18123 = ~v_16892;
assign v_18124 = v_16892;
assign v_18125 = ~v_1331;
assign v_18126 = ~v_16896;
assign v_18127 = v_16896;
assign v_18128 = ~v_1335;
assign v_18129 = ~v_16900;
assign v_18130 = v_16900;
assign v_18131 = ~v_16903;
assign v_18132 = ~v_1340;
assign v_18133 = v_1340;
assign v_18134 = ~v_16907;
assign v_18135 = ~v_1344;
assign v_18136 = v_1344;
assign v_18137 = ~v_16911;
assign v_18138 = ~v_1348;
assign v_18139 = v_1348;
assign v_18140 = ~v_16915;
assign v_18141 = ~v_1352;
assign v_18142 = v_1352;
assign v_18143 = ~v_16919;
assign v_18144 = ~v_1356;
assign v_18145 = v_1356;
assign v_18146 = ~v_16923;
assign v_18147 = ~v_1360;
assign v_18148 = v_1360;
assign v_18149 = ~v_16927;
assign v_18150 = ~v_1364;
assign v_18151 = v_1364;
assign v_18152 = ~v_16931;
assign v_18153 = ~v_1368;
assign v_18154 = v_1368;
assign v_18155 = ~v_16935;
assign v_18156 = ~v_1372;
assign v_18157 = v_1372;
assign v_18158 = ~v_16939;
assign v_18159 = ~v_1376;
assign v_18160 = v_1376;
assign v_18161 = ~v_16943;
assign v_18162 = ~v_1380;
assign v_18163 = v_1380;
assign v_18164 = ~v_16947;
assign v_18165 = ~v_1384;
assign v_18166 = v_1384;
assign v_18167 = ~v_16951;
assign v_18168 = ~v_1388;
assign v_18169 = v_18168;
assign v_18171 = v_18170;
assign v_18173 = v_18165 & v_18172;
assign v_18175 = v_16947;
assign v_18177 = v_18174 & v_18176;
assign v_18179 = v_18162 & v_18178;
assign v_18181 = v_16943;
assign v_18183 = v_18180 & v_18182;
assign v_18185 = v_18159 & v_18184;
assign v_18187 = v_16939;
assign v_18189 = v_18186 & v_18188;
assign v_18191 = v_18156 & v_18190;
assign v_18193 = v_16935;
assign v_18195 = v_18192 & v_18194;
assign v_18197 = v_18153 & v_18196;
assign v_18199 = v_16931;
assign v_18201 = v_18198 & v_18200;
assign v_18203 = v_18150 & v_18202;
assign v_18205 = v_16927;
assign v_18207 = v_18204 & v_18206;
assign v_18209 = v_18147 & v_18208;
assign v_18211 = v_16923;
assign v_18213 = v_18210 & v_18212;
assign v_18215 = v_18144 & v_18214;
assign v_18217 = v_16919;
assign v_18219 = v_18216 & v_18218;
assign v_18221 = v_18141 & v_18220;
assign v_18223 = v_16915;
assign v_18225 = v_18222 & v_18224;
assign v_18227 = v_18138 & v_18226;
assign v_18229 = v_16911;
assign v_18231 = v_18228 & v_18230;
assign v_18233 = v_18135 & v_18232;
assign v_18235 = v_16907;
assign v_18237 = v_18234 & v_18236;
assign v_18239 = v_18132 & v_18238;
assign v_18241 = v_16903;
assign v_18243 = v_18240 & v_18242;
assign v_18245 = v_18129 & v_18244;
assign v_18247 = v_1335;
assign v_18249 = v_18246 & v_18248;
assign v_18251 = v_18126 & v_18250;
assign v_18253 = v_1331;
assign v_18255 = v_18252 & v_18254;
assign v_18257 = v_18123 & v_18256;
assign v_18259 = v_1327;
assign v_18261 = v_18258 & v_18260;
assign v_18263 = v_18120 & v_18262;
assign v_18265 = v_1323;
assign v_18267 = v_18264 & v_18266;
assign v_18268 = v_18267;
assign v_18270 = v_16951;
assign v_18271 = v_1388;
assign v_18272 = v_18271;
assign v_18273 = v_18270 & v_18272;
assign v_18274 = v_18273;
assign v_18275 = v_18165 & v_18274;
assign v_18277 = v_18175 & v_18276;
assign v_18278 = v_18164 & v_18274;
assign v_18280 = v_18162 & v_18279;
assign v_18282 = v_18181 & v_18281;
assign v_18283 = v_18161 & v_18279;
assign v_18285 = v_18159 & v_18284;
assign v_18287 = v_18187 & v_18286;
assign v_18288 = v_18158 & v_18284;
assign v_18290 = v_18156 & v_18289;
assign v_18292 = v_18193 & v_18291;
assign v_18293 = v_18155 & v_18289;
assign v_18295 = v_18153 & v_18294;
assign v_18297 = v_18199 & v_18296;
assign v_18298 = v_18152 & v_18294;
assign v_18300 = v_18150 & v_18299;
assign v_18302 = v_18205 & v_18301;
assign v_18303 = v_18149 & v_18299;
assign v_18305 = v_18147 & v_18304;
assign v_18307 = v_18211 & v_18306;
assign v_18308 = v_18146 & v_18304;
assign v_18310 = v_18144 & v_18309;
assign v_18312 = v_18217 & v_18311;
assign v_18313 = v_18143 & v_18309;
assign v_18315 = v_18141 & v_18314;
assign v_18317 = v_18223 & v_18316;
assign v_18318 = v_18140 & v_18314;
assign v_18320 = v_18138 & v_18319;
assign v_18322 = v_18229 & v_18321;
assign v_18323 = v_18137 & v_18319;
assign v_18325 = v_18135 & v_18324;
assign v_18327 = v_18235 & v_18326;
assign v_18328 = v_18134 & v_18324;
assign v_18330 = v_18132 & v_18329;
assign v_18332 = v_18241 & v_18331;
assign v_18333 = v_18131 & v_18329;
assign v_18335 = v_18129 & v_18334;
assign v_18337 = v_18247 & v_18336;
assign v_18338 = v_18128 & v_18334;
assign v_18340 = v_18126 & v_18339;
assign v_18342 = v_18253 & v_18341;
assign v_18343 = v_18125 & v_18339;
assign v_18345 = v_18123 & v_18344;
assign v_18347 = v_18259 & v_18346;
assign v_18348 = v_18122 & v_18344;
assign v_18350 = v_18120 & v_18349;
assign v_18352 = v_18265 & v_18351;
assign v_18353 = v_18119 & v_18349;
assign v_18355 = v_18354;
assign v_18357 = v_18269 & v_18356;
assign v_18358 = v_18357;
assign v_18360 = v_18359;
assign v_18362 = ~v_1583;
assign v_18363 = ~v_16888;
assign v_18364 = v_16888;
assign v_18365 = ~v_1587;
assign v_18366 = ~v_16892;
assign v_18367 = v_16892;
assign v_18368 = ~v_1591;
assign v_18369 = ~v_16896;
assign v_18370 = v_16896;
assign v_18371 = ~v_1595;
assign v_18372 = ~v_16900;
assign v_18373 = v_16900;
assign v_18374 = ~v_16903;
assign v_18375 = ~v_1600;
assign v_18376 = v_1600;
assign v_18377 = ~v_16907;
assign v_18378 = ~v_1604;
assign v_18379 = v_1604;
assign v_18380 = ~v_16911;
assign v_18381 = ~v_1608;
assign v_18382 = v_1608;
assign v_18383 = ~v_16915;
assign v_18384 = ~v_1612;
assign v_18385 = v_1612;
assign v_18386 = ~v_16919;
assign v_18387 = ~v_1616;
assign v_18388 = v_1616;
assign v_18389 = ~v_16923;
assign v_18390 = ~v_1620;
assign v_18391 = v_1620;
assign v_18392 = ~v_16927;
assign v_18393 = ~v_1624;
assign v_18394 = v_1624;
assign v_18395 = ~v_16931;
assign v_18396 = ~v_1628;
assign v_18397 = v_1628;
assign v_18398 = ~v_16935;
assign v_18399 = ~v_1632;
assign v_18400 = v_1632;
assign v_18401 = ~v_16939;
assign v_18402 = ~v_1636;
assign v_18403 = v_1636;
assign v_18404 = ~v_16943;
assign v_18405 = ~v_1640;
assign v_18406 = v_1640;
assign v_18407 = ~v_16947;
assign v_18408 = ~v_1644;
assign v_18409 = v_1644;
assign v_18410 = ~v_16951;
assign v_18411 = ~v_1648;
assign v_18412 = v_18411;
assign v_18414 = v_18413;
assign v_18416 = v_18408 & v_18415;
assign v_18418 = v_16947;
assign v_18420 = v_18417 & v_18419;
assign v_18422 = v_18405 & v_18421;
assign v_18424 = v_16943;
assign v_18426 = v_18423 & v_18425;
assign v_18428 = v_18402 & v_18427;
assign v_18430 = v_16939;
assign v_18432 = v_18429 & v_18431;
assign v_18434 = v_18399 & v_18433;
assign v_18436 = v_16935;
assign v_18438 = v_18435 & v_18437;
assign v_18440 = v_18396 & v_18439;
assign v_18442 = v_16931;
assign v_18444 = v_18441 & v_18443;
assign v_18446 = v_18393 & v_18445;
assign v_18448 = v_16927;
assign v_18450 = v_18447 & v_18449;
assign v_18452 = v_18390 & v_18451;
assign v_18454 = v_16923;
assign v_18456 = v_18453 & v_18455;
assign v_18458 = v_18387 & v_18457;
assign v_18460 = v_16919;
assign v_18462 = v_18459 & v_18461;
assign v_18464 = v_18384 & v_18463;
assign v_18466 = v_16915;
assign v_18468 = v_18465 & v_18467;
assign v_18470 = v_18381 & v_18469;
assign v_18472 = v_16911;
assign v_18474 = v_18471 & v_18473;
assign v_18476 = v_18378 & v_18475;
assign v_18478 = v_16907;
assign v_18480 = v_18477 & v_18479;
assign v_18482 = v_18375 & v_18481;
assign v_18484 = v_16903;
assign v_18486 = v_18483 & v_18485;
assign v_18488 = v_18372 & v_18487;
assign v_18490 = v_1595;
assign v_18492 = v_18489 & v_18491;
assign v_18494 = v_18369 & v_18493;
assign v_18496 = v_1591;
assign v_18498 = v_18495 & v_18497;
assign v_18500 = v_18366 & v_18499;
assign v_18502 = v_1587;
assign v_18504 = v_18501 & v_18503;
assign v_18506 = v_18363 & v_18505;
assign v_18508 = v_1583;
assign v_18510 = v_18507 & v_18509;
assign v_18511 = v_18510;
assign v_18513 = v_16951;
assign v_18514 = v_1648;
assign v_18515 = v_18514;
assign v_18516 = v_18513 & v_18515;
assign v_18517 = v_18516;
assign v_18518 = v_18408 & v_18517;
assign v_18520 = v_18418 & v_18519;
assign v_18521 = v_18407 & v_18517;
assign v_18523 = v_18405 & v_18522;
assign v_18525 = v_18424 & v_18524;
assign v_18526 = v_18404 & v_18522;
assign v_18528 = v_18402 & v_18527;
assign v_18530 = v_18430 & v_18529;
assign v_18531 = v_18401 & v_18527;
assign v_18533 = v_18399 & v_18532;
assign v_18535 = v_18436 & v_18534;
assign v_18536 = v_18398 & v_18532;
assign v_18538 = v_18396 & v_18537;
assign v_18540 = v_18442 & v_18539;
assign v_18541 = v_18395 & v_18537;
assign v_18543 = v_18393 & v_18542;
assign v_18545 = v_18448 & v_18544;
assign v_18546 = v_18392 & v_18542;
assign v_18548 = v_18390 & v_18547;
assign v_18550 = v_18454 & v_18549;
assign v_18551 = v_18389 & v_18547;
assign v_18553 = v_18387 & v_18552;
assign v_18555 = v_18460 & v_18554;
assign v_18556 = v_18386 & v_18552;
assign v_18558 = v_18384 & v_18557;
assign v_18560 = v_18466 & v_18559;
assign v_18561 = v_18383 & v_18557;
assign v_18563 = v_18381 & v_18562;
assign v_18565 = v_18472 & v_18564;
assign v_18566 = v_18380 & v_18562;
assign v_18568 = v_18378 & v_18567;
assign v_18570 = v_18478 & v_18569;
assign v_18571 = v_18377 & v_18567;
assign v_18573 = v_18375 & v_18572;
assign v_18575 = v_18484 & v_18574;
assign v_18576 = v_18374 & v_18572;
assign v_18578 = v_18372 & v_18577;
assign v_18580 = v_18490 & v_18579;
assign v_18581 = v_18371 & v_18577;
assign v_18583 = v_18369 & v_18582;
assign v_18585 = v_18496 & v_18584;
assign v_18586 = v_18368 & v_18582;
assign v_18588 = v_18366 & v_18587;
assign v_18590 = v_18502 & v_18589;
assign v_18591 = v_18365 & v_18587;
assign v_18593 = v_18363 & v_18592;
assign v_18595 = v_18508 & v_18594;
assign v_18596 = v_18362 & v_18592;
assign v_18598 = v_18597;
assign v_18600 = v_18512 & v_18599;
assign v_18601 = v_18600;
assign v_18603 = v_18602;
assign v_18605 = ~v_1843;
assign v_18606 = ~v_16888;
assign v_18607 = v_16888;
assign v_18608 = ~v_1847;
assign v_18609 = ~v_16892;
assign v_18610 = v_16892;
assign v_18611 = ~v_1851;
assign v_18612 = ~v_16896;
assign v_18613 = v_16896;
assign v_18614 = ~v_1855;
assign v_18615 = ~v_16900;
assign v_18616 = v_16900;
assign v_18617 = ~v_16903;
assign v_18618 = ~v_1860;
assign v_18619 = v_1860;
assign v_18620 = ~v_16907;
assign v_18621 = ~v_1864;
assign v_18622 = v_1864;
assign v_18623 = ~v_16911;
assign v_18624 = ~v_1868;
assign v_18625 = v_1868;
assign v_18626 = ~v_16915;
assign v_18627 = ~v_1872;
assign v_18628 = v_1872;
assign v_18629 = ~v_16919;
assign v_18630 = ~v_1876;
assign v_18631 = v_1876;
assign v_18632 = ~v_16923;
assign v_18633 = ~v_1880;
assign v_18634 = v_1880;
assign v_18635 = ~v_16927;
assign v_18636 = ~v_1884;
assign v_18637 = v_1884;
assign v_18638 = ~v_16931;
assign v_18639 = ~v_1888;
assign v_18640 = v_1888;
assign v_18641 = ~v_16935;
assign v_18642 = ~v_1892;
assign v_18643 = v_1892;
assign v_18644 = ~v_16939;
assign v_18645 = ~v_1896;
assign v_18646 = v_1896;
assign v_18647 = ~v_16943;
assign v_18648 = ~v_1900;
assign v_18649 = v_1900;
assign v_18650 = ~v_16947;
assign v_18651 = ~v_1904;
assign v_18652 = v_1904;
assign v_18653 = ~v_16951;
assign v_18654 = ~v_1908;
assign v_18655 = v_18654;
assign v_18657 = v_18656;
assign v_18659 = v_18651 & v_18658;
assign v_18661 = v_16947;
assign v_18663 = v_18660 & v_18662;
assign v_18665 = v_18648 & v_18664;
assign v_18667 = v_16943;
assign v_18669 = v_18666 & v_18668;
assign v_18671 = v_18645 & v_18670;
assign v_18673 = v_16939;
assign v_18675 = v_18672 & v_18674;
assign v_18677 = v_18642 & v_18676;
assign v_18679 = v_16935;
assign v_18681 = v_18678 & v_18680;
assign v_18683 = v_18639 & v_18682;
assign v_18685 = v_16931;
assign v_18687 = v_18684 & v_18686;
assign v_18689 = v_18636 & v_18688;
assign v_18691 = v_16927;
assign v_18693 = v_18690 & v_18692;
assign v_18695 = v_18633 & v_18694;
assign v_18697 = v_16923;
assign v_18699 = v_18696 & v_18698;
assign v_18701 = v_18630 & v_18700;
assign v_18703 = v_16919;
assign v_18705 = v_18702 & v_18704;
assign v_18707 = v_18627 & v_18706;
assign v_18709 = v_16915;
assign v_18711 = v_18708 & v_18710;
assign v_18713 = v_18624 & v_18712;
assign v_18715 = v_16911;
assign v_18717 = v_18714 & v_18716;
assign v_18719 = v_18621 & v_18718;
assign v_18721 = v_16907;
assign v_18723 = v_18720 & v_18722;
assign v_18725 = v_18618 & v_18724;
assign v_18727 = v_16903;
assign v_18729 = v_18726 & v_18728;
assign v_18731 = v_18615 & v_18730;
assign v_18733 = v_1855;
assign v_18735 = v_18732 & v_18734;
assign v_18737 = v_18612 & v_18736;
assign v_18739 = v_1851;
assign v_18741 = v_18738 & v_18740;
assign v_18743 = v_18609 & v_18742;
assign v_18745 = v_1847;
assign v_18747 = v_18744 & v_18746;
assign v_18749 = v_18606 & v_18748;
assign v_18751 = v_1843;
assign v_18753 = v_18750 & v_18752;
assign v_18754 = v_18753;
assign v_18756 = v_16951;
assign v_18757 = v_1908;
assign v_18758 = v_18757;
assign v_18759 = v_18756 & v_18758;
assign v_18760 = v_18759;
assign v_18761 = v_18651 & v_18760;
assign v_18763 = v_18661 & v_18762;
assign v_18764 = v_18650 & v_18760;
assign v_18766 = v_18648 & v_18765;
assign v_18768 = v_18667 & v_18767;
assign v_18769 = v_18647 & v_18765;
assign v_18771 = v_18645 & v_18770;
assign v_18773 = v_18673 & v_18772;
assign v_18774 = v_18644 & v_18770;
assign v_18776 = v_18642 & v_18775;
assign v_18778 = v_18679 & v_18777;
assign v_18779 = v_18641 & v_18775;
assign v_18781 = v_18639 & v_18780;
assign v_18783 = v_18685 & v_18782;
assign v_18784 = v_18638 & v_18780;
assign v_18786 = v_18636 & v_18785;
assign v_18788 = v_18691 & v_18787;
assign v_18789 = v_18635 & v_18785;
assign v_18791 = v_18633 & v_18790;
assign v_18793 = v_18697 & v_18792;
assign v_18794 = v_18632 & v_18790;
assign v_18796 = v_18630 & v_18795;
assign v_18798 = v_18703 & v_18797;
assign v_18799 = v_18629 & v_18795;
assign v_18801 = v_18627 & v_18800;
assign v_18803 = v_18709 & v_18802;
assign v_18804 = v_18626 & v_18800;
assign v_18806 = v_18624 & v_18805;
assign v_18808 = v_18715 & v_18807;
assign v_18809 = v_18623 & v_18805;
assign v_18811 = v_18621 & v_18810;
assign v_18813 = v_18721 & v_18812;
assign v_18814 = v_18620 & v_18810;
assign v_18816 = v_18618 & v_18815;
assign v_18818 = v_18727 & v_18817;
assign v_18819 = v_18617 & v_18815;
assign v_18821 = v_18615 & v_18820;
assign v_18823 = v_18733 & v_18822;
assign v_18824 = v_18614 & v_18820;
assign v_18826 = v_18612 & v_18825;
assign v_18828 = v_18739 & v_18827;
assign v_18829 = v_18611 & v_18825;
assign v_18831 = v_18609 & v_18830;
assign v_18833 = v_18745 & v_18832;
assign v_18834 = v_18608 & v_18830;
assign v_18836 = v_18606 & v_18835;
assign v_18838 = v_18751 & v_18837;
assign v_18839 = v_18605 & v_18835;
assign v_18841 = v_18840;
assign v_18843 = v_18755 & v_18842;
assign v_18844 = v_18843;
assign v_18846 = v_18845;
assign v_18848 = ~v_2103;
assign v_18849 = ~v_16888;
assign v_18850 = v_16888;
assign v_18851 = ~v_2107;
assign v_18852 = ~v_16892;
assign v_18853 = v_16892;
assign v_18854 = ~v_2111;
assign v_18855 = ~v_16896;
assign v_18856 = v_16896;
assign v_18857 = ~v_2115;
assign v_18858 = ~v_16900;
assign v_18859 = v_16900;
assign v_18860 = ~v_16903;
assign v_18861 = ~v_2120;
assign v_18862 = v_2120;
assign v_18863 = ~v_16907;
assign v_18864 = ~v_2124;
assign v_18865 = v_2124;
assign v_18866 = ~v_16911;
assign v_18867 = ~v_2128;
assign v_18868 = v_2128;
assign v_18869 = ~v_16915;
assign v_18870 = ~v_2132;
assign v_18871 = v_2132;
assign v_18872 = ~v_16919;
assign v_18873 = ~v_2136;
assign v_18874 = v_2136;
assign v_18875 = ~v_16923;
assign v_18876 = ~v_2140;
assign v_18877 = v_2140;
assign v_18878 = ~v_16927;
assign v_18879 = ~v_2144;
assign v_18880 = v_2144;
assign v_18881 = ~v_16931;
assign v_18882 = ~v_2148;
assign v_18883 = v_2148;
assign v_18884 = ~v_16935;
assign v_18885 = ~v_2152;
assign v_18886 = v_2152;
assign v_18887 = ~v_16939;
assign v_18888 = ~v_2156;
assign v_18889 = v_2156;
assign v_18890 = ~v_16943;
assign v_18891 = ~v_2160;
assign v_18892 = v_2160;
assign v_18893 = ~v_16947;
assign v_18894 = ~v_2164;
assign v_18895 = v_2164;
assign v_18896 = ~v_16951;
assign v_18897 = ~v_2168;
assign v_18898 = v_18897;
assign v_18900 = v_18899;
assign v_18902 = v_18894 & v_18901;
assign v_18904 = v_16947;
assign v_18906 = v_18903 & v_18905;
assign v_18908 = v_18891 & v_18907;
assign v_18910 = v_16943;
assign v_18912 = v_18909 & v_18911;
assign v_18914 = v_18888 & v_18913;
assign v_18916 = v_16939;
assign v_18918 = v_18915 & v_18917;
assign v_18920 = v_18885 & v_18919;
assign v_18922 = v_16935;
assign v_18924 = v_18921 & v_18923;
assign v_18926 = v_18882 & v_18925;
assign v_18928 = v_16931;
assign v_18930 = v_18927 & v_18929;
assign v_18932 = v_18879 & v_18931;
assign v_18934 = v_16927;
assign v_18936 = v_18933 & v_18935;
assign v_18938 = v_18876 & v_18937;
assign v_18940 = v_16923;
assign v_18942 = v_18939 & v_18941;
assign v_18944 = v_18873 & v_18943;
assign v_18946 = v_16919;
assign v_18948 = v_18945 & v_18947;
assign v_18950 = v_18870 & v_18949;
assign v_18952 = v_16915;
assign v_18954 = v_18951 & v_18953;
assign v_18956 = v_18867 & v_18955;
assign v_18958 = v_16911;
assign v_18960 = v_18957 & v_18959;
assign v_18962 = v_18864 & v_18961;
assign v_18964 = v_16907;
assign v_18966 = v_18963 & v_18965;
assign v_18968 = v_18861 & v_18967;
assign v_18970 = v_16903;
assign v_18972 = v_18969 & v_18971;
assign v_18974 = v_18858 & v_18973;
assign v_18976 = v_2115;
assign v_18978 = v_18975 & v_18977;
assign v_18980 = v_18855 & v_18979;
assign v_18982 = v_2111;
assign v_18984 = v_18981 & v_18983;
assign v_18986 = v_18852 & v_18985;
assign v_18988 = v_2107;
assign v_18990 = v_18987 & v_18989;
assign v_18992 = v_18849 & v_18991;
assign v_18994 = v_2103;
assign v_18996 = v_18993 & v_18995;
assign v_18997 = v_18996;
assign v_18999 = v_16951;
assign v_19000 = v_2168;
assign v_19001 = v_19000;
assign v_19002 = v_18999 & v_19001;
assign v_19003 = v_19002;
assign v_19004 = v_18894 & v_19003;
assign v_19006 = v_18904 & v_19005;
assign v_19007 = v_18893 & v_19003;
assign v_19009 = v_18891 & v_19008;
assign v_19011 = v_18910 & v_19010;
assign v_19012 = v_18890 & v_19008;
assign v_19014 = v_18888 & v_19013;
assign v_19016 = v_18916 & v_19015;
assign v_19017 = v_18887 & v_19013;
assign v_19019 = v_18885 & v_19018;
assign v_19021 = v_18922 & v_19020;
assign v_19022 = v_18884 & v_19018;
assign v_19024 = v_18882 & v_19023;
assign v_19026 = v_18928 & v_19025;
assign v_19027 = v_18881 & v_19023;
assign v_19029 = v_18879 & v_19028;
assign v_19031 = v_18934 & v_19030;
assign v_19032 = v_18878 & v_19028;
assign v_19034 = v_18876 & v_19033;
assign v_19036 = v_18940 & v_19035;
assign v_19037 = v_18875 & v_19033;
assign v_19039 = v_18873 & v_19038;
assign v_19041 = v_18946 & v_19040;
assign v_19042 = v_18872 & v_19038;
assign v_19044 = v_18870 & v_19043;
assign v_19046 = v_18952 & v_19045;
assign v_19047 = v_18869 & v_19043;
assign v_19049 = v_18867 & v_19048;
assign v_19051 = v_18958 & v_19050;
assign v_19052 = v_18866 & v_19048;
assign v_19054 = v_18864 & v_19053;
assign v_19056 = v_18964 & v_19055;
assign v_19057 = v_18863 & v_19053;
assign v_19059 = v_18861 & v_19058;
assign v_19061 = v_18970 & v_19060;
assign v_19062 = v_18860 & v_19058;
assign v_19064 = v_18858 & v_19063;
assign v_19066 = v_18976 & v_19065;
assign v_19067 = v_18857 & v_19063;
assign v_19069 = v_18855 & v_19068;
assign v_19071 = v_18982 & v_19070;
assign v_19072 = v_18854 & v_19068;
assign v_19074 = v_18852 & v_19073;
assign v_19076 = v_18988 & v_19075;
assign v_19077 = v_18851 & v_19073;
assign v_19079 = v_18849 & v_19078;
assign v_19081 = v_18994 & v_19080;
assign v_19082 = v_18848 & v_19078;
assign v_19084 = v_19083;
assign v_19086 = v_18998 & v_19085;
assign v_19087 = v_19086;
assign v_19089 = v_19088;
assign v_19091 = ~v_2363;
assign v_19092 = ~v_16888;
assign v_19093 = v_16888;
assign v_19094 = ~v_2367;
assign v_19095 = ~v_16892;
assign v_19096 = v_16892;
assign v_19097 = ~v_2371;
assign v_19098 = ~v_16896;
assign v_19099 = v_16896;
assign v_19100 = ~v_2375;
assign v_19101 = ~v_16900;
assign v_19102 = v_16900;
assign v_19103 = ~v_16903;
assign v_19104 = ~v_2380;
assign v_19105 = v_2380;
assign v_19106 = ~v_16907;
assign v_19107 = ~v_2384;
assign v_19108 = v_2384;
assign v_19109 = ~v_16911;
assign v_19110 = ~v_2388;
assign v_19111 = v_2388;
assign v_19112 = ~v_16915;
assign v_19113 = ~v_2392;
assign v_19114 = v_2392;
assign v_19115 = ~v_16919;
assign v_19116 = ~v_2396;
assign v_19117 = v_2396;
assign v_19118 = ~v_16923;
assign v_19119 = ~v_2400;
assign v_19120 = v_2400;
assign v_19121 = ~v_16927;
assign v_19122 = ~v_2404;
assign v_19123 = v_2404;
assign v_19124 = ~v_16931;
assign v_19125 = ~v_2408;
assign v_19126 = v_2408;
assign v_19127 = ~v_16935;
assign v_19128 = ~v_2412;
assign v_19129 = v_2412;
assign v_19130 = ~v_16939;
assign v_19131 = ~v_2416;
assign v_19132 = v_2416;
assign v_19133 = ~v_16943;
assign v_19134 = ~v_2420;
assign v_19135 = v_2420;
assign v_19136 = ~v_16947;
assign v_19137 = ~v_2424;
assign v_19138 = v_2424;
assign v_19139 = ~v_16951;
assign v_19140 = ~v_2428;
assign v_19141 = v_19140;
assign v_19143 = v_19142;
assign v_19145 = v_19137 & v_19144;
assign v_19147 = v_16947;
assign v_19149 = v_19146 & v_19148;
assign v_19151 = v_19134 & v_19150;
assign v_19153 = v_16943;
assign v_19155 = v_19152 & v_19154;
assign v_19157 = v_19131 & v_19156;
assign v_19159 = v_16939;
assign v_19161 = v_19158 & v_19160;
assign v_19163 = v_19128 & v_19162;
assign v_19165 = v_16935;
assign v_19167 = v_19164 & v_19166;
assign v_19169 = v_19125 & v_19168;
assign v_19171 = v_16931;
assign v_19173 = v_19170 & v_19172;
assign v_19175 = v_19122 & v_19174;
assign v_19177 = v_16927;
assign v_19179 = v_19176 & v_19178;
assign v_19181 = v_19119 & v_19180;
assign v_19183 = v_16923;
assign v_19185 = v_19182 & v_19184;
assign v_19187 = v_19116 & v_19186;
assign v_19189 = v_16919;
assign v_19191 = v_19188 & v_19190;
assign v_19193 = v_19113 & v_19192;
assign v_19195 = v_16915;
assign v_19197 = v_19194 & v_19196;
assign v_19199 = v_19110 & v_19198;
assign v_19201 = v_16911;
assign v_19203 = v_19200 & v_19202;
assign v_19205 = v_19107 & v_19204;
assign v_19207 = v_16907;
assign v_19209 = v_19206 & v_19208;
assign v_19211 = v_19104 & v_19210;
assign v_19213 = v_16903;
assign v_19215 = v_19212 & v_19214;
assign v_19217 = v_19101 & v_19216;
assign v_19219 = v_2375;
assign v_19221 = v_19218 & v_19220;
assign v_19223 = v_19098 & v_19222;
assign v_19225 = v_2371;
assign v_19227 = v_19224 & v_19226;
assign v_19229 = v_19095 & v_19228;
assign v_19231 = v_2367;
assign v_19233 = v_19230 & v_19232;
assign v_19235 = v_19092 & v_19234;
assign v_19237 = v_2363;
assign v_19239 = v_19236 & v_19238;
assign v_19240 = v_19239;
assign v_19242 = v_16951;
assign v_19243 = v_2428;
assign v_19244 = v_19243;
assign v_19245 = v_19242 & v_19244;
assign v_19246 = v_19245;
assign v_19247 = v_19137 & v_19246;
assign v_19249 = v_19147 & v_19248;
assign v_19250 = v_19136 & v_19246;
assign v_19252 = v_19134 & v_19251;
assign v_19254 = v_19153 & v_19253;
assign v_19255 = v_19133 & v_19251;
assign v_19257 = v_19131 & v_19256;
assign v_19259 = v_19159 & v_19258;
assign v_19260 = v_19130 & v_19256;
assign v_19262 = v_19128 & v_19261;
assign v_19264 = v_19165 & v_19263;
assign v_19265 = v_19127 & v_19261;
assign v_19267 = v_19125 & v_19266;
assign v_19269 = v_19171 & v_19268;
assign v_19270 = v_19124 & v_19266;
assign v_19272 = v_19122 & v_19271;
assign v_19274 = v_19177 & v_19273;
assign v_19275 = v_19121 & v_19271;
assign v_19277 = v_19119 & v_19276;
assign v_19279 = v_19183 & v_19278;
assign v_19280 = v_19118 & v_19276;
assign v_19282 = v_19116 & v_19281;
assign v_19284 = v_19189 & v_19283;
assign v_19285 = v_19115 & v_19281;
assign v_19287 = v_19113 & v_19286;
assign v_19289 = v_19195 & v_19288;
assign v_19290 = v_19112 & v_19286;
assign v_19292 = v_19110 & v_19291;
assign v_19294 = v_19201 & v_19293;
assign v_19295 = v_19109 & v_19291;
assign v_19297 = v_19107 & v_19296;
assign v_19299 = v_19207 & v_19298;
assign v_19300 = v_19106 & v_19296;
assign v_19302 = v_19104 & v_19301;
assign v_19304 = v_19213 & v_19303;
assign v_19305 = v_19103 & v_19301;
assign v_19307 = v_19101 & v_19306;
assign v_19309 = v_19219 & v_19308;
assign v_19310 = v_19100 & v_19306;
assign v_19312 = v_19098 & v_19311;
assign v_19314 = v_19225 & v_19313;
assign v_19315 = v_19097 & v_19311;
assign v_19317 = v_19095 & v_19316;
assign v_19319 = v_19231 & v_19318;
assign v_19320 = v_19094 & v_19316;
assign v_19322 = v_19092 & v_19321;
assign v_19324 = v_19237 & v_19323;
assign v_19325 = v_19091 & v_19321;
assign v_19327 = v_19326;
assign v_19329 = v_19241 & v_19328;
assign v_19330 = v_19329;
assign v_19332 = v_19331;
assign v_19334 = ~v_2623;
assign v_19335 = ~v_16888;
assign v_19336 = v_16888;
assign v_19337 = ~v_2627;
assign v_19338 = ~v_16892;
assign v_19339 = v_16892;
assign v_19340 = ~v_2631;
assign v_19341 = ~v_16896;
assign v_19342 = v_16896;
assign v_19343 = ~v_2635;
assign v_19344 = ~v_16900;
assign v_19345 = v_16900;
assign v_19346 = ~v_16903;
assign v_19347 = ~v_2640;
assign v_19348 = v_2640;
assign v_19349 = ~v_16907;
assign v_19350 = ~v_2644;
assign v_19351 = v_2644;
assign v_19352 = ~v_16911;
assign v_19353 = ~v_2648;
assign v_19354 = v_2648;
assign v_19355 = ~v_16915;
assign v_19356 = ~v_2652;
assign v_19357 = v_2652;
assign v_19358 = ~v_16919;
assign v_19359 = ~v_2656;
assign v_19360 = v_2656;
assign v_19361 = ~v_16923;
assign v_19362 = ~v_2660;
assign v_19363 = v_2660;
assign v_19364 = ~v_16927;
assign v_19365 = ~v_2664;
assign v_19366 = v_2664;
assign v_19367 = ~v_16931;
assign v_19368 = ~v_2668;
assign v_19369 = v_2668;
assign v_19370 = ~v_16935;
assign v_19371 = ~v_2672;
assign v_19372 = v_2672;
assign v_19373 = ~v_16939;
assign v_19374 = ~v_2676;
assign v_19375 = v_2676;
assign v_19376 = ~v_16943;
assign v_19377 = ~v_2680;
assign v_19378 = v_2680;
assign v_19379 = ~v_16947;
assign v_19380 = ~v_2684;
assign v_19381 = v_2684;
assign v_19382 = ~v_16951;
assign v_19383 = ~v_2688;
assign v_19384 = v_19383;
assign v_19386 = v_19385;
assign v_19388 = v_19380 & v_19387;
assign v_19390 = v_16947;
assign v_19392 = v_19389 & v_19391;
assign v_19394 = v_19377 & v_19393;
assign v_19396 = v_16943;
assign v_19398 = v_19395 & v_19397;
assign v_19400 = v_19374 & v_19399;
assign v_19402 = v_16939;
assign v_19404 = v_19401 & v_19403;
assign v_19406 = v_19371 & v_19405;
assign v_19408 = v_16935;
assign v_19410 = v_19407 & v_19409;
assign v_19412 = v_19368 & v_19411;
assign v_19414 = v_16931;
assign v_19416 = v_19413 & v_19415;
assign v_19418 = v_19365 & v_19417;
assign v_19420 = v_16927;
assign v_19422 = v_19419 & v_19421;
assign v_19424 = v_19362 & v_19423;
assign v_19426 = v_16923;
assign v_19428 = v_19425 & v_19427;
assign v_19430 = v_19359 & v_19429;
assign v_19432 = v_16919;
assign v_19434 = v_19431 & v_19433;
assign v_19436 = v_19356 & v_19435;
assign v_19438 = v_16915;
assign v_19440 = v_19437 & v_19439;
assign v_19442 = v_19353 & v_19441;
assign v_19444 = v_16911;
assign v_19446 = v_19443 & v_19445;
assign v_19448 = v_19350 & v_19447;
assign v_19450 = v_16907;
assign v_19452 = v_19449 & v_19451;
assign v_19454 = v_19347 & v_19453;
assign v_19456 = v_16903;
assign v_19458 = v_19455 & v_19457;
assign v_19460 = v_19344 & v_19459;
assign v_19462 = v_2635;
assign v_19464 = v_19461 & v_19463;
assign v_19466 = v_19341 & v_19465;
assign v_19468 = v_2631;
assign v_19470 = v_19467 & v_19469;
assign v_19472 = v_19338 & v_19471;
assign v_19474 = v_2627;
assign v_19476 = v_19473 & v_19475;
assign v_19478 = v_19335 & v_19477;
assign v_19480 = v_2623;
assign v_19482 = v_19479 & v_19481;
assign v_19483 = v_19482;
assign v_19485 = v_16951;
assign v_19486 = v_2688;
assign v_19487 = v_19486;
assign v_19488 = v_19485 & v_19487;
assign v_19489 = v_19488;
assign v_19490 = v_19380 & v_19489;
assign v_19492 = v_19390 & v_19491;
assign v_19493 = v_19379 & v_19489;
assign v_19495 = v_19377 & v_19494;
assign v_19497 = v_19396 & v_19496;
assign v_19498 = v_19376 & v_19494;
assign v_19500 = v_19374 & v_19499;
assign v_19502 = v_19402 & v_19501;
assign v_19503 = v_19373 & v_19499;
assign v_19505 = v_19371 & v_19504;
assign v_19507 = v_19408 & v_19506;
assign v_19508 = v_19370 & v_19504;
assign v_19510 = v_19368 & v_19509;
assign v_19512 = v_19414 & v_19511;
assign v_19513 = v_19367 & v_19509;
assign v_19515 = v_19365 & v_19514;
assign v_19517 = v_19420 & v_19516;
assign v_19518 = v_19364 & v_19514;
assign v_19520 = v_19362 & v_19519;
assign v_19522 = v_19426 & v_19521;
assign v_19523 = v_19361 & v_19519;
assign v_19525 = v_19359 & v_19524;
assign v_19527 = v_19432 & v_19526;
assign v_19528 = v_19358 & v_19524;
assign v_19530 = v_19356 & v_19529;
assign v_19532 = v_19438 & v_19531;
assign v_19533 = v_19355 & v_19529;
assign v_19535 = v_19353 & v_19534;
assign v_19537 = v_19444 & v_19536;
assign v_19538 = v_19352 & v_19534;
assign v_19540 = v_19350 & v_19539;
assign v_19542 = v_19450 & v_19541;
assign v_19543 = v_19349 & v_19539;
assign v_19545 = v_19347 & v_19544;
assign v_19547 = v_19456 & v_19546;
assign v_19548 = v_19346 & v_19544;
assign v_19550 = v_19344 & v_19549;
assign v_19552 = v_19462 & v_19551;
assign v_19553 = v_19343 & v_19549;
assign v_19555 = v_19341 & v_19554;
assign v_19557 = v_19468 & v_19556;
assign v_19558 = v_19340 & v_19554;
assign v_19560 = v_19338 & v_19559;
assign v_19562 = v_19474 & v_19561;
assign v_19563 = v_19337 & v_19559;
assign v_19565 = v_19335 & v_19564;
assign v_19567 = v_19480 & v_19566;
assign v_19568 = v_19334 & v_19564;
assign v_19570 = v_19569;
assign v_19572 = v_19484 & v_19571;
assign v_19573 = v_19572;
assign v_19575 = v_19574;
assign v_19577 = ~v_2883;
assign v_19578 = ~v_16888;
assign v_19579 = v_16888;
assign v_19580 = ~v_2887;
assign v_19581 = ~v_16892;
assign v_19582 = v_16892;
assign v_19583 = ~v_2891;
assign v_19584 = ~v_16896;
assign v_19585 = v_16896;
assign v_19586 = ~v_2895;
assign v_19587 = ~v_16900;
assign v_19588 = v_16900;
assign v_19589 = ~v_16903;
assign v_19590 = ~v_2900;
assign v_19591 = v_2900;
assign v_19592 = ~v_16907;
assign v_19593 = ~v_2904;
assign v_19594 = v_2904;
assign v_19595 = ~v_16911;
assign v_19596 = ~v_2908;
assign v_19597 = v_2908;
assign v_19598 = ~v_16915;
assign v_19599 = ~v_2912;
assign v_19600 = v_2912;
assign v_19601 = ~v_16919;
assign v_19602 = ~v_2916;
assign v_19603 = v_2916;
assign v_19604 = ~v_16923;
assign v_19605 = ~v_2920;
assign v_19606 = v_2920;
assign v_19607 = ~v_16927;
assign v_19608 = ~v_2924;
assign v_19609 = v_2924;
assign v_19610 = ~v_16931;
assign v_19611 = ~v_2928;
assign v_19612 = v_2928;
assign v_19613 = ~v_16935;
assign v_19614 = ~v_2932;
assign v_19615 = v_2932;
assign v_19616 = ~v_16939;
assign v_19617 = ~v_2936;
assign v_19618 = v_2936;
assign v_19619 = ~v_16943;
assign v_19620 = ~v_2940;
assign v_19621 = v_2940;
assign v_19622 = ~v_16947;
assign v_19623 = ~v_2944;
assign v_19624 = v_2944;
assign v_19625 = ~v_16951;
assign v_19626 = ~v_2948;
assign v_19627 = v_19626;
assign v_19629 = v_19628;
assign v_19631 = v_19623 & v_19630;
assign v_19633 = v_16947;
assign v_19635 = v_19632 & v_19634;
assign v_19637 = v_19620 & v_19636;
assign v_19639 = v_16943;
assign v_19641 = v_19638 & v_19640;
assign v_19643 = v_19617 & v_19642;
assign v_19645 = v_16939;
assign v_19647 = v_19644 & v_19646;
assign v_19649 = v_19614 & v_19648;
assign v_19651 = v_16935;
assign v_19653 = v_19650 & v_19652;
assign v_19655 = v_19611 & v_19654;
assign v_19657 = v_16931;
assign v_19659 = v_19656 & v_19658;
assign v_19661 = v_19608 & v_19660;
assign v_19663 = v_16927;
assign v_19665 = v_19662 & v_19664;
assign v_19667 = v_19605 & v_19666;
assign v_19669 = v_16923;
assign v_19671 = v_19668 & v_19670;
assign v_19673 = v_19602 & v_19672;
assign v_19675 = v_16919;
assign v_19677 = v_19674 & v_19676;
assign v_19679 = v_19599 & v_19678;
assign v_19681 = v_16915;
assign v_19683 = v_19680 & v_19682;
assign v_19685 = v_19596 & v_19684;
assign v_19687 = v_16911;
assign v_19689 = v_19686 & v_19688;
assign v_19691 = v_19593 & v_19690;
assign v_19693 = v_16907;
assign v_19695 = v_19692 & v_19694;
assign v_19697 = v_19590 & v_19696;
assign v_19699 = v_16903;
assign v_19701 = v_19698 & v_19700;
assign v_19703 = v_19587 & v_19702;
assign v_19705 = v_2895;
assign v_19707 = v_19704 & v_19706;
assign v_19709 = v_19584 & v_19708;
assign v_19711 = v_2891;
assign v_19713 = v_19710 & v_19712;
assign v_19715 = v_19581 & v_19714;
assign v_19717 = v_2887;
assign v_19719 = v_19716 & v_19718;
assign v_19721 = v_19578 & v_19720;
assign v_19723 = v_2883;
assign v_19725 = v_19722 & v_19724;
assign v_19726 = v_19725;
assign v_19728 = v_16951;
assign v_19729 = v_2948;
assign v_19730 = v_19729;
assign v_19731 = v_19728 & v_19730;
assign v_19732 = v_19731;
assign v_19733 = v_19623 & v_19732;
assign v_19735 = v_19633 & v_19734;
assign v_19736 = v_19622 & v_19732;
assign v_19738 = v_19620 & v_19737;
assign v_19740 = v_19639 & v_19739;
assign v_19741 = v_19619 & v_19737;
assign v_19743 = v_19617 & v_19742;
assign v_19745 = v_19645 & v_19744;
assign v_19746 = v_19616 & v_19742;
assign v_19748 = v_19614 & v_19747;
assign v_19750 = v_19651 & v_19749;
assign v_19751 = v_19613 & v_19747;
assign v_19753 = v_19611 & v_19752;
assign v_19755 = v_19657 & v_19754;
assign v_19756 = v_19610 & v_19752;
assign v_19758 = v_19608 & v_19757;
assign v_19760 = v_19663 & v_19759;
assign v_19761 = v_19607 & v_19757;
assign v_19763 = v_19605 & v_19762;
assign v_19765 = v_19669 & v_19764;
assign v_19766 = v_19604 & v_19762;
assign v_19768 = v_19602 & v_19767;
assign v_19770 = v_19675 & v_19769;
assign v_19771 = v_19601 & v_19767;
assign v_19773 = v_19599 & v_19772;
assign v_19775 = v_19681 & v_19774;
assign v_19776 = v_19598 & v_19772;
assign v_19778 = v_19596 & v_19777;
assign v_19780 = v_19687 & v_19779;
assign v_19781 = v_19595 & v_19777;
assign v_19783 = v_19593 & v_19782;
assign v_19785 = v_19693 & v_19784;
assign v_19786 = v_19592 & v_19782;
assign v_19788 = v_19590 & v_19787;
assign v_19790 = v_19699 & v_19789;
assign v_19791 = v_19589 & v_19787;
assign v_19793 = v_19587 & v_19792;
assign v_19795 = v_19705 & v_19794;
assign v_19796 = v_19586 & v_19792;
assign v_19798 = v_19584 & v_19797;
assign v_19800 = v_19711 & v_19799;
assign v_19801 = v_19583 & v_19797;
assign v_19803 = v_19581 & v_19802;
assign v_19805 = v_19717 & v_19804;
assign v_19806 = v_19580 & v_19802;
assign v_19808 = v_19578 & v_19807;
assign v_19810 = v_19723 & v_19809;
assign v_19811 = v_19577 & v_19807;
assign v_19813 = v_19812;
assign v_19815 = v_19727 & v_19814;
assign v_19816 = v_19815;
assign v_19818 = v_19817;
assign v_19820 = ~v_3143;
assign v_19821 = ~v_16888;
assign v_19822 = v_16888;
assign v_19823 = ~v_3147;
assign v_19824 = ~v_16892;
assign v_19825 = v_16892;
assign v_19826 = ~v_3151;
assign v_19827 = ~v_16896;
assign v_19828 = v_16896;
assign v_19829 = ~v_3155;
assign v_19830 = ~v_16900;
assign v_19831 = v_16900;
assign v_19832 = ~v_16903;
assign v_19833 = ~v_3160;
assign v_19834 = v_3160;
assign v_19835 = ~v_16907;
assign v_19836 = ~v_3164;
assign v_19837 = v_3164;
assign v_19838 = ~v_16911;
assign v_19839 = ~v_3168;
assign v_19840 = v_3168;
assign v_19841 = ~v_16915;
assign v_19842 = ~v_3172;
assign v_19843 = v_3172;
assign v_19844 = ~v_16919;
assign v_19845 = ~v_3176;
assign v_19846 = v_3176;
assign v_19847 = ~v_16923;
assign v_19848 = ~v_3180;
assign v_19849 = v_3180;
assign v_19850 = ~v_16927;
assign v_19851 = ~v_3184;
assign v_19852 = v_3184;
assign v_19853 = ~v_16931;
assign v_19854 = ~v_3188;
assign v_19855 = v_3188;
assign v_19856 = ~v_16935;
assign v_19857 = ~v_3192;
assign v_19858 = v_3192;
assign v_19859 = ~v_16939;
assign v_19860 = ~v_3196;
assign v_19861 = v_3196;
assign v_19862 = ~v_16943;
assign v_19863 = ~v_3200;
assign v_19864 = v_3200;
assign v_19865 = ~v_16947;
assign v_19866 = ~v_3204;
assign v_19867 = v_3204;
assign v_19868 = ~v_16951;
assign v_19869 = ~v_3208;
assign v_19870 = v_19869;
assign v_19872 = v_19871;
assign v_19874 = v_19866 & v_19873;
assign v_19876 = v_16947;
assign v_19878 = v_19875 & v_19877;
assign v_19880 = v_19863 & v_19879;
assign v_19882 = v_16943;
assign v_19884 = v_19881 & v_19883;
assign v_19886 = v_19860 & v_19885;
assign v_19888 = v_16939;
assign v_19890 = v_19887 & v_19889;
assign v_19892 = v_19857 & v_19891;
assign v_19894 = v_16935;
assign v_19896 = v_19893 & v_19895;
assign v_19898 = v_19854 & v_19897;
assign v_19900 = v_16931;
assign v_19902 = v_19899 & v_19901;
assign v_19904 = v_19851 & v_19903;
assign v_19906 = v_16927;
assign v_19908 = v_19905 & v_19907;
assign v_19910 = v_19848 & v_19909;
assign v_19912 = v_16923;
assign v_19914 = v_19911 & v_19913;
assign v_19916 = v_19845 & v_19915;
assign v_19918 = v_16919;
assign v_19920 = v_19917 & v_19919;
assign v_19922 = v_19842 & v_19921;
assign v_19924 = v_16915;
assign v_19926 = v_19923 & v_19925;
assign v_19928 = v_19839 & v_19927;
assign v_19930 = v_16911;
assign v_19932 = v_19929 & v_19931;
assign v_19934 = v_19836 & v_19933;
assign v_19936 = v_16907;
assign v_19938 = v_19935 & v_19937;
assign v_19940 = v_19833 & v_19939;
assign v_19942 = v_16903;
assign v_19944 = v_19941 & v_19943;
assign v_19946 = v_19830 & v_19945;
assign v_19948 = v_3155;
assign v_19950 = v_19947 & v_19949;
assign v_19952 = v_19827 & v_19951;
assign v_19954 = v_3151;
assign v_19956 = v_19953 & v_19955;
assign v_19958 = v_19824 & v_19957;
assign v_19960 = v_3147;
assign v_19962 = v_19959 & v_19961;
assign v_19964 = v_19821 & v_19963;
assign v_19966 = v_3143;
assign v_19968 = v_19965 & v_19967;
assign v_19969 = v_19968;
assign v_19971 = v_16951;
assign v_19972 = v_3208;
assign v_19973 = v_19972;
assign v_19974 = v_19971 & v_19973;
assign v_19975 = v_19974;
assign v_19976 = v_19866 & v_19975;
assign v_19978 = v_19876 & v_19977;
assign v_19979 = v_19865 & v_19975;
assign v_19981 = v_19863 & v_19980;
assign v_19983 = v_19882 & v_19982;
assign v_19984 = v_19862 & v_19980;
assign v_19986 = v_19860 & v_19985;
assign v_19988 = v_19888 & v_19987;
assign v_19989 = v_19859 & v_19985;
assign v_19991 = v_19857 & v_19990;
assign v_19993 = v_19894 & v_19992;
assign v_19994 = v_19856 & v_19990;
assign v_19996 = v_19854 & v_19995;
assign v_19998 = v_19900 & v_19997;
assign v_19999 = v_19853 & v_19995;
assign v_20001 = v_19851 & v_20000;
assign v_20003 = v_19906 & v_20002;
assign v_20004 = v_19850 & v_20000;
assign v_20006 = v_19848 & v_20005;
assign v_20008 = v_19912 & v_20007;
assign v_20009 = v_19847 & v_20005;
assign v_20011 = v_19845 & v_20010;
assign v_20013 = v_19918 & v_20012;
assign v_20014 = v_19844 & v_20010;
assign v_20016 = v_19842 & v_20015;
assign v_20018 = v_19924 & v_20017;
assign v_20019 = v_19841 & v_20015;
assign v_20021 = v_19839 & v_20020;
assign v_20023 = v_19930 & v_20022;
assign v_20024 = v_19838 & v_20020;
assign v_20026 = v_19836 & v_20025;
assign v_20028 = v_19936 & v_20027;
assign v_20029 = v_19835 & v_20025;
assign v_20031 = v_19833 & v_20030;
assign v_20033 = v_19942 & v_20032;
assign v_20034 = v_19832 & v_20030;
assign v_20036 = v_19830 & v_20035;
assign v_20038 = v_19948 & v_20037;
assign v_20039 = v_19829 & v_20035;
assign v_20041 = v_19827 & v_20040;
assign v_20043 = v_19954 & v_20042;
assign v_20044 = v_19826 & v_20040;
assign v_20046 = v_19824 & v_20045;
assign v_20048 = v_19960 & v_20047;
assign v_20049 = v_19823 & v_20045;
assign v_20051 = v_19821 & v_20050;
assign v_20053 = v_19966 & v_20052;
assign v_20054 = v_19820 & v_20050;
assign v_20056 = v_20055;
assign v_20058 = v_19970 & v_20057;
assign v_20059 = v_20058;
assign v_20061 = v_20060;
assign v_20063 = ~v_3403;
assign v_20064 = ~v_16888;
assign v_20065 = v_16888;
assign v_20066 = ~v_3407;
assign v_20067 = ~v_16892;
assign v_20068 = v_16892;
assign v_20069 = ~v_3411;
assign v_20070 = ~v_16896;
assign v_20071 = v_16896;
assign v_20072 = ~v_3415;
assign v_20073 = ~v_16900;
assign v_20074 = v_16900;
assign v_20075 = ~v_16903;
assign v_20076 = ~v_3420;
assign v_20077 = v_3420;
assign v_20078 = ~v_16907;
assign v_20079 = ~v_3424;
assign v_20080 = v_3424;
assign v_20081 = ~v_16911;
assign v_20082 = ~v_3428;
assign v_20083 = v_3428;
assign v_20084 = ~v_16915;
assign v_20085 = ~v_3432;
assign v_20086 = v_3432;
assign v_20087 = ~v_16919;
assign v_20088 = ~v_3436;
assign v_20089 = v_3436;
assign v_20090 = ~v_16923;
assign v_20091 = ~v_3440;
assign v_20092 = v_3440;
assign v_20093 = ~v_16927;
assign v_20094 = ~v_3444;
assign v_20095 = v_3444;
assign v_20096 = ~v_16931;
assign v_20097 = ~v_3448;
assign v_20098 = v_3448;
assign v_20099 = ~v_16935;
assign v_20100 = ~v_3452;
assign v_20101 = v_3452;
assign v_20102 = ~v_16939;
assign v_20103 = ~v_3456;
assign v_20104 = v_3456;
assign v_20105 = ~v_16943;
assign v_20106 = ~v_3460;
assign v_20107 = v_3460;
assign v_20108 = ~v_16947;
assign v_20109 = ~v_3464;
assign v_20110 = v_3464;
assign v_20111 = ~v_16951;
assign v_20112 = ~v_3468;
assign v_20113 = v_20112;
assign v_20115 = v_20114;
assign v_20117 = v_20109 & v_20116;
assign v_20119 = v_16947;
assign v_20121 = v_20118 & v_20120;
assign v_20123 = v_20106 & v_20122;
assign v_20125 = v_16943;
assign v_20127 = v_20124 & v_20126;
assign v_20129 = v_20103 & v_20128;
assign v_20131 = v_16939;
assign v_20133 = v_20130 & v_20132;
assign v_20135 = v_20100 & v_20134;
assign v_20137 = v_16935;
assign v_20139 = v_20136 & v_20138;
assign v_20141 = v_20097 & v_20140;
assign v_20143 = v_16931;
assign v_20145 = v_20142 & v_20144;
assign v_20147 = v_20094 & v_20146;
assign v_20149 = v_16927;
assign v_20151 = v_20148 & v_20150;
assign v_20153 = v_20091 & v_20152;
assign v_20155 = v_16923;
assign v_20157 = v_20154 & v_20156;
assign v_20159 = v_20088 & v_20158;
assign v_20161 = v_16919;
assign v_20163 = v_20160 & v_20162;
assign v_20165 = v_20085 & v_20164;
assign v_20167 = v_16915;
assign v_20169 = v_20166 & v_20168;
assign v_20171 = v_20082 & v_20170;
assign v_20173 = v_16911;
assign v_20175 = v_20172 & v_20174;
assign v_20177 = v_20079 & v_20176;
assign v_20179 = v_16907;
assign v_20181 = v_20178 & v_20180;
assign v_20183 = v_20076 & v_20182;
assign v_20185 = v_16903;
assign v_20187 = v_20184 & v_20186;
assign v_20189 = v_20073 & v_20188;
assign v_20191 = v_3415;
assign v_20193 = v_20190 & v_20192;
assign v_20195 = v_20070 & v_20194;
assign v_20197 = v_3411;
assign v_20199 = v_20196 & v_20198;
assign v_20201 = v_20067 & v_20200;
assign v_20203 = v_3407;
assign v_20205 = v_20202 & v_20204;
assign v_20207 = v_20064 & v_20206;
assign v_20209 = v_3403;
assign v_20211 = v_20208 & v_20210;
assign v_20212 = v_20211;
assign v_20214 = v_16951;
assign v_20215 = v_3468;
assign v_20216 = v_20215;
assign v_20217 = v_20214 & v_20216;
assign v_20218 = v_20217;
assign v_20219 = v_20109 & v_20218;
assign v_20221 = v_20119 & v_20220;
assign v_20222 = v_20108 & v_20218;
assign v_20224 = v_20106 & v_20223;
assign v_20226 = v_20125 & v_20225;
assign v_20227 = v_20105 & v_20223;
assign v_20229 = v_20103 & v_20228;
assign v_20231 = v_20131 & v_20230;
assign v_20232 = v_20102 & v_20228;
assign v_20234 = v_20100 & v_20233;
assign v_20236 = v_20137 & v_20235;
assign v_20237 = v_20099 & v_20233;
assign v_20239 = v_20097 & v_20238;
assign v_20241 = v_20143 & v_20240;
assign v_20242 = v_20096 & v_20238;
assign v_20244 = v_20094 & v_20243;
assign v_20246 = v_20149 & v_20245;
assign v_20247 = v_20093 & v_20243;
assign v_20249 = v_20091 & v_20248;
assign v_20251 = v_20155 & v_20250;
assign v_20252 = v_20090 & v_20248;
assign v_20254 = v_20088 & v_20253;
assign v_20256 = v_20161 & v_20255;
assign v_20257 = v_20087 & v_20253;
assign v_20259 = v_20085 & v_20258;
assign v_20261 = v_20167 & v_20260;
assign v_20262 = v_20084 & v_20258;
assign v_20264 = v_20082 & v_20263;
assign v_20266 = v_20173 & v_20265;
assign v_20267 = v_20081 & v_20263;
assign v_20269 = v_20079 & v_20268;
assign v_20271 = v_20179 & v_20270;
assign v_20272 = v_20078 & v_20268;
assign v_20274 = v_20076 & v_20273;
assign v_20276 = v_20185 & v_20275;
assign v_20277 = v_20075 & v_20273;
assign v_20279 = v_20073 & v_20278;
assign v_20281 = v_20191 & v_20280;
assign v_20282 = v_20072 & v_20278;
assign v_20284 = v_20070 & v_20283;
assign v_20286 = v_20197 & v_20285;
assign v_20287 = v_20069 & v_20283;
assign v_20289 = v_20067 & v_20288;
assign v_20291 = v_20203 & v_20290;
assign v_20292 = v_20066 & v_20288;
assign v_20294 = v_20064 & v_20293;
assign v_20296 = v_20209 & v_20295;
assign v_20297 = v_20063 & v_20293;
assign v_20299 = v_20298;
assign v_20301 = v_20213 & v_20300;
assign v_20302 = v_20301;
assign v_20304 = v_20303;
assign v_20306 = ~v_3663;
assign v_20307 = ~v_16888;
assign v_20308 = v_16888;
assign v_20309 = ~v_3667;
assign v_20310 = ~v_16892;
assign v_20311 = v_16892;
assign v_20312 = ~v_3671;
assign v_20313 = ~v_16896;
assign v_20314 = v_16896;
assign v_20315 = ~v_3675;
assign v_20316 = ~v_16900;
assign v_20317 = v_16900;
assign v_20318 = ~v_16903;
assign v_20319 = ~v_3680;
assign v_20320 = v_3680;
assign v_20321 = ~v_16907;
assign v_20322 = ~v_3684;
assign v_20323 = v_3684;
assign v_20324 = ~v_16911;
assign v_20325 = ~v_3688;
assign v_20326 = v_3688;
assign v_20327 = ~v_16915;
assign v_20328 = ~v_3692;
assign v_20329 = v_3692;
assign v_20330 = ~v_16919;
assign v_20331 = ~v_3696;
assign v_20332 = v_3696;
assign v_20333 = ~v_16923;
assign v_20334 = ~v_3700;
assign v_20335 = v_3700;
assign v_20336 = ~v_16927;
assign v_20337 = ~v_3704;
assign v_20338 = v_3704;
assign v_20339 = ~v_16931;
assign v_20340 = ~v_3708;
assign v_20341 = v_3708;
assign v_20342 = ~v_16935;
assign v_20343 = ~v_3712;
assign v_20344 = v_3712;
assign v_20345 = ~v_16939;
assign v_20346 = ~v_3716;
assign v_20347 = v_3716;
assign v_20348 = ~v_16943;
assign v_20349 = ~v_3720;
assign v_20350 = v_3720;
assign v_20351 = ~v_16947;
assign v_20352 = ~v_3724;
assign v_20353 = v_3724;
assign v_20354 = ~v_16951;
assign v_20355 = ~v_3728;
assign v_20356 = v_20355;
assign v_20358 = v_20357;
assign v_20360 = v_20352 & v_20359;
assign v_20362 = v_16947;
assign v_20364 = v_20361 & v_20363;
assign v_20366 = v_20349 & v_20365;
assign v_20368 = v_16943;
assign v_20370 = v_20367 & v_20369;
assign v_20372 = v_20346 & v_20371;
assign v_20374 = v_16939;
assign v_20376 = v_20373 & v_20375;
assign v_20378 = v_20343 & v_20377;
assign v_20380 = v_16935;
assign v_20382 = v_20379 & v_20381;
assign v_20384 = v_20340 & v_20383;
assign v_20386 = v_16931;
assign v_20388 = v_20385 & v_20387;
assign v_20390 = v_20337 & v_20389;
assign v_20392 = v_16927;
assign v_20394 = v_20391 & v_20393;
assign v_20396 = v_20334 & v_20395;
assign v_20398 = v_16923;
assign v_20400 = v_20397 & v_20399;
assign v_20402 = v_20331 & v_20401;
assign v_20404 = v_16919;
assign v_20406 = v_20403 & v_20405;
assign v_20408 = v_20328 & v_20407;
assign v_20410 = v_16915;
assign v_20412 = v_20409 & v_20411;
assign v_20414 = v_20325 & v_20413;
assign v_20416 = v_16911;
assign v_20418 = v_20415 & v_20417;
assign v_20420 = v_20322 & v_20419;
assign v_20422 = v_16907;
assign v_20424 = v_20421 & v_20423;
assign v_20426 = v_20319 & v_20425;
assign v_20428 = v_16903;
assign v_20430 = v_20427 & v_20429;
assign v_20432 = v_20316 & v_20431;
assign v_20434 = v_3675;
assign v_20436 = v_20433 & v_20435;
assign v_20438 = v_20313 & v_20437;
assign v_20440 = v_3671;
assign v_20442 = v_20439 & v_20441;
assign v_20444 = v_20310 & v_20443;
assign v_20446 = v_3667;
assign v_20448 = v_20445 & v_20447;
assign v_20450 = v_20307 & v_20449;
assign v_20452 = v_3663;
assign v_20454 = v_20451 & v_20453;
assign v_20455 = v_20454;
assign v_20457 = v_16951;
assign v_20458 = v_3728;
assign v_20459 = v_20458;
assign v_20460 = v_20457 & v_20459;
assign v_20461 = v_20460;
assign v_20462 = v_20352 & v_20461;
assign v_20464 = v_20362 & v_20463;
assign v_20465 = v_20351 & v_20461;
assign v_20467 = v_20349 & v_20466;
assign v_20469 = v_20368 & v_20468;
assign v_20470 = v_20348 & v_20466;
assign v_20472 = v_20346 & v_20471;
assign v_20474 = v_20374 & v_20473;
assign v_20475 = v_20345 & v_20471;
assign v_20477 = v_20343 & v_20476;
assign v_20479 = v_20380 & v_20478;
assign v_20480 = v_20342 & v_20476;
assign v_20482 = v_20340 & v_20481;
assign v_20484 = v_20386 & v_20483;
assign v_20485 = v_20339 & v_20481;
assign v_20487 = v_20337 & v_20486;
assign v_20489 = v_20392 & v_20488;
assign v_20490 = v_20336 & v_20486;
assign v_20492 = v_20334 & v_20491;
assign v_20494 = v_20398 & v_20493;
assign v_20495 = v_20333 & v_20491;
assign v_20497 = v_20331 & v_20496;
assign v_20499 = v_20404 & v_20498;
assign v_20500 = v_20330 & v_20496;
assign v_20502 = v_20328 & v_20501;
assign v_20504 = v_20410 & v_20503;
assign v_20505 = v_20327 & v_20501;
assign v_20507 = v_20325 & v_20506;
assign v_20509 = v_20416 & v_20508;
assign v_20510 = v_20324 & v_20506;
assign v_20512 = v_20322 & v_20511;
assign v_20514 = v_20422 & v_20513;
assign v_20515 = v_20321 & v_20511;
assign v_20517 = v_20319 & v_20516;
assign v_20519 = v_20428 & v_20518;
assign v_20520 = v_20318 & v_20516;
assign v_20522 = v_20316 & v_20521;
assign v_20524 = v_20434 & v_20523;
assign v_20525 = v_20315 & v_20521;
assign v_20527 = v_20313 & v_20526;
assign v_20529 = v_20440 & v_20528;
assign v_20530 = v_20312 & v_20526;
assign v_20532 = v_20310 & v_20531;
assign v_20534 = v_20446 & v_20533;
assign v_20535 = v_20309 & v_20531;
assign v_20537 = v_20307 & v_20536;
assign v_20539 = v_20452 & v_20538;
assign v_20540 = v_20306 & v_20536;
assign v_20542 = v_20541;
assign v_20544 = v_20456 & v_20543;
assign v_20545 = v_20544;
assign v_20547 = v_20546;
assign v_20549 = ~v_3923;
assign v_20550 = ~v_16888;
assign v_20551 = v_16888;
assign v_20552 = ~v_3927;
assign v_20553 = ~v_16892;
assign v_20554 = v_16892;
assign v_20555 = ~v_3931;
assign v_20556 = ~v_16896;
assign v_20557 = v_16896;
assign v_20558 = ~v_3935;
assign v_20559 = ~v_16900;
assign v_20560 = v_16900;
assign v_20561 = ~v_16903;
assign v_20562 = ~v_3940;
assign v_20563 = v_3940;
assign v_20564 = ~v_16907;
assign v_20565 = ~v_3944;
assign v_20566 = v_3944;
assign v_20567 = ~v_16911;
assign v_20568 = ~v_3948;
assign v_20569 = v_3948;
assign v_20570 = ~v_16915;
assign v_20571 = ~v_3952;
assign v_20572 = v_3952;
assign v_20573 = ~v_16919;
assign v_20574 = ~v_3956;
assign v_20575 = v_3956;
assign v_20576 = ~v_16923;
assign v_20577 = ~v_3960;
assign v_20578 = v_3960;
assign v_20579 = ~v_16927;
assign v_20580 = ~v_3964;
assign v_20581 = v_3964;
assign v_20582 = ~v_16931;
assign v_20583 = ~v_3968;
assign v_20584 = v_3968;
assign v_20585 = ~v_16935;
assign v_20586 = ~v_3972;
assign v_20587 = v_3972;
assign v_20588 = ~v_16939;
assign v_20589 = ~v_3976;
assign v_20590 = v_3976;
assign v_20591 = ~v_16943;
assign v_20592 = ~v_3980;
assign v_20593 = v_3980;
assign v_20594 = ~v_16947;
assign v_20595 = ~v_3984;
assign v_20596 = v_3984;
assign v_20597 = ~v_16951;
assign v_20598 = ~v_3988;
assign v_20599 = v_20598;
assign v_20601 = v_20600;
assign v_20603 = v_20595 & v_20602;
assign v_20605 = v_16947;
assign v_20607 = v_20604 & v_20606;
assign v_20609 = v_20592 & v_20608;
assign v_20611 = v_16943;
assign v_20613 = v_20610 & v_20612;
assign v_20615 = v_20589 & v_20614;
assign v_20617 = v_16939;
assign v_20619 = v_20616 & v_20618;
assign v_20621 = v_20586 & v_20620;
assign v_20623 = v_16935;
assign v_20625 = v_20622 & v_20624;
assign v_20627 = v_20583 & v_20626;
assign v_20629 = v_16931;
assign v_20631 = v_20628 & v_20630;
assign v_20633 = v_20580 & v_20632;
assign v_20635 = v_16927;
assign v_20637 = v_20634 & v_20636;
assign v_20639 = v_20577 & v_20638;
assign v_20641 = v_16923;
assign v_20643 = v_20640 & v_20642;
assign v_20645 = v_20574 & v_20644;
assign v_20647 = v_16919;
assign v_20649 = v_20646 & v_20648;
assign v_20651 = v_20571 & v_20650;
assign v_20653 = v_16915;
assign v_20655 = v_20652 & v_20654;
assign v_20657 = v_20568 & v_20656;
assign v_20659 = v_16911;
assign v_20661 = v_20658 & v_20660;
assign v_20663 = v_20565 & v_20662;
assign v_20665 = v_16907;
assign v_20667 = v_20664 & v_20666;
assign v_20669 = v_20562 & v_20668;
assign v_20671 = v_16903;
assign v_20673 = v_20670 & v_20672;
assign v_20675 = v_20559 & v_20674;
assign v_20677 = v_3935;
assign v_20679 = v_20676 & v_20678;
assign v_20681 = v_20556 & v_20680;
assign v_20683 = v_3931;
assign v_20685 = v_20682 & v_20684;
assign v_20687 = v_20553 & v_20686;
assign v_20689 = v_3927;
assign v_20691 = v_20688 & v_20690;
assign v_20693 = v_20550 & v_20692;
assign v_20695 = v_3923;
assign v_20697 = v_20694 & v_20696;
assign v_20698 = v_20697;
assign v_20700 = v_16951;
assign v_20701 = v_3988;
assign v_20702 = v_20701;
assign v_20703 = v_20700 & v_20702;
assign v_20704 = v_20703;
assign v_20705 = v_20595 & v_20704;
assign v_20707 = v_20605 & v_20706;
assign v_20708 = v_20594 & v_20704;
assign v_20710 = v_20592 & v_20709;
assign v_20712 = v_20611 & v_20711;
assign v_20713 = v_20591 & v_20709;
assign v_20715 = v_20589 & v_20714;
assign v_20717 = v_20617 & v_20716;
assign v_20718 = v_20588 & v_20714;
assign v_20720 = v_20586 & v_20719;
assign v_20722 = v_20623 & v_20721;
assign v_20723 = v_20585 & v_20719;
assign v_20725 = v_20583 & v_20724;
assign v_20727 = v_20629 & v_20726;
assign v_20728 = v_20582 & v_20724;
assign v_20730 = v_20580 & v_20729;
assign v_20732 = v_20635 & v_20731;
assign v_20733 = v_20579 & v_20729;
assign v_20735 = v_20577 & v_20734;
assign v_20737 = v_20641 & v_20736;
assign v_20738 = v_20576 & v_20734;
assign v_20740 = v_20574 & v_20739;
assign v_20742 = v_20647 & v_20741;
assign v_20743 = v_20573 & v_20739;
assign v_20745 = v_20571 & v_20744;
assign v_20747 = v_20653 & v_20746;
assign v_20748 = v_20570 & v_20744;
assign v_20750 = v_20568 & v_20749;
assign v_20752 = v_20659 & v_20751;
assign v_20753 = v_20567 & v_20749;
assign v_20755 = v_20565 & v_20754;
assign v_20757 = v_20665 & v_20756;
assign v_20758 = v_20564 & v_20754;
assign v_20760 = v_20562 & v_20759;
assign v_20762 = v_20671 & v_20761;
assign v_20763 = v_20561 & v_20759;
assign v_20765 = v_20559 & v_20764;
assign v_20767 = v_20677 & v_20766;
assign v_20768 = v_20558 & v_20764;
assign v_20770 = v_20556 & v_20769;
assign v_20772 = v_20683 & v_20771;
assign v_20773 = v_20555 & v_20769;
assign v_20775 = v_20553 & v_20774;
assign v_20777 = v_20689 & v_20776;
assign v_20778 = v_20552 & v_20774;
assign v_20780 = v_20550 & v_20779;
assign v_20782 = v_20695 & v_20781;
assign v_20783 = v_20549 & v_20779;
assign v_20785 = v_20784;
assign v_20787 = v_20699 & v_20786;
assign v_20788 = v_20787;
assign v_20790 = v_20789;
assign v_20791 = ~v_4182;
assign v_20792 = ~v_16888;
assign v_20793 = v_16888;
assign v_20794 = ~v_4186;
assign v_20795 = ~v_16892;
assign v_20796 = v_16892;
assign v_20797 = ~v_4190;
assign v_20798 = ~v_16896;
assign v_20799 = v_16896;
assign v_20800 = ~v_4194;
assign v_20801 = ~v_16900;
assign v_20802 = v_16900;
assign v_20803 = ~v_16903;
assign v_20804 = ~v_4199;
assign v_20805 = v_4199;
assign v_20806 = ~v_16907;
assign v_20807 = ~v_4203;
assign v_20808 = v_4203;
assign v_20809 = ~v_16911;
assign v_20810 = ~v_4207;
assign v_20811 = v_4207;
assign v_20812 = ~v_16915;
assign v_20813 = ~v_4211;
assign v_20814 = v_4211;
assign v_20815 = ~v_16919;
assign v_20816 = ~v_4215;
assign v_20817 = v_4215;
assign v_20818 = ~v_16923;
assign v_20819 = ~v_4219;
assign v_20820 = v_4219;
assign v_20821 = ~v_16927;
assign v_20822 = ~v_4223;
assign v_20823 = v_4223;
assign v_20824 = ~v_16931;
assign v_20825 = ~v_4227;
assign v_20826 = v_4227;
assign v_20827 = ~v_16935;
assign v_20828 = ~v_4231;
assign v_20829 = v_4231;
assign v_20830 = ~v_16939;
assign v_20831 = ~v_4235;
assign v_20832 = v_4235;
assign v_20833 = ~v_16943;
assign v_20834 = ~v_4239;
assign v_20835 = v_4239;
assign v_20836 = ~v_16947;
assign v_20837 = ~v_4243;
assign v_20838 = v_4243;
assign v_20839 = ~v_16951;
assign v_20840 = ~v_4247;
assign v_20841 = v_20840;
assign v_20843 = v_20842;
assign v_20845 = v_20837 & v_20844;
assign v_20847 = v_16947;
assign v_20849 = v_20846 & v_20848;
assign v_20851 = v_20834 & v_20850;
assign v_20853 = v_16943;
assign v_20855 = v_20852 & v_20854;
assign v_20857 = v_20831 & v_20856;
assign v_20859 = v_16939;
assign v_20861 = v_20858 & v_20860;
assign v_20863 = v_20828 & v_20862;
assign v_20865 = v_16935;
assign v_20867 = v_20864 & v_20866;
assign v_20869 = v_20825 & v_20868;
assign v_20871 = v_16931;
assign v_20873 = v_20870 & v_20872;
assign v_20875 = v_20822 & v_20874;
assign v_20877 = v_16927;
assign v_20879 = v_20876 & v_20878;
assign v_20881 = v_20819 & v_20880;
assign v_20883 = v_16923;
assign v_20885 = v_20882 & v_20884;
assign v_20887 = v_20816 & v_20886;
assign v_20889 = v_16919;
assign v_20891 = v_20888 & v_20890;
assign v_20893 = v_20813 & v_20892;
assign v_20895 = v_16915;
assign v_20897 = v_20894 & v_20896;
assign v_20899 = v_20810 & v_20898;
assign v_20901 = v_16911;
assign v_20903 = v_20900 & v_20902;
assign v_20905 = v_20807 & v_20904;
assign v_20907 = v_16907;
assign v_20909 = v_20906 & v_20908;
assign v_20911 = v_20804 & v_20910;
assign v_20913 = v_16903;
assign v_20915 = v_20912 & v_20914;
assign v_20917 = v_20801 & v_20916;
assign v_20919 = v_4194;
assign v_20921 = v_20918 & v_20920;
assign v_20923 = v_20798 & v_20922;
assign v_20925 = v_4190;
assign v_20927 = v_20924 & v_20926;
assign v_20929 = v_20795 & v_20928;
assign v_20931 = v_4186;
assign v_20933 = v_20930 & v_20932;
assign v_20935 = v_20792 & v_20934;
assign v_20937 = v_4182;
assign v_20939 = v_20936 & v_20938;
assign v_20941 = ~v_20940;
assign v_20943 = v_16951;
assign v_20944 = v_4247;
assign v_20945 = v_20944;
assign v_20946 = v_20943 & v_20945;
assign v_20947 = v_20946;
assign v_20948 = v_20837 & v_20947;
assign v_20950 = v_20847 & v_20949;
assign v_20951 = v_20836 & v_20947;
assign v_20953 = v_20834 & v_20952;
assign v_20955 = v_20853 & v_20954;
assign v_20956 = v_20833 & v_20952;
assign v_20958 = v_20831 & v_20957;
assign v_20960 = v_20859 & v_20959;
assign v_20961 = v_20830 & v_20957;
assign v_20963 = v_20828 & v_20962;
assign v_20965 = v_20865 & v_20964;
assign v_20966 = v_20827 & v_20962;
assign v_20968 = v_20825 & v_20967;
assign v_20970 = v_20871 & v_20969;
assign v_20971 = v_20824 & v_20967;
assign v_20973 = v_20822 & v_20972;
assign v_20975 = v_20877 & v_20974;
assign v_20976 = v_20821 & v_20972;
assign v_20978 = v_20819 & v_20977;
assign v_20980 = v_20883 & v_20979;
assign v_20981 = v_20818 & v_20977;
assign v_20983 = v_20816 & v_20982;
assign v_20985 = v_20889 & v_20984;
assign v_20986 = v_20815 & v_20982;
assign v_20988 = v_20813 & v_20987;
assign v_20990 = v_20895 & v_20989;
assign v_20991 = v_20812 & v_20987;
assign v_20993 = v_20810 & v_20992;
assign v_20995 = v_20901 & v_20994;
assign v_20996 = v_20809 & v_20992;
assign v_20998 = v_20807 & v_20997;
assign v_21000 = v_20907 & v_20999;
assign v_21001 = v_20806 & v_20997;
assign v_21003 = v_20804 & v_21002;
assign v_21005 = v_20913 & v_21004;
assign v_21006 = v_20803 & v_21002;
assign v_21008 = v_20801 & v_21007;
assign v_21010 = v_20919 & v_21009;
assign v_21011 = v_20800 & v_21007;
assign v_21013 = v_20798 & v_21012;
assign v_21015 = v_20925 & v_21014;
assign v_21016 = v_20797 & v_21012;
assign v_21018 = v_20795 & v_21017;
assign v_21020 = v_20931 & v_21019;
assign v_21021 = v_20794 & v_21017;
assign v_21023 = v_20792 & v_21022;
assign v_21025 = v_20937 & v_21024;
assign v_21026 = v_20791 & v_21022;
assign v_21028 = v_20940;
assign v_21030 = v_20942 & v_21029;
assign v_21031 = v_21030;
assign v_21033 = v_21032;
assign v_21035 = ~v_6;
assign v_21037 = ~v_21036;
assign v_21038 = v_21036;
assign v_21039 = ~v_13;
assign v_21041 = ~v_21040;
assign v_21042 = v_21040;
assign v_21043 = ~v_18;
assign v_21045 = ~v_21044;
assign v_21046 = v_21044;
assign v_21047 = ~v_23;
assign v_21049 = ~v_21048;
assign v_21050 = v_21048;
assign v_21052 = ~v_21051;
assign v_21053 = ~v_30;
assign v_21054 = v_30;
assign v_21056 = ~v_21055;
assign v_21057 = ~v_35;
assign v_21058 = v_35;
assign v_21060 = ~v_21059;
assign v_21061 = ~v_40;
assign v_21062 = v_40;
assign v_21064 = ~v_21063;
assign v_21065 = ~v_45;
assign v_21066 = v_45;
assign v_21068 = ~v_21067;
assign v_21069 = ~v_50;
assign v_21070 = v_50;
assign v_21072 = ~v_21071;
assign v_21073 = ~v_55;
assign v_21074 = v_55;
assign v_21076 = ~v_21075;
assign v_21077 = ~v_60;
assign v_21078 = v_60;
assign v_21080 = ~v_21079;
assign v_21081 = ~v_65;
assign v_21082 = v_65;
assign v_21084 = ~v_21083;
assign v_21085 = ~v_70;
assign v_21086 = v_70;
assign v_21088 = ~v_21087;
assign v_21089 = ~v_75;
assign v_21090 = v_75;
assign v_21092 = ~v_21091;
assign v_21093 = ~v_80;
assign v_21094 = v_80;
assign v_21096 = ~v_21095;
assign v_21097 = ~v_85;
assign v_21098 = v_85;
assign v_21100 = ~v_21099;
assign v_21101 = ~v_90;
assign v_21102 = v_21101;
assign v_21104 = v_21103;
assign v_21106 = v_21097 & v_21105;
assign v_21108 = v_21095;
assign v_21110 = v_21107 & v_21109;
assign v_21112 = v_21093 & v_21111;
assign v_21114 = v_21091;
assign v_21116 = v_21113 & v_21115;
assign v_21118 = v_21089 & v_21117;
assign v_21120 = v_21087;
assign v_21122 = v_21119 & v_21121;
assign v_21124 = v_21085 & v_21123;
assign v_21126 = v_21083;
assign v_21128 = v_21125 & v_21127;
assign v_21130 = v_21081 & v_21129;
assign v_21132 = v_21079;
assign v_21134 = v_21131 & v_21133;
assign v_21136 = v_21077 & v_21135;
assign v_21138 = v_21075;
assign v_21140 = v_21137 & v_21139;
assign v_21142 = v_21073 & v_21141;
assign v_21144 = v_21071;
assign v_21146 = v_21143 & v_21145;
assign v_21148 = v_21069 & v_21147;
assign v_21150 = v_21067;
assign v_21152 = v_21149 & v_21151;
assign v_21154 = v_21065 & v_21153;
assign v_21156 = v_21063;
assign v_21158 = v_21155 & v_21157;
assign v_21160 = v_21061 & v_21159;
assign v_21162 = v_21059;
assign v_21164 = v_21161 & v_21163;
assign v_21166 = v_21057 & v_21165;
assign v_21168 = v_21055;
assign v_21170 = v_21167 & v_21169;
assign v_21172 = v_21053 & v_21171;
assign v_21174 = v_21051;
assign v_21176 = v_21173 & v_21175;
assign v_21178 = v_21049 & v_21177;
assign v_21180 = v_23;
assign v_21182 = v_21179 & v_21181;
assign v_21184 = v_21045 & v_21183;
assign v_21186 = v_18;
assign v_21188 = v_21185 & v_21187;
assign v_21190 = v_21041 & v_21189;
assign v_21192 = v_13;
assign v_21194 = v_21191 & v_21193;
assign v_21196 = v_21037 & v_21195;
assign v_21198 = v_6;
assign v_21200 = v_21197 & v_21199;
assign v_21201 = v_21200;
assign v_21203 = v_21099;
assign v_21204 = v_90;
assign v_21205 = v_21204;
assign v_21206 = v_21203 & v_21205;
assign v_21207 = v_21206;
assign v_21208 = v_21097 & v_21207;
assign v_21210 = v_21108 & v_21209;
assign v_21211 = v_21096 & v_21207;
assign v_21213 = v_21093 & v_21212;
assign v_21215 = v_21114 & v_21214;
assign v_21216 = v_21092 & v_21212;
assign v_21218 = v_21089 & v_21217;
assign v_21220 = v_21120 & v_21219;
assign v_21221 = v_21088 & v_21217;
assign v_21223 = v_21085 & v_21222;
assign v_21225 = v_21126 & v_21224;
assign v_21226 = v_21084 & v_21222;
assign v_21228 = v_21081 & v_21227;
assign v_21230 = v_21132 & v_21229;
assign v_21231 = v_21080 & v_21227;
assign v_21233 = v_21077 & v_21232;
assign v_21235 = v_21138 & v_21234;
assign v_21236 = v_21076 & v_21232;
assign v_21238 = v_21073 & v_21237;
assign v_21240 = v_21144 & v_21239;
assign v_21241 = v_21072 & v_21237;
assign v_21243 = v_21069 & v_21242;
assign v_21245 = v_21150 & v_21244;
assign v_21246 = v_21068 & v_21242;
assign v_21248 = v_21065 & v_21247;
assign v_21250 = v_21156 & v_21249;
assign v_21251 = v_21064 & v_21247;
assign v_21253 = v_21061 & v_21252;
assign v_21255 = v_21162 & v_21254;
assign v_21256 = v_21060 & v_21252;
assign v_21258 = v_21057 & v_21257;
assign v_21260 = v_21168 & v_21259;
assign v_21261 = v_21056 & v_21257;
assign v_21263 = v_21053 & v_21262;
assign v_21265 = v_21174 & v_21264;
assign v_21266 = v_21052 & v_21262;
assign v_21268 = v_21049 & v_21267;
assign v_21270 = v_21180 & v_21269;
assign v_21271 = v_21047 & v_21267;
assign v_21273 = v_21045 & v_21272;
assign v_21275 = v_21186 & v_21274;
assign v_21276 = v_21043 & v_21272;
assign v_21278 = v_21041 & v_21277;
assign v_21280 = v_21192 & v_21279;
assign v_21281 = v_21039 & v_21277;
assign v_21283 = v_21037 & v_21282;
assign v_21285 = v_21198 & v_21284;
assign v_21286 = v_21035 & v_21282;
assign v_21288 = v_21287;
assign v_21290 = v_21202 & v_21289;
assign v_21291 = v_21290;
assign v_21293 = v_21292;
assign v_21295 = ~v_283;
assign v_21296 = ~v_21036;
assign v_21297 = v_21036;
assign v_21298 = ~v_287;
assign v_21299 = ~v_21040;
assign v_21300 = v_21040;
assign v_21301 = ~v_291;
assign v_21302 = ~v_21044;
assign v_21303 = v_21044;
assign v_21304 = ~v_295;
assign v_21305 = ~v_21048;
assign v_21306 = v_21048;
assign v_21307 = ~v_21051;
assign v_21308 = ~v_300;
assign v_21309 = v_300;
assign v_21310 = ~v_21055;
assign v_21311 = ~v_304;
assign v_21312 = v_304;
assign v_21313 = ~v_21059;
assign v_21314 = ~v_308;
assign v_21315 = v_308;
assign v_21316 = ~v_21063;
assign v_21317 = ~v_312;
assign v_21318 = v_312;
assign v_21319 = ~v_21067;
assign v_21320 = ~v_316;
assign v_21321 = v_316;
assign v_21322 = ~v_21071;
assign v_21323 = ~v_320;
assign v_21324 = v_320;
assign v_21325 = ~v_21075;
assign v_21326 = ~v_324;
assign v_21327 = v_324;
assign v_21328 = ~v_21079;
assign v_21329 = ~v_328;
assign v_21330 = v_328;
assign v_21331 = ~v_21083;
assign v_21332 = ~v_332;
assign v_21333 = v_332;
assign v_21334 = ~v_21087;
assign v_21335 = ~v_336;
assign v_21336 = v_336;
assign v_21337 = ~v_21091;
assign v_21338 = ~v_340;
assign v_21339 = v_340;
assign v_21340 = ~v_21095;
assign v_21341 = ~v_344;
assign v_21342 = v_344;
assign v_21343 = ~v_21099;
assign v_21344 = ~v_348;
assign v_21345 = v_21344;
assign v_21347 = v_21346;
assign v_21349 = v_21341 & v_21348;
assign v_21351 = v_21095;
assign v_21353 = v_21350 & v_21352;
assign v_21355 = v_21338 & v_21354;
assign v_21357 = v_21091;
assign v_21359 = v_21356 & v_21358;
assign v_21361 = v_21335 & v_21360;
assign v_21363 = v_21087;
assign v_21365 = v_21362 & v_21364;
assign v_21367 = v_21332 & v_21366;
assign v_21369 = v_21083;
assign v_21371 = v_21368 & v_21370;
assign v_21373 = v_21329 & v_21372;
assign v_21375 = v_21079;
assign v_21377 = v_21374 & v_21376;
assign v_21379 = v_21326 & v_21378;
assign v_21381 = v_21075;
assign v_21383 = v_21380 & v_21382;
assign v_21385 = v_21323 & v_21384;
assign v_21387 = v_21071;
assign v_21389 = v_21386 & v_21388;
assign v_21391 = v_21320 & v_21390;
assign v_21393 = v_21067;
assign v_21395 = v_21392 & v_21394;
assign v_21397 = v_21317 & v_21396;
assign v_21399 = v_21063;
assign v_21401 = v_21398 & v_21400;
assign v_21403 = v_21314 & v_21402;
assign v_21405 = v_21059;
assign v_21407 = v_21404 & v_21406;
assign v_21409 = v_21311 & v_21408;
assign v_21411 = v_21055;
assign v_21413 = v_21410 & v_21412;
assign v_21415 = v_21308 & v_21414;
assign v_21417 = v_21051;
assign v_21419 = v_21416 & v_21418;
assign v_21421 = v_21305 & v_21420;
assign v_21423 = v_295;
assign v_21425 = v_21422 & v_21424;
assign v_21427 = v_21302 & v_21426;
assign v_21429 = v_291;
assign v_21431 = v_21428 & v_21430;
assign v_21433 = v_21299 & v_21432;
assign v_21435 = v_287;
assign v_21437 = v_21434 & v_21436;
assign v_21439 = v_21296 & v_21438;
assign v_21441 = v_283;
assign v_21443 = v_21440 & v_21442;
assign v_21444 = v_21443;
assign v_21446 = v_21099;
assign v_21447 = v_348;
assign v_21448 = v_21447;
assign v_21449 = v_21446 & v_21448;
assign v_21450 = v_21449;
assign v_21451 = v_21341 & v_21450;
assign v_21453 = v_21351 & v_21452;
assign v_21454 = v_21340 & v_21450;
assign v_21456 = v_21338 & v_21455;
assign v_21458 = v_21357 & v_21457;
assign v_21459 = v_21337 & v_21455;
assign v_21461 = v_21335 & v_21460;
assign v_21463 = v_21363 & v_21462;
assign v_21464 = v_21334 & v_21460;
assign v_21466 = v_21332 & v_21465;
assign v_21468 = v_21369 & v_21467;
assign v_21469 = v_21331 & v_21465;
assign v_21471 = v_21329 & v_21470;
assign v_21473 = v_21375 & v_21472;
assign v_21474 = v_21328 & v_21470;
assign v_21476 = v_21326 & v_21475;
assign v_21478 = v_21381 & v_21477;
assign v_21479 = v_21325 & v_21475;
assign v_21481 = v_21323 & v_21480;
assign v_21483 = v_21387 & v_21482;
assign v_21484 = v_21322 & v_21480;
assign v_21486 = v_21320 & v_21485;
assign v_21488 = v_21393 & v_21487;
assign v_21489 = v_21319 & v_21485;
assign v_21491 = v_21317 & v_21490;
assign v_21493 = v_21399 & v_21492;
assign v_21494 = v_21316 & v_21490;
assign v_21496 = v_21314 & v_21495;
assign v_21498 = v_21405 & v_21497;
assign v_21499 = v_21313 & v_21495;
assign v_21501 = v_21311 & v_21500;
assign v_21503 = v_21411 & v_21502;
assign v_21504 = v_21310 & v_21500;
assign v_21506 = v_21308 & v_21505;
assign v_21508 = v_21417 & v_21507;
assign v_21509 = v_21307 & v_21505;
assign v_21511 = v_21305 & v_21510;
assign v_21513 = v_21423 & v_21512;
assign v_21514 = v_21304 & v_21510;
assign v_21516 = v_21302 & v_21515;
assign v_21518 = v_21429 & v_21517;
assign v_21519 = v_21301 & v_21515;
assign v_21521 = v_21299 & v_21520;
assign v_21523 = v_21435 & v_21522;
assign v_21524 = v_21298 & v_21520;
assign v_21526 = v_21296 & v_21525;
assign v_21528 = v_21441 & v_21527;
assign v_21529 = v_21295 & v_21525;
assign v_21531 = v_21530;
assign v_21533 = v_21445 & v_21532;
assign v_21534 = v_21533;
assign v_21536 = v_21535;
assign v_21538 = ~v_543;
assign v_21539 = ~v_21036;
assign v_21540 = v_21036;
assign v_21541 = ~v_547;
assign v_21542 = ~v_21040;
assign v_21543 = v_21040;
assign v_21544 = ~v_551;
assign v_21545 = ~v_21044;
assign v_21546 = v_21044;
assign v_21547 = ~v_555;
assign v_21548 = ~v_21048;
assign v_21549 = v_21048;
assign v_21550 = ~v_21051;
assign v_21551 = ~v_560;
assign v_21552 = v_560;
assign v_21553 = ~v_21055;
assign v_21554 = ~v_564;
assign v_21555 = v_564;
assign v_21556 = ~v_21059;
assign v_21557 = ~v_568;
assign v_21558 = v_568;
assign v_21559 = ~v_21063;
assign v_21560 = ~v_572;
assign v_21561 = v_572;
assign v_21562 = ~v_21067;
assign v_21563 = ~v_576;
assign v_21564 = v_576;
assign v_21565 = ~v_21071;
assign v_21566 = ~v_580;
assign v_21567 = v_580;
assign v_21568 = ~v_21075;
assign v_21569 = ~v_584;
assign v_21570 = v_584;
assign v_21571 = ~v_21079;
assign v_21572 = ~v_588;
assign v_21573 = v_588;
assign v_21574 = ~v_21083;
assign v_21575 = ~v_592;
assign v_21576 = v_592;
assign v_21577 = ~v_21087;
assign v_21578 = ~v_596;
assign v_21579 = v_596;
assign v_21580 = ~v_21091;
assign v_21581 = ~v_600;
assign v_21582 = v_600;
assign v_21583 = ~v_21095;
assign v_21584 = ~v_604;
assign v_21585 = v_604;
assign v_21586 = ~v_21099;
assign v_21587 = ~v_608;
assign v_21588 = v_21587;
assign v_21590 = v_21589;
assign v_21592 = v_21584 & v_21591;
assign v_21594 = v_21095;
assign v_21596 = v_21593 & v_21595;
assign v_21598 = v_21581 & v_21597;
assign v_21600 = v_21091;
assign v_21602 = v_21599 & v_21601;
assign v_21604 = v_21578 & v_21603;
assign v_21606 = v_21087;
assign v_21608 = v_21605 & v_21607;
assign v_21610 = v_21575 & v_21609;
assign v_21612 = v_21083;
assign v_21614 = v_21611 & v_21613;
assign v_21616 = v_21572 & v_21615;
assign v_21618 = v_21079;
assign v_21620 = v_21617 & v_21619;
assign v_21622 = v_21569 & v_21621;
assign v_21624 = v_21075;
assign v_21626 = v_21623 & v_21625;
assign v_21628 = v_21566 & v_21627;
assign v_21630 = v_21071;
assign v_21632 = v_21629 & v_21631;
assign v_21634 = v_21563 & v_21633;
assign v_21636 = v_21067;
assign v_21638 = v_21635 & v_21637;
assign v_21640 = v_21560 & v_21639;
assign v_21642 = v_21063;
assign v_21644 = v_21641 & v_21643;
assign v_21646 = v_21557 & v_21645;
assign v_21648 = v_21059;
assign v_21650 = v_21647 & v_21649;
assign v_21652 = v_21554 & v_21651;
assign v_21654 = v_21055;
assign v_21656 = v_21653 & v_21655;
assign v_21658 = v_21551 & v_21657;
assign v_21660 = v_21051;
assign v_21662 = v_21659 & v_21661;
assign v_21664 = v_21548 & v_21663;
assign v_21666 = v_555;
assign v_21668 = v_21665 & v_21667;
assign v_21670 = v_21545 & v_21669;
assign v_21672 = v_551;
assign v_21674 = v_21671 & v_21673;
assign v_21676 = v_21542 & v_21675;
assign v_21678 = v_547;
assign v_21680 = v_21677 & v_21679;
assign v_21682 = v_21539 & v_21681;
assign v_21684 = v_543;
assign v_21686 = v_21683 & v_21685;
assign v_21687 = v_21686;
assign v_21689 = v_21099;
assign v_21690 = v_608;
assign v_21691 = v_21690;
assign v_21692 = v_21689 & v_21691;
assign v_21693 = v_21692;
assign v_21694 = v_21584 & v_21693;
assign v_21696 = v_21594 & v_21695;
assign v_21697 = v_21583 & v_21693;
assign v_21699 = v_21581 & v_21698;
assign v_21701 = v_21600 & v_21700;
assign v_21702 = v_21580 & v_21698;
assign v_21704 = v_21578 & v_21703;
assign v_21706 = v_21606 & v_21705;
assign v_21707 = v_21577 & v_21703;
assign v_21709 = v_21575 & v_21708;
assign v_21711 = v_21612 & v_21710;
assign v_21712 = v_21574 & v_21708;
assign v_21714 = v_21572 & v_21713;
assign v_21716 = v_21618 & v_21715;
assign v_21717 = v_21571 & v_21713;
assign v_21719 = v_21569 & v_21718;
assign v_21721 = v_21624 & v_21720;
assign v_21722 = v_21568 & v_21718;
assign v_21724 = v_21566 & v_21723;
assign v_21726 = v_21630 & v_21725;
assign v_21727 = v_21565 & v_21723;
assign v_21729 = v_21563 & v_21728;
assign v_21731 = v_21636 & v_21730;
assign v_21732 = v_21562 & v_21728;
assign v_21734 = v_21560 & v_21733;
assign v_21736 = v_21642 & v_21735;
assign v_21737 = v_21559 & v_21733;
assign v_21739 = v_21557 & v_21738;
assign v_21741 = v_21648 & v_21740;
assign v_21742 = v_21556 & v_21738;
assign v_21744 = v_21554 & v_21743;
assign v_21746 = v_21654 & v_21745;
assign v_21747 = v_21553 & v_21743;
assign v_21749 = v_21551 & v_21748;
assign v_21751 = v_21660 & v_21750;
assign v_21752 = v_21550 & v_21748;
assign v_21754 = v_21548 & v_21753;
assign v_21756 = v_21666 & v_21755;
assign v_21757 = v_21547 & v_21753;
assign v_21759 = v_21545 & v_21758;
assign v_21761 = v_21672 & v_21760;
assign v_21762 = v_21544 & v_21758;
assign v_21764 = v_21542 & v_21763;
assign v_21766 = v_21678 & v_21765;
assign v_21767 = v_21541 & v_21763;
assign v_21769 = v_21539 & v_21768;
assign v_21771 = v_21684 & v_21770;
assign v_21772 = v_21538 & v_21768;
assign v_21774 = v_21773;
assign v_21776 = v_21688 & v_21775;
assign v_21777 = v_21776;
assign v_21779 = v_21778;
assign v_21781 = ~v_803;
assign v_21782 = ~v_21036;
assign v_21783 = v_21036;
assign v_21784 = ~v_807;
assign v_21785 = ~v_21040;
assign v_21786 = v_21040;
assign v_21787 = ~v_811;
assign v_21788 = ~v_21044;
assign v_21789 = v_21044;
assign v_21790 = ~v_815;
assign v_21791 = ~v_21048;
assign v_21792 = v_21048;
assign v_21793 = ~v_21051;
assign v_21794 = ~v_820;
assign v_21795 = v_820;
assign v_21796 = ~v_21055;
assign v_21797 = ~v_824;
assign v_21798 = v_824;
assign v_21799 = ~v_21059;
assign v_21800 = ~v_828;
assign v_21801 = v_828;
assign v_21802 = ~v_21063;
assign v_21803 = ~v_832;
assign v_21804 = v_832;
assign v_21805 = ~v_21067;
assign v_21806 = ~v_836;
assign v_21807 = v_836;
assign v_21808 = ~v_21071;
assign v_21809 = ~v_840;
assign v_21810 = v_840;
assign v_21811 = ~v_21075;
assign v_21812 = ~v_844;
assign v_21813 = v_844;
assign v_21814 = ~v_21079;
assign v_21815 = ~v_848;
assign v_21816 = v_848;
assign v_21817 = ~v_21083;
assign v_21818 = ~v_852;
assign v_21819 = v_852;
assign v_21820 = ~v_21087;
assign v_21821 = ~v_856;
assign v_21822 = v_856;
assign v_21823 = ~v_21091;
assign v_21824 = ~v_860;
assign v_21825 = v_860;
assign v_21826 = ~v_21095;
assign v_21827 = ~v_864;
assign v_21828 = v_864;
assign v_21829 = ~v_21099;
assign v_21830 = ~v_868;
assign v_21831 = v_21830;
assign v_21833 = v_21832;
assign v_21835 = v_21827 & v_21834;
assign v_21837 = v_21095;
assign v_21839 = v_21836 & v_21838;
assign v_21841 = v_21824 & v_21840;
assign v_21843 = v_21091;
assign v_21845 = v_21842 & v_21844;
assign v_21847 = v_21821 & v_21846;
assign v_21849 = v_21087;
assign v_21851 = v_21848 & v_21850;
assign v_21853 = v_21818 & v_21852;
assign v_21855 = v_21083;
assign v_21857 = v_21854 & v_21856;
assign v_21859 = v_21815 & v_21858;
assign v_21861 = v_21079;
assign v_21863 = v_21860 & v_21862;
assign v_21865 = v_21812 & v_21864;
assign v_21867 = v_21075;
assign v_21869 = v_21866 & v_21868;
assign v_21871 = v_21809 & v_21870;
assign v_21873 = v_21071;
assign v_21875 = v_21872 & v_21874;
assign v_21877 = v_21806 & v_21876;
assign v_21879 = v_21067;
assign v_21881 = v_21878 & v_21880;
assign v_21883 = v_21803 & v_21882;
assign v_21885 = v_21063;
assign v_21887 = v_21884 & v_21886;
assign v_21889 = v_21800 & v_21888;
assign v_21891 = v_21059;
assign v_21893 = v_21890 & v_21892;
assign v_21895 = v_21797 & v_21894;
assign v_21897 = v_21055;
assign v_21899 = v_21896 & v_21898;
assign v_21901 = v_21794 & v_21900;
assign v_21903 = v_21051;
assign v_21905 = v_21902 & v_21904;
assign v_21907 = v_21791 & v_21906;
assign v_21909 = v_815;
assign v_21911 = v_21908 & v_21910;
assign v_21913 = v_21788 & v_21912;
assign v_21915 = v_811;
assign v_21917 = v_21914 & v_21916;
assign v_21919 = v_21785 & v_21918;
assign v_21921 = v_807;
assign v_21923 = v_21920 & v_21922;
assign v_21925 = v_21782 & v_21924;
assign v_21927 = v_803;
assign v_21929 = v_21926 & v_21928;
assign v_21930 = v_21929;
assign v_21932 = v_21099;
assign v_21933 = v_868;
assign v_21934 = v_21933;
assign v_21935 = v_21932 & v_21934;
assign v_21936 = v_21935;
assign v_21937 = v_21827 & v_21936;
assign v_21939 = v_21837 & v_21938;
assign v_21940 = v_21826 & v_21936;
assign v_21942 = v_21824 & v_21941;
assign v_21944 = v_21843 & v_21943;
assign v_21945 = v_21823 & v_21941;
assign v_21947 = v_21821 & v_21946;
assign v_21949 = v_21849 & v_21948;
assign v_21950 = v_21820 & v_21946;
assign v_21952 = v_21818 & v_21951;
assign v_21954 = v_21855 & v_21953;
assign v_21955 = v_21817 & v_21951;
assign v_21957 = v_21815 & v_21956;
assign v_21959 = v_21861 & v_21958;
assign v_21960 = v_21814 & v_21956;
assign v_21962 = v_21812 & v_21961;
assign v_21964 = v_21867 & v_21963;
assign v_21965 = v_21811 & v_21961;
assign v_21967 = v_21809 & v_21966;
assign v_21969 = v_21873 & v_21968;
assign v_21970 = v_21808 & v_21966;
assign v_21972 = v_21806 & v_21971;
assign v_21974 = v_21879 & v_21973;
assign v_21975 = v_21805 & v_21971;
assign v_21977 = v_21803 & v_21976;
assign v_21979 = v_21885 & v_21978;
assign v_21980 = v_21802 & v_21976;
assign v_21982 = v_21800 & v_21981;
assign v_21984 = v_21891 & v_21983;
assign v_21985 = v_21799 & v_21981;
assign v_21987 = v_21797 & v_21986;
assign v_21989 = v_21897 & v_21988;
assign v_21990 = v_21796 & v_21986;
assign v_21992 = v_21794 & v_21991;
assign v_21994 = v_21903 & v_21993;
assign v_21995 = v_21793 & v_21991;
assign v_21997 = v_21791 & v_21996;
assign v_21999 = v_21909 & v_21998;
assign v_22000 = v_21790 & v_21996;
assign v_22002 = v_21788 & v_22001;
assign v_22004 = v_21915 & v_22003;
assign v_22005 = v_21787 & v_22001;
assign v_22007 = v_21785 & v_22006;
assign v_22009 = v_21921 & v_22008;
assign v_22010 = v_21784 & v_22006;
assign v_22012 = v_21782 & v_22011;
assign v_22014 = v_21927 & v_22013;
assign v_22015 = v_21781 & v_22011;
assign v_22017 = v_22016;
assign v_22019 = v_21931 & v_22018;
assign v_22020 = v_22019;
assign v_22022 = v_22021;
assign v_22024 = ~v_1063;
assign v_22025 = ~v_21036;
assign v_22026 = v_21036;
assign v_22027 = ~v_1067;
assign v_22028 = ~v_21040;
assign v_22029 = v_21040;
assign v_22030 = ~v_1071;
assign v_22031 = ~v_21044;
assign v_22032 = v_21044;
assign v_22033 = ~v_1075;
assign v_22034 = ~v_21048;
assign v_22035 = v_21048;
assign v_22036 = ~v_21051;
assign v_22037 = ~v_1080;
assign v_22038 = v_1080;
assign v_22039 = ~v_21055;
assign v_22040 = ~v_1084;
assign v_22041 = v_1084;
assign v_22042 = ~v_21059;
assign v_22043 = ~v_1088;
assign v_22044 = v_1088;
assign v_22045 = ~v_21063;
assign v_22046 = ~v_1092;
assign v_22047 = v_1092;
assign v_22048 = ~v_21067;
assign v_22049 = ~v_1096;
assign v_22050 = v_1096;
assign v_22051 = ~v_21071;
assign v_22052 = ~v_1100;
assign v_22053 = v_1100;
assign v_22054 = ~v_21075;
assign v_22055 = ~v_1104;
assign v_22056 = v_1104;
assign v_22057 = ~v_21079;
assign v_22058 = ~v_1108;
assign v_22059 = v_1108;
assign v_22060 = ~v_21083;
assign v_22061 = ~v_1112;
assign v_22062 = v_1112;
assign v_22063 = ~v_21087;
assign v_22064 = ~v_1116;
assign v_22065 = v_1116;
assign v_22066 = ~v_21091;
assign v_22067 = ~v_1120;
assign v_22068 = v_1120;
assign v_22069 = ~v_21095;
assign v_22070 = ~v_1124;
assign v_22071 = v_1124;
assign v_22072 = ~v_21099;
assign v_22073 = ~v_1128;
assign v_22074 = v_22073;
assign v_22076 = v_22075;
assign v_22078 = v_22070 & v_22077;
assign v_22080 = v_21095;
assign v_22082 = v_22079 & v_22081;
assign v_22084 = v_22067 & v_22083;
assign v_22086 = v_21091;
assign v_22088 = v_22085 & v_22087;
assign v_22090 = v_22064 & v_22089;
assign v_22092 = v_21087;
assign v_22094 = v_22091 & v_22093;
assign v_22096 = v_22061 & v_22095;
assign v_22098 = v_21083;
assign v_22100 = v_22097 & v_22099;
assign v_22102 = v_22058 & v_22101;
assign v_22104 = v_21079;
assign v_22106 = v_22103 & v_22105;
assign v_22108 = v_22055 & v_22107;
assign v_22110 = v_21075;
assign v_22112 = v_22109 & v_22111;
assign v_22114 = v_22052 & v_22113;
assign v_22116 = v_21071;
assign v_22118 = v_22115 & v_22117;
assign v_22120 = v_22049 & v_22119;
assign v_22122 = v_21067;
assign v_22124 = v_22121 & v_22123;
assign v_22126 = v_22046 & v_22125;
assign v_22128 = v_21063;
assign v_22130 = v_22127 & v_22129;
assign v_22132 = v_22043 & v_22131;
assign v_22134 = v_21059;
assign v_22136 = v_22133 & v_22135;
assign v_22138 = v_22040 & v_22137;
assign v_22140 = v_21055;
assign v_22142 = v_22139 & v_22141;
assign v_22144 = v_22037 & v_22143;
assign v_22146 = v_21051;
assign v_22148 = v_22145 & v_22147;
assign v_22150 = v_22034 & v_22149;
assign v_22152 = v_1075;
assign v_22154 = v_22151 & v_22153;
assign v_22156 = v_22031 & v_22155;
assign v_22158 = v_1071;
assign v_22160 = v_22157 & v_22159;
assign v_22162 = v_22028 & v_22161;
assign v_22164 = v_1067;
assign v_22166 = v_22163 & v_22165;
assign v_22168 = v_22025 & v_22167;
assign v_22170 = v_1063;
assign v_22172 = v_22169 & v_22171;
assign v_22173 = v_22172;
assign v_22175 = v_21099;
assign v_22176 = v_1128;
assign v_22177 = v_22176;
assign v_22178 = v_22175 & v_22177;
assign v_22179 = v_22178;
assign v_22180 = v_22070 & v_22179;
assign v_22182 = v_22080 & v_22181;
assign v_22183 = v_22069 & v_22179;
assign v_22185 = v_22067 & v_22184;
assign v_22187 = v_22086 & v_22186;
assign v_22188 = v_22066 & v_22184;
assign v_22190 = v_22064 & v_22189;
assign v_22192 = v_22092 & v_22191;
assign v_22193 = v_22063 & v_22189;
assign v_22195 = v_22061 & v_22194;
assign v_22197 = v_22098 & v_22196;
assign v_22198 = v_22060 & v_22194;
assign v_22200 = v_22058 & v_22199;
assign v_22202 = v_22104 & v_22201;
assign v_22203 = v_22057 & v_22199;
assign v_22205 = v_22055 & v_22204;
assign v_22207 = v_22110 & v_22206;
assign v_22208 = v_22054 & v_22204;
assign v_22210 = v_22052 & v_22209;
assign v_22212 = v_22116 & v_22211;
assign v_22213 = v_22051 & v_22209;
assign v_22215 = v_22049 & v_22214;
assign v_22217 = v_22122 & v_22216;
assign v_22218 = v_22048 & v_22214;
assign v_22220 = v_22046 & v_22219;
assign v_22222 = v_22128 & v_22221;
assign v_22223 = v_22045 & v_22219;
assign v_22225 = v_22043 & v_22224;
assign v_22227 = v_22134 & v_22226;
assign v_22228 = v_22042 & v_22224;
assign v_22230 = v_22040 & v_22229;
assign v_22232 = v_22140 & v_22231;
assign v_22233 = v_22039 & v_22229;
assign v_22235 = v_22037 & v_22234;
assign v_22237 = v_22146 & v_22236;
assign v_22238 = v_22036 & v_22234;
assign v_22240 = v_22034 & v_22239;
assign v_22242 = v_22152 & v_22241;
assign v_22243 = v_22033 & v_22239;
assign v_22245 = v_22031 & v_22244;
assign v_22247 = v_22158 & v_22246;
assign v_22248 = v_22030 & v_22244;
assign v_22250 = v_22028 & v_22249;
assign v_22252 = v_22164 & v_22251;
assign v_22253 = v_22027 & v_22249;
assign v_22255 = v_22025 & v_22254;
assign v_22257 = v_22170 & v_22256;
assign v_22258 = v_22024 & v_22254;
assign v_22260 = v_22259;
assign v_22262 = v_22174 & v_22261;
assign v_22263 = v_22262;
assign v_22265 = v_22264;
assign v_22267 = ~v_1323;
assign v_22268 = ~v_21036;
assign v_22269 = v_21036;
assign v_22270 = ~v_1327;
assign v_22271 = ~v_21040;
assign v_22272 = v_21040;
assign v_22273 = ~v_1331;
assign v_22274 = ~v_21044;
assign v_22275 = v_21044;
assign v_22276 = ~v_1335;
assign v_22277 = ~v_21048;
assign v_22278 = v_21048;
assign v_22279 = ~v_21051;
assign v_22280 = ~v_1340;
assign v_22281 = v_1340;
assign v_22282 = ~v_21055;
assign v_22283 = ~v_1344;
assign v_22284 = v_1344;
assign v_22285 = ~v_21059;
assign v_22286 = ~v_1348;
assign v_22287 = v_1348;
assign v_22288 = ~v_21063;
assign v_22289 = ~v_1352;
assign v_22290 = v_1352;
assign v_22291 = ~v_21067;
assign v_22292 = ~v_1356;
assign v_22293 = v_1356;
assign v_22294 = ~v_21071;
assign v_22295 = ~v_1360;
assign v_22296 = v_1360;
assign v_22297 = ~v_21075;
assign v_22298 = ~v_1364;
assign v_22299 = v_1364;
assign v_22300 = ~v_21079;
assign v_22301 = ~v_1368;
assign v_22302 = v_1368;
assign v_22303 = ~v_21083;
assign v_22304 = ~v_1372;
assign v_22305 = v_1372;
assign v_22306 = ~v_21087;
assign v_22307 = ~v_1376;
assign v_22308 = v_1376;
assign v_22309 = ~v_21091;
assign v_22310 = ~v_1380;
assign v_22311 = v_1380;
assign v_22312 = ~v_21095;
assign v_22313 = ~v_1384;
assign v_22314 = v_1384;
assign v_22315 = ~v_21099;
assign v_22316 = ~v_1388;
assign v_22317 = v_22316;
assign v_22319 = v_22318;
assign v_22321 = v_22313 & v_22320;
assign v_22323 = v_21095;
assign v_22325 = v_22322 & v_22324;
assign v_22327 = v_22310 & v_22326;
assign v_22329 = v_21091;
assign v_22331 = v_22328 & v_22330;
assign v_22333 = v_22307 & v_22332;
assign v_22335 = v_21087;
assign v_22337 = v_22334 & v_22336;
assign v_22339 = v_22304 & v_22338;
assign v_22341 = v_21083;
assign v_22343 = v_22340 & v_22342;
assign v_22345 = v_22301 & v_22344;
assign v_22347 = v_21079;
assign v_22349 = v_22346 & v_22348;
assign v_22351 = v_22298 & v_22350;
assign v_22353 = v_21075;
assign v_22355 = v_22352 & v_22354;
assign v_22357 = v_22295 & v_22356;
assign v_22359 = v_21071;
assign v_22361 = v_22358 & v_22360;
assign v_22363 = v_22292 & v_22362;
assign v_22365 = v_21067;
assign v_22367 = v_22364 & v_22366;
assign v_22369 = v_22289 & v_22368;
assign v_22371 = v_21063;
assign v_22373 = v_22370 & v_22372;
assign v_22375 = v_22286 & v_22374;
assign v_22377 = v_21059;
assign v_22379 = v_22376 & v_22378;
assign v_22381 = v_22283 & v_22380;
assign v_22383 = v_21055;
assign v_22385 = v_22382 & v_22384;
assign v_22387 = v_22280 & v_22386;
assign v_22389 = v_21051;
assign v_22391 = v_22388 & v_22390;
assign v_22393 = v_22277 & v_22392;
assign v_22395 = v_1335;
assign v_22397 = v_22394 & v_22396;
assign v_22399 = v_22274 & v_22398;
assign v_22401 = v_1331;
assign v_22403 = v_22400 & v_22402;
assign v_22405 = v_22271 & v_22404;
assign v_22407 = v_1327;
assign v_22409 = v_22406 & v_22408;
assign v_22411 = v_22268 & v_22410;
assign v_22413 = v_1323;
assign v_22415 = v_22412 & v_22414;
assign v_22416 = v_22415;
assign v_22418 = v_21099;
assign v_22419 = v_1388;
assign v_22420 = v_22419;
assign v_22421 = v_22418 & v_22420;
assign v_22422 = v_22421;
assign v_22423 = v_22313 & v_22422;
assign v_22425 = v_22323 & v_22424;
assign v_22426 = v_22312 & v_22422;
assign v_22428 = v_22310 & v_22427;
assign v_22430 = v_22329 & v_22429;
assign v_22431 = v_22309 & v_22427;
assign v_22433 = v_22307 & v_22432;
assign v_22435 = v_22335 & v_22434;
assign v_22436 = v_22306 & v_22432;
assign v_22438 = v_22304 & v_22437;
assign v_22440 = v_22341 & v_22439;
assign v_22441 = v_22303 & v_22437;
assign v_22443 = v_22301 & v_22442;
assign v_22445 = v_22347 & v_22444;
assign v_22446 = v_22300 & v_22442;
assign v_22448 = v_22298 & v_22447;
assign v_22450 = v_22353 & v_22449;
assign v_22451 = v_22297 & v_22447;
assign v_22453 = v_22295 & v_22452;
assign v_22455 = v_22359 & v_22454;
assign v_22456 = v_22294 & v_22452;
assign v_22458 = v_22292 & v_22457;
assign v_22460 = v_22365 & v_22459;
assign v_22461 = v_22291 & v_22457;
assign v_22463 = v_22289 & v_22462;
assign v_22465 = v_22371 & v_22464;
assign v_22466 = v_22288 & v_22462;
assign v_22468 = v_22286 & v_22467;
assign v_22470 = v_22377 & v_22469;
assign v_22471 = v_22285 & v_22467;
assign v_22473 = v_22283 & v_22472;
assign v_22475 = v_22383 & v_22474;
assign v_22476 = v_22282 & v_22472;
assign v_22478 = v_22280 & v_22477;
assign v_22480 = v_22389 & v_22479;
assign v_22481 = v_22279 & v_22477;
assign v_22483 = v_22277 & v_22482;
assign v_22485 = v_22395 & v_22484;
assign v_22486 = v_22276 & v_22482;
assign v_22488 = v_22274 & v_22487;
assign v_22490 = v_22401 & v_22489;
assign v_22491 = v_22273 & v_22487;
assign v_22493 = v_22271 & v_22492;
assign v_22495 = v_22407 & v_22494;
assign v_22496 = v_22270 & v_22492;
assign v_22498 = v_22268 & v_22497;
assign v_22500 = v_22413 & v_22499;
assign v_22501 = v_22267 & v_22497;
assign v_22503 = v_22502;
assign v_22505 = v_22417 & v_22504;
assign v_22506 = v_22505;
assign v_22508 = v_22507;
assign v_22510 = ~v_1583;
assign v_22511 = ~v_21036;
assign v_22512 = v_21036;
assign v_22513 = ~v_1587;
assign v_22514 = ~v_21040;
assign v_22515 = v_21040;
assign v_22516 = ~v_1591;
assign v_22517 = ~v_21044;
assign v_22518 = v_21044;
assign v_22519 = ~v_1595;
assign v_22520 = ~v_21048;
assign v_22521 = v_21048;
assign v_22522 = ~v_21051;
assign v_22523 = ~v_1600;
assign v_22524 = v_1600;
assign v_22525 = ~v_21055;
assign v_22526 = ~v_1604;
assign v_22527 = v_1604;
assign v_22528 = ~v_21059;
assign v_22529 = ~v_1608;
assign v_22530 = v_1608;
assign v_22531 = ~v_21063;
assign v_22532 = ~v_1612;
assign v_22533 = v_1612;
assign v_22534 = ~v_21067;
assign v_22535 = ~v_1616;
assign v_22536 = v_1616;
assign v_22537 = ~v_21071;
assign v_22538 = ~v_1620;
assign v_22539 = v_1620;
assign v_22540 = ~v_21075;
assign v_22541 = ~v_1624;
assign v_22542 = v_1624;
assign v_22543 = ~v_21079;
assign v_22544 = ~v_1628;
assign v_22545 = v_1628;
assign v_22546 = ~v_21083;
assign v_22547 = ~v_1632;
assign v_22548 = v_1632;
assign v_22549 = ~v_21087;
assign v_22550 = ~v_1636;
assign v_22551 = v_1636;
assign v_22552 = ~v_21091;
assign v_22553 = ~v_1640;
assign v_22554 = v_1640;
assign v_22555 = ~v_21095;
assign v_22556 = ~v_1644;
assign v_22557 = v_1644;
assign v_22558 = ~v_21099;
assign v_22559 = ~v_1648;
assign v_22560 = v_22559;
assign v_22562 = v_22561;
assign v_22564 = v_22556 & v_22563;
assign v_22566 = v_21095;
assign v_22568 = v_22565 & v_22567;
assign v_22570 = v_22553 & v_22569;
assign v_22572 = v_21091;
assign v_22574 = v_22571 & v_22573;
assign v_22576 = v_22550 & v_22575;
assign v_22578 = v_21087;
assign v_22580 = v_22577 & v_22579;
assign v_22582 = v_22547 & v_22581;
assign v_22584 = v_21083;
assign v_22586 = v_22583 & v_22585;
assign v_22588 = v_22544 & v_22587;
assign v_22590 = v_21079;
assign v_22592 = v_22589 & v_22591;
assign v_22594 = v_22541 & v_22593;
assign v_22596 = v_21075;
assign v_22598 = v_22595 & v_22597;
assign v_22600 = v_22538 & v_22599;
assign v_22602 = v_21071;
assign v_22604 = v_22601 & v_22603;
assign v_22606 = v_22535 & v_22605;
assign v_22608 = v_21067;
assign v_22610 = v_22607 & v_22609;
assign v_22612 = v_22532 & v_22611;
assign v_22614 = v_21063;
assign v_22616 = v_22613 & v_22615;
assign v_22618 = v_22529 & v_22617;
assign v_22620 = v_21059;
assign v_22622 = v_22619 & v_22621;
assign v_22624 = v_22526 & v_22623;
assign v_22626 = v_21055;
assign v_22628 = v_22625 & v_22627;
assign v_22630 = v_22523 & v_22629;
assign v_22632 = v_21051;
assign v_22634 = v_22631 & v_22633;
assign v_22636 = v_22520 & v_22635;
assign v_22638 = v_1595;
assign v_22640 = v_22637 & v_22639;
assign v_22642 = v_22517 & v_22641;
assign v_22644 = v_1591;
assign v_22646 = v_22643 & v_22645;
assign v_22648 = v_22514 & v_22647;
assign v_22650 = v_1587;
assign v_22652 = v_22649 & v_22651;
assign v_22654 = v_22511 & v_22653;
assign v_22656 = v_1583;
assign v_22658 = v_22655 & v_22657;
assign v_22659 = v_22658;
assign v_22661 = v_21099;
assign v_22662 = v_1648;
assign v_22663 = v_22662;
assign v_22664 = v_22661 & v_22663;
assign v_22665 = v_22664;
assign v_22666 = v_22556 & v_22665;
assign v_22668 = v_22566 & v_22667;
assign v_22669 = v_22555 & v_22665;
assign v_22671 = v_22553 & v_22670;
assign v_22673 = v_22572 & v_22672;
assign v_22674 = v_22552 & v_22670;
assign v_22676 = v_22550 & v_22675;
assign v_22678 = v_22578 & v_22677;
assign v_22679 = v_22549 & v_22675;
assign v_22681 = v_22547 & v_22680;
assign v_22683 = v_22584 & v_22682;
assign v_22684 = v_22546 & v_22680;
assign v_22686 = v_22544 & v_22685;
assign v_22688 = v_22590 & v_22687;
assign v_22689 = v_22543 & v_22685;
assign v_22691 = v_22541 & v_22690;
assign v_22693 = v_22596 & v_22692;
assign v_22694 = v_22540 & v_22690;
assign v_22696 = v_22538 & v_22695;
assign v_22698 = v_22602 & v_22697;
assign v_22699 = v_22537 & v_22695;
assign v_22701 = v_22535 & v_22700;
assign v_22703 = v_22608 & v_22702;
assign v_22704 = v_22534 & v_22700;
assign v_22706 = v_22532 & v_22705;
assign v_22708 = v_22614 & v_22707;
assign v_22709 = v_22531 & v_22705;
assign v_22711 = v_22529 & v_22710;
assign v_22713 = v_22620 & v_22712;
assign v_22714 = v_22528 & v_22710;
assign v_22716 = v_22526 & v_22715;
assign v_22718 = v_22626 & v_22717;
assign v_22719 = v_22525 & v_22715;
assign v_22721 = v_22523 & v_22720;
assign v_22723 = v_22632 & v_22722;
assign v_22724 = v_22522 & v_22720;
assign v_22726 = v_22520 & v_22725;
assign v_22728 = v_22638 & v_22727;
assign v_22729 = v_22519 & v_22725;
assign v_22731 = v_22517 & v_22730;
assign v_22733 = v_22644 & v_22732;
assign v_22734 = v_22516 & v_22730;
assign v_22736 = v_22514 & v_22735;
assign v_22738 = v_22650 & v_22737;
assign v_22739 = v_22513 & v_22735;
assign v_22741 = v_22511 & v_22740;
assign v_22743 = v_22656 & v_22742;
assign v_22744 = v_22510 & v_22740;
assign v_22746 = v_22745;
assign v_22748 = v_22660 & v_22747;
assign v_22749 = v_22748;
assign v_22751 = v_22750;
assign v_22753 = ~v_1843;
assign v_22754 = ~v_21036;
assign v_22755 = v_21036;
assign v_22756 = ~v_1847;
assign v_22757 = ~v_21040;
assign v_22758 = v_21040;
assign v_22759 = ~v_1851;
assign v_22760 = ~v_21044;
assign v_22761 = v_21044;
assign v_22762 = ~v_1855;
assign v_22763 = ~v_21048;
assign v_22764 = v_21048;
assign v_22765 = ~v_21051;
assign v_22766 = ~v_1860;
assign v_22767 = v_1860;
assign v_22768 = ~v_21055;
assign v_22769 = ~v_1864;
assign v_22770 = v_1864;
assign v_22771 = ~v_21059;
assign v_22772 = ~v_1868;
assign v_22773 = v_1868;
assign v_22774 = ~v_21063;
assign v_22775 = ~v_1872;
assign v_22776 = v_1872;
assign v_22777 = ~v_21067;
assign v_22778 = ~v_1876;
assign v_22779 = v_1876;
assign v_22780 = ~v_21071;
assign v_22781 = ~v_1880;
assign v_22782 = v_1880;
assign v_22783 = ~v_21075;
assign v_22784 = ~v_1884;
assign v_22785 = v_1884;
assign v_22786 = ~v_21079;
assign v_22787 = ~v_1888;
assign v_22788 = v_1888;
assign v_22789 = ~v_21083;
assign v_22790 = ~v_1892;
assign v_22791 = v_1892;
assign v_22792 = ~v_21087;
assign v_22793 = ~v_1896;
assign v_22794 = v_1896;
assign v_22795 = ~v_21091;
assign v_22796 = ~v_1900;
assign v_22797 = v_1900;
assign v_22798 = ~v_21095;
assign v_22799 = ~v_1904;
assign v_22800 = v_1904;
assign v_22801 = ~v_21099;
assign v_22802 = ~v_1908;
assign v_22803 = v_22802;
assign v_22805 = v_22804;
assign v_22807 = v_22799 & v_22806;
assign v_22809 = v_21095;
assign v_22811 = v_22808 & v_22810;
assign v_22813 = v_22796 & v_22812;
assign v_22815 = v_21091;
assign v_22817 = v_22814 & v_22816;
assign v_22819 = v_22793 & v_22818;
assign v_22821 = v_21087;
assign v_22823 = v_22820 & v_22822;
assign v_22825 = v_22790 & v_22824;
assign v_22827 = v_21083;
assign v_22829 = v_22826 & v_22828;
assign v_22831 = v_22787 & v_22830;
assign v_22833 = v_21079;
assign v_22835 = v_22832 & v_22834;
assign v_22837 = v_22784 & v_22836;
assign v_22839 = v_21075;
assign v_22841 = v_22838 & v_22840;
assign v_22843 = v_22781 & v_22842;
assign v_22845 = v_21071;
assign v_22847 = v_22844 & v_22846;
assign v_22849 = v_22778 & v_22848;
assign v_22851 = v_21067;
assign v_22853 = v_22850 & v_22852;
assign v_22855 = v_22775 & v_22854;
assign v_22857 = v_21063;
assign v_22859 = v_22856 & v_22858;
assign v_22861 = v_22772 & v_22860;
assign v_22863 = v_21059;
assign v_22865 = v_22862 & v_22864;
assign v_22867 = v_22769 & v_22866;
assign v_22869 = v_21055;
assign v_22871 = v_22868 & v_22870;
assign v_22873 = v_22766 & v_22872;
assign v_22875 = v_21051;
assign v_22877 = v_22874 & v_22876;
assign v_22879 = v_22763 & v_22878;
assign v_22881 = v_1855;
assign v_22883 = v_22880 & v_22882;
assign v_22885 = v_22760 & v_22884;
assign v_22887 = v_1851;
assign v_22889 = v_22886 & v_22888;
assign v_22891 = v_22757 & v_22890;
assign v_22893 = v_1847;
assign v_22895 = v_22892 & v_22894;
assign v_22897 = v_22754 & v_22896;
assign v_22899 = v_1843;
assign v_22901 = v_22898 & v_22900;
assign v_22902 = v_22901;
assign v_22904 = v_21099;
assign v_22905 = v_1908;
assign v_22906 = v_22905;
assign v_22907 = v_22904 & v_22906;
assign v_22908 = v_22907;
assign v_22909 = v_22799 & v_22908;
assign v_22911 = v_22809 & v_22910;
assign v_22912 = v_22798 & v_22908;
assign v_22914 = v_22796 & v_22913;
assign v_22916 = v_22815 & v_22915;
assign v_22917 = v_22795 & v_22913;
assign v_22919 = v_22793 & v_22918;
assign v_22921 = v_22821 & v_22920;
assign v_22922 = v_22792 & v_22918;
assign v_22924 = v_22790 & v_22923;
assign v_22926 = v_22827 & v_22925;
assign v_22927 = v_22789 & v_22923;
assign v_22929 = v_22787 & v_22928;
assign v_22931 = v_22833 & v_22930;
assign v_22932 = v_22786 & v_22928;
assign v_22934 = v_22784 & v_22933;
assign v_22936 = v_22839 & v_22935;
assign v_22937 = v_22783 & v_22933;
assign v_22939 = v_22781 & v_22938;
assign v_22941 = v_22845 & v_22940;
assign v_22942 = v_22780 & v_22938;
assign v_22944 = v_22778 & v_22943;
assign v_22946 = v_22851 & v_22945;
assign v_22947 = v_22777 & v_22943;
assign v_22949 = v_22775 & v_22948;
assign v_22951 = v_22857 & v_22950;
assign v_22952 = v_22774 & v_22948;
assign v_22954 = v_22772 & v_22953;
assign v_22956 = v_22863 & v_22955;
assign v_22957 = v_22771 & v_22953;
assign v_22959 = v_22769 & v_22958;
assign v_22961 = v_22869 & v_22960;
assign v_22962 = v_22768 & v_22958;
assign v_22964 = v_22766 & v_22963;
assign v_22966 = v_22875 & v_22965;
assign v_22967 = v_22765 & v_22963;
assign v_22969 = v_22763 & v_22968;
assign v_22971 = v_22881 & v_22970;
assign v_22972 = v_22762 & v_22968;
assign v_22974 = v_22760 & v_22973;
assign v_22976 = v_22887 & v_22975;
assign v_22977 = v_22759 & v_22973;
assign v_22979 = v_22757 & v_22978;
assign v_22981 = v_22893 & v_22980;
assign v_22982 = v_22756 & v_22978;
assign v_22984 = v_22754 & v_22983;
assign v_22986 = v_22899 & v_22985;
assign v_22987 = v_22753 & v_22983;
assign v_22989 = v_22988;
assign v_22991 = v_22903 & v_22990;
assign v_22992 = v_22991;
assign v_22994 = v_22993;
assign v_22996 = ~v_2103;
assign v_22997 = ~v_21036;
assign v_22998 = v_21036;
assign v_22999 = ~v_2107;
assign v_23000 = ~v_21040;
assign v_23001 = v_21040;
assign v_23002 = ~v_2111;
assign v_23003 = ~v_21044;
assign v_23004 = v_21044;
assign v_23005 = ~v_2115;
assign v_23006 = ~v_21048;
assign v_23007 = v_21048;
assign v_23008 = ~v_21051;
assign v_23009 = ~v_2120;
assign v_23010 = v_2120;
assign v_23011 = ~v_21055;
assign v_23012 = ~v_2124;
assign v_23013 = v_2124;
assign v_23014 = ~v_21059;
assign v_23015 = ~v_2128;
assign v_23016 = v_2128;
assign v_23017 = ~v_21063;
assign v_23018 = ~v_2132;
assign v_23019 = v_2132;
assign v_23020 = ~v_21067;
assign v_23021 = ~v_2136;
assign v_23022 = v_2136;
assign v_23023 = ~v_21071;
assign v_23024 = ~v_2140;
assign v_23025 = v_2140;
assign v_23026 = ~v_21075;
assign v_23027 = ~v_2144;
assign v_23028 = v_2144;
assign v_23029 = ~v_21079;
assign v_23030 = ~v_2148;
assign v_23031 = v_2148;
assign v_23032 = ~v_21083;
assign v_23033 = ~v_2152;
assign v_23034 = v_2152;
assign v_23035 = ~v_21087;
assign v_23036 = ~v_2156;
assign v_23037 = v_2156;
assign v_23038 = ~v_21091;
assign v_23039 = ~v_2160;
assign v_23040 = v_2160;
assign v_23041 = ~v_21095;
assign v_23042 = ~v_2164;
assign v_23043 = v_2164;
assign v_23044 = ~v_21099;
assign v_23045 = ~v_2168;
assign v_23046 = v_23045;
assign v_23048 = v_23047;
assign v_23050 = v_23042 & v_23049;
assign v_23052 = v_21095;
assign v_23054 = v_23051 & v_23053;
assign v_23056 = v_23039 & v_23055;
assign v_23058 = v_21091;
assign v_23060 = v_23057 & v_23059;
assign v_23062 = v_23036 & v_23061;
assign v_23064 = v_21087;
assign v_23066 = v_23063 & v_23065;
assign v_23068 = v_23033 & v_23067;
assign v_23070 = v_21083;
assign v_23072 = v_23069 & v_23071;
assign v_23074 = v_23030 & v_23073;
assign v_23076 = v_21079;
assign v_23078 = v_23075 & v_23077;
assign v_23080 = v_23027 & v_23079;
assign v_23082 = v_21075;
assign v_23084 = v_23081 & v_23083;
assign v_23086 = v_23024 & v_23085;
assign v_23088 = v_21071;
assign v_23090 = v_23087 & v_23089;
assign v_23092 = v_23021 & v_23091;
assign v_23094 = v_21067;
assign v_23096 = v_23093 & v_23095;
assign v_23098 = v_23018 & v_23097;
assign v_23100 = v_21063;
assign v_23102 = v_23099 & v_23101;
assign v_23104 = v_23015 & v_23103;
assign v_23106 = v_21059;
assign v_23108 = v_23105 & v_23107;
assign v_23110 = v_23012 & v_23109;
assign v_23112 = v_21055;
assign v_23114 = v_23111 & v_23113;
assign v_23116 = v_23009 & v_23115;
assign v_23118 = v_21051;
assign v_23120 = v_23117 & v_23119;
assign v_23122 = v_23006 & v_23121;
assign v_23124 = v_2115;
assign v_23126 = v_23123 & v_23125;
assign v_23128 = v_23003 & v_23127;
assign v_23130 = v_2111;
assign v_23132 = v_23129 & v_23131;
assign v_23134 = v_23000 & v_23133;
assign v_23136 = v_2107;
assign v_23138 = v_23135 & v_23137;
assign v_23140 = v_22997 & v_23139;
assign v_23142 = v_2103;
assign v_23144 = v_23141 & v_23143;
assign v_23145 = v_23144;
assign v_23147 = v_21099;
assign v_23148 = v_2168;
assign v_23149 = v_23148;
assign v_23150 = v_23147 & v_23149;
assign v_23151 = v_23150;
assign v_23152 = v_23042 & v_23151;
assign v_23154 = v_23052 & v_23153;
assign v_23155 = v_23041 & v_23151;
assign v_23157 = v_23039 & v_23156;
assign v_23159 = v_23058 & v_23158;
assign v_23160 = v_23038 & v_23156;
assign v_23162 = v_23036 & v_23161;
assign v_23164 = v_23064 & v_23163;
assign v_23165 = v_23035 & v_23161;
assign v_23167 = v_23033 & v_23166;
assign v_23169 = v_23070 & v_23168;
assign v_23170 = v_23032 & v_23166;
assign v_23172 = v_23030 & v_23171;
assign v_23174 = v_23076 & v_23173;
assign v_23175 = v_23029 & v_23171;
assign v_23177 = v_23027 & v_23176;
assign v_23179 = v_23082 & v_23178;
assign v_23180 = v_23026 & v_23176;
assign v_23182 = v_23024 & v_23181;
assign v_23184 = v_23088 & v_23183;
assign v_23185 = v_23023 & v_23181;
assign v_23187 = v_23021 & v_23186;
assign v_23189 = v_23094 & v_23188;
assign v_23190 = v_23020 & v_23186;
assign v_23192 = v_23018 & v_23191;
assign v_23194 = v_23100 & v_23193;
assign v_23195 = v_23017 & v_23191;
assign v_23197 = v_23015 & v_23196;
assign v_23199 = v_23106 & v_23198;
assign v_23200 = v_23014 & v_23196;
assign v_23202 = v_23012 & v_23201;
assign v_23204 = v_23112 & v_23203;
assign v_23205 = v_23011 & v_23201;
assign v_23207 = v_23009 & v_23206;
assign v_23209 = v_23118 & v_23208;
assign v_23210 = v_23008 & v_23206;
assign v_23212 = v_23006 & v_23211;
assign v_23214 = v_23124 & v_23213;
assign v_23215 = v_23005 & v_23211;
assign v_23217 = v_23003 & v_23216;
assign v_23219 = v_23130 & v_23218;
assign v_23220 = v_23002 & v_23216;
assign v_23222 = v_23000 & v_23221;
assign v_23224 = v_23136 & v_23223;
assign v_23225 = v_22999 & v_23221;
assign v_23227 = v_22997 & v_23226;
assign v_23229 = v_23142 & v_23228;
assign v_23230 = v_22996 & v_23226;
assign v_23232 = v_23231;
assign v_23234 = v_23146 & v_23233;
assign v_23235 = v_23234;
assign v_23237 = v_23236;
assign v_23239 = ~v_2363;
assign v_23240 = ~v_21036;
assign v_23241 = v_21036;
assign v_23242 = ~v_2367;
assign v_23243 = ~v_21040;
assign v_23244 = v_21040;
assign v_23245 = ~v_2371;
assign v_23246 = ~v_21044;
assign v_23247 = v_21044;
assign v_23248 = ~v_2375;
assign v_23249 = ~v_21048;
assign v_23250 = v_21048;
assign v_23251 = ~v_21051;
assign v_23252 = ~v_2380;
assign v_23253 = v_2380;
assign v_23254 = ~v_21055;
assign v_23255 = ~v_2384;
assign v_23256 = v_2384;
assign v_23257 = ~v_21059;
assign v_23258 = ~v_2388;
assign v_23259 = v_2388;
assign v_23260 = ~v_21063;
assign v_23261 = ~v_2392;
assign v_23262 = v_2392;
assign v_23263 = ~v_21067;
assign v_23264 = ~v_2396;
assign v_23265 = v_2396;
assign v_23266 = ~v_21071;
assign v_23267 = ~v_2400;
assign v_23268 = v_2400;
assign v_23269 = ~v_21075;
assign v_23270 = ~v_2404;
assign v_23271 = v_2404;
assign v_23272 = ~v_21079;
assign v_23273 = ~v_2408;
assign v_23274 = v_2408;
assign v_23275 = ~v_21083;
assign v_23276 = ~v_2412;
assign v_23277 = v_2412;
assign v_23278 = ~v_21087;
assign v_23279 = ~v_2416;
assign v_23280 = v_2416;
assign v_23281 = ~v_21091;
assign v_23282 = ~v_2420;
assign v_23283 = v_2420;
assign v_23284 = ~v_21095;
assign v_23285 = ~v_2424;
assign v_23286 = v_2424;
assign v_23287 = ~v_21099;
assign v_23288 = ~v_2428;
assign v_23289 = v_23288;
assign v_23291 = v_23290;
assign v_23293 = v_23285 & v_23292;
assign v_23295 = v_21095;
assign v_23297 = v_23294 & v_23296;
assign v_23299 = v_23282 & v_23298;
assign v_23301 = v_21091;
assign v_23303 = v_23300 & v_23302;
assign v_23305 = v_23279 & v_23304;
assign v_23307 = v_21087;
assign v_23309 = v_23306 & v_23308;
assign v_23311 = v_23276 & v_23310;
assign v_23313 = v_21083;
assign v_23315 = v_23312 & v_23314;
assign v_23317 = v_23273 & v_23316;
assign v_23319 = v_21079;
assign v_23321 = v_23318 & v_23320;
assign v_23323 = v_23270 & v_23322;
assign v_23325 = v_21075;
assign v_23327 = v_23324 & v_23326;
assign v_23329 = v_23267 & v_23328;
assign v_23331 = v_21071;
assign v_23333 = v_23330 & v_23332;
assign v_23335 = v_23264 & v_23334;
assign v_23337 = v_21067;
assign v_23339 = v_23336 & v_23338;
assign v_23341 = v_23261 & v_23340;
assign v_23343 = v_21063;
assign v_23345 = v_23342 & v_23344;
assign v_23347 = v_23258 & v_23346;
assign v_23349 = v_21059;
assign v_23351 = v_23348 & v_23350;
assign v_23353 = v_23255 & v_23352;
assign v_23355 = v_21055;
assign v_23357 = v_23354 & v_23356;
assign v_23359 = v_23252 & v_23358;
assign v_23361 = v_21051;
assign v_23363 = v_23360 & v_23362;
assign v_23365 = v_23249 & v_23364;
assign v_23367 = v_2375;
assign v_23369 = v_23366 & v_23368;
assign v_23371 = v_23246 & v_23370;
assign v_23373 = v_2371;
assign v_23375 = v_23372 & v_23374;
assign v_23377 = v_23243 & v_23376;
assign v_23379 = v_2367;
assign v_23381 = v_23378 & v_23380;
assign v_23383 = v_23240 & v_23382;
assign v_23385 = v_2363;
assign v_23387 = v_23384 & v_23386;
assign v_23388 = v_23387;
assign v_23390 = v_21099;
assign v_23391 = v_2428;
assign v_23392 = v_23391;
assign v_23393 = v_23390 & v_23392;
assign v_23394 = v_23393;
assign v_23395 = v_23285 & v_23394;
assign v_23397 = v_23295 & v_23396;
assign v_23398 = v_23284 & v_23394;
assign v_23400 = v_23282 & v_23399;
assign v_23402 = v_23301 & v_23401;
assign v_23403 = v_23281 & v_23399;
assign v_23405 = v_23279 & v_23404;
assign v_23407 = v_23307 & v_23406;
assign v_23408 = v_23278 & v_23404;
assign v_23410 = v_23276 & v_23409;
assign v_23412 = v_23313 & v_23411;
assign v_23413 = v_23275 & v_23409;
assign v_23415 = v_23273 & v_23414;
assign v_23417 = v_23319 & v_23416;
assign v_23418 = v_23272 & v_23414;
assign v_23420 = v_23270 & v_23419;
assign v_23422 = v_23325 & v_23421;
assign v_23423 = v_23269 & v_23419;
assign v_23425 = v_23267 & v_23424;
assign v_23427 = v_23331 & v_23426;
assign v_23428 = v_23266 & v_23424;
assign v_23430 = v_23264 & v_23429;
assign v_23432 = v_23337 & v_23431;
assign v_23433 = v_23263 & v_23429;
assign v_23435 = v_23261 & v_23434;
assign v_23437 = v_23343 & v_23436;
assign v_23438 = v_23260 & v_23434;
assign v_23440 = v_23258 & v_23439;
assign v_23442 = v_23349 & v_23441;
assign v_23443 = v_23257 & v_23439;
assign v_23445 = v_23255 & v_23444;
assign v_23447 = v_23355 & v_23446;
assign v_23448 = v_23254 & v_23444;
assign v_23450 = v_23252 & v_23449;
assign v_23452 = v_23361 & v_23451;
assign v_23453 = v_23251 & v_23449;
assign v_23455 = v_23249 & v_23454;
assign v_23457 = v_23367 & v_23456;
assign v_23458 = v_23248 & v_23454;
assign v_23460 = v_23246 & v_23459;
assign v_23462 = v_23373 & v_23461;
assign v_23463 = v_23245 & v_23459;
assign v_23465 = v_23243 & v_23464;
assign v_23467 = v_23379 & v_23466;
assign v_23468 = v_23242 & v_23464;
assign v_23470 = v_23240 & v_23469;
assign v_23472 = v_23385 & v_23471;
assign v_23473 = v_23239 & v_23469;
assign v_23475 = v_23474;
assign v_23477 = v_23389 & v_23476;
assign v_23478 = v_23477;
assign v_23480 = v_23479;
assign v_23482 = ~v_2623;
assign v_23483 = ~v_21036;
assign v_23484 = v_21036;
assign v_23485 = ~v_2627;
assign v_23486 = ~v_21040;
assign v_23487 = v_21040;
assign v_23488 = ~v_2631;
assign v_23489 = ~v_21044;
assign v_23490 = v_21044;
assign v_23491 = ~v_2635;
assign v_23492 = ~v_21048;
assign v_23493 = v_21048;
assign v_23494 = ~v_21051;
assign v_23495 = ~v_2640;
assign v_23496 = v_2640;
assign v_23497 = ~v_21055;
assign v_23498 = ~v_2644;
assign v_23499 = v_2644;
assign v_23500 = ~v_21059;
assign v_23501 = ~v_2648;
assign v_23502 = v_2648;
assign v_23503 = ~v_21063;
assign v_23504 = ~v_2652;
assign v_23505 = v_2652;
assign v_23506 = ~v_21067;
assign v_23507 = ~v_2656;
assign v_23508 = v_2656;
assign v_23509 = ~v_21071;
assign v_23510 = ~v_2660;
assign v_23511 = v_2660;
assign v_23512 = ~v_21075;
assign v_23513 = ~v_2664;
assign v_23514 = v_2664;
assign v_23515 = ~v_21079;
assign v_23516 = ~v_2668;
assign v_23517 = v_2668;
assign v_23518 = ~v_21083;
assign v_23519 = ~v_2672;
assign v_23520 = v_2672;
assign v_23521 = ~v_21087;
assign v_23522 = ~v_2676;
assign v_23523 = v_2676;
assign v_23524 = ~v_21091;
assign v_23525 = ~v_2680;
assign v_23526 = v_2680;
assign v_23527 = ~v_21095;
assign v_23528 = ~v_2684;
assign v_23529 = v_2684;
assign v_23530 = ~v_21099;
assign v_23531 = ~v_2688;
assign v_23532 = v_23531;
assign v_23534 = v_23533;
assign v_23536 = v_23528 & v_23535;
assign v_23538 = v_21095;
assign v_23540 = v_23537 & v_23539;
assign v_23542 = v_23525 & v_23541;
assign v_23544 = v_21091;
assign v_23546 = v_23543 & v_23545;
assign v_23548 = v_23522 & v_23547;
assign v_23550 = v_21087;
assign v_23552 = v_23549 & v_23551;
assign v_23554 = v_23519 & v_23553;
assign v_23556 = v_21083;
assign v_23558 = v_23555 & v_23557;
assign v_23560 = v_23516 & v_23559;
assign v_23562 = v_21079;
assign v_23564 = v_23561 & v_23563;
assign v_23566 = v_23513 & v_23565;
assign v_23568 = v_21075;
assign v_23570 = v_23567 & v_23569;
assign v_23572 = v_23510 & v_23571;
assign v_23574 = v_21071;
assign v_23576 = v_23573 & v_23575;
assign v_23578 = v_23507 & v_23577;
assign v_23580 = v_21067;
assign v_23582 = v_23579 & v_23581;
assign v_23584 = v_23504 & v_23583;
assign v_23586 = v_21063;
assign v_23588 = v_23585 & v_23587;
assign v_23590 = v_23501 & v_23589;
assign v_23592 = v_21059;
assign v_23594 = v_23591 & v_23593;
assign v_23596 = v_23498 & v_23595;
assign v_23598 = v_21055;
assign v_23600 = v_23597 & v_23599;
assign v_23602 = v_23495 & v_23601;
assign v_23604 = v_21051;
assign v_23606 = v_23603 & v_23605;
assign v_23608 = v_23492 & v_23607;
assign v_23610 = v_2635;
assign v_23612 = v_23609 & v_23611;
assign v_23614 = v_23489 & v_23613;
assign v_23616 = v_2631;
assign v_23618 = v_23615 & v_23617;
assign v_23620 = v_23486 & v_23619;
assign v_23622 = v_2627;
assign v_23624 = v_23621 & v_23623;
assign v_23626 = v_23483 & v_23625;
assign v_23628 = v_2623;
assign v_23630 = v_23627 & v_23629;
assign v_23631 = v_23630;
assign v_23633 = v_21099;
assign v_23634 = v_2688;
assign v_23635 = v_23634;
assign v_23636 = v_23633 & v_23635;
assign v_23637 = v_23636;
assign v_23638 = v_23528 & v_23637;
assign v_23640 = v_23538 & v_23639;
assign v_23641 = v_23527 & v_23637;
assign v_23643 = v_23525 & v_23642;
assign v_23645 = v_23544 & v_23644;
assign v_23646 = v_23524 & v_23642;
assign v_23648 = v_23522 & v_23647;
assign v_23650 = v_23550 & v_23649;
assign v_23651 = v_23521 & v_23647;
assign v_23653 = v_23519 & v_23652;
assign v_23655 = v_23556 & v_23654;
assign v_23656 = v_23518 & v_23652;
assign v_23658 = v_23516 & v_23657;
assign v_23660 = v_23562 & v_23659;
assign v_23661 = v_23515 & v_23657;
assign v_23663 = v_23513 & v_23662;
assign v_23665 = v_23568 & v_23664;
assign v_23666 = v_23512 & v_23662;
assign v_23668 = v_23510 & v_23667;
assign v_23670 = v_23574 & v_23669;
assign v_23671 = v_23509 & v_23667;
assign v_23673 = v_23507 & v_23672;
assign v_23675 = v_23580 & v_23674;
assign v_23676 = v_23506 & v_23672;
assign v_23678 = v_23504 & v_23677;
assign v_23680 = v_23586 & v_23679;
assign v_23681 = v_23503 & v_23677;
assign v_23683 = v_23501 & v_23682;
assign v_23685 = v_23592 & v_23684;
assign v_23686 = v_23500 & v_23682;
assign v_23688 = v_23498 & v_23687;
assign v_23690 = v_23598 & v_23689;
assign v_23691 = v_23497 & v_23687;
assign v_23693 = v_23495 & v_23692;
assign v_23695 = v_23604 & v_23694;
assign v_23696 = v_23494 & v_23692;
assign v_23698 = v_23492 & v_23697;
assign v_23700 = v_23610 & v_23699;
assign v_23701 = v_23491 & v_23697;
assign v_23703 = v_23489 & v_23702;
assign v_23705 = v_23616 & v_23704;
assign v_23706 = v_23488 & v_23702;
assign v_23708 = v_23486 & v_23707;
assign v_23710 = v_23622 & v_23709;
assign v_23711 = v_23485 & v_23707;
assign v_23713 = v_23483 & v_23712;
assign v_23715 = v_23628 & v_23714;
assign v_23716 = v_23482 & v_23712;
assign v_23718 = v_23717;
assign v_23720 = v_23632 & v_23719;
assign v_23721 = v_23720;
assign v_23723 = v_23722;
assign v_23725 = ~v_2883;
assign v_23726 = ~v_21036;
assign v_23727 = v_21036;
assign v_23728 = ~v_2887;
assign v_23729 = ~v_21040;
assign v_23730 = v_21040;
assign v_23731 = ~v_2891;
assign v_23732 = ~v_21044;
assign v_23733 = v_21044;
assign v_23734 = ~v_2895;
assign v_23735 = ~v_21048;
assign v_23736 = v_21048;
assign v_23737 = ~v_21051;
assign v_23738 = ~v_2900;
assign v_23739 = v_2900;
assign v_23740 = ~v_21055;
assign v_23741 = ~v_2904;
assign v_23742 = v_2904;
assign v_23743 = ~v_21059;
assign v_23744 = ~v_2908;
assign v_23745 = v_2908;
assign v_23746 = ~v_21063;
assign v_23747 = ~v_2912;
assign v_23748 = v_2912;
assign v_23749 = ~v_21067;
assign v_23750 = ~v_2916;
assign v_23751 = v_2916;
assign v_23752 = ~v_21071;
assign v_23753 = ~v_2920;
assign v_23754 = v_2920;
assign v_23755 = ~v_21075;
assign v_23756 = ~v_2924;
assign v_23757 = v_2924;
assign v_23758 = ~v_21079;
assign v_23759 = ~v_2928;
assign v_23760 = v_2928;
assign v_23761 = ~v_21083;
assign v_23762 = ~v_2932;
assign v_23763 = v_2932;
assign v_23764 = ~v_21087;
assign v_23765 = ~v_2936;
assign v_23766 = v_2936;
assign v_23767 = ~v_21091;
assign v_23768 = ~v_2940;
assign v_23769 = v_2940;
assign v_23770 = ~v_21095;
assign v_23771 = ~v_2944;
assign v_23772 = v_2944;
assign v_23773 = ~v_21099;
assign v_23774 = ~v_2948;
assign v_23775 = v_23774;
assign v_23777 = v_23776;
assign v_23779 = v_23771 & v_23778;
assign v_23781 = v_21095;
assign v_23783 = v_23780 & v_23782;
assign v_23785 = v_23768 & v_23784;
assign v_23787 = v_21091;
assign v_23789 = v_23786 & v_23788;
assign v_23791 = v_23765 & v_23790;
assign v_23793 = v_21087;
assign v_23795 = v_23792 & v_23794;
assign v_23797 = v_23762 & v_23796;
assign v_23799 = v_21083;
assign v_23801 = v_23798 & v_23800;
assign v_23803 = v_23759 & v_23802;
assign v_23805 = v_21079;
assign v_23807 = v_23804 & v_23806;
assign v_23809 = v_23756 & v_23808;
assign v_23811 = v_21075;
assign v_23813 = v_23810 & v_23812;
assign v_23815 = v_23753 & v_23814;
assign v_23817 = v_21071;
assign v_23819 = v_23816 & v_23818;
assign v_23821 = v_23750 & v_23820;
assign v_23823 = v_21067;
assign v_23825 = v_23822 & v_23824;
assign v_23827 = v_23747 & v_23826;
assign v_23829 = v_21063;
assign v_23831 = v_23828 & v_23830;
assign v_23833 = v_23744 & v_23832;
assign v_23835 = v_21059;
assign v_23837 = v_23834 & v_23836;
assign v_23839 = v_23741 & v_23838;
assign v_23841 = v_21055;
assign v_23843 = v_23840 & v_23842;
assign v_23845 = v_23738 & v_23844;
assign v_23847 = v_21051;
assign v_23849 = v_23846 & v_23848;
assign v_23851 = v_23735 & v_23850;
assign v_23853 = v_2895;
assign v_23855 = v_23852 & v_23854;
assign v_23857 = v_23732 & v_23856;
assign v_23859 = v_2891;
assign v_23861 = v_23858 & v_23860;
assign v_23863 = v_23729 & v_23862;
assign v_23865 = v_2887;
assign v_23867 = v_23864 & v_23866;
assign v_23869 = v_23726 & v_23868;
assign v_23871 = v_2883;
assign v_23873 = v_23870 & v_23872;
assign v_23874 = v_23873;
assign v_23876 = v_21099;
assign v_23877 = v_2948;
assign v_23878 = v_23877;
assign v_23879 = v_23876 & v_23878;
assign v_23880 = v_23879;
assign v_23881 = v_23771 & v_23880;
assign v_23883 = v_23781 & v_23882;
assign v_23884 = v_23770 & v_23880;
assign v_23886 = v_23768 & v_23885;
assign v_23888 = v_23787 & v_23887;
assign v_23889 = v_23767 & v_23885;
assign v_23891 = v_23765 & v_23890;
assign v_23893 = v_23793 & v_23892;
assign v_23894 = v_23764 & v_23890;
assign v_23896 = v_23762 & v_23895;
assign v_23898 = v_23799 & v_23897;
assign v_23899 = v_23761 & v_23895;
assign v_23901 = v_23759 & v_23900;
assign v_23903 = v_23805 & v_23902;
assign v_23904 = v_23758 & v_23900;
assign v_23906 = v_23756 & v_23905;
assign v_23908 = v_23811 & v_23907;
assign v_23909 = v_23755 & v_23905;
assign v_23911 = v_23753 & v_23910;
assign v_23913 = v_23817 & v_23912;
assign v_23914 = v_23752 & v_23910;
assign v_23916 = v_23750 & v_23915;
assign v_23918 = v_23823 & v_23917;
assign v_23919 = v_23749 & v_23915;
assign v_23921 = v_23747 & v_23920;
assign v_23923 = v_23829 & v_23922;
assign v_23924 = v_23746 & v_23920;
assign v_23926 = v_23744 & v_23925;
assign v_23928 = v_23835 & v_23927;
assign v_23929 = v_23743 & v_23925;
assign v_23931 = v_23741 & v_23930;
assign v_23933 = v_23841 & v_23932;
assign v_23934 = v_23740 & v_23930;
assign v_23936 = v_23738 & v_23935;
assign v_23938 = v_23847 & v_23937;
assign v_23939 = v_23737 & v_23935;
assign v_23941 = v_23735 & v_23940;
assign v_23943 = v_23853 & v_23942;
assign v_23944 = v_23734 & v_23940;
assign v_23946 = v_23732 & v_23945;
assign v_23948 = v_23859 & v_23947;
assign v_23949 = v_23731 & v_23945;
assign v_23951 = v_23729 & v_23950;
assign v_23953 = v_23865 & v_23952;
assign v_23954 = v_23728 & v_23950;
assign v_23956 = v_23726 & v_23955;
assign v_23958 = v_23871 & v_23957;
assign v_23959 = v_23725 & v_23955;
assign v_23961 = v_23960;
assign v_23963 = v_23875 & v_23962;
assign v_23964 = v_23963;
assign v_23966 = v_23965;
assign v_23968 = ~v_3143;
assign v_23969 = ~v_21036;
assign v_23970 = v_21036;
assign v_23971 = ~v_3147;
assign v_23972 = ~v_21040;
assign v_23973 = v_21040;
assign v_23974 = ~v_3151;
assign v_23975 = ~v_21044;
assign v_23976 = v_21044;
assign v_23977 = ~v_3155;
assign v_23978 = ~v_21048;
assign v_23979 = v_21048;
assign v_23980 = ~v_21051;
assign v_23981 = ~v_3160;
assign v_23982 = v_3160;
assign v_23983 = ~v_21055;
assign v_23984 = ~v_3164;
assign v_23985 = v_3164;
assign v_23986 = ~v_21059;
assign v_23987 = ~v_3168;
assign v_23988 = v_3168;
assign v_23989 = ~v_21063;
assign v_23990 = ~v_3172;
assign v_23991 = v_3172;
assign v_23992 = ~v_21067;
assign v_23993 = ~v_3176;
assign v_23994 = v_3176;
assign v_23995 = ~v_21071;
assign v_23996 = ~v_3180;
assign v_23997 = v_3180;
assign v_23998 = ~v_21075;
assign v_23999 = ~v_3184;
assign v_24000 = v_3184;
assign v_24001 = ~v_21079;
assign v_24002 = ~v_3188;
assign v_24003 = v_3188;
assign v_24004 = ~v_21083;
assign v_24005 = ~v_3192;
assign v_24006 = v_3192;
assign v_24007 = ~v_21087;
assign v_24008 = ~v_3196;
assign v_24009 = v_3196;
assign v_24010 = ~v_21091;
assign v_24011 = ~v_3200;
assign v_24012 = v_3200;
assign v_24013 = ~v_21095;
assign v_24014 = ~v_3204;
assign v_24015 = v_3204;
assign v_24016 = ~v_21099;
assign v_24017 = ~v_3208;
assign v_24018 = v_24017;
assign v_24020 = v_24019;
assign v_24022 = v_24014 & v_24021;
assign v_24024 = v_21095;
assign v_24026 = v_24023 & v_24025;
assign v_24028 = v_24011 & v_24027;
assign v_24030 = v_21091;
assign v_24032 = v_24029 & v_24031;
assign v_24034 = v_24008 & v_24033;
assign v_24036 = v_21087;
assign v_24038 = v_24035 & v_24037;
assign v_24040 = v_24005 & v_24039;
assign v_24042 = v_21083;
assign v_24044 = v_24041 & v_24043;
assign v_24046 = v_24002 & v_24045;
assign v_24048 = v_21079;
assign v_24050 = v_24047 & v_24049;
assign v_24052 = v_23999 & v_24051;
assign v_24054 = v_21075;
assign v_24056 = v_24053 & v_24055;
assign v_24058 = v_23996 & v_24057;
assign v_24060 = v_21071;
assign v_24062 = v_24059 & v_24061;
assign v_24064 = v_23993 & v_24063;
assign v_24066 = v_21067;
assign v_24068 = v_24065 & v_24067;
assign v_24070 = v_23990 & v_24069;
assign v_24072 = v_21063;
assign v_24074 = v_24071 & v_24073;
assign v_24076 = v_23987 & v_24075;
assign v_24078 = v_21059;
assign v_24080 = v_24077 & v_24079;
assign v_24082 = v_23984 & v_24081;
assign v_24084 = v_21055;
assign v_24086 = v_24083 & v_24085;
assign v_24088 = v_23981 & v_24087;
assign v_24090 = v_21051;
assign v_24092 = v_24089 & v_24091;
assign v_24094 = v_23978 & v_24093;
assign v_24096 = v_3155;
assign v_24098 = v_24095 & v_24097;
assign v_24100 = v_23975 & v_24099;
assign v_24102 = v_3151;
assign v_24104 = v_24101 & v_24103;
assign v_24106 = v_23972 & v_24105;
assign v_24108 = v_3147;
assign v_24110 = v_24107 & v_24109;
assign v_24112 = v_23969 & v_24111;
assign v_24114 = v_3143;
assign v_24116 = v_24113 & v_24115;
assign v_24117 = v_24116;
assign v_24119 = v_21099;
assign v_24120 = v_3208;
assign v_24121 = v_24120;
assign v_24122 = v_24119 & v_24121;
assign v_24123 = v_24122;
assign v_24124 = v_24014 & v_24123;
assign v_24126 = v_24024 & v_24125;
assign v_24127 = v_24013 & v_24123;
assign v_24129 = v_24011 & v_24128;
assign v_24131 = v_24030 & v_24130;
assign v_24132 = v_24010 & v_24128;
assign v_24134 = v_24008 & v_24133;
assign v_24136 = v_24036 & v_24135;
assign v_24137 = v_24007 & v_24133;
assign v_24139 = v_24005 & v_24138;
assign v_24141 = v_24042 & v_24140;
assign v_24142 = v_24004 & v_24138;
assign v_24144 = v_24002 & v_24143;
assign v_24146 = v_24048 & v_24145;
assign v_24147 = v_24001 & v_24143;
assign v_24149 = v_23999 & v_24148;
assign v_24151 = v_24054 & v_24150;
assign v_24152 = v_23998 & v_24148;
assign v_24154 = v_23996 & v_24153;
assign v_24156 = v_24060 & v_24155;
assign v_24157 = v_23995 & v_24153;
assign v_24159 = v_23993 & v_24158;
assign v_24161 = v_24066 & v_24160;
assign v_24162 = v_23992 & v_24158;
assign v_24164 = v_23990 & v_24163;
assign v_24166 = v_24072 & v_24165;
assign v_24167 = v_23989 & v_24163;
assign v_24169 = v_23987 & v_24168;
assign v_24171 = v_24078 & v_24170;
assign v_24172 = v_23986 & v_24168;
assign v_24174 = v_23984 & v_24173;
assign v_24176 = v_24084 & v_24175;
assign v_24177 = v_23983 & v_24173;
assign v_24179 = v_23981 & v_24178;
assign v_24181 = v_24090 & v_24180;
assign v_24182 = v_23980 & v_24178;
assign v_24184 = v_23978 & v_24183;
assign v_24186 = v_24096 & v_24185;
assign v_24187 = v_23977 & v_24183;
assign v_24189 = v_23975 & v_24188;
assign v_24191 = v_24102 & v_24190;
assign v_24192 = v_23974 & v_24188;
assign v_24194 = v_23972 & v_24193;
assign v_24196 = v_24108 & v_24195;
assign v_24197 = v_23971 & v_24193;
assign v_24199 = v_23969 & v_24198;
assign v_24201 = v_24114 & v_24200;
assign v_24202 = v_23968 & v_24198;
assign v_24204 = v_24203;
assign v_24206 = v_24118 & v_24205;
assign v_24207 = v_24206;
assign v_24209 = v_24208;
assign v_24211 = ~v_3403;
assign v_24212 = ~v_21036;
assign v_24213 = v_21036;
assign v_24214 = ~v_3407;
assign v_24215 = ~v_21040;
assign v_24216 = v_21040;
assign v_24217 = ~v_3411;
assign v_24218 = ~v_21044;
assign v_24219 = v_21044;
assign v_24220 = ~v_3415;
assign v_24221 = ~v_21048;
assign v_24222 = v_21048;
assign v_24223 = ~v_21051;
assign v_24224 = ~v_3420;
assign v_24225 = v_3420;
assign v_24226 = ~v_21055;
assign v_24227 = ~v_3424;
assign v_24228 = v_3424;
assign v_24229 = ~v_21059;
assign v_24230 = ~v_3428;
assign v_24231 = v_3428;
assign v_24232 = ~v_21063;
assign v_24233 = ~v_3432;
assign v_24234 = v_3432;
assign v_24235 = ~v_21067;
assign v_24236 = ~v_3436;
assign v_24237 = v_3436;
assign v_24238 = ~v_21071;
assign v_24239 = ~v_3440;
assign v_24240 = v_3440;
assign v_24241 = ~v_21075;
assign v_24242 = ~v_3444;
assign v_24243 = v_3444;
assign v_24244 = ~v_21079;
assign v_24245 = ~v_3448;
assign v_24246 = v_3448;
assign v_24247 = ~v_21083;
assign v_24248 = ~v_3452;
assign v_24249 = v_3452;
assign v_24250 = ~v_21087;
assign v_24251 = ~v_3456;
assign v_24252 = v_3456;
assign v_24253 = ~v_21091;
assign v_24254 = ~v_3460;
assign v_24255 = v_3460;
assign v_24256 = ~v_21095;
assign v_24257 = ~v_3464;
assign v_24258 = v_3464;
assign v_24259 = ~v_21099;
assign v_24260 = ~v_3468;
assign v_24261 = v_24260;
assign v_24263 = v_24262;
assign v_24265 = v_24257 & v_24264;
assign v_24267 = v_21095;
assign v_24269 = v_24266 & v_24268;
assign v_24271 = v_24254 & v_24270;
assign v_24273 = v_21091;
assign v_24275 = v_24272 & v_24274;
assign v_24277 = v_24251 & v_24276;
assign v_24279 = v_21087;
assign v_24281 = v_24278 & v_24280;
assign v_24283 = v_24248 & v_24282;
assign v_24285 = v_21083;
assign v_24287 = v_24284 & v_24286;
assign v_24289 = v_24245 & v_24288;
assign v_24291 = v_21079;
assign v_24293 = v_24290 & v_24292;
assign v_24295 = v_24242 & v_24294;
assign v_24297 = v_21075;
assign v_24299 = v_24296 & v_24298;
assign v_24301 = v_24239 & v_24300;
assign v_24303 = v_21071;
assign v_24305 = v_24302 & v_24304;
assign v_24307 = v_24236 & v_24306;
assign v_24309 = v_21067;
assign v_24311 = v_24308 & v_24310;
assign v_24313 = v_24233 & v_24312;
assign v_24315 = v_21063;
assign v_24317 = v_24314 & v_24316;
assign v_24319 = v_24230 & v_24318;
assign v_24321 = v_21059;
assign v_24323 = v_24320 & v_24322;
assign v_24325 = v_24227 & v_24324;
assign v_24327 = v_21055;
assign v_24329 = v_24326 & v_24328;
assign v_24331 = v_24224 & v_24330;
assign v_24333 = v_21051;
assign v_24335 = v_24332 & v_24334;
assign v_24337 = v_24221 & v_24336;
assign v_24339 = v_3415;
assign v_24341 = v_24338 & v_24340;
assign v_24343 = v_24218 & v_24342;
assign v_24345 = v_3411;
assign v_24347 = v_24344 & v_24346;
assign v_24349 = v_24215 & v_24348;
assign v_24351 = v_3407;
assign v_24353 = v_24350 & v_24352;
assign v_24355 = v_24212 & v_24354;
assign v_24357 = v_3403;
assign v_24359 = v_24356 & v_24358;
assign v_24360 = v_24359;
assign v_24362 = v_21099;
assign v_24363 = v_3468;
assign v_24364 = v_24363;
assign v_24365 = v_24362 & v_24364;
assign v_24366 = v_24365;
assign v_24367 = v_24257 & v_24366;
assign v_24369 = v_24267 & v_24368;
assign v_24370 = v_24256 & v_24366;
assign v_24372 = v_24254 & v_24371;
assign v_24374 = v_24273 & v_24373;
assign v_24375 = v_24253 & v_24371;
assign v_24377 = v_24251 & v_24376;
assign v_24379 = v_24279 & v_24378;
assign v_24380 = v_24250 & v_24376;
assign v_24382 = v_24248 & v_24381;
assign v_24384 = v_24285 & v_24383;
assign v_24385 = v_24247 & v_24381;
assign v_24387 = v_24245 & v_24386;
assign v_24389 = v_24291 & v_24388;
assign v_24390 = v_24244 & v_24386;
assign v_24392 = v_24242 & v_24391;
assign v_24394 = v_24297 & v_24393;
assign v_24395 = v_24241 & v_24391;
assign v_24397 = v_24239 & v_24396;
assign v_24399 = v_24303 & v_24398;
assign v_24400 = v_24238 & v_24396;
assign v_24402 = v_24236 & v_24401;
assign v_24404 = v_24309 & v_24403;
assign v_24405 = v_24235 & v_24401;
assign v_24407 = v_24233 & v_24406;
assign v_24409 = v_24315 & v_24408;
assign v_24410 = v_24232 & v_24406;
assign v_24412 = v_24230 & v_24411;
assign v_24414 = v_24321 & v_24413;
assign v_24415 = v_24229 & v_24411;
assign v_24417 = v_24227 & v_24416;
assign v_24419 = v_24327 & v_24418;
assign v_24420 = v_24226 & v_24416;
assign v_24422 = v_24224 & v_24421;
assign v_24424 = v_24333 & v_24423;
assign v_24425 = v_24223 & v_24421;
assign v_24427 = v_24221 & v_24426;
assign v_24429 = v_24339 & v_24428;
assign v_24430 = v_24220 & v_24426;
assign v_24432 = v_24218 & v_24431;
assign v_24434 = v_24345 & v_24433;
assign v_24435 = v_24217 & v_24431;
assign v_24437 = v_24215 & v_24436;
assign v_24439 = v_24351 & v_24438;
assign v_24440 = v_24214 & v_24436;
assign v_24442 = v_24212 & v_24441;
assign v_24444 = v_24357 & v_24443;
assign v_24445 = v_24211 & v_24441;
assign v_24447 = v_24446;
assign v_24449 = v_24361 & v_24448;
assign v_24450 = v_24449;
assign v_24452 = v_24451;
assign v_24454 = ~v_3663;
assign v_24455 = ~v_21036;
assign v_24456 = v_21036;
assign v_24457 = ~v_3667;
assign v_24458 = ~v_21040;
assign v_24459 = v_21040;
assign v_24460 = ~v_3671;
assign v_24461 = ~v_21044;
assign v_24462 = v_21044;
assign v_24463 = ~v_3675;
assign v_24464 = ~v_21048;
assign v_24465 = v_21048;
assign v_24466 = ~v_21051;
assign v_24467 = ~v_3680;
assign v_24468 = v_3680;
assign v_24469 = ~v_21055;
assign v_24470 = ~v_3684;
assign v_24471 = v_3684;
assign v_24472 = ~v_21059;
assign v_24473 = ~v_3688;
assign v_24474 = v_3688;
assign v_24475 = ~v_21063;
assign v_24476 = ~v_3692;
assign v_24477 = v_3692;
assign v_24478 = ~v_21067;
assign v_24479 = ~v_3696;
assign v_24480 = v_3696;
assign v_24481 = ~v_21071;
assign v_24482 = ~v_3700;
assign v_24483 = v_3700;
assign v_24484 = ~v_21075;
assign v_24485 = ~v_3704;
assign v_24486 = v_3704;
assign v_24487 = ~v_21079;
assign v_24488 = ~v_3708;
assign v_24489 = v_3708;
assign v_24490 = ~v_21083;
assign v_24491 = ~v_3712;
assign v_24492 = v_3712;
assign v_24493 = ~v_21087;
assign v_24494 = ~v_3716;
assign v_24495 = v_3716;
assign v_24496 = ~v_21091;
assign v_24497 = ~v_3720;
assign v_24498 = v_3720;
assign v_24499 = ~v_21095;
assign v_24500 = ~v_3724;
assign v_24501 = v_3724;
assign v_24502 = ~v_21099;
assign v_24503 = ~v_3728;
assign v_24504 = v_24503;
assign v_24506 = v_24505;
assign v_24508 = v_24500 & v_24507;
assign v_24510 = v_21095;
assign v_24512 = v_24509 & v_24511;
assign v_24514 = v_24497 & v_24513;
assign v_24516 = v_21091;
assign v_24518 = v_24515 & v_24517;
assign v_24520 = v_24494 & v_24519;
assign v_24522 = v_21087;
assign v_24524 = v_24521 & v_24523;
assign v_24526 = v_24491 & v_24525;
assign v_24528 = v_21083;
assign v_24530 = v_24527 & v_24529;
assign v_24532 = v_24488 & v_24531;
assign v_24534 = v_21079;
assign v_24536 = v_24533 & v_24535;
assign v_24538 = v_24485 & v_24537;
assign v_24540 = v_21075;
assign v_24542 = v_24539 & v_24541;
assign v_24544 = v_24482 & v_24543;
assign v_24546 = v_21071;
assign v_24548 = v_24545 & v_24547;
assign v_24550 = v_24479 & v_24549;
assign v_24552 = v_21067;
assign v_24554 = v_24551 & v_24553;
assign v_24556 = v_24476 & v_24555;
assign v_24558 = v_21063;
assign v_24560 = v_24557 & v_24559;
assign v_24562 = v_24473 & v_24561;
assign v_24564 = v_21059;
assign v_24566 = v_24563 & v_24565;
assign v_24568 = v_24470 & v_24567;
assign v_24570 = v_21055;
assign v_24572 = v_24569 & v_24571;
assign v_24574 = v_24467 & v_24573;
assign v_24576 = v_21051;
assign v_24578 = v_24575 & v_24577;
assign v_24580 = v_24464 & v_24579;
assign v_24582 = v_3675;
assign v_24584 = v_24581 & v_24583;
assign v_24586 = v_24461 & v_24585;
assign v_24588 = v_3671;
assign v_24590 = v_24587 & v_24589;
assign v_24592 = v_24458 & v_24591;
assign v_24594 = v_3667;
assign v_24596 = v_24593 & v_24595;
assign v_24598 = v_24455 & v_24597;
assign v_24600 = v_3663;
assign v_24602 = v_24599 & v_24601;
assign v_24603 = v_24602;
assign v_24605 = v_21099;
assign v_24606 = v_3728;
assign v_24607 = v_24606;
assign v_24608 = v_24605 & v_24607;
assign v_24609 = v_24608;
assign v_24610 = v_24500 & v_24609;
assign v_24612 = v_24510 & v_24611;
assign v_24613 = v_24499 & v_24609;
assign v_24615 = v_24497 & v_24614;
assign v_24617 = v_24516 & v_24616;
assign v_24618 = v_24496 & v_24614;
assign v_24620 = v_24494 & v_24619;
assign v_24622 = v_24522 & v_24621;
assign v_24623 = v_24493 & v_24619;
assign v_24625 = v_24491 & v_24624;
assign v_24627 = v_24528 & v_24626;
assign v_24628 = v_24490 & v_24624;
assign v_24630 = v_24488 & v_24629;
assign v_24632 = v_24534 & v_24631;
assign v_24633 = v_24487 & v_24629;
assign v_24635 = v_24485 & v_24634;
assign v_24637 = v_24540 & v_24636;
assign v_24638 = v_24484 & v_24634;
assign v_24640 = v_24482 & v_24639;
assign v_24642 = v_24546 & v_24641;
assign v_24643 = v_24481 & v_24639;
assign v_24645 = v_24479 & v_24644;
assign v_24647 = v_24552 & v_24646;
assign v_24648 = v_24478 & v_24644;
assign v_24650 = v_24476 & v_24649;
assign v_24652 = v_24558 & v_24651;
assign v_24653 = v_24475 & v_24649;
assign v_24655 = v_24473 & v_24654;
assign v_24657 = v_24564 & v_24656;
assign v_24658 = v_24472 & v_24654;
assign v_24660 = v_24470 & v_24659;
assign v_24662 = v_24570 & v_24661;
assign v_24663 = v_24469 & v_24659;
assign v_24665 = v_24467 & v_24664;
assign v_24667 = v_24576 & v_24666;
assign v_24668 = v_24466 & v_24664;
assign v_24670 = v_24464 & v_24669;
assign v_24672 = v_24582 & v_24671;
assign v_24673 = v_24463 & v_24669;
assign v_24675 = v_24461 & v_24674;
assign v_24677 = v_24588 & v_24676;
assign v_24678 = v_24460 & v_24674;
assign v_24680 = v_24458 & v_24679;
assign v_24682 = v_24594 & v_24681;
assign v_24683 = v_24457 & v_24679;
assign v_24685 = v_24455 & v_24684;
assign v_24687 = v_24600 & v_24686;
assign v_24688 = v_24454 & v_24684;
assign v_24690 = v_24689;
assign v_24692 = v_24604 & v_24691;
assign v_24693 = v_24692;
assign v_24695 = v_24694;
assign v_24697 = ~v_3923;
assign v_24698 = ~v_21036;
assign v_24699 = v_21036;
assign v_24700 = ~v_3927;
assign v_24701 = ~v_21040;
assign v_24702 = v_21040;
assign v_24703 = ~v_3931;
assign v_24704 = ~v_21044;
assign v_24705 = v_21044;
assign v_24706 = ~v_3935;
assign v_24707 = ~v_21048;
assign v_24708 = v_21048;
assign v_24709 = ~v_21051;
assign v_24710 = ~v_3940;
assign v_24711 = v_3940;
assign v_24712 = ~v_21055;
assign v_24713 = ~v_3944;
assign v_24714 = v_3944;
assign v_24715 = ~v_21059;
assign v_24716 = ~v_3948;
assign v_24717 = v_3948;
assign v_24718 = ~v_21063;
assign v_24719 = ~v_3952;
assign v_24720 = v_3952;
assign v_24721 = ~v_21067;
assign v_24722 = ~v_3956;
assign v_24723 = v_3956;
assign v_24724 = ~v_21071;
assign v_24725 = ~v_3960;
assign v_24726 = v_3960;
assign v_24727 = ~v_21075;
assign v_24728 = ~v_3964;
assign v_24729 = v_3964;
assign v_24730 = ~v_21079;
assign v_24731 = ~v_3968;
assign v_24732 = v_3968;
assign v_24733 = ~v_21083;
assign v_24734 = ~v_3972;
assign v_24735 = v_3972;
assign v_24736 = ~v_21087;
assign v_24737 = ~v_3976;
assign v_24738 = v_3976;
assign v_24739 = ~v_21091;
assign v_24740 = ~v_3980;
assign v_24741 = v_3980;
assign v_24742 = ~v_21095;
assign v_24743 = ~v_3984;
assign v_24744 = v_3984;
assign v_24745 = ~v_21099;
assign v_24746 = ~v_3988;
assign v_24747 = v_24746;
assign v_24749 = v_24748;
assign v_24751 = v_24743 & v_24750;
assign v_24753 = v_21095;
assign v_24755 = v_24752 & v_24754;
assign v_24757 = v_24740 & v_24756;
assign v_24759 = v_21091;
assign v_24761 = v_24758 & v_24760;
assign v_24763 = v_24737 & v_24762;
assign v_24765 = v_21087;
assign v_24767 = v_24764 & v_24766;
assign v_24769 = v_24734 & v_24768;
assign v_24771 = v_21083;
assign v_24773 = v_24770 & v_24772;
assign v_24775 = v_24731 & v_24774;
assign v_24777 = v_21079;
assign v_24779 = v_24776 & v_24778;
assign v_24781 = v_24728 & v_24780;
assign v_24783 = v_21075;
assign v_24785 = v_24782 & v_24784;
assign v_24787 = v_24725 & v_24786;
assign v_24789 = v_21071;
assign v_24791 = v_24788 & v_24790;
assign v_24793 = v_24722 & v_24792;
assign v_24795 = v_21067;
assign v_24797 = v_24794 & v_24796;
assign v_24799 = v_24719 & v_24798;
assign v_24801 = v_21063;
assign v_24803 = v_24800 & v_24802;
assign v_24805 = v_24716 & v_24804;
assign v_24807 = v_21059;
assign v_24809 = v_24806 & v_24808;
assign v_24811 = v_24713 & v_24810;
assign v_24813 = v_21055;
assign v_24815 = v_24812 & v_24814;
assign v_24817 = v_24710 & v_24816;
assign v_24819 = v_21051;
assign v_24821 = v_24818 & v_24820;
assign v_24823 = v_24707 & v_24822;
assign v_24825 = v_3935;
assign v_24827 = v_24824 & v_24826;
assign v_24829 = v_24704 & v_24828;
assign v_24831 = v_3931;
assign v_24833 = v_24830 & v_24832;
assign v_24835 = v_24701 & v_24834;
assign v_24837 = v_3927;
assign v_24839 = v_24836 & v_24838;
assign v_24841 = v_24698 & v_24840;
assign v_24843 = v_3923;
assign v_24845 = v_24842 & v_24844;
assign v_24846 = v_24845;
assign v_24848 = v_21099;
assign v_24849 = v_3988;
assign v_24850 = v_24849;
assign v_24851 = v_24848 & v_24850;
assign v_24852 = v_24851;
assign v_24853 = v_24743 & v_24852;
assign v_24855 = v_24753 & v_24854;
assign v_24856 = v_24742 & v_24852;
assign v_24858 = v_24740 & v_24857;
assign v_24860 = v_24759 & v_24859;
assign v_24861 = v_24739 & v_24857;
assign v_24863 = v_24737 & v_24862;
assign v_24865 = v_24765 & v_24864;
assign v_24866 = v_24736 & v_24862;
assign v_24868 = v_24734 & v_24867;
assign v_24870 = v_24771 & v_24869;
assign v_24871 = v_24733 & v_24867;
assign v_24873 = v_24731 & v_24872;
assign v_24875 = v_24777 & v_24874;
assign v_24876 = v_24730 & v_24872;
assign v_24878 = v_24728 & v_24877;
assign v_24880 = v_24783 & v_24879;
assign v_24881 = v_24727 & v_24877;
assign v_24883 = v_24725 & v_24882;
assign v_24885 = v_24789 & v_24884;
assign v_24886 = v_24724 & v_24882;
assign v_24888 = v_24722 & v_24887;
assign v_24890 = v_24795 & v_24889;
assign v_24891 = v_24721 & v_24887;
assign v_24893 = v_24719 & v_24892;
assign v_24895 = v_24801 & v_24894;
assign v_24896 = v_24718 & v_24892;
assign v_24898 = v_24716 & v_24897;
assign v_24900 = v_24807 & v_24899;
assign v_24901 = v_24715 & v_24897;
assign v_24903 = v_24713 & v_24902;
assign v_24905 = v_24813 & v_24904;
assign v_24906 = v_24712 & v_24902;
assign v_24908 = v_24710 & v_24907;
assign v_24910 = v_24819 & v_24909;
assign v_24911 = v_24709 & v_24907;
assign v_24913 = v_24707 & v_24912;
assign v_24915 = v_24825 & v_24914;
assign v_24916 = v_24706 & v_24912;
assign v_24918 = v_24704 & v_24917;
assign v_24920 = v_24831 & v_24919;
assign v_24921 = v_24703 & v_24917;
assign v_24923 = v_24701 & v_24922;
assign v_24925 = v_24837 & v_24924;
assign v_24926 = v_24700 & v_24922;
assign v_24928 = v_24698 & v_24927;
assign v_24930 = v_24843 & v_24929;
assign v_24931 = v_24697 & v_24927;
assign v_24933 = v_24932;
assign v_24935 = v_24847 & v_24934;
assign v_24936 = v_24935;
assign v_24938 = v_24937;
assign v_24939 = ~v_4182;
assign v_24940 = ~v_21036;
assign v_24941 = v_21036;
assign v_24942 = ~v_4186;
assign v_24943 = ~v_21040;
assign v_24944 = v_21040;
assign v_24945 = ~v_4190;
assign v_24946 = ~v_21044;
assign v_24947 = v_21044;
assign v_24948 = ~v_4194;
assign v_24949 = ~v_21048;
assign v_24950 = v_21048;
assign v_24951 = ~v_21051;
assign v_24952 = ~v_4199;
assign v_24953 = v_4199;
assign v_24954 = ~v_21055;
assign v_24955 = ~v_4203;
assign v_24956 = v_4203;
assign v_24957 = ~v_21059;
assign v_24958 = ~v_4207;
assign v_24959 = v_4207;
assign v_24960 = ~v_21063;
assign v_24961 = ~v_4211;
assign v_24962 = v_4211;
assign v_24963 = ~v_21067;
assign v_24964 = ~v_4215;
assign v_24965 = v_4215;
assign v_24966 = ~v_21071;
assign v_24967 = ~v_4219;
assign v_24968 = v_4219;
assign v_24969 = ~v_21075;
assign v_24970 = ~v_4223;
assign v_24971 = v_4223;
assign v_24972 = ~v_21079;
assign v_24973 = ~v_4227;
assign v_24974 = v_4227;
assign v_24975 = ~v_21083;
assign v_24976 = ~v_4231;
assign v_24977 = v_4231;
assign v_24978 = ~v_21087;
assign v_24979 = ~v_4235;
assign v_24980 = v_4235;
assign v_24981 = ~v_21091;
assign v_24982 = ~v_4239;
assign v_24983 = v_4239;
assign v_24984 = ~v_21095;
assign v_24985 = ~v_4243;
assign v_24986 = v_4243;
assign v_24987 = ~v_21099;
assign v_24988 = ~v_4247;
assign v_24989 = v_24988;
assign v_24991 = v_24990;
assign v_24993 = v_24985 & v_24992;
assign v_24995 = v_21095;
assign v_24997 = v_24994 & v_24996;
assign v_24999 = v_24982 & v_24998;
assign v_25001 = v_21091;
assign v_25003 = v_25000 & v_25002;
assign v_25005 = v_24979 & v_25004;
assign v_25007 = v_21087;
assign v_25009 = v_25006 & v_25008;
assign v_25011 = v_24976 & v_25010;
assign v_25013 = v_21083;
assign v_25015 = v_25012 & v_25014;
assign v_25017 = v_24973 & v_25016;
assign v_25019 = v_21079;
assign v_25021 = v_25018 & v_25020;
assign v_25023 = v_24970 & v_25022;
assign v_25025 = v_21075;
assign v_25027 = v_25024 & v_25026;
assign v_25029 = v_24967 & v_25028;
assign v_25031 = v_21071;
assign v_25033 = v_25030 & v_25032;
assign v_25035 = v_24964 & v_25034;
assign v_25037 = v_21067;
assign v_25039 = v_25036 & v_25038;
assign v_25041 = v_24961 & v_25040;
assign v_25043 = v_21063;
assign v_25045 = v_25042 & v_25044;
assign v_25047 = v_24958 & v_25046;
assign v_25049 = v_21059;
assign v_25051 = v_25048 & v_25050;
assign v_25053 = v_24955 & v_25052;
assign v_25055 = v_21055;
assign v_25057 = v_25054 & v_25056;
assign v_25059 = v_24952 & v_25058;
assign v_25061 = v_21051;
assign v_25063 = v_25060 & v_25062;
assign v_25065 = v_24949 & v_25064;
assign v_25067 = v_4194;
assign v_25069 = v_25066 & v_25068;
assign v_25071 = v_24946 & v_25070;
assign v_25073 = v_4190;
assign v_25075 = v_25072 & v_25074;
assign v_25077 = v_24943 & v_25076;
assign v_25079 = v_4186;
assign v_25081 = v_25078 & v_25080;
assign v_25083 = v_24940 & v_25082;
assign v_25085 = v_4182;
assign v_25087 = v_25084 & v_25086;
assign v_25089 = ~v_25088;
assign v_25091 = v_21099;
assign v_25092 = v_4247;
assign v_25093 = v_25092;
assign v_25094 = v_25091 & v_25093;
assign v_25095 = v_25094;
assign v_25096 = v_24985 & v_25095;
assign v_25098 = v_24995 & v_25097;
assign v_25099 = v_24984 & v_25095;
assign v_25101 = v_24982 & v_25100;
assign v_25103 = v_25001 & v_25102;
assign v_25104 = v_24981 & v_25100;
assign v_25106 = v_24979 & v_25105;
assign v_25108 = v_25007 & v_25107;
assign v_25109 = v_24978 & v_25105;
assign v_25111 = v_24976 & v_25110;
assign v_25113 = v_25013 & v_25112;
assign v_25114 = v_24975 & v_25110;
assign v_25116 = v_24973 & v_25115;
assign v_25118 = v_25019 & v_25117;
assign v_25119 = v_24972 & v_25115;
assign v_25121 = v_24970 & v_25120;
assign v_25123 = v_25025 & v_25122;
assign v_25124 = v_24969 & v_25120;
assign v_25126 = v_24967 & v_25125;
assign v_25128 = v_25031 & v_25127;
assign v_25129 = v_24966 & v_25125;
assign v_25131 = v_24964 & v_25130;
assign v_25133 = v_25037 & v_25132;
assign v_25134 = v_24963 & v_25130;
assign v_25136 = v_24961 & v_25135;
assign v_25138 = v_25043 & v_25137;
assign v_25139 = v_24960 & v_25135;
assign v_25141 = v_24958 & v_25140;
assign v_25143 = v_25049 & v_25142;
assign v_25144 = v_24957 & v_25140;
assign v_25146 = v_24955 & v_25145;
assign v_25148 = v_25055 & v_25147;
assign v_25149 = v_24954 & v_25145;
assign v_25151 = v_24952 & v_25150;
assign v_25153 = v_25061 & v_25152;
assign v_25154 = v_24951 & v_25150;
assign v_25156 = v_24949 & v_25155;
assign v_25158 = v_25067 & v_25157;
assign v_25159 = v_24948 & v_25155;
assign v_25161 = v_24946 & v_25160;
assign v_25163 = v_25073 & v_25162;
assign v_25164 = v_24945 & v_25160;
assign v_25166 = v_24943 & v_25165;
assign v_25168 = v_25079 & v_25167;
assign v_25169 = v_24942 & v_25165;
assign v_25171 = v_24940 & v_25170;
assign v_25173 = v_25085 & v_25172;
assign v_25174 = v_24939 & v_25170;
assign v_25176 = v_25088;
assign v_25178 = v_25090 & v_25177;
assign v_25179 = v_25178;
assign v_25181 = v_25180;
assign v_25183 = ~v_6;
assign v_25185 = ~v_25184;
assign v_25186 = v_25184;
assign v_25187 = ~v_13;
assign v_25189 = ~v_25188;
assign v_25190 = v_25188;
assign v_25191 = ~v_18;
assign v_25193 = ~v_25192;
assign v_25194 = v_25192;
assign v_25195 = ~v_23;
assign v_25197 = ~v_25196;
assign v_25198 = v_25196;
assign v_25200 = ~v_25199;
assign v_25201 = ~v_30;
assign v_25202 = v_30;
assign v_25204 = ~v_25203;
assign v_25205 = ~v_35;
assign v_25206 = v_35;
assign v_25208 = ~v_25207;
assign v_25209 = ~v_40;
assign v_25210 = v_40;
assign v_25212 = ~v_25211;
assign v_25213 = ~v_45;
assign v_25214 = v_45;
assign v_25216 = ~v_25215;
assign v_25217 = ~v_50;
assign v_25218 = v_50;
assign v_25220 = ~v_25219;
assign v_25221 = ~v_55;
assign v_25222 = v_55;
assign v_25224 = ~v_25223;
assign v_25225 = ~v_60;
assign v_25226 = v_60;
assign v_25228 = ~v_25227;
assign v_25229 = ~v_65;
assign v_25230 = v_65;
assign v_25232 = ~v_25231;
assign v_25233 = ~v_70;
assign v_25234 = v_70;
assign v_25236 = ~v_25235;
assign v_25237 = ~v_75;
assign v_25238 = v_75;
assign v_25240 = ~v_25239;
assign v_25241 = ~v_80;
assign v_25242 = v_80;
assign v_25244 = ~v_25243;
assign v_25245 = ~v_85;
assign v_25246 = v_85;
assign v_25248 = ~v_25247;
assign v_25249 = ~v_90;
assign v_25250 = v_25249;
assign v_25252 = v_25251;
assign v_25254 = v_25245 & v_25253;
assign v_25256 = v_25243;
assign v_25258 = v_25255 & v_25257;
assign v_25260 = v_25241 & v_25259;
assign v_25262 = v_25239;
assign v_25264 = v_25261 & v_25263;
assign v_25266 = v_25237 & v_25265;
assign v_25268 = v_25235;
assign v_25270 = v_25267 & v_25269;
assign v_25272 = v_25233 & v_25271;
assign v_25274 = v_25231;
assign v_25276 = v_25273 & v_25275;
assign v_25278 = v_25229 & v_25277;
assign v_25280 = v_25227;
assign v_25282 = v_25279 & v_25281;
assign v_25284 = v_25225 & v_25283;
assign v_25286 = v_25223;
assign v_25288 = v_25285 & v_25287;
assign v_25290 = v_25221 & v_25289;
assign v_25292 = v_25219;
assign v_25294 = v_25291 & v_25293;
assign v_25296 = v_25217 & v_25295;
assign v_25298 = v_25215;
assign v_25300 = v_25297 & v_25299;
assign v_25302 = v_25213 & v_25301;
assign v_25304 = v_25211;
assign v_25306 = v_25303 & v_25305;
assign v_25308 = v_25209 & v_25307;
assign v_25310 = v_25207;
assign v_25312 = v_25309 & v_25311;
assign v_25314 = v_25205 & v_25313;
assign v_25316 = v_25203;
assign v_25318 = v_25315 & v_25317;
assign v_25320 = v_25201 & v_25319;
assign v_25322 = v_25199;
assign v_25324 = v_25321 & v_25323;
assign v_25326 = v_25197 & v_25325;
assign v_25328 = v_23;
assign v_25330 = v_25327 & v_25329;
assign v_25332 = v_25193 & v_25331;
assign v_25334 = v_18;
assign v_25336 = v_25333 & v_25335;
assign v_25338 = v_25189 & v_25337;
assign v_25340 = v_13;
assign v_25342 = v_25339 & v_25341;
assign v_25344 = v_25185 & v_25343;
assign v_25346 = v_6;
assign v_25348 = v_25345 & v_25347;
assign v_25349 = v_25348;
assign v_25351 = v_25247;
assign v_25352 = v_90;
assign v_25353 = v_25352;
assign v_25354 = v_25351 & v_25353;
assign v_25355 = v_25354;
assign v_25356 = v_25245 & v_25355;
assign v_25358 = v_25256 & v_25357;
assign v_25359 = v_25244 & v_25355;
assign v_25361 = v_25241 & v_25360;
assign v_25363 = v_25262 & v_25362;
assign v_25364 = v_25240 & v_25360;
assign v_25366 = v_25237 & v_25365;
assign v_25368 = v_25268 & v_25367;
assign v_25369 = v_25236 & v_25365;
assign v_25371 = v_25233 & v_25370;
assign v_25373 = v_25274 & v_25372;
assign v_25374 = v_25232 & v_25370;
assign v_25376 = v_25229 & v_25375;
assign v_25378 = v_25280 & v_25377;
assign v_25379 = v_25228 & v_25375;
assign v_25381 = v_25225 & v_25380;
assign v_25383 = v_25286 & v_25382;
assign v_25384 = v_25224 & v_25380;
assign v_25386 = v_25221 & v_25385;
assign v_25388 = v_25292 & v_25387;
assign v_25389 = v_25220 & v_25385;
assign v_25391 = v_25217 & v_25390;
assign v_25393 = v_25298 & v_25392;
assign v_25394 = v_25216 & v_25390;
assign v_25396 = v_25213 & v_25395;
assign v_25398 = v_25304 & v_25397;
assign v_25399 = v_25212 & v_25395;
assign v_25401 = v_25209 & v_25400;
assign v_25403 = v_25310 & v_25402;
assign v_25404 = v_25208 & v_25400;
assign v_25406 = v_25205 & v_25405;
assign v_25408 = v_25316 & v_25407;
assign v_25409 = v_25204 & v_25405;
assign v_25411 = v_25201 & v_25410;
assign v_25413 = v_25322 & v_25412;
assign v_25414 = v_25200 & v_25410;
assign v_25416 = v_25197 & v_25415;
assign v_25418 = v_25328 & v_25417;
assign v_25419 = v_25195 & v_25415;
assign v_25421 = v_25193 & v_25420;
assign v_25423 = v_25334 & v_25422;
assign v_25424 = v_25191 & v_25420;
assign v_25426 = v_25189 & v_25425;
assign v_25428 = v_25340 & v_25427;
assign v_25429 = v_25187 & v_25425;
assign v_25431 = v_25185 & v_25430;
assign v_25433 = v_25346 & v_25432;
assign v_25434 = v_25183 & v_25430;
assign v_25436 = v_25435;
assign v_25438 = v_25350 & v_25437;
assign v_25439 = v_25438;
assign v_25441 = v_25440;
assign v_25443 = ~v_283;
assign v_25444 = ~v_25184;
assign v_25445 = v_25184;
assign v_25446 = ~v_287;
assign v_25447 = ~v_25188;
assign v_25448 = v_25188;
assign v_25449 = ~v_291;
assign v_25450 = ~v_25192;
assign v_25451 = v_25192;
assign v_25452 = ~v_295;
assign v_25453 = ~v_25196;
assign v_25454 = v_25196;
assign v_25455 = ~v_25199;
assign v_25456 = ~v_300;
assign v_25457 = v_300;
assign v_25458 = ~v_25203;
assign v_25459 = ~v_304;
assign v_25460 = v_304;
assign v_25461 = ~v_25207;
assign v_25462 = ~v_308;
assign v_25463 = v_308;
assign v_25464 = ~v_25211;
assign v_25465 = ~v_312;
assign v_25466 = v_312;
assign v_25467 = ~v_25215;
assign v_25468 = ~v_316;
assign v_25469 = v_316;
assign v_25470 = ~v_25219;
assign v_25471 = ~v_320;
assign v_25472 = v_320;
assign v_25473 = ~v_25223;
assign v_25474 = ~v_324;
assign v_25475 = v_324;
assign v_25476 = ~v_25227;
assign v_25477 = ~v_328;
assign v_25478 = v_328;
assign v_25479 = ~v_25231;
assign v_25480 = ~v_332;
assign v_25481 = v_332;
assign v_25482 = ~v_25235;
assign v_25483 = ~v_336;
assign v_25484 = v_336;
assign v_25485 = ~v_25239;
assign v_25486 = ~v_340;
assign v_25487 = v_340;
assign v_25488 = ~v_25243;
assign v_25489 = ~v_344;
assign v_25490 = v_344;
assign v_25491 = ~v_25247;
assign v_25492 = ~v_348;
assign v_25493 = v_25492;
assign v_25495 = v_25494;
assign v_25497 = v_25489 & v_25496;
assign v_25499 = v_25243;
assign v_25501 = v_25498 & v_25500;
assign v_25503 = v_25486 & v_25502;
assign v_25505 = v_25239;
assign v_25507 = v_25504 & v_25506;
assign v_25509 = v_25483 & v_25508;
assign v_25511 = v_25235;
assign v_25513 = v_25510 & v_25512;
assign v_25515 = v_25480 & v_25514;
assign v_25517 = v_25231;
assign v_25519 = v_25516 & v_25518;
assign v_25521 = v_25477 & v_25520;
assign v_25523 = v_25227;
assign v_25525 = v_25522 & v_25524;
assign v_25527 = v_25474 & v_25526;
assign v_25529 = v_25223;
assign v_25531 = v_25528 & v_25530;
assign v_25533 = v_25471 & v_25532;
assign v_25535 = v_25219;
assign v_25537 = v_25534 & v_25536;
assign v_25539 = v_25468 & v_25538;
assign v_25541 = v_25215;
assign v_25543 = v_25540 & v_25542;
assign v_25545 = v_25465 & v_25544;
assign v_25547 = v_25211;
assign v_25549 = v_25546 & v_25548;
assign v_25551 = v_25462 & v_25550;
assign v_25553 = v_25207;
assign v_25555 = v_25552 & v_25554;
assign v_25557 = v_25459 & v_25556;
assign v_25559 = v_25203;
assign v_25561 = v_25558 & v_25560;
assign v_25563 = v_25456 & v_25562;
assign v_25565 = v_25199;
assign v_25567 = v_25564 & v_25566;
assign v_25569 = v_25453 & v_25568;
assign v_25571 = v_295;
assign v_25573 = v_25570 & v_25572;
assign v_25575 = v_25450 & v_25574;
assign v_25577 = v_291;
assign v_25579 = v_25576 & v_25578;
assign v_25581 = v_25447 & v_25580;
assign v_25583 = v_287;
assign v_25585 = v_25582 & v_25584;
assign v_25587 = v_25444 & v_25586;
assign v_25589 = v_283;
assign v_25591 = v_25588 & v_25590;
assign v_25592 = v_25591;
assign v_25594 = v_25247;
assign v_25595 = v_348;
assign v_25596 = v_25595;
assign v_25597 = v_25594 & v_25596;
assign v_25598 = v_25597;
assign v_25599 = v_25489 & v_25598;
assign v_25601 = v_25499 & v_25600;
assign v_25602 = v_25488 & v_25598;
assign v_25604 = v_25486 & v_25603;
assign v_25606 = v_25505 & v_25605;
assign v_25607 = v_25485 & v_25603;
assign v_25609 = v_25483 & v_25608;
assign v_25611 = v_25511 & v_25610;
assign v_25612 = v_25482 & v_25608;
assign v_25614 = v_25480 & v_25613;
assign v_25616 = v_25517 & v_25615;
assign v_25617 = v_25479 & v_25613;
assign v_25619 = v_25477 & v_25618;
assign v_25621 = v_25523 & v_25620;
assign v_25622 = v_25476 & v_25618;
assign v_25624 = v_25474 & v_25623;
assign v_25626 = v_25529 & v_25625;
assign v_25627 = v_25473 & v_25623;
assign v_25629 = v_25471 & v_25628;
assign v_25631 = v_25535 & v_25630;
assign v_25632 = v_25470 & v_25628;
assign v_25634 = v_25468 & v_25633;
assign v_25636 = v_25541 & v_25635;
assign v_25637 = v_25467 & v_25633;
assign v_25639 = v_25465 & v_25638;
assign v_25641 = v_25547 & v_25640;
assign v_25642 = v_25464 & v_25638;
assign v_25644 = v_25462 & v_25643;
assign v_25646 = v_25553 & v_25645;
assign v_25647 = v_25461 & v_25643;
assign v_25649 = v_25459 & v_25648;
assign v_25651 = v_25559 & v_25650;
assign v_25652 = v_25458 & v_25648;
assign v_25654 = v_25456 & v_25653;
assign v_25656 = v_25565 & v_25655;
assign v_25657 = v_25455 & v_25653;
assign v_25659 = v_25453 & v_25658;
assign v_25661 = v_25571 & v_25660;
assign v_25662 = v_25452 & v_25658;
assign v_25664 = v_25450 & v_25663;
assign v_25666 = v_25577 & v_25665;
assign v_25667 = v_25449 & v_25663;
assign v_25669 = v_25447 & v_25668;
assign v_25671 = v_25583 & v_25670;
assign v_25672 = v_25446 & v_25668;
assign v_25674 = v_25444 & v_25673;
assign v_25676 = v_25589 & v_25675;
assign v_25677 = v_25443 & v_25673;
assign v_25679 = v_25678;
assign v_25681 = v_25593 & v_25680;
assign v_25682 = v_25681;
assign v_25684 = v_25683;
assign v_25686 = ~v_543;
assign v_25687 = ~v_25184;
assign v_25688 = v_25184;
assign v_25689 = ~v_547;
assign v_25690 = ~v_25188;
assign v_25691 = v_25188;
assign v_25692 = ~v_551;
assign v_25693 = ~v_25192;
assign v_25694 = v_25192;
assign v_25695 = ~v_555;
assign v_25696 = ~v_25196;
assign v_25697 = v_25196;
assign v_25698 = ~v_25199;
assign v_25699 = ~v_560;
assign v_25700 = v_560;
assign v_25701 = ~v_25203;
assign v_25702 = ~v_564;
assign v_25703 = v_564;
assign v_25704 = ~v_25207;
assign v_25705 = ~v_568;
assign v_25706 = v_568;
assign v_25707 = ~v_25211;
assign v_25708 = ~v_572;
assign v_25709 = v_572;
assign v_25710 = ~v_25215;
assign v_25711 = ~v_576;
assign v_25712 = v_576;
assign v_25713 = ~v_25219;
assign v_25714 = ~v_580;
assign v_25715 = v_580;
assign v_25716 = ~v_25223;
assign v_25717 = ~v_584;
assign v_25718 = v_584;
assign v_25719 = ~v_25227;
assign v_25720 = ~v_588;
assign v_25721 = v_588;
assign v_25722 = ~v_25231;
assign v_25723 = ~v_592;
assign v_25724 = v_592;
assign v_25725 = ~v_25235;
assign v_25726 = ~v_596;
assign v_25727 = v_596;
assign v_25728 = ~v_25239;
assign v_25729 = ~v_600;
assign v_25730 = v_600;
assign v_25731 = ~v_25243;
assign v_25732 = ~v_604;
assign v_25733 = v_604;
assign v_25734 = ~v_25247;
assign v_25735 = ~v_608;
assign v_25736 = v_25735;
assign v_25738 = v_25737;
assign v_25740 = v_25732 & v_25739;
assign v_25742 = v_25243;
assign v_25744 = v_25741 & v_25743;
assign v_25746 = v_25729 & v_25745;
assign v_25748 = v_25239;
assign v_25750 = v_25747 & v_25749;
assign v_25752 = v_25726 & v_25751;
assign v_25754 = v_25235;
assign v_25756 = v_25753 & v_25755;
assign v_25758 = v_25723 & v_25757;
assign v_25760 = v_25231;
assign v_25762 = v_25759 & v_25761;
assign v_25764 = v_25720 & v_25763;
assign v_25766 = v_25227;
assign v_25768 = v_25765 & v_25767;
assign v_25770 = v_25717 & v_25769;
assign v_25772 = v_25223;
assign v_25774 = v_25771 & v_25773;
assign v_25776 = v_25714 & v_25775;
assign v_25778 = v_25219;
assign v_25780 = v_25777 & v_25779;
assign v_25782 = v_25711 & v_25781;
assign v_25784 = v_25215;
assign v_25786 = v_25783 & v_25785;
assign v_25788 = v_25708 & v_25787;
assign v_25790 = v_25211;
assign v_25792 = v_25789 & v_25791;
assign v_25794 = v_25705 & v_25793;
assign v_25796 = v_25207;
assign v_25798 = v_25795 & v_25797;
assign v_25800 = v_25702 & v_25799;
assign v_25802 = v_25203;
assign v_25804 = v_25801 & v_25803;
assign v_25806 = v_25699 & v_25805;
assign v_25808 = v_25199;
assign v_25810 = v_25807 & v_25809;
assign v_25812 = v_25696 & v_25811;
assign v_25814 = v_555;
assign v_25816 = v_25813 & v_25815;
assign v_25818 = v_25693 & v_25817;
assign v_25820 = v_551;
assign v_25822 = v_25819 & v_25821;
assign v_25824 = v_25690 & v_25823;
assign v_25826 = v_547;
assign v_25828 = v_25825 & v_25827;
assign v_25830 = v_25687 & v_25829;
assign v_25832 = v_543;
assign v_25834 = v_25831 & v_25833;
assign v_25835 = v_25834;
assign v_25837 = v_25247;
assign v_25838 = v_608;
assign v_25839 = v_25838;
assign v_25840 = v_25837 & v_25839;
assign v_25841 = v_25840;
assign v_25842 = v_25732 & v_25841;
assign v_25844 = v_25742 & v_25843;
assign v_25845 = v_25731 & v_25841;
assign v_25847 = v_25729 & v_25846;
assign v_25849 = v_25748 & v_25848;
assign v_25850 = v_25728 & v_25846;
assign v_25852 = v_25726 & v_25851;
assign v_25854 = v_25754 & v_25853;
assign v_25855 = v_25725 & v_25851;
assign v_25857 = v_25723 & v_25856;
assign v_25859 = v_25760 & v_25858;
assign v_25860 = v_25722 & v_25856;
assign v_25862 = v_25720 & v_25861;
assign v_25864 = v_25766 & v_25863;
assign v_25865 = v_25719 & v_25861;
assign v_25867 = v_25717 & v_25866;
assign v_25869 = v_25772 & v_25868;
assign v_25870 = v_25716 & v_25866;
assign v_25872 = v_25714 & v_25871;
assign v_25874 = v_25778 & v_25873;
assign v_25875 = v_25713 & v_25871;
assign v_25877 = v_25711 & v_25876;
assign v_25879 = v_25784 & v_25878;
assign v_25880 = v_25710 & v_25876;
assign v_25882 = v_25708 & v_25881;
assign v_25884 = v_25790 & v_25883;
assign v_25885 = v_25707 & v_25881;
assign v_25887 = v_25705 & v_25886;
assign v_25889 = v_25796 & v_25888;
assign v_25890 = v_25704 & v_25886;
assign v_25892 = v_25702 & v_25891;
assign v_25894 = v_25802 & v_25893;
assign v_25895 = v_25701 & v_25891;
assign v_25897 = v_25699 & v_25896;
assign v_25899 = v_25808 & v_25898;
assign v_25900 = v_25698 & v_25896;
assign v_25902 = v_25696 & v_25901;
assign v_25904 = v_25814 & v_25903;
assign v_25905 = v_25695 & v_25901;
assign v_25907 = v_25693 & v_25906;
assign v_25909 = v_25820 & v_25908;
assign v_25910 = v_25692 & v_25906;
assign v_25912 = v_25690 & v_25911;
assign v_25914 = v_25826 & v_25913;
assign v_25915 = v_25689 & v_25911;
assign v_25917 = v_25687 & v_25916;
assign v_25919 = v_25832 & v_25918;
assign v_25920 = v_25686 & v_25916;
assign v_25922 = v_25921;
assign v_25924 = v_25836 & v_25923;
assign v_25925 = v_25924;
assign v_25927 = v_25926;
assign v_25929 = ~v_803;
assign v_25930 = ~v_25184;
assign v_25931 = v_25184;
assign v_25932 = ~v_807;
assign v_25933 = ~v_25188;
assign v_25934 = v_25188;
assign v_25935 = ~v_811;
assign v_25936 = ~v_25192;
assign v_25937 = v_25192;
assign v_25938 = ~v_815;
assign v_25939 = ~v_25196;
assign v_25940 = v_25196;
assign v_25941 = ~v_25199;
assign v_25942 = ~v_820;
assign v_25943 = v_820;
assign v_25944 = ~v_25203;
assign v_25945 = ~v_824;
assign v_25946 = v_824;
assign v_25947 = ~v_25207;
assign v_25948 = ~v_828;
assign v_25949 = v_828;
assign v_25950 = ~v_25211;
assign v_25951 = ~v_832;
assign v_25952 = v_832;
assign v_25953 = ~v_25215;
assign v_25954 = ~v_836;
assign v_25955 = v_836;
assign v_25956 = ~v_25219;
assign v_25957 = ~v_840;
assign v_25958 = v_840;
assign v_25959 = ~v_25223;
assign v_25960 = ~v_844;
assign v_25961 = v_844;
assign v_25962 = ~v_25227;
assign v_25963 = ~v_848;
assign v_25964 = v_848;
assign v_25965 = ~v_25231;
assign v_25966 = ~v_852;
assign v_25967 = v_852;
assign v_25968 = ~v_25235;
assign v_25969 = ~v_856;
assign v_25970 = v_856;
assign v_25971 = ~v_25239;
assign v_25972 = ~v_860;
assign v_25973 = v_860;
assign v_25974 = ~v_25243;
assign v_25975 = ~v_864;
assign v_25976 = v_864;
assign v_25977 = ~v_25247;
assign v_25978 = ~v_868;
assign v_25979 = v_25978;
assign v_25981 = v_25980;
assign v_25983 = v_25975 & v_25982;
assign v_25985 = v_25243;
assign v_25987 = v_25984 & v_25986;
assign v_25989 = v_25972 & v_25988;
assign v_25991 = v_25239;
assign v_25993 = v_25990 & v_25992;
assign v_25995 = v_25969 & v_25994;
assign v_25997 = v_25235;
assign v_25999 = v_25996 & v_25998;
assign v_26001 = v_25966 & v_26000;
assign v_26003 = v_25231;
assign v_26005 = v_26002 & v_26004;
assign v_26007 = v_25963 & v_26006;
assign v_26009 = v_25227;
assign v_26011 = v_26008 & v_26010;
assign v_26013 = v_25960 & v_26012;
assign v_26015 = v_25223;
assign v_26017 = v_26014 & v_26016;
assign v_26019 = v_25957 & v_26018;
assign v_26021 = v_25219;
assign v_26023 = v_26020 & v_26022;
assign v_26025 = v_25954 & v_26024;
assign v_26027 = v_25215;
assign v_26029 = v_26026 & v_26028;
assign v_26031 = v_25951 & v_26030;
assign v_26033 = v_25211;
assign v_26035 = v_26032 & v_26034;
assign v_26037 = v_25948 & v_26036;
assign v_26039 = v_25207;
assign v_26041 = v_26038 & v_26040;
assign v_26043 = v_25945 & v_26042;
assign v_26045 = v_25203;
assign v_26047 = v_26044 & v_26046;
assign v_26049 = v_25942 & v_26048;
assign v_26051 = v_25199;
assign v_26053 = v_26050 & v_26052;
assign v_26055 = v_25939 & v_26054;
assign v_26057 = v_815;
assign v_26059 = v_26056 & v_26058;
assign v_26061 = v_25936 & v_26060;
assign v_26063 = v_811;
assign v_26065 = v_26062 & v_26064;
assign v_26067 = v_25933 & v_26066;
assign v_26069 = v_807;
assign v_26071 = v_26068 & v_26070;
assign v_26073 = v_25930 & v_26072;
assign v_26075 = v_803;
assign v_26077 = v_26074 & v_26076;
assign v_26078 = v_26077;
assign v_26080 = v_25247;
assign v_26081 = v_868;
assign v_26082 = v_26081;
assign v_26083 = v_26080 & v_26082;
assign v_26084 = v_26083;
assign v_26085 = v_25975 & v_26084;
assign v_26087 = v_25985 & v_26086;
assign v_26088 = v_25974 & v_26084;
assign v_26090 = v_25972 & v_26089;
assign v_26092 = v_25991 & v_26091;
assign v_26093 = v_25971 & v_26089;
assign v_26095 = v_25969 & v_26094;
assign v_26097 = v_25997 & v_26096;
assign v_26098 = v_25968 & v_26094;
assign v_26100 = v_25966 & v_26099;
assign v_26102 = v_26003 & v_26101;
assign v_26103 = v_25965 & v_26099;
assign v_26105 = v_25963 & v_26104;
assign v_26107 = v_26009 & v_26106;
assign v_26108 = v_25962 & v_26104;
assign v_26110 = v_25960 & v_26109;
assign v_26112 = v_26015 & v_26111;
assign v_26113 = v_25959 & v_26109;
assign v_26115 = v_25957 & v_26114;
assign v_26117 = v_26021 & v_26116;
assign v_26118 = v_25956 & v_26114;
assign v_26120 = v_25954 & v_26119;
assign v_26122 = v_26027 & v_26121;
assign v_26123 = v_25953 & v_26119;
assign v_26125 = v_25951 & v_26124;
assign v_26127 = v_26033 & v_26126;
assign v_26128 = v_25950 & v_26124;
assign v_26130 = v_25948 & v_26129;
assign v_26132 = v_26039 & v_26131;
assign v_26133 = v_25947 & v_26129;
assign v_26135 = v_25945 & v_26134;
assign v_26137 = v_26045 & v_26136;
assign v_26138 = v_25944 & v_26134;
assign v_26140 = v_25942 & v_26139;
assign v_26142 = v_26051 & v_26141;
assign v_26143 = v_25941 & v_26139;
assign v_26145 = v_25939 & v_26144;
assign v_26147 = v_26057 & v_26146;
assign v_26148 = v_25938 & v_26144;
assign v_26150 = v_25936 & v_26149;
assign v_26152 = v_26063 & v_26151;
assign v_26153 = v_25935 & v_26149;
assign v_26155 = v_25933 & v_26154;
assign v_26157 = v_26069 & v_26156;
assign v_26158 = v_25932 & v_26154;
assign v_26160 = v_25930 & v_26159;
assign v_26162 = v_26075 & v_26161;
assign v_26163 = v_25929 & v_26159;
assign v_26165 = v_26164;
assign v_26167 = v_26079 & v_26166;
assign v_26168 = v_26167;
assign v_26170 = v_26169;
assign v_26172 = ~v_1063;
assign v_26173 = ~v_25184;
assign v_26174 = v_25184;
assign v_26175 = ~v_1067;
assign v_26176 = ~v_25188;
assign v_26177 = v_25188;
assign v_26178 = ~v_1071;
assign v_26179 = ~v_25192;
assign v_26180 = v_25192;
assign v_26181 = ~v_1075;
assign v_26182 = ~v_25196;
assign v_26183 = v_25196;
assign v_26184 = ~v_25199;
assign v_26185 = ~v_1080;
assign v_26186 = v_1080;
assign v_26187 = ~v_25203;
assign v_26188 = ~v_1084;
assign v_26189 = v_1084;
assign v_26190 = ~v_25207;
assign v_26191 = ~v_1088;
assign v_26192 = v_1088;
assign v_26193 = ~v_25211;
assign v_26194 = ~v_1092;
assign v_26195 = v_1092;
assign v_26196 = ~v_25215;
assign v_26197 = ~v_1096;
assign v_26198 = v_1096;
assign v_26199 = ~v_25219;
assign v_26200 = ~v_1100;
assign v_26201 = v_1100;
assign v_26202 = ~v_25223;
assign v_26203 = ~v_1104;
assign v_26204 = v_1104;
assign v_26205 = ~v_25227;
assign v_26206 = ~v_1108;
assign v_26207 = v_1108;
assign v_26208 = ~v_25231;
assign v_26209 = ~v_1112;
assign v_26210 = v_1112;
assign v_26211 = ~v_25235;
assign v_26212 = ~v_1116;
assign v_26213 = v_1116;
assign v_26214 = ~v_25239;
assign v_26215 = ~v_1120;
assign v_26216 = v_1120;
assign v_26217 = ~v_25243;
assign v_26218 = ~v_1124;
assign v_26219 = v_1124;
assign v_26220 = ~v_25247;
assign v_26221 = ~v_1128;
assign v_26222 = v_26221;
assign v_26224 = v_26223;
assign v_26226 = v_26218 & v_26225;
assign v_26228 = v_25243;
assign v_26230 = v_26227 & v_26229;
assign v_26232 = v_26215 & v_26231;
assign v_26234 = v_25239;
assign v_26236 = v_26233 & v_26235;
assign v_26238 = v_26212 & v_26237;
assign v_26240 = v_25235;
assign v_26242 = v_26239 & v_26241;
assign v_26244 = v_26209 & v_26243;
assign v_26246 = v_25231;
assign v_26248 = v_26245 & v_26247;
assign v_26250 = v_26206 & v_26249;
assign v_26252 = v_25227;
assign v_26254 = v_26251 & v_26253;
assign v_26256 = v_26203 & v_26255;
assign v_26258 = v_25223;
assign v_26260 = v_26257 & v_26259;
assign v_26262 = v_26200 & v_26261;
assign v_26264 = v_25219;
assign v_26266 = v_26263 & v_26265;
assign v_26268 = v_26197 & v_26267;
assign v_26270 = v_25215;
assign v_26272 = v_26269 & v_26271;
assign v_26274 = v_26194 & v_26273;
assign v_26276 = v_25211;
assign v_26278 = v_26275 & v_26277;
assign v_26280 = v_26191 & v_26279;
assign v_26282 = v_25207;
assign v_26284 = v_26281 & v_26283;
assign v_26286 = v_26188 & v_26285;
assign v_26288 = v_25203;
assign v_26290 = v_26287 & v_26289;
assign v_26292 = v_26185 & v_26291;
assign v_26294 = v_25199;
assign v_26296 = v_26293 & v_26295;
assign v_26298 = v_26182 & v_26297;
assign v_26300 = v_1075;
assign v_26302 = v_26299 & v_26301;
assign v_26304 = v_26179 & v_26303;
assign v_26306 = v_1071;
assign v_26308 = v_26305 & v_26307;
assign v_26310 = v_26176 & v_26309;
assign v_26312 = v_1067;
assign v_26314 = v_26311 & v_26313;
assign v_26316 = v_26173 & v_26315;
assign v_26318 = v_1063;
assign v_26320 = v_26317 & v_26319;
assign v_26321 = v_26320;
assign v_26323 = v_25247;
assign v_26324 = v_1128;
assign v_26325 = v_26324;
assign v_26326 = v_26323 & v_26325;
assign v_26327 = v_26326;
assign v_26328 = v_26218 & v_26327;
assign v_26330 = v_26228 & v_26329;
assign v_26331 = v_26217 & v_26327;
assign v_26333 = v_26215 & v_26332;
assign v_26335 = v_26234 & v_26334;
assign v_26336 = v_26214 & v_26332;
assign v_26338 = v_26212 & v_26337;
assign v_26340 = v_26240 & v_26339;
assign v_26341 = v_26211 & v_26337;
assign v_26343 = v_26209 & v_26342;
assign v_26345 = v_26246 & v_26344;
assign v_26346 = v_26208 & v_26342;
assign v_26348 = v_26206 & v_26347;
assign v_26350 = v_26252 & v_26349;
assign v_26351 = v_26205 & v_26347;
assign v_26353 = v_26203 & v_26352;
assign v_26355 = v_26258 & v_26354;
assign v_26356 = v_26202 & v_26352;
assign v_26358 = v_26200 & v_26357;
assign v_26360 = v_26264 & v_26359;
assign v_26361 = v_26199 & v_26357;
assign v_26363 = v_26197 & v_26362;
assign v_26365 = v_26270 & v_26364;
assign v_26366 = v_26196 & v_26362;
assign v_26368 = v_26194 & v_26367;
assign v_26370 = v_26276 & v_26369;
assign v_26371 = v_26193 & v_26367;
assign v_26373 = v_26191 & v_26372;
assign v_26375 = v_26282 & v_26374;
assign v_26376 = v_26190 & v_26372;
assign v_26378 = v_26188 & v_26377;
assign v_26380 = v_26288 & v_26379;
assign v_26381 = v_26187 & v_26377;
assign v_26383 = v_26185 & v_26382;
assign v_26385 = v_26294 & v_26384;
assign v_26386 = v_26184 & v_26382;
assign v_26388 = v_26182 & v_26387;
assign v_26390 = v_26300 & v_26389;
assign v_26391 = v_26181 & v_26387;
assign v_26393 = v_26179 & v_26392;
assign v_26395 = v_26306 & v_26394;
assign v_26396 = v_26178 & v_26392;
assign v_26398 = v_26176 & v_26397;
assign v_26400 = v_26312 & v_26399;
assign v_26401 = v_26175 & v_26397;
assign v_26403 = v_26173 & v_26402;
assign v_26405 = v_26318 & v_26404;
assign v_26406 = v_26172 & v_26402;
assign v_26408 = v_26407;
assign v_26410 = v_26322 & v_26409;
assign v_26411 = v_26410;
assign v_26413 = v_26412;
assign v_26415 = ~v_1323;
assign v_26416 = ~v_25184;
assign v_26417 = v_25184;
assign v_26418 = ~v_1327;
assign v_26419 = ~v_25188;
assign v_26420 = v_25188;
assign v_26421 = ~v_1331;
assign v_26422 = ~v_25192;
assign v_26423 = v_25192;
assign v_26424 = ~v_1335;
assign v_26425 = ~v_25196;
assign v_26426 = v_25196;
assign v_26427 = ~v_25199;
assign v_26428 = ~v_1340;
assign v_26429 = v_1340;
assign v_26430 = ~v_25203;
assign v_26431 = ~v_1344;
assign v_26432 = v_1344;
assign v_26433 = ~v_25207;
assign v_26434 = ~v_1348;
assign v_26435 = v_1348;
assign v_26436 = ~v_25211;
assign v_26437 = ~v_1352;
assign v_26438 = v_1352;
assign v_26439 = ~v_25215;
assign v_26440 = ~v_1356;
assign v_26441 = v_1356;
assign v_26442 = ~v_25219;
assign v_26443 = ~v_1360;
assign v_26444 = v_1360;
assign v_26445 = ~v_25223;
assign v_26446 = ~v_1364;
assign v_26447 = v_1364;
assign v_26448 = ~v_25227;
assign v_26449 = ~v_1368;
assign v_26450 = v_1368;
assign v_26451 = ~v_25231;
assign v_26452 = ~v_1372;
assign v_26453 = v_1372;
assign v_26454 = ~v_25235;
assign v_26455 = ~v_1376;
assign v_26456 = v_1376;
assign v_26457 = ~v_25239;
assign v_26458 = ~v_1380;
assign v_26459 = v_1380;
assign v_26460 = ~v_25243;
assign v_26461 = ~v_1384;
assign v_26462 = v_1384;
assign v_26463 = ~v_25247;
assign v_26464 = ~v_1388;
assign v_26465 = v_26464;
assign v_26467 = v_26466;
assign v_26469 = v_26461 & v_26468;
assign v_26471 = v_25243;
assign v_26473 = v_26470 & v_26472;
assign v_26475 = v_26458 & v_26474;
assign v_26477 = v_25239;
assign v_26479 = v_26476 & v_26478;
assign v_26481 = v_26455 & v_26480;
assign v_26483 = v_25235;
assign v_26485 = v_26482 & v_26484;
assign v_26487 = v_26452 & v_26486;
assign v_26489 = v_25231;
assign v_26491 = v_26488 & v_26490;
assign v_26493 = v_26449 & v_26492;
assign v_26495 = v_25227;
assign v_26497 = v_26494 & v_26496;
assign v_26499 = v_26446 & v_26498;
assign v_26501 = v_25223;
assign v_26503 = v_26500 & v_26502;
assign v_26505 = v_26443 & v_26504;
assign v_26507 = v_25219;
assign v_26509 = v_26506 & v_26508;
assign v_26511 = v_26440 & v_26510;
assign v_26513 = v_25215;
assign v_26515 = v_26512 & v_26514;
assign v_26517 = v_26437 & v_26516;
assign v_26519 = v_25211;
assign v_26521 = v_26518 & v_26520;
assign v_26523 = v_26434 & v_26522;
assign v_26525 = v_25207;
assign v_26527 = v_26524 & v_26526;
assign v_26529 = v_26431 & v_26528;
assign v_26531 = v_25203;
assign v_26533 = v_26530 & v_26532;
assign v_26535 = v_26428 & v_26534;
assign v_26537 = v_25199;
assign v_26539 = v_26536 & v_26538;
assign v_26541 = v_26425 & v_26540;
assign v_26543 = v_1335;
assign v_26545 = v_26542 & v_26544;
assign v_26547 = v_26422 & v_26546;
assign v_26549 = v_1331;
assign v_26551 = v_26548 & v_26550;
assign v_26553 = v_26419 & v_26552;
assign v_26555 = v_1327;
assign v_26557 = v_26554 & v_26556;
assign v_26559 = v_26416 & v_26558;
assign v_26561 = v_1323;
assign v_26563 = v_26560 & v_26562;
assign v_26564 = v_26563;
assign v_26566 = v_25247;
assign v_26567 = v_1388;
assign v_26568 = v_26567;
assign v_26569 = v_26566 & v_26568;
assign v_26570 = v_26569;
assign v_26571 = v_26461 & v_26570;
assign v_26573 = v_26471 & v_26572;
assign v_26574 = v_26460 & v_26570;
assign v_26576 = v_26458 & v_26575;
assign v_26578 = v_26477 & v_26577;
assign v_26579 = v_26457 & v_26575;
assign v_26581 = v_26455 & v_26580;
assign v_26583 = v_26483 & v_26582;
assign v_26584 = v_26454 & v_26580;
assign v_26586 = v_26452 & v_26585;
assign v_26588 = v_26489 & v_26587;
assign v_26589 = v_26451 & v_26585;
assign v_26591 = v_26449 & v_26590;
assign v_26593 = v_26495 & v_26592;
assign v_26594 = v_26448 & v_26590;
assign v_26596 = v_26446 & v_26595;
assign v_26598 = v_26501 & v_26597;
assign v_26599 = v_26445 & v_26595;
assign v_26601 = v_26443 & v_26600;
assign v_26603 = v_26507 & v_26602;
assign v_26604 = v_26442 & v_26600;
assign v_26606 = v_26440 & v_26605;
assign v_26608 = v_26513 & v_26607;
assign v_26609 = v_26439 & v_26605;
assign v_26611 = v_26437 & v_26610;
assign v_26613 = v_26519 & v_26612;
assign v_26614 = v_26436 & v_26610;
assign v_26616 = v_26434 & v_26615;
assign v_26618 = v_26525 & v_26617;
assign v_26619 = v_26433 & v_26615;
assign v_26621 = v_26431 & v_26620;
assign v_26623 = v_26531 & v_26622;
assign v_26624 = v_26430 & v_26620;
assign v_26626 = v_26428 & v_26625;
assign v_26628 = v_26537 & v_26627;
assign v_26629 = v_26427 & v_26625;
assign v_26631 = v_26425 & v_26630;
assign v_26633 = v_26543 & v_26632;
assign v_26634 = v_26424 & v_26630;
assign v_26636 = v_26422 & v_26635;
assign v_26638 = v_26549 & v_26637;
assign v_26639 = v_26421 & v_26635;
assign v_26641 = v_26419 & v_26640;
assign v_26643 = v_26555 & v_26642;
assign v_26644 = v_26418 & v_26640;
assign v_26646 = v_26416 & v_26645;
assign v_26648 = v_26561 & v_26647;
assign v_26649 = v_26415 & v_26645;
assign v_26651 = v_26650;
assign v_26653 = v_26565 & v_26652;
assign v_26654 = v_26653;
assign v_26656 = v_26655;
assign v_26658 = ~v_1583;
assign v_26659 = ~v_25184;
assign v_26660 = v_25184;
assign v_26661 = ~v_1587;
assign v_26662 = ~v_25188;
assign v_26663 = v_25188;
assign v_26664 = ~v_1591;
assign v_26665 = ~v_25192;
assign v_26666 = v_25192;
assign v_26667 = ~v_1595;
assign v_26668 = ~v_25196;
assign v_26669 = v_25196;
assign v_26670 = ~v_25199;
assign v_26671 = ~v_1600;
assign v_26672 = v_1600;
assign v_26673 = ~v_25203;
assign v_26674 = ~v_1604;
assign v_26675 = v_1604;
assign v_26676 = ~v_25207;
assign v_26677 = ~v_1608;
assign v_26678 = v_1608;
assign v_26679 = ~v_25211;
assign v_26680 = ~v_1612;
assign v_26681 = v_1612;
assign v_26682 = ~v_25215;
assign v_26683 = ~v_1616;
assign v_26684 = v_1616;
assign v_26685 = ~v_25219;
assign v_26686 = ~v_1620;
assign v_26687 = v_1620;
assign v_26688 = ~v_25223;
assign v_26689 = ~v_1624;
assign v_26690 = v_1624;
assign v_26691 = ~v_25227;
assign v_26692 = ~v_1628;
assign v_26693 = v_1628;
assign v_26694 = ~v_25231;
assign v_26695 = ~v_1632;
assign v_26696 = v_1632;
assign v_26697 = ~v_25235;
assign v_26698 = ~v_1636;
assign v_26699 = v_1636;
assign v_26700 = ~v_25239;
assign v_26701 = ~v_1640;
assign v_26702 = v_1640;
assign v_26703 = ~v_25243;
assign v_26704 = ~v_1644;
assign v_26705 = v_1644;
assign v_26706 = ~v_25247;
assign v_26707 = ~v_1648;
assign v_26708 = v_26707;
assign v_26710 = v_26709;
assign v_26712 = v_26704 & v_26711;
assign v_26714 = v_25243;
assign v_26716 = v_26713 & v_26715;
assign v_26718 = v_26701 & v_26717;
assign v_26720 = v_25239;
assign v_26722 = v_26719 & v_26721;
assign v_26724 = v_26698 & v_26723;
assign v_26726 = v_25235;
assign v_26728 = v_26725 & v_26727;
assign v_26730 = v_26695 & v_26729;
assign v_26732 = v_25231;
assign v_26734 = v_26731 & v_26733;
assign v_26736 = v_26692 & v_26735;
assign v_26738 = v_25227;
assign v_26740 = v_26737 & v_26739;
assign v_26742 = v_26689 & v_26741;
assign v_26744 = v_25223;
assign v_26746 = v_26743 & v_26745;
assign v_26748 = v_26686 & v_26747;
assign v_26750 = v_25219;
assign v_26752 = v_26749 & v_26751;
assign v_26754 = v_26683 & v_26753;
assign v_26756 = v_25215;
assign v_26758 = v_26755 & v_26757;
assign v_26760 = v_26680 & v_26759;
assign v_26762 = v_25211;
assign v_26764 = v_26761 & v_26763;
assign v_26766 = v_26677 & v_26765;
assign v_26768 = v_25207;
assign v_26770 = v_26767 & v_26769;
assign v_26772 = v_26674 & v_26771;
assign v_26774 = v_25203;
assign v_26776 = v_26773 & v_26775;
assign v_26778 = v_26671 & v_26777;
assign v_26780 = v_25199;
assign v_26782 = v_26779 & v_26781;
assign v_26784 = v_26668 & v_26783;
assign v_26786 = v_1595;
assign v_26788 = v_26785 & v_26787;
assign v_26790 = v_26665 & v_26789;
assign v_26792 = v_1591;
assign v_26794 = v_26791 & v_26793;
assign v_26796 = v_26662 & v_26795;
assign v_26798 = v_1587;
assign v_26800 = v_26797 & v_26799;
assign v_26802 = v_26659 & v_26801;
assign v_26804 = v_1583;
assign v_26806 = v_26803 & v_26805;
assign v_26807 = v_26806;
assign v_26809 = v_25247;
assign v_26810 = v_1648;
assign v_26811 = v_26810;
assign v_26812 = v_26809 & v_26811;
assign v_26813 = v_26812;
assign v_26814 = v_26704 & v_26813;
assign v_26816 = v_26714 & v_26815;
assign v_26817 = v_26703 & v_26813;
assign v_26819 = v_26701 & v_26818;
assign v_26821 = v_26720 & v_26820;
assign v_26822 = v_26700 & v_26818;
assign v_26824 = v_26698 & v_26823;
assign v_26826 = v_26726 & v_26825;
assign v_26827 = v_26697 & v_26823;
assign v_26829 = v_26695 & v_26828;
assign v_26831 = v_26732 & v_26830;
assign v_26832 = v_26694 & v_26828;
assign v_26834 = v_26692 & v_26833;
assign v_26836 = v_26738 & v_26835;
assign v_26837 = v_26691 & v_26833;
assign v_26839 = v_26689 & v_26838;
assign v_26841 = v_26744 & v_26840;
assign v_26842 = v_26688 & v_26838;
assign v_26844 = v_26686 & v_26843;
assign v_26846 = v_26750 & v_26845;
assign v_26847 = v_26685 & v_26843;
assign v_26849 = v_26683 & v_26848;
assign v_26851 = v_26756 & v_26850;
assign v_26852 = v_26682 & v_26848;
assign v_26854 = v_26680 & v_26853;
assign v_26856 = v_26762 & v_26855;
assign v_26857 = v_26679 & v_26853;
assign v_26859 = v_26677 & v_26858;
assign v_26861 = v_26768 & v_26860;
assign v_26862 = v_26676 & v_26858;
assign v_26864 = v_26674 & v_26863;
assign v_26866 = v_26774 & v_26865;
assign v_26867 = v_26673 & v_26863;
assign v_26869 = v_26671 & v_26868;
assign v_26871 = v_26780 & v_26870;
assign v_26872 = v_26670 & v_26868;
assign v_26874 = v_26668 & v_26873;
assign v_26876 = v_26786 & v_26875;
assign v_26877 = v_26667 & v_26873;
assign v_26879 = v_26665 & v_26878;
assign v_26881 = v_26792 & v_26880;
assign v_26882 = v_26664 & v_26878;
assign v_26884 = v_26662 & v_26883;
assign v_26886 = v_26798 & v_26885;
assign v_26887 = v_26661 & v_26883;
assign v_26889 = v_26659 & v_26888;
assign v_26891 = v_26804 & v_26890;
assign v_26892 = v_26658 & v_26888;
assign v_26894 = v_26893;
assign v_26896 = v_26808 & v_26895;
assign v_26897 = v_26896;
assign v_26899 = v_26898;
assign v_26901 = ~v_1843;
assign v_26902 = ~v_25184;
assign v_26903 = v_25184;
assign v_26904 = ~v_1847;
assign v_26905 = ~v_25188;
assign v_26906 = v_25188;
assign v_26907 = ~v_1851;
assign v_26908 = ~v_25192;
assign v_26909 = v_25192;
assign v_26910 = ~v_1855;
assign v_26911 = ~v_25196;
assign v_26912 = v_25196;
assign v_26913 = ~v_25199;
assign v_26914 = ~v_1860;
assign v_26915 = v_1860;
assign v_26916 = ~v_25203;
assign v_26917 = ~v_1864;
assign v_26918 = v_1864;
assign v_26919 = ~v_25207;
assign v_26920 = ~v_1868;
assign v_26921 = v_1868;
assign v_26922 = ~v_25211;
assign v_26923 = ~v_1872;
assign v_26924 = v_1872;
assign v_26925 = ~v_25215;
assign v_26926 = ~v_1876;
assign v_26927 = v_1876;
assign v_26928 = ~v_25219;
assign v_26929 = ~v_1880;
assign v_26930 = v_1880;
assign v_26931 = ~v_25223;
assign v_26932 = ~v_1884;
assign v_26933 = v_1884;
assign v_26934 = ~v_25227;
assign v_26935 = ~v_1888;
assign v_26936 = v_1888;
assign v_26937 = ~v_25231;
assign v_26938 = ~v_1892;
assign v_26939 = v_1892;
assign v_26940 = ~v_25235;
assign v_26941 = ~v_1896;
assign v_26942 = v_1896;
assign v_26943 = ~v_25239;
assign v_26944 = ~v_1900;
assign v_26945 = v_1900;
assign v_26946 = ~v_25243;
assign v_26947 = ~v_1904;
assign v_26948 = v_1904;
assign v_26949 = ~v_25247;
assign v_26950 = ~v_1908;
assign v_26951 = v_26950;
assign v_26953 = v_26952;
assign v_26955 = v_26947 & v_26954;
assign v_26957 = v_25243;
assign v_26959 = v_26956 & v_26958;
assign v_26961 = v_26944 & v_26960;
assign v_26963 = v_25239;
assign v_26965 = v_26962 & v_26964;
assign v_26967 = v_26941 & v_26966;
assign v_26969 = v_25235;
assign v_26971 = v_26968 & v_26970;
assign v_26973 = v_26938 & v_26972;
assign v_26975 = v_25231;
assign v_26977 = v_26974 & v_26976;
assign v_26979 = v_26935 & v_26978;
assign v_26981 = v_25227;
assign v_26983 = v_26980 & v_26982;
assign v_26985 = v_26932 & v_26984;
assign v_26987 = v_25223;
assign v_26989 = v_26986 & v_26988;
assign v_26991 = v_26929 & v_26990;
assign v_26993 = v_25219;
assign v_26995 = v_26992 & v_26994;
assign v_26997 = v_26926 & v_26996;
assign v_26999 = v_25215;
assign v_27001 = v_26998 & v_27000;
assign v_27003 = v_26923 & v_27002;
assign v_27005 = v_25211;
assign v_27007 = v_27004 & v_27006;
assign v_27009 = v_26920 & v_27008;
assign v_27011 = v_25207;
assign v_27013 = v_27010 & v_27012;
assign v_27015 = v_26917 & v_27014;
assign v_27017 = v_25203;
assign v_27019 = v_27016 & v_27018;
assign v_27021 = v_26914 & v_27020;
assign v_27023 = v_25199;
assign v_27025 = v_27022 & v_27024;
assign v_27027 = v_26911 & v_27026;
assign v_27029 = v_1855;
assign v_27031 = v_27028 & v_27030;
assign v_27033 = v_26908 & v_27032;
assign v_27035 = v_1851;
assign v_27037 = v_27034 & v_27036;
assign v_27039 = v_26905 & v_27038;
assign v_27041 = v_1847;
assign v_27043 = v_27040 & v_27042;
assign v_27045 = v_26902 & v_27044;
assign v_27047 = v_1843;
assign v_27049 = v_27046 & v_27048;
assign v_27050 = v_27049;
assign v_27052 = v_25247;
assign v_27053 = v_1908;
assign v_27054 = v_27053;
assign v_27055 = v_27052 & v_27054;
assign v_27056 = v_27055;
assign v_27057 = v_26947 & v_27056;
assign v_27059 = v_26957 & v_27058;
assign v_27060 = v_26946 & v_27056;
assign v_27062 = v_26944 & v_27061;
assign v_27064 = v_26963 & v_27063;
assign v_27065 = v_26943 & v_27061;
assign v_27067 = v_26941 & v_27066;
assign v_27069 = v_26969 & v_27068;
assign v_27070 = v_26940 & v_27066;
assign v_27072 = v_26938 & v_27071;
assign v_27074 = v_26975 & v_27073;
assign v_27075 = v_26937 & v_27071;
assign v_27077 = v_26935 & v_27076;
assign v_27079 = v_26981 & v_27078;
assign v_27080 = v_26934 & v_27076;
assign v_27082 = v_26932 & v_27081;
assign v_27084 = v_26987 & v_27083;
assign v_27085 = v_26931 & v_27081;
assign v_27087 = v_26929 & v_27086;
assign v_27089 = v_26993 & v_27088;
assign v_27090 = v_26928 & v_27086;
assign v_27092 = v_26926 & v_27091;
assign v_27094 = v_26999 & v_27093;
assign v_27095 = v_26925 & v_27091;
assign v_27097 = v_26923 & v_27096;
assign v_27099 = v_27005 & v_27098;
assign v_27100 = v_26922 & v_27096;
assign v_27102 = v_26920 & v_27101;
assign v_27104 = v_27011 & v_27103;
assign v_27105 = v_26919 & v_27101;
assign v_27107 = v_26917 & v_27106;
assign v_27109 = v_27017 & v_27108;
assign v_27110 = v_26916 & v_27106;
assign v_27112 = v_26914 & v_27111;
assign v_27114 = v_27023 & v_27113;
assign v_27115 = v_26913 & v_27111;
assign v_27117 = v_26911 & v_27116;
assign v_27119 = v_27029 & v_27118;
assign v_27120 = v_26910 & v_27116;
assign v_27122 = v_26908 & v_27121;
assign v_27124 = v_27035 & v_27123;
assign v_27125 = v_26907 & v_27121;
assign v_27127 = v_26905 & v_27126;
assign v_27129 = v_27041 & v_27128;
assign v_27130 = v_26904 & v_27126;
assign v_27132 = v_26902 & v_27131;
assign v_27134 = v_27047 & v_27133;
assign v_27135 = v_26901 & v_27131;
assign v_27137 = v_27136;
assign v_27139 = v_27051 & v_27138;
assign v_27140 = v_27139;
assign v_27142 = v_27141;
assign v_27144 = ~v_2103;
assign v_27145 = ~v_25184;
assign v_27146 = v_25184;
assign v_27147 = ~v_2107;
assign v_27148 = ~v_25188;
assign v_27149 = v_25188;
assign v_27150 = ~v_2111;
assign v_27151 = ~v_25192;
assign v_27152 = v_25192;
assign v_27153 = ~v_2115;
assign v_27154 = ~v_25196;
assign v_27155 = v_25196;
assign v_27156 = ~v_25199;
assign v_27157 = ~v_2120;
assign v_27158 = v_2120;
assign v_27159 = ~v_25203;
assign v_27160 = ~v_2124;
assign v_27161 = v_2124;
assign v_27162 = ~v_25207;
assign v_27163 = ~v_2128;
assign v_27164 = v_2128;
assign v_27165 = ~v_25211;
assign v_27166 = ~v_2132;
assign v_27167 = v_2132;
assign v_27168 = ~v_25215;
assign v_27169 = ~v_2136;
assign v_27170 = v_2136;
assign v_27171 = ~v_25219;
assign v_27172 = ~v_2140;
assign v_27173 = v_2140;
assign v_27174 = ~v_25223;
assign v_27175 = ~v_2144;
assign v_27176 = v_2144;
assign v_27177 = ~v_25227;
assign v_27178 = ~v_2148;
assign v_27179 = v_2148;
assign v_27180 = ~v_25231;
assign v_27181 = ~v_2152;
assign v_27182 = v_2152;
assign v_27183 = ~v_25235;
assign v_27184 = ~v_2156;
assign v_27185 = v_2156;
assign v_27186 = ~v_25239;
assign v_27187 = ~v_2160;
assign v_27188 = v_2160;
assign v_27189 = ~v_25243;
assign v_27190 = ~v_2164;
assign v_27191 = v_2164;
assign v_27192 = ~v_25247;
assign v_27193 = ~v_2168;
assign v_27194 = v_27193;
assign v_27196 = v_27195;
assign v_27198 = v_27190 & v_27197;
assign v_27200 = v_25243;
assign v_27202 = v_27199 & v_27201;
assign v_27204 = v_27187 & v_27203;
assign v_27206 = v_25239;
assign v_27208 = v_27205 & v_27207;
assign v_27210 = v_27184 & v_27209;
assign v_27212 = v_25235;
assign v_27214 = v_27211 & v_27213;
assign v_27216 = v_27181 & v_27215;
assign v_27218 = v_25231;
assign v_27220 = v_27217 & v_27219;
assign v_27222 = v_27178 & v_27221;
assign v_27224 = v_25227;
assign v_27226 = v_27223 & v_27225;
assign v_27228 = v_27175 & v_27227;
assign v_27230 = v_25223;
assign v_27232 = v_27229 & v_27231;
assign v_27234 = v_27172 & v_27233;
assign v_27236 = v_25219;
assign v_27238 = v_27235 & v_27237;
assign v_27240 = v_27169 & v_27239;
assign v_27242 = v_25215;
assign v_27244 = v_27241 & v_27243;
assign v_27246 = v_27166 & v_27245;
assign v_27248 = v_25211;
assign v_27250 = v_27247 & v_27249;
assign v_27252 = v_27163 & v_27251;
assign v_27254 = v_25207;
assign v_27256 = v_27253 & v_27255;
assign v_27258 = v_27160 & v_27257;
assign v_27260 = v_25203;
assign v_27262 = v_27259 & v_27261;
assign v_27264 = v_27157 & v_27263;
assign v_27266 = v_25199;
assign v_27268 = v_27265 & v_27267;
assign v_27270 = v_27154 & v_27269;
assign v_27272 = v_2115;
assign v_27274 = v_27271 & v_27273;
assign v_27276 = v_27151 & v_27275;
assign v_27278 = v_2111;
assign v_27280 = v_27277 & v_27279;
assign v_27282 = v_27148 & v_27281;
assign v_27284 = v_2107;
assign v_27286 = v_27283 & v_27285;
assign v_27288 = v_27145 & v_27287;
assign v_27290 = v_2103;
assign v_27292 = v_27289 & v_27291;
assign v_27293 = v_27292;
assign v_27295 = v_25247;
assign v_27296 = v_2168;
assign v_27297 = v_27296;
assign v_27298 = v_27295 & v_27297;
assign v_27299 = v_27298;
assign v_27300 = v_27190 & v_27299;
assign v_27302 = v_27200 & v_27301;
assign v_27303 = v_27189 & v_27299;
assign v_27305 = v_27187 & v_27304;
assign v_27307 = v_27206 & v_27306;
assign v_27308 = v_27186 & v_27304;
assign v_27310 = v_27184 & v_27309;
assign v_27312 = v_27212 & v_27311;
assign v_27313 = v_27183 & v_27309;
assign v_27315 = v_27181 & v_27314;
assign v_27317 = v_27218 & v_27316;
assign v_27318 = v_27180 & v_27314;
assign v_27320 = v_27178 & v_27319;
assign v_27322 = v_27224 & v_27321;
assign v_27323 = v_27177 & v_27319;
assign v_27325 = v_27175 & v_27324;
assign v_27327 = v_27230 & v_27326;
assign v_27328 = v_27174 & v_27324;
assign v_27330 = v_27172 & v_27329;
assign v_27332 = v_27236 & v_27331;
assign v_27333 = v_27171 & v_27329;
assign v_27335 = v_27169 & v_27334;
assign v_27337 = v_27242 & v_27336;
assign v_27338 = v_27168 & v_27334;
assign v_27340 = v_27166 & v_27339;
assign v_27342 = v_27248 & v_27341;
assign v_27343 = v_27165 & v_27339;
assign v_27345 = v_27163 & v_27344;
assign v_27347 = v_27254 & v_27346;
assign v_27348 = v_27162 & v_27344;
assign v_27350 = v_27160 & v_27349;
assign v_27352 = v_27260 & v_27351;
assign v_27353 = v_27159 & v_27349;
assign v_27355 = v_27157 & v_27354;
assign v_27357 = v_27266 & v_27356;
assign v_27358 = v_27156 & v_27354;
assign v_27360 = v_27154 & v_27359;
assign v_27362 = v_27272 & v_27361;
assign v_27363 = v_27153 & v_27359;
assign v_27365 = v_27151 & v_27364;
assign v_27367 = v_27278 & v_27366;
assign v_27368 = v_27150 & v_27364;
assign v_27370 = v_27148 & v_27369;
assign v_27372 = v_27284 & v_27371;
assign v_27373 = v_27147 & v_27369;
assign v_27375 = v_27145 & v_27374;
assign v_27377 = v_27290 & v_27376;
assign v_27378 = v_27144 & v_27374;
assign v_27380 = v_27379;
assign v_27382 = v_27294 & v_27381;
assign v_27383 = v_27382;
assign v_27385 = v_27384;
assign v_27387 = ~v_2363;
assign v_27388 = ~v_25184;
assign v_27389 = v_25184;
assign v_27390 = ~v_2367;
assign v_27391 = ~v_25188;
assign v_27392 = v_25188;
assign v_27393 = ~v_2371;
assign v_27394 = ~v_25192;
assign v_27395 = v_25192;
assign v_27396 = ~v_2375;
assign v_27397 = ~v_25196;
assign v_27398 = v_25196;
assign v_27399 = ~v_25199;
assign v_27400 = ~v_2380;
assign v_27401 = v_2380;
assign v_27402 = ~v_25203;
assign v_27403 = ~v_2384;
assign v_27404 = v_2384;
assign v_27405 = ~v_25207;
assign v_27406 = ~v_2388;
assign v_27407 = v_2388;
assign v_27408 = ~v_25211;
assign v_27409 = ~v_2392;
assign v_27410 = v_2392;
assign v_27411 = ~v_25215;
assign v_27412 = ~v_2396;
assign v_27413 = v_2396;
assign v_27414 = ~v_25219;
assign v_27415 = ~v_2400;
assign v_27416 = v_2400;
assign v_27417 = ~v_25223;
assign v_27418 = ~v_2404;
assign v_27419 = v_2404;
assign v_27420 = ~v_25227;
assign v_27421 = ~v_2408;
assign v_27422 = v_2408;
assign v_27423 = ~v_25231;
assign v_27424 = ~v_2412;
assign v_27425 = v_2412;
assign v_27426 = ~v_25235;
assign v_27427 = ~v_2416;
assign v_27428 = v_2416;
assign v_27429 = ~v_25239;
assign v_27430 = ~v_2420;
assign v_27431 = v_2420;
assign v_27432 = ~v_25243;
assign v_27433 = ~v_2424;
assign v_27434 = v_2424;
assign v_27435 = ~v_25247;
assign v_27436 = ~v_2428;
assign v_27437 = v_27436;
assign v_27439 = v_27438;
assign v_27441 = v_27433 & v_27440;
assign v_27443 = v_25243;
assign v_27445 = v_27442 & v_27444;
assign v_27447 = v_27430 & v_27446;
assign v_27449 = v_25239;
assign v_27451 = v_27448 & v_27450;
assign v_27453 = v_27427 & v_27452;
assign v_27455 = v_25235;
assign v_27457 = v_27454 & v_27456;
assign v_27459 = v_27424 & v_27458;
assign v_27461 = v_25231;
assign v_27463 = v_27460 & v_27462;
assign v_27465 = v_27421 & v_27464;
assign v_27467 = v_25227;
assign v_27469 = v_27466 & v_27468;
assign v_27471 = v_27418 & v_27470;
assign v_27473 = v_25223;
assign v_27475 = v_27472 & v_27474;
assign v_27477 = v_27415 & v_27476;
assign v_27479 = v_25219;
assign v_27481 = v_27478 & v_27480;
assign v_27483 = v_27412 & v_27482;
assign v_27485 = v_25215;
assign v_27487 = v_27484 & v_27486;
assign v_27489 = v_27409 & v_27488;
assign v_27491 = v_25211;
assign v_27493 = v_27490 & v_27492;
assign v_27495 = v_27406 & v_27494;
assign v_27497 = v_25207;
assign v_27499 = v_27496 & v_27498;
assign v_27501 = v_27403 & v_27500;
assign v_27503 = v_25203;
assign v_27505 = v_27502 & v_27504;
assign v_27507 = v_27400 & v_27506;
assign v_27509 = v_25199;
assign v_27511 = v_27508 & v_27510;
assign v_27513 = v_27397 & v_27512;
assign v_27515 = v_2375;
assign v_27517 = v_27514 & v_27516;
assign v_27519 = v_27394 & v_27518;
assign v_27521 = v_2371;
assign v_27523 = v_27520 & v_27522;
assign v_27525 = v_27391 & v_27524;
assign v_27527 = v_2367;
assign v_27529 = v_27526 & v_27528;
assign v_27531 = v_27388 & v_27530;
assign v_27533 = v_2363;
assign v_27535 = v_27532 & v_27534;
assign v_27536 = v_27535;
assign v_27538 = v_25247;
assign v_27539 = v_2428;
assign v_27540 = v_27539;
assign v_27541 = v_27538 & v_27540;
assign v_27542 = v_27541;
assign v_27543 = v_27433 & v_27542;
assign v_27545 = v_27443 & v_27544;
assign v_27546 = v_27432 & v_27542;
assign v_27548 = v_27430 & v_27547;
assign v_27550 = v_27449 & v_27549;
assign v_27551 = v_27429 & v_27547;
assign v_27553 = v_27427 & v_27552;
assign v_27555 = v_27455 & v_27554;
assign v_27556 = v_27426 & v_27552;
assign v_27558 = v_27424 & v_27557;
assign v_27560 = v_27461 & v_27559;
assign v_27561 = v_27423 & v_27557;
assign v_27563 = v_27421 & v_27562;
assign v_27565 = v_27467 & v_27564;
assign v_27566 = v_27420 & v_27562;
assign v_27568 = v_27418 & v_27567;
assign v_27570 = v_27473 & v_27569;
assign v_27571 = v_27417 & v_27567;
assign v_27573 = v_27415 & v_27572;
assign v_27575 = v_27479 & v_27574;
assign v_27576 = v_27414 & v_27572;
assign v_27578 = v_27412 & v_27577;
assign v_27580 = v_27485 & v_27579;
assign v_27581 = v_27411 & v_27577;
assign v_27583 = v_27409 & v_27582;
assign v_27585 = v_27491 & v_27584;
assign v_27586 = v_27408 & v_27582;
assign v_27588 = v_27406 & v_27587;
assign v_27590 = v_27497 & v_27589;
assign v_27591 = v_27405 & v_27587;
assign v_27593 = v_27403 & v_27592;
assign v_27595 = v_27503 & v_27594;
assign v_27596 = v_27402 & v_27592;
assign v_27598 = v_27400 & v_27597;
assign v_27600 = v_27509 & v_27599;
assign v_27601 = v_27399 & v_27597;
assign v_27603 = v_27397 & v_27602;
assign v_27605 = v_27515 & v_27604;
assign v_27606 = v_27396 & v_27602;
assign v_27608 = v_27394 & v_27607;
assign v_27610 = v_27521 & v_27609;
assign v_27611 = v_27393 & v_27607;
assign v_27613 = v_27391 & v_27612;
assign v_27615 = v_27527 & v_27614;
assign v_27616 = v_27390 & v_27612;
assign v_27618 = v_27388 & v_27617;
assign v_27620 = v_27533 & v_27619;
assign v_27621 = v_27387 & v_27617;
assign v_27623 = v_27622;
assign v_27625 = v_27537 & v_27624;
assign v_27626 = v_27625;
assign v_27628 = v_27627;
assign v_27630 = ~v_2623;
assign v_27631 = ~v_25184;
assign v_27632 = v_25184;
assign v_27633 = ~v_2627;
assign v_27634 = ~v_25188;
assign v_27635 = v_25188;
assign v_27636 = ~v_2631;
assign v_27637 = ~v_25192;
assign v_27638 = v_25192;
assign v_27639 = ~v_2635;
assign v_27640 = ~v_25196;
assign v_27641 = v_25196;
assign v_27642 = ~v_25199;
assign v_27643 = ~v_2640;
assign v_27644 = v_2640;
assign v_27645 = ~v_25203;
assign v_27646 = ~v_2644;
assign v_27647 = v_2644;
assign v_27648 = ~v_25207;
assign v_27649 = ~v_2648;
assign v_27650 = v_2648;
assign v_27651 = ~v_25211;
assign v_27652 = ~v_2652;
assign v_27653 = v_2652;
assign v_27654 = ~v_25215;
assign v_27655 = ~v_2656;
assign v_27656 = v_2656;
assign v_27657 = ~v_25219;
assign v_27658 = ~v_2660;
assign v_27659 = v_2660;
assign v_27660 = ~v_25223;
assign v_27661 = ~v_2664;
assign v_27662 = v_2664;
assign v_27663 = ~v_25227;
assign v_27664 = ~v_2668;
assign v_27665 = v_2668;
assign v_27666 = ~v_25231;
assign v_27667 = ~v_2672;
assign v_27668 = v_2672;
assign v_27669 = ~v_25235;
assign v_27670 = ~v_2676;
assign v_27671 = v_2676;
assign v_27672 = ~v_25239;
assign v_27673 = ~v_2680;
assign v_27674 = v_2680;
assign v_27675 = ~v_25243;
assign v_27676 = ~v_2684;
assign v_27677 = v_2684;
assign v_27678 = ~v_25247;
assign v_27679 = ~v_2688;
assign v_27680 = v_27679;
assign v_27682 = v_27681;
assign v_27684 = v_27676 & v_27683;
assign v_27686 = v_25243;
assign v_27688 = v_27685 & v_27687;
assign v_27690 = v_27673 & v_27689;
assign v_27692 = v_25239;
assign v_27694 = v_27691 & v_27693;
assign v_27696 = v_27670 & v_27695;
assign v_27698 = v_25235;
assign v_27700 = v_27697 & v_27699;
assign v_27702 = v_27667 & v_27701;
assign v_27704 = v_25231;
assign v_27706 = v_27703 & v_27705;
assign v_27708 = v_27664 & v_27707;
assign v_27710 = v_25227;
assign v_27712 = v_27709 & v_27711;
assign v_27714 = v_27661 & v_27713;
assign v_27716 = v_25223;
assign v_27718 = v_27715 & v_27717;
assign v_27720 = v_27658 & v_27719;
assign v_27722 = v_25219;
assign v_27724 = v_27721 & v_27723;
assign v_27726 = v_27655 & v_27725;
assign v_27728 = v_25215;
assign v_27730 = v_27727 & v_27729;
assign v_27732 = v_27652 & v_27731;
assign v_27734 = v_25211;
assign v_27736 = v_27733 & v_27735;
assign v_27738 = v_27649 & v_27737;
assign v_27740 = v_25207;
assign v_27742 = v_27739 & v_27741;
assign v_27744 = v_27646 & v_27743;
assign v_27746 = v_25203;
assign v_27748 = v_27745 & v_27747;
assign v_27750 = v_27643 & v_27749;
assign v_27752 = v_25199;
assign v_27754 = v_27751 & v_27753;
assign v_27756 = v_27640 & v_27755;
assign v_27758 = v_2635;
assign v_27760 = v_27757 & v_27759;
assign v_27762 = v_27637 & v_27761;
assign v_27764 = v_2631;
assign v_27766 = v_27763 & v_27765;
assign v_27768 = v_27634 & v_27767;
assign v_27770 = v_2627;
assign v_27772 = v_27769 & v_27771;
assign v_27774 = v_27631 & v_27773;
assign v_27776 = v_2623;
assign v_27778 = v_27775 & v_27777;
assign v_27779 = v_27778;
assign v_27781 = v_25247;
assign v_27782 = v_2688;
assign v_27783 = v_27782;
assign v_27784 = v_27781 & v_27783;
assign v_27785 = v_27784;
assign v_27786 = v_27676 & v_27785;
assign v_27788 = v_27686 & v_27787;
assign v_27789 = v_27675 & v_27785;
assign v_27791 = v_27673 & v_27790;
assign v_27793 = v_27692 & v_27792;
assign v_27794 = v_27672 & v_27790;
assign v_27796 = v_27670 & v_27795;
assign v_27798 = v_27698 & v_27797;
assign v_27799 = v_27669 & v_27795;
assign v_27801 = v_27667 & v_27800;
assign v_27803 = v_27704 & v_27802;
assign v_27804 = v_27666 & v_27800;
assign v_27806 = v_27664 & v_27805;
assign v_27808 = v_27710 & v_27807;
assign v_27809 = v_27663 & v_27805;
assign v_27811 = v_27661 & v_27810;
assign v_27813 = v_27716 & v_27812;
assign v_27814 = v_27660 & v_27810;
assign v_27816 = v_27658 & v_27815;
assign v_27818 = v_27722 & v_27817;
assign v_27819 = v_27657 & v_27815;
assign v_27821 = v_27655 & v_27820;
assign v_27823 = v_27728 & v_27822;
assign v_27824 = v_27654 & v_27820;
assign v_27826 = v_27652 & v_27825;
assign v_27828 = v_27734 & v_27827;
assign v_27829 = v_27651 & v_27825;
assign v_27831 = v_27649 & v_27830;
assign v_27833 = v_27740 & v_27832;
assign v_27834 = v_27648 & v_27830;
assign v_27836 = v_27646 & v_27835;
assign v_27838 = v_27746 & v_27837;
assign v_27839 = v_27645 & v_27835;
assign v_27841 = v_27643 & v_27840;
assign v_27843 = v_27752 & v_27842;
assign v_27844 = v_27642 & v_27840;
assign v_27846 = v_27640 & v_27845;
assign v_27848 = v_27758 & v_27847;
assign v_27849 = v_27639 & v_27845;
assign v_27851 = v_27637 & v_27850;
assign v_27853 = v_27764 & v_27852;
assign v_27854 = v_27636 & v_27850;
assign v_27856 = v_27634 & v_27855;
assign v_27858 = v_27770 & v_27857;
assign v_27859 = v_27633 & v_27855;
assign v_27861 = v_27631 & v_27860;
assign v_27863 = v_27776 & v_27862;
assign v_27864 = v_27630 & v_27860;
assign v_27866 = v_27865;
assign v_27868 = v_27780 & v_27867;
assign v_27869 = v_27868;
assign v_27871 = v_27870;
assign v_27873 = ~v_2883;
assign v_27874 = ~v_25184;
assign v_27875 = v_25184;
assign v_27876 = ~v_2887;
assign v_27877 = ~v_25188;
assign v_27878 = v_25188;
assign v_27879 = ~v_2891;
assign v_27880 = ~v_25192;
assign v_27881 = v_25192;
assign v_27882 = ~v_2895;
assign v_27883 = ~v_25196;
assign v_27884 = v_25196;
assign v_27885 = ~v_25199;
assign v_27886 = ~v_2900;
assign v_27887 = v_2900;
assign v_27888 = ~v_25203;
assign v_27889 = ~v_2904;
assign v_27890 = v_2904;
assign v_27891 = ~v_25207;
assign v_27892 = ~v_2908;
assign v_27893 = v_2908;
assign v_27894 = ~v_25211;
assign v_27895 = ~v_2912;
assign v_27896 = v_2912;
assign v_27897 = ~v_25215;
assign v_27898 = ~v_2916;
assign v_27899 = v_2916;
assign v_27900 = ~v_25219;
assign v_27901 = ~v_2920;
assign v_27902 = v_2920;
assign v_27903 = ~v_25223;
assign v_27904 = ~v_2924;
assign v_27905 = v_2924;
assign v_27906 = ~v_25227;
assign v_27907 = ~v_2928;
assign v_27908 = v_2928;
assign v_27909 = ~v_25231;
assign v_27910 = ~v_2932;
assign v_27911 = v_2932;
assign v_27912 = ~v_25235;
assign v_27913 = ~v_2936;
assign v_27914 = v_2936;
assign v_27915 = ~v_25239;
assign v_27916 = ~v_2940;
assign v_27917 = v_2940;
assign v_27918 = ~v_25243;
assign v_27919 = ~v_2944;
assign v_27920 = v_2944;
assign v_27921 = ~v_25247;
assign v_27922 = ~v_2948;
assign v_27923 = v_27922;
assign v_27925 = v_27924;
assign v_27927 = v_27919 & v_27926;
assign v_27929 = v_25243;
assign v_27931 = v_27928 & v_27930;
assign v_27933 = v_27916 & v_27932;
assign v_27935 = v_25239;
assign v_27937 = v_27934 & v_27936;
assign v_27939 = v_27913 & v_27938;
assign v_27941 = v_25235;
assign v_27943 = v_27940 & v_27942;
assign v_27945 = v_27910 & v_27944;
assign v_27947 = v_25231;
assign v_27949 = v_27946 & v_27948;
assign v_27951 = v_27907 & v_27950;
assign v_27953 = v_25227;
assign v_27955 = v_27952 & v_27954;
assign v_27957 = v_27904 & v_27956;
assign v_27959 = v_25223;
assign v_27961 = v_27958 & v_27960;
assign v_27963 = v_27901 & v_27962;
assign v_27965 = v_25219;
assign v_27967 = v_27964 & v_27966;
assign v_27969 = v_27898 & v_27968;
assign v_27971 = v_25215;
assign v_27973 = v_27970 & v_27972;
assign v_27975 = v_27895 & v_27974;
assign v_27977 = v_25211;
assign v_27979 = v_27976 & v_27978;
assign v_27981 = v_27892 & v_27980;
assign v_27983 = v_25207;
assign v_27985 = v_27982 & v_27984;
assign v_27987 = v_27889 & v_27986;
assign v_27989 = v_25203;
assign v_27991 = v_27988 & v_27990;
assign v_27993 = v_27886 & v_27992;
assign v_27995 = v_25199;
assign v_27997 = v_27994 & v_27996;
assign v_27999 = v_27883 & v_27998;
assign v_28001 = v_2895;
assign v_28003 = v_28000 & v_28002;
assign v_28005 = v_27880 & v_28004;
assign v_28007 = v_2891;
assign v_28009 = v_28006 & v_28008;
assign v_28011 = v_27877 & v_28010;
assign v_28013 = v_2887;
assign v_28015 = v_28012 & v_28014;
assign v_28017 = v_27874 & v_28016;
assign v_28019 = v_2883;
assign v_28021 = v_28018 & v_28020;
assign v_28022 = v_28021;
assign v_28024 = v_25247;
assign v_28025 = v_2948;
assign v_28026 = v_28025;
assign v_28027 = v_28024 & v_28026;
assign v_28028 = v_28027;
assign v_28029 = v_27919 & v_28028;
assign v_28031 = v_27929 & v_28030;
assign v_28032 = v_27918 & v_28028;
assign v_28034 = v_27916 & v_28033;
assign v_28036 = v_27935 & v_28035;
assign v_28037 = v_27915 & v_28033;
assign v_28039 = v_27913 & v_28038;
assign v_28041 = v_27941 & v_28040;
assign v_28042 = v_27912 & v_28038;
assign v_28044 = v_27910 & v_28043;
assign v_28046 = v_27947 & v_28045;
assign v_28047 = v_27909 & v_28043;
assign v_28049 = v_27907 & v_28048;
assign v_28051 = v_27953 & v_28050;
assign v_28052 = v_27906 & v_28048;
assign v_28054 = v_27904 & v_28053;
assign v_28056 = v_27959 & v_28055;
assign v_28057 = v_27903 & v_28053;
assign v_28059 = v_27901 & v_28058;
assign v_28061 = v_27965 & v_28060;
assign v_28062 = v_27900 & v_28058;
assign v_28064 = v_27898 & v_28063;
assign v_28066 = v_27971 & v_28065;
assign v_28067 = v_27897 & v_28063;
assign v_28069 = v_27895 & v_28068;
assign v_28071 = v_27977 & v_28070;
assign v_28072 = v_27894 & v_28068;
assign v_28074 = v_27892 & v_28073;
assign v_28076 = v_27983 & v_28075;
assign v_28077 = v_27891 & v_28073;
assign v_28079 = v_27889 & v_28078;
assign v_28081 = v_27989 & v_28080;
assign v_28082 = v_27888 & v_28078;
assign v_28084 = v_27886 & v_28083;
assign v_28086 = v_27995 & v_28085;
assign v_28087 = v_27885 & v_28083;
assign v_28089 = v_27883 & v_28088;
assign v_28091 = v_28001 & v_28090;
assign v_28092 = v_27882 & v_28088;
assign v_28094 = v_27880 & v_28093;
assign v_28096 = v_28007 & v_28095;
assign v_28097 = v_27879 & v_28093;
assign v_28099 = v_27877 & v_28098;
assign v_28101 = v_28013 & v_28100;
assign v_28102 = v_27876 & v_28098;
assign v_28104 = v_27874 & v_28103;
assign v_28106 = v_28019 & v_28105;
assign v_28107 = v_27873 & v_28103;
assign v_28109 = v_28108;
assign v_28111 = v_28023 & v_28110;
assign v_28112 = v_28111;
assign v_28114 = v_28113;
assign v_28116 = ~v_3143;
assign v_28117 = ~v_25184;
assign v_28118 = v_25184;
assign v_28119 = ~v_3147;
assign v_28120 = ~v_25188;
assign v_28121 = v_25188;
assign v_28122 = ~v_3151;
assign v_28123 = ~v_25192;
assign v_28124 = v_25192;
assign v_28125 = ~v_3155;
assign v_28126 = ~v_25196;
assign v_28127 = v_25196;
assign v_28128 = ~v_25199;
assign v_28129 = ~v_3160;
assign v_28130 = v_3160;
assign v_28131 = ~v_25203;
assign v_28132 = ~v_3164;
assign v_28133 = v_3164;
assign v_28134 = ~v_25207;
assign v_28135 = ~v_3168;
assign v_28136 = v_3168;
assign v_28137 = ~v_25211;
assign v_28138 = ~v_3172;
assign v_28139 = v_3172;
assign v_28140 = ~v_25215;
assign v_28141 = ~v_3176;
assign v_28142 = v_3176;
assign v_28143 = ~v_25219;
assign v_28144 = ~v_3180;
assign v_28145 = v_3180;
assign v_28146 = ~v_25223;
assign v_28147 = ~v_3184;
assign v_28148 = v_3184;
assign v_28149 = ~v_25227;
assign v_28150 = ~v_3188;
assign v_28151 = v_3188;
assign v_28152 = ~v_25231;
assign v_28153 = ~v_3192;
assign v_28154 = v_3192;
assign v_28155 = ~v_25235;
assign v_28156 = ~v_3196;
assign v_28157 = v_3196;
assign v_28158 = ~v_25239;
assign v_28159 = ~v_3200;
assign v_28160 = v_3200;
assign v_28161 = ~v_25243;
assign v_28162 = ~v_3204;
assign v_28163 = v_3204;
assign v_28164 = ~v_25247;
assign v_28165 = ~v_3208;
assign v_28166 = v_28165;
assign v_28168 = v_28167;
assign v_28170 = v_28162 & v_28169;
assign v_28172 = v_25243;
assign v_28174 = v_28171 & v_28173;
assign v_28176 = v_28159 & v_28175;
assign v_28178 = v_25239;
assign v_28180 = v_28177 & v_28179;
assign v_28182 = v_28156 & v_28181;
assign v_28184 = v_25235;
assign v_28186 = v_28183 & v_28185;
assign v_28188 = v_28153 & v_28187;
assign v_28190 = v_25231;
assign v_28192 = v_28189 & v_28191;
assign v_28194 = v_28150 & v_28193;
assign v_28196 = v_25227;
assign v_28198 = v_28195 & v_28197;
assign v_28200 = v_28147 & v_28199;
assign v_28202 = v_25223;
assign v_28204 = v_28201 & v_28203;
assign v_28206 = v_28144 & v_28205;
assign v_28208 = v_25219;
assign v_28210 = v_28207 & v_28209;
assign v_28212 = v_28141 & v_28211;
assign v_28214 = v_25215;
assign v_28216 = v_28213 & v_28215;
assign v_28218 = v_28138 & v_28217;
assign v_28220 = v_25211;
assign v_28222 = v_28219 & v_28221;
assign v_28224 = v_28135 & v_28223;
assign v_28226 = v_25207;
assign v_28228 = v_28225 & v_28227;
assign v_28230 = v_28132 & v_28229;
assign v_28232 = v_25203;
assign v_28234 = v_28231 & v_28233;
assign v_28236 = v_28129 & v_28235;
assign v_28238 = v_25199;
assign v_28240 = v_28237 & v_28239;
assign v_28242 = v_28126 & v_28241;
assign v_28244 = v_3155;
assign v_28246 = v_28243 & v_28245;
assign v_28248 = v_28123 & v_28247;
assign v_28250 = v_3151;
assign v_28252 = v_28249 & v_28251;
assign v_28254 = v_28120 & v_28253;
assign v_28256 = v_3147;
assign v_28258 = v_28255 & v_28257;
assign v_28260 = v_28117 & v_28259;
assign v_28262 = v_3143;
assign v_28264 = v_28261 & v_28263;
assign v_28265 = v_28264;
assign v_28267 = v_25247;
assign v_28268 = v_3208;
assign v_28269 = v_28268;
assign v_28270 = v_28267 & v_28269;
assign v_28271 = v_28270;
assign v_28272 = v_28162 & v_28271;
assign v_28274 = v_28172 & v_28273;
assign v_28275 = v_28161 & v_28271;
assign v_28277 = v_28159 & v_28276;
assign v_28279 = v_28178 & v_28278;
assign v_28280 = v_28158 & v_28276;
assign v_28282 = v_28156 & v_28281;
assign v_28284 = v_28184 & v_28283;
assign v_28285 = v_28155 & v_28281;
assign v_28287 = v_28153 & v_28286;
assign v_28289 = v_28190 & v_28288;
assign v_28290 = v_28152 & v_28286;
assign v_28292 = v_28150 & v_28291;
assign v_28294 = v_28196 & v_28293;
assign v_28295 = v_28149 & v_28291;
assign v_28297 = v_28147 & v_28296;
assign v_28299 = v_28202 & v_28298;
assign v_28300 = v_28146 & v_28296;
assign v_28302 = v_28144 & v_28301;
assign v_28304 = v_28208 & v_28303;
assign v_28305 = v_28143 & v_28301;
assign v_28307 = v_28141 & v_28306;
assign v_28309 = v_28214 & v_28308;
assign v_28310 = v_28140 & v_28306;
assign v_28312 = v_28138 & v_28311;
assign v_28314 = v_28220 & v_28313;
assign v_28315 = v_28137 & v_28311;
assign v_28317 = v_28135 & v_28316;
assign v_28319 = v_28226 & v_28318;
assign v_28320 = v_28134 & v_28316;
assign v_28322 = v_28132 & v_28321;
assign v_28324 = v_28232 & v_28323;
assign v_28325 = v_28131 & v_28321;
assign v_28327 = v_28129 & v_28326;
assign v_28329 = v_28238 & v_28328;
assign v_28330 = v_28128 & v_28326;
assign v_28332 = v_28126 & v_28331;
assign v_28334 = v_28244 & v_28333;
assign v_28335 = v_28125 & v_28331;
assign v_28337 = v_28123 & v_28336;
assign v_28339 = v_28250 & v_28338;
assign v_28340 = v_28122 & v_28336;
assign v_28342 = v_28120 & v_28341;
assign v_28344 = v_28256 & v_28343;
assign v_28345 = v_28119 & v_28341;
assign v_28347 = v_28117 & v_28346;
assign v_28349 = v_28262 & v_28348;
assign v_28350 = v_28116 & v_28346;
assign v_28352 = v_28351;
assign v_28354 = v_28266 & v_28353;
assign v_28355 = v_28354;
assign v_28357 = v_28356;
assign v_28359 = ~v_3403;
assign v_28360 = ~v_25184;
assign v_28361 = v_25184;
assign v_28362 = ~v_3407;
assign v_28363 = ~v_25188;
assign v_28364 = v_25188;
assign v_28365 = ~v_3411;
assign v_28366 = ~v_25192;
assign v_28367 = v_25192;
assign v_28368 = ~v_3415;
assign v_28369 = ~v_25196;
assign v_28370 = v_25196;
assign v_28371 = ~v_25199;
assign v_28372 = ~v_3420;
assign v_28373 = v_3420;
assign v_28374 = ~v_25203;
assign v_28375 = ~v_3424;
assign v_28376 = v_3424;
assign v_28377 = ~v_25207;
assign v_28378 = ~v_3428;
assign v_28379 = v_3428;
assign v_28380 = ~v_25211;
assign v_28381 = ~v_3432;
assign v_28382 = v_3432;
assign v_28383 = ~v_25215;
assign v_28384 = ~v_3436;
assign v_28385 = v_3436;
assign v_28386 = ~v_25219;
assign v_28387 = ~v_3440;
assign v_28388 = v_3440;
assign v_28389 = ~v_25223;
assign v_28390 = ~v_3444;
assign v_28391 = v_3444;
assign v_28392 = ~v_25227;
assign v_28393 = ~v_3448;
assign v_28394 = v_3448;
assign v_28395 = ~v_25231;
assign v_28396 = ~v_3452;
assign v_28397 = v_3452;
assign v_28398 = ~v_25235;
assign v_28399 = ~v_3456;
assign v_28400 = v_3456;
assign v_28401 = ~v_25239;
assign v_28402 = ~v_3460;
assign v_28403 = v_3460;
assign v_28404 = ~v_25243;
assign v_28405 = ~v_3464;
assign v_28406 = v_3464;
assign v_28407 = ~v_25247;
assign v_28408 = ~v_3468;
assign v_28409 = v_28408;
assign v_28411 = v_28410;
assign v_28413 = v_28405 & v_28412;
assign v_28415 = v_25243;
assign v_28417 = v_28414 & v_28416;
assign v_28419 = v_28402 & v_28418;
assign v_28421 = v_25239;
assign v_28423 = v_28420 & v_28422;
assign v_28425 = v_28399 & v_28424;
assign v_28427 = v_25235;
assign v_28429 = v_28426 & v_28428;
assign v_28431 = v_28396 & v_28430;
assign v_28433 = v_25231;
assign v_28435 = v_28432 & v_28434;
assign v_28437 = v_28393 & v_28436;
assign v_28439 = v_25227;
assign v_28441 = v_28438 & v_28440;
assign v_28443 = v_28390 & v_28442;
assign v_28445 = v_25223;
assign v_28447 = v_28444 & v_28446;
assign v_28449 = v_28387 & v_28448;
assign v_28451 = v_25219;
assign v_28453 = v_28450 & v_28452;
assign v_28455 = v_28384 & v_28454;
assign v_28457 = v_25215;
assign v_28459 = v_28456 & v_28458;
assign v_28461 = v_28381 & v_28460;
assign v_28463 = v_25211;
assign v_28465 = v_28462 & v_28464;
assign v_28467 = v_28378 & v_28466;
assign v_28469 = v_25207;
assign v_28471 = v_28468 & v_28470;
assign v_28473 = v_28375 & v_28472;
assign v_28475 = v_25203;
assign v_28477 = v_28474 & v_28476;
assign v_28479 = v_28372 & v_28478;
assign v_28481 = v_25199;
assign v_28483 = v_28480 & v_28482;
assign v_28485 = v_28369 & v_28484;
assign v_28487 = v_3415;
assign v_28489 = v_28486 & v_28488;
assign v_28491 = v_28366 & v_28490;
assign v_28493 = v_3411;
assign v_28495 = v_28492 & v_28494;
assign v_28497 = v_28363 & v_28496;
assign v_28499 = v_3407;
assign v_28501 = v_28498 & v_28500;
assign v_28503 = v_28360 & v_28502;
assign v_28505 = v_3403;
assign v_28507 = v_28504 & v_28506;
assign v_28508 = v_28507;
assign v_28510 = v_25247;
assign v_28511 = v_3468;
assign v_28512 = v_28511;
assign v_28513 = v_28510 & v_28512;
assign v_28514 = v_28513;
assign v_28515 = v_28405 & v_28514;
assign v_28517 = v_28415 & v_28516;
assign v_28518 = v_28404 & v_28514;
assign v_28520 = v_28402 & v_28519;
assign v_28522 = v_28421 & v_28521;
assign v_28523 = v_28401 & v_28519;
assign v_28525 = v_28399 & v_28524;
assign v_28527 = v_28427 & v_28526;
assign v_28528 = v_28398 & v_28524;
assign v_28530 = v_28396 & v_28529;
assign v_28532 = v_28433 & v_28531;
assign v_28533 = v_28395 & v_28529;
assign v_28535 = v_28393 & v_28534;
assign v_28537 = v_28439 & v_28536;
assign v_28538 = v_28392 & v_28534;
assign v_28540 = v_28390 & v_28539;
assign v_28542 = v_28445 & v_28541;
assign v_28543 = v_28389 & v_28539;
assign v_28545 = v_28387 & v_28544;
assign v_28547 = v_28451 & v_28546;
assign v_28548 = v_28386 & v_28544;
assign v_28550 = v_28384 & v_28549;
assign v_28552 = v_28457 & v_28551;
assign v_28553 = v_28383 & v_28549;
assign v_28555 = v_28381 & v_28554;
assign v_28557 = v_28463 & v_28556;
assign v_28558 = v_28380 & v_28554;
assign v_28560 = v_28378 & v_28559;
assign v_28562 = v_28469 & v_28561;
assign v_28563 = v_28377 & v_28559;
assign v_28565 = v_28375 & v_28564;
assign v_28567 = v_28475 & v_28566;
assign v_28568 = v_28374 & v_28564;
assign v_28570 = v_28372 & v_28569;
assign v_28572 = v_28481 & v_28571;
assign v_28573 = v_28371 & v_28569;
assign v_28575 = v_28369 & v_28574;
assign v_28577 = v_28487 & v_28576;
assign v_28578 = v_28368 & v_28574;
assign v_28580 = v_28366 & v_28579;
assign v_28582 = v_28493 & v_28581;
assign v_28583 = v_28365 & v_28579;
assign v_28585 = v_28363 & v_28584;
assign v_28587 = v_28499 & v_28586;
assign v_28588 = v_28362 & v_28584;
assign v_28590 = v_28360 & v_28589;
assign v_28592 = v_28505 & v_28591;
assign v_28593 = v_28359 & v_28589;
assign v_28595 = v_28594;
assign v_28597 = v_28509 & v_28596;
assign v_28598 = v_28597;
assign v_28600 = v_28599;
assign v_28602 = ~v_3663;
assign v_28603 = ~v_25184;
assign v_28604 = v_25184;
assign v_28605 = ~v_3667;
assign v_28606 = ~v_25188;
assign v_28607 = v_25188;
assign v_28608 = ~v_3671;
assign v_28609 = ~v_25192;
assign v_28610 = v_25192;
assign v_28611 = ~v_3675;
assign v_28612 = ~v_25196;
assign v_28613 = v_25196;
assign v_28614 = ~v_25199;
assign v_28615 = ~v_3680;
assign v_28616 = v_3680;
assign v_28617 = ~v_25203;
assign v_28618 = ~v_3684;
assign v_28619 = v_3684;
assign v_28620 = ~v_25207;
assign v_28621 = ~v_3688;
assign v_28622 = v_3688;
assign v_28623 = ~v_25211;
assign v_28624 = ~v_3692;
assign v_28625 = v_3692;
assign v_28626 = ~v_25215;
assign v_28627 = ~v_3696;
assign v_28628 = v_3696;
assign v_28629 = ~v_25219;
assign v_28630 = ~v_3700;
assign v_28631 = v_3700;
assign v_28632 = ~v_25223;
assign v_28633 = ~v_3704;
assign v_28634 = v_3704;
assign v_28635 = ~v_25227;
assign v_28636 = ~v_3708;
assign v_28637 = v_3708;
assign v_28638 = ~v_25231;
assign v_28639 = ~v_3712;
assign v_28640 = v_3712;
assign v_28641 = ~v_25235;
assign v_28642 = ~v_3716;
assign v_28643 = v_3716;
assign v_28644 = ~v_25239;
assign v_28645 = ~v_3720;
assign v_28646 = v_3720;
assign v_28647 = ~v_25243;
assign v_28648 = ~v_3724;
assign v_28649 = v_3724;
assign v_28650 = ~v_25247;
assign v_28651 = ~v_3728;
assign v_28652 = v_28651;
assign v_28654 = v_28653;
assign v_28656 = v_28648 & v_28655;
assign v_28658 = v_25243;
assign v_28660 = v_28657 & v_28659;
assign v_28662 = v_28645 & v_28661;
assign v_28664 = v_25239;
assign v_28666 = v_28663 & v_28665;
assign v_28668 = v_28642 & v_28667;
assign v_28670 = v_25235;
assign v_28672 = v_28669 & v_28671;
assign v_28674 = v_28639 & v_28673;
assign v_28676 = v_25231;
assign v_28678 = v_28675 & v_28677;
assign v_28680 = v_28636 & v_28679;
assign v_28682 = v_25227;
assign v_28684 = v_28681 & v_28683;
assign v_28686 = v_28633 & v_28685;
assign v_28688 = v_25223;
assign v_28690 = v_28687 & v_28689;
assign v_28692 = v_28630 & v_28691;
assign v_28694 = v_25219;
assign v_28696 = v_28693 & v_28695;
assign v_28698 = v_28627 & v_28697;
assign v_28700 = v_25215;
assign v_28702 = v_28699 & v_28701;
assign v_28704 = v_28624 & v_28703;
assign v_28706 = v_25211;
assign v_28708 = v_28705 & v_28707;
assign v_28710 = v_28621 & v_28709;
assign v_28712 = v_25207;
assign v_28714 = v_28711 & v_28713;
assign v_28716 = v_28618 & v_28715;
assign v_28718 = v_25203;
assign v_28720 = v_28717 & v_28719;
assign v_28722 = v_28615 & v_28721;
assign v_28724 = v_25199;
assign v_28726 = v_28723 & v_28725;
assign v_28728 = v_28612 & v_28727;
assign v_28730 = v_3675;
assign v_28732 = v_28729 & v_28731;
assign v_28734 = v_28609 & v_28733;
assign v_28736 = v_3671;
assign v_28738 = v_28735 & v_28737;
assign v_28740 = v_28606 & v_28739;
assign v_28742 = v_3667;
assign v_28744 = v_28741 & v_28743;
assign v_28746 = v_28603 & v_28745;
assign v_28748 = v_3663;
assign v_28750 = v_28747 & v_28749;
assign v_28751 = v_28750;
assign v_28753 = v_25247;
assign v_28754 = v_3728;
assign v_28755 = v_28754;
assign v_28756 = v_28753 & v_28755;
assign v_28757 = v_28756;
assign v_28758 = v_28648 & v_28757;
assign v_28760 = v_28658 & v_28759;
assign v_28761 = v_28647 & v_28757;
assign v_28763 = v_28645 & v_28762;
assign v_28765 = v_28664 & v_28764;
assign v_28766 = v_28644 & v_28762;
assign v_28768 = v_28642 & v_28767;
assign v_28770 = v_28670 & v_28769;
assign v_28771 = v_28641 & v_28767;
assign v_28773 = v_28639 & v_28772;
assign v_28775 = v_28676 & v_28774;
assign v_28776 = v_28638 & v_28772;
assign v_28778 = v_28636 & v_28777;
assign v_28780 = v_28682 & v_28779;
assign v_28781 = v_28635 & v_28777;
assign v_28783 = v_28633 & v_28782;
assign v_28785 = v_28688 & v_28784;
assign v_28786 = v_28632 & v_28782;
assign v_28788 = v_28630 & v_28787;
assign v_28790 = v_28694 & v_28789;
assign v_28791 = v_28629 & v_28787;
assign v_28793 = v_28627 & v_28792;
assign v_28795 = v_28700 & v_28794;
assign v_28796 = v_28626 & v_28792;
assign v_28798 = v_28624 & v_28797;
assign v_28800 = v_28706 & v_28799;
assign v_28801 = v_28623 & v_28797;
assign v_28803 = v_28621 & v_28802;
assign v_28805 = v_28712 & v_28804;
assign v_28806 = v_28620 & v_28802;
assign v_28808 = v_28618 & v_28807;
assign v_28810 = v_28718 & v_28809;
assign v_28811 = v_28617 & v_28807;
assign v_28813 = v_28615 & v_28812;
assign v_28815 = v_28724 & v_28814;
assign v_28816 = v_28614 & v_28812;
assign v_28818 = v_28612 & v_28817;
assign v_28820 = v_28730 & v_28819;
assign v_28821 = v_28611 & v_28817;
assign v_28823 = v_28609 & v_28822;
assign v_28825 = v_28736 & v_28824;
assign v_28826 = v_28608 & v_28822;
assign v_28828 = v_28606 & v_28827;
assign v_28830 = v_28742 & v_28829;
assign v_28831 = v_28605 & v_28827;
assign v_28833 = v_28603 & v_28832;
assign v_28835 = v_28748 & v_28834;
assign v_28836 = v_28602 & v_28832;
assign v_28838 = v_28837;
assign v_28840 = v_28752 & v_28839;
assign v_28841 = v_28840;
assign v_28843 = v_28842;
assign v_28845 = ~v_3923;
assign v_28846 = ~v_25184;
assign v_28847 = v_25184;
assign v_28848 = ~v_3927;
assign v_28849 = ~v_25188;
assign v_28850 = v_25188;
assign v_28851 = ~v_3931;
assign v_28852 = ~v_25192;
assign v_28853 = v_25192;
assign v_28854 = ~v_3935;
assign v_28855 = ~v_25196;
assign v_28856 = v_25196;
assign v_28857 = ~v_25199;
assign v_28858 = ~v_3940;
assign v_28859 = v_3940;
assign v_28860 = ~v_25203;
assign v_28861 = ~v_3944;
assign v_28862 = v_3944;
assign v_28863 = ~v_25207;
assign v_28864 = ~v_3948;
assign v_28865 = v_3948;
assign v_28866 = ~v_25211;
assign v_28867 = ~v_3952;
assign v_28868 = v_3952;
assign v_28869 = ~v_25215;
assign v_28870 = ~v_3956;
assign v_28871 = v_3956;
assign v_28872 = ~v_25219;
assign v_28873 = ~v_3960;
assign v_28874 = v_3960;
assign v_28875 = ~v_25223;
assign v_28876 = ~v_3964;
assign v_28877 = v_3964;
assign v_28878 = ~v_25227;
assign v_28879 = ~v_3968;
assign v_28880 = v_3968;
assign v_28881 = ~v_25231;
assign v_28882 = ~v_3972;
assign v_28883 = v_3972;
assign v_28884 = ~v_25235;
assign v_28885 = ~v_3976;
assign v_28886 = v_3976;
assign v_28887 = ~v_25239;
assign v_28888 = ~v_3980;
assign v_28889 = v_3980;
assign v_28890 = ~v_25243;
assign v_28891 = ~v_3984;
assign v_28892 = v_3984;
assign v_28893 = ~v_25247;
assign v_28894 = ~v_3988;
assign v_28895 = v_28894;
assign v_28897 = v_28896;
assign v_28899 = v_28891 & v_28898;
assign v_28901 = v_25243;
assign v_28903 = v_28900 & v_28902;
assign v_28905 = v_28888 & v_28904;
assign v_28907 = v_25239;
assign v_28909 = v_28906 & v_28908;
assign v_28911 = v_28885 & v_28910;
assign v_28913 = v_25235;
assign v_28915 = v_28912 & v_28914;
assign v_28917 = v_28882 & v_28916;
assign v_28919 = v_25231;
assign v_28921 = v_28918 & v_28920;
assign v_28923 = v_28879 & v_28922;
assign v_28925 = v_25227;
assign v_28927 = v_28924 & v_28926;
assign v_28929 = v_28876 & v_28928;
assign v_28931 = v_25223;
assign v_28933 = v_28930 & v_28932;
assign v_28935 = v_28873 & v_28934;
assign v_28937 = v_25219;
assign v_28939 = v_28936 & v_28938;
assign v_28941 = v_28870 & v_28940;
assign v_28943 = v_25215;
assign v_28945 = v_28942 & v_28944;
assign v_28947 = v_28867 & v_28946;
assign v_28949 = v_25211;
assign v_28951 = v_28948 & v_28950;
assign v_28953 = v_28864 & v_28952;
assign v_28955 = v_25207;
assign v_28957 = v_28954 & v_28956;
assign v_28959 = v_28861 & v_28958;
assign v_28961 = v_25203;
assign v_28963 = v_28960 & v_28962;
assign v_28965 = v_28858 & v_28964;
assign v_28967 = v_25199;
assign v_28969 = v_28966 & v_28968;
assign v_28971 = v_28855 & v_28970;
assign v_28973 = v_3935;
assign v_28975 = v_28972 & v_28974;
assign v_28977 = v_28852 & v_28976;
assign v_28979 = v_3931;
assign v_28981 = v_28978 & v_28980;
assign v_28983 = v_28849 & v_28982;
assign v_28985 = v_3927;
assign v_28987 = v_28984 & v_28986;
assign v_28989 = v_28846 & v_28988;
assign v_28991 = v_3923;
assign v_28993 = v_28990 & v_28992;
assign v_28994 = v_28993;
assign v_28996 = v_25247;
assign v_28997 = v_3988;
assign v_28998 = v_28997;
assign v_28999 = v_28996 & v_28998;
assign v_29000 = v_28999;
assign v_29001 = v_28891 & v_29000;
assign v_29003 = v_28901 & v_29002;
assign v_29004 = v_28890 & v_29000;
assign v_29006 = v_28888 & v_29005;
assign v_29008 = v_28907 & v_29007;
assign v_29009 = v_28887 & v_29005;
assign v_29011 = v_28885 & v_29010;
assign v_29013 = v_28913 & v_29012;
assign v_29014 = v_28884 & v_29010;
assign v_29016 = v_28882 & v_29015;
assign v_29018 = v_28919 & v_29017;
assign v_29019 = v_28881 & v_29015;
assign v_29021 = v_28879 & v_29020;
assign v_29023 = v_28925 & v_29022;
assign v_29024 = v_28878 & v_29020;
assign v_29026 = v_28876 & v_29025;
assign v_29028 = v_28931 & v_29027;
assign v_29029 = v_28875 & v_29025;
assign v_29031 = v_28873 & v_29030;
assign v_29033 = v_28937 & v_29032;
assign v_29034 = v_28872 & v_29030;
assign v_29036 = v_28870 & v_29035;
assign v_29038 = v_28943 & v_29037;
assign v_29039 = v_28869 & v_29035;
assign v_29041 = v_28867 & v_29040;
assign v_29043 = v_28949 & v_29042;
assign v_29044 = v_28866 & v_29040;
assign v_29046 = v_28864 & v_29045;
assign v_29048 = v_28955 & v_29047;
assign v_29049 = v_28863 & v_29045;
assign v_29051 = v_28861 & v_29050;
assign v_29053 = v_28961 & v_29052;
assign v_29054 = v_28860 & v_29050;
assign v_29056 = v_28858 & v_29055;
assign v_29058 = v_28967 & v_29057;
assign v_29059 = v_28857 & v_29055;
assign v_29061 = v_28855 & v_29060;
assign v_29063 = v_28973 & v_29062;
assign v_29064 = v_28854 & v_29060;
assign v_29066 = v_28852 & v_29065;
assign v_29068 = v_28979 & v_29067;
assign v_29069 = v_28851 & v_29065;
assign v_29071 = v_28849 & v_29070;
assign v_29073 = v_28985 & v_29072;
assign v_29074 = v_28848 & v_29070;
assign v_29076 = v_28846 & v_29075;
assign v_29078 = v_28991 & v_29077;
assign v_29079 = v_28845 & v_29075;
assign v_29081 = v_29080;
assign v_29083 = v_28995 & v_29082;
assign v_29084 = v_29083;
assign v_29086 = v_29085;
assign v_29087 = ~v_4182;
assign v_29088 = ~v_25184;
assign v_29089 = v_25184;
assign v_29090 = ~v_4186;
assign v_29091 = ~v_25188;
assign v_29092 = v_25188;
assign v_29093 = ~v_4190;
assign v_29094 = ~v_25192;
assign v_29095 = v_25192;
assign v_29096 = ~v_4194;
assign v_29097 = ~v_25196;
assign v_29098 = v_25196;
assign v_29099 = ~v_25199;
assign v_29100 = ~v_4199;
assign v_29101 = v_4199;
assign v_29102 = ~v_25203;
assign v_29103 = ~v_4203;
assign v_29104 = v_4203;
assign v_29105 = ~v_25207;
assign v_29106 = ~v_4207;
assign v_29107 = v_4207;
assign v_29108 = ~v_25211;
assign v_29109 = ~v_4211;
assign v_29110 = v_4211;
assign v_29111 = ~v_25215;
assign v_29112 = ~v_4215;
assign v_29113 = v_4215;
assign v_29114 = ~v_25219;
assign v_29115 = ~v_4219;
assign v_29116 = v_4219;
assign v_29117 = ~v_25223;
assign v_29118 = ~v_4223;
assign v_29119 = v_4223;
assign v_29120 = ~v_25227;
assign v_29121 = ~v_4227;
assign v_29122 = v_4227;
assign v_29123 = ~v_25231;
assign v_29124 = ~v_4231;
assign v_29125 = v_4231;
assign v_29126 = ~v_25235;
assign v_29127 = ~v_4235;
assign v_29128 = v_4235;
assign v_29129 = ~v_25239;
assign v_29130 = ~v_4239;
assign v_29131 = v_4239;
assign v_29132 = ~v_25243;
assign v_29133 = ~v_4243;
assign v_29134 = v_4243;
assign v_29135 = ~v_25247;
assign v_29136 = ~v_4247;
assign v_29137 = v_29136;
assign v_29139 = v_29138;
assign v_29141 = v_29133 & v_29140;
assign v_29143 = v_25243;
assign v_29145 = v_29142 & v_29144;
assign v_29147 = v_29130 & v_29146;
assign v_29149 = v_25239;
assign v_29151 = v_29148 & v_29150;
assign v_29153 = v_29127 & v_29152;
assign v_29155 = v_25235;
assign v_29157 = v_29154 & v_29156;
assign v_29159 = v_29124 & v_29158;
assign v_29161 = v_25231;
assign v_29163 = v_29160 & v_29162;
assign v_29165 = v_29121 & v_29164;
assign v_29167 = v_25227;
assign v_29169 = v_29166 & v_29168;
assign v_29171 = v_29118 & v_29170;
assign v_29173 = v_25223;
assign v_29175 = v_29172 & v_29174;
assign v_29177 = v_29115 & v_29176;
assign v_29179 = v_25219;
assign v_29181 = v_29178 & v_29180;
assign v_29183 = v_29112 & v_29182;
assign v_29185 = v_25215;
assign v_29187 = v_29184 & v_29186;
assign v_29189 = v_29109 & v_29188;
assign v_29191 = v_25211;
assign v_29193 = v_29190 & v_29192;
assign v_29195 = v_29106 & v_29194;
assign v_29197 = v_25207;
assign v_29199 = v_29196 & v_29198;
assign v_29201 = v_29103 & v_29200;
assign v_29203 = v_25203;
assign v_29205 = v_29202 & v_29204;
assign v_29207 = v_29100 & v_29206;
assign v_29209 = v_25199;
assign v_29211 = v_29208 & v_29210;
assign v_29213 = v_29097 & v_29212;
assign v_29215 = v_4194;
assign v_29217 = v_29214 & v_29216;
assign v_29219 = v_29094 & v_29218;
assign v_29221 = v_4190;
assign v_29223 = v_29220 & v_29222;
assign v_29225 = v_29091 & v_29224;
assign v_29227 = v_4186;
assign v_29229 = v_29226 & v_29228;
assign v_29231 = v_29088 & v_29230;
assign v_29233 = v_4182;
assign v_29235 = v_29232 & v_29234;
assign v_29237 = ~v_29236;
assign v_29239 = v_25247;
assign v_29240 = v_4247;
assign v_29241 = v_29240;
assign v_29242 = v_29239 & v_29241;
assign v_29243 = v_29242;
assign v_29244 = v_29133 & v_29243;
assign v_29246 = v_29143 & v_29245;
assign v_29247 = v_29132 & v_29243;
assign v_29249 = v_29130 & v_29248;
assign v_29251 = v_29149 & v_29250;
assign v_29252 = v_29129 & v_29248;
assign v_29254 = v_29127 & v_29253;
assign v_29256 = v_29155 & v_29255;
assign v_29257 = v_29126 & v_29253;
assign v_29259 = v_29124 & v_29258;
assign v_29261 = v_29161 & v_29260;
assign v_29262 = v_29123 & v_29258;
assign v_29264 = v_29121 & v_29263;
assign v_29266 = v_29167 & v_29265;
assign v_29267 = v_29120 & v_29263;
assign v_29269 = v_29118 & v_29268;
assign v_29271 = v_29173 & v_29270;
assign v_29272 = v_29117 & v_29268;
assign v_29274 = v_29115 & v_29273;
assign v_29276 = v_29179 & v_29275;
assign v_29277 = v_29114 & v_29273;
assign v_29279 = v_29112 & v_29278;
assign v_29281 = v_29185 & v_29280;
assign v_29282 = v_29111 & v_29278;
assign v_29284 = v_29109 & v_29283;
assign v_29286 = v_29191 & v_29285;
assign v_29287 = v_29108 & v_29283;
assign v_29289 = v_29106 & v_29288;
assign v_29291 = v_29197 & v_29290;
assign v_29292 = v_29105 & v_29288;
assign v_29294 = v_29103 & v_29293;
assign v_29296 = v_29203 & v_29295;
assign v_29297 = v_29102 & v_29293;
assign v_29299 = v_29100 & v_29298;
assign v_29301 = v_29209 & v_29300;
assign v_29302 = v_29099 & v_29298;
assign v_29304 = v_29097 & v_29303;
assign v_29306 = v_29215 & v_29305;
assign v_29307 = v_29096 & v_29303;
assign v_29309 = v_29094 & v_29308;
assign v_29311 = v_29221 & v_29310;
assign v_29312 = v_29093 & v_29308;
assign v_29314 = v_29091 & v_29313;
assign v_29316 = v_29227 & v_29315;
assign v_29317 = v_29090 & v_29313;
assign v_29319 = v_29088 & v_29318;
assign v_29321 = v_29233 & v_29320;
assign v_29322 = v_29087 & v_29318;
assign v_29324 = v_29236;
assign v_29326 = v_29238 & v_29325;
assign v_29327 = v_29326;
assign v_29329 = v_29328;
assign v_29331 = ~v_6;
assign v_29333 = ~v_29332;
assign v_29334 = v_29332;
assign v_29335 = ~v_13;
assign v_29337 = ~v_29336;
assign v_29338 = v_29336;
assign v_29339 = ~v_18;
assign v_29341 = ~v_29340;
assign v_29342 = v_29340;
assign v_29343 = ~v_23;
assign v_29345 = ~v_29344;
assign v_29346 = v_29344;
assign v_29348 = ~v_29347;
assign v_29349 = ~v_30;
assign v_29350 = v_30;
assign v_29352 = ~v_29351;
assign v_29353 = ~v_35;
assign v_29354 = v_35;
assign v_29356 = ~v_29355;
assign v_29357 = ~v_40;
assign v_29358 = v_40;
assign v_29360 = ~v_29359;
assign v_29361 = ~v_45;
assign v_29362 = v_45;
assign v_29364 = ~v_29363;
assign v_29365 = ~v_50;
assign v_29366 = v_50;
assign v_29368 = ~v_29367;
assign v_29369 = ~v_55;
assign v_29370 = v_55;
assign v_29372 = ~v_29371;
assign v_29373 = ~v_60;
assign v_29374 = v_60;
assign v_29376 = ~v_29375;
assign v_29377 = ~v_65;
assign v_29378 = v_65;
assign v_29380 = ~v_29379;
assign v_29381 = ~v_70;
assign v_29382 = v_70;
assign v_29384 = ~v_29383;
assign v_29385 = ~v_75;
assign v_29386 = v_75;
assign v_29388 = ~v_29387;
assign v_29389 = ~v_80;
assign v_29390 = v_80;
assign v_29392 = ~v_29391;
assign v_29393 = ~v_85;
assign v_29394 = v_85;
assign v_29396 = ~v_29395;
assign v_29397 = ~v_90;
assign v_29398 = v_29397;
assign v_29400 = v_29399;
assign v_29402 = v_29393 & v_29401;
assign v_29404 = v_29391;
assign v_29406 = v_29403 & v_29405;
assign v_29408 = v_29389 & v_29407;
assign v_29410 = v_29387;
assign v_29412 = v_29409 & v_29411;
assign v_29414 = v_29385 & v_29413;
assign v_29416 = v_29383;
assign v_29418 = v_29415 & v_29417;
assign v_29420 = v_29381 & v_29419;
assign v_29422 = v_29379;
assign v_29424 = v_29421 & v_29423;
assign v_29426 = v_29377 & v_29425;
assign v_29428 = v_29375;
assign v_29430 = v_29427 & v_29429;
assign v_29432 = v_29373 & v_29431;
assign v_29434 = v_29371;
assign v_29436 = v_29433 & v_29435;
assign v_29438 = v_29369 & v_29437;
assign v_29440 = v_29367;
assign v_29442 = v_29439 & v_29441;
assign v_29444 = v_29365 & v_29443;
assign v_29446 = v_29363;
assign v_29448 = v_29445 & v_29447;
assign v_29450 = v_29361 & v_29449;
assign v_29452 = v_29359;
assign v_29454 = v_29451 & v_29453;
assign v_29456 = v_29357 & v_29455;
assign v_29458 = v_29355;
assign v_29460 = v_29457 & v_29459;
assign v_29462 = v_29353 & v_29461;
assign v_29464 = v_29351;
assign v_29466 = v_29463 & v_29465;
assign v_29468 = v_29349 & v_29467;
assign v_29470 = v_29347;
assign v_29472 = v_29469 & v_29471;
assign v_29474 = v_29345 & v_29473;
assign v_29476 = v_23;
assign v_29478 = v_29475 & v_29477;
assign v_29480 = v_29341 & v_29479;
assign v_29482 = v_18;
assign v_29484 = v_29481 & v_29483;
assign v_29486 = v_29337 & v_29485;
assign v_29488 = v_13;
assign v_29490 = v_29487 & v_29489;
assign v_29492 = v_29333 & v_29491;
assign v_29494 = v_6;
assign v_29496 = v_29493 & v_29495;
assign v_29497 = v_29496;
assign v_29499 = v_29395;
assign v_29500 = v_90;
assign v_29501 = v_29500;
assign v_29502 = v_29499 & v_29501;
assign v_29503 = v_29502;
assign v_29504 = v_29393 & v_29503;
assign v_29506 = v_29404 & v_29505;
assign v_29507 = v_29392 & v_29503;
assign v_29509 = v_29389 & v_29508;
assign v_29511 = v_29410 & v_29510;
assign v_29512 = v_29388 & v_29508;
assign v_29514 = v_29385 & v_29513;
assign v_29516 = v_29416 & v_29515;
assign v_29517 = v_29384 & v_29513;
assign v_29519 = v_29381 & v_29518;
assign v_29521 = v_29422 & v_29520;
assign v_29522 = v_29380 & v_29518;
assign v_29524 = v_29377 & v_29523;
assign v_29526 = v_29428 & v_29525;
assign v_29527 = v_29376 & v_29523;
assign v_29529 = v_29373 & v_29528;
assign v_29531 = v_29434 & v_29530;
assign v_29532 = v_29372 & v_29528;
assign v_29534 = v_29369 & v_29533;
assign v_29536 = v_29440 & v_29535;
assign v_29537 = v_29368 & v_29533;
assign v_29539 = v_29365 & v_29538;
assign v_29541 = v_29446 & v_29540;
assign v_29542 = v_29364 & v_29538;
assign v_29544 = v_29361 & v_29543;
assign v_29546 = v_29452 & v_29545;
assign v_29547 = v_29360 & v_29543;
assign v_29549 = v_29357 & v_29548;
assign v_29551 = v_29458 & v_29550;
assign v_29552 = v_29356 & v_29548;
assign v_29554 = v_29353 & v_29553;
assign v_29556 = v_29464 & v_29555;
assign v_29557 = v_29352 & v_29553;
assign v_29559 = v_29349 & v_29558;
assign v_29561 = v_29470 & v_29560;
assign v_29562 = v_29348 & v_29558;
assign v_29564 = v_29345 & v_29563;
assign v_29566 = v_29476 & v_29565;
assign v_29567 = v_29343 & v_29563;
assign v_29569 = v_29341 & v_29568;
assign v_29571 = v_29482 & v_29570;
assign v_29572 = v_29339 & v_29568;
assign v_29574 = v_29337 & v_29573;
assign v_29576 = v_29488 & v_29575;
assign v_29577 = v_29335 & v_29573;
assign v_29579 = v_29333 & v_29578;
assign v_29581 = v_29494 & v_29580;
assign v_29582 = v_29331 & v_29578;
assign v_29584 = v_29583;
assign v_29586 = v_29498 & v_29585;
assign v_29587 = v_29586;
assign v_29589 = v_29588;
assign v_29591 = ~v_283;
assign v_29592 = ~v_29332;
assign v_29593 = v_29332;
assign v_29594 = ~v_287;
assign v_29595 = ~v_29336;
assign v_29596 = v_29336;
assign v_29597 = ~v_291;
assign v_29598 = ~v_29340;
assign v_29599 = v_29340;
assign v_29600 = ~v_295;
assign v_29601 = ~v_29344;
assign v_29602 = v_29344;
assign v_29603 = ~v_29347;
assign v_29604 = ~v_300;
assign v_29605 = v_300;
assign v_29606 = ~v_29351;
assign v_29607 = ~v_304;
assign v_29608 = v_304;
assign v_29609 = ~v_29355;
assign v_29610 = ~v_308;
assign v_29611 = v_308;
assign v_29612 = ~v_29359;
assign v_29613 = ~v_312;
assign v_29614 = v_312;
assign v_29615 = ~v_29363;
assign v_29616 = ~v_316;
assign v_29617 = v_316;
assign v_29618 = ~v_29367;
assign v_29619 = ~v_320;
assign v_29620 = v_320;
assign v_29621 = ~v_29371;
assign v_29622 = ~v_324;
assign v_29623 = v_324;
assign v_29624 = ~v_29375;
assign v_29625 = ~v_328;
assign v_29626 = v_328;
assign v_29627 = ~v_29379;
assign v_29628 = ~v_332;
assign v_29629 = v_332;
assign v_29630 = ~v_29383;
assign v_29631 = ~v_336;
assign v_29632 = v_336;
assign v_29633 = ~v_29387;
assign v_29634 = ~v_340;
assign v_29635 = v_340;
assign v_29636 = ~v_29391;
assign v_29637 = ~v_344;
assign v_29638 = v_344;
assign v_29639 = ~v_29395;
assign v_29640 = ~v_348;
assign v_29641 = v_29640;
assign v_29643 = v_29642;
assign v_29645 = v_29637 & v_29644;
assign v_29647 = v_29391;
assign v_29649 = v_29646 & v_29648;
assign v_29651 = v_29634 & v_29650;
assign v_29653 = v_29387;
assign v_29655 = v_29652 & v_29654;
assign v_29657 = v_29631 & v_29656;
assign v_29659 = v_29383;
assign v_29661 = v_29658 & v_29660;
assign v_29663 = v_29628 & v_29662;
assign v_29665 = v_29379;
assign v_29667 = v_29664 & v_29666;
assign v_29669 = v_29625 & v_29668;
assign v_29671 = v_29375;
assign v_29673 = v_29670 & v_29672;
assign v_29675 = v_29622 & v_29674;
assign v_29677 = v_29371;
assign v_29679 = v_29676 & v_29678;
assign v_29681 = v_29619 & v_29680;
assign v_29683 = v_29367;
assign v_29685 = v_29682 & v_29684;
assign v_29687 = v_29616 & v_29686;
assign v_29689 = v_29363;
assign v_29691 = v_29688 & v_29690;
assign v_29693 = v_29613 & v_29692;
assign v_29695 = v_29359;
assign v_29697 = v_29694 & v_29696;
assign v_29699 = v_29610 & v_29698;
assign v_29701 = v_29355;
assign v_29703 = v_29700 & v_29702;
assign v_29705 = v_29607 & v_29704;
assign v_29707 = v_29351;
assign v_29709 = v_29706 & v_29708;
assign v_29711 = v_29604 & v_29710;
assign v_29713 = v_29347;
assign v_29715 = v_29712 & v_29714;
assign v_29717 = v_29601 & v_29716;
assign v_29719 = v_295;
assign v_29721 = v_29718 & v_29720;
assign v_29723 = v_29598 & v_29722;
assign v_29725 = v_291;
assign v_29727 = v_29724 & v_29726;
assign v_29729 = v_29595 & v_29728;
assign v_29731 = v_287;
assign v_29733 = v_29730 & v_29732;
assign v_29735 = v_29592 & v_29734;
assign v_29737 = v_283;
assign v_29739 = v_29736 & v_29738;
assign v_29740 = v_29739;
assign v_29742 = v_29395;
assign v_29743 = v_348;
assign v_29744 = v_29743;
assign v_29745 = v_29742 & v_29744;
assign v_29746 = v_29745;
assign v_29747 = v_29637 & v_29746;
assign v_29749 = v_29647 & v_29748;
assign v_29750 = v_29636 & v_29746;
assign v_29752 = v_29634 & v_29751;
assign v_29754 = v_29653 & v_29753;
assign v_29755 = v_29633 & v_29751;
assign v_29757 = v_29631 & v_29756;
assign v_29759 = v_29659 & v_29758;
assign v_29760 = v_29630 & v_29756;
assign v_29762 = v_29628 & v_29761;
assign v_29764 = v_29665 & v_29763;
assign v_29765 = v_29627 & v_29761;
assign v_29767 = v_29625 & v_29766;
assign v_29769 = v_29671 & v_29768;
assign v_29770 = v_29624 & v_29766;
assign v_29772 = v_29622 & v_29771;
assign v_29774 = v_29677 & v_29773;
assign v_29775 = v_29621 & v_29771;
assign v_29777 = v_29619 & v_29776;
assign v_29779 = v_29683 & v_29778;
assign v_29780 = v_29618 & v_29776;
assign v_29782 = v_29616 & v_29781;
assign v_29784 = v_29689 & v_29783;
assign v_29785 = v_29615 & v_29781;
assign v_29787 = v_29613 & v_29786;
assign v_29789 = v_29695 & v_29788;
assign v_29790 = v_29612 & v_29786;
assign v_29792 = v_29610 & v_29791;
assign v_29794 = v_29701 & v_29793;
assign v_29795 = v_29609 & v_29791;
assign v_29797 = v_29607 & v_29796;
assign v_29799 = v_29707 & v_29798;
assign v_29800 = v_29606 & v_29796;
assign v_29802 = v_29604 & v_29801;
assign v_29804 = v_29713 & v_29803;
assign v_29805 = v_29603 & v_29801;
assign v_29807 = v_29601 & v_29806;
assign v_29809 = v_29719 & v_29808;
assign v_29810 = v_29600 & v_29806;
assign v_29812 = v_29598 & v_29811;
assign v_29814 = v_29725 & v_29813;
assign v_29815 = v_29597 & v_29811;
assign v_29817 = v_29595 & v_29816;
assign v_29819 = v_29731 & v_29818;
assign v_29820 = v_29594 & v_29816;
assign v_29822 = v_29592 & v_29821;
assign v_29824 = v_29737 & v_29823;
assign v_29825 = v_29591 & v_29821;
assign v_29827 = v_29826;
assign v_29829 = v_29741 & v_29828;
assign v_29830 = v_29829;
assign v_29832 = v_29831;
assign v_29834 = ~v_543;
assign v_29835 = ~v_29332;
assign v_29836 = v_29332;
assign v_29837 = ~v_547;
assign v_29838 = ~v_29336;
assign v_29839 = v_29336;
assign v_29840 = ~v_551;
assign v_29841 = ~v_29340;
assign v_29842 = v_29340;
assign v_29843 = ~v_555;
assign v_29844 = ~v_29344;
assign v_29845 = v_29344;
assign v_29846 = ~v_29347;
assign v_29847 = ~v_560;
assign v_29848 = v_560;
assign v_29849 = ~v_29351;
assign v_29850 = ~v_564;
assign v_29851 = v_564;
assign v_29852 = ~v_29355;
assign v_29853 = ~v_568;
assign v_29854 = v_568;
assign v_29855 = ~v_29359;
assign v_29856 = ~v_572;
assign v_29857 = v_572;
assign v_29858 = ~v_29363;
assign v_29859 = ~v_576;
assign v_29860 = v_576;
assign v_29861 = ~v_29367;
assign v_29862 = ~v_580;
assign v_29863 = v_580;
assign v_29864 = ~v_29371;
assign v_29865 = ~v_584;
assign v_29866 = v_584;
assign v_29867 = ~v_29375;
assign v_29868 = ~v_588;
assign v_29869 = v_588;
assign v_29870 = ~v_29379;
assign v_29871 = ~v_592;
assign v_29872 = v_592;
assign v_29873 = ~v_29383;
assign v_29874 = ~v_596;
assign v_29875 = v_596;
assign v_29876 = ~v_29387;
assign v_29877 = ~v_600;
assign v_29878 = v_600;
assign v_29879 = ~v_29391;
assign v_29880 = ~v_604;
assign v_29881 = v_604;
assign v_29882 = ~v_29395;
assign v_29883 = ~v_608;
assign v_29884 = v_29883;
assign v_29886 = v_29885;
assign v_29888 = v_29880 & v_29887;
assign v_29890 = v_29391;
assign v_29892 = v_29889 & v_29891;
assign v_29894 = v_29877 & v_29893;
assign v_29896 = v_29387;
assign v_29898 = v_29895 & v_29897;
assign v_29900 = v_29874 & v_29899;
assign v_29902 = v_29383;
assign v_29904 = v_29901 & v_29903;
assign v_29906 = v_29871 & v_29905;
assign v_29908 = v_29379;
assign v_29910 = v_29907 & v_29909;
assign v_29912 = v_29868 & v_29911;
assign v_29914 = v_29375;
assign v_29916 = v_29913 & v_29915;
assign v_29918 = v_29865 & v_29917;
assign v_29920 = v_29371;
assign v_29922 = v_29919 & v_29921;
assign v_29924 = v_29862 & v_29923;
assign v_29926 = v_29367;
assign v_29928 = v_29925 & v_29927;
assign v_29930 = v_29859 & v_29929;
assign v_29932 = v_29363;
assign v_29934 = v_29931 & v_29933;
assign v_29936 = v_29856 & v_29935;
assign v_29938 = v_29359;
assign v_29940 = v_29937 & v_29939;
assign v_29942 = v_29853 & v_29941;
assign v_29944 = v_29355;
assign v_29946 = v_29943 & v_29945;
assign v_29948 = v_29850 & v_29947;
assign v_29950 = v_29351;
assign v_29952 = v_29949 & v_29951;
assign v_29954 = v_29847 & v_29953;
assign v_29956 = v_29347;
assign v_29958 = v_29955 & v_29957;
assign v_29960 = v_29844 & v_29959;
assign v_29962 = v_555;
assign v_29964 = v_29961 & v_29963;
assign v_29966 = v_29841 & v_29965;
assign v_29968 = v_551;
assign v_29970 = v_29967 & v_29969;
assign v_29972 = v_29838 & v_29971;
assign v_29974 = v_547;
assign v_29976 = v_29973 & v_29975;
assign v_29978 = v_29835 & v_29977;
assign v_29980 = v_543;
assign v_29982 = v_29979 & v_29981;
assign v_29983 = v_29982;
assign v_29985 = v_29395;
assign v_29986 = v_608;
assign v_29987 = v_29986;
assign v_29988 = v_29985 & v_29987;
assign v_29989 = v_29988;
assign v_29990 = v_29880 & v_29989;
assign v_29992 = v_29890 & v_29991;
assign v_29993 = v_29879 & v_29989;
assign v_29995 = v_29877 & v_29994;
assign v_29997 = v_29896 & v_29996;
assign v_29998 = v_29876 & v_29994;
assign v_30000 = v_29874 & v_29999;
assign v_30002 = v_29902 & v_30001;
assign v_30003 = v_29873 & v_29999;
assign v_30005 = v_29871 & v_30004;
assign v_30007 = v_29908 & v_30006;
assign v_30008 = v_29870 & v_30004;
assign v_30010 = v_29868 & v_30009;
assign v_30012 = v_29914 & v_30011;
assign v_30013 = v_29867 & v_30009;
assign v_30015 = v_29865 & v_30014;
assign v_30017 = v_29920 & v_30016;
assign v_30018 = v_29864 & v_30014;
assign v_30020 = v_29862 & v_30019;
assign v_30022 = v_29926 & v_30021;
assign v_30023 = v_29861 & v_30019;
assign v_30025 = v_29859 & v_30024;
assign v_30027 = v_29932 & v_30026;
assign v_30028 = v_29858 & v_30024;
assign v_30030 = v_29856 & v_30029;
assign v_30032 = v_29938 & v_30031;
assign v_30033 = v_29855 & v_30029;
assign v_30035 = v_29853 & v_30034;
assign v_30037 = v_29944 & v_30036;
assign v_30038 = v_29852 & v_30034;
assign v_30040 = v_29850 & v_30039;
assign v_30042 = v_29950 & v_30041;
assign v_30043 = v_29849 & v_30039;
assign v_30045 = v_29847 & v_30044;
assign v_30047 = v_29956 & v_30046;
assign v_30048 = v_29846 & v_30044;
assign v_30050 = v_29844 & v_30049;
assign v_30052 = v_29962 & v_30051;
assign v_30053 = v_29843 & v_30049;
assign v_30055 = v_29841 & v_30054;
assign v_30057 = v_29968 & v_30056;
assign v_30058 = v_29840 & v_30054;
assign v_30060 = v_29838 & v_30059;
assign v_30062 = v_29974 & v_30061;
assign v_30063 = v_29837 & v_30059;
assign v_30065 = v_29835 & v_30064;
assign v_30067 = v_29980 & v_30066;
assign v_30068 = v_29834 & v_30064;
assign v_30070 = v_30069;
assign v_30072 = v_29984 & v_30071;
assign v_30073 = v_30072;
assign v_30075 = v_30074;
assign v_30077 = ~v_803;
assign v_30078 = ~v_29332;
assign v_30079 = v_29332;
assign v_30080 = ~v_807;
assign v_30081 = ~v_29336;
assign v_30082 = v_29336;
assign v_30083 = ~v_811;
assign v_30084 = ~v_29340;
assign v_30085 = v_29340;
assign v_30086 = ~v_815;
assign v_30087 = ~v_29344;
assign v_30088 = v_29344;
assign v_30089 = ~v_29347;
assign v_30090 = ~v_820;
assign v_30091 = v_820;
assign v_30092 = ~v_29351;
assign v_30093 = ~v_824;
assign v_30094 = v_824;
assign v_30095 = ~v_29355;
assign v_30096 = ~v_828;
assign v_30097 = v_828;
assign v_30098 = ~v_29359;
assign v_30099 = ~v_832;
assign v_30100 = v_832;
assign v_30101 = ~v_29363;
assign v_30102 = ~v_836;
assign v_30103 = v_836;
assign v_30104 = ~v_29367;
assign v_30105 = ~v_840;
assign v_30106 = v_840;
assign v_30107 = ~v_29371;
assign v_30108 = ~v_844;
assign v_30109 = v_844;
assign v_30110 = ~v_29375;
assign v_30111 = ~v_848;
assign v_30112 = v_848;
assign v_30113 = ~v_29379;
assign v_30114 = ~v_852;
assign v_30115 = v_852;
assign v_30116 = ~v_29383;
assign v_30117 = ~v_856;
assign v_30118 = v_856;
assign v_30119 = ~v_29387;
assign v_30120 = ~v_860;
assign v_30121 = v_860;
assign v_30122 = ~v_29391;
assign v_30123 = ~v_864;
assign v_30124 = v_864;
assign v_30125 = ~v_29395;
assign v_30126 = ~v_868;
assign v_30127 = v_30126;
assign v_30129 = v_30128;
assign v_30131 = v_30123 & v_30130;
assign v_30133 = v_29391;
assign v_30135 = v_30132 & v_30134;
assign v_30137 = v_30120 & v_30136;
assign v_30139 = v_29387;
assign v_30141 = v_30138 & v_30140;
assign v_30143 = v_30117 & v_30142;
assign v_30145 = v_29383;
assign v_30147 = v_30144 & v_30146;
assign v_30149 = v_30114 & v_30148;
assign v_30151 = v_29379;
assign v_30153 = v_30150 & v_30152;
assign v_30155 = v_30111 & v_30154;
assign v_30157 = v_29375;
assign v_30159 = v_30156 & v_30158;
assign v_30161 = v_30108 & v_30160;
assign v_30163 = v_29371;
assign v_30165 = v_30162 & v_30164;
assign v_30167 = v_30105 & v_30166;
assign v_30169 = v_29367;
assign v_30171 = v_30168 & v_30170;
assign v_30173 = v_30102 & v_30172;
assign v_30175 = v_29363;
assign v_30177 = v_30174 & v_30176;
assign v_30179 = v_30099 & v_30178;
assign v_30181 = v_29359;
assign v_30183 = v_30180 & v_30182;
assign v_30185 = v_30096 & v_30184;
assign v_30187 = v_29355;
assign v_30189 = v_30186 & v_30188;
assign v_30191 = v_30093 & v_30190;
assign v_30193 = v_29351;
assign v_30195 = v_30192 & v_30194;
assign v_30197 = v_30090 & v_30196;
assign v_30199 = v_29347;
assign v_30201 = v_30198 & v_30200;
assign v_30203 = v_30087 & v_30202;
assign v_30205 = v_815;
assign v_30207 = v_30204 & v_30206;
assign v_30209 = v_30084 & v_30208;
assign v_30211 = v_811;
assign v_30213 = v_30210 & v_30212;
assign v_30215 = v_30081 & v_30214;
assign v_30217 = v_807;
assign v_30219 = v_30216 & v_30218;
assign v_30221 = v_30078 & v_30220;
assign v_30223 = v_803;
assign v_30225 = v_30222 & v_30224;
assign v_30226 = v_30225;
assign v_30228 = v_29395;
assign v_30229 = v_868;
assign v_30230 = v_30229;
assign v_30231 = v_30228 & v_30230;
assign v_30232 = v_30231;
assign v_30233 = v_30123 & v_30232;
assign v_30235 = v_30133 & v_30234;
assign v_30236 = v_30122 & v_30232;
assign v_30238 = v_30120 & v_30237;
assign v_30240 = v_30139 & v_30239;
assign v_30241 = v_30119 & v_30237;
assign v_30243 = v_30117 & v_30242;
assign v_30245 = v_30145 & v_30244;
assign v_30246 = v_30116 & v_30242;
assign v_30248 = v_30114 & v_30247;
assign v_30250 = v_30151 & v_30249;
assign v_30251 = v_30113 & v_30247;
assign v_30253 = v_30111 & v_30252;
assign v_30255 = v_30157 & v_30254;
assign v_30256 = v_30110 & v_30252;
assign v_30258 = v_30108 & v_30257;
assign v_30260 = v_30163 & v_30259;
assign v_30261 = v_30107 & v_30257;
assign v_30263 = v_30105 & v_30262;
assign v_30265 = v_30169 & v_30264;
assign v_30266 = v_30104 & v_30262;
assign v_30268 = v_30102 & v_30267;
assign v_30270 = v_30175 & v_30269;
assign v_30271 = v_30101 & v_30267;
assign v_30273 = v_30099 & v_30272;
assign v_30275 = v_30181 & v_30274;
assign v_30276 = v_30098 & v_30272;
assign v_30278 = v_30096 & v_30277;
assign v_30280 = v_30187 & v_30279;
assign v_30281 = v_30095 & v_30277;
assign v_30283 = v_30093 & v_30282;
assign v_30285 = v_30193 & v_30284;
assign v_30286 = v_30092 & v_30282;
assign v_30288 = v_30090 & v_30287;
assign v_30290 = v_30199 & v_30289;
assign v_30291 = v_30089 & v_30287;
assign v_30293 = v_30087 & v_30292;
assign v_30295 = v_30205 & v_30294;
assign v_30296 = v_30086 & v_30292;
assign v_30298 = v_30084 & v_30297;
assign v_30300 = v_30211 & v_30299;
assign v_30301 = v_30083 & v_30297;
assign v_30303 = v_30081 & v_30302;
assign v_30305 = v_30217 & v_30304;
assign v_30306 = v_30080 & v_30302;
assign v_30308 = v_30078 & v_30307;
assign v_30310 = v_30223 & v_30309;
assign v_30311 = v_30077 & v_30307;
assign v_30313 = v_30312;
assign v_30315 = v_30227 & v_30314;
assign v_30316 = v_30315;
assign v_30318 = v_30317;
assign v_30320 = ~v_1063;
assign v_30321 = ~v_29332;
assign v_30322 = v_29332;
assign v_30323 = ~v_1067;
assign v_30324 = ~v_29336;
assign v_30325 = v_29336;
assign v_30326 = ~v_1071;
assign v_30327 = ~v_29340;
assign v_30328 = v_29340;
assign v_30329 = ~v_1075;
assign v_30330 = ~v_29344;
assign v_30331 = v_29344;
assign v_30332 = ~v_29347;
assign v_30333 = ~v_1080;
assign v_30334 = v_1080;
assign v_30335 = ~v_29351;
assign v_30336 = ~v_1084;
assign v_30337 = v_1084;
assign v_30338 = ~v_29355;
assign v_30339 = ~v_1088;
assign v_30340 = v_1088;
assign v_30341 = ~v_29359;
assign v_30342 = ~v_1092;
assign v_30343 = v_1092;
assign v_30344 = ~v_29363;
assign v_30345 = ~v_1096;
assign v_30346 = v_1096;
assign v_30347 = ~v_29367;
assign v_30348 = ~v_1100;
assign v_30349 = v_1100;
assign v_30350 = ~v_29371;
assign v_30351 = ~v_1104;
assign v_30352 = v_1104;
assign v_30353 = ~v_29375;
assign v_30354 = ~v_1108;
assign v_30355 = v_1108;
assign v_30356 = ~v_29379;
assign v_30357 = ~v_1112;
assign v_30358 = v_1112;
assign v_30359 = ~v_29383;
assign v_30360 = ~v_1116;
assign v_30361 = v_1116;
assign v_30362 = ~v_29387;
assign v_30363 = ~v_1120;
assign v_30364 = v_1120;
assign v_30365 = ~v_29391;
assign v_30366 = ~v_1124;
assign v_30367 = v_1124;
assign v_30368 = ~v_29395;
assign v_30369 = ~v_1128;
assign v_30370 = v_30369;
assign v_30372 = v_30371;
assign v_30374 = v_30366 & v_30373;
assign v_30376 = v_29391;
assign v_30378 = v_30375 & v_30377;
assign v_30380 = v_30363 & v_30379;
assign v_30382 = v_29387;
assign v_30384 = v_30381 & v_30383;
assign v_30386 = v_30360 & v_30385;
assign v_30388 = v_29383;
assign v_30390 = v_30387 & v_30389;
assign v_30392 = v_30357 & v_30391;
assign v_30394 = v_29379;
assign v_30396 = v_30393 & v_30395;
assign v_30398 = v_30354 & v_30397;
assign v_30400 = v_29375;
assign v_30402 = v_30399 & v_30401;
assign v_30404 = v_30351 & v_30403;
assign v_30406 = v_29371;
assign v_30408 = v_30405 & v_30407;
assign v_30410 = v_30348 & v_30409;
assign v_30412 = v_29367;
assign v_30414 = v_30411 & v_30413;
assign v_30416 = v_30345 & v_30415;
assign v_30418 = v_29363;
assign v_30420 = v_30417 & v_30419;
assign v_30422 = v_30342 & v_30421;
assign v_30424 = v_29359;
assign v_30426 = v_30423 & v_30425;
assign v_30428 = v_30339 & v_30427;
assign v_30430 = v_29355;
assign v_30432 = v_30429 & v_30431;
assign v_30434 = v_30336 & v_30433;
assign v_30436 = v_29351;
assign v_30438 = v_30435 & v_30437;
assign v_30440 = v_30333 & v_30439;
assign v_30442 = v_29347;
assign v_30444 = v_30441 & v_30443;
assign v_30446 = v_30330 & v_30445;
assign v_30448 = v_1075;
assign v_30450 = v_30447 & v_30449;
assign v_30452 = v_30327 & v_30451;
assign v_30454 = v_1071;
assign v_30456 = v_30453 & v_30455;
assign v_30458 = v_30324 & v_30457;
assign v_30460 = v_1067;
assign v_30462 = v_30459 & v_30461;
assign v_30464 = v_30321 & v_30463;
assign v_30466 = v_1063;
assign v_30468 = v_30465 & v_30467;
assign v_30469 = v_30468;
assign v_30471 = v_29395;
assign v_30472 = v_1128;
assign v_30473 = v_30472;
assign v_30474 = v_30471 & v_30473;
assign v_30475 = v_30474;
assign v_30476 = v_30366 & v_30475;
assign v_30478 = v_30376 & v_30477;
assign v_30479 = v_30365 & v_30475;
assign v_30481 = v_30363 & v_30480;
assign v_30483 = v_30382 & v_30482;
assign v_30484 = v_30362 & v_30480;
assign v_30486 = v_30360 & v_30485;
assign v_30488 = v_30388 & v_30487;
assign v_30489 = v_30359 & v_30485;
assign v_30491 = v_30357 & v_30490;
assign v_30493 = v_30394 & v_30492;
assign v_30494 = v_30356 & v_30490;
assign v_30496 = v_30354 & v_30495;
assign v_30498 = v_30400 & v_30497;
assign v_30499 = v_30353 & v_30495;
assign v_30501 = v_30351 & v_30500;
assign v_30503 = v_30406 & v_30502;
assign v_30504 = v_30350 & v_30500;
assign v_30506 = v_30348 & v_30505;
assign v_30508 = v_30412 & v_30507;
assign v_30509 = v_30347 & v_30505;
assign v_30511 = v_30345 & v_30510;
assign v_30513 = v_30418 & v_30512;
assign v_30514 = v_30344 & v_30510;
assign v_30516 = v_30342 & v_30515;
assign v_30518 = v_30424 & v_30517;
assign v_30519 = v_30341 & v_30515;
assign v_30521 = v_30339 & v_30520;
assign v_30523 = v_30430 & v_30522;
assign v_30524 = v_30338 & v_30520;
assign v_30526 = v_30336 & v_30525;
assign v_30528 = v_30436 & v_30527;
assign v_30529 = v_30335 & v_30525;
assign v_30531 = v_30333 & v_30530;
assign v_30533 = v_30442 & v_30532;
assign v_30534 = v_30332 & v_30530;
assign v_30536 = v_30330 & v_30535;
assign v_30538 = v_30448 & v_30537;
assign v_30539 = v_30329 & v_30535;
assign v_30541 = v_30327 & v_30540;
assign v_30543 = v_30454 & v_30542;
assign v_30544 = v_30326 & v_30540;
assign v_30546 = v_30324 & v_30545;
assign v_30548 = v_30460 & v_30547;
assign v_30549 = v_30323 & v_30545;
assign v_30551 = v_30321 & v_30550;
assign v_30553 = v_30466 & v_30552;
assign v_30554 = v_30320 & v_30550;
assign v_30556 = v_30555;
assign v_30558 = v_30470 & v_30557;
assign v_30559 = v_30558;
assign v_30561 = v_30560;
assign v_30563 = ~v_1323;
assign v_30564 = ~v_29332;
assign v_30565 = v_29332;
assign v_30566 = ~v_1327;
assign v_30567 = ~v_29336;
assign v_30568 = v_29336;
assign v_30569 = ~v_1331;
assign v_30570 = ~v_29340;
assign v_30571 = v_29340;
assign v_30572 = ~v_1335;
assign v_30573 = ~v_29344;
assign v_30574 = v_29344;
assign v_30575 = ~v_29347;
assign v_30576 = ~v_1340;
assign v_30577 = v_1340;
assign v_30578 = ~v_29351;
assign v_30579 = ~v_1344;
assign v_30580 = v_1344;
assign v_30581 = ~v_29355;
assign v_30582 = ~v_1348;
assign v_30583 = v_1348;
assign v_30584 = ~v_29359;
assign v_30585 = ~v_1352;
assign v_30586 = v_1352;
assign v_30587 = ~v_29363;
assign v_30588 = ~v_1356;
assign v_30589 = v_1356;
assign v_30590 = ~v_29367;
assign v_30591 = ~v_1360;
assign v_30592 = v_1360;
assign v_30593 = ~v_29371;
assign v_30594 = ~v_1364;
assign v_30595 = v_1364;
assign v_30596 = ~v_29375;
assign v_30597 = ~v_1368;
assign v_30598 = v_1368;
assign v_30599 = ~v_29379;
assign v_30600 = ~v_1372;
assign v_30601 = v_1372;
assign v_30602 = ~v_29383;
assign v_30603 = ~v_1376;
assign v_30604 = v_1376;
assign v_30605 = ~v_29387;
assign v_30606 = ~v_1380;
assign v_30607 = v_1380;
assign v_30608 = ~v_29391;
assign v_30609 = ~v_1384;
assign v_30610 = v_1384;
assign v_30611 = ~v_29395;
assign v_30612 = ~v_1388;
assign v_30613 = v_30612;
assign v_30615 = v_30614;
assign v_30617 = v_30609 & v_30616;
assign v_30619 = v_29391;
assign v_30621 = v_30618 & v_30620;
assign v_30623 = v_30606 & v_30622;
assign v_30625 = v_29387;
assign v_30627 = v_30624 & v_30626;
assign v_30629 = v_30603 & v_30628;
assign v_30631 = v_29383;
assign v_30633 = v_30630 & v_30632;
assign v_30635 = v_30600 & v_30634;
assign v_30637 = v_29379;
assign v_30639 = v_30636 & v_30638;
assign v_30641 = v_30597 & v_30640;
assign v_30643 = v_29375;
assign v_30645 = v_30642 & v_30644;
assign v_30647 = v_30594 & v_30646;
assign v_30649 = v_29371;
assign v_30651 = v_30648 & v_30650;
assign v_30653 = v_30591 & v_30652;
assign v_30655 = v_29367;
assign v_30657 = v_30654 & v_30656;
assign v_30659 = v_30588 & v_30658;
assign v_30661 = v_29363;
assign v_30663 = v_30660 & v_30662;
assign v_30665 = v_30585 & v_30664;
assign v_30667 = v_29359;
assign v_30669 = v_30666 & v_30668;
assign v_30671 = v_30582 & v_30670;
assign v_30673 = v_29355;
assign v_30675 = v_30672 & v_30674;
assign v_30677 = v_30579 & v_30676;
assign v_30679 = v_29351;
assign v_30681 = v_30678 & v_30680;
assign v_30683 = v_30576 & v_30682;
assign v_30685 = v_29347;
assign v_30687 = v_30684 & v_30686;
assign v_30689 = v_30573 & v_30688;
assign v_30691 = v_1335;
assign v_30693 = v_30690 & v_30692;
assign v_30695 = v_30570 & v_30694;
assign v_30697 = v_1331;
assign v_30699 = v_30696 & v_30698;
assign v_30701 = v_30567 & v_30700;
assign v_30703 = v_1327;
assign v_30705 = v_30702 & v_30704;
assign v_30707 = v_30564 & v_30706;
assign v_30709 = v_1323;
assign v_30711 = v_30708 & v_30710;
assign v_30712 = v_30711;
assign v_30714 = v_29395;
assign v_30715 = v_1388;
assign v_30716 = v_30715;
assign v_30717 = v_30714 & v_30716;
assign v_30718 = v_30717;
assign v_30719 = v_30609 & v_30718;
assign v_30721 = v_30619 & v_30720;
assign v_30722 = v_30608 & v_30718;
assign v_30724 = v_30606 & v_30723;
assign v_30726 = v_30625 & v_30725;
assign v_30727 = v_30605 & v_30723;
assign v_30729 = v_30603 & v_30728;
assign v_30731 = v_30631 & v_30730;
assign v_30732 = v_30602 & v_30728;
assign v_30734 = v_30600 & v_30733;
assign v_30736 = v_30637 & v_30735;
assign v_30737 = v_30599 & v_30733;
assign v_30739 = v_30597 & v_30738;
assign v_30741 = v_30643 & v_30740;
assign v_30742 = v_30596 & v_30738;
assign v_30744 = v_30594 & v_30743;
assign v_30746 = v_30649 & v_30745;
assign v_30747 = v_30593 & v_30743;
assign v_30749 = v_30591 & v_30748;
assign v_30751 = v_30655 & v_30750;
assign v_30752 = v_30590 & v_30748;
assign v_30754 = v_30588 & v_30753;
assign v_30756 = v_30661 & v_30755;
assign v_30757 = v_30587 & v_30753;
assign v_30759 = v_30585 & v_30758;
assign v_30761 = v_30667 & v_30760;
assign v_30762 = v_30584 & v_30758;
assign v_30764 = v_30582 & v_30763;
assign v_30766 = v_30673 & v_30765;
assign v_30767 = v_30581 & v_30763;
assign v_30769 = v_30579 & v_30768;
assign v_30771 = v_30679 & v_30770;
assign v_30772 = v_30578 & v_30768;
assign v_30774 = v_30576 & v_30773;
assign v_30776 = v_30685 & v_30775;
assign v_30777 = v_30575 & v_30773;
assign v_30779 = v_30573 & v_30778;
assign v_30781 = v_30691 & v_30780;
assign v_30782 = v_30572 & v_30778;
assign v_30784 = v_30570 & v_30783;
assign v_30786 = v_30697 & v_30785;
assign v_30787 = v_30569 & v_30783;
assign v_30789 = v_30567 & v_30788;
assign v_30791 = v_30703 & v_30790;
assign v_30792 = v_30566 & v_30788;
assign v_30794 = v_30564 & v_30793;
assign v_30796 = v_30709 & v_30795;
assign v_30797 = v_30563 & v_30793;
assign v_30799 = v_30798;
assign v_30801 = v_30713 & v_30800;
assign v_30802 = v_30801;
assign v_30804 = v_30803;
assign v_30806 = ~v_1583;
assign v_30807 = ~v_29332;
assign v_30808 = v_29332;
assign v_30809 = ~v_1587;
assign v_30810 = ~v_29336;
assign v_30811 = v_29336;
assign v_30812 = ~v_1591;
assign v_30813 = ~v_29340;
assign v_30814 = v_29340;
assign v_30815 = ~v_1595;
assign v_30816 = ~v_29344;
assign v_30817 = v_29344;
assign v_30818 = ~v_29347;
assign v_30819 = ~v_1600;
assign v_30820 = v_1600;
assign v_30821 = ~v_29351;
assign v_30822 = ~v_1604;
assign v_30823 = v_1604;
assign v_30824 = ~v_29355;
assign v_30825 = ~v_1608;
assign v_30826 = v_1608;
assign v_30827 = ~v_29359;
assign v_30828 = ~v_1612;
assign v_30829 = v_1612;
assign v_30830 = ~v_29363;
assign v_30831 = ~v_1616;
assign v_30832 = v_1616;
assign v_30833 = ~v_29367;
assign v_30834 = ~v_1620;
assign v_30835 = v_1620;
assign v_30836 = ~v_29371;
assign v_30837 = ~v_1624;
assign v_30838 = v_1624;
assign v_30839 = ~v_29375;
assign v_30840 = ~v_1628;
assign v_30841 = v_1628;
assign v_30842 = ~v_29379;
assign v_30843 = ~v_1632;
assign v_30844 = v_1632;
assign v_30845 = ~v_29383;
assign v_30846 = ~v_1636;
assign v_30847 = v_1636;
assign v_30848 = ~v_29387;
assign v_30849 = ~v_1640;
assign v_30850 = v_1640;
assign v_30851 = ~v_29391;
assign v_30852 = ~v_1644;
assign v_30853 = v_1644;
assign v_30854 = ~v_29395;
assign v_30855 = ~v_1648;
assign v_30856 = v_30855;
assign v_30858 = v_30857;
assign v_30860 = v_30852 & v_30859;
assign v_30862 = v_29391;
assign v_30864 = v_30861 & v_30863;
assign v_30866 = v_30849 & v_30865;
assign v_30868 = v_29387;
assign v_30870 = v_30867 & v_30869;
assign v_30872 = v_30846 & v_30871;
assign v_30874 = v_29383;
assign v_30876 = v_30873 & v_30875;
assign v_30878 = v_30843 & v_30877;
assign v_30880 = v_29379;
assign v_30882 = v_30879 & v_30881;
assign v_30884 = v_30840 & v_30883;
assign v_30886 = v_29375;
assign v_30888 = v_30885 & v_30887;
assign v_30890 = v_30837 & v_30889;
assign v_30892 = v_29371;
assign v_30894 = v_30891 & v_30893;
assign v_30896 = v_30834 & v_30895;
assign v_30898 = v_29367;
assign v_30900 = v_30897 & v_30899;
assign v_30902 = v_30831 & v_30901;
assign v_30904 = v_29363;
assign v_30906 = v_30903 & v_30905;
assign v_30908 = v_30828 & v_30907;
assign v_30910 = v_29359;
assign v_30912 = v_30909 & v_30911;
assign v_30914 = v_30825 & v_30913;
assign v_30916 = v_29355;
assign v_30918 = v_30915 & v_30917;
assign v_30920 = v_30822 & v_30919;
assign v_30922 = v_29351;
assign v_30924 = v_30921 & v_30923;
assign v_30926 = v_30819 & v_30925;
assign v_30928 = v_29347;
assign v_30930 = v_30927 & v_30929;
assign v_30932 = v_30816 & v_30931;
assign v_30934 = v_1595;
assign v_30936 = v_30933 & v_30935;
assign v_30938 = v_30813 & v_30937;
assign v_30940 = v_1591;
assign v_30942 = v_30939 & v_30941;
assign v_30944 = v_30810 & v_30943;
assign v_30946 = v_1587;
assign v_30948 = v_30945 & v_30947;
assign v_30950 = v_30807 & v_30949;
assign v_30952 = v_1583;
assign v_30954 = v_30951 & v_30953;
assign v_30955 = v_30954;
assign v_30957 = v_29395;
assign v_30958 = v_1648;
assign v_30959 = v_30958;
assign v_30960 = v_30957 & v_30959;
assign v_30961 = v_30960;
assign v_30962 = v_30852 & v_30961;
assign v_30964 = v_30862 & v_30963;
assign v_30965 = v_30851 & v_30961;
assign v_30967 = v_30849 & v_30966;
assign v_30969 = v_30868 & v_30968;
assign v_30970 = v_30848 & v_30966;
assign v_30972 = v_30846 & v_30971;
assign v_30974 = v_30874 & v_30973;
assign v_30975 = v_30845 & v_30971;
assign v_30977 = v_30843 & v_30976;
assign v_30979 = v_30880 & v_30978;
assign v_30980 = v_30842 & v_30976;
assign v_30982 = v_30840 & v_30981;
assign v_30984 = v_30886 & v_30983;
assign v_30985 = v_30839 & v_30981;
assign v_30987 = v_30837 & v_30986;
assign v_30989 = v_30892 & v_30988;
assign v_30990 = v_30836 & v_30986;
assign v_30992 = v_30834 & v_30991;
assign v_30994 = v_30898 & v_30993;
assign v_30995 = v_30833 & v_30991;
assign v_30997 = v_30831 & v_30996;
assign v_30999 = v_30904 & v_30998;
assign v_31000 = v_30830 & v_30996;
assign v_31002 = v_30828 & v_31001;
assign v_31004 = v_30910 & v_31003;
assign v_31005 = v_30827 & v_31001;
assign v_31007 = v_30825 & v_31006;
assign v_31009 = v_30916 & v_31008;
assign v_31010 = v_30824 & v_31006;
assign v_31012 = v_30822 & v_31011;
assign v_31014 = v_30922 & v_31013;
assign v_31015 = v_30821 & v_31011;
assign v_31017 = v_30819 & v_31016;
assign v_31019 = v_30928 & v_31018;
assign v_31020 = v_30818 & v_31016;
assign v_31022 = v_30816 & v_31021;
assign v_31024 = v_30934 & v_31023;
assign v_31025 = v_30815 & v_31021;
assign v_31027 = v_30813 & v_31026;
assign v_31029 = v_30940 & v_31028;
assign v_31030 = v_30812 & v_31026;
assign v_31032 = v_30810 & v_31031;
assign v_31034 = v_30946 & v_31033;
assign v_31035 = v_30809 & v_31031;
assign v_31037 = v_30807 & v_31036;
assign v_31039 = v_30952 & v_31038;
assign v_31040 = v_30806 & v_31036;
assign v_31042 = v_31041;
assign v_31044 = v_30956 & v_31043;
assign v_31045 = v_31044;
assign v_31047 = v_31046;
assign v_31049 = ~v_1843;
assign v_31050 = ~v_29332;
assign v_31051 = v_29332;
assign v_31052 = ~v_1847;
assign v_31053 = ~v_29336;
assign v_31054 = v_29336;
assign v_31055 = ~v_1851;
assign v_31056 = ~v_29340;
assign v_31057 = v_29340;
assign v_31058 = ~v_1855;
assign v_31059 = ~v_29344;
assign v_31060 = v_29344;
assign v_31061 = ~v_29347;
assign v_31062 = ~v_1860;
assign v_31063 = v_1860;
assign v_31064 = ~v_29351;
assign v_31065 = ~v_1864;
assign v_31066 = v_1864;
assign v_31067 = ~v_29355;
assign v_31068 = ~v_1868;
assign v_31069 = v_1868;
assign v_31070 = ~v_29359;
assign v_31071 = ~v_1872;
assign v_31072 = v_1872;
assign v_31073 = ~v_29363;
assign v_31074 = ~v_1876;
assign v_31075 = v_1876;
assign v_31076 = ~v_29367;
assign v_31077 = ~v_1880;
assign v_31078 = v_1880;
assign v_31079 = ~v_29371;
assign v_31080 = ~v_1884;
assign v_31081 = v_1884;
assign v_31082 = ~v_29375;
assign v_31083 = ~v_1888;
assign v_31084 = v_1888;
assign v_31085 = ~v_29379;
assign v_31086 = ~v_1892;
assign v_31087 = v_1892;
assign v_31088 = ~v_29383;
assign v_31089 = ~v_1896;
assign v_31090 = v_1896;
assign v_31091 = ~v_29387;
assign v_31092 = ~v_1900;
assign v_31093 = v_1900;
assign v_31094 = ~v_29391;
assign v_31095 = ~v_1904;
assign v_31096 = v_1904;
assign v_31097 = ~v_29395;
assign v_31098 = ~v_1908;
assign v_31099 = v_31098;
assign v_31101 = v_31100;
assign v_31103 = v_31095 & v_31102;
assign v_31105 = v_29391;
assign v_31107 = v_31104 & v_31106;
assign v_31109 = v_31092 & v_31108;
assign v_31111 = v_29387;
assign v_31113 = v_31110 & v_31112;
assign v_31115 = v_31089 & v_31114;
assign v_31117 = v_29383;
assign v_31119 = v_31116 & v_31118;
assign v_31121 = v_31086 & v_31120;
assign v_31123 = v_29379;
assign v_31125 = v_31122 & v_31124;
assign v_31127 = v_31083 & v_31126;
assign v_31129 = v_29375;
assign v_31131 = v_31128 & v_31130;
assign v_31133 = v_31080 & v_31132;
assign v_31135 = v_29371;
assign v_31137 = v_31134 & v_31136;
assign v_31139 = v_31077 & v_31138;
assign v_31141 = v_29367;
assign v_31143 = v_31140 & v_31142;
assign v_31145 = v_31074 & v_31144;
assign v_31147 = v_29363;
assign v_31149 = v_31146 & v_31148;
assign v_31151 = v_31071 & v_31150;
assign v_31153 = v_29359;
assign v_31155 = v_31152 & v_31154;
assign v_31157 = v_31068 & v_31156;
assign v_31159 = v_29355;
assign v_31161 = v_31158 & v_31160;
assign v_31163 = v_31065 & v_31162;
assign v_31165 = v_29351;
assign v_31167 = v_31164 & v_31166;
assign v_31169 = v_31062 & v_31168;
assign v_31171 = v_29347;
assign v_31173 = v_31170 & v_31172;
assign v_31175 = v_31059 & v_31174;
assign v_31177 = v_1855;
assign v_31179 = v_31176 & v_31178;
assign v_31181 = v_31056 & v_31180;
assign v_31183 = v_1851;
assign v_31185 = v_31182 & v_31184;
assign v_31187 = v_31053 & v_31186;
assign v_31189 = v_1847;
assign v_31191 = v_31188 & v_31190;
assign v_31193 = v_31050 & v_31192;
assign v_31195 = v_1843;
assign v_31197 = v_31194 & v_31196;
assign v_31198 = v_31197;
assign v_31200 = v_29395;
assign v_31201 = v_1908;
assign v_31202 = v_31201;
assign v_31203 = v_31200 & v_31202;
assign v_31204 = v_31203;
assign v_31205 = v_31095 & v_31204;
assign v_31207 = v_31105 & v_31206;
assign v_31208 = v_31094 & v_31204;
assign v_31210 = v_31092 & v_31209;
assign v_31212 = v_31111 & v_31211;
assign v_31213 = v_31091 & v_31209;
assign v_31215 = v_31089 & v_31214;
assign v_31217 = v_31117 & v_31216;
assign v_31218 = v_31088 & v_31214;
assign v_31220 = v_31086 & v_31219;
assign v_31222 = v_31123 & v_31221;
assign v_31223 = v_31085 & v_31219;
assign v_31225 = v_31083 & v_31224;
assign v_31227 = v_31129 & v_31226;
assign v_31228 = v_31082 & v_31224;
assign v_31230 = v_31080 & v_31229;
assign v_31232 = v_31135 & v_31231;
assign v_31233 = v_31079 & v_31229;
assign v_31235 = v_31077 & v_31234;
assign v_31237 = v_31141 & v_31236;
assign v_31238 = v_31076 & v_31234;
assign v_31240 = v_31074 & v_31239;
assign v_31242 = v_31147 & v_31241;
assign v_31243 = v_31073 & v_31239;
assign v_31245 = v_31071 & v_31244;
assign v_31247 = v_31153 & v_31246;
assign v_31248 = v_31070 & v_31244;
assign v_31250 = v_31068 & v_31249;
assign v_31252 = v_31159 & v_31251;
assign v_31253 = v_31067 & v_31249;
assign v_31255 = v_31065 & v_31254;
assign v_31257 = v_31165 & v_31256;
assign v_31258 = v_31064 & v_31254;
assign v_31260 = v_31062 & v_31259;
assign v_31262 = v_31171 & v_31261;
assign v_31263 = v_31061 & v_31259;
assign v_31265 = v_31059 & v_31264;
assign v_31267 = v_31177 & v_31266;
assign v_31268 = v_31058 & v_31264;
assign v_31270 = v_31056 & v_31269;
assign v_31272 = v_31183 & v_31271;
assign v_31273 = v_31055 & v_31269;
assign v_31275 = v_31053 & v_31274;
assign v_31277 = v_31189 & v_31276;
assign v_31278 = v_31052 & v_31274;
assign v_31280 = v_31050 & v_31279;
assign v_31282 = v_31195 & v_31281;
assign v_31283 = v_31049 & v_31279;
assign v_31285 = v_31284;
assign v_31287 = v_31199 & v_31286;
assign v_31288 = v_31287;
assign v_31290 = v_31289;
assign v_31292 = ~v_2103;
assign v_31293 = ~v_29332;
assign v_31294 = v_29332;
assign v_31295 = ~v_2107;
assign v_31296 = ~v_29336;
assign v_31297 = v_29336;
assign v_31298 = ~v_2111;
assign v_31299 = ~v_29340;
assign v_31300 = v_29340;
assign v_31301 = ~v_2115;
assign v_31302 = ~v_29344;
assign v_31303 = v_29344;
assign v_31304 = ~v_29347;
assign v_31305 = ~v_2120;
assign v_31306 = v_2120;
assign v_31307 = ~v_29351;
assign v_31308 = ~v_2124;
assign v_31309 = v_2124;
assign v_31310 = ~v_29355;
assign v_31311 = ~v_2128;
assign v_31312 = v_2128;
assign v_31313 = ~v_29359;
assign v_31314 = ~v_2132;
assign v_31315 = v_2132;
assign v_31316 = ~v_29363;
assign v_31317 = ~v_2136;
assign v_31318 = v_2136;
assign v_31319 = ~v_29367;
assign v_31320 = ~v_2140;
assign v_31321 = v_2140;
assign v_31322 = ~v_29371;
assign v_31323 = ~v_2144;
assign v_31324 = v_2144;
assign v_31325 = ~v_29375;
assign v_31326 = ~v_2148;
assign v_31327 = v_2148;
assign v_31328 = ~v_29379;
assign v_31329 = ~v_2152;
assign v_31330 = v_2152;
assign v_31331 = ~v_29383;
assign v_31332 = ~v_2156;
assign v_31333 = v_2156;
assign v_31334 = ~v_29387;
assign v_31335 = ~v_2160;
assign v_31336 = v_2160;
assign v_31337 = ~v_29391;
assign v_31338 = ~v_2164;
assign v_31339 = v_2164;
assign v_31340 = ~v_29395;
assign v_31341 = ~v_2168;
assign v_31342 = v_31341;
assign v_31344 = v_31343;
assign v_31346 = v_31338 & v_31345;
assign v_31348 = v_29391;
assign v_31350 = v_31347 & v_31349;
assign v_31352 = v_31335 & v_31351;
assign v_31354 = v_29387;
assign v_31356 = v_31353 & v_31355;
assign v_31358 = v_31332 & v_31357;
assign v_31360 = v_29383;
assign v_31362 = v_31359 & v_31361;
assign v_31364 = v_31329 & v_31363;
assign v_31366 = v_29379;
assign v_31368 = v_31365 & v_31367;
assign v_31370 = v_31326 & v_31369;
assign v_31372 = v_29375;
assign v_31374 = v_31371 & v_31373;
assign v_31376 = v_31323 & v_31375;
assign v_31378 = v_29371;
assign v_31380 = v_31377 & v_31379;
assign v_31382 = v_31320 & v_31381;
assign v_31384 = v_29367;
assign v_31386 = v_31383 & v_31385;
assign v_31388 = v_31317 & v_31387;
assign v_31390 = v_29363;
assign v_31392 = v_31389 & v_31391;
assign v_31394 = v_31314 & v_31393;
assign v_31396 = v_29359;
assign v_31398 = v_31395 & v_31397;
assign v_31400 = v_31311 & v_31399;
assign v_31402 = v_29355;
assign v_31404 = v_31401 & v_31403;
assign v_31406 = v_31308 & v_31405;
assign v_31408 = v_29351;
assign v_31410 = v_31407 & v_31409;
assign v_31412 = v_31305 & v_31411;
assign v_31414 = v_29347;
assign v_31416 = v_31413 & v_31415;
assign v_31418 = v_31302 & v_31417;
assign v_31420 = v_2115;
assign v_31422 = v_31419 & v_31421;
assign v_31424 = v_31299 & v_31423;
assign v_31426 = v_2111;
assign v_31428 = v_31425 & v_31427;
assign v_31430 = v_31296 & v_31429;
assign v_31432 = v_2107;
assign v_31434 = v_31431 & v_31433;
assign v_31436 = v_31293 & v_31435;
assign v_31438 = v_2103;
assign v_31440 = v_31437 & v_31439;
assign v_31441 = v_31440;
assign v_31443 = v_29395;
assign v_31444 = v_2168;
assign v_31445 = v_31444;
assign v_31446 = v_31443 & v_31445;
assign v_31447 = v_31446;
assign v_31448 = v_31338 & v_31447;
assign v_31450 = v_31348 & v_31449;
assign v_31451 = v_31337 & v_31447;
assign v_31453 = v_31335 & v_31452;
assign v_31455 = v_31354 & v_31454;
assign v_31456 = v_31334 & v_31452;
assign v_31458 = v_31332 & v_31457;
assign v_31460 = v_31360 & v_31459;
assign v_31461 = v_31331 & v_31457;
assign v_31463 = v_31329 & v_31462;
assign v_31465 = v_31366 & v_31464;
assign v_31466 = v_31328 & v_31462;
assign v_31468 = v_31326 & v_31467;
assign v_31470 = v_31372 & v_31469;
assign v_31471 = v_31325 & v_31467;
assign v_31473 = v_31323 & v_31472;
assign v_31475 = v_31378 & v_31474;
assign v_31476 = v_31322 & v_31472;
assign v_31478 = v_31320 & v_31477;
assign v_31480 = v_31384 & v_31479;
assign v_31481 = v_31319 & v_31477;
assign v_31483 = v_31317 & v_31482;
assign v_31485 = v_31390 & v_31484;
assign v_31486 = v_31316 & v_31482;
assign v_31488 = v_31314 & v_31487;
assign v_31490 = v_31396 & v_31489;
assign v_31491 = v_31313 & v_31487;
assign v_31493 = v_31311 & v_31492;
assign v_31495 = v_31402 & v_31494;
assign v_31496 = v_31310 & v_31492;
assign v_31498 = v_31308 & v_31497;
assign v_31500 = v_31408 & v_31499;
assign v_31501 = v_31307 & v_31497;
assign v_31503 = v_31305 & v_31502;
assign v_31505 = v_31414 & v_31504;
assign v_31506 = v_31304 & v_31502;
assign v_31508 = v_31302 & v_31507;
assign v_31510 = v_31420 & v_31509;
assign v_31511 = v_31301 & v_31507;
assign v_31513 = v_31299 & v_31512;
assign v_31515 = v_31426 & v_31514;
assign v_31516 = v_31298 & v_31512;
assign v_31518 = v_31296 & v_31517;
assign v_31520 = v_31432 & v_31519;
assign v_31521 = v_31295 & v_31517;
assign v_31523 = v_31293 & v_31522;
assign v_31525 = v_31438 & v_31524;
assign v_31526 = v_31292 & v_31522;
assign v_31528 = v_31527;
assign v_31530 = v_31442 & v_31529;
assign v_31531 = v_31530;
assign v_31533 = v_31532;
assign v_31535 = ~v_2363;
assign v_31536 = ~v_29332;
assign v_31537 = v_29332;
assign v_31538 = ~v_2367;
assign v_31539 = ~v_29336;
assign v_31540 = v_29336;
assign v_31541 = ~v_2371;
assign v_31542 = ~v_29340;
assign v_31543 = v_29340;
assign v_31544 = ~v_2375;
assign v_31545 = ~v_29344;
assign v_31546 = v_29344;
assign v_31547 = ~v_29347;
assign v_31548 = ~v_2380;
assign v_31549 = v_2380;
assign v_31550 = ~v_29351;
assign v_31551 = ~v_2384;
assign v_31552 = v_2384;
assign v_31553 = ~v_29355;
assign v_31554 = ~v_2388;
assign v_31555 = v_2388;
assign v_31556 = ~v_29359;
assign v_31557 = ~v_2392;
assign v_31558 = v_2392;
assign v_31559 = ~v_29363;
assign v_31560 = ~v_2396;
assign v_31561 = v_2396;
assign v_31562 = ~v_29367;
assign v_31563 = ~v_2400;
assign v_31564 = v_2400;
assign v_31565 = ~v_29371;
assign v_31566 = ~v_2404;
assign v_31567 = v_2404;
assign v_31568 = ~v_29375;
assign v_31569 = ~v_2408;
assign v_31570 = v_2408;
assign v_31571 = ~v_29379;
assign v_31572 = ~v_2412;
assign v_31573 = v_2412;
assign v_31574 = ~v_29383;
assign v_31575 = ~v_2416;
assign v_31576 = v_2416;
assign v_31577 = ~v_29387;
assign v_31578 = ~v_2420;
assign v_31579 = v_2420;
assign v_31580 = ~v_29391;
assign v_31581 = ~v_2424;
assign v_31582 = v_2424;
assign v_31583 = ~v_29395;
assign v_31584 = ~v_2428;
assign v_31585 = v_31584;
assign v_31587 = v_31586;
assign v_31589 = v_31581 & v_31588;
assign v_31591 = v_29391;
assign v_31593 = v_31590 & v_31592;
assign v_31595 = v_31578 & v_31594;
assign v_31597 = v_29387;
assign v_31599 = v_31596 & v_31598;
assign v_31601 = v_31575 & v_31600;
assign v_31603 = v_29383;
assign v_31605 = v_31602 & v_31604;
assign v_31607 = v_31572 & v_31606;
assign v_31609 = v_29379;
assign v_31611 = v_31608 & v_31610;
assign v_31613 = v_31569 & v_31612;
assign v_31615 = v_29375;
assign v_31617 = v_31614 & v_31616;
assign v_31619 = v_31566 & v_31618;
assign v_31621 = v_29371;
assign v_31623 = v_31620 & v_31622;
assign v_31625 = v_31563 & v_31624;
assign v_31627 = v_29367;
assign v_31629 = v_31626 & v_31628;
assign v_31631 = v_31560 & v_31630;
assign v_31633 = v_29363;
assign v_31635 = v_31632 & v_31634;
assign v_31637 = v_31557 & v_31636;
assign v_31639 = v_29359;
assign v_31641 = v_31638 & v_31640;
assign v_31643 = v_31554 & v_31642;
assign v_31645 = v_29355;
assign v_31647 = v_31644 & v_31646;
assign v_31649 = v_31551 & v_31648;
assign v_31651 = v_29351;
assign v_31653 = v_31650 & v_31652;
assign v_31655 = v_31548 & v_31654;
assign v_31657 = v_29347;
assign v_31659 = v_31656 & v_31658;
assign v_31661 = v_31545 & v_31660;
assign v_31663 = v_2375;
assign v_31665 = v_31662 & v_31664;
assign v_31667 = v_31542 & v_31666;
assign v_31669 = v_2371;
assign v_31671 = v_31668 & v_31670;
assign v_31673 = v_31539 & v_31672;
assign v_31675 = v_2367;
assign v_31677 = v_31674 & v_31676;
assign v_31679 = v_31536 & v_31678;
assign v_31681 = v_2363;
assign v_31683 = v_31680 & v_31682;
assign v_31684 = v_31683;
assign v_31686 = v_29395;
assign v_31687 = v_2428;
assign v_31688 = v_31687;
assign v_31689 = v_31686 & v_31688;
assign v_31690 = v_31689;
assign v_31691 = v_31581 & v_31690;
assign v_31693 = v_31591 & v_31692;
assign v_31694 = v_31580 & v_31690;
assign v_31696 = v_31578 & v_31695;
assign v_31698 = v_31597 & v_31697;
assign v_31699 = v_31577 & v_31695;
assign v_31701 = v_31575 & v_31700;
assign v_31703 = v_31603 & v_31702;
assign v_31704 = v_31574 & v_31700;
assign v_31706 = v_31572 & v_31705;
assign v_31708 = v_31609 & v_31707;
assign v_31709 = v_31571 & v_31705;
assign v_31711 = v_31569 & v_31710;
assign v_31713 = v_31615 & v_31712;
assign v_31714 = v_31568 & v_31710;
assign v_31716 = v_31566 & v_31715;
assign v_31718 = v_31621 & v_31717;
assign v_31719 = v_31565 & v_31715;
assign v_31721 = v_31563 & v_31720;
assign v_31723 = v_31627 & v_31722;
assign v_31724 = v_31562 & v_31720;
assign v_31726 = v_31560 & v_31725;
assign v_31728 = v_31633 & v_31727;
assign v_31729 = v_31559 & v_31725;
assign v_31731 = v_31557 & v_31730;
assign v_31733 = v_31639 & v_31732;
assign v_31734 = v_31556 & v_31730;
assign v_31736 = v_31554 & v_31735;
assign v_31738 = v_31645 & v_31737;
assign v_31739 = v_31553 & v_31735;
assign v_31741 = v_31551 & v_31740;
assign v_31743 = v_31651 & v_31742;
assign v_31744 = v_31550 & v_31740;
assign v_31746 = v_31548 & v_31745;
assign v_31748 = v_31657 & v_31747;
assign v_31749 = v_31547 & v_31745;
assign v_31751 = v_31545 & v_31750;
assign v_31753 = v_31663 & v_31752;
assign v_31754 = v_31544 & v_31750;
assign v_31756 = v_31542 & v_31755;
assign v_31758 = v_31669 & v_31757;
assign v_31759 = v_31541 & v_31755;
assign v_31761 = v_31539 & v_31760;
assign v_31763 = v_31675 & v_31762;
assign v_31764 = v_31538 & v_31760;
assign v_31766 = v_31536 & v_31765;
assign v_31768 = v_31681 & v_31767;
assign v_31769 = v_31535 & v_31765;
assign v_31771 = v_31770;
assign v_31773 = v_31685 & v_31772;
assign v_31774 = v_31773;
assign v_31776 = v_31775;
assign v_31778 = ~v_2623;
assign v_31779 = ~v_29332;
assign v_31780 = v_29332;
assign v_31781 = ~v_2627;
assign v_31782 = ~v_29336;
assign v_31783 = v_29336;
assign v_31784 = ~v_2631;
assign v_31785 = ~v_29340;
assign v_31786 = v_29340;
assign v_31787 = ~v_2635;
assign v_31788 = ~v_29344;
assign v_31789 = v_29344;
assign v_31790 = ~v_29347;
assign v_31791 = ~v_2640;
assign v_31792 = v_2640;
assign v_31793 = ~v_29351;
assign v_31794 = ~v_2644;
assign v_31795 = v_2644;
assign v_31796 = ~v_29355;
assign v_31797 = ~v_2648;
assign v_31798 = v_2648;
assign v_31799 = ~v_29359;
assign v_31800 = ~v_2652;
assign v_31801 = v_2652;
assign v_31802 = ~v_29363;
assign v_31803 = ~v_2656;
assign v_31804 = v_2656;
assign v_31805 = ~v_29367;
assign v_31806 = ~v_2660;
assign v_31807 = v_2660;
assign v_31808 = ~v_29371;
assign v_31809 = ~v_2664;
assign v_31810 = v_2664;
assign v_31811 = ~v_29375;
assign v_31812 = ~v_2668;
assign v_31813 = v_2668;
assign v_31814 = ~v_29379;
assign v_31815 = ~v_2672;
assign v_31816 = v_2672;
assign v_31817 = ~v_29383;
assign v_31818 = ~v_2676;
assign v_31819 = v_2676;
assign v_31820 = ~v_29387;
assign v_31821 = ~v_2680;
assign v_31822 = v_2680;
assign v_31823 = ~v_29391;
assign v_31824 = ~v_2684;
assign v_31825 = v_2684;
assign v_31826 = ~v_29395;
assign v_31827 = ~v_2688;
assign v_31828 = v_31827;
assign v_31830 = v_31829;
assign v_31832 = v_31824 & v_31831;
assign v_31834 = v_29391;
assign v_31836 = v_31833 & v_31835;
assign v_31838 = v_31821 & v_31837;
assign v_31840 = v_29387;
assign v_31842 = v_31839 & v_31841;
assign v_31844 = v_31818 & v_31843;
assign v_31846 = v_29383;
assign v_31848 = v_31845 & v_31847;
assign v_31850 = v_31815 & v_31849;
assign v_31852 = v_29379;
assign v_31854 = v_31851 & v_31853;
assign v_31856 = v_31812 & v_31855;
assign v_31858 = v_29375;
assign v_31860 = v_31857 & v_31859;
assign v_31862 = v_31809 & v_31861;
assign v_31864 = v_29371;
assign v_31866 = v_31863 & v_31865;
assign v_31868 = v_31806 & v_31867;
assign v_31870 = v_29367;
assign v_31872 = v_31869 & v_31871;
assign v_31874 = v_31803 & v_31873;
assign v_31876 = v_29363;
assign v_31878 = v_31875 & v_31877;
assign v_31880 = v_31800 & v_31879;
assign v_31882 = v_29359;
assign v_31884 = v_31881 & v_31883;
assign v_31886 = v_31797 & v_31885;
assign v_31888 = v_29355;
assign v_31890 = v_31887 & v_31889;
assign v_31892 = v_31794 & v_31891;
assign v_31894 = v_29351;
assign v_31896 = v_31893 & v_31895;
assign v_31898 = v_31791 & v_31897;
assign v_31900 = v_29347;
assign v_31902 = v_31899 & v_31901;
assign v_31904 = v_31788 & v_31903;
assign v_31906 = v_2635;
assign v_31908 = v_31905 & v_31907;
assign v_31910 = v_31785 & v_31909;
assign v_31912 = v_2631;
assign v_31914 = v_31911 & v_31913;
assign v_31916 = v_31782 & v_31915;
assign v_31918 = v_2627;
assign v_31920 = v_31917 & v_31919;
assign v_31922 = v_31779 & v_31921;
assign v_31924 = v_2623;
assign v_31926 = v_31923 & v_31925;
assign v_31927 = v_31926;
assign v_31929 = v_29395;
assign v_31930 = v_2688;
assign v_31931 = v_31930;
assign v_31932 = v_31929 & v_31931;
assign v_31933 = v_31932;
assign v_31934 = v_31824 & v_31933;
assign v_31936 = v_31834 & v_31935;
assign v_31937 = v_31823 & v_31933;
assign v_31939 = v_31821 & v_31938;
assign v_31941 = v_31840 & v_31940;
assign v_31942 = v_31820 & v_31938;
assign v_31944 = v_31818 & v_31943;
assign v_31946 = v_31846 & v_31945;
assign v_31947 = v_31817 & v_31943;
assign v_31949 = v_31815 & v_31948;
assign v_31951 = v_31852 & v_31950;
assign v_31952 = v_31814 & v_31948;
assign v_31954 = v_31812 & v_31953;
assign v_31956 = v_31858 & v_31955;
assign v_31957 = v_31811 & v_31953;
assign v_31959 = v_31809 & v_31958;
assign v_31961 = v_31864 & v_31960;
assign v_31962 = v_31808 & v_31958;
assign v_31964 = v_31806 & v_31963;
assign v_31966 = v_31870 & v_31965;
assign v_31967 = v_31805 & v_31963;
assign v_31969 = v_31803 & v_31968;
assign v_31971 = v_31876 & v_31970;
assign v_31972 = v_31802 & v_31968;
assign v_31974 = v_31800 & v_31973;
assign v_31976 = v_31882 & v_31975;
assign v_31977 = v_31799 & v_31973;
assign v_31979 = v_31797 & v_31978;
assign v_31981 = v_31888 & v_31980;
assign v_31982 = v_31796 & v_31978;
assign v_31984 = v_31794 & v_31983;
assign v_31986 = v_31894 & v_31985;
assign v_31987 = v_31793 & v_31983;
assign v_31989 = v_31791 & v_31988;
assign v_31991 = v_31900 & v_31990;
assign v_31992 = v_31790 & v_31988;
assign v_31994 = v_31788 & v_31993;
assign v_31996 = v_31906 & v_31995;
assign v_31997 = v_31787 & v_31993;
assign v_31999 = v_31785 & v_31998;
assign v_32001 = v_31912 & v_32000;
assign v_32002 = v_31784 & v_31998;
assign v_32004 = v_31782 & v_32003;
assign v_32006 = v_31918 & v_32005;
assign v_32007 = v_31781 & v_32003;
assign v_32009 = v_31779 & v_32008;
assign v_32011 = v_31924 & v_32010;
assign v_32012 = v_31778 & v_32008;
assign v_32014 = v_32013;
assign v_32016 = v_31928 & v_32015;
assign v_32017 = v_32016;
assign v_32019 = v_32018;
assign v_32021 = ~v_2883;
assign v_32022 = ~v_29332;
assign v_32023 = v_29332;
assign v_32024 = ~v_2887;
assign v_32025 = ~v_29336;
assign v_32026 = v_29336;
assign v_32027 = ~v_2891;
assign v_32028 = ~v_29340;
assign v_32029 = v_29340;
assign v_32030 = ~v_2895;
assign v_32031 = ~v_29344;
assign v_32032 = v_29344;
assign v_32033 = ~v_29347;
assign v_32034 = ~v_2900;
assign v_32035 = v_2900;
assign v_32036 = ~v_29351;
assign v_32037 = ~v_2904;
assign v_32038 = v_2904;
assign v_32039 = ~v_29355;
assign v_32040 = ~v_2908;
assign v_32041 = v_2908;
assign v_32042 = ~v_29359;
assign v_32043 = ~v_2912;
assign v_32044 = v_2912;
assign v_32045 = ~v_29363;
assign v_32046 = ~v_2916;
assign v_32047 = v_2916;
assign v_32048 = ~v_29367;
assign v_32049 = ~v_2920;
assign v_32050 = v_2920;
assign v_32051 = ~v_29371;
assign v_32052 = ~v_2924;
assign v_32053 = v_2924;
assign v_32054 = ~v_29375;
assign v_32055 = ~v_2928;
assign v_32056 = v_2928;
assign v_32057 = ~v_29379;
assign v_32058 = ~v_2932;
assign v_32059 = v_2932;
assign v_32060 = ~v_29383;
assign v_32061 = ~v_2936;
assign v_32062 = v_2936;
assign v_32063 = ~v_29387;
assign v_32064 = ~v_2940;
assign v_32065 = v_2940;
assign v_32066 = ~v_29391;
assign v_32067 = ~v_2944;
assign v_32068 = v_2944;
assign v_32069 = ~v_29395;
assign v_32070 = ~v_2948;
assign v_32071 = v_32070;
assign v_32073 = v_32072;
assign v_32075 = v_32067 & v_32074;
assign v_32077 = v_29391;
assign v_32079 = v_32076 & v_32078;
assign v_32081 = v_32064 & v_32080;
assign v_32083 = v_29387;
assign v_32085 = v_32082 & v_32084;
assign v_32087 = v_32061 & v_32086;
assign v_32089 = v_29383;
assign v_32091 = v_32088 & v_32090;
assign v_32093 = v_32058 & v_32092;
assign v_32095 = v_29379;
assign v_32097 = v_32094 & v_32096;
assign v_32099 = v_32055 & v_32098;
assign v_32101 = v_29375;
assign v_32103 = v_32100 & v_32102;
assign v_32105 = v_32052 & v_32104;
assign v_32107 = v_29371;
assign v_32109 = v_32106 & v_32108;
assign v_32111 = v_32049 & v_32110;
assign v_32113 = v_29367;
assign v_32115 = v_32112 & v_32114;
assign v_32117 = v_32046 & v_32116;
assign v_32119 = v_29363;
assign v_32121 = v_32118 & v_32120;
assign v_32123 = v_32043 & v_32122;
assign v_32125 = v_29359;
assign v_32127 = v_32124 & v_32126;
assign v_32129 = v_32040 & v_32128;
assign v_32131 = v_29355;
assign v_32133 = v_32130 & v_32132;
assign v_32135 = v_32037 & v_32134;
assign v_32137 = v_29351;
assign v_32139 = v_32136 & v_32138;
assign v_32141 = v_32034 & v_32140;
assign v_32143 = v_29347;
assign v_32145 = v_32142 & v_32144;
assign v_32147 = v_32031 & v_32146;
assign v_32149 = v_2895;
assign v_32151 = v_32148 & v_32150;
assign v_32153 = v_32028 & v_32152;
assign v_32155 = v_2891;
assign v_32157 = v_32154 & v_32156;
assign v_32159 = v_32025 & v_32158;
assign v_32161 = v_2887;
assign v_32163 = v_32160 & v_32162;
assign v_32165 = v_32022 & v_32164;
assign v_32167 = v_2883;
assign v_32169 = v_32166 & v_32168;
assign v_32170 = v_32169;
assign v_32172 = v_29395;
assign v_32173 = v_2948;
assign v_32174 = v_32173;
assign v_32175 = v_32172 & v_32174;
assign v_32176 = v_32175;
assign v_32177 = v_32067 & v_32176;
assign v_32179 = v_32077 & v_32178;
assign v_32180 = v_32066 & v_32176;
assign v_32182 = v_32064 & v_32181;
assign v_32184 = v_32083 & v_32183;
assign v_32185 = v_32063 & v_32181;
assign v_32187 = v_32061 & v_32186;
assign v_32189 = v_32089 & v_32188;
assign v_32190 = v_32060 & v_32186;
assign v_32192 = v_32058 & v_32191;
assign v_32194 = v_32095 & v_32193;
assign v_32195 = v_32057 & v_32191;
assign v_32197 = v_32055 & v_32196;
assign v_32199 = v_32101 & v_32198;
assign v_32200 = v_32054 & v_32196;
assign v_32202 = v_32052 & v_32201;
assign v_32204 = v_32107 & v_32203;
assign v_32205 = v_32051 & v_32201;
assign v_32207 = v_32049 & v_32206;
assign v_32209 = v_32113 & v_32208;
assign v_32210 = v_32048 & v_32206;
assign v_32212 = v_32046 & v_32211;
assign v_32214 = v_32119 & v_32213;
assign v_32215 = v_32045 & v_32211;
assign v_32217 = v_32043 & v_32216;
assign v_32219 = v_32125 & v_32218;
assign v_32220 = v_32042 & v_32216;
assign v_32222 = v_32040 & v_32221;
assign v_32224 = v_32131 & v_32223;
assign v_32225 = v_32039 & v_32221;
assign v_32227 = v_32037 & v_32226;
assign v_32229 = v_32137 & v_32228;
assign v_32230 = v_32036 & v_32226;
assign v_32232 = v_32034 & v_32231;
assign v_32234 = v_32143 & v_32233;
assign v_32235 = v_32033 & v_32231;
assign v_32237 = v_32031 & v_32236;
assign v_32239 = v_32149 & v_32238;
assign v_32240 = v_32030 & v_32236;
assign v_32242 = v_32028 & v_32241;
assign v_32244 = v_32155 & v_32243;
assign v_32245 = v_32027 & v_32241;
assign v_32247 = v_32025 & v_32246;
assign v_32249 = v_32161 & v_32248;
assign v_32250 = v_32024 & v_32246;
assign v_32252 = v_32022 & v_32251;
assign v_32254 = v_32167 & v_32253;
assign v_32255 = v_32021 & v_32251;
assign v_32257 = v_32256;
assign v_32259 = v_32171 & v_32258;
assign v_32260 = v_32259;
assign v_32262 = v_32261;
assign v_32264 = ~v_3143;
assign v_32265 = ~v_29332;
assign v_32266 = v_29332;
assign v_32267 = ~v_3147;
assign v_32268 = ~v_29336;
assign v_32269 = v_29336;
assign v_32270 = ~v_3151;
assign v_32271 = ~v_29340;
assign v_32272 = v_29340;
assign v_32273 = ~v_3155;
assign v_32274 = ~v_29344;
assign v_32275 = v_29344;
assign v_32276 = ~v_29347;
assign v_32277 = ~v_3160;
assign v_32278 = v_3160;
assign v_32279 = ~v_29351;
assign v_32280 = ~v_3164;
assign v_32281 = v_3164;
assign v_32282 = ~v_29355;
assign v_32283 = ~v_3168;
assign v_32284 = v_3168;
assign v_32285 = ~v_29359;
assign v_32286 = ~v_3172;
assign v_32287 = v_3172;
assign v_32288 = ~v_29363;
assign v_32289 = ~v_3176;
assign v_32290 = v_3176;
assign v_32291 = ~v_29367;
assign v_32292 = ~v_3180;
assign v_32293 = v_3180;
assign v_32294 = ~v_29371;
assign v_32295 = ~v_3184;
assign v_32296 = v_3184;
assign v_32297 = ~v_29375;
assign v_32298 = ~v_3188;
assign v_32299 = v_3188;
assign v_32300 = ~v_29379;
assign v_32301 = ~v_3192;
assign v_32302 = v_3192;
assign v_32303 = ~v_29383;
assign v_32304 = ~v_3196;
assign v_32305 = v_3196;
assign v_32306 = ~v_29387;
assign v_32307 = ~v_3200;
assign v_32308 = v_3200;
assign v_32309 = ~v_29391;
assign v_32310 = ~v_3204;
assign v_32311 = v_3204;
assign v_32312 = ~v_29395;
assign v_32313 = ~v_3208;
assign v_32314 = v_32313;
assign v_32316 = v_32315;
assign v_32318 = v_32310 & v_32317;
assign v_32320 = v_29391;
assign v_32322 = v_32319 & v_32321;
assign v_32324 = v_32307 & v_32323;
assign v_32326 = v_29387;
assign v_32328 = v_32325 & v_32327;
assign v_32330 = v_32304 & v_32329;
assign v_32332 = v_29383;
assign v_32334 = v_32331 & v_32333;
assign v_32336 = v_32301 & v_32335;
assign v_32338 = v_29379;
assign v_32340 = v_32337 & v_32339;
assign v_32342 = v_32298 & v_32341;
assign v_32344 = v_29375;
assign v_32346 = v_32343 & v_32345;
assign v_32348 = v_32295 & v_32347;
assign v_32350 = v_29371;
assign v_32352 = v_32349 & v_32351;
assign v_32354 = v_32292 & v_32353;
assign v_32356 = v_29367;
assign v_32358 = v_32355 & v_32357;
assign v_32360 = v_32289 & v_32359;
assign v_32362 = v_29363;
assign v_32364 = v_32361 & v_32363;
assign v_32366 = v_32286 & v_32365;
assign v_32368 = v_29359;
assign v_32370 = v_32367 & v_32369;
assign v_32372 = v_32283 & v_32371;
assign v_32374 = v_29355;
assign v_32376 = v_32373 & v_32375;
assign v_32378 = v_32280 & v_32377;
assign v_32380 = v_29351;
assign v_32382 = v_32379 & v_32381;
assign v_32384 = v_32277 & v_32383;
assign v_32386 = v_29347;
assign v_32388 = v_32385 & v_32387;
assign v_32390 = v_32274 & v_32389;
assign v_32392 = v_3155;
assign v_32394 = v_32391 & v_32393;
assign v_32396 = v_32271 & v_32395;
assign v_32398 = v_3151;
assign v_32400 = v_32397 & v_32399;
assign v_32402 = v_32268 & v_32401;
assign v_32404 = v_3147;
assign v_32406 = v_32403 & v_32405;
assign v_32408 = v_32265 & v_32407;
assign v_32410 = v_3143;
assign v_32412 = v_32409 & v_32411;
assign v_32413 = v_32412;
assign v_32415 = v_29395;
assign v_32416 = v_3208;
assign v_32417 = v_32416;
assign v_32418 = v_32415 & v_32417;
assign v_32419 = v_32418;
assign v_32420 = v_32310 & v_32419;
assign v_32422 = v_32320 & v_32421;
assign v_32423 = v_32309 & v_32419;
assign v_32425 = v_32307 & v_32424;
assign v_32427 = v_32326 & v_32426;
assign v_32428 = v_32306 & v_32424;
assign v_32430 = v_32304 & v_32429;
assign v_32432 = v_32332 & v_32431;
assign v_32433 = v_32303 & v_32429;
assign v_32435 = v_32301 & v_32434;
assign v_32437 = v_32338 & v_32436;
assign v_32438 = v_32300 & v_32434;
assign v_32440 = v_32298 & v_32439;
assign v_32442 = v_32344 & v_32441;
assign v_32443 = v_32297 & v_32439;
assign v_32445 = v_32295 & v_32444;
assign v_32447 = v_32350 & v_32446;
assign v_32448 = v_32294 & v_32444;
assign v_32450 = v_32292 & v_32449;
assign v_32452 = v_32356 & v_32451;
assign v_32453 = v_32291 & v_32449;
assign v_32455 = v_32289 & v_32454;
assign v_32457 = v_32362 & v_32456;
assign v_32458 = v_32288 & v_32454;
assign v_32460 = v_32286 & v_32459;
assign v_32462 = v_32368 & v_32461;
assign v_32463 = v_32285 & v_32459;
assign v_32465 = v_32283 & v_32464;
assign v_32467 = v_32374 & v_32466;
assign v_32468 = v_32282 & v_32464;
assign v_32470 = v_32280 & v_32469;
assign v_32472 = v_32380 & v_32471;
assign v_32473 = v_32279 & v_32469;
assign v_32475 = v_32277 & v_32474;
assign v_32477 = v_32386 & v_32476;
assign v_32478 = v_32276 & v_32474;
assign v_32480 = v_32274 & v_32479;
assign v_32482 = v_32392 & v_32481;
assign v_32483 = v_32273 & v_32479;
assign v_32485 = v_32271 & v_32484;
assign v_32487 = v_32398 & v_32486;
assign v_32488 = v_32270 & v_32484;
assign v_32490 = v_32268 & v_32489;
assign v_32492 = v_32404 & v_32491;
assign v_32493 = v_32267 & v_32489;
assign v_32495 = v_32265 & v_32494;
assign v_32497 = v_32410 & v_32496;
assign v_32498 = v_32264 & v_32494;
assign v_32500 = v_32499;
assign v_32502 = v_32414 & v_32501;
assign v_32503 = v_32502;
assign v_32505 = v_32504;
assign v_32507 = ~v_3403;
assign v_32508 = ~v_29332;
assign v_32509 = v_29332;
assign v_32510 = ~v_3407;
assign v_32511 = ~v_29336;
assign v_32512 = v_29336;
assign v_32513 = ~v_3411;
assign v_32514 = ~v_29340;
assign v_32515 = v_29340;
assign v_32516 = ~v_3415;
assign v_32517 = ~v_29344;
assign v_32518 = v_29344;
assign v_32519 = ~v_29347;
assign v_32520 = ~v_3420;
assign v_32521 = v_3420;
assign v_32522 = ~v_29351;
assign v_32523 = ~v_3424;
assign v_32524 = v_3424;
assign v_32525 = ~v_29355;
assign v_32526 = ~v_3428;
assign v_32527 = v_3428;
assign v_32528 = ~v_29359;
assign v_32529 = ~v_3432;
assign v_32530 = v_3432;
assign v_32531 = ~v_29363;
assign v_32532 = ~v_3436;
assign v_32533 = v_3436;
assign v_32534 = ~v_29367;
assign v_32535 = ~v_3440;
assign v_32536 = v_3440;
assign v_32537 = ~v_29371;
assign v_32538 = ~v_3444;
assign v_32539 = v_3444;
assign v_32540 = ~v_29375;
assign v_32541 = ~v_3448;
assign v_32542 = v_3448;
assign v_32543 = ~v_29379;
assign v_32544 = ~v_3452;
assign v_32545 = v_3452;
assign v_32546 = ~v_29383;
assign v_32547 = ~v_3456;
assign v_32548 = v_3456;
assign v_32549 = ~v_29387;
assign v_32550 = ~v_3460;
assign v_32551 = v_3460;
assign v_32552 = ~v_29391;
assign v_32553 = ~v_3464;
assign v_32554 = v_3464;
assign v_32555 = ~v_29395;
assign v_32556 = ~v_3468;
assign v_32557 = v_32556;
assign v_32559 = v_32558;
assign v_32561 = v_32553 & v_32560;
assign v_32563 = v_29391;
assign v_32565 = v_32562 & v_32564;
assign v_32567 = v_32550 & v_32566;
assign v_32569 = v_29387;
assign v_32571 = v_32568 & v_32570;
assign v_32573 = v_32547 & v_32572;
assign v_32575 = v_29383;
assign v_32577 = v_32574 & v_32576;
assign v_32579 = v_32544 & v_32578;
assign v_32581 = v_29379;
assign v_32583 = v_32580 & v_32582;
assign v_32585 = v_32541 & v_32584;
assign v_32587 = v_29375;
assign v_32589 = v_32586 & v_32588;
assign v_32591 = v_32538 & v_32590;
assign v_32593 = v_29371;
assign v_32595 = v_32592 & v_32594;
assign v_32597 = v_32535 & v_32596;
assign v_32599 = v_29367;
assign v_32601 = v_32598 & v_32600;
assign v_32603 = v_32532 & v_32602;
assign v_32605 = v_29363;
assign v_32607 = v_32604 & v_32606;
assign v_32609 = v_32529 & v_32608;
assign v_32611 = v_29359;
assign v_32613 = v_32610 & v_32612;
assign v_32615 = v_32526 & v_32614;
assign v_32617 = v_29355;
assign v_32619 = v_32616 & v_32618;
assign v_32621 = v_32523 & v_32620;
assign v_32623 = v_29351;
assign v_32625 = v_32622 & v_32624;
assign v_32627 = v_32520 & v_32626;
assign v_32629 = v_29347;
assign v_32631 = v_32628 & v_32630;
assign v_32633 = v_32517 & v_32632;
assign v_32635 = v_3415;
assign v_32637 = v_32634 & v_32636;
assign v_32639 = v_32514 & v_32638;
assign v_32641 = v_3411;
assign v_32643 = v_32640 & v_32642;
assign v_32645 = v_32511 & v_32644;
assign v_32647 = v_3407;
assign v_32649 = v_32646 & v_32648;
assign v_32651 = v_32508 & v_32650;
assign v_32653 = v_3403;
assign v_32655 = v_32652 & v_32654;
assign v_32656 = v_32655;
assign v_32658 = v_29395;
assign v_32659 = v_3468;
assign v_32660 = v_32659;
assign v_32661 = v_32658 & v_32660;
assign v_32662 = v_32661;
assign v_32663 = v_32553 & v_32662;
assign v_32665 = v_32563 & v_32664;
assign v_32666 = v_32552 & v_32662;
assign v_32668 = v_32550 & v_32667;
assign v_32670 = v_32569 & v_32669;
assign v_32671 = v_32549 & v_32667;
assign v_32673 = v_32547 & v_32672;
assign v_32675 = v_32575 & v_32674;
assign v_32676 = v_32546 & v_32672;
assign v_32678 = v_32544 & v_32677;
assign v_32680 = v_32581 & v_32679;
assign v_32681 = v_32543 & v_32677;
assign v_32683 = v_32541 & v_32682;
assign v_32685 = v_32587 & v_32684;
assign v_32686 = v_32540 & v_32682;
assign v_32688 = v_32538 & v_32687;
assign v_32690 = v_32593 & v_32689;
assign v_32691 = v_32537 & v_32687;
assign v_32693 = v_32535 & v_32692;
assign v_32695 = v_32599 & v_32694;
assign v_32696 = v_32534 & v_32692;
assign v_32698 = v_32532 & v_32697;
assign v_32700 = v_32605 & v_32699;
assign v_32701 = v_32531 & v_32697;
assign v_32703 = v_32529 & v_32702;
assign v_32705 = v_32611 & v_32704;
assign v_32706 = v_32528 & v_32702;
assign v_32708 = v_32526 & v_32707;
assign v_32710 = v_32617 & v_32709;
assign v_32711 = v_32525 & v_32707;
assign v_32713 = v_32523 & v_32712;
assign v_32715 = v_32623 & v_32714;
assign v_32716 = v_32522 & v_32712;
assign v_32718 = v_32520 & v_32717;
assign v_32720 = v_32629 & v_32719;
assign v_32721 = v_32519 & v_32717;
assign v_32723 = v_32517 & v_32722;
assign v_32725 = v_32635 & v_32724;
assign v_32726 = v_32516 & v_32722;
assign v_32728 = v_32514 & v_32727;
assign v_32730 = v_32641 & v_32729;
assign v_32731 = v_32513 & v_32727;
assign v_32733 = v_32511 & v_32732;
assign v_32735 = v_32647 & v_32734;
assign v_32736 = v_32510 & v_32732;
assign v_32738 = v_32508 & v_32737;
assign v_32740 = v_32653 & v_32739;
assign v_32741 = v_32507 & v_32737;
assign v_32743 = v_32742;
assign v_32745 = v_32657 & v_32744;
assign v_32746 = v_32745;
assign v_32748 = v_32747;
assign v_32750 = ~v_3663;
assign v_32751 = ~v_29332;
assign v_32752 = v_29332;
assign v_32753 = ~v_3667;
assign v_32754 = ~v_29336;
assign v_32755 = v_29336;
assign v_32756 = ~v_3671;
assign v_32757 = ~v_29340;
assign v_32758 = v_29340;
assign v_32759 = ~v_3675;
assign v_32760 = ~v_29344;
assign v_32761 = v_29344;
assign v_32762 = ~v_29347;
assign v_32763 = ~v_3680;
assign v_32764 = v_3680;
assign v_32765 = ~v_29351;
assign v_32766 = ~v_3684;
assign v_32767 = v_3684;
assign v_32768 = ~v_29355;
assign v_32769 = ~v_3688;
assign v_32770 = v_3688;
assign v_32771 = ~v_29359;
assign v_32772 = ~v_3692;
assign v_32773 = v_3692;
assign v_32774 = ~v_29363;
assign v_32775 = ~v_3696;
assign v_32776 = v_3696;
assign v_32777 = ~v_29367;
assign v_32778 = ~v_3700;
assign v_32779 = v_3700;
assign v_32780 = ~v_29371;
assign v_32781 = ~v_3704;
assign v_32782 = v_3704;
assign v_32783 = ~v_29375;
assign v_32784 = ~v_3708;
assign v_32785 = v_3708;
assign v_32786 = ~v_29379;
assign v_32787 = ~v_3712;
assign v_32788 = v_3712;
assign v_32789 = ~v_29383;
assign v_32790 = ~v_3716;
assign v_32791 = v_3716;
assign v_32792 = ~v_29387;
assign v_32793 = ~v_3720;
assign v_32794 = v_3720;
assign v_32795 = ~v_29391;
assign v_32796 = ~v_3724;
assign v_32797 = v_3724;
assign v_32798 = ~v_29395;
assign v_32799 = ~v_3728;
assign v_32800 = v_32799;
assign v_32802 = v_32801;
assign v_32804 = v_32796 & v_32803;
assign v_32806 = v_29391;
assign v_32808 = v_32805 & v_32807;
assign v_32810 = v_32793 & v_32809;
assign v_32812 = v_29387;
assign v_32814 = v_32811 & v_32813;
assign v_32816 = v_32790 & v_32815;
assign v_32818 = v_29383;
assign v_32820 = v_32817 & v_32819;
assign v_32822 = v_32787 & v_32821;
assign v_32824 = v_29379;
assign v_32826 = v_32823 & v_32825;
assign v_32828 = v_32784 & v_32827;
assign v_32830 = v_29375;
assign v_32832 = v_32829 & v_32831;
assign v_32834 = v_32781 & v_32833;
assign v_32836 = v_29371;
assign v_32838 = v_32835 & v_32837;
assign v_32840 = v_32778 & v_32839;
assign v_32842 = v_29367;
assign v_32844 = v_32841 & v_32843;
assign v_32846 = v_32775 & v_32845;
assign v_32848 = v_29363;
assign v_32850 = v_32847 & v_32849;
assign v_32852 = v_32772 & v_32851;
assign v_32854 = v_29359;
assign v_32856 = v_32853 & v_32855;
assign v_32858 = v_32769 & v_32857;
assign v_32860 = v_29355;
assign v_32862 = v_32859 & v_32861;
assign v_32864 = v_32766 & v_32863;
assign v_32866 = v_29351;
assign v_32868 = v_32865 & v_32867;
assign v_32870 = v_32763 & v_32869;
assign v_32872 = v_29347;
assign v_32874 = v_32871 & v_32873;
assign v_32876 = v_32760 & v_32875;
assign v_32878 = v_3675;
assign v_32880 = v_32877 & v_32879;
assign v_32882 = v_32757 & v_32881;
assign v_32884 = v_3671;
assign v_32886 = v_32883 & v_32885;
assign v_32888 = v_32754 & v_32887;
assign v_32890 = v_3667;
assign v_32892 = v_32889 & v_32891;
assign v_32894 = v_32751 & v_32893;
assign v_32896 = v_3663;
assign v_32898 = v_32895 & v_32897;
assign v_32899 = v_32898;
assign v_32901 = v_29395;
assign v_32902 = v_3728;
assign v_32903 = v_32902;
assign v_32904 = v_32901 & v_32903;
assign v_32905 = v_32904;
assign v_32906 = v_32796 & v_32905;
assign v_32908 = v_32806 & v_32907;
assign v_32909 = v_32795 & v_32905;
assign v_32911 = v_32793 & v_32910;
assign v_32913 = v_32812 & v_32912;
assign v_32914 = v_32792 & v_32910;
assign v_32916 = v_32790 & v_32915;
assign v_32918 = v_32818 & v_32917;
assign v_32919 = v_32789 & v_32915;
assign v_32921 = v_32787 & v_32920;
assign v_32923 = v_32824 & v_32922;
assign v_32924 = v_32786 & v_32920;
assign v_32926 = v_32784 & v_32925;
assign v_32928 = v_32830 & v_32927;
assign v_32929 = v_32783 & v_32925;
assign v_32931 = v_32781 & v_32930;
assign v_32933 = v_32836 & v_32932;
assign v_32934 = v_32780 & v_32930;
assign v_32936 = v_32778 & v_32935;
assign v_32938 = v_32842 & v_32937;
assign v_32939 = v_32777 & v_32935;
assign v_32941 = v_32775 & v_32940;
assign v_32943 = v_32848 & v_32942;
assign v_32944 = v_32774 & v_32940;
assign v_32946 = v_32772 & v_32945;
assign v_32948 = v_32854 & v_32947;
assign v_32949 = v_32771 & v_32945;
assign v_32951 = v_32769 & v_32950;
assign v_32953 = v_32860 & v_32952;
assign v_32954 = v_32768 & v_32950;
assign v_32956 = v_32766 & v_32955;
assign v_32958 = v_32866 & v_32957;
assign v_32959 = v_32765 & v_32955;
assign v_32961 = v_32763 & v_32960;
assign v_32963 = v_32872 & v_32962;
assign v_32964 = v_32762 & v_32960;
assign v_32966 = v_32760 & v_32965;
assign v_32968 = v_32878 & v_32967;
assign v_32969 = v_32759 & v_32965;
assign v_32971 = v_32757 & v_32970;
assign v_32973 = v_32884 & v_32972;
assign v_32974 = v_32756 & v_32970;
assign v_32976 = v_32754 & v_32975;
assign v_32978 = v_32890 & v_32977;
assign v_32979 = v_32753 & v_32975;
assign v_32981 = v_32751 & v_32980;
assign v_32983 = v_32896 & v_32982;
assign v_32984 = v_32750 & v_32980;
assign v_32986 = v_32985;
assign v_32988 = v_32900 & v_32987;
assign v_32989 = v_32988;
assign v_32991 = v_32990;
assign v_32993 = ~v_3923;
assign v_32994 = ~v_29332;
assign v_32995 = v_29332;
assign v_32996 = ~v_3927;
assign v_32997 = ~v_29336;
assign v_32998 = v_29336;
assign v_32999 = ~v_3931;
assign v_33000 = ~v_29340;
assign v_33001 = v_29340;
assign v_33002 = ~v_3935;
assign v_33003 = ~v_29344;
assign v_33004 = v_29344;
assign v_33005 = ~v_29347;
assign v_33006 = ~v_3940;
assign v_33007 = v_3940;
assign v_33008 = ~v_29351;
assign v_33009 = ~v_3944;
assign v_33010 = v_3944;
assign v_33011 = ~v_29355;
assign v_33012 = ~v_3948;
assign v_33013 = v_3948;
assign v_33014 = ~v_29359;
assign v_33015 = ~v_3952;
assign v_33016 = v_3952;
assign v_33017 = ~v_29363;
assign v_33018 = ~v_3956;
assign v_33019 = v_3956;
assign v_33020 = ~v_29367;
assign v_33021 = ~v_3960;
assign v_33022 = v_3960;
assign v_33023 = ~v_29371;
assign v_33024 = ~v_3964;
assign v_33025 = v_3964;
assign v_33026 = ~v_29375;
assign v_33027 = ~v_3968;
assign v_33028 = v_3968;
assign v_33029 = ~v_29379;
assign v_33030 = ~v_3972;
assign v_33031 = v_3972;
assign v_33032 = ~v_29383;
assign v_33033 = ~v_3976;
assign v_33034 = v_3976;
assign v_33035 = ~v_29387;
assign v_33036 = ~v_3980;
assign v_33037 = v_3980;
assign v_33038 = ~v_29391;
assign v_33039 = ~v_3984;
assign v_33040 = v_3984;
assign v_33041 = ~v_29395;
assign v_33042 = ~v_3988;
assign v_33043 = v_33042;
assign v_33045 = v_33044;
assign v_33047 = v_33039 & v_33046;
assign v_33049 = v_29391;
assign v_33051 = v_33048 & v_33050;
assign v_33053 = v_33036 & v_33052;
assign v_33055 = v_29387;
assign v_33057 = v_33054 & v_33056;
assign v_33059 = v_33033 & v_33058;
assign v_33061 = v_29383;
assign v_33063 = v_33060 & v_33062;
assign v_33065 = v_33030 & v_33064;
assign v_33067 = v_29379;
assign v_33069 = v_33066 & v_33068;
assign v_33071 = v_33027 & v_33070;
assign v_33073 = v_29375;
assign v_33075 = v_33072 & v_33074;
assign v_33077 = v_33024 & v_33076;
assign v_33079 = v_29371;
assign v_33081 = v_33078 & v_33080;
assign v_33083 = v_33021 & v_33082;
assign v_33085 = v_29367;
assign v_33087 = v_33084 & v_33086;
assign v_33089 = v_33018 & v_33088;
assign v_33091 = v_29363;
assign v_33093 = v_33090 & v_33092;
assign v_33095 = v_33015 & v_33094;
assign v_33097 = v_29359;
assign v_33099 = v_33096 & v_33098;
assign v_33101 = v_33012 & v_33100;
assign v_33103 = v_29355;
assign v_33105 = v_33102 & v_33104;
assign v_33107 = v_33009 & v_33106;
assign v_33109 = v_29351;
assign v_33111 = v_33108 & v_33110;
assign v_33113 = v_33006 & v_33112;
assign v_33115 = v_29347;
assign v_33117 = v_33114 & v_33116;
assign v_33119 = v_33003 & v_33118;
assign v_33121 = v_3935;
assign v_33123 = v_33120 & v_33122;
assign v_33125 = v_33000 & v_33124;
assign v_33127 = v_3931;
assign v_33129 = v_33126 & v_33128;
assign v_33131 = v_32997 & v_33130;
assign v_33133 = v_3927;
assign v_33135 = v_33132 & v_33134;
assign v_33137 = v_32994 & v_33136;
assign v_33139 = v_3923;
assign v_33141 = v_33138 & v_33140;
assign v_33142 = v_33141;
assign v_33144 = v_29395;
assign v_33145 = v_3988;
assign v_33146 = v_33145;
assign v_33147 = v_33144 & v_33146;
assign v_33148 = v_33147;
assign v_33149 = v_33039 & v_33148;
assign v_33151 = v_33049 & v_33150;
assign v_33152 = v_33038 & v_33148;
assign v_33154 = v_33036 & v_33153;
assign v_33156 = v_33055 & v_33155;
assign v_33157 = v_33035 & v_33153;
assign v_33159 = v_33033 & v_33158;
assign v_33161 = v_33061 & v_33160;
assign v_33162 = v_33032 & v_33158;
assign v_33164 = v_33030 & v_33163;
assign v_33166 = v_33067 & v_33165;
assign v_33167 = v_33029 & v_33163;
assign v_33169 = v_33027 & v_33168;
assign v_33171 = v_33073 & v_33170;
assign v_33172 = v_33026 & v_33168;
assign v_33174 = v_33024 & v_33173;
assign v_33176 = v_33079 & v_33175;
assign v_33177 = v_33023 & v_33173;
assign v_33179 = v_33021 & v_33178;
assign v_33181 = v_33085 & v_33180;
assign v_33182 = v_33020 & v_33178;
assign v_33184 = v_33018 & v_33183;
assign v_33186 = v_33091 & v_33185;
assign v_33187 = v_33017 & v_33183;
assign v_33189 = v_33015 & v_33188;
assign v_33191 = v_33097 & v_33190;
assign v_33192 = v_33014 & v_33188;
assign v_33194 = v_33012 & v_33193;
assign v_33196 = v_33103 & v_33195;
assign v_33197 = v_33011 & v_33193;
assign v_33199 = v_33009 & v_33198;
assign v_33201 = v_33109 & v_33200;
assign v_33202 = v_33008 & v_33198;
assign v_33204 = v_33006 & v_33203;
assign v_33206 = v_33115 & v_33205;
assign v_33207 = v_33005 & v_33203;
assign v_33209 = v_33003 & v_33208;
assign v_33211 = v_33121 & v_33210;
assign v_33212 = v_33002 & v_33208;
assign v_33214 = v_33000 & v_33213;
assign v_33216 = v_33127 & v_33215;
assign v_33217 = v_32999 & v_33213;
assign v_33219 = v_32997 & v_33218;
assign v_33221 = v_33133 & v_33220;
assign v_33222 = v_32996 & v_33218;
assign v_33224 = v_32994 & v_33223;
assign v_33226 = v_33139 & v_33225;
assign v_33227 = v_32993 & v_33223;
assign v_33229 = v_33228;
assign v_33231 = v_33143 & v_33230;
assign v_33232 = v_33231;
assign v_33234 = v_33233;
assign v_33235 = ~v_4182;
assign v_33236 = ~v_29332;
assign v_33237 = v_29332;
assign v_33238 = ~v_4186;
assign v_33239 = ~v_29336;
assign v_33240 = v_29336;
assign v_33241 = ~v_4190;
assign v_33242 = ~v_29340;
assign v_33243 = v_29340;
assign v_33244 = ~v_4194;
assign v_33245 = ~v_29344;
assign v_33246 = v_29344;
assign v_33247 = ~v_29347;
assign v_33248 = ~v_4199;
assign v_33249 = v_4199;
assign v_33250 = ~v_29351;
assign v_33251 = ~v_4203;
assign v_33252 = v_4203;
assign v_33253 = ~v_29355;
assign v_33254 = ~v_4207;
assign v_33255 = v_4207;
assign v_33256 = ~v_29359;
assign v_33257 = ~v_4211;
assign v_33258 = v_4211;
assign v_33259 = ~v_29363;
assign v_33260 = ~v_4215;
assign v_33261 = v_4215;
assign v_33262 = ~v_29367;
assign v_33263 = ~v_4219;
assign v_33264 = v_4219;
assign v_33265 = ~v_29371;
assign v_33266 = ~v_4223;
assign v_33267 = v_4223;
assign v_33268 = ~v_29375;
assign v_33269 = ~v_4227;
assign v_33270 = v_4227;
assign v_33271 = ~v_29379;
assign v_33272 = ~v_4231;
assign v_33273 = v_4231;
assign v_33274 = ~v_29383;
assign v_33275 = ~v_4235;
assign v_33276 = v_4235;
assign v_33277 = ~v_29387;
assign v_33278 = ~v_4239;
assign v_33279 = v_4239;
assign v_33280 = ~v_29391;
assign v_33281 = ~v_4243;
assign v_33282 = v_4243;
assign v_33283 = ~v_29395;
assign v_33284 = ~v_4247;
assign v_33285 = v_33284;
assign v_33287 = v_33286;
assign v_33289 = v_33281 & v_33288;
assign v_33291 = v_29391;
assign v_33293 = v_33290 & v_33292;
assign v_33295 = v_33278 & v_33294;
assign v_33297 = v_29387;
assign v_33299 = v_33296 & v_33298;
assign v_33301 = v_33275 & v_33300;
assign v_33303 = v_29383;
assign v_33305 = v_33302 & v_33304;
assign v_33307 = v_33272 & v_33306;
assign v_33309 = v_29379;
assign v_33311 = v_33308 & v_33310;
assign v_33313 = v_33269 & v_33312;
assign v_33315 = v_29375;
assign v_33317 = v_33314 & v_33316;
assign v_33319 = v_33266 & v_33318;
assign v_33321 = v_29371;
assign v_33323 = v_33320 & v_33322;
assign v_33325 = v_33263 & v_33324;
assign v_33327 = v_29367;
assign v_33329 = v_33326 & v_33328;
assign v_33331 = v_33260 & v_33330;
assign v_33333 = v_29363;
assign v_33335 = v_33332 & v_33334;
assign v_33337 = v_33257 & v_33336;
assign v_33339 = v_29359;
assign v_33341 = v_33338 & v_33340;
assign v_33343 = v_33254 & v_33342;
assign v_33345 = v_29355;
assign v_33347 = v_33344 & v_33346;
assign v_33349 = v_33251 & v_33348;
assign v_33351 = v_29351;
assign v_33353 = v_33350 & v_33352;
assign v_33355 = v_33248 & v_33354;
assign v_33357 = v_29347;
assign v_33359 = v_33356 & v_33358;
assign v_33361 = v_33245 & v_33360;
assign v_33363 = v_4194;
assign v_33365 = v_33362 & v_33364;
assign v_33367 = v_33242 & v_33366;
assign v_33369 = v_4190;
assign v_33371 = v_33368 & v_33370;
assign v_33373 = v_33239 & v_33372;
assign v_33375 = v_4186;
assign v_33377 = v_33374 & v_33376;
assign v_33379 = v_33236 & v_33378;
assign v_33381 = v_4182;
assign v_33383 = v_33380 & v_33382;
assign v_33385 = ~v_33384;
assign v_33387 = v_29395;
assign v_33388 = v_4247;
assign v_33389 = v_33388;
assign v_33390 = v_33387 & v_33389;
assign v_33391 = v_33390;
assign v_33392 = v_33281 & v_33391;
assign v_33394 = v_33291 & v_33393;
assign v_33395 = v_33280 & v_33391;
assign v_33397 = v_33278 & v_33396;
assign v_33399 = v_33297 & v_33398;
assign v_33400 = v_33277 & v_33396;
assign v_33402 = v_33275 & v_33401;
assign v_33404 = v_33303 & v_33403;
assign v_33405 = v_33274 & v_33401;
assign v_33407 = v_33272 & v_33406;
assign v_33409 = v_33309 & v_33408;
assign v_33410 = v_33271 & v_33406;
assign v_33412 = v_33269 & v_33411;
assign v_33414 = v_33315 & v_33413;
assign v_33415 = v_33268 & v_33411;
assign v_33417 = v_33266 & v_33416;
assign v_33419 = v_33321 & v_33418;
assign v_33420 = v_33265 & v_33416;
assign v_33422 = v_33263 & v_33421;
assign v_33424 = v_33327 & v_33423;
assign v_33425 = v_33262 & v_33421;
assign v_33427 = v_33260 & v_33426;
assign v_33429 = v_33333 & v_33428;
assign v_33430 = v_33259 & v_33426;
assign v_33432 = v_33257 & v_33431;
assign v_33434 = v_33339 & v_33433;
assign v_33435 = v_33256 & v_33431;
assign v_33437 = v_33254 & v_33436;
assign v_33439 = v_33345 & v_33438;
assign v_33440 = v_33253 & v_33436;
assign v_33442 = v_33251 & v_33441;
assign v_33444 = v_33351 & v_33443;
assign v_33445 = v_33250 & v_33441;
assign v_33447 = v_33248 & v_33446;
assign v_33449 = v_33357 & v_33448;
assign v_33450 = v_33247 & v_33446;
assign v_33452 = v_33245 & v_33451;
assign v_33454 = v_33363 & v_33453;
assign v_33455 = v_33244 & v_33451;
assign v_33457 = v_33242 & v_33456;
assign v_33459 = v_33369 & v_33458;
assign v_33460 = v_33241 & v_33456;
assign v_33462 = v_33239 & v_33461;
assign v_33464 = v_33375 & v_33463;
assign v_33465 = v_33238 & v_33461;
assign v_33467 = v_33236 & v_33466;
assign v_33469 = v_33381 & v_33468;
assign v_33470 = v_33235 & v_33466;
assign v_33472 = v_33384;
assign v_33474 = v_33386 & v_33473;
assign v_33475 = v_33474;
assign v_33477 = v_33476;
assign v_33479 = ~v_6;
assign v_33481 = ~v_33480;
assign v_33482 = v_33480;
assign v_33483 = ~v_13;
assign v_33485 = ~v_33484;
assign v_33486 = v_33484;
assign v_33487 = ~v_18;
assign v_33489 = ~v_33488;
assign v_33490 = v_33488;
assign v_33491 = ~v_23;
assign v_33493 = ~v_33492;
assign v_33494 = v_33492;
assign v_33496 = ~v_33495;
assign v_33497 = ~v_30;
assign v_33498 = v_30;
assign v_33500 = ~v_33499;
assign v_33501 = ~v_35;
assign v_33502 = v_35;
assign v_33504 = ~v_33503;
assign v_33505 = ~v_40;
assign v_33506 = v_40;
assign v_33508 = ~v_33507;
assign v_33509 = ~v_45;
assign v_33510 = v_45;
assign v_33512 = ~v_33511;
assign v_33513 = ~v_50;
assign v_33514 = v_50;
assign v_33516 = ~v_33515;
assign v_33517 = ~v_55;
assign v_33518 = v_55;
assign v_33520 = ~v_33519;
assign v_33521 = ~v_60;
assign v_33522 = v_60;
assign v_33524 = ~v_33523;
assign v_33525 = ~v_65;
assign v_33526 = v_65;
assign v_33528 = ~v_33527;
assign v_33529 = ~v_70;
assign v_33530 = v_70;
assign v_33532 = ~v_33531;
assign v_33533 = ~v_75;
assign v_33534 = v_75;
assign v_33536 = ~v_33535;
assign v_33537 = ~v_80;
assign v_33538 = v_80;
assign v_33540 = ~v_33539;
assign v_33541 = ~v_85;
assign v_33542 = v_85;
assign v_33544 = ~v_33543;
assign v_33545 = ~v_90;
assign v_33546 = v_33545;
assign v_33548 = v_33547;
assign v_33550 = v_33541 & v_33549;
assign v_33552 = v_33539;
assign v_33554 = v_33551 & v_33553;
assign v_33556 = v_33537 & v_33555;
assign v_33558 = v_33535;
assign v_33560 = v_33557 & v_33559;
assign v_33562 = v_33533 & v_33561;
assign v_33564 = v_33531;
assign v_33566 = v_33563 & v_33565;
assign v_33568 = v_33529 & v_33567;
assign v_33570 = v_33527;
assign v_33572 = v_33569 & v_33571;
assign v_33574 = v_33525 & v_33573;
assign v_33576 = v_33523;
assign v_33578 = v_33575 & v_33577;
assign v_33580 = v_33521 & v_33579;
assign v_33582 = v_33519;
assign v_33584 = v_33581 & v_33583;
assign v_33586 = v_33517 & v_33585;
assign v_33588 = v_33515;
assign v_33590 = v_33587 & v_33589;
assign v_33592 = v_33513 & v_33591;
assign v_33594 = v_33511;
assign v_33596 = v_33593 & v_33595;
assign v_33598 = v_33509 & v_33597;
assign v_33600 = v_33507;
assign v_33602 = v_33599 & v_33601;
assign v_33604 = v_33505 & v_33603;
assign v_33606 = v_33503;
assign v_33608 = v_33605 & v_33607;
assign v_33610 = v_33501 & v_33609;
assign v_33612 = v_33499;
assign v_33614 = v_33611 & v_33613;
assign v_33616 = v_33497 & v_33615;
assign v_33618 = v_33495;
assign v_33620 = v_33617 & v_33619;
assign v_33622 = v_33493 & v_33621;
assign v_33624 = v_23;
assign v_33626 = v_33623 & v_33625;
assign v_33628 = v_33489 & v_33627;
assign v_33630 = v_18;
assign v_33632 = v_33629 & v_33631;
assign v_33634 = v_33485 & v_33633;
assign v_33636 = v_13;
assign v_33638 = v_33635 & v_33637;
assign v_33640 = v_33481 & v_33639;
assign v_33642 = v_6;
assign v_33644 = v_33641 & v_33643;
assign v_33645 = v_33644;
assign v_33647 = v_33543;
assign v_33648 = v_90;
assign v_33649 = v_33648;
assign v_33650 = v_33647 & v_33649;
assign v_33651 = v_33650;
assign v_33652 = v_33541 & v_33651;
assign v_33654 = v_33552 & v_33653;
assign v_33655 = v_33540 & v_33651;
assign v_33657 = v_33537 & v_33656;
assign v_33659 = v_33558 & v_33658;
assign v_33660 = v_33536 & v_33656;
assign v_33662 = v_33533 & v_33661;
assign v_33664 = v_33564 & v_33663;
assign v_33665 = v_33532 & v_33661;
assign v_33667 = v_33529 & v_33666;
assign v_33669 = v_33570 & v_33668;
assign v_33670 = v_33528 & v_33666;
assign v_33672 = v_33525 & v_33671;
assign v_33674 = v_33576 & v_33673;
assign v_33675 = v_33524 & v_33671;
assign v_33677 = v_33521 & v_33676;
assign v_33679 = v_33582 & v_33678;
assign v_33680 = v_33520 & v_33676;
assign v_33682 = v_33517 & v_33681;
assign v_33684 = v_33588 & v_33683;
assign v_33685 = v_33516 & v_33681;
assign v_33687 = v_33513 & v_33686;
assign v_33689 = v_33594 & v_33688;
assign v_33690 = v_33512 & v_33686;
assign v_33692 = v_33509 & v_33691;
assign v_33694 = v_33600 & v_33693;
assign v_33695 = v_33508 & v_33691;
assign v_33697 = v_33505 & v_33696;
assign v_33699 = v_33606 & v_33698;
assign v_33700 = v_33504 & v_33696;
assign v_33702 = v_33501 & v_33701;
assign v_33704 = v_33612 & v_33703;
assign v_33705 = v_33500 & v_33701;
assign v_33707 = v_33497 & v_33706;
assign v_33709 = v_33618 & v_33708;
assign v_33710 = v_33496 & v_33706;
assign v_33712 = v_33493 & v_33711;
assign v_33714 = v_33624 & v_33713;
assign v_33715 = v_33491 & v_33711;
assign v_33717 = v_33489 & v_33716;
assign v_33719 = v_33630 & v_33718;
assign v_33720 = v_33487 & v_33716;
assign v_33722 = v_33485 & v_33721;
assign v_33724 = v_33636 & v_33723;
assign v_33725 = v_33483 & v_33721;
assign v_33727 = v_33481 & v_33726;
assign v_33729 = v_33642 & v_33728;
assign v_33730 = v_33479 & v_33726;
assign v_33732 = v_33731;
assign v_33734 = v_33646 & v_33733;
assign v_33735 = v_33734;
assign v_33737 = v_33736;
assign v_33739 = ~v_283;
assign v_33740 = ~v_33480;
assign v_33741 = v_33480;
assign v_33742 = ~v_287;
assign v_33743 = ~v_33484;
assign v_33744 = v_33484;
assign v_33745 = ~v_291;
assign v_33746 = ~v_33488;
assign v_33747 = v_33488;
assign v_33748 = ~v_295;
assign v_33749 = ~v_33492;
assign v_33750 = v_33492;
assign v_33751 = ~v_33495;
assign v_33752 = ~v_300;
assign v_33753 = v_300;
assign v_33754 = ~v_33499;
assign v_33755 = ~v_304;
assign v_33756 = v_304;
assign v_33757 = ~v_33503;
assign v_33758 = ~v_308;
assign v_33759 = v_308;
assign v_33760 = ~v_33507;
assign v_33761 = ~v_312;
assign v_33762 = v_312;
assign v_33763 = ~v_33511;
assign v_33764 = ~v_316;
assign v_33765 = v_316;
assign v_33766 = ~v_33515;
assign v_33767 = ~v_320;
assign v_33768 = v_320;
assign v_33769 = ~v_33519;
assign v_33770 = ~v_324;
assign v_33771 = v_324;
assign v_33772 = ~v_33523;
assign v_33773 = ~v_328;
assign v_33774 = v_328;
assign v_33775 = ~v_33527;
assign v_33776 = ~v_332;
assign v_33777 = v_332;
assign v_33778 = ~v_33531;
assign v_33779 = ~v_336;
assign v_33780 = v_336;
assign v_33781 = ~v_33535;
assign v_33782 = ~v_340;
assign v_33783 = v_340;
assign v_33784 = ~v_33539;
assign v_33785 = ~v_344;
assign v_33786 = v_344;
assign v_33787 = ~v_33543;
assign v_33788 = ~v_348;
assign v_33789 = v_33788;
assign v_33791 = v_33790;
assign v_33793 = v_33785 & v_33792;
assign v_33795 = v_33539;
assign v_33797 = v_33794 & v_33796;
assign v_33799 = v_33782 & v_33798;
assign v_33801 = v_33535;
assign v_33803 = v_33800 & v_33802;
assign v_33805 = v_33779 & v_33804;
assign v_33807 = v_33531;
assign v_33809 = v_33806 & v_33808;
assign v_33811 = v_33776 & v_33810;
assign v_33813 = v_33527;
assign v_33815 = v_33812 & v_33814;
assign v_33817 = v_33773 & v_33816;
assign v_33819 = v_33523;
assign v_33821 = v_33818 & v_33820;
assign v_33823 = v_33770 & v_33822;
assign v_33825 = v_33519;
assign v_33827 = v_33824 & v_33826;
assign v_33829 = v_33767 & v_33828;
assign v_33831 = v_33515;
assign v_33833 = v_33830 & v_33832;
assign v_33835 = v_33764 & v_33834;
assign v_33837 = v_33511;
assign v_33839 = v_33836 & v_33838;
assign v_33841 = v_33761 & v_33840;
assign v_33843 = v_33507;
assign v_33845 = v_33842 & v_33844;
assign v_33847 = v_33758 & v_33846;
assign v_33849 = v_33503;
assign v_33851 = v_33848 & v_33850;
assign v_33853 = v_33755 & v_33852;
assign v_33855 = v_33499;
assign v_33857 = v_33854 & v_33856;
assign v_33859 = v_33752 & v_33858;
assign v_33861 = v_33495;
assign v_33863 = v_33860 & v_33862;
assign v_33865 = v_33749 & v_33864;
assign v_33867 = v_295;
assign v_33869 = v_33866 & v_33868;
assign v_33871 = v_33746 & v_33870;
assign v_33873 = v_291;
assign v_33875 = v_33872 & v_33874;
assign v_33877 = v_33743 & v_33876;
assign v_33879 = v_287;
assign v_33881 = v_33878 & v_33880;
assign v_33883 = v_33740 & v_33882;
assign v_33885 = v_283;
assign v_33887 = v_33884 & v_33886;
assign v_33888 = v_33887;
assign v_33890 = v_33543;
assign v_33891 = v_348;
assign v_33892 = v_33891;
assign v_33893 = v_33890 & v_33892;
assign v_33894 = v_33893;
assign v_33895 = v_33785 & v_33894;
assign v_33897 = v_33795 & v_33896;
assign v_33898 = v_33784 & v_33894;
assign v_33900 = v_33782 & v_33899;
assign v_33902 = v_33801 & v_33901;
assign v_33903 = v_33781 & v_33899;
assign v_33905 = v_33779 & v_33904;
assign v_33907 = v_33807 & v_33906;
assign v_33908 = v_33778 & v_33904;
assign v_33910 = v_33776 & v_33909;
assign v_33912 = v_33813 & v_33911;
assign v_33913 = v_33775 & v_33909;
assign v_33915 = v_33773 & v_33914;
assign v_33917 = v_33819 & v_33916;
assign v_33918 = v_33772 & v_33914;
assign v_33920 = v_33770 & v_33919;
assign v_33922 = v_33825 & v_33921;
assign v_33923 = v_33769 & v_33919;
assign v_33925 = v_33767 & v_33924;
assign v_33927 = v_33831 & v_33926;
assign v_33928 = v_33766 & v_33924;
assign v_33930 = v_33764 & v_33929;
assign v_33932 = v_33837 & v_33931;
assign v_33933 = v_33763 & v_33929;
assign v_33935 = v_33761 & v_33934;
assign v_33937 = v_33843 & v_33936;
assign v_33938 = v_33760 & v_33934;
assign v_33940 = v_33758 & v_33939;
assign v_33942 = v_33849 & v_33941;
assign v_33943 = v_33757 & v_33939;
assign v_33945 = v_33755 & v_33944;
assign v_33947 = v_33855 & v_33946;
assign v_33948 = v_33754 & v_33944;
assign v_33950 = v_33752 & v_33949;
assign v_33952 = v_33861 & v_33951;
assign v_33953 = v_33751 & v_33949;
assign v_33955 = v_33749 & v_33954;
assign v_33957 = v_33867 & v_33956;
assign v_33958 = v_33748 & v_33954;
assign v_33960 = v_33746 & v_33959;
assign v_33962 = v_33873 & v_33961;
assign v_33963 = v_33745 & v_33959;
assign v_33965 = v_33743 & v_33964;
assign v_33967 = v_33879 & v_33966;
assign v_33968 = v_33742 & v_33964;
assign v_33970 = v_33740 & v_33969;
assign v_33972 = v_33885 & v_33971;
assign v_33973 = v_33739 & v_33969;
assign v_33975 = v_33974;
assign v_33977 = v_33889 & v_33976;
assign v_33978 = v_33977;
assign v_33980 = v_33979;
assign v_33982 = ~v_543;
assign v_33983 = ~v_33480;
assign v_33984 = v_33480;
assign v_33985 = ~v_547;
assign v_33986 = ~v_33484;
assign v_33987 = v_33484;
assign v_33988 = ~v_551;
assign v_33989 = ~v_33488;
assign v_33990 = v_33488;
assign v_33991 = ~v_555;
assign v_33992 = ~v_33492;
assign v_33993 = v_33492;
assign v_33994 = ~v_33495;
assign v_33995 = ~v_560;
assign v_33996 = v_560;
assign v_33997 = ~v_33499;
assign v_33998 = ~v_564;
assign v_33999 = v_564;
assign v_34000 = ~v_33503;
assign v_34001 = ~v_568;
assign v_34002 = v_568;
assign v_34003 = ~v_33507;
assign v_34004 = ~v_572;
assign v_34005 = v_572;
assign v_34006 = ~v_33511;
assign v_34007 = ~v_576;
assign v_34008 = v_576;
assign v_34009 = ~v_33515;
assign v_34010 = ~v_580;
assign v_34011 = v_580;
assign v_34012 = ~v_33519;
assign v_34013 = ~v_584;
assign v_34014 = v_584;
assign v_34015 = ~v_33523;
assign v_34016 = ~v_588;
assign v_34017 = v_588;
assign v_34018 = ~v_33527;
assign v_34019 = ~v_592;
assign v_34020 = v_592;
assign v_34021 = ~v_33531;
assign v_34022 = ~v_596;
assign v_34023 = v_596;
assign v_34024 = ~v_33535;
assign v_34025 = ~v_600;
assign v_34026 = v_600;
assign v_34027 = ~v_33539;
assign v_34028 = ~v_604;
assign v_34029 = v_604;
assign v_34030 = ~v_33543;
assign v_34031 = ~v_608;
assign v_34032 = v_34031;
assign v_34034 = v_34033;
assign v_34036 = v_34028 & v_34035;
assign v_34038 = v_33539;
assign v_34040 = v_34037 & v_34039;
assign v_34042 = v_34025 & v_34041;
assign v_34044 = v_33535;
assign v_34046 = v_34043 & v_34045;
assign v_34048 = v_34022 & v_34047;
assign v_34050 = v_33531;
assign v_34052 = v_34049 & v_34051;
assign v_34054 = v_34019 & v_34053;
assign v_34056 = v_33527;
assign v_34058 = v_34055 & v_34057;
assign v_34060 = v_34016 & v_34059;
assign v_34062 = v_33523;
assign v_34064 = v_34061 & v_34063;
assign v_34066 = v_34013 & v_34065;
assign v_34068 = v_33519;
assign v_34070 = v_34067 & v_34069;
assign v_34072 = v_34010 & v_34071;
assign v_34074 = v_33515;
assign v_34076 = v_34073 & v_34075;
assign v_34078 = v_34007 & v_34077;
assign v_34080 = v_33511;
assign v_34082 = v_34079 & v_34081;
assign v_34084 = v_34004 & v_34083;
assign v_34086 = v_33507;
assign v_34088 = v_34085 & v_34087;
assign v_34090 = v_34001 & v_34089;
assign v_34092 = v_33503;
assign v_34094 = v_34091 & v_34093;
assign v_34096 = v_33998 & v_34095;
assign v_34098 = v_33499;
assign v_34100 = v_34097 & v_34099;
assign v_34102 = v_33995 & v_34101;
assign v_34104 = v_33495;
assign v_34106 = v_34103 & v_34105;
assign v_34108 = v_33992 & v_34107;
assign v_34110 = v_555;
assign v_34112 = v_34109 & v_34111;
assign v_34114 = v_33989 & v_34113;
assign v_34116 = v_551;
assign v_34118 = v_34115 & v_34117;
assign v_34120 = v_33986 & v_34119;
assign v_34122 = v_547;
assign v_34124 = v_34121 & v_34123;
assign v_34126 = v_33983 & v_34125;
assign v_34128 = v_543;
assign v_34130 = v_34127 & v_34129;
assign v_34131 = v_34130;
assign v_34133 = v_33543;
assign v_34134 = v_608;
assign v_34135 = v_34134;
assign v_34136 = v_34133 & v_34135;
assign v_34137 = v_34136;
assign v_34138 = v_34028 & v_34137;
assign v_34140 = v_34038 & v_34139;
assign v_34141 = v_34027 & v_34137;
assign v_34143 = v_34025 & v_34142;
assign v_34145 = v_34044 & v_34144;
assign v_34146 = v_34024 & v_34142;
assign v_34148 = v_34022 & v_34147;
assign v_34150 = v_34050 & v_34149;
assign v_34151 = v_34021 & v_34147;
assign v_34153 = v_34019 & v_34152;
assign v_34155 = v_34056 & v_34154;
assign v_34156 = v_34018 & v_34152;
assign v_34158 = v_34016 & v_34157;
assign v_34160 = v_34062 & v_34159;
assign v_34161 = v_34015 & v_34157;
assign v_34163 = v_34013 & v_34162;
assign v_34165 = v_34068 & v_34164;
assign v_34166 = v_34012 & v_34162;
assign v_34168 = v_34010 & v_34167;
assign v_34170 = v_34074 & v_34169;
assign v_34171 = v_34009 & v_34167;
assign v_34173 = v_34007 & v_34172;
assign v_34175 = v_34080 & v_34174;
assign v_34176 = v_34006 & v_34172;
assign v_34178 = v_34004 & v_34177;
assign v_34180 = v_34086 & v_34179;
assign v_34181 = v_34003 & v_34177;
assign v_34183 = v_34001 & v_34182;
assign v_34185 = v_34092 & v_34184;
assign v_34186 = v_34000 & v_34182;
assign v_34188 = v_33998 & v_34187;
assign v_34190 = v_34098 & v_34189;
assign v_34191 = v_33997 & v_34187;
assign v_34193 = v_33995 & v_34192;
assign v_34195 = v_34104 & v_34194;
assign v_34196 = v_33994 & v_34192;
assign v_34198 = v_33992 & v_34197;
assign v_34200 = v_34110 & v_34199;
assign v_34201 = v_33991 & v_34197;
assign v_34203 = v_33989 & v_34202;
assign v_34205 = v_34116 & v_34204;
assign v_34206 = v_33988 & v_34202;
assign v_34208 = v_33986 & v_34207;
assign v_34210 = v_34122 & v_34209;
assign v_34211 = v_33985 & v_34207;
assign v_34213 = v_33983 & v_34212;
assign v_34215 = v_34128 & v_34214;
assign v_34216 = v_33982 & v_34212;
assign v_34218 = v_34217;
assign v_34220 = v_34132 & v_34219;
assign v_34221 = v_34220;
assign v_34223 = v_34222;
assign v_34225 = ~v_803;
assign v_34226 = ~v_33480;
assign v_34227 = v_33480;
assign v_34228 = ~v_807;
assign v_34229 = ~v_33484;
assign v_34230 = v_33484;
assign v_34231 = ~v_811;
assign v_34232 = ~v_33488;
assign v_34233 = v_33488;
assign v_34234 = ~v_815;
assign v_34235 = ~v_33492;
assign v_34236 = v_33492;
assign v_34237 = ~v_33495;
assign v_34238 = ~v_820;
assign v_34239 = v_820;
assign v_34240 = ~v_33499;
assign v_34241 = ~v_824;
assign v_34242 = v_824;
assign v_34243 = ~v_33503;
assign v_34244 = ~v_828;
assign v_34245 = v_828;
assign v_34246 = ~v_33507;
assign v_34247 = ~v_832;
assign v_34248 = v_832;
assign v_34249 = ~v_33511;
assign v_34250 = ~v_836;
assign v_34251 = v_836;
assign v_34252 = ~v_33515;
assign v_34253 = ~v_840;
assign v_34254 = v_840;
assign v_34255 = ~v_33519;
assign v_34256 = ~v_844;
assign v_34257 = v_844;
assign v_34258 = ~v_33523;
assign v_34259 = ~v_848;
assign v_34260 = v_848;
assign v_34261 = ~v_33527;
assign v_34262 = ~v_852;
assign v_34263 = v_852;
assign v_34264 = ~v_33531;
assign v_34265 = ~v_856;
assign v_34266 = v_856;
assign v_34267 = ~v_33535;
assign v_34268 = ~v_860;
assign v_34269 = v_860;
assign v_34270 = ~v_33539;
assign v_34271 = ~v_864;
assign v_34272 = v_864;
assign v_34273 = ~v_33543;
assign v_34274 = ~v_868;
assign v_34275 = v_34274;
assign v_34277 = v_34276;
assign v_34279 = v_34271 & v_34278;
assign v_34281 = v_33539;
assign v_34283 = v_34280 & v_34282;
assign v_34285 = v_34268 & v_34284;
assign v_34287 = v_33535;
assign v_34289 = v_34286 & v_34288;
assign v_34291 = v_34265 & v_34290;
assign v_34293 = v_33531;
assign v_34295 = v_34292 & v_34294;
assign v_34297 = v_34262 & v_34296;
assign v_34299 = v_33527;
assign v_34301 = v_34298 & v_34300;
assign v_34303 = v_34259 & v_34302;
assign v_34305 = v_33523;
assign v_34307 = v_34304 & v_34306;
assign v_34309 = v_34256 & v_34308;
assign v_34311 = v_33519;
assign v_34313 = v_34310 & v_34312;
assign v_34315 = v_34253 & v_34314;
assign v_34317 = v_33515;
assign v_34319 = v_34316 & v_34318;
assign v_34321 = v_34250 & v_34320;
assign v_34323 = v_33511;
assign v_34325 = v_34322 & v_34324;
assign v_34327 = v_34247 & v_34326;
assign v_34329 = v_33507;
assign v_34331 = v_34328 & v_34330;
assign v_34333 = v_34244 & v_34332;
assign v_34335 = v_33503;
assign v_34337 = v_34334 & v_34336;
assign v_34339 = v_34241 & v_34338;
assign v_34341 = v_33499;
assign v_34343 = v_34340 & v_34342;
assign v_34345 = v_34238 & v_34344;
assign v_34347 = v_33495;
assign v_34349 = v_34346 & v_34348;
assign v_34351 = v_34235 & v_34350;
assign v_34353 = v_815;
assign v_34355 = v_34352 & v_34354;
assign v_34357 = v_34232 & v_34356;
assign v_34359 = v_811;
assign v_34361 = v_34358 & v_34360;
assign v_34363 = v_34229 & v_34362;
assign v_34365 = v_807;
assign v_34367 = v_34364 & v_34366;
assign v_34369 = v_34226 & v_34368;
assign v_34371 = v_803;
assign v_34373 = v_34370 & v_34372;
assign v_34374 = v_34373;
assign v_34376 = v_33543;
assign v_34377 = v_868;
assign v_34378 = v_34377;
assign v_34379 = v_34376 & v_34378;
assign v_34380 = v_34379;
assign v_34381 = v_34271 & v_34380;
assign v_34383 = v_34281 & v_34382;
assign v_34384 = v_34270 & v_34380;
assign v_34386 = v_34268 & v_34385;
assign v_34388 = v_34287 & v_34387;
assign v_34389 = v_34267 & v_34385;
assign v_34391 = v_34265 & v_34390;
assign v_34393 = v_34293 & v_34392;
assign v_34394 = v_34264 & v_34390;
assign v_34396 = v_34262 & v_34395;
assign v_34398 = v_34299 & v_34397;
assign v_34399 = v_34261 & v_34395;
assign v_34401 = v_34259 & v_34400;
assign v_34403 = v_34305 & v_34402;
assign v_34404 = v_34258 & v_34400;
assign v_34406 = v_34256 & v_34405;
assign v_34408 = v_34311 & v_34407;
assign v_34409 = v_34255 & v_34405;
assign v_34411 = v_34253 & v_34410;
assign v_34413 = v_34317 & v_34412;
assign v_34414 = v_34252 & v_34410;
assign v_34416 = v_34250 & v_34415;
assign v_34418 = v_34323 & v_34417;
assign v_34419 = v_34249 & v_34415;
assign v_34421 = v_34247 & v_34420;
assign v_34423 = v_34329 & v_34422;
assign v_34424 = v_34246 & v_34420;
assign v_34426 = v_34244 & v_34425;
assign v_34428 = v_34335 & v_34427;
assign v_34429 = v_34243 & v_34425;
assign v_34431 = v_34241 & v_34430;
assign v_34433 = v_34341 & v_34432;
assign v_34434 = v_34240 & v_34430;
assign v_34436 = v_34238 & v_34435;
assign v_34438 = v_34347 & v_34437;
assign v_34439 = v_34237 & v_34435;
assign v_34441 = v_34235 & v_34440;
assign v_34443 = v_34353 & v_34442;
assign v_34444 = v_34234 & v_34440;
assign v_34446 = v_34232 & v_34445;
assign v_34448 = v_34359 & v_34447;
assign v_34449 = v_34231 & v_34445;
assign v_34451 = v_34229 & v_34450;
assign v_34453 = v_34365 & v_34452;
assign v_34454 = v_34228 & v_34450;
assign v_34456 = v_34226 & v_34455;
assign v_34458 = v_34371 & v_34457;
assign v_34459 = v_34225 & v_34455;
assign v_34461 = v_34460;
assign v_34463 = v_34375 & v_34462;
assign v_34464 = v_34463;
assign v_34466 = v_34465;
assign v_34468 = ~v_1063;
assign v_34469 = ~v_33480;
assign v_34470 = v_33480;
assign v_34471 = ~v_1067;
assign v_34472 = ~v_33484;
assign v_34473 = v_33484;
assign v_34474 = ~v_1071;
assign v_34475 = ~v_33488;
assign v_34476 = v_33488;
assign v_34477 = ~v_1075;
assign v_34478 = ~v_33492;
assign v_34479 = v_33492;
assign v_34480 = ~v_33495;
assign v_34481 = ~v_1080;
assign v_34482 = v_1080;
assign v_34483 = ~v_33499;
assign v_34484 = ~v_1084;
assign v_34485 = v_1084;
assign v_34486 = ~v_33503;
assign v_34487 = ~v_1088;
assign v_34488 = v_1088;
assign v_34489 = ~v_33507;
assign v_34490 = ~v_1092;
assign v_34491 = v_1092;
assign v_34492 = ~v_33511;
assign v_34493 = ~v_1096;
assign v_34494 = v_1096;
assign v_34495 = ~v_33515;
assign v_34496 = ~v_1100;
assign v_34497 = v_1100;
assign v_34498 = ~v_33519;
assign v_34499 = ~v_1104;
assign v_34500 = v_1104;
assign v_34501 = ~v_33523;
assign v_34502 = ~v_1108;
assign v_34503 = v_1108;
assign v_34504 = ~v_33527;
assign v_34505 = ~v_1112;
assign v_34506 = v_1112;
assign v_34507 = ~v_33531;
assign v_34508 = ~v_1116;
assign v_34509 = v_1116;
assign v_34510 = ~v_33535;
assign v_34511 = ~v_1120;
assign v_34512 = v_1120;
assign v_34513 = ~v_33539;
assign v_34514 = ~v_1124;
assign v_34515 = v_1124;
assign v_34516 = ~v_33543;
assign v_34517 = ~v_1128;
assign v_34518 = v_34517;
assign v_34520 = v_34519;
assign v_34522 = v_34514 & v_34521;
assign v_34524 = v_33539;
assign v_34526 = v_34523 & v_34525;
assign v_34528 = v_34511 & v_34527;
assign v_34530 = v_33535;
assign v_34532 = v_34529 & v_34531;
assign v_34534 = v_34508 & v_34533;
assign v_34536 = v_33531;
assign v_34538 = v_34535 & v_34537;
assign v_34540 = v_34505 & v_34539;
assign v_34542 = v_33527;
assign v_34544 = v_34541 & v_34543;
assign v_34546 = v_34502 & v_34545;
assign v_34548 = v_33523;
assign v_34550 = v_34547 & v_34549;
assign v_34552 = v_34499 & v_34551;
assign v_34554 = v_33519;
assign v_34556 = v_34553 & v_34555;
assign v_34558 = v_34496 & v_34557;
assign v_34560 = v_33515;
assign v_34562 = v_34559 & v_34561;
assign v_34564 = v_34493 & v_34563;
assign v_34566 = v_33511;
assign v_34568 = v_34565 & v_34567;
assign v_34570 = v_34490 & v_34569;
assign v_34572 = v_33507;
assign v_34574 = v_34571 & v_34573;
assign v_34576 = v_34487 & v_34575;
assign v_34578 = v_33503;
assign v_34580 = v_34577 & v_34579;
assign v_34582 = v_34484 & v_34581;
assign v_34584 = v_33499;
assign v_34586 = v_34583 & v_34585;
assign v_34588 = v_34481 & v_34587;
assign v_34590 = v_33495;
assign v_34592 = v_34589 & v_34591;
assign v_34594 = v_34478 & v_34593;
assign v_34596 = v_1075;
assign v_34598 = v_34595 & v_34597;
assign v_34600 = v_34475 & v_34599;
assign v_34602 = v_1071;
assign v_34604 = v_34601 & v_34603;
assign v_34606 = v_34472 & v_34605;
assign v_34608 = v_1067;
assign v_34610 = v_34607 & v_34609;
assign v_34612 = v_34469 & v_34611;
assign v_34614 = v_1063;
assign v_34616 = v_34613 & v_34615;
assign v_34617 = v_34616;
assign v_34619 = v_33543;
assign v_34620 = v_1128;
assign v_34621 = v_34620;
assign v_34622 = v_34619 & v_34621;
assign v_34623 = v_34622;
assign v_34624 = v_34514 & v_34623;
assign v_34626 = v_34524 & v_34625;
assign v_34627 = v_34513 & v_34623;
assign v_34629 = v_34511 & v_34628;
assign v_34631 = v_34530 & v_34630;
assign v_34632 = v_34510 & v_34628;
assign v_34634 = v_34508 & v_34633;
assign v_34636 = v_34536 & v_34635;
assign v_34637 = v_34507 & v_34633;
assign v_34639 = v_34505 & v_34638;
assign v_34641 = v_34542 & v_34640;
assign v_34642 = v_34504 & v_34638;
assign v_34644 = v_34502 & v_34643;
assign v_34646 = v_34548 & v_34645;
assign v_34647 = v_34501 & v_34643;
assign v_34649 = v_34499 & v_34648;
assign v_34651 = v_34554 & v_34650;
assign v_34652 = v_34498 & v_34648;
assign v_34654 = v_34496 & v_34653;
assign v_34656 = v_34560 & v_34655;
assign v_34657 = v_34495 & v_34653;
assign v_34659 = v_34493 & v_34658;
assign v_34661 = v_34566 & v_34660;
assign v_34662 = v_34492 & v_34658;
assign v_34664 = v_34490 & v_34663;
assign v_34666 = v_34572 & v_34665;
assign v_34667 = v_34489 & v_34663;
assign v_34669 = v_34487 & v_34668;
assign v_34671 = v_34578 & v_34670;
assign v_34672 = v_34486 & v_34668;
assign v_34674 = v_34484 & v_34673;
assign v_34676 = v_34584 & v_34675;
assign v_34677 = v_34483 & v_34673;
assign v_34679 = v_34481 & v_34678;
assign v_34681 = v_34590 & v_34680;
assign v_34682 = v_34480 & v_34678;
assign v_34684 = v_34478 & v_34683;
assign v_34686 = v_34596 & v_34685;
assign v_34687 = v_34477 & v_34683;
assign v_34689 = v_34475 & v_34688;
assign v_34691 = v_34602 & v_34690;
assign v_34692 = v_34474 & v_34688;
assign v_34694 = v_34472 & v_34693;
assign v_34696 = v_34608 & v_34695;
assign v_34697 = v_34471 & v_34693;
assign v_34699 = v_34469 & v_34698;
assign v_34701 = v_34614 & v_34700;
assign v_34702 = v_34468 & v_34698;
assign v_34704 = v_34703;
assign v_34706 = v_34618 & v_34705;
assign v_34707 = v_34706;
assign v_34709 = v_34708;
assign v_34711 = ~v_1323;
assign v_34712 = ~v_33480;
assign v_34713 = v_33480;
assign v_34714 = ~v_1327;
assign v_34715 = ~v_33484;
assign v_34716 = v_33484;
assign v_34717 = ~v_1331;
assign v_34718 = ~v_33488;
assign v_34719 = v_33488;
assign v_34720 = ~v_1335;
assign v_34721 = ~v_33492;
assign v_34722 = v_33492;
assign v_34723 = ~v_33495;
assign v_34724 = ~v_1340;
assign v_34725 = v_1340;
assign v_34726 = ~v_33499;
assign v_34727 = ~v_1344;
assign v_34728 = v_1344;
assign v_34729 = ~v_33503;
assign v_34730 = ~v_1348;
assign v_34731 = v_1348;
assign v_34732 = ~v_33507;
assign v_34733 = ~v_1352;
assign v_34734 = v_1352;
assign v_34735 = ~v_33511;
assign v_34736 = ~v_1356;
assign v_34737 = v_1356;
assign v_34738 = ~v_33515;
assign v_34739 = ~v_1360;
assign v_34740 = v_1360;
assign v_34741 = ~v_33519;
assign v_34742 = ~v_1364;
assign v_34743 = v_1364;
assign v_34744 = ~v_33523;
assign v_34745 = ~v_1368;
assign v_34746 = v_1368;
assign v_34747 = ~v_33527;
assign v_34748 = ~v_1372;
assign v_34749 = v_1372;
assign v_34750 = ~v_33531;
assign v_34751 = ~v_1376;
assign v_34752 = v_1376;
assign v_34753 = ~v_33535;
assign v_34754 = ~v_1380;
assign v_34755 = v_1380;
assign v_34756 = ~v_33539;
assign v_34757 = ~v_1384;
assign v_34758 = v_1384;
assign v_34759 = ~v_33543;
assign v_34760 = ~v_1388;
assign v_34761 = v_34760;
assign v_34763 = v_34762;
assign v_34765 = v_34757 & v_34764;
assign v_34767 = v_33539;
assign v_34769 = v_34766 & v_34768;
assign v_34771 = v_34754 & v_34770;
assign v_34773 = v_33535;
assign v_34775 = v_34772 & v_34774;
assign v_34777 = v_34751 & v_34776;
assign v_34779 = v_33531;
assign v_34781 = v_34778 & v_34780;
assign v_34783 = v_34748 & v_34782;
assign v_34785 = v_33527;
assign v_34787 = v_34784 & v_34786;
assign v_34789 = v_34745 & v_34788;
assign v_34791 = v_33523;
assign v_34793 = v_34790 & v_34792;
assign v_34795 = v_34742 & v_34794;
assign v_34797 = v_33519;
assign v_34799 = v_34796 & v_34798;
assign v_34801 = v_34739 & v_34800;
assign v_34803 = v_33515;
assign v_34805 = v_34802 & v_34804;
assign v_34807 = v_34736 & v_34806;
assign v_34809 = v_33511;
assign v_34811 = v_34808 & v_34810;
assign v_34813 = v_34733 & v_34812;
assign v_34815 = v_33507;
assign v_34817 = v_34814 & v_34816;
assign v_34819 = v_34730 & v_34818;
assign v_34821 = v_33503;
assign v_34823 = v_34820 & v_34822;
assign v_34825 = v_34727 & v_34824;
assign v_34827 = v_33499;
assign v_34829 = v_34826 & v_34828;
assign v_34831 = v_34724 & v_34830;
assign v_34833 = v_33495;
assign v_34835 = v_34832 & v_34834;
assign v_34837 = v_34721 & v_34836;
assign v_34839 = v_1335;
assign v_34841 = v_34838 & v_34840;
assign v_34843 = v_34718 & v_34842;
assign v_34845 = v_1331;
assign v_34847 = v_34844 & v_34846;
assign v_34849 = v_34715 & v_34848;
assign v_34851 = v_1327;
assign v_34853 = v_34850 & v_34852;
assign v_34855 = v_34712 & v_34854;
assign v_34857 = v_1323;
assign v_34859 = v_34856 & v_34858;
assign v_34860 = v_34859;
assign v_34862 = v_33543;
assign v_34863 = v_1388;
assign v_34864 = v_34863;
assign v_34865 = v_34862 & v_34864;
assign v_34866 = v_34865;
assign v_34867 = v_34757 & v_34866;
assign v_34869 = v_34767 & v_34868;
assign v_34870 = v_34756 & v_34866;
assign v_34872 = v_34754 & v_34871;
assign v_34874 = v_34773 & v_34873;
assign v_34875 = v_34753 & v_34871;
assign v_34877 = v_34751 & v_34876;
assign v_34879 = v_34779 & v_34878;
assign v_34880 = v_34750 & v_34876;
assign v_34882 = v_34748 & v_34881;
assign v_34884 = v_34785 & v_34883;
assign v_34885 = v_34747 & v_34881;
assign v_34887 = v_34745 & v_34886;
assign v_34889 = v_34791 & v_34888;
assign v_34890 = v_34744 & v_34886;
assign v_34892 = v_34742 & v_34891;
assign v_34894 = v_34797 & v_34893;
assign v_34895 = v_34741 & v_34891;
assign v_34897 = v_34739 & v_34896;
assign v_34899 = v_34803 & v_34898;
assign v_34900 = v_34738 & v_34896;
assign v_34902 = v_34736 & v_34901;
assign v_34904 = v_34809 & v_34903;
assign v_34905 = v_34735 & v_34901;
assign v_34907 = v_34733 & v_34906;
assign v_34909 = v_34815 & v_34908;
assign v_34910 = v_34732 & v_34906;
assign v_34912 = v_34730 & v_34911;
assign v_34914 = v_34821 & v_34913;
assign v_34915 = v_34729 & v_34911;
assign v_34917 = v_34727 & v_34916;
assign v_34919 = v_34827 & v_34918;
assign v_34920 = v_34726 & v_34916;
assign v_34922 = v_34724 & v_34921;
assign v_34924 = v_34833 & v_34923;
assign v_34925 = v_34723 & v_34921;
assign v_34927 = v_34721 & v_34926;
assign v_34929 = v_34839 & v_34928;
assign v_34930 = v_34720 & v_34926;
assign v_34932 = v_34718 & v_34931;
assign v_34934 = v_34845 & v_34933;
assign v_34935 = v_34717 & v_34931;
assign v_34937 = v_34715 & v_34936;
assign v_34939 = v_34851 & v_34938;
assign v_34940 = v_34714 & v_34936;
assign v_34942 = v_34712 & v_34941;
assign v_34944 = v_34857 & v_34943;
assign v_34945 = v_34711 & v_34941;
assign v_34947 = v_34946;
assign v_34949 = v_34861 & v_34948;
assign v_34950 = v_34949;
assign v_34952 = v_34951;
assign v_34954 = ~v_1583;
assign v_34955 = ~v_33480;
assign v_34956 = v_33480;
assign v_34957 = ~v_1587;
assign v_34958 = ~v_33484;
assign v_34959 = v_33484;
assign v_34960 = ~v_1591;
assign v_34961 = ~v_33488;
assign v_34962 = v_33488;
assign v_34963 = ~v_1595;
assign v_34964 = ~v_33492;
assign v_34965 = v_33492;
assign v_34966 = ~v_33495;
assign v_34967 = ~v_1600;
assign v_34968 = v_1600;
assign v_34969 = ~v_33499;
assign v_34970 = ~v_1604;
assign v_34971 = v_1604;
assign v_34972 = ~v_33503;
assign v_34973 = ~v_1608;
assign v_34974 = v_1608;
assign v_34975 = ~v_33507;
assign v_34976 = ~v_1612;
assign v_34977 = v_1612;
assign v_34978 = ~v_33511;
assign v_34979 = ~v_1616;
assign v_34980 = v_1616;
assign v_34981 = ~v_33515;
assign v_34982 = ~v_1620;
assign v_34983 = v_1620;
assign v_34984 = ~v_33519;
assign v_34985 = ~v_1624;
assign v_34986 = v_1624;
assign v_34987 = ~v_33523;
assign v_34988 = ~v_1628;
assign v_34989 = v_1628;
assign v_34990 = ~v_33527;
assign v_34991 = ~v_1632;
assign v_34992 = v_1632;
assign v_34993 = ~v_33531;
assign v_34994 = ~v_1636;
assign v_34995 = v_1636;
assign v_34996 = ~v_33535;
assign v_34997 = ~v_1640;
assign v_34998 = v_1640;
assign v_34999 = ~v_33539;
assign v_35000 = ~v_1644;
assign v_35001 = v_1644;
assign v_35002 = ~v_33543;
assign v_35003 = ~v_1648;
assign v_35004 = v_35003;
assign v_35006 = v_35005;
assign v_35008 = v_35000 & v_35007;
assign v_35010 = v_33539;
assign v_35012 = v_35009 & v_35011;
assign v_35014 = v_34997 & v_35013;
assign v_35016 = v_33535;
assign v_35018 = v_35015 & v_35017;
assign v_35020 = v_34994 & v_35019;
assign v_35022 = v_33531;
assign v_35024 = v_35021 & v_35023;
assign v_35026 = v_34991 & v_35025;
assign v_35028 = v_33527;
assign v_35030 = v_35027 & v_35029;
assign v_35032 = v_34988 & v_35031;
assign v_35034 = v_33523;
assign v_35036 = v_35033 & v_35035;
assign v_35038 = v_34985 & v_35037;
assign v_35040 = v_33519;
assign v_35042 = v_35039 & v_35041;
assign v_35044 = v_34982 & v_35043;
assign v_35046 = v_33515;
assign v_35048 = v_35045 & v_35047;
assign v_35050 = v_34979 & v_35049;
assign v_35052 = v_33511;
assign v_35054 = v_35051 & v_35053;
assign v_35056 = v_34976 & v_35055;
assign v_35058 = v_33507;
assign v_35060 = v_35057 & v_35059;
assign v_35062 = v_34973 & v_35061;
assign v_35064 = v_33503;
assign v_35066 = v_35063 & v_35065;
assign v_35068 = v_34970 & v_35067;
assign v_35070 = v_33499;
assign v_35072 = v_35069 & v_35071;
assign v_35074 = v_34967 & v_35073;
assign v_35076 = v_33495;
assign v_35078 = v_35075 & v_35077;
assign v_35080 = v_34964 & v_35079;
assign v_35082 = v_1595;
assign v_35084 = v_35081 & v_35083;
assign v_35086 = v_34961 & v_35085;
assign v_35088 = v_1591;
assign v_35090 = v_35087 & v_35089;
assign v_35092 = v_34958 & v_35091;
assign v_35094 = v_1587;
assign v_35096 = v_35093 & v_35095;
assign v_35098 = v_34955 & v_35097;
assign v_35100 = v_1583;
assign v_35102 = v_35099 & v_35101;
assign v_35103 = v_35102;
assign v_35105 = v_33543;
assign v_35106 = v_1648;
assign v_35107 = v_35106;
assign v_35108 = v_35105 & v_35107;
assign v_35109 = v_35108;
assign v_35110 = v_35000 & v_35109;
assign v_35112 = v_35010 & v_35111;
assign v_35113 = v_34999 & v_35109;
assign v_35115 = v_34997 & v_35114;
assign v_35117 = v_35016 & v_35116;
assign v_35118 = v_34996 & v_35114;
assign v_35120 = v_34994 & v_35119;
assign v_35122 = v_35022 & v_35121;
assign v_35123 = v_34993 & v_35119;
assign v_35125 = v_34991 & v_35124;
assign v_35127 = v_35028 & v_35126;
assign v_35128 = v_34990 & v_35124;
assign v_35130 = v_34988 & v_35129;
assign v_35132 = v_35034 & v_35131;
assign v_35133 = v_34987 & v_35129;
assign v_35135 = v_34985 & v_35134;
assign v_35137 = v_35040 & v_35136;
assign v_35138 = v_34984 & v_35134;
assign v_35140 = v_34982 & v_35139;
assign v_35142 = v_35046 & v_35141;
assign v_35143 = v_34981 & v_35139;
assign v_35145 = v_34979 & v_35144;
assign v_35147 = v_35052 & v_35146;
assign v_35148 = v_34978 & v_35144;
assign v_35150 = v_34976 & v_35149;
assign v_35152 = v_35058 & v_35151;
assign v_35153 = v_34975 & v_35149;
assign v_35155 = v_34973 & v_35154;
assign v_35157 = v_35064 & v_35156;
assign v_35158 = v_34972 & v_35154;
assign v_35160 = v_34970 & v_35159;
assign v_35162 = v_35070 & v_35161;
assign v_35163 = v_34969 & v_35159;
assign v_35165 = v_34967 & v_35164;
assign v_35167 = v_35076 & v_35166;
assign v_35168 = v_34966 & v_35164;
assign v_35170 = v_34964 & v_35169;
assign v_35172 = v_35082 & v_35171;
assign v_35173 = v_34963 & v_35169;
assign v_35175 = v_34961 & v_35174;
assign v_35177 = v_35088 & v_35176;
assign v_35178 = v_34960 & v_35174;
assign v_35180 = v_34958 & v_35179;
assign v_35182 = v_35094 & v_35181;
assign v_35183 = v_34957 & v_35179;
assign v_35185 = v_34955 & v_35184;
assign v_35187 = v_35100 & v_35186;
assign v_35188 = v_34954 & v_35184;
assign v_35190 = v_35189;
assign v_35192 = v_35104 & v_35191;
assign v_35193 = v_35192;
assign v_35195 = v_35194;
assign v_35197 = ~v_1843;
assign v_35198 = ~v_33480;
assign v_35199 = v_33480;
assign v_35200 = ~v_1847;
assign v_35201 = ~v_33484;
assign v_35202 = v_33484;
assign v_35203 = ~v_1851;
assign v_35204 = ~v_33488;
assign v_35205 = v_33488;
assign v_35206 = ~v_1855;
assign v_35207 = ~v_33492;
assign v_35208 = v_33492;
assign v_35209 = ~v_33495;
assign v_35210 = ~v_1860;
assign v_35211 = v_1860;
assign v_35212 = ~v_33499;
assign v_35213 = ~v_1864;
assign v_35214 = v_1864;
assign v_35215 = ~v_33503;
assign v_35216 = ~v_1868;
assign v_35217 = v_1868;
assign v_35218 = ~v_33507;
assign v_35219 = ~v_1872;
assign v_35220 = v_1872;
assign v_35221 = ~v_33511;
assign v_35222 = ~v_1876;
assign v_35223 = v_1876;
assign v_35224 = ~v_33515;
assign v_35225 = ~v_1880;
assign v_35226 = v_1880;
assign v_35227 = ~v_33519;
assign v_35228 = ~v_1884;
assign v_35229 = v_1884;
assign v_35230 = ~v_33523;
assign v_35231 = ~v_1888;
assign v_35232 = v_1888;
assign v_35233 = ~v_33527;
assign v_35234 = ~v_1892;
assign v_35235 = v_1892;
assign v_35236 = ~v_33531;
assign v_35237 = ~v_1896;
assign v_35238 = v_1896;
assign v_35239 = ~v_33535;
assign v_35240 = ~v_1900;
assign v_35241 = v_1900;
assign v_35242 = ~v_33539;
assign v_35243 = ~v_1904;
assign v_35244 = v_1904;
assign v_35245 = ~v_33543;
assign v_35246 = ~v_1908;
assign v_35247 = v_35246;
assign v_35249 = v_35248;
assign v_35251 = v_35243 & v_35250;
assign v_35253 = v_33539;
assign v_35255 = v_35252 & v_35254;
assign v_35257 = v_35240 & v_35256;
assign v_35259 = v_33535;
assign v_35261 = v_35258 & v_35260;
assign v_35263 = v_35237 & v_35262;
assign v_35265 = v_33531;
assign v_35267 = v_35264 & v_35266;
assign v_35269 = v_35234 & v_35268;
assign v_35271 = v_33527;
assign v_35273 = v_35270 & v_35272;
assign v_35275 = v_35231 & v_35274;
assign v_35277 = v_33523;
assign v_35279 = v_35276 & v_35278;
assign v_35281 = v_35228 & v_35280;
assign v_35283 = v_33519;
assign v_35285 = v_35282 & v_35284;
assign v_35287 = v_35225 & v_35286;
assign v_35289 = v_33515;
assign v_35291 = v_35288 & v_35290;
assign v_35293 = v_35222 & v_35292;
assign v_35295 = v_33511;
assign v_35297 = v_35294 & v_35296;
assign v_35299 = v_35219 & v_35298;
assign v_35301 = v_33507;
assign v_35303 = v_35300 & v_35302;
assign v_35305 = v_35216 & v_35304;
assign v_35307 = v_33503;
assign v_35309 = v_35306 & v_35308;
assign v_35311 = v_35213 & v_35310;
assign v_35313 = v_33499;
assign v_35315 = v_35312 & v_35314;
assign v_35317 = v_35210 & v_35316;
assign v_35319 = v_33495;
assign v_35321 = v_35318 & v_35320;
assign v_35323 = v_35207 & v_35322;
assign v_35325 = v_1855;
assign v_35327 = v_35324 & v_35326;
assign v_35329 = v_35204 & v_35328;
assign v_35331 = v_1851;
assign v_35333 = v_35330 & v_35332;
assign v_35335 = v_35201 & v_35334;
assign v_35337 = v_1847;
assign v_35339 = v_35336 & v_35338;
assign v_35341 = v_35198 & v_35340;
assign v_35343 = v_1843;
assign v_35345 = v_35342 & v_35344;
assign v_35346 = v_35345;
assign v_35348 = v_33543;
assign v_35349 = v_1908;
assign v_35350 = v_35349;
assign v_35351 = v_35348 & v_35350;
assign v_35352 = v_35351;
assign v_35353 = v_35243 & v_35352;
assign v_35355 = v_35253 & v_35354;
assign v_35356 = v_35242 & v_35352;
assign v_35358 = v_35240 & v_35357;
assign v_35360 = v_35259 & v_35359;
assign v_35361 = v_35239 & v_35357;
assign v_35363 = v_35237 & v_35362;
assign v_35365 = v_35265 & v_35364;
assign v_35366 = v_35236 & v_35362;
assign v_35368 = v_35234 & v_35367;
assign v_35370 = v_35271 & v_35369;
assign v_35371 = v_35233 & v_35367;
assign v_35373 = v_35231 & v_35372;
assign v_35375 = v_35277 & v_35374;
assign v_35376 = v_35230 & v_35372;
assign v_35378 = v_35228 & v_35377;
assign v_35380 = v_35283 & v_35379;
assign v_35381 = v_35227 & v_35377;
assign v_35383 = v_35225 & v_35382;
assign v_35385 = v_35289 & v_35384;
assign v_35386 = v_35224 & v_35382;
assign v_35388 = v_35222 & v_35387;
assign v_35390 = v_35295 & v_35389;
assign v_35391 = v_35221 & v_35387;
assign v_35393 = v_35219 & v_35392;
assign v_35395 = v_35301 & v_35394;
assign v_35396 = v_35218 & v_35392;
assign v_35398 = v_35216 & v_35397;
assign v_35400 = v_35307 & v_35399;
assign v_35401 = v_35215 & v_35397;
assign v_35403 = v_35213 & v_35402;
assign v_35405 = v_35313 & v_35404;
assign v_35406 = v_35212 & v_35402;
assign v_35408 = v_35210 & v_35407;
assign v_35410 = v_35319 & v_35409;
assign v_35411 = v_35209 & v_35407;
assign v_35413 = v_35207 & v_35412;
assign v_35415 = v_35325 & v_35414;
assign v_35416 = v_35206 & v_35412;
assign v_35418 = v_35204 & v_35417;
assign v_35420 = v_35331 & v_35419;
assign v_35421 = v_35203 & v_35417;
assign v_35423 = v_35201 & v_35422;
assign v_35425 = v_35337 & v_35424;
assign v_35426 = v_35200 & v_35422;
assign v_35428 = v_35198 & v_35427;
assign v_35430 = v_35343 & v_35429;
assign v_35431 = v_35197 & v_35427;
assign v_35433 = v_35432;
assign v_35435 = v_35347 & v_35434;
assign v_35436 = v_35435;
assign v_35438 = v_35437;
assign v_35440 = ~v_2103;
assign v_35441 = ~v_33480;
assign v_35442 = v_33480;
assign v_35443 = ~v_2107;
assign v_35444 = ~v_33484;
assign v_35445 = v_33484;
assign v_35446 = ~v_2111;
assign v_35447 = ~v_33488;
assign v_35448 = v_33488;
assign v_35449 = ~v_2115;
assign v_35450 = ~v_33492;
assign v_35451 = v_33492;
assign v_35452 = ~v_33495;
assign v_35453 = ~v_2120;
assign v_35454 = v_2120;
assign v_35455 = ~v_33499;
assign v_35456 = ~v_2124;
assign v_35457 = v_2124;
assign v_35458 = ~v_33503;
assign v_35459 = ~v_2128;
assign v_35460 = v_2128;
assign v_35461 = ~v_33507;
assign v_35462 = ~v_2132;
assign v_35463 = v_2132;
assign v_35464 = ~v_33511;
assign v_35465 = ~v_2136;
assign v_35466 = v_2136;
assign v_35467 = ~v_33515;
assign v_35468 = ~v_2140;
assign v_35469 = v_2140;
assign v_35470 = ~v_33519;
assign v_35471 = ~v_2144;
assign v_35472 = v_2144;
assign v_35473 = ~v_33523;
assign v_35474 = ~v_2148;
assign v_35475 = v_2148;
assign v_35476 = ~v_33527;
assign v_35477 = ~v_2152;
assign v_35478 = v_2152;
assign v_35479 = ~v_33531;
assign v_35480 = ~v_2156;
assign v_35481 = v_2156;
assign v_35482 = ~v_33535;
assign v_35483 = ~v_2160;
assign v_35484 = v_2160;
assign v_35485 = ~v_33539;
assign v_35486 = ~v_2164;
assign v_35487 = v_2164;
assign v_35488 = ~v_33543;
assign v_35489 = ~v_2168;
assign v_35490 = v_35489;
assign v_35492 = v_35491;
assign v_35494 = v_35486 & v_35493;
assign v_35496 = v_33539;
assign v_35498 = v_35495 & v_35497;
assign v_35500 = v_35483 & v_35499;
assign v_35502 = v_33535;
assign v_35504 = v_35501 & v_35503;
assign v_35506 = v_35480 & v_35505;
assign v_35508 = v_33531;
assign v_35510 = v_35507 & v_35509;
assign v_35512 = v_35477 & v_35511;
assign v_35514 = v_33527;
assign v_35516 = v_35513 & v_35515;
assign v_35518 = v_35474 & v_35517;
assign v_35520 = v_33523;
assign v_35522 = v_35519 & v_35521;
assign v_35524 = v_35471 & v_35523;
assign v_35526 = v_33519;
assign v_35528 = v_35525 & v_35527;
assign v_35530 = v_35468 & v_35529;
assign v_35532 = v_33515;
assign v_35534 = v_35531 & v_35533;
assign v_35536 = v_35465 & v_35535;
assign v_35538 = v_33511;
assign v_35540 = v_35537 & v_35539;
assign v_35542 = v_35462 & v_35541;
assign v_35544 = v_33507;
assign v_35546 = v_35543 & v_35545;
assign v_35548 = v_35459 & v_35547;
assign v_35550 = v_33503;
assign v_35552 = v_35549 & v_35551;
assign v_35554 = v_35456 & v_35553;
assign v_35556 = v_33499;
assign v_35558 = v_35555 & v_35557;
assign v_35560 = v_35453 & v_35559;
assign v_35562 = v_33495;
assign v_35564 = v_35561 & v_35563;
assign v_35566 = v_35450 & v_35565;
assign v_35568 = v_2115;
assign v_35570 = v_35567 & v_35569;
assign v_35572 = v_35447 & v_35571;
assign v_35574 = v_2111;
assign v_35576 = v_35573 & v_35575;
assign v_35578 = v_35444 & v_35577;
assign v_35580 = v_2107;
assign v_35582 = v_35579 & v_35581;
assign v_35584 = v_35441 & v_35583;
assign v_35586 = v_2103;
assign v_35588 = v_35585 & v_35587;
assign v_35589 = v_35588;
assign v_35591 = v_33543;
assign v_35592 = v_2168;
assign v_35593 = v_35592;
assign v_35594 = v_35591 & v_35593;
assign v_35595 = v_35594;
assign v_35596 = v_35486 & v_35595;
assign v_35598 = v_35496 & v_35597;
assign v_35599 = v_35485 & v_35595;
assign v_35601 = v_35483 & v_35600;
assign v_35603 = v_35502 & v_35602;
assign v_35604 = v_35482 & v_35600;
assign v_35606 = v_35480 & v_35605;
assign v_35608 = v_35508 & v_35607;
assign v_35609 = v_35479 & v_35605;
assign v_35611 = v_35477 & v_35610;
assign v_35613 = v_35514 & v_35612;
assign v_35614 = v_35476 & v_35610;
assign v_35616 = v_35474 & v_35615;
assign v_35618 = v_35520 & v_35617;
assign v_35619 = v_35473 & v_35615;
assign v_35621 = v_35471 & v_35620;
assign v_35623 = v_35526 & v_35622;
assign v_35624 = v_35470 & v_35620;
assign v_35626 = v_35468 & v_35625;
assign v_35628 = v_35532 & v_35627;
assign v_35629 = v_35467 & v_35625;
assign v_35631 = v_35465 & v_35630;
assign v_35633 = v_35538 & v_35632;
assign v_35634 = v_35464 & v_35630;
assign v_35636 = v_35462 & v_35635;
assign v_35638 = v_35544 & v_35637;
assign v_35639 = v_35461 & v_35635;
assign v_35641 = v_35459 & v_35640;
assign v_35643 = v_35550 & v_35642;
assign v_35644 = v_35458 & v_35640;
assign v_35646 = v_35456 & v_35645;
assign v_35648 = v_35556 & v_35647;
assign v_35649 = v_35455 & v_35645;
assign v_35651 = v_35453 & v_35650;
assign v_35653 = v_35562 & v_35652;
assign v_35654 = v_35452 & v_35650;
assign v_35656 = v_35450 & v_35655;
assign v_35658 = v_35568 & v_35657;
assign v_35659 = v_35449 & v_35655;
assign v_35661 = v_35447 & v_35660;
assign v_35663 = v_35574 & v_35662;
assign v_35664 = v_35446 & v_35660;
assign v_35666 = v_35444 & v_35665;
assign v_35668 = v_35580 & v_35667;
assign v_35669 = v_35443 & v_35665;
assign v_35671 = v_35441 & v_35670;
assign v_35673 = v_35586 & v_35672;
assign v_35674 = v_35440 & v_35670;
assign v_35676 = v_35675;
assign v_35678 = v_35590 & v_35677;
assign v_35679 = v_35678;
assign v_35681 = v_35680;
assign v_35683 = ~v_2363;
assign v_35684 = ~v_33480;
assign v_35685 = v_33480;
assign v_35686 = ~v_2367;
assign v_35687 = ~v_33484;
assign v_35688 = v_33484;
assign v_35689 = ~v_2371;
assign v_35690 = ~v_33488;
assign v_35691 = v_33488;
assign v_35692 = ~v_2375;
assign v_35693 = ~v_33492;
assign v_35694 = v_33492;
assign v_35695 = ~v_33495;
assign v_35696 = ~v_2380;
assign v_35697 = v_2380;
assign v_35698 = ~v_33499;
assign v_35699 = ~v_2384;
assign v_35700 = v_2384;
assign v_35701 = ~v_33503;
assign v_35702 = ~v_2388;
assign v_35703 = v_2388;
assign v_35704 = ~v_33507;
assign v_35705 = ~v_2392;
assign v_35706 = v_2392;
assign v_35707 = ~v_33511;
assign v_35708 = ~v_2396;
assign v_35709 = v_2396;
assign v_35710 = ~v_33515;
assign v_35711 = ~v_2400;
assign v_35712 = v_2400;
assign v_35713 = ~v_33519;
assign v_35714 = ~v_2404;
assign v_35715 = v_2404;
assign v_35716 = ~v_33523;
assign v_35717 = ~v_2408;
assign v_35718 = v_2408;
assign v_35719 = ~v_33527;
assign v_35720 = ~v_2412;
assign v_35721 = v_2412;
assign v_35722 = ~v_33531;
assign v_35723 = ~v_2416;
assign v_35724 = v_2416;
assign v_35725 = ~v_33535;
assign v_35726 = ~v_2420;
assign v_35727 = v_2420;
assign v_35728 = ~v_33539;
assign v_35729 = ~v_2424;
assign v_35730 = v_2424;
assign v_35731 = ~v_33543;
assign v_35732 = ~v_2428;
assign v_35733 = v_35732;
assign v_35735 = v_35734;
assign v_35737 = v_35729 & v_35736;
assign v_35739 = v_33539;
assign v_35741 = v_35738 & v_35740;
assign v_35743 = v_35726 & v_35742;
assign v_35745 = v_33535;
assign v_35747 = v_35744 & v_35746;
assign v_35749 = v_35723 & v_35748;
assign v_35751 = v_33531;
assign v_35753 = v_35750 & v_35752;
assign v_35755 = v_35720 & v_35754;
assign v_35757 = v_33527;
assign v_35759 = v_35756 & v_35758;
assign v_35761 = v_35717 & v_35760;
assign v_35763 = v_33523;
assign v_35765 = v_35762 & v_35764;
assign v_35767 = v_35714 & v_35766;
assign v_35769 = v_33519;
assign v_35771 = v_35768 & v_35770;
assign v_35773 = v_35711 & v_35772;
assign v_35775 = v_33515;
assign v_35777 = v_35774 & v_35776;
assign v_35779 = v_35708 & v_35778;
assign v_35781 = v_33511;
assign v_35783 = v_35780 & v_35782;
assign v_35785 = v_35705 & v_35784;
assign v_35787 = v_33507;
assign v_35789 = v_35786 & v_35788;
assign v_35791 = v_35702 & v_35790;
assign v_35793 = v_33503;
assign v_35795 = v_35792 & v_35794;
assign v_35797 = v_35699 & v_35796;
assign v_35799 = v_33499;
assign v_35801 = v_35798 & v_35800;
assign v_35803 = v_35696 & v_35802;
assign v_35805 = v_33495;
assign v_35807 = v_35804 & v_35806;
assign v_35809 = v_35693 & v_35808;
assign v_35811 = v_2375;
assign v_35813 = v_35810 & v_35812;
assign v_35815 = v_35690 & v_35814;
assign v_35817 = v_2371;
assign v_35819 = v_35816 & v_35818;
assign v_35821 = v_35687 & v_35820;
assign v_35823 = v_2367;
assign v_35825 = v_35822 & v_35824;
assign v_35827 = v_35684 & v_35826;
assign v_35829 = v_2363;
assign v_35831 = v_35828 & v_35830;
assign v_35832 = v_35831;
assign v_35834 = v_33543;
assign v_35835 = v_2428;
assign v_35836 = v_35835;
assign v_35837 = v_35834 & v_35836;
assign v_35838 = v_35837;
assign v_35839 = v_35729 & v_35838;
assign v_35841 = v_35739 & v_35840;
assign v_35842 = v_35728 & v_35838;
assign v_35844 = v_35726 & v_35843;
assign v_35846 = v_35745 & v_35845;
assign v_35847 = v_35725 & v_35843;
assign v_35849 = v_35723 & v_35848;
assign v_35851 = v_35751 & v_35850;
assign v_35852 = v_35722 & v_35848;
assign v_35854 = v_35720 & v_35853;
assign v_35856 = v_35757 & v_35855;
assign v_35857 = v_35719 & v_35853;
assign v_35859 = v_35717 & v_35858;
assign v_35861 = v_35763 & v_35860;
assign v_35862 = v_35716 & v_35858;
assign v_35864 = v_35714 & v_35863;
assign v_35866 = v_35769 & v_35865;
assign v_35867 = v_35713 & v_35863;
assign v_35869 = v_35711 & v_35868;
assign v_35871 = v_35775 & v_35870;
assign v_35872 = v_35710 & v_35868;
assign v_35874 = v_35708 & v_35873;
assign v_35876 = v_35781 & v_35875;
assign v_35877 = v_35707 & v_35873;
assign v_35879 = v_35705 & v_35878;
assign v_35881 = v_35787 & v_35880;
assign v_35882 = v_35704 & v_35878;
assign v_35884 = v_35702 & v_35883;
assign v_35886 = v_35793 & v_35885;
assign v_35887 = v_35701 & v_35883;
assign v_35889 = v_35699 & v_35888;
assign v_35891 = v_35799 & v_35890;
assign v_35892 = v_35698 & v_35888;
assign v_35894 = v_35696 & v_35893;
assign v_35896 = v_35805 & v_35895;
assign v_35897 = v_35695 & v_35893;
assign v_35899 = v_35693 & v_35898;
assign v_35901 = v_35811 & v_35900;
assign v_35902 = v_35692 & v_35898;
assign v_35904 = v_35690 & v_35903;
assign v_35906 = v_35817 & v_35905;
assign v_35907 = v_35689 & v_35903;
assign v_35909 = v_35687 & v_35908;
assign v_35911 = v_35823 & v_35910;
assign v_35912 = v_35686 & v_35908;
assign v_35914 = v_35684 & v_35913;
assign v_35916 = v_35829 & v_35915;
assign v_35917 = v_35683 & v_35913;
assign v_35919 = v_35918;
assign v_35921 = v_35833 & v_35920;
assign v_35922 = v_35921;
assign v_35924 = v_35923;
assign v_35926 = ~v_2623;
assign v_35927 = ~v_33480;
assign v_35928 = v_33480;
assign v_35929 = ~v_2627;
assign v_35930 = ~v_33484;
assign v_35931 = v_33484;
assign v_35932 = ~v_2631;
assign v_35933 = ~v_33488;
assign v_35934 = v_33488;
assign v_35935 = ~v_2635;
assign v_35936 = ~v_33492;
assign v_35937 = v_33492;
assign v_35938 = ~v_33495;
assign v_35939 = ~v_2640;
assign v_35940 = v_2640;
assign v_35941 = ~v_33499;
assign v_35942 = ~v_2644;
assign v_35943 = v_2644;
assign v_35944 = ~v_33503;
assign v_35945 = ~v_2648;
assign v_35946 = v_2648;
assign v_35947 = ~v_33507;
assign v_35948 = ~v_2652;
assign v_35949 = v_2652;
assign v_35950 = ~v_33511;
assign v_35951 = ~v_2656;
assign v_35952 = v_2656;
assign v_35953 = ~v_33515;
assign v_35954 = ~v_2660;
assign v_35955 = v_2660;
assign v_35956 = ~v_33519;
assign v_35957 = ~v_2664;
assign v_35958 = v_2664;
assign v_35959 = ~v_33523;
assign v_35960 = ~v_2668;
assign v_35961 = v_2668;
assign v_35962 = ~v_33527;
assign v_35963 = ~v_2672;
assign v_35964 = v_2672;
assign v_35965 = ~v_33531;
assign v_35966 = ~v_2676;
assign v_35967 = v_2676;
assign v_35968 = ~v_33535;
assign v_35969 = ~v_2680;
assign v_35970 = v_2680;
assign v_35971 = ~v_33539;
assign v_35972 = ~v_2684;
assign v_35973 = v_2684;
assign v_35974 = ~v_33543;
assign v_35975 = ~v_2688;
assign v_35976 = v_35975;
assign v_35978 = v_35977;
assign v_35980 = v_35972 & v_35979;
assign v_35982 = v_33539;
assign v_35984 = v_35981 & v_35983;
assign v_35986 = v_35969 & v_35985;
assign v_35988 = v_33535;
assign v_35990 = v_35987 & v_35989;
assign v_35992 = v_35966 & v_35991;
assign v_35994 = v_33531;
assign v_35996 = v_35993 & v_35995;
assign v_35998 = v_35963 & v_35997;
assign v_36000 = v_33527;
assign v_36002 = v_35999 & v_36001;
assign v_36004 = v_35960 & v_36003;
assign v_36006 = v_33523;
assign v_36008 = v_36005 & v_36007;
assign v_36010 = v_35957 & v_36009;
assign v_36012 = v_33519;
assign v_36014 = v_36011 & v_36013;
assign v_36016 = v_35954 & v_36015;
assign v_36018 = v_33515;
assign v_36020 = v_36017 & v_36019;
assign v_36022 = v_35951 & v_36021;
assign v_36024 = v_33511;
assign v_36026 = v_36023 & v_36025;
assign v_36028 = v_35948 & v_36027;
assign v_36030 = v_33507;
assign v_36032 = v_36029 & v_36031;
assign v_36034 = v_35945 & v_36033;
assign v_36036 = v_33503;
assign v_36038 = v_36035 & v_36037;
assign v_36040 = v_35942 & v_36039;
assign v_36042 = v_33499;
assign v_36044 = v_36041 & v_36043;
assign v_36046 = v_35939 & v_36045;
assign v_36048 = v_33495;
assign v_36050 = v_36047 & v_36049;
assign v_36052 = v_35936 & v_36051;
assign v_36054 = v_2635;
assign v_36056 = v_36053 & v_36055;
assign v_36058 = v_35933 & v_36057;
assign v_36060 = v_2631;
assign v_36062 = v_36059 & v_36061;
assign v_36064 = v_35930 & v_36063;
assign v_36066 = v_2627;
assign v_36068 = v_36065 & v_36067;
assign v_36070 = v_35927 & v_36069;
assign v_36072 = v_2623;
assign v_36074 = v_36071 & v_36073;
assign v_36075 = v_36074;
assign v_36077 = v_33543;
assign v_36078 = v_2688;
assign v_36079 = v_36078;
assign v_36080 = v_36077 & v_36079;
assign v_36081 = v_36080;
assign v_36082 = v_35972 & v_36081;
assign v_36084 = v_35982 & v_36083;
assign v_36085 = v_35971 & v_36081;
assign v_36087 = v_35969 & v_36086;
assign v_36089 = v_35988 & v_36088;
assign v_36090 = v_35968 & v_36086;
assign v_36092 = v_35966 & v_36091;
assign v_36094 = v_35994 & v_36093;
assign v_36095 = v_35965 & v_36091;
assign v_36097 = v_35963 & v_36096;
assign v_36099 = v_36000 & v_36098;
assign v_36100 = v_35962 & v_36096;
assign v_36102 = v_35960 & v_36101;
assign v_36104 = v_36006 & v_36103;
assign v_36105 = v_35959 & v_36101;
assign v_36107 = v_35957 & v_36106;
assign v_36109 = v_36012 & v_36108;
assign v_36110 = v_35956 & v_36106;
assign v_36112 = v_35954 & v_36111;
assign v_36114 = v_36018 & v_36113;
assign v_36115 = v_35953 & v_36111;
assign v_36117 = v_35951 & v_36116;
assign v_36119 = v_36024 & v_36118;
assign v_36120 = v_35950 & v_36116;
assign v_36122 = v_35948 & v_36121;
assign v_36124 = v_36030 & v_36123;
assign v_36125 = v_35947 & v_36121;
assign v_36127 = v_35945 & v_36126;
assign v_36129 = v_36036 & v_36128;
assign v_36130 = v_35944 & v_36126;
assign v_36132 = v_35942 & v_36131;
assign v_36134 = v_36042 & v_36133;
assign v_36135 = v_35941 & v_36131;
assign v_36137 = v_35939 & v_36136;
assign v_36139 = v_36048 & v_36138;
assign v_36140 = v_35938 & v_36136;
assign v_36142 = v_35936 & v_36141;
assign v_36144 = v_36054 & v_36143;
assign v_36145 = v_35935 & v_36141;
assign v_36147 = v_35933 & v_36146;
assign v_36149 = v_36060 & v_36148;
assign v_36150 = v_35932 & v_36146;
assign v_36152 = v_35930 & v_36151;
assign v_36154 = v_36066 & v_36153;
assign v_36155 = v_35929 & v_36151;
assign v_36157 = v_35927 & v_36156;
assign v_36159 = v_36072 & v_36158;
assign v_36160 = v_35926 & v_36156;
assign v_36162 = v_36161;
assign v_36164 = v_36076 & v_36163;
assign v_36165 = v_36164;
assign v_36167 = v_36166;
assign v_36169 = ~v_2883;
assign v_36170 = ~v_33480;
assign v_36171 = v_33480;
assign v_36172 = ~v_2887;
assign v_36173 = ~v_33484;
assign v_36174 = v_33484;
assign v_36175 = ~v_2891;
assign v_36176 = ~v_33488;
assign v_36177 = v_33488;
assign v_36178 = ~v_2895;
assign v_36179 = ~v_33492;
assign v_36180 = v_33492;
assign v_36181 = ~v_33495;
assign v_36182 = ~v_2900;
assign v_36183 = v_2900;
assign v_36184 = ~v_33499;
assign v_36185 = ~v_2904;
assign v_36186 = v_2904;
assign v_36187 = ~v_33503;
assign v_36188 = ~v_2908;
assign v_36189 = v_2908;
assign v_36190 = ~v_33507;
assign v_36191 = ~v_2912;
assign v_36192 = v_2912;
assign v_36193 = ~v_33511;
assign v_36194 = ~v_2916;
assign v_36195 = v_2916;
assign v_36196 = ~v_33515;
assign v_36197 = ~v_2920;
assign v_36198 = v_2920;
assign v_36199 = ~v_33519;
assign v_36200 = ~v_2924;
assign v_36201 = v_2924;
assign v_36202 = ~v_33523;
assign v_36203 = ~v_2928;
assign v_36204 = v_2928;
assign v_36205 = ~v_33527;
assign v_36206 = ~v_2932;
assign v_36207 = v_2932;
assign v_36208 = ~v_33531;
assign v_36209 = ~v_2936;
assign v_36210 = v_2936;
assign v_36211 = ~v_33535;
assign v_36212 = ~v_2940;
assign v_36213 = v_2940;
assign v_36214 = ~v_33539;
assign v_36215 = ~v_2944;
assign v_36216 = v_2944;
assign v_36217 = ~v_33543;
assign v_36218 = ~v_2948;
assign v_36219 = v_36218;
assign v_36221 = v_36220;
assign v_36223 = v_36215 & v_36222;
assign v_36225 = v_33539;
assign v_36227 = v_36224 & v_36226;
assign v_36229 = v_36212 & v_36228;
assign v_36231 = v_33535;
assign v_36233 = v_36230 & v_36232;
assign v_36235 = v_36209 & v_36234;
assign v_36237 = v_33531;
assign v_36239 = v_36236 & v_36238;
assign v_36241 = v_36206 & v_36240;
assign v_36243 = v_33527;
assign v_36245 = v_36242 & v_36244;
assign v_36247 = v_36203 & v_36246;
assign v_36249 = v_33523;
assign v_36251 = v_36248 & v_36250;
assign v_36253 = v_36200 & v_36252;
assign v_36255 = v_33519;
assign v_36257 = v_36254 & v_36256;
assign v_36259 = v_36197 & v_36258;
assign v_36261 = v_33515;
assign v_36263 = v_36260 & v_36262;
assign v_36265 = v_36194 & v_36264;
assign v_36267 = v_33511;
assign v_36269 = v_36266 & v_36268;
assign v_36271 = v_36191 & v_36270;
assign v_36273 = v_33507;
assign v_36275 = v_36272 & v_36274;
assign v_36277 = v_36188 & v_36276;
assign v_36279 = v_33503;
assign v_36281 = v_36278 & v_36280;
assign v_36283 = v_36185 & v_36282;
assign v_36285 = v_33499;
assign v_36287 = v_36284 & v_36286;
assign v_36289 = v_36182 & v_36288;
assign v_36291 = v_33495;
assign v_36293 = v_36290 & v_36292;
assign v_36295 = v_36179 & v_36294;
assign v_36297 = v_2895;
assign v_36299 = v_36296 & v_36298;
assign v_36301 = v_36176 & v_36300;
assign v_36303 = v_2891;
assign v_36305 = v_36302 & v_36304;
assign v_36307 = v_36173 & v_36306;
assign v_36309 = v_2887;
assign v_36311 = v_36308 & v_36310;
assign v_36313 = v_36170 & v_36312;
assign v_36315 = v_2883;
assign v_36317 = v_36314 & v_36316;
assign v_36318 = v_36317;
assign v_36320 = v_33543;
assign v_36321 = v_2948;
assign v_36322 = v_36321;
assign v_36323 = v_36320 & v_36322;
assign v_36324 = v_36323;
assign v_36325 = v_36215 & v_36324;
assign v_36327 = v_36225 & v_36326;
assign v_36328 = v_36214 & v_36324;
assign v_36330 = v_36212 & v_36329;
assign v_36332 = v_36231 & v_36331;
assign v_36333 = v_36211 & v_36329;
assign v_36335 = v_36209 & v_36334;
assign v_36337 = v_36237 & v_36336;
assign v_36338 = v_36208 & v_36334;
assign v_36340 = v_36206 & v_36339;
assign v_36342 = v_36243 & v_36341;
assign v_36343 = v_36205 & v_36339;
assign v_36345 = v_36203 & v_36344;
assign v_36347 = v_36249 & v_36346;
assign v_36348 = v_36202 & v_36344;
assign v_36350 = v_36200 & v_36349;
assign v_36352 = v_36255 & v_36351;
assign v_36353 = v_36199 & v_36349;
assign v_36355 = v_36197 & v_36354;
assign v_36357 = v_36261 & v_36356;
assign v_36358 = v_36196 & v_36354;
assign v_36360 = v_36194 & v_36359;
assign v_36362 = v_36267 & v_36361;
assign v_36363 = v_36193 & v_36359;
assign v_36365 = v_36191 & v_36364;
assign v_36367 = v_36273 & v_36366;
assign v_36368 = v_36190 & v_36364;
assign v_36370 = v_36188 & v_36369;
assign v_36372 = v_36279 & v_36371;
assign v_36373 = v_36187 & v_36369;
assign v_36375 = v_36185 & v_36374;
assign v_36377 = v_36285 & v_36376;
assign v_36378 = v_36184 & v_36374;
assign v_36380 = v_36182 & v_36379;
assign v_36382 = v_36291 & v_36381;
assign v_36383 = v_36181 & v_36379;
assign v_36385 = v_36179 & v_36384;
assign v_36387 = v_36297 & v_36386;
assign v_36388 = v_36178 & v_36384;
assign v_36390 = v_36176 & v_36389;
assign v_36392 = v_36303 & v_36391;
assign v_36393 = v_36175 & v_36389;
assign v_36395 = v_36173 & v_36394;
assign v_36397 = v_36309 & v_36396;
assign v_36398 = v_36172 & v_36394;
assign v_36400 = v_36170 & v_36399;
assign v_36402 = v_36315 & v_36401;
assign v_36403 = v_36169 & v_36399;
assign v_36405 = v_36404;
assign v_36407 = v_36319 & v_36406;
assign v_36408 = v_36407;
assign v_36410 = v_36409;
assign v_36412 = ~v_3143;
assign v_36413 = ~v_33480;
assign v_36414 = v_33480;
assign v_36415 = ~v_3147;
assign v_36416 = ~v_33484;
assign v_36417 = v_33484;
assign v_36418 = ~v_3151;
assign v_36419 = ~v_33488;
assign v_36420 = v_33488;
assign v_36421 = ~v_3155;
assign v_36422 = ~v_33492;
assign v_36423 = v_33492;
assign v_36424 = ~v_33495;
assign v_36425 = ~v_3160;
assign v_36426 = v_3160;
assign v_36427 = ~v_33499;
assign v_36428 = ~v_3164;
assign v_36429 = v_3164;
assign v_36430 = ~v_33503;
assign v_36431 = ~v_3168;
assign v_36432 = v_3168;
assign v_36433 = ~v_33507;
assign v_36434 = ~v_3172;
assign v_36435 = v_3172;
assign v_36436 = ~v_33511;
assign v_36437 = ~v_3176;
assign v_36438 = v_3176;
assign v_36439 = ~v_33515;
assign v_36440 = ~v_3180;
assign v_36441 = v_3180;
assign v_36442 = ~v_33519;
assign v_36443 = ~v_3184;
assign v_36444 = v_3184;
assign v_36445 = ~v_33523;
assign v_36446 = ~v_3188;
assign v_36447 = v_3188;
assign v_36448 = ~v_33527;
assign v_36449 = ~v_3192;
assign v_36450 = v_3192;
assign v_36451 = ~v_33531;
assign v_36452 = ~v_3196;
assign v_36453 = v_3196;
assign v_36454 = ~v_33535;
assign v_36455 = ~v_3200;
assign v_36456 = v_3200;
assign v_36457 = ~v_33539;
assign v_36458 = ~v_3204;
assign v_36459 = v_3204;
assign v_36460 = ~v_33543;
assign v_36461 = ~v_3208;
assign v_36462 = v_36461;
assign v_36464 = v_36463;
assign v_36466 = v_36458 & v_36465;
assign v_36468 = v_33539;
assign v_36470 = v_36467 & v_36469;
assign v_36472 = v_36455 & v_36471;
assign v_36474 = v_33535;
assign v_36476 = v_36473 & v_36475;
assign v_36478 = v_36452 & v_36477;
assign v_36480 = v_33531;
assign v_36482 = v_36479 & v_36481;
assign v_36484 = v_36449 & v_36483;
assign v_36486 = v_33527;
assign v_36488 = v_36485 & v_36487;
assign v_36490 = v_36446 & v_36489;
assign v_36492 = v_33523;
assign v_36494 = v_36491 & v_36493;
assign v_36496 = v_36443 & v_36495;
assign v_36498 = v_33519;
assign v_36500 = v_36497 & v_36499;
assign v_36502 = v_36440 & v_36501;
assign v_36504 = v_33515;
assign v_36506 = v_36503 & v_36505;
assign v_36508 = v_36437 & v_36507;
assign v_36510 = v_33511;
assign v_36512 = v_36509 & v_36511;
assign v_36514 = v_36434 & v_36513;
assign v_36516 = v_33507;
assign v_36518 = v_36515 & v_36517;
assign v_36520 = v_36431 & v_36519;
assign v_36522 = v_33503;
assign v_36524 = v_36521 & v_36523;
assign v_36526 = v_36428 & v_36525;
assign v_36528 = v_33499;
assign v_36530 = v_36527 & v_36529;
assign v_36532 = v_36425 & v_36531;
assign v_36534 = v_33495;
assign v_36536 = v_36533 & v_36535;
assign v_36538 = v_36422 & v_36537;
assign v_36540 = v_3155;
assign v_36542 = v_36539 & v_36541;
assign v_36544 = v_36419 & v_36543;
assign v_36546 = v_3151;
assign v_36548 = v_36545 & v_36547;
assign v_36550 = v_36416 & v_36549;
assign v_36552 = v_3147;
assign v_36554 = v_36551 & v_36553;
assign v_36556 = v_36413 & v_36555;
assign v_36558 = v_3143;
assign v_36560 = v_36557 & v_36559;
assign v_36561 = v_36560;
assign v_36563 = v_33543;
assign v_36564 = v_3208;
assign v_36565 = v_36564;
assign v_36566 = v_36563 & v_36565;
assign v_36567 = v_36566;
assign v_36568 = v_36458 & v_36567;
assign v_36570 = v_36468 & v_36569;
assign v_36571 = v_36457 & v_36567;
assign v_36573 = v_36455 & v_36572;
assign v_36575 = v_36474 & v_36574;
assign v_36576 = v_36454 & v_36572;
assign v_36578 = v_36452 & v_36577;
assign v_36580 = v_36480 & v_36579;
assign v_36581 = v_36451 & v_36577;
assign v_36583 = v_36449 & v_36582;
assign v_36585 = v_36486 & v_36584;
assign v_36586 = v_36448 & v_36582;
assign v_36588 = v_36446 & v_36587;
assign v_36590 = v_36492 & v_36589;
assign v_36591 = v_36445 & v_36587;
assign v_36593 = v_36443 & v_36592;
assign v_36595 = v_36498 & v_36594;
assign v_36596 = v_36442 & v_36592;
assign v_36598 = v_36440 & v_36597;
assign v_36600 = v_36504 & v_36599;
assign v_36601 = v_36439 & v_36597;
assign v_36603 = v_36437 & v_36602;
assign v_36605 = v_36510 & v_36604;
assign v_36606 = v_36436 & v_36602;
assign v_36608 = v_36434 & v_36607;
assign v_36610 = v_36516 & v_36609;
assign v_36611 = v_36433 & v_36607;
assign v_36613 = v_36431 & v_36612;
assign v_36615 = v_36522 & v_36614;
assign v_36616 = v_36430 & v_36612;
assign v_36618 = v_36428 & v_36617;
assign v_36620 = v_36528 & v_36619;
assign v_36621 = v_36427 & v_36617;
assign v_36623 = v_36425 & v_36622;
assign v_36625 = v_36534 & v_36624;
assign v_36626 = v_36424 & v_36622;
assign v_36628 = v_36422 & v_36627;
assign v_36630 = v_36540 & v_36629;
assign v_36631 = v_36421 & v_36627;
assign v_36633 = v_36419 & v_36632;
assign v_36635 = v_36546 & v_36634;
assign v_36636 = v_36418 & v_36632;
assign v_36638 = v_36416 & v_36637;
assign v_36640 = v_36552 & v_36639;
assign v_36641 = v_36415 & v_36637;
assign v_36643 = v_36413 & v_36642;
assign v_36645 = v_36558 & v_36644;
assign v_36646 = v_36412 & v_36642;
assign v_36648 = v_36647;
assign v_36650 = v_36562 & v_36649;
assign v_36651 = v_36650;
assign v_36653 = v_36652;
assign v_36655 = ~v_3403;
assign v_36656 = ~v_33480;
assign v_36657 = v_33480;
assign v_36658 = ~v_3407;
assign v_36659 = ~v_33484;
assign v_36660 = v_33484;
assign v_36661 = ~v_3411;
assign v_36662 = ~v_33488;
assign v_36663 = v_33488;
assign v_36664 = ~v_3415;
assign v_36665 = ~v_33492;
assign v_36666 = v_33492;
assign v_36667 = ~v_33495;
assign v_36668 = ~v_3420;
assign v_36669 = v_3420;
assign v_36670 = ~v_33499;
assign v_36671 = ~v_3424;
assign v_36672 = v_3424;
assign v_36673 = ~v_33503;
assign v_36674 = ~v_3428;
assign v_36675 = v_3428;
assign v_36676 = ~v_33507;
assign v_36677 = ~v_3432;
assign v_36678 = v_3432;
assign v_36679 = ~v_33511;
assign v_36680 = ~v_3436;
assign v_36681 = v_3436;
assign v_36682 = ~v_33515;
assign v_36683 = ~v_3440;
assign v_36684 = v_3440;
assign v_36685 = ~v_33519;
assign v_36686 = ~v_3444;
assign v_36687 = v_3444;
assign v_36688 = ~v_33523;
assign v_36689 = ~v_3448;
assign v_36690 = v_3448;
assign v_36691 = ~v_33527;
assign v_36692 = ~v_3452;
assign v_36693 = v_3452;
assign v_36694 = ~v_33531;
assign v_36695 = ~v_3456;
assign v_36696 = v_3456;
assign v_36697 = ~v_33535;
assign v_36698 = ~v_3460;
assign v_36699 = v_3460;
assign v_36700 = ~v_33539;
assign v_36701 = ~v_3464;
assign v_36702 = v_3464;
assign v_36703 = ~v_33543;
assign v_36704 = ~v_3468;
assign v_36705 = v_36704;
assign v_36707 = v_36706;
assign v_36709 = v_36701 & v_36708;
assign v_36711 = v_33539;
assign v_36713 = v_36710 & v_36712;
assign v_36715 = v_36698 & v_36714;
assign v_36717 = v_33535;
assign v_36719 = v_36716 & v_36718;
assign v_36721 = v_36695 & v_36720;
assign v_36723 = v_33531;
assign v_36725 = v_36722 & v_36724;
assign v_36727 = v_36692 & v_36726;
assign v_36729 = v_33527;
assign v_36731 = v_36728 & v_36730;
assign v_36733 = v_36689 & v_36732;
assign v_36735 = v_33523;
assign v_36737 = v_36734 & v_36736;
assign v_36739 = v_36686 & v_36738;
assign v_36741 = v_33519;
assign v_36743 = v_36740 & v_36742;
assign v_36745 = v_36683 & v_36744;
assign v_36747 = v_33515;
assign v_36749 = v_36746 & v_36748;
assign v_36751 = v_36680 & v_36750;
assign v_36753 = v_33511;
assign v_36755 = v_36752 & v_36754;
assign v_36757 = v_36677 & v_36756;
assign v_36759 = v_33507;
assign v_36761 = v_36758 & v_36760;
assign v_36763 = v_36674 & v_36762;
assign v_36765 = v_33503;
assign v_36767 = v_36764 & v_36766;
assign v_36769 = v_36671 & v_36768;
assign v_36771 = v_33499;
assign v_36773 = v_36770 & v_36772;
assign v_36775 = v_36668 & v_36774;
assign v_36777 = v_33495;
assign v_36779 = v_36776 & v_36778;
assign v_36781 = v_36665 & v_36780;
assign v_36783 = v_3415;
assign v_36785 = v_36782 & v_36784;
assign v_36787 = v_36662 & v_36786;
assign v_36789 = v_3411;
assign v_36791 = v_36788 & v_36790;
assign v_36793 = v_36659 & v_36792;
assign v_36795 = v_3407;
assign v_36797 = v_36794 & v_36796;
assign v_36799 = v_36656 & v_36798;
assign v_36801 = v_3403;
assign v_36803 = v_36800 & v_36802;
assign v_36804 = v_36803;
assign v_36806 = v_33543;
assign v_36807 = v_3468;
assign v_36808 = v_36807;
assign v_36809 = v_36806 & v_36808;
assign v_36810 = v_36809;
assign v_36811 = v_36701 & v_36810;
assign v_36813 = v_36711 & v_36812;
assign v_36814 = v_36700 & v_36810;
assign v_36816 = v_36698 & v_36815;
assign v_36818 = v_36717 & v_36817;
assign v_36819 = v_36697 & v_36815;
assign v_36821 = v_36695 & v_36820;
assign v_36823 = v_36723 & v_36822;
assign v_36824 = v_36694 & v_36820;
assign v_36826 = v_36692 & v_36825;
assign v_36828 = v_36729 & v_36827;
assign v_36829 = v_36691 & v_36825;
assign v_36831 = v_36689 & v_36830;
assign v_36833 = v_36735 & v_36832;
assign v_36834 = v_36688 & v_36830;
assign v_36836 = v_36686 & v_36835;
assign v_36838 = v_36741 & v_36837;
assign v_36839 = v_36685 & v_36835;
assign v_36841 = v_36683 & v_36840;
assign v_36843 = v_36747 & v_36842;
assign v_36844 = v_36682 & v_36840;
assign v_36846 = v_36680 & v_36845;
assign v_36848 = v_36753 & v_36847;
assign v_36849 = v_36679 & v_36845;
assign v_36851 = v_36677 & v_36850;
assign v_36853 = v_36759 & v_36852;
assign v_36854 = v_36676 & v_36850;
assign v_36856 = v_36674 & v_36855;
assign v_36858 = v_36765 & v_36857;
assign v_36859 = v_36673 & v_36855;
assign v_36861 = v_36671 & v_36860;
assign v_36863 = v_36771 & v_36862;
assign v_36864 = v_36670 & v_36860;
assign v_36866 = v_36668 & v_36865;
assign v_36868 = v_36777 & v_36867;
assign v_36869 = v_36667 & v_36865;
assign v_36871 = v_36665 & v_36870;
assign v_36873 = v_36783 & v_36872;
assign v_36874 = v_36664 & v_36870;
assign v_36876 = v_36662 & v_36875;
assign v_36878 = v_36789 & v_36877;
assign v_36879 = v_36661 & v_36875;
assign v_36881 = v_36659 & v_36880;
assign v_36883 = v_36795 & v_36882;
assign v_36884 = v_36658 & v_36880;
assign v_36886 = v_36656 & v_36885;
assign v_36888 = v_36801 & v_36887;
assign v_36889 = v_36655 & v_36885;
assign v_36891 = v_36890;
assign v_36893 = v_36805 & v_36892;
assign v_36894 = v_36893;
assign v_36896 = v_36895;
assign v_36898 = ~v_3663;
assign v_36899 = ~v_33480;
assign v_36900 = v_33480;
assign v_36901 = ~v_3667;
assign v_36902 = ~v_33484;
assign v_36903 = v_33484;
assign v_36904 = ~v_3671;
assign v_36905 = ~v_33488;
assign v_36906 = v_33488;
assign v_36907 = ~v_3675;
assign v_36908 = ~v_33492;
assign v_36909 = v_33492;
assign v_36910 = ~v_33495;
assign v_36911 = ~v_3680;
assign v_36912 = v_3680;
assign v_36913 = ~v_33499;
assign v_36914 = ~v_3684;
assign v_36915 = v_3684;
assign v_36916 = ~v_33503;
assign v_36917 = ~v_3688;
assign v_36918 = v_3688;
assign v_36919 = ~v_33507;
assign v_36920 = ~v_3692;
assign v_36921 = v_3692;
assign v_36922 = ~v_33511;
assign v_36923 = ~v_3696;
assign v_36924 = v_3696;
assign v_36925 = ~v_33515;
assign v_36926 = ~v_3700;
assign v_36927 = v_3700;
assign v_36928 = ~v_33519;
assign v_36929 = ~v_3704;
assign v_36930 = v_3704;
assign v_36931 = ~v_33523;
assign v_36932 = ~v_3708;
assign v_36933 = v_3708;
assign v_36934 = ~v_33527;
assign v_36935 = ~v_3712;
assign v_36936 = v_3712;
assign v_36937 = ~v_33531;
assign v_36938 = ~v_3716;
assign v_36939 = v_3716;
assign v_36940 = ~v_33535;
assign v_36941 = ~v_3720;
assign v_36942 = v_3720;
assign v_36943 = ~v_33539;
assign v_36944 = ~v_3724;
assign v_36945 = v_3724;
assign v_36946 = ~v_33543;
assign v_36947 = ~v_3728;
assign v_36948 = v_36947;
assign v_36950 = v_36949;
assign v_36952 = v_36944 & v_36951;
assign v_36954 = v_33539;
assign v_36956 = v_36953 & v_36955;
assign v_36958 = v_36941 & v_36957;
assign v_36960 = v_33535;
assign v_36962 = v_36959 & v_36961;
assign v_36964 = v_36938 & v_36963;
assign v_36966 = v_33531;
assign v_36968 = v_36965 & v_36967;
assign v_36970 = v_36935 & v_36969;
assign v_36972 = v_33527;
assign v_36974 = v_36971 & v_36973;
assign v_36976 = v_36932 & v_36975;
assign v_36978 = v_33523;
assign v_36980 = v_36977 & v_36979;
assign v_36982 = v_36929 & v_36981;
assign v_36984 = v_33519;
assign v_36986 = v_36983 & v_36985;
assign v_36988 = v_36926 & v_36987;
assign v_36990 = v_33515;
assign v_36992 = v_36989 & v_36991;
assign v_36994 = v_36923 & v_36993;
assign v_36996 = v_33511;
assign v_36998 = v_36995 & v_36997;
assign v_37000 = v_36920 & v_36999;
assign v_37002 = v_33507;
assign v_37004 = v_37001 & v_37003;
assign v_37006 = v_36917 & v_37005;
assign v_37008 = v_33503;
assign v_37010 = v_37007 & v_37009;
assign v_37012 = v_36914 & v_37011;
assign v_37014 = v_33499;
assign v_37016 = v_37013 & v_37015;
assign v_37018 = v_36911 & v_37017;
assign v_37020 = v_33495;
assign v_37022 = v_37019 & v_37021;
assign v_37024 = v_36908 & v_37023;
assign v_37026 = v_3675;
assign v_37028 = v_37025 & v_37027;
assign v_37030 = v_36905 & v_37029;
assign v_37032 = v_3671;
assign v_37034 = v_37031 & v_37033;
assign v_37036 = v_36902 & v_37035;
assign v_37038 = v_3667;
assign v_37040 = v_37037 & v_37039;
assign v_37042 = v_36899 & v_37041;
assign v_37044 = v_3663;
assign v_37046 = v_37043 & v_37045;
assign v_37047 = v_37046;
assign v_37049 = v_33543;
assign v_37050 = v_3728;
assign v_37051 = v_37050;
assign v_37052 = v_37049 & v_37051;
assign v_37053 = v_37052;
assign v_37054 = v_36944 & v_37053;
assign v_37056 = v_36954 & v_37055;
assign v_37057 = v_36943 & v_37053;
assign v_37059 = v_36941 & v_37058;
assign v_37061 = v_36960 & v_37060;
assign v_37062 = v_36940 & v_37058;
assign v_37064 = v_36938 & v_37063;
assign v_37066 = v_36966 & v_37065;
assign v_37067 = v_36937 & v_37063;
assign v_37069 = v_36935 & v_37068;
assign v_37071 = v_36972 & v_37070;
assign v_37072 = v_36934 & v_37068;
assign v_37074 = v_36932 & v_37073;
assign v_37076 = v_36978 & v_37075;
assign v_37077 = v_36931 & v_37073;
assign v_37079 = v_36929 & v_37078;
assign v_37081 = v_36984 & v_37080;
assign v_37082 = v_36928 & v_37078;
assign v_37084 = v_36926 & v_37083;
assign v_37086 = v_36990 & v_37085;
assign v_37087 = v_36925 & v_37083;
assign v_37089 = v_36923 & v_37088;
assign v_37091 = v_36996 & v_37090;
assign v_37092 = v_36922 & v_37088;
assign v_37094 = v_36920 & v_37093;
assign v_37096 = v_37002 & v_37095;
assign v_37097 = v_36919 & v_37093;
assign v_37099 = v_36917 & v_37098;
assign v_37101 = v_37008 & v_37100;
assign v_37102 = v_36916 & v_37098;
assign v_37104 = v_36914 & v_37103;
assign v_37106 = v_37014 & v_37105;
assign v_37107 = v_36913 & v_37103;
assign v_37109 = v_36911 & v_37108;
assign v_37111 = v_37020 & v_37110;
assign v_37112 = v_36910 & v_37108;
assign v_37114 = v_36908 & v_37113;
assign v_37116 = v_37026 & v_37115;
assign v_37117 = v_36907 & v_37113;
assign v_37119 = v_36905 & v_37118;
assign v_37121 = v_37032 & v_37120;
assign v_37122 = v_36904 & v_37118;
assign v_37124 = v_36902 & v_37123;
assign v_37126 = v_37038 & v_37125;
assign v_37127 = v_36901 & v_37123;
assign v_37129 = v_36899 & v_37128;
assign v_37131 = v_37044 & v_37130;
assign v_37132 = v_36898 & v_37128;
assign v_37134 = v_37133;
assign v_37136 = v_37048 & v_37135;
assign v_37137 = v_37136;
assign v_37139 = v_37138;
assign v_37141 = ~v_3923;
assign v_37142 = ~v_33480;
assign v_37143 = v_33480;
assign v_37144 = ~v_3927;
assign v_37145 = ~v_33484;
assign v_37146 = v_33484;
assign v_37147 = ~v_3931;
assign v_37148 = ~v_33488;
assign v_37149 = v_33488;
assign v_37150 = ~v_3935;
assign v_37151 = ~v_33492;
assign v_37152 = v_33492;
assign v_37153 = ~v_33495;
assign v_37154 = ~v_3940;
assign v_37155 = v_3940;
assign v_37156 = ~v_33499;
assign v_37157 = ~v_3944;
assign v_37158 = v_3944;
assign v_37159 = ~v_33503;
assign v_37160 = ~v_3948;
assign v_37161 = v_3948;
assign v_37162 = ~v_33507;
assign v_37163 = ~v_3952;
assign v_37164 = v_3952;
assign v_37165 = ~v_33511;
assign v_37166 = ~v_3956;
assign v_37167 = v_3956;
assign v_37168 = ~v_33515;
assign v_37169 = ~v_3960;
assign v_37170 = v_3960;
assign v_37171 = ~v_33519;
assign v_37172 = ~v_3964;
assign v_37173 = v_3964;
assign v_37174 = ~v_33523;
assign v_37175 = ~v_3968;
assign v_37176 = v_3968;
assign v_37177 = ~v_33527;
assign v_37178 = ~v_3972;
assign v_37179 = v_3972;
assign v_37180 = ~v_33531;
assign v_37181 = ~v_3976;
assign v_37182 = v_3976;
assign v_37183 = ~v_33535;
assign v_37184 = ~v_3980;
assign v_37185 = v_3980;
assign v_37186 = ~v_33539;
assign v_37187 = ~v_3984;
assign v_37188 = v_3984;
assign v_37189 = ~v_33543;
assign v_37190 = ~v_3988;
assign v_37191 = v_37190;
assign v_37193 = v_37192;
assign v_37195 = v_37187 & v_37194;
assign v_37197 = v_33539;
assign v_37199 = v_37196 & v_37198;
assign v_37201 = v_37184 & v_37200;
assign v_37203 = v_33535;
assign v_37205 = v_37202 & v_37204;
assign v_37207 = v_37181 & v_37206;
assign v_37209 = v_33531;
assign v_37211 = v_37208 & v_37210;
assign v_37213 = v_37178 & v_37212;
assign v_37215 = v_33527;
assign v_37217 = v_37214 & v_37216;
assign v_37219 = v_37175 & v_37218;
assign v_37221 = v_33523;
assign v_37223 = v_37220 & v_37222;
assign v_37225 = v_37172 & v_37224;
assign v_37227 = v_33519;
assign v_37229 = v_37226 & v_37228;
assign v_37231 = v_37169 & v_37230;
assign v_37233 = v_33515;
assign v_37235 = v_37232 & v_37234;
assign v_37237 = v_37166 & v_37236;
assign v_37239 = v_33511;
assign v_37241 = v_37238 & v_37240;
assign v_37243 = v_37163 & v_37242;
assign v_37245 = v_33507;
assign v_37247 = v_37244 & v_37246;
assign v_37249 = v_37160 & v_37248;
assign v_37251 = v_33503;
assign v_37253 = v_37250 & v_37252;
assign v_37255 = v_37157 & v_37254;
assign v_37257 = v_33499;
assign v_37259 = v_37256 & v_37258;
assign v_37261 = v_37154 & v_37260;
assign v_37263 = v_33495;
assign v_37265 = v_37262 & v_37264;
assign v_37267 = v_37151 & v_37266;
assign v_37269 = v_3935;
assign v_37271 = v_37268 & v_37270;
assign v_37273 = v_37148 & v_37272;
assign v_37275 = v_3931;
assign v_37277 = v_37274 & v_37276;
assign v_37279 = v_37145 & v_37278;
assign v_37281 = v_3927;
assign v_37283 = v_37280 & v_37282;
assign v_37285 = v_37142 & v_37284;
assign v_37287 = v_3923;
assign v_37289 = v_37286 & v_37288;
assign v_37290 = v_37289;
assign v_37292 = v_33543;
assign v_37293 = v_3988;
assign v_37294 = v_37293;
assign v_37295 = v_37292 & v_37294;
assign v_37296 = v_37295;
assign v_37297 = v_37187 & v_37296;
assign v_37299 = v_37197 & v_37298;
assign v_37300 = v_37186 & v_37296;
assign v_37302 = v_37184 & v_37301;
assign v_37304 = v_37203 & v_37303;
assign v_37305 = v_37183 & v_37301;
assign v_37307 = v_37181 & v_37306;
assign v_37309 = v_37209 & v_37308;
assign v_37310 = v_37180 & v_37306;
assign v_37312 = v_37178 & v_37311;
assign v_37314 = v_37215 & v_37313;
assign v_37315 = v_37177 & v_37311;
assign v_37317 = v_37175 & v_37316;
assign v_37319 = v_37221 & v_37318;
assign v_37320 = v_37174 & v_37316;
assign v_37322 = v_37172 & v_37321;
assign v_37324 = v_37227 & v_37323;
assign v_37325 = v_37171 & v_37321;
assign v_37327 = v_37169 & v_37326;
assign v_37329 = v_37233 & v_37328;
assign v_37330 = v_37168 & v_37326;
assign v_37332 = v_37166 & v_37331;
assign v_37334 = v_37239 & v_37333;
assign v_37335 = v_37165 & v_37331;
assign v_37337 = v_37163 & v_37336;
assign v_37339 = v_37245 & v_37338;
assign v_37340 = v_37162 & v_37336;
assign v_37342 = v_37160 & v_37341;
assign v_37344 = v_37251 & v_37343;
assign v_37345 = v_37159 & v_37341;
assign v_37347 = v_37157 & v_37346;
assign v_37349 = v_37257 & v_37348;
assign v_37350 = v_37156 & v_37346;
assign v_37352 = v_37154 & v_37351;
assign v_37354 = v_37263 & v_37353;
assign v_37355 = v_37153 & v_37351;
assign v_37357 = v_37151 & v_37356;
assign v_37359 = v_37269 & v_37358;
assign v_37360 = v_37150 & v_37356;
assign v_37362 = v_37148 & v_37361;
assign v_37364 = v_37275 & v_37363;
assign v_37365 = v_37147 & v_37361;
assign v_37367 = v_37145 & v_37366;
assign v_37369 = v_37281 & v_37368;
assign v_37370 = v_37144 & v_37366;
assign v_37372 = v_37142 & v_37371;
assign v_37374 = v_37287 & v_37373;
assign v_37375 = v_37141 & v_37371;
assign v_37377 = v_37376;
assign v_37379 = v_37291 & v_37378;
assign v_37380 = v_37379;
assign v_37382 = v_37381;
assign v_37383 = ~v_4182;
assign v_37384 = ~v_33480;
assign v_37385 = v_33480;
assign v_37386 = ~v_4186;
assign v_37387 = ~v_33484;
assign v_37388 = v_33484;
assign v_37389 = ~v_4190;
assign v_37390 = ~v_33488;
assign v_37391 = v_33488;
assign v_37392 = ~v_4194;
assign v_37393 = ~v_33492;
assign v_37394 = v_33492;
assign v_37395 = ~v_33495;
assign v_37396 = ~v_4199;
assign v_37397 = v_4199;
assign v_37398 = ~v_33499;
assign v_37399 = ~v_4203;
assign v_37400 = v_4203;
assign v_37401 = ~v_33503;
assign v_37402 = ~v_4207;
assign v_37403 = v_4207;
assign v_37404 = ~v_33507;
assign v_37405 = ~v_4211;
assign v_37406 = v_4211;
assign v_37407 = ~v_33511;
assign v_37408 = ~v_4215;
assign v_37409 = v_4215;
assign v_37410 = ~v_33515;
assign v_37411 = ~v_4219;
assign v_37412 = v_4219;
assign v_37413 = ~v_33519;
assign v_37414 = ~v_4223;
assign v_37415 = v_4223;
assign v_37416 = ~v_33523;
assign v_37417 = ~v_4227;
assign v_37418 = v_4227;
assign v_37419 = ~v_33527;
assign v_37420 = ~v_4231;
assign v_37421 = v_4231;
assign v_37422 = ~v_33531;
assign v_37423 = ~v_4235;
assign v_37424 = v_4235;
assign v_37425 = ~v_33535;
assign v_37426 = ~v_4239;
assign v_37427 = v_4239;
assign v_37428 = ~v_33539;
assign v_37429 = ~v_4243;
assign v_37430 = v_4243;
assign v_37431 = ~v_33543;
assign v_37432 = ~v_4247;
assign v_37433 = v_37432;
assign v_37435 = v_37434;
assign v_37437 = v_37429 & v_37436;
assign v_37439 = v_33539;
assign v_37441 = v_37438 & v_37440;
assign v_37443 = v_37426 & v_37442;
assign v_37445 = v_33535;
assign v_37447 = v_37444 & v_37446;
assign v_37449 = v_37423 & v_37448;
assign v_37451 = v_33531;
assign v_37453 = v_37450 & v_37452;
assign v_37455 = v_37420 & v_37454;
assign v_37457 = v_33527;
assign v_37459 = v_37456 & v_37458;
assign v_37461 = v_37417 & v_37460;
assign v_37463 = v_33523;
assign v_37465 = v_37462 & v_37464;
assign v_37467 = v_37414 & v_37466;
assign v_37469 = v_33519;
assign v_37471 = v_37468 & v_37470;
assign v_37473 = v_37411 & v_37472;
assign v_37475 = v_33515;
assign v_37477 = v_37474 & v_37476;
assign v_37479 = v_37408 & v_37478;
assign v_37481 = v_33511;
assign v_37483 = v_37480 & v_37482;
assign v_37485 = v_37405 & v_37484;
assign v_37487 = v_33507;
assign v_37489 = v_37486 & v_37488;
assign v_37491 = v_37402 & v_37490;
assign v_37493 = v_33503;
assign v_37495 = v_37492 & v_37494;
assign v_37497 = v_37399 & v_37496;
assign v_37499 = v_33499;
assign v_37501 = v_37498 & v_37500;
assign v_37503 = v_37396 & v_37502;
assign v_37505 = v_33495;
assign v_37507 = v_37504 & v_37506;
assign v_37509 = v_37393 & v_37508;
assign v_37511 = v_4194;
assign v_37513 = v_37510 & v_37512;
assign v_37515 = v_37390 & v_37514;
assign v_37517 = v_4190;
assign v_37519 = v_37516 & v_37518;
assign v_37521 = v_37387 & v_37520;
assign v_37523 = v_4186;
assign v_37525 = v_37522 & v_37524;
assign v_37527 = v_37384 & v_37526;
assign v_37529 = v_4182;
assign v_37531 = v_37528 & v_37530;
assign v_37533 = ~v_37532;
assign v_37535 = v_33543;
assign v_37536 = v_4247;
assign v_37537 = v_37536;
assign v_37538 = v_37535 & v_37537;
assign v_37539 = v_37538;
assign v_37540 = v_37429 & v_37539;
assign v_37542 = v_37439 & v_37541;
assign v_37543 = v_37428 & v_37539;
assign v_37545 = v_37426 & v_37544;
assign v_37547 = v_37445 & v_37546;
assign v_37548 = v_37425 & v_37544;
assign v_37550 = v_37423 & v_37549;
assign v_37552 = v_37451 & v_37551;
assign v_37553 = v_37422 & v_37549;
assign v_37555 = v_37420 & v_37554;
assign v_37557 = v_37457 & v_37556;
assign v_37558 = v_37419 & v_37554;
assign v_37560 = v_37417 & v_37559;
assign v_37562 = v_37463 & v_37561;
assign v_37563 = v_37416 & v_37559;
assign v_37565 = v_37414 & v_37564;
assign v_37567 = v_37469 & v_37566;
assign v_37568 = v_37413 & v_37564;
assign v_37570 = v_37411 & v_37569;
assign v_37572 = v_37475 & v_37571;
assign v_37573 = v_37410 & v_37569;
assign v_37575 = v_37408 & v_37574;
assign v_37577 = v_37481 & v_37576;
assign v_37578 = v_37407 & v_37574;
assign v_37580 = v_37405 & v_37579;
assign v_37582 = v_37487 & v_37581;
assign v_37583 = v_37404 & v_37579;
assign v_37585 = v_37402 & v_37584;
assign v_37587 = v_37493 & v_37586;
assign v_37588 = v_37401 & v_37584;
assign v_37590 = v_37399 & v_37589;
assign v_37592 = v_37499 & v_37591;
assign v_37593 = v_37398 & v_37589;
assign v_37595 = v_37396 & v_37594;
assign v_37597 = v_37505 & v_37596;
assign v_37598 = v_37395 & v_37594;
assign v_37600 = v_37393 & v_37599;
assign v_37602 = v_37511 & v_37601;
assign v_37603 = v_37392 & v_37599;
assign v_37605 = v_37390 & v_37604;
assign v_37607 = v_37517 & v_37606;
assign v_37608 = v_37389 & v_37604;
assign v_37610 = v_37387 & v_37609;
assign v_37612 = v_37523 & v_37611;
assign v_37613 = v_37386 & v_37609;
assign v_37615 = v_37384 & v_37614;
assign v_37617 = v_37529 & v_37616;
assign v_37618 = v_37383 & v_37614;
assign v_37620 = v_37532;
assign v_37622 = v_37534 & v_37621;
assign v_37623 = v_37622;
assign v_37625 = v_37624;
assign v_37627 = ~v_6;
assign v_37629 = ~v_37628;
assign v_37630 = v_37628;
assign v_37631 = ~v_13;
assign v_37633 = ~v_37632;
assign v_37634 = v_37632;
assign v_37635 = ~v_18;
assign v_37637 = ~v_37636;
assign v_37638 = v_37636;
assign v_37639 = ~v_23;
assign v_37641 = ~v_37640;
assign v_37642 = v_37640;
assign v_37644 = ~v_37643;
assign v_37645 = ~v_30;
assign v_37646 = v_30;
assign v_37648 = ~v_37647;
assign v_37649 = ~v_35;
assign v_37650 = v_35;
assign v_37652 = ~v_37651;
assign v_37653 = ~v_40;
assign v_37654 = v_40;
assign v_37656 = ~v_37655;
assign v_37657 = ~v_45;
assign v_37658 = v_45;
assign v_37660 = ~v_37659;
assign v_37661 = ~v_50;
assign v_37662 = v_50;
assign v_37664 = ~v_37663;
assign v_37665 = ~v_55;
assign v_37666 = v_55;
assign v_37668 = ~v_37667;
assign v_37669 = ~v_60;
assign v_37670 = v_60;
assign v_37672 = ~v_37671;
assign v_37673 = ~v_65;
assign v_37674 = v_65;
assign v_37676 = ~v_37675;
assign v_37677 = ~v_70;
assign v_37678 = v_70;
assign v_37680 = ~v_37679;
assign v_37681 = ~v_75;
assign v_37682 = v_75;
assign v_37684 = ~v_37683;
assign v_37685 = ~v_80;
assign v_37686 = v_80;
assign v_37688 = ~v_37687;
assign v_37689 = ~v_85;
assign v_37690 = v_85;
assign v_37692 = ~v_37691;
assign v_37693 = ~v_90;
assign v_37694 = v_37693;
assign v_37696 = v_37695;
assign v_37698 = v_37689 & v_37697;
assign v_37700 = v_37687;
assign v_37702 = v_37699 & v_37701;
assign v_37704 = v_37685 & v_37703;
assign v_37706 = v_37683;
assign v_37708 = v_37705 & v_37707;
assign v_37710 = v_37681 & v_37709;
assign v_37712 = v_37679;
assign v_37714 = v_37711 & v_37713;
assign v_37716 = v_37677 & v_37715;
assign v_37718 = v_37675;
assign v_37720 = v_37717 & v_37719;
assign v_37722 = v_37673 & v_37721;
assign v_37724 = v_37671;
assign v_37726 = v_37723 & v_37725;
assign v_37728 = v_37669 & v_37727;
assign v_37730 = v_37667;
assign v_37732 = v_37729 & v_37731;
assign v_37734 = v_37665 & v_37733;
assign v_37736 = v_37663;
assign v_37738 = v_37735 & v_37737;
assign v_37740 = v_37661 & v_37739;
assign v_37742 = v_37659;
assign v_37744 = v_37741 & v_37743;
assign v_37746 = v_37657 & v_37745;
assign v_37748 = v_37655;
assign v_37750 = v_37747 & v_37749;
assign v_37752 = v_37653 & v_37751;
assign v_37754 = v_37651;
assign v_37756 = v_37753 & v_37755;
assign v_37758 = v_37649 & v_37757;
assign v_37760 = v_37647;
assign v_37762 = v_37759 & v_37761;
assign v_37764 = v_37645 & v_37763;
assign v_37766 = v_37643;
assign v_37768 = v_37765 & v_37767;
assign v_37770 = v_37641 & v_37769;
assign v_37772 = v_23;
assign v_37774 = v_37771 & v_37773;
assign v_37776 = v_37637 & v_37775;
assign v_37778 = v_18;
assign v_37780 = v_37777 & v_37779;
assign v_37782 = v_37633 & v_37781;
assign v_37784 = v_13;
assign v_37786 = v_37783 & v_37785;
assign v_37788 = v_37629 & v_37787;
assign v_37790 = v_6;
assign v_37792 = v_37789 & v_37791;
assign v_37793 = v_37792;
assign v_37795 = v_37691;
assign v_37796 = v_90;
assign v_37797 = v_37796;
assign v_37798 = v_37795 & v_37797;
assign v_37799 = v_37798;
assign v_37800 = v_37689 & v_37799;
assign v_37802 = v_37700 & v_37801;
assign v_37803 = v_37688 & v_37799;
assign v_37805 = v_37685 & v_37804;
assign v_37807 = v_37706 & v_37806;
assign v_37808 = v_37684 & v_37804;
assign v_37810 = v_37681 & v_37809;
assign v_37812 = v_37712 & v_37811;
assign v_37813 = v_37680 & v_37809;
assign v_37815 = v_37677 & v_37814;
assign v_37817 = v_37718 & v_37816;
assign v_37818 = v_37676 & v_37814;
assign v_37820 = v_37673 & v_37819;
assign v_37822 = v_37724 & v_37821;
assign v_37823 = v_37672 & v_37819;
assign v_37825 = v_37669 & v_37824;
assign v_37827 = v_37730 & v_37826;
assign v_37828 = v_37668 & v_37824;
assign v_37830 = v_37665 & v_37829;
assign v_37832 = v_37736 & v_37831;
assign v_37833 = v_37664 & v_37829;
assign v_37835 = v_37661 & v_37834;
assign v_37837 = v_37742 & v_37836;
assign v_37838 = v_37660 & v_37834;
assign v_37840 = v_37657 & v_37839;
assign v_37842 = v_37748 & v_37841;
assign v_37843 = v_37656 & v_37839;
assign v_37845 = v_37653 & v_37844;
assign v_37847 = v_37754 & v_37846;
assign v_37848 = v_37652 & v_37844;
assign v_37850 = v_37649 & v_37849;
assign v_37852 = v_37760 & v_37851;
assign v_37853 = v_37648 & v_37849;
assign v_37855 = v_37645 & v_37854;
assign v_37857 = v_37766 & v_37856;
assign v_37858 = v_37644 & v_37854;
assign v_37860 = v_37641 & v_37859;
assign v_37862 = v_37772 & v_37861;
assign v_37863 = v_37639 & v_37859;
assign v_37865 = v_37637 & v_37864;
assign v_37867 = v_37778 & v_37866;
assign v_37868 = v_37635 & v_37864;
assign v_37870 = v_37633 & v_37869;
assign v_37872 = v_37784 & v_37871;
assign v_37873 = v_37631 & v_37869;
assign v_37875 = v_37629 & v_37874;
assign v_37877 = v_37790 & v_37876;
assign v_37878 = v_37627 & v_37874;
assign v_37880 = v_37879;
assign v_37882 = v_37794 & v_37881;
assign v_37883 = v_37882;
assign v_37885 = v_37884;
assign v_37887 = ~v_283;
assign v_37888 = ~v_37628;
assign v_37889 = v_37628;
assign v_37890 = ~v_287;
assign v_37891 = ~v_37632;
assign v_37892 = v_37632;
assign v_37893 = ~v_291;
assign v_37894 = ~v_37636;
assign v_37895 = v_37636;
assign v_37896 = ~v_295;
assign v_37897 = ~v_37640;
assign v_37898 = v_37640;
assign v_37899 = ~v_37643;
assign v_37900 = ~v_300;
assign v_37901 = v_300;
assign v_37902 = ~v_37647;
assign v_37903 = ~v_304;
assign v_37904 = v_304;
assign v_37905 = ~v_37651;
assign v_37906 = ~v_308;
assign v_37907 = v_308;
assign v_37908 = ~v_37655;
assign v_37909 = ~v_312;
assign v_37910 = v_312;
assign v_37911 = ~v_37659;
assign v_37912 = ~v_316;
assign v_37913 = v_316;
assign v_37914 = ~v_37663;
assign v_37915 = ~v_320;
assign v_37916 = v_320;
assign v_37917 = ~v_37667;
assign v_37918 = ~v_324;
assign v_37919 = v_324;
assign v_37920 = ~v_37671;
assign v_37921 = ~v_328;
assign v_37922 = v_328;
assign v_37923 = ~v_37675;
assign v_37924 = ~v_332;
assign v_37925 = v_332;
assign v_37926 = ~v_37679;
assign v_37927 = ~v_336;
assign v_37928 = v_336;
assign v_37929 = ~v_37683;
assign v_37930 = ~v_340;
assign v_37931 = v_340;
assign v_37932 = ~v_37687;
assign v_37933 = ~v_344;
assign v_37934 = v_344;
assign v_37935 = ~v_37691;
assign v_37936 = ~v_348;
assign v_37937 = v_37936;
assign v_37939 = v_37938;
assign v_37941 = v_37933 & v_37940;
assign v_37943 = v_37687;
assign v_37945 = v_37942 & v_37944;
assign v_37947 = v_37930 & v_37946;
assign v_37949 = v_37683;
assign v_37951 = v_37948 & v_37950;
assign v_37953 = v_37927 & v_37952;
assign v_37955 = v_37679;
assign v_37957 = v_37954 & v_37956;
assign v_37959 = v_37924 & v_37958;
assign v_37961 = v_37675;
assign v_37963 = v_37960 & v_37962;
assign v_37965 = v_37921 & v_37964;
assign v_37967 = v_37671;
assign v_37969 = v_37966 & v_37968;
assign v_37971 = v_37918 & v_37970;
assign v_37973 = v_37667;
assign v_37975 = v_37972 & v_37974;
assign v_37977 = v_37915 & v_37976;
assign v_37979 = v_37663;
assign v_37981 = v_37978 & v_37980;
assign v_37983 = v_37912 & v_37982;
assign v_37985 = v_37659;
assign v_37987 = v_37984 & v_37986;
assign v_37989 = v_37909 & v_37988;
assign v_37991 = v_37655;
assign v_37993 = v_37990 & v_37992;
assign v_37995 = v_37906 & v_37994;
assign v_37997 = v_37651;
assign v_37999 = v_37996 & v_37998;
assign v_38001 = v_37903 & v_38000;
assign v_38003 = v_37647;
assign v_38005 = v_38002 & v_38004;
assign v_38007 = v_37900 & v_38006;
assign v_38009 = v_37643;
assign v_38011 = v_38008 & v_38010;
assign v_38013 = v_37897 & v_38012;
assign v_38015 = v_295;
assign v_38017 = v_38014 & v_38016;
assign v_38019 = v_37894 & v_38018;
assign v_38021 = v_291;
assign v_38023 = v_38020 & v_38022;
assign v_38025 = v_37891 & v_38024;
assign v_38027 = v_287;
assign v_38029 = v_38026 & v_38028;
assign v_38031 = v_37888 & v_38030;
assign v_38033 = v_283;
assign v_38035 = v_38032 & v_38034;
assign v_38036 = v_38035;
assign v_38038 = v_37691;
assign v_38039 = v_348;
assign v_38040 = v_38039;
assign v_38041 = v_38038 & v_38040;
assign v_38042 = v_38041;
assign v_38043 = v_37933 & v_38042;
assign v_38045 = v_37943 & v_38044;
assign v_38046 = v_37932 & v_38042;
assign v_38048 = v_37930 & v_38047;
assign v_38050 = v_37949 & v_38049;
assign v_38051 = v_37929 & v_38047;
assign v_38053 = v_37927 & v_38052;
assign v_38055 = v_37955 & v_38054;
assign v_38056 = v_37926 & v_38052;
assign v_38058 = v_37924 & v_38057;
assign v_38060 = v_37961 & v_38059;
assign v_38061 = v_37923 & v_38057;
assign v_38063 = v_37921 & v_38062;
assign v_38065 = v_37967 & v_38064;
assign v_38066 = v_37920 & v_38062;
assign v_38068 = v_37918 & v_38067;
assign v_38070 = v_37973 & v_38069;
assign v_38071 = v_37917 & v_38067;
assign v_38073 = v_37915 & v_38072;
assign v_38075 = v_37979 & v_38074;
assign v_38076 = v_37914 & v_38072;
assign v_38078 = v_37912 & v_38077;
assign v_38080 = v_37985 & v_38079;
assign v_38081 = v_37911 & v_38077;
assign v_38083 = v_37909 & v_38082;
assign v_38085 = v_37991 & v_38084;
assign v_38086 = v_37908 & v_38082;
assign v_38088 = v_37906 & v_38087;
assign v_38090 = v_37997 & v_38089;
assign v_38091 = v_37905 & v_38087;
assign v_38093 = v_37903 & v_38092;
assign v_38095 = v_38003 & v_38094;
assign v_38096 = v_37902 & v_38092;
assign v_38098 = v_37900 & v_38097;
assign v_38100 = v_38009 & v_38099;
assign v_38101 = v_37899 & v_38097;
assign v_38103 = v_37897 & v_38102;
assign v_38105 = v_38015 & v_38104;
assign v_38106 = v_37896 & v_38102;
assign v_38108 = v_37894 & v_38107;
assign v_38110 = v_38021 & v_38109;
assign v_38111 = v_37893 & v_38107;
assign v_38113 = v_37891 & v_38112;
assign v_38115 = v_38027 & v_38114;
assign v_38116 = v_37890 & v_38112;
assign v_38118 = v_37888 & v_38117;
assign v_38120 = v_38033 & v_38119;
assign v_38121 = v_37887 & v_38117;
assign v_38123 = v_38122;
assign v_38125 = v_38037 & v_38124;
assign v_38126 = v_38125;
assign v_38128 = v_38127;
assign v_38130 = ~v_543;
assign v_38131 = ~v_37628;
assign v_38132 = v_37628;
assign v_38133 = ~v_547;
assign v_38134 = ~v_37632;
assign v_38135 = v_37632;
assign v_38136 = ~v_551;
assign v_38137 = ~v_37636;
assign v_38138 = v_37636;
assign v_38139 = ~v_555;
assign v_38140 = ~v_37640;
assign v_38141 = v_37640;
assign v_38142 = ~v_37643;
assign v_38143 = ~v_560;
assign v_38144 = v_560;
assign v_38145 = ~v_37647;
assign v_38146 = ~v_564;
assign v_38147 = v_564;
assign v_38148 = ~v_37651;
assign v_38149 = ~v_568;
assign v_38150 = v_568;
assign v_38151 = ~v_37655;
assign v_38152 = ~v_572;
assign v_38153 = v_572;
assign v_38154 = ~v_37659;
assign v_38155 = ~v_576;
assign v_38156 = v_576;
assign v_38157 = ~v_37663;
assign v_38158 = ~v_580;
assign v_38159 = v_580;
assign v_38160 = ~v_37667;
assign v_38161 = ~v_584;
assign v_38162 = v_584;
assign v_38163 = ~v_37671;
assign v_38164 = ~v_588;
assign v_38165 = v_588;
assign v_38166 = ~v_37675;
assign v_38167 = ~v_592;
assign v_38168 = v_592;
assign v_38169 = ~v_37679;
assign v_38170 = ~v_596;
assign v_38171 = v_596;
assign v_38172 = ~v_37683;
assign v_38173 = ~v_600;
assign v_38174 = v_600;
assign v_38175 = ~v_37687;
assign v_38176 = ~v_604;
assign v_38177 = v_604;
assign v_38178 = ~v_37691;
assign v_38179 = ~v_608;
assign v_38180 = v_38179;
assign v_38182 = v_38181;
assign v_38184 = v_38176 & v_38183;
assign v_38186 = v_37687;
assign v_38188 = v_38185 & v_38187;
assign v_38190 = v_38173 & v_38189;
assign v_38192 = v_37683;
assign v_38194 = v_38191 & v_38193;
assign v_38196 = v_38170 & v_38195;
assign v_38198 = v_37679;
assign v_38200 = v_38197 & v_38199;
assign v_38202 = v_38167 & v_38201;
assign v_38204 = v_37675;
assign v_38206 = v_38203 & v_38205;
assign v_38208 = v_38164 & v_38207;
assign v_38210 = v_37671;
assign v_38212 = v_38209 & v_38211;
assign v_38214 = v_38161 & v_38213;
assign v_38216 = v_37667;
assign v_38218 = v_38215 & v_38217;
assign v_38220 = v_38158 & v_38219;
assign v_38222 = v_37663;
assign v_38224 = v_38221 & v_38223;
assign v_38226 = v_38155 & v_38225;
assign v_38228 = v_37659;
assign v_38230 = v_38227 & v_38229;
assign v_38232 = v_38152 & v_38231;
assign v_38234 = v_37655;
assign v_38236 = v_38233 & v_38235;
assign v_38238 = v_38149 & v_38237;
assign v_38240 = v_37651;
assign v_38242 = v_38239 & v_38241;
assign v_38244 = v_38146 & v_38243;
assign v_38246 = v_37647;
assign v_38248 = v_38245 & v_38247;
assign v_38250 = v_38143 & v_38249;
assign v_38252 = v_37643;
assign v_38254 = v_38251 & v_38253;
assign v_38256 = v_38140 & v_38255;
assign v_38258 = v_555;
assign v_38260 = v_38257 & v_38259;
assign v_38262 = v_38137 & v_38261;
assign v_38264 = v_551;
assign v_38266 = v_38263 & v_38265;
assign v_38268 = v_38134 & v_38267;
assign v_38270 = v_547;
assign v_38272 = v_38269 & v_38271;
assign v_38274 = v_38131 & v_38273;
assign v_38276 = v_543;
assign v_38278 = v_38275 & v_38277;
assign v_38279 = v_38278;
assign v_38281 = v_37691;
assign v_38282 = v_608;
assign v_38283 = v_38282;
assign v_38284 = v_38281 & v_38283;
assign v_38285 = v_38284;
assign v_38286 = v_38176 & v_38285;
assign v_38288 = v_38186 & v_38287;
assign v_38289 = v_38175 & v_38285;
assign v_38291 = v_38173 & v_38290;
assign v_38293 = v_38192 & v_38292;
assign v_38294 = v_38172 & v_38290;
assign v_38296 = v_38170 & v_38295;
assign v_38298 = v_38198 & v_38297;
assign v_38299 = v_38169 & v_38295;
assign v_38301 = v_38167 & v_38300;
assign v_38303 = v_38204 & v_38302;
assign v_38304 = v_38166 & v_38300;
assign v_38306 = v_38164 & v_38305;
assign v_38308 = v_38210 & v_38307;
assign v_38309 = v_38163 & v_38305;
assign v_38311 = v_38161 & v_38310;
assign v_38313 = v_38216 & v_38312;
assign v_38314 = v_38160 & v_38310;
assign v_38316 = v_38158 & v_38315;
assign v_38318 = v_38222 & v_38317;
assign v_38319 = v_38157 & v_38315;
assign v_38321 = v_38155 & v_38320;
assign v_38323 = v_38228 & v_38322;
assign v_38324 = v_38154 & v_38320;
assign v_38326 = v_38152 & v_38325;
assign v_38328 = v_38234 & v_38327;
assign v_38329 = v_38151 & v_38325;
assign v_38331 = v_38149 & v_38330;
assign v_38333 = v_38240 & v_38332;
assign v_38334 = v_38148 & v_38330;
assign v_38336 = v_38146 & v_38335;
assign v_38338 = v_38246 & v_38337;
assign v_38339 = v_38145 & v_38335;
assign v_38341 = v_38143 & v_38340;
assign v_38343 = v_38252 & v_38342;
assign v_38344 = v_38142 & v_38340;
assign v_38346 = v_38140 & v_38345;
assign v_38348 = v_38258 & v_38347;
assign v_38349 = v_38139 & v_38345;
assign v_38351 = v_38137 & v_38350;
assign v_38353 = v_38264 & v_38352;
assign v_38354 = v_38136 & v_38350;
assign v_38356 = v_38134 & v_38355;
assign v_38358 = v_38270 & v_38357;
assign v_38359 = v_38133 & v_38355;
assign v_38361 = v_38131 & v_38360;
assign v_38363 = v_38276 & v_38362;
assign v_38364 = v_38130 & v_38360;
assign v_38366 = v_38365;
assign v_38368 = v_38280 & v_38367;
assign v_38369 = v_38368;
assign v_38371 = v_38370;
assign v_38373 = ~v_803;
assign v_38374 = ~v_37628;
assign v_38375 = v_37628;
assign v_38376 = ~v_807;
assign v_38377 = ~v_37632;
assign v_38378 = v_37632;
assign v_38379 = ~v_811;
assign v_38380 = ~v_37636;
assign v_38381 = v_37636;
assign v_38382 = ~v_815;
assign v_38383 = ~v_37640;
assign v_38384 = v_37640;
assign v_38385 = ~v_37643;
assign v_38386 = ~v_820;
assign v_38387 = v_820;
assign v_38388 = ~v_37647;
assign v_38389 = ~v_824;
assign v_38390 = v_824;
assign v_38391 = ~v_37651;
assign v_38392 = ~v_828;
assign v_38393 = v_828;
assign v_38394 = ~v_37655;
assign v_38395 = ~v_832;
assign v_38396 = v_832;
assign v_38397 = ~v_37659;
assign v_38398 = ~v_836;
assign v_38399 = v_836;
assign v_38400 = ~v_37663;
assign v_38401 = ~v_840;
assign v_38402 = v_840;
assign v_38403 = ~v_37667;
assign v_38404 = ~v_844;
assign v_38405 = v_844;
assign v_38406 = ~v_37671;
assign v_38407 = ~v_848;
assign v_38408 = v_848;
assign v_38409 = ~v_37675;
assign v_38410 = ~v_852;
assign v_38411 = v_852;
assign v_38412 = ~v_37679;
assign v_38413 = ~v_856;
assign v_38414 = v_856;
assign v_38415 = ~v_37683;
assign v_38416 = ~v_860;
assign v_38417 = v_860;
assign v_38418 = ~v_37687;
assign v_38419 = ~v_864;
assign v_38420 = v_864;
assign v_38421 = ~v_37691;
assign v_38422 = ~v_868;
assign v_38423 = v_38422;
assign v_38425 = v_38424;
assign v_38427 = v_38419 & v_38426;
assign v_38429 = v_37687;
assign v_38431 = v_38428 & v_38430;
assign v_38433 = v_38416 & v_38432;
assign v_38435 = v_37683;
assign v_38437 = v_38434 & v_38436;
assign v_38439 = v_38413 & v_38438;
assign v_38441 = v_37679;
assign v_38443 = v_38440 & v_38442;
assign v_38445 = v_38410 & v_38444;
assign v_38447 = v_37675;
assign v_38449 = v_38446 & v_38448;
assign v_38451 = v_38407 & v_38450;
assign v_38453 = v_37671;
assign v_38455 = v_38452 & v_38454;
assign v_38457 = v_38404 & v_38456;
assign v_38459 = v_37667;
assign v_38461 = v_38458 & v_38460;
assign v_38463 = v_38401 & v_38462;
assign v_38465 = v_37663;
assign v_38467 = v_38464 & v_38466;
assign v_38469 = v_38398 & v_38468;
assign v_38471 = v_37659;
assign v_38473 = v_38470 & v_38472;
assign v_38475 = v_38395 & v_38474;
assign v_38477 = v_37655;
assign v_38479 = v_38476 & v_38478;
assign v_38481 = v_38392 & v_38480;
assign v_38483 = v_37651;
assign v_38485 = v_38482 & v_38484;
assign v_38487 = v_38389 & v_38486;
assign v_38489 = v_37647;
assign v_38491 = v_38488 & v_38490;
assign v_38493 = v_38386 & v_38492;
assign v_38495 = v_37643;
assign v_38497 = v_38494 & v_38496;
assign v_38499 = v_38383 & v_38498;
assign v_38501 = v_815;
assign v_38503 = v_38500 & v_38502;
assign v_38505 = v_38380 & v_38504;
assign v_38507 = v_811;
assign v_38509 = v_38506 & v_38508;
assign v_38511 = v_38377 & v_38510;
assign v_38513 = v_807;
assign v_38515 = v_38512 & v_38514;
assign v_38517 = v_38374 & v_38516;
assign v_38519 = v_803;
assign v_38521 = v_38518 & v_38520;
assign v_38522 = v_38521;
assign v_38524 = v_37691;
assign v_38525 = v_868;
assign v_38526 = v_38525;
assign v_38527 = v_38524 & v_38526;
assign v_38528 = v_38527;
assign v_38529 = v_38419 & v_38528;
assign v_38531 = v_38429 & v_38530;
assign v_38532 = v_38418 & v_38528;
assign v_38534 = v_38416 & v_38533;
assign v_38536 = v_38435 & v_38535;
assign v_38537 = v_38415 & v_38533;
assign v_38539 = v_38413 & v_38538;
assign v_38541 = v_38441 & v_38540;
assign v_38542 = v_38412 & v_38538;
assign v_38544 = v_38410 & v_38543;
assign v_38546 = v_38447 & v_38545;
assign v_38547 = v_38409 & v_38543;
assign v_38549 = v_38407 & v_38548;
assign v_38551 = v_38453 & v_38550;
assign v_38552 = v_38406 & v_38548;
assign v_38554 = v_38404 & v_38553;
assign v_38556 = v_38459 & v_38555;
assign v_38557 = v_38403 & v_38553;
assign v_38559 = v_38401 & v_38558;
assign v_38561 = v_38465 & v_38560;
assign v_38562 = v_38400 & v_38558;
assign v_38564 = v_38398 & v_38563;
assign v_38566 = v_38471 & v_38565;
assign v_38567 = v_38397 & v_38563;
assign v_38569 = v_38395 & v_38568;
assign v_38571 = v_38477 & v_38570;
assign v_38572 = v_38394 & v_38568;
assign v_38574 = v_38392 & v_38573;
assign v_38576 = v_38483 & v_38575;
assign v_38577 = v_38391 & v_38573;
assign v_38579 = v_38389 & v_38578;
assign v_38581 = v_38489 & v_38580;
assign v_38582 = v_38388 & v_38578;
assign v_38584 = v_38386 & v_38583;
assign v_38586 = v_38495 & v_38585;
assign v_38587 = v_38385 & v_38583;
assign v_38589 = v_38383 & v_38588;
assign v_38591 = v_38501 & v_38590;
assign v_38592 = v_38382 & v_38588;
assign v_38594 = v_38380 & v_38593;
assign v_38596 = v_38507 & v_38595;
assign v_38597 = v_38379 & v_38593;
assign v_38599 = v_38377 & v_38598;
assign v_38601 = v_38513 & v_38600;
assign v_38602 = v_38376 & v_38598;
assign v_38604 = v_38374 & v_38603;
assign v_38606 = v_38519 & v_38605;
assign v_38607 = v_38373 & v_38603;
assign v_38609 = v_38608;
assign v_38611 = v_38523 & v_38610;
assign v_38612 = v_38611;
assign v_38614 = v_38613;
assign v_38616 = ~v_1063;
assign v_38617 = ~v_37628;
assign v_38618 = v_37628;
assign v_38619 = ~v_1067;
assign v_38620 = ~v_37632;
assign v_38621 = v_37632;
assign v_38622 = ~v_1071;
assign v_38623 = ~v_37636;
assign v_38624 = v_37636;
assign v_38625 = ~v_1075;
assign v_38626 = ~v_37640;
assign v_38627 = v_37640;
assign v_38628 = ~v_37643;
assign v_38629 = ~v_1080;
assign v_38630 = v_1080;
assign v_38631 = ~v_37647;
assign v_38632 = ~v_1084;
assign v_38633 = v_1084;
assign v_38634 = ~v_37651;
assign v_38635 = ~v_1088;
assign v_38636 = v_1088;
assign v_38637 = ~v_37655;
assign v_38638 = ~v_1092;
assign v_38639 = v_1092;
assign v_38640 = ~v_37659;
assign v_38641 = ~v_1096;
assign v_38642 = v_1096;
assign v_38643 = ~v_37663;
assign v_38644 = ~v_1100;
assign v_38645 = v_1100;
assign v_38646 = ~v_37667;
assign v_38647 = ~v_1104;
assign v_38648 = v_1104;
assign v_38649 = ~v_37671;
assign v_38650 = ~v_1108;
assign v_38651 = v_1108;
assign v_38652 = ~v_37675;
assign v_38653 = ~v_1112;
assign v_38654 = v_1112;
assign v_38655 = ~v_37679;
assign v_38656 = ~v_1116;
assign v_38657 = v_1116;
assign v_38658 = ~v_37683;
assign v_38659 = ~v_1120;
assign v_38660 = v_1120;
assign v_38661 = ~v_37687;
assign v_38662 = ~v_1124;
assign v_38663 = v_1124;
assign v_38664 = ~v_37691;
assign v_38665 = ~v_1128;
assign v_38666 = v_38665;
assign v_38668 = v_38667;
assign v_38670 = v_38662 & v_38669;
assign v_38672 = v_37687;
assign v_38674 = v_38671 & v_38673;
assign v_38676 = v_38659 & v_38675;
assign v_38678 = v_37683;
assign v_38680 = v_38677 & v_38679;
assign v_38682 = v_38656 & v_38681;
assign v_38684 = v_37679;
assign v_38686 = v_38683 & v_38685;
assign v_38688 = v_38653 & v_38687;
assign v_38690 = v_37675;
assign v_38692 = v_38689 & v_38691;
assign v_38694 = v_38650 & v_38693;
assign v_38696 = v_37671;
assign v_38698 = v_38695 & v_38697;
assign v_38700 = v_38647 & v_38699;
assign v_38702 = v_37667;
assign v_38704 = v_38701 & v_38703;
assign v_38706 = v_38644 & v_38705;
assign v_38708 = v_37663;
assign v_38710 = v_38707 & v_38709;
assign v_38712 = v_38641 & v_38711;
assign v_38714 = v_37659;
assign v_38716 = v_38713 & v_38715;
assign v_38718 = v_38638 & v_38717;
assign v_38720 = v_37655;
assign v_38722 = v_38719 & v_38721;
assign v_38724 = v_38635 & v_38723;
assign v_38726 = v_37651;
assign v_38728 = v_38725 & v_38727;
assign v_38730 = v_38632 & v_38729;
assign v_38732 = v_37647;
assign v_38734 = v_38731 & v_38733;
assign v_38736 = v_38629 & v_38735;
assign v_38738 = v_37643;
assign v_38740 = v_38737 & v_38739;
assign v_38742 = v_38626 & v_38741;
assign v_38744 = v_1075;
assign v_38746 = v_38743 & v_38745;
assign v_38748 = v_38623 & v_38747;
assign v_38750 = v_1071;
assign v_38752 = v_38749 & v_38751;
assign v_38754 = v_38620 & v_38753;
assign v_38756 = v_1067;
assign v_38758 = v_38755 & v_38757;
assign v_38760 = v_38617 & v_38759;
assign v_38762 = v_1063;
assign v_38764 = v_38761 & v_38763;
assign v_38765 = v_38764;
assign v_38767 = v_37691;
assign v_38768 = v_1128;
assign v_38769 = v_38768;
assign v_38770 = v_38767 & v_38769;
assign v_38771 = v_38770;
assign v_38772 = v_38662 & v_38771;
assign v_38774 = v_38672 & v_38773;
assign v_38775 = v_38661 & v_38771;
assign v_38777 = v_38659 & v_38776;
assign v_38779 = v_38678 & v_38778;
assign v_38780 = v_38658 & v_38776;
assign v_38782 = v_38656 & v_38781;
assign v_38784 = v_38684 & v_38783;
assign v_38785 = v_38655 & v_38781;
assign v_38787 = v_38653 & v_38786;
assign v_38789 = v_38690 & v_38788;
assign v_38790 = v_38652 & v_38786;
assign v_38792 = v_38650 & v_38791;
assign v_38794 = v_38696 & v_38793;
assign v_38795 = v_38649 & v_38791;
assign v_38797 = v_38647 & v_38796;
assign v_38799 = v_38702 & v_38798;
assign v_38800 = v_38646 & v_38796;
assign v_38802 = v_38644 & v_38801;
assign v_38804 = v_38708 & v_38803;
assign v_38805 = v_38643 & v_38801;
assign v_38807 = v_38641 & v_38806;
assign v_38809 = v_38714 & v_38808;
assign v_38810 = v_38640 & v_38806;
assign v_38812 = v_38638 & v_38811;
assign v_38814 = v_38720 & v_38813;
assign v_38815 = v_38637 & v_38811;
assign v_38817 = v_38635 & v_38816;
assign v_38819 = v_38726 & v_38818;
assign v_38820 = v_38634 & v_38816;
assign v_38822 = v_38632 & v_38821;
assign v_38824 = v_38732 & v_38823;
assign v_38825 = v_38631 & v_38821;
assign v_38827 = v_38629 & v_38826;
assign v_38829 = v_38738 & v_38828;
assign v_38830 = v_38628 & v_38826;
assign v_38832 = v_38626 & v_38831;
assign v_38834 = v_38744 & v_38833;
assign v_38835 = v_38625 & v_38831;
assign v_38837 = v_38623 & v_38836;
assign v_38839 = v_38750 & v_38838;
assign v_38840 = v_38622 & v_38836;
assign v_38842 = v_38620 & v_38841;
assign v_38844 = v_38756 & v_38843;
assign v_38845 = v_38619 & v_38841;
assign v_38847 = v_38617 & v_38846;
assign v_38849 = v_38762 & v_38848;
assign v_38850 = v_38616 & v_38846;
assign v_38852 = v_38851;
assign v_38854 = v_38766 & v_38853;
assign v_38855 = v_38854;
assign v_38857 = v_38856;
assign v_38859 = ~v_1323;
assign v_38860 = ~v_37628;
assign v_38861 = v_37628;
assign v_38862 = ~v_1327;
assign v_38863 = ~v_37632;
assign v_38864 = v_37632;
assign v_38865 = ~v_1331;
assign v_38866 = ~v_37636;
assign v_38867 = v_37636;
assign v_38868 = ~v_1335;
assign v_38869 = ~v_37640;
assign v_38870 = v_37640;
assign v_38871 = ~v_37643;
assign v_38872 = ~v_1340;
assign v_38873 = v_1340;
assign v_38874 = ~v_37647;
assign v_38875 = ~v_1344;
assign v_38876 = v_1344;
assign v_38877 = ~v_37651;
assign v_38878 = ~v_1348;
assign v_38879 = v_1348;
assign v_38880 = ~v_37655;
assign v_38881 = ~v_1352;
assign v_38882 = v_1352;
assign v_38883 = ~v_37659;
assign v_38884 = ~v_1356;
assign v_38885 = v_1356;
assign v_38886 = ~v_37663;
assign v_38887 = ~v_1360;
assign v_38888 = v_1360;
assign v_38889 = ~v_37667;
assign v_38890 = ~v_1364;
assign v_38891 = v_1364;
assign v_38892 = ~v_37671;
assign v_38893 = ~v_1368;
assign v_38894 = v_1368;
assign v_38895 = ~v_37675;
assign v_38896 = ~v_1372;
assign v_38897 = v_1372;
assign v_38898 = ~v_37679;
assign v_38899 = ~v_1376;
assign v_38900 = v_1376;
assign v_38901 = ~v_37683;
assign v_38902 = ~v_1380;
assign v_38903 = v_1380;
assign v_38904 = ~v_37687;
assign v_38905 = ~v_1384;
assign v_38906 = v_1384;
assign v_38907 = ~v_37691;
assign v_38908 = ~v_1388;
assign v_38909 = v_38908;
assign v_38911 = v_38910;
assign v_38913 = v_38905 & v_38912;
assign v_38915 = v_37687;
assign v_38917 = v_38914 & v_38916;
assign v_38919 = v_38902 & v_38918;
assign v_38921 = v_37683;
assign v_38923 = v_38920 & v_38922;
assign v_38925 = v_38899 & v_38924;
assign v_38927 = v_37679;
assign v_38929 = v_38926 & v_38928;
assign v_38931 = v_38896 & v_38930;
assign v_38933 = v_37675;
assign v_38935 = v_38932 & v_38934;
assign v_38937 = v_38893 & v_38936;
assign v_38939 = v_37671;
assign v_38941 = v_38938 & v_38940;
assign v_38943 = v_38890 & v_38942;
assign v_38945 = v_37667;
assign v_38947 = v_38944 & v_38946;
assign v_38949 = v_38887 & v_38948;
assign v_38951 = v_37663;
assign v_38953 = v_38950 & v_38952;
assign v_38955 = v_38884 & v_38954;
assign v_38957 = v_37659;
assign v_38959 = v_38956 & v_38958;
assign v_38961 = v_38881 & v_38960;
assign v_38963 = v_37655;
assign v_38965 = v_38962 & v_38964;
assign v_38967 = v_38878 & v_38966;
assign v_38969 = v_37651;
assign v_38971 = v_38968 & v_38970;
assign v_38973 = v_38875 & v_38972;
assign v_38975 = v_37647;
assign v_38977 = v_38974 & v_38976;
assign v_38979 = v_38872 & v_38978;
assign v_38981 = v_37643;
assign v_38983 = v_38980 & v_38982;
assign v_38985 = v_38869 & v_38984;
assign v_38987 = v_1335;
assign v_38989 = v_38986 & v_38988;
assign v_38991 = v_38866 & v_38990;
assign v_38993 = v_1331;
assign v_38995 = v_38992 & v_38994;
assign v_38997 = v_38863 & v_38996;
assign v_38999 = v_1327;
assign v_39001 = v_38998 & v_39000;
assign v_39003 = v_38860 & v_39002;
assign v_39005 = v_1323;
assign v_39007 = v_39004 & v_39006;
assign v_39008 = v_39007;
assign v_39010 = v_37691;
assign v_39011 = v_1388;
assign v_39012 = v_39011;
assign v_39013 = v_39010 & v_39012;
assign v_39014 = v_39013;
assign v_39015 = v_38905 & v_39014;
assign v_39017 = v_38915 & v_39016;
assign v_39018 = v_38904 & v_39014;
assign v_39020 = v_38902 & v_39019;
assign v_39022 = v_38921 & v_39021;
assign v_39023 = v_38901 & v_39019;
assign v_39025 = v_38899 & v_39024;
assign v_39027 = v_38927 & v_39026;
assign v_39028 = v_38898 & v_39024;
assign v_39030 = v_38896 & v_39029;
assign v_39032 = v_38933 & v_39031;
assign v_39033 = v_38895 & v_39029;
assign v_39035 = v_38893 & v_39034;
assign v_39037 = v_38939 & v_39036;
assign v_39038 = v_38892 & v_39034;
assign v_39040 = v_38890 & v_39039;
assign v_39042 = v_38945 & v_39041;
assign v_39043 = v_38889 & v_39039;
assign v_39045 = v_38887 & v_39044;
assign v_39047 = v_38951 & v_39046;
assign v_39048 = v_38886 & v_39044;
assign v_39050 = v_38884 & v_39049;
assign v_39052 = v_38957 & v_39051;
assign v_39053 = v_38883 & v_39049;
assign v_39055 = v_38881 & v_39054;
assign v_39057 = v_38963 & v_39056;
assign v_39058 = v_38880 & v_39054;
assign v_39060 = v_38878 & v_39059;
assign v_39062 = v_38969 & v_39061;
assign v_39063 = v_38877 & v_39059;
assign v_39065 = v_38875 & v_39064;
assign v_39067 = v_38975 & v_39066;
assign v_39068 = v_38874 & v_39064;
assign v_39070 = v_38872 & v_39069;
assign v_39072 = v_38981 & v_39071;
assign v_39073 = v_38871 & v_39069;
assign v_39075 = v_38869 & v_39074;
assign v_39077 = v_38987 & v_39076;
assign v_39078 = v_38868 & v_39074;
assign v_39080 = v_38866 & v_39079;
assign v_39082 = v_38993 & v_39081;
assign v_39083 = v_38865 & v_39079;
assign v_39085 = v_38863 & v_39084;
assign v_39087 = v_38999 & v_39086;
assign v_39088 = v_38862 & v_39084;
assign v_39090 = v_38860 & v_39089;
assign v_39092 = v_39005 & v_39091;
assign v_39093 = v_38859 & v_39089;
assign v_39095 = v_39094;
assign v_39097 = v_39009 & v_39096;
assign v_39098 = v_39097;
assign v_39100 = v_39099;
assign v_39102 = ~v_1583;
assign v_39103 = ~v_37628;
assign v_39104 = v_37628;
assign v_39105 = ~v_1587;
assign v_39106 = ~v_37632;
assign v_39107 = v_37632;
assign v_39108 = ~v_1591;
assign v_39109 = ~v_37636;
assign v_39110 = v_37636;
assign v_39111 = ~v_1595;
assign v_39112 = ~v_37640;
assign v_39113 = v_37640;
assign v_39114 = ~v_37643;
assign v_39115 = ~v_1600;
assign v_39116 = v_1600;
assign v_39117 = ~v_37647;
assign v_39118 = ~v_1604;
assign v_39119 = v_1604;
assign v_39120 = ~v_37651;
assign v_39121 = ~v_1608;
assign v_39122 = v_1608;
assign v_39123 = ~v_37655;
assign v_39124 = ~v_1612;
assign v_39125 = v_1612;
assign v_39126 = ~v_37659;
assign v_39127 = ~v_1616;
assign v_39128 = v_1616;
assign v_39129 = ~v_37663;
assign v_39130 = ~v_1620;
assign v_39131 = v_1620;
assign v_39132 = ~v_37667;
assign v_39133 = ~v_1624;
assign v_39134 = v_1624;
assign v_39135 = ~v_37671;
assign v_39136 = ~v_1628;
assign v_39137 = v_1628;
assign v_39138 = ~v_37675;
assign v_39139 = ~v_1632;
assign v_39140 = v_1632;
assign v_39141 = ~v_37679;
assign v_39142 = ~v_1636;
assign v_39143 = v_1636;
assign v_39144 = ~v_37683;
assign v_39145 = ~v_1640;
assign v_39146 = v_1640;
assign v_39147 = ~v_37687;
assign v_39148 = ~v_1644;
assign v_39149 = v_1644;
assign v_39150 = ~v_37691;
assign v_39151 = ~v_1648;
assign v_39152 = v_39151;
assign v_39154 = v_39153;
assign v_39156 = v_39148 & v_39155;
assign v_39158 = v_37687;
assign v_39160 = v_39157 & v_39159;
assign v_39162 = v_39145 & v_39161;
assign v_39164 = v_37683;
assign v_39166 = v_39163 & v_39165;
assign v_39168 = v_39142 & v_39167;
assign v_39170 = v_37679;
assign v_39172 = v_39169 & v_39171;
assign v_39174 = v_39139 & v_39173;
assign v_39176 = v_37675;
assign v_39178 = v_39175 & v_39177;
assign v_39180 = v_39136 & v_39179;
assign v_39182 = v_37671;
assign v_39184 = v_39181 & v_39183;
assign v_39186 = v_39133 & v_39185;
assign v_39188 = v_37667;
assign v_39190 = v_39187 & v_39189;
assign v_39192 = v_39130 & v_39191;
assign v_39194 = v_37663;
assign v_39196 = v_39193 & v_39195;
assign v_39198 = v_39127 & v_39197;
assign v_39200 = v_37659;
assign v_39202 = v_39199 & v_39201;
assign v_39204 = v_39124 & v_39203;
assign v_39206 = v_37655;
assign v_39208 = v_39205 & v_39207;
assign v_39210 = v_39121 & v_39209;
assign v_39212 = v_37651;
assign v_39214 = v_39211 & v_39213;
assign v_39216 = v_39118 & v_39215;
assign v_39218 = v_37647;
assign v_39220 = v_39217 & v_39219;
assign v_39222 = v_39115 & v_39221;
assign v_39224 = v_37643;
assign v_39226 = v_39223 & v_39225;
assign v_39228 = v_39112 & v_39227;
assign v_39230 = v_1595;
assign v_39232 = v_39229 & v_39231;
assign v_39234 = v_39109 & v_39233;
assign v_39236 = v_1591;
assign v_39238 = v_39235 & v_39237;
assign v_39240 = v_39106 & v_39239;
assign v_39242 = v_1587;
assign v_39244 = v_39241 & v_39243;
assign v_39246 = v_39103 & v_39245;
assign v_39248 = v_1583;
assign v_39250 = v_39247 & v_39249;
assign v_39251 = v_39250;
assign v_39253 = v_37691;
assign v_39254 = v_1648;
assign v_39255 = v_39254;
assign v_39256 = v_39253 & v_39255;
assign v_39257 = v_39256;
assign v_39258 = v_39148 & v_39257;
assign v_39260 = v_39158 & v_39259;
assign v_39261 = v_39147 & v_39257;
assign v_39263 = v_39145 & v_39262;
assign v_39265 = v_39164 & v_39264;
assign v_39266 = v_39144 & v_39262;
assign v_39268 = v_39142 & v_39267;
assign v_39270 = v_39170 & v_39269;
assign v_39271 = v_39141 & v_39267;
assign v_39273 = v_39139 & v_39272;
assign v_39275 = v_39176 & v_39274;
assign v_39276 = v_39138 & v_39272;
assign v_39278 = v_39136 & v_39277;
assign v_39280 = v_39182 & v_39279;
assign v_39281 = v_39135 & v_39277;
assign v_39283 = v_39133 & v_39282;
assign v_39285 = v_39188 & v_39284;
assign v_39286 = v_39132 & v_39282;
assign v_39288 = v_39130 & v_39287;
assign v_39290 = v_39194 & v_39289;
assign v_39291 = v_39129 & v_39287;
assign v_39293 = v_39127 & v_39292;
assign v_39295 = v_39200 & v_39294;
assign v_39296 = v_39126 & v_39292;
assign v_39298 = v_39124 & v_39297;
assign v_39300 = v_39206 & v_39299;
assign v_39301 = v_39123 & v_39297;
assign v_39303 = v_39121 & v_39302;
assign v_39305 = v_39212 & v_39304;
assign v_39306 = v_39120 & v_39302;
assign v_39308 = v_39118 & v_39307;
assign v_39310 = v_39218 & v_39309;
assign v_39311 = v_39117 & v_39307;
assign v_39313 = v_39115 & v_39312;
assign v_39315 = v_39224 & v_39314;
assign v_39316 = v_39114 & v_39312;
assign v_39318 = v_39112 & v_39317;
assign v_39320 = v_39230 & v_39319;
assign v_39321 = v_39111 & v_39317;
assign v_39323 = v_39109 & v_39322;
assign v_39325 = v_39236 & v_39324;
assign v_39326 = v_39108 & v_39322;
assign v_39328 = v_39106 & v_39327;
assign v_39330 = v_39242 & v_39329;
assign v_39331 = v_39105 & v_39327;
assign v_39333 = v_39103 & v_39332;
assign v_39335 = v_39248 & v_39334;
assign v_39336 = v_39102 & v_39332;
assign v_39338 = v_39337;
assign v_39340 = v_39252 & v_39339;
assign v_39341 = v_39340;
assign v_39343 = v_39342;
assign v_39345 = ~v_1843;
assign v_39346 = ~v_37628;
assign v_39347 = v_37628;
assign v_39348 = ~v_1847;
assign v_39349 = ~v_37632;
assign v_39350 = v_37632;
assign v_39351 = ~v_1851;
assign v_39352 = ~v_37636;
assign v_39353 = v_37636;
assign v_39354 = ~v_1855;
assign v_39355 = ~v_37640;
assign v_39356 = v_37640;
assign v_39357 = ~v_37643;
assign v_39358 = ~v_1860;
assign v_39359 = v_1860;
assign v_39360 = ~v_37647;
assign v_39361 = ~v_1864;
assign v_39362 = v_1864;
assign v_39363 = ~v_37651;
assign v_39364 = ~v_1868;
assign v_39365 = v_1868;
assign v_39366 = ~v_37655;
assign v_39367 = ~v_1872;
assign v_39368 = v_1872;
assign v_39369 = ~v_37659;
assign v_39370 = ~v_1876;
assign v_39371 = v_1876;
assign v_39372 = ~v_37663;
assign v_39373 = ~v_1880;
assign v_39374 = v_1880;
assign v_39375 = ~v_37667;
assign v_39376 = ~v_1884;
assign v_39377 = v_1884;
assign v_39378 = ~v_37671;
assign v_39379 = ~v_1888;
assign v_39380 = v_1888;
assign v_39381 = ~v_37675;
assign v_39382 = ~v_1892;
assign v_39383 = v_1892;
assign v_39384 = ~v_37679;
assign v_39385 = ~v_1896;
assign v_39386 = v_1896;
assign v_39387 = ~v_37683;
assign v_39388 = ~v_1900;
assign v_39389 = v_1900;
assign v_39390 = ~v_37687;
assign v_39391 = ~v_1904;
assign v_39392 = v_1904;
assign v_39393 = ~v_37691;
assign v_39394 = ~v_1908;
assign v_39395 = v_39394;
assign v_39397 = v_39396;
assign v_39399 = v_39391 & v_39398;
assign v_39401 = v_37687;
assign v_39403 = v_39400 & v_39402;
assign v_39405 = v_39388 & v_39404;
assign v_39407 = v_37683;
assign v_39409 = v_39406 & v_39408;
assign v_39411 = v_39385 & v_39410;
assign v_39413 = v_37679;
assign v_39415 = v_39412 & v_39414;
assign v_39417 = v_39382 & v_39416;
assign v_39419 = v_37675;
assign v_39421 = v_39418 & v_39420;
assign v_39423 = v_39379 & v_39422;
assign v_39425 = v_37671;
assign v_39427 = v_39424 & v_39426;
assign v_39429 = v_39376 & v_39428;
assign v_39431 = v_37667;
assign v_39433 = v_39430 & v_39432;
assign v_39435 = v_39373 & v_39434;
assign v_39437 = v_37663;
assign v_39439 = v_39436 & v_39438;
assign v_39441 = v_39370 & v_39440;
assign v_39443 = v_37659;
assign v_39445 = v_39442 & v_39444;
assign v_39447 = v_39367 & v_39446;
assign v_39449 = v_37655;
assign v_39451 = v_39448 & v_39450;
assign v_39453 = v_39364 & v_39452;
assign v_39455 = v_37651;
assign v_39457 = v_39454 & v_39456;
assign v_39459 = v_39361 & v_39458;
assign v_39461 = v_37647;
assign v_39463 = v_39460 & v_39462;
assign v_39465 = v_39358 & v_39464;
assign v_39467 = v_37643;
assign v_39469 = v_39466 & v_39468;
assign v_39471 = v_39355 & v_39470;
assign v_39473 = v_1855;
assign v_39475 = v_39472 & v_39474;
assign v_39477 = v_39352 & v_39476;
assign v_39479 = v_1851;
assign v_39481 = v_39478 & v_39480;
assign v_39483 = v_39349 & v_39482;
assign v_39485 = v_1847;
assign v_39487 = v_39484 & v_39486;
assign v_39489 = v_39346 & v_39488;
assign v_39491 = v_1843;
assign v_39493 = v_39490 & v_39492;
assign v_39494 = v_39493;
assign v_39496 = v_37691;
assign v_39497 = v_1908;
assign v_39498 = v_39497;
assign v_39499 = v_39496 & v_39498;
assign v_39500 = v_39499;
assign v_39501 = v_39391 & v_39500;
assign v_39503 = v_39401 & v_39502;
assign v_39504 = v_39390 & v_39500;
assign v_39506 = v_39388 & v_39505;
assign v_39508 = v_39407 & v_39507;
assign v_39509 = v_39387 & v_39505;
assign v_39511 = v_39385 & v_39510;
assign v_39513 = v_39413 & v_39512;
assign v_39514 = v_39384 & v_39510;
assign v_39516 = v_39382 & v_39515;
assign v_39518 = v_39419 & v_39517;
assign v_39519 = v_39381 & v_39515;
assign v_39521 = v_39379 & v_39520;
assign v_39523 = v_39425 & v_39522;
assign v_39524 = v_39378 & v_39520;
assign v_39526 = v_39376 & v_39525;
assign v_39528 = v_39431 & v_39527;
assign v_39529 = v_39375 & v_39525;
assign v_39531 = v_39373 & v_39530;
assign v_39533 = v_39437 & v_39532;
assign v_39534 = v_39372 & v_39530;
assign v_39536 = v_39370 & v_39535;
assign v_39538 = v_39443 & v_39537;
assign v_39539 = v_39369 & v_39535;
assign v_39541 = v_39367 & v_39540;
assign v_39543 = v_39449 & v_39542;
assign v_39544 = v_39366 & v_39540;
assign v_39546 = v_39364 & v_39545;
assign v_39548 = v_39455 & v_39547;
assign v_39549 = v_39363 & v_39545;
assign v_39551 = v_39361 & v_39550;
assign v_39553 = v_39461 & v_39552;
assign v_39554 = v_39360 & v_39550;
assign v_39556 = v_39358 & v_39555;
assign v_39558 = v_39467 & v_39557;
assign v_39559 = v_39357 & v_39555;
assign v_39561 = v_39355 & v_39560;
assign v_39563 = v_39473 & v_39562;
assign v_39564 = v_39354 & v_39560;
assign v_39566 = v_39352 & v_39565;
assign v_39568 = v_39479 & v_39567;
assign v_39569 = v_39351 & v_39565;
assign v_39571 = v_39349 & v_39570;
assign v_39573 = v_39485 & v_39572;
assign v_39574 = v_39348 & v_39570;
assign v_39576 = v_39346 & v_39575;
assign v_39578 = v_39491 & v_39577;
assign v_39579 = v_39345 & v_39575;
assign v_39581 = v_39580;
assign v_39583 = v_39495 & v_39582;
assign v_39584 = v_39583;
assign v_39586 = v_39585;
assign v_39588 = ~v_2103;
assign v_39589 = ~v_37628;
assign v_39590 = v_37628;
assign v_39591 = ~v_2107;
assign v_39592 = ~v_37632;
assign v_39593 = v_37632;
assign v_39594 = ~v_2111;
assign v_39595 = ~v_37636;
assign v_39596 = v_37636;
assign v_39597 = ~v_2115;
assign v_39598 = ~v_37640;
assign v_39599 = v_37640;
assign v_39600 = ~v_37643;
assign v_39601 = ~v_2120;
assign v_39602 = v_2120;
assign v_39603 = ~v_37647;
assign v_39604 = ~v_2124;
assign v_39605 = v_2124;
assign v_39606 = ~v_37651;
assign v_39607 = ~v_2128;
assign v_39608 = v_2128;
assign v_39609 = ~v_37655;
assign v_39610 = ~v_2132;
assign v_39611 = v_2132;
assign v_39612 = ~v_37659;
assign v_39613 = ~v_2136;
assign v_39614 = v_2136;
assign v_39615 = ~v_37663;
assign v_39616 = ~v_2140;
assign v_39617 = v_2140;
assign v_39618 = ~v_37667;
assign v_39619 = ~v_2144;
assign v_39620 = v_2144;
assign v_39621 = ~v_37671;
assign v_39622 = ~v_2148;
assign v_39623 = v_2148;
assign v_39624 = ~v_37675;
assign v_39625 = ~v_2152;
assign v_39626 = v_2152;
assign v_39627 = ~v_37679;
assign v_39628 = ~v_2156;
assign v_39629 = v_2156;
assign v_39630 = ~v_37683;
assign v_39631 = ~v_2160;
assign v_39632 = v_2160;
assign v_39633 = ~v_37687;
assign v_39634 = ~v_2164;
assign v_39635 = v_2164;
assign v_39636 = ~v_37691;
assign v_39637 = ~v_2168;
assign v_39638 = v_39637;
assign v_39640 = v_39639;
assign v_39642 = v_39634 & v_39641;
assign v_39644 = v_37687;
assign v_39646 = v_39643 & v_39645;
assign v_39648 = v_39631 & v_39647;
assign v_39650 = v_37683;
assign v_39652 = v_39649 & v_39651;
assign v_39654 = v_39628 & v_39653;
assign v_39656 = v_37679;
assign v_39658 = v_39655 & v_39657;
assign v_39660 = v_39625 & v_39659;
assign v_39662 = v_37675;
assign v_39664 = v_39661 & v_39663;
assign v_39666 = v_39622 & v_39665;
assign v_39668 = v_37671;
assign v_39670 = v_39667 & v_39669;
assign v_39672 = v_39619 & v_39671;
assign v_39674 = v_37667;
assign v_39676 = v_39673 & v_39675;
assign v_39678 = v_39616 & v_39677;
assign v_39680 = v_37663;
assign v_39682 = v_39679 & v_39681;
assign v_39684 = v_39613 & v_39683;
assign v_39686 = v_37659;
assign v_39688 = v_39685 & v_39687;
assign v_39690 = v_39610 & v_39689;
assign v_39692 = v_37655;
assign v_39694 = v_39691 & v_39693;
assign v_39696 = v_39607 & v_39695;
assign v_39698 = v_37651;
assign v_39700 = v_39697 & v_39699;
assign v_39702 = v_39604 & v_39701;
assign v_39704 = v_37647;
assign v_39706 = v_39703 & v_39705;
assign v_39708 = v_39601 & v_39707;
assign v_39710 = v_37643;
assign v_39712 = v_39709 & v_39711;
assign v_39714 = v_39598 & v_39713;
assign v_39716 = v_2115;
assign v_39718 = v_39715 & v_39717;
assign v_39720 = v_39595 & v_39719;
assign v_39722 = v_2111;
assign v_39724 = v_39721 & v_39723;
assign v_39726 = v_39592 & v_39725;
assign v_39728 = v_2107;
assign v_39730 = v_39727 & v_39729;
assign v_39732 = v_39589 & v_39731;
assign v_39734 = v_2103;
assign v_39736 = v_39733 & v_39735;
assign v_39737 = v_39736;
assign v_39739 = v_37691;
assign v_39740 = v_2168;
assign v_39741 = v_39740;
assign v_39742 = v_39739 & v_39741;
assign v_39743 = v_39742;
assign v_39744 = v_39634 & v_39743;
assign v_39746 = v_39644 & v_39745;
assign v_39747 = v_39633 & v_39743;
assign v_39749 = v_39631 & v_39748;
assign v_39751 = v_39650 & v_39750;
assign v_39752 = v_39630 & v_39748;
assign v_39754 = v_39628 & v_39753;
assign v_39756 = v_39656 & v_39755;
assign v_39757 = v_39627 & v_39753;
assign v_39759 = v_39625 & v_39758;
assign v_39761 = v_39662 & v_39760;
assign v_39762 = v_39624 & v_39758;
assign v_39764 = v_39622 & v_39763;
assign v_39766 = v_39668 & v_39765;
assign v_39767 = v_39621 & v_39763;
assign v_39769 = v_39619 & v_39768;
assign v_39771 = v_39674 & v_39770;
assign v_39772 = v_39618 & v_39768;
assign v_39774 = v_39616 & v_39773;
assign v_39776 = v_39680 & v_39775;
assign v_39777 = v_39615 & v_39773;
assign v_39779 = v_39613 & v_39778;
assign v_39781 = v_39686 & v_39780;
assign v_39782 = v_39612 & v_39778;
assign v_39784 = v_39610 & v_39783;
assign v_39786 = v_39692 & v_39785;
assign v_39787 = v_39609 & v_39783;
assign v_39789 = v_39607 & v_39788;
assign v_39791 = v_39698 & v_39790;
assign v_39792 = v_39606 & v_39788;
assign v_39794 = v_39604 & v_39793;
assign v_39796 = v_39704 & v_39795;
assign v_39797 = v_39603 & v_39793;
assign v_39799 = v_39601 & v_39798;
assign v_39801 = v_39710 & v_39800;
assign v_39802 = v_39600 & v_39798;
assign v_39804 = v_39598 & v_39803;
assign v_39806 = v_39716 & v_39805;
assign v_39807 = v_39597 & v_39803;
assign v_39809 = v_39595 & v_39808;
assign v_39811 = v_39722 & v_39810;
assign v_39812 = v_39594 & v_39808;
assign v_39814 = v_39592 & v_39813;
assign v_39816 = v_39728 & v_39815;
assign v_39817 = v_39591 & v_39813;
assign v_39819 = v_39589 & v_39818;
assign v_39821 = v_39734 & v_39820;
assign v_39822 = v_39588 & v_39818;
assign v_39824 = v_39823;
assign v_39826 = v_39738 & v_39825;
assign v_39827 = v_39826;
assign v_39829 = v_39828;
assign v_39831 = ~v_2363;
assign v_39832 = ~v_37628;
assign v_39833 = v_37628;
assign v_39834 = ~v_2367;
assign v_39835 = ~v_37632;
assign v_39836 = v_37632;
assign v_39837 = ~v_2371;
assign v_39838 = ~v_37636;
assign v_39839 = v_37636;
assign v_39840 = ~v_2375;
assign v_39841 = ~v_37640;
assign v_39842 = v_37640;
assign v_39843 = ~v_37643;
assign v_39844 = ~v_2380;
assign v_39845 = v_2380;
assign v_39846 = ~v_37647;
assign v_39847 = ~v_2384;
assign v_39848 = v_2384;
assign v_39849 = ~v_37651;
assign v_39850 = ~v_2388;
assign v_39851 = v_2388;
assign v_39852 = ~v_37655;
assign v_39853 = ~v_2392;
assign v_39854 = v_2392;
assign v_39855 = ~v_37659;
assign v_39856 = ~v_2396;
assign v_39857 = v_2396;
assign v_39858 = ~v_37663;
assign v_39859 = ~v_2400;
assign v_39860 = v_2400;
assign v_39861 = ~v_37667;
assign v_39862 = ~v_2404;
assign v_39863 = v_2404;
assign v_39864 = ~v_37671;
assign v_39865 = ~v_2408;
assign v_39866 = v_2408;
assign v_39867 = ~v_37675;
assign v_39868 = ~v_2412;
assign v_39869 = v_2412;
assign v_39870 = ~v_37679;
assign v_39871 = ~v_2416;
assign v_39872 = v_2416;
assign v_39873 = ~v_37683;
assign v_39874 = ~v_2420;
assign v_39875 = v_2420;
assign v_39876 = ~v_37687;
assign v_39877 = ~v_2424;
assign v_39878 = v_2424;
assign v_39879 = ~v_37691;
assign v_39880 = ~v_2428;
assign v_39881 = v_39880;
assign v_39883 = v_39882;
assign v_39885 = v_39877 & v_39884;
assign v_39887 = v_37687;
assign v_39889 = v_39886 & v_39888;
assign v_39891 = v_39874 & v_39890;
assign v_39893 = v_37683;
assign v_39895 = v_39892 & v_39894;
assign v_39897 = v_39871 & v_39896;
assign v_39899 = v_37679;
assign v_39901 = v_39898 & v_39900;
assign v_39903 = v_39868 & v_39902;
assign v_39905 = v_37675;
assign v_39907 = v_39904 & v_39906;
assign v_39909 = v_39865 & v_39908;
assign v_39911 = v_37671;
assign v_39913 = v_39910 & v_39912;
assign v_39915 = v_39862 & v_39914;
assign v_39917 = v_37667;
assign v_39919 = v_39916 & v_39918;
assign v_39921 = v_39859 & v_39920;
assign v_39923 = v_37663;
assign v_39925 = v_39922 & v_39924;
assign v_39927 = v_39856 & v_39926;
assign v_39929 = v_37659;
assign v_39931 = v_39928 & v_39930;
assign v_39933 = v_39853 & v_39932;
assign v_39935 = v_37655;
assign v_39937 = v_39934 & v_39936;
assign v_39939 = v_39850 & v_39938;
assign v_39941 = v_37651;
assign v_39943 = v_39940 & v_39942;
assign v_39945 = v_39847 & v_39944;
assign v_39947 = v_37647;
assign v_39949 = v_39946 & v_39948;
assign v_39951 = v_39844 & v_39950;
assign v_39953 = v_37643;
assign v_39955 = v_39952 & v_39954;
assign v_39957 = v_39841 & v_39956;
assign v_39959 = v_2375;
assign v_39961 = v_39958 & v_39960;
assign v_39963 = v_39838 & v_39962;
assign v_39965 = v_2371;
assign v_39967 = v_39964 & v_39966;
assign v_39969 = v_39835 & v_39968;
assign v_39971 = v_2367;
assign v_39973 = v_39970 & v_39972;
assign v_39975 = v_39832 & v_39974;
assign v_39977 = v_2363;
assign v_39979 = v_39976 & v_39978;
assign v_39980 = v_39979;
assign v_39982 = v_37691;
assign v_39983 = v_2428;
assign v_39984 = v_39983;
assign v_39985 = v_39982 & v_39984;
assign v_39986 = v_39985;
assign v_39987 = v_39877 & v_39986;
assign v_39989 = v_39887 & v_39988;
assign v_39990 = v_39876 & v_39986;
assign v_39992 = v_39874 & v_39991;
assign v_39994 = v_39893 & v_39993;
assign v_39995 = v_39873 & v_39991;
assign v_39997 = v_39871 & v_39996;
assign v_39999 = v_39899 & v_39998;
assign v_40000 = v_39870 & v_39996;
assign v_40002 = v_39868 & v_40001;
assign v_40004 = v_39905 & v_40003;
assign v_40005 = v_39867 & v_40001;
assign v_40007 = v_39865 & v_40006;
assign v_40009 = v_39911 & v_40008;
assign v_40010 = v_39864 & v_40006;
assign v_40012 = v_39862 & v_40011;
assign v_40014 = v_39917 & v_40013;
assign v_40015 = v_39861 & v_40011;
assign v_40017 = v_39859 & v_40016;
assign v_40019 = v_39923 & v_40018;
assign v_40020 = v_39858 & v_40016;
assign v_40022 = v_39856 & v_40021;
assign v_40024 = v_39929 & v_40023;
assign v_40025 = v_39855 & v_40021;
assign v_40027 = v_39853 & v_40026;
assign v_40029 = v_39935 & v_40028;
assign v_40030 = v_39852 & v_40026;
assign v_40032 = v_39850 & v_40031;
assign v_40034 = v_39941 & v_40033;
assign v_40035 = v_39849 & v_40031;
assign v_40037 = v_39847 & v_40036;
assign v_40039 = v_39947 & v_40038;
assign v_40040 = v_39846 & v_40036;
assign v_40042 = v_39844 & v_40041;
assign v_40044 = v_39953 & v_40043;
assign v_40045 = v_39843 & v_40041;
assign v_40047 = v_39841 & v_40046;
assign v_40049 = v_39959 & v_40048;
assign v_40050 = v_39840 & v_40046;
assign v_40052 = v_39838 & v_40051;
assign v_40054 = v_39965 & v_40053;
assign v_40055 = v_39837 & v_40051;
assign v_40057 = v_39835 & v_40056;
assign v_40059 = v_39971 & v_40058;
assign v_40060 = v_39834 & v_40056;
assign v_40062 = v_39832 & v_40061;
assign v_40064 = v_39977 & v_40063;
assign v_40065 = v_39831 & v_40061;
assign v_40067 = v_40066;
assign v_40069 = v_39981 & v_40068;
assign v_40070 = v_40069;
assign v_40072 = v_40071;
assign v_40074 = ~v_2623;
assign v_40075 = ~v_37628;
assign v_40076 = v_37628;
assign v_40077 = ~v_2627;
assign v_40078 = ~v_37632;
assign v_40079 = v_37632;
assign v_40080 = ~v_2631;
assign v_40081 = ~v_37636;
assign v_40082 = v_37636;
assign v_40083 = ~v_2635;
assign v_40084 = ~v_37640;
assign v_40085 = v_37640;
assign v_40086 = ~v_37643;
assign v_40087 = ~v_2640;
assign v_40088 = v_2640;
assign v_40089 = ~v_37647;
assign v_40090 = ~v_2644;
assign v_40091 = v_2644;
assign v_40092 = ~v_37651;
assign v_40093 = ~v_2648;
assign v_40094 = v_2648;
assign v_40095 = ~v_37655;
assign v_40096 = ~v_2652;
assign v_40097 = v_2652;
assign v_40098 = ~v_37659;
assign v_40099 = ~v_2656;
assign v_40100 = v_2656;
assign v_40101 = ~v_37663;
assign v_40102 = ~v_2660;
assign v_40103 = v_2660;
assign v_40104 = ~v_37667;
assign v_40105 = ~v_2664;
assign v_40106 = v_2664;
assign v_40107 = ~v_37671;
assign v_40108 = ~v_2668;
assign v_40109 = v_2668;
assign v_40110 = ~v_37675;
assign v_40111 = ~v_2672;
assign v_40112 = v_2672;
assign v_40113 = ~v_37679;
assign v_40114 = ~v_2676;
assign v_40115 = v_2676;
assign v_40116 = ~v_37683;
assign v_40117 = ~v_2680;
assign v_40118 = v_2680;
assign v_40119 = ~v_37687;
assign v_40120 = ~v_2684;
assign v_40121 = v_2684;
assign v_40122 = ~v_37691;
assign v_40123 = ~v_2688;
assign v_40124 = v_40123;
assign v_40126 = v_40125;
assign v_40128 = v_40120 & v_40127;
assign v_40130 = v_37687;
assign v_40132 = v_40129 & v_40131;
assign v_40134 = v_40117 & v_40133;
assign v_40136 = v_37683;
assign v_40138 = v_40135 & v_40137;
assign v_40140 = v_40114 & v_40139;
assign v_40142 = v_37679;
assign v_40144 = v_40141 & v_40143;
assign v_40146 = v_40111 & v_40145;
assign v_40148 = v_37675;
assign v_40150 = v_40147 & v_40149;
assign v_40152 = v_40108 & v_40151;
assign v_40154 = v_37671;
assign v_40156 = v_40153 & v_40155;
assign v_40158 = v_40105 & v_40157;
assign v_40160 = v_37667;
assign v_40162 = v_40159 & v_40161;
assign v_40164 = v_40102 & v_40163;
assign v_40166 = v_37663;
assign v_40168 = v_40165 & v_40167;
assign v_40170 = v_40099 & v_40169;
assign v_40172 = v_37659;
assign v_40174 = v_40171 & v_40173;
assign v_40176 = v_40096 & v_40175;
assign v_40178 = v_37655;
assign v_40180 = v_40177 & v_40179;
assign v_40182 = v_40093 & v_40181;
assign v_40184 = v_37651;
assign v_40186 = v_40183 & v_40185;
assign v_40188 = v_40090 & v_40187;
assign v_40190 = v_37647;
assign v_40192 = v_40189 & v_40191;
assign v_40194 = v_40087 & v_40193;
assign v_40196 = v_37643;
assign v_40198 = v_40195 & v_40197;
assign v_40200 = v_40084 & v_40199;
assign v_40202 = v_2635;
assign v_40204 = v_40201 & v_40203;
assign v_40206 = v_40081 & v_40205;
assign v_40208 = v_2631;
assign v_40210 = v_40207 & v_40209;
assign v_40212 = v_40078 & v_40211;
assign v_40214 = v_2627;
assign v_40216 = v_40213 & v_40215;
assign v_40218 = v_40075 & v_40217;
assign v_40220 = v_2623;
assign v_40222 = v_40219 & v_40221;
assign v_40223 = v_40222;
assign v_40225 = v_37691;
assign v_40226 = v_2688;
assign v_40227 = v_40226;
assign v_40228 = v_40225 & v_40227;
assign v_40229 = v_40228;
assign v_40230 = v_40120 & v_40229;
assign v_40232 = v_40130 & v_40231;
assign v_40233 = v_40119 & v_40229;
assign v_40235 = v_40117 & v_40234;
assign v_40237 = v_40136 & v_40236;
assign v_40238 = v_40116 & v_40234;
assign v_40240 = v_40114 & v_40239;
assign v_40242 = v_40142 & v_40241;
assign v_40243 = v_40113 & v_40239;
assign v_40245 = v_40111 & v_40244;
assign v_40247 = v_40148 & v_40246;
assign v_40248 = v_40110 & v_40244;
assign v_40250 = v_40108 & v_40249;
assign v_40252 = v_40154 & v_40251;
assign v_40253 = v_40107 & v_40249;
assign v_40255 = v_40105 & v_40254;
assign v_40257 = v_40160 & v_40256;
assign v_40258 = v_40104 & v_40254;
assign v_40260 = v_40102 & v_40259;
assign v_40262 = v_40166 & v_40261;
assign v_40263 = v_40101 & v_40259;
assign v_40265 = v_40099 & v_40264;
assign v_40267 = v_40172 & v_40266;
assign v_40268 = v_40098 & v_40264;
assign v_40270 = v_40096 & v_40269;
assign v_40272 = v_40178 & v_40271;
assign v_40273 = v_40095 & v_40269;
assign v_40275 = v_40093 & v_40274;
assign v_40277 = v_40184 & v_40276;
assign v_40278 = v_40092 & v_40274;
assign v_40280 = v_40090 & v_40279;
assign v_40282 = v_40190 & v_40281;
assign v_40283 = v_40089 & v_40279;
assign v_40285 = v_40087 & v_40284;
assign v_40287 = v_40196 & v_40286;
assign v_40288 = v_40086 & v_40284;
assign v_40290 = v_40084 & v_40289;
assign v_40292 = v_40202 & v_40291;
assign v_40293 = v_40083 & v_40289;
assign v_40295 = v_40081 & v_40294;
assign v_40297 = v_40208 & v_40296;
assign v_40298 = v_40080 & v_40294;
assign v_40300 = v_40078 & v_40299;
assign v_40302 = v_40214 & v_40301;
assign v_40303 = v_40077 & v_40299;
assign v_40305 = v_40075 & v_40304;
assign v_40307 = v_40220 & v_40306;
assign v_40308 = v_40074 & v_40304;
assign v_40310 = v_40309;
assign v_40312 = v_40224 & v_40311;
assign v_40313 = v_40312;
assign v_40315 = v_40314;
assign v_40317 = ~v_2883;
assign v_40318 = ~v_37628;
assign v_40319 = v_37628;
assign v_40320 = ~v_2887;
assign v_40321 = ~v_37632;
assign v_40322 = v_37632;
assign v_40323 = ~v_2891;
assign v_40324 = ~v_37636;
assign v_40325 = v_37636;
assign v_40326 = ~v_2895;
assign v_40327 = ~v_37640;
assign v_40328 = v_37640;
assign v_40329 = ~v_37643;
assign v_40330 = ~v_2900;
assign v_40331 = v_2900;
assign v_40332 = ~v_37647;
assign v_40333 = ~v_2904;
assign v_40334 = v_2904;
assign v_40335 = ~v_37651;
assign v_40336 = ~v_2908;
assign v_40337 = v_2908;
assign v_40338 = ~v_37655;
assign v_40339 = ~v_2912;
assign v_40340 = v_2912;
assign v_40341 = ~v_37659;
assign v_40342 = ~v_2916;
assign v_40343 = v_2916;
assign v_40344 = ~v_37663;
assign v_40345 = ~v_2920;
assign v_40346 = v_2920;
assign v_40347 = ~v_37667;
assign v_40348 = ~v_2924;
assign v_40349 = v_2924;
assign v_40350 = ~v_37671;
assign v_40351 = ~v_2928;
assign v_40352 = v_2928;
assign v_40353 = ~v_37675;
assign v_40354 = ~v_2932;
assign v_40355 = v_2932;
assign v_40356 = ~v_37679;
assign v_40357 = ~v_2936;
assign v_40358 = v_2936;
assign v_40359 = ~v_37683;
assign v_40360 = ~v_2940;
assign v_40361 = v_2940;
assign v_40362 = ~v_37687;
assign v_40363 = ~v_2944;
assign v_40364 = v_2944;
assign v_40365 = ~v_37691;
assign v_40366 = ~v_2948;
assign v_40367 = v_40366;
assign v_40369 = v_40368;
assign v_40371 = v_40363 & v_40370;
assign v_40373 = v_37687;
assign v_40375 = v_40372 & v_40374;
assign v_40377 = v_40360 & v_40376;
assign v_40379 = v_37683;
assign v_40381 = v_40378 & v_40380;
assign v_40383 = v_40357 & v_40382;
assign v_40385 = v_37679;
assign v_40387 = v_40384 & v_40386;
assign v_40389 = v_40354 & v_40388;
assign v_40391 = v_37675;
assign v_40393 = v_40390 & v_40392;
assign v_40395 = v_40351 & v_40394;
assign v_40397 = v_37671;
assign v_40399 = v_40396 & v_40398;
assign v_40401 = v_40348 & v_40400;
assign v_40403 = v_37667;
assign v_40405 = v_40402 & v_40404;
assign v_40407 = v_40345 & v_40406;
assign v_40409 = v_37663;
assign v_40411 = v_40408 & v_40410;
assign v_40413 = v_40342 & v_40412;
assign v_40415 = v_37659;
assign v_40417 = v_40414 & v_40416;
assign v_40419 = v_40339 & v_40418;
assign v_40421 = v_37655;
assign v_40423 = v_40420 & v_40422;
assign v_40425 = v_40336 & v_40424;
assign v_40427 = v_37651;
assign v_40429 = v_40426 & v_40428;
assign v_40431 = v_40333 & v_40430;
assign v_40433 = v_37647;
assign v_40435 = v_40432 & v_40434;
assign v_40437 = v_40330 & v_40436;
assign v_40439 = v_37643;
assign v_40441 = v_40438 & v_40440;
assign v_40443 = v_40327 & v_40442;
assign v_40445 = v_2895;
assign v_40447 = v_40444 & v_40446;
assign v_40449 = v_40324 & v_40448;
assign v_40451 = v_2891;
assign v_40453 = v_40450 & v_40452;
assign v_40455 = v_40321 & v_40454;
assign v_40457 = v_2887;
assign v_40459 = v_40456 & v_40458;
assign v_40461 = v_40318 & v_40460;
assign v_40463 = v_2883;
assign v_40465 = v_40462 & v_40464;
assign v_40466 = v_40465;
assign v_40468 = v_37691;
assign v_40469 = v_2948;
assign v_40470 = v_40469;
assign v_40471 = v_40468 & v_40470;
assign v_40472 = v_40471;
assign v_40473 = v_40363 & v_40472;
assign v_40475 = v_40373 & v_40474;
assign v_40476 = v_40362 & v_40472;
assign v_40478 = v_40360 & v_40477;
assign v_40480 = v_40379 & v_40479;
assign v_40481 = v_40359 & v_40477;
assign v_40483 = v_40357 & v_40482;
assign v_40485 = v_40385 & v_40484;
assign v_40486 = v_40356 & v_40482;
assign v_40488 = v_40354 & v_40487;
assign v_40490 = v_40391 & v_40489;
assign v_40491 = v_40353 & v_40487;
assign v_40493 = v_40351 & v_40492;
assign v_40495 = v_40397 & v_40494;
assign v_40496 = v_40350 & v_40492;
assign v_40498 = v_40348 & v_40497;
assign v_40500 = v_40403 & v_40499;
assign v_40501 = v_40347 & v_40497;
assign v_40503 = v_40345 & v_40502;
assign v_40505 = v_40409 & v_40504;
assign v_40506 = v_40344 & v_40502;
assign v_40508 = v_40342 & v_40507;
assign v_40510 = v_40415 & v_40509;
assign v_40511 = v_40341 & v_40507;
assign v_40513 = v_40339 & v_40512;
assign v_40515 = v_40421 & v_40514;
assign v_40516 = v_40338 & v_40512;
assign v_40518 = v_40336 & v_40517;
assign v_40520 = v_40427 & v_40519;
assign v_40521 = v_40335 & v_40517;
assign v_40523 = v_40333 & v_40522;
assign v_40525 = v_40433 & v_40524;
assign v_40526 = v_40332 & v_40522;
assign v_40528 = v_40330 & v_40527;
assign v_40530 = v_40439 & v_40529;
assign v_40531 = v_40329 & v_40527;
assign v_40533 = v_40327 & v_40532;
assign v_40535 = v_40445 & v_40534;
assign v_40536 = v_40326 & v_40532;
assign v_40538 = v_40324 & v_40537;
assign v_40540 = v_40451 & v_40539;
assign v_40541 = v_40323 & v_40537;
assign v_40543 = v_40321 & v_40542;
assign v_40545 = v_40457 & v_40544;
assign v_40546 = v_40320 & v_40542;
assign v_40548 = v_40318 & v_40547;
assign v_40550 = v_40463 & v_40549;
assign v_40551 = v_40317 & v_40547;
assign v_40553 = v_40552;
assign v_40555 = v_40467 & v_40554;
assign v_40556 = v_40555;
assign v_40558 = v_40557;
assign v_40560 = ~v_3143;
assign v_40561 = ~v_37628;
assign v_40562 = v_37628;
assign v_40563 = ~v_3147;
assign v_40564 = ~v_37632;
assign v_40565 = v_37632;
assign v_40566 = ~v_3151;
assign v_40567 = ~v_37636;
assign v_40568 = v_37636;
assign v_40569 = ~v_3155;
assign v_40570 = ~v_37640;
assign v_40571 = v_37640;
assign v_40572 = ~v_37643;
assign v_40573 = ~v_3160;
assign v_40574 = v_3160;
assign v_40575 = ~v_37647;
assign v_40576 = ~v_3164;
assign v_40577 = v_3164;
assign v_40578 = ~v_37651;
assign v_40579 = ~v_3168;
assign v_40580 = v_3168;
assign v_40581 = ~v_37655;
assign v_40582 = ~v_3172;
assign v_40583 = v_3172;
assign v_40584 = ~v_37659;
assign v_40585 = ~v_3176;
assign v_40586 = v_3176;
assign v_40587 = ~v_37663;
assign v_40588 = ~v_3180;
assign v_40589 = v_3180;
assign v_40590 = ~v_37667;
assign v_40591 = ~v_3184;
assign v_40592 = v_3184;
assign v_40593 = ~v_37671;
assign v_40594 = ~v_3188;
assign v_40595 = v_3188;
assign v_40596 = ~v_37675;
assign v_40597 = ~v_3192;
assign v_40598 = v_3192;
assign v_40599 = ~v_37679;
assign v_40600 = ~v_3196;
assign v_40601 = v_3196;
assign v_40602 = ~v_37683;
assign v_40603 = ~v_3200;
assign v_40604 = v_3200;
assign v_40605 = ~v_37687;
assign v_40606 = ~v_3204;
assign v_40607 = v_3204;
assign v_40608 = ~v_37691;
assign v_40609 = ~v_3208;
assign v_40610 = v_40609;
assign v_40612 = v_40611;
assign v_40614 = v_40606 & v_40613;
assign v_40616 = v_37687;
assign v_40618 = v_40615 & v_40617;
assign v_40620 = v_40603 & v_40619;
assign v_40622 = v_37683;
assign v_40624 = v_40621 & v_40623;
assign v_40626 = v_40600 & v_40625;
assign v_40628 = v_37679;
assign v_40630 = v_40627 & v_40629;
assign v_40632 = v_40597 & v_40631;
assign v_40634 = v_37675;
assign v_40636 = v_40633 & v_40635;
assign v_40638 = v_40594 & v_40637;
assign v_40640 = v_37671;
assign v_40642 = v_40639 & v_40641;
assign v_40644 = v_40591 & v_40643;
assign v_40646 = v_37667;
assign v_40648 = v_40645 & v_40647;
assign v_40650 = v_40588 & v_40649;
assign v_40652 = v_37663;
assign v_40654 = v_40651 & v_40653;
assign v_40656 = v_40585 & v_40655;
assign v_40658 = v_37659;
assign v_40660 = v_40657 & v_40659;
assign v_40662 = v_40582 & v_40661;
assign v_40664 = v_37655;
assign v_40666 = v_40663 & v_40665;
assign v_40668 = v_40579 & v_40667;
assign v_40670 = v_37651;
assign v_40672 = v_40669 & v_40671;
assign v_40674 = v_40576 & v_40673;
assign v_40676 = v_37647;
assign v_40678 = v_40675 & v_40677;
assign v_40680 = v_40573 & v_40679;
assign v_40682 = v_37643;
assign v_40684 = v_40681 & v_40683;
assign v_40686 = v_40570 & v_40685;
assign v_40688 = v_3155;
assign v_40690 = v_40687 & v_40689;
assign v_40692 = v_40567 & v_40691;
assign v_40694 = v_3151;
assign v_40696 = v_40693 & v_40695;
assign v_40698 = v_40564 & v_40697;
assign v_40700 = v_3147;
assign v_40702 = v_40699 & v_40701;
assign v_40704 = v_40561 & v_40703;
assign v_40706 = v_3143;
assign v_40708 = v_40705 & v_40707;
assign v_40709 = v_40708;
assign v_40711 = v_37691;
assign v_40712 = v_3208;
assign v_40713 = v_40712;
assign v_40714 = v_40711 & v_40713;
assign v_40715 = v_40714;
assign v_40716 = v_40606 & v_40715;
assign v_40718 = v_40616 & v_40717;
assign v_40719 = v_40605 & v_40715;
assign v_40721 = v_40603 & v_40720;
assign v_40723 = v_40622 & v_40722;
assign v_40724 = v_40602 & v_40720;
assign v_40726 = v_40600 & v_40725;
assign v_40728 = v_40628 & v_40727;
assign v_40729 = v_40599 & v_40725;
assign v_40731 = v_40597 & v_40730;
assign v_40733 = v_40634 & v_40732;
assign v_40734 = v_40596 & v_40730;
assign v_40736 = v_40594 & v_40735;
assign v_40738 = v_40640 & v_40737;
assign v_40739 = v_40593 & v_40735;
assign v_40741 = v_40591 & v_40740;
assign v_40743 = v_40646 & v_40742;
assign v_40744 = v_40590 & v_40740;
assign v_40746 = v_40588 & v_40745;
assign v_40748 = v_40652 & v_40747;
assign v_40749 = v_40587 & v_40745;
assign v_40751 = v_40585 & v_40750;
assign v_40753 = v_40658 & v_40752;
assign v_40754 = v_40584 & v_40750;
assign v_40756 = v_40582 & v_40755;
assign v_40758 = v_40664 & v_40757;
assign v_40759 = v_40581 & v_40755;
assign v_40761 = v_40579 & v_40760;
assign v_40763 = v_40670 & v_40762;
assign v_40764 = v_40578 & v_40760;
assign v_40766 = v_40576 & v_40765;
assign v_40768 = v_40676 & v_40767;
assign v_40769 = v_40575 & v_40765;
assign v_40771 = v_40573 & v_40770;
assign v_40773 = v_40682 & v_40772;
assign v_40774 = v_40572 & v_40770;
assign v_40776 = v_40570 & v_40775;
assign v_40778 = v_40688 & v_40777;
assign v_40779 = v_40569 & v_40775;
assign v_40781 = v_40567 & v_40780;
assign v_40783 = v_40694 & v_40782;
assign v_40784 = v_40566 & v_40780;
assign v_40786 = v_40564 & v_40785;
assign v_40788 = v_40700 & v_40787;
assign v_40789 = v_40563 & v_40785;
assign v_40791 = v_40561 & v_40790;
assign v_40793 = v_40706 & v_40792;
assign v_40794 = v_40560 & v_40790;
assign v_40796 = v_40795;
assign v_40798 = v_40710 & v_40797;
assign v_40799 = v_40798;
assign v_40801 = v_40800;
assign v_40803 = ~v_3403;
assign v_40804 = ~v_37628;
assign v_40805 = v_37628;
assign v_40806 = ~v_3407;
assign v_40807 = ~v_37632;
assign v_40808 = v_37632;
assign v_40809 = ~v_3411;
assign v_40810 = ~v_37636;
assign v_40811 = v_37636;
assign v_40812 = ~v_3415;
assign v_40813 = ~v_37640;
assign v_40814 = v_37640;
assign v_40815 = ~v_37643;
assign v_40816 = ~v_3420;
assign v_40817 = v_3420;
assign v_40818 = ~v_37647;
assign v_40819 = ~v_3424;
assign v_40820 = v_3424;
assign v_40821 = ~v_37651;
assign v_40822 = ~v_3428;
assign v_40823 = v_3428;
assign v_40824 = ~v_37655;
assign v_40825 = ~v_3432;
assign v_40826 = v_3432;
assign v_40827 = ~v_37659;
assign v_40828 = ~v_3436;
assign v_40829 = v_3436;
assign v_40830 = ~v_37663;
assign v_40831 = ~v_3440;
assign v_40832 = v_3440;
assign v_40833 = ~v_37667;
assign v_40834 = ~v_3444;
assign v_40835 = v_3444;
assign v_40836 = ~v_37671;
assign v_40837 = ~v_3448;
assign v_40838 = v_3448;
assign v_40839 = ~v_37675;
assign v_40840 = ~v_3452;
assign v_40841 = v_3452;
assign v_40842 = ~v_37679;
assign v_40843 = ~v_3456;
assign v_40844 = v_3456;
assign v_40845 = ~v_37683;
assign v_40846 = ~v_3460;
assign v_40847 = v_3460;
assign v_40848 = ~v_37687;
assign v_40849 = ~v_3464;
assign v_40850 = v_3464;
assign v_40851 = ~v_37691;
assign v_40852 = ~v_3468;
assign v_40853 = v_40852;
assign v_40855 = v_40854;
assign v_40857 = v_40849 & v_40856;
assign v_40859 = v_37687;
assign v_40861 = v_40858 & v_40860;
assign v_40863 = v_40846 & v_40862;
assign v_40865 = v_37683;
assign v_40867 = v_40864 & v_40866;
assign v_40869 = v_40843 & v_40868;
assign v_40871 = v_37679;
assign v_40873 = v_40870 & v_40872;
assign v_40875 = v_40840 & v_40874;
assign v_40877 = v_37675;
assign v_40879 = v_40876 & v_40878;
assign v_40881 = v_40837 & v_40880;
assign v_40883 = v_37671;
assign v_40885 = v_40882 & v_40884;
assign v_40887 = v_40834 & v_40886;
assign v_40889 = v_37667;
assign v_40891 = v_40888 & v_40890;
assign v_40893 = v_40831 & v_40892;
assign v_40895 = v_37663;
assign v_40897 = v_40894 & v_40896;
assign v_40899 = v_40828 & v_40898;
assign v_40901 = v_37659;
assign v_40903 = v_40900 & v_40902;
assign v_40905 = v_40825 & v_40904;
assign v_40907 = v_37655;
assign v_40909 = v_40906 & v_40908;
assign v_40911 = v_40822 & v_40910;
assign v_40913 = v_37651;
assign v_40915 = v_40912 & v_40914;
assign v_40917 = v_40819 & v_40916;
assign v_40919 = v_37647;
assign v_40921 = v_40918 & v_40920;
assign v_40923 = v_40816 & v_40922;
assign v_40925 = v_37643;
assign v_40927 = v_40924 & v_40926;
assign v_40929 = v_40813 & v_40928;
assign v_40931 = v_3415;
assign v_40933 = v_40930 & v_40932;
assign v_40935 = v_40810 & v_40934;
assign v_40937 = v_3411;
assign v_40939 = v_40936 & v_40938;
assign v_40941 = v_40807 & v_40940;
assign v_40943 = v_3407;
assign v_40945 = v_40942 & v_40944;
assign v_40947 = v_40804 & v_40946;
assign v_40949 = v_3403;
assign v_40951 = v_40948 & v_40950;
assign v_40952 = v_40951;
assign v_40954 = v_37691;
assign v_40955 = v_3468;
assign v_40956 = v_40955;
assign v_40957 = v_40954 & v_40956;
assign v_40958 = v_40957;
assign v_40959 = v_40849 & v_40958;
assign v_40961 = v_40859 & v_40960;
assign v_40962 = v_40848 & v_40958;
assign v_40964 = v_40846 & v_40963;
assign v_40966 = v_40865 & v_40965;
assign v_40967 = v_40845 & v_40963;
assign v_40969 = v_40843 & v_40968;
assign v_40971 = v_40871 & v_40970;
assign v_40972 = v_40842 & v_40968;
assign v_40974 = v_40840 & v_40973;
assign v_40976 = v_40877 & v_40975;
assign v_40977 = v_40839 & v_40973;
assign v_40979 = v_40837 & v_40978;
assign v_40981 = v_40883 & v_40980;
assign v_40982 = v_40836 & v_40978;
assign v_40984 = v_40834 & v_40983;
assign v_40986 = v_40889 & v_40985;
assign v_40987 = v_40833 & v_40983;
assign v_40989 = v_40831 & v_40988;
assign v_40991 = v_40895 & v_40990;
assign v_40992 = v_40830 & v_40988;
assign v_40994 = v_40828 & v_40993;
assign v_40996 = v_40901 & v_40995;
assign v_40997 = v_40827 & v_40993;
assign v_40999 = v_40825 & v_40998;
assign v_41001 = v_40907 & v_41000;
assign v_41002 = v_40824 & v_40998;
assign v_41004 = v_40822 & v_41003;
assign v_41006 = v_40913 & v_41005;
assign v_41007 = v_40821 & v_41003;
assign v_41009 = v_40819 & v_41008;
assign v_41011 = v_40919 & v_41010;
assign v_41012 = v_40818 & v_41008;
assign v_41014 = v_40816 & v_41013;
assign v_41016 = v_40925 & v_41015;
assign v_41017 = v_40815 & v_41013;
assign v_41019 = v_40813 & v_41018;
assign v_41021 = v_40931 & v_41020;
assign v_41022 = v_40812 & v_41018;
assign v_41024 = v_40810 & v_41023;
assign v_41026 = v_40937 & v_41025;
assign v_41027 = v_40809 & v_41023;
assign v_41029 = v_40807 & v_41028;
assign v_41031 = v_40943 & v_41030;
assign v_41032 = v_40806 & v_41028;
assign v_41034 = v_40804 & v_41033;
assign v_41036 = v_40949 & v_41035;
assign v_41037 = v_40803 & v_41033;
assign v_41039 = v_41038;
assign v_41041 = v_40953 & v_41040;
assign v_41042 = v_41041;
assign v_41044 = v_41043;
assign v_41046 = ~v_3663;
assign v_41047 = ~v_37628;
assign v_41048 = v_37628;
assign v_41049 = ~v_3667;
assign v_41050 = ~v_37632;
assign v_41051 = v_37632;
assign v_41052 = ~v_3671;
assign v_41053 = ~v_37636;
assign v_41054 = v_37636;
assign v_41055 = ~v_3675;
assign v_41056 = ~v_37640;
assign v_41057 = v_37640;
assign v_41058 = ~v_37643;
assign v_41059 = ~v_3680;
assign v_41060 = v_3680;
assign v_41061 = ~v_37647;
assign v_41062 = ~v_3684;
assign v_41063 = v_3684;
assign v_41064 = ~v_37651;
assign v_41065 = ~v_3688;
assign v_41066 = v_3688;
assign v_41067 = ~v_37655;
assign v_41068 = ~v_3692;
assign v_41069 = v_3692;
assign v_41070 = ~v_37659;
assign v_41071 = ~v_3696;
assign v_41072 = v_3696;
assign v_41073 = ~v_37663;
assign v_41074 = ~v_3700;
assign v_41075 = v_3700;
assign v_41076 = ~v_37667;
assign v_41077 = ~v_3704;
assign v_41078 = v_3704;
assign v_41079 = ~v_37671;
assign v_41080 = ~v_3708;
assign v_41081 = v_3708;
assign v_41082 = ~v_37675;
assign v_41083 = ~v_3712;
assign v_41084 = v_3712;
assign v_41085 = ~v_37679;
assign v_41086 = ~v_3716;
assign v_41087 = v_3716;
assign v_41088 = ~v_37683;
assign v_41089 = ~v_3720;
assign v_41090 = v_3720;
assign v_41091 = ~v_37687;
assign v_41092 = ~v_3724;
assign v_41093 = v_3724;
assign v_41094 = ~v_37691;
assign v_41095 = ~v_3728;
assign v_41096 = v_41095;
assign v_41098 = v_41097;
assign v_41100 = v_41092 & v_41099;
assign v_41102 = v_37687;
assign v_41104 = v_41101 & v_41103;
assign v_41106 = v_41089 & v_41105;
assign v_41108 = v_37683;
assign v_41110 = v_41107 & v_41109;
assign v_41112 = v_41086 & v_41111;
assign v_41114 = v_37679;
assign v_41116 = v_41113 & v_41115;
assign v_41118 = v_41083 & v_41117;
assign v_41120 = v_37675;
assign v_41122 = v_41119 & v_41121;
assign v_41124 = v_41080 & v_41123;
assign v_41126 = v_37671;
assign v_41128 = v_41125 & v_41127;
assign v_41130 = v_41077 & v_41129;
assign v_41132 = v_37667;
assign v_41134 = v_41131 & v_41133;
assign v_41136 = v_41074 & v_41135;
assign v_41138 = v_37663;
assign v_41140 = v_41137 & v_41139;
assign v_41142 = v_41071 & v_41141;
assign v_41144 = v_37659;
assign v_41146 = v_41143 & v_41145;
assign v_41148 = v_41068 & v_41147;
assign v_41150 = v_37655;
assign v_41152 = v_41149 & v_41151;
assign v_41154 = v_41065 & v_41153;
assign v_41156 = v_37651;
assign v_41158 = v_41155 & v_41157;
assign v_41160 = v_41062 & v_41159;
assign v_41162 = v_37647;
assign v_41164 = v_41161 & v_41163;
assign v_41166 = v_41059 & v_41165;
assign v_41168 = v_37643;
assign v_41170 = v_41167 & v_41169;
assign v_41172 = v_41056 & v_41171;
assign v_41174 = v_3675;
assign v_41176 = v_41173 & v_41175;
assign v_41178 = v_41053 & v_41177;
assign v_41180 = v_3671;
assign v_41182 = v_41179 & v_41181;
assign v_41184 = v_41050 & v_41183;
assign v_41186 = v_3667;
assign v_41188 = v_41185 & v_41187;
assign v_41190 = v_41047 & v_41189;
assign v_41192 = v_3663;
assign v_41194 = v_41191 & v_41193;
assign v_41195 = v_41194;
assign v_41197 = v_37691;
assign v_41198 = v_3728;
assign v_41199 = v_41198;
assign v_41200 = v_41197 & v_41199;
assign v_41201 = v_41200;
assign v_41202 = v_41092 & v_41201;
assign v_41204 = v_41102 & v_41203;
assign v_41205 = v_41091 & v_41201;
assign v_41207 = v_41089 & v_41206;
assign v_41209 = v_41108 & v_41208;
assign v_41210 = v_41088 & v_41206;
assign v_41212 = v_41086 & v_41211;
assign v_41214 = v_41114 & v_41213;
assign v_41215 = v_41085 & v_41211;
assign v_41217 = v_41083 & v_41216;
assign v_41219 = v_41120 & v_41218;
assign v_41220 = v_41082 & v_41216;
assign v_41222 = v_41080 & v_41221;
assign v_41224 = v_41126 & v_41223;
assign v_41225 = v_41079 & v_41221;
assign v_41227 = v_41077 & v_41226;
assign v_41229 = v_41132 & v_41228;
assign v_41230 = v_41076 & v_41226;
assign v_41232 = v_41074 & v_41231;
assign v_41234 = v_41138 & v_41233;
assign v_41235 = v_41073 & v_41231;
assign v_41237 = v_41071 & v_41236;
assign v_41239 = v_41144 & v_41238;
assign v_41240 = v_41070 & v_41236;
assign v_41242 = v_41068 & v_41241;
assign v_41244 = v_41150 & v_41243;
assign v_41245 = v_41067 & v_41241;
assign v_41247 = v_41065 & v_41246;
assign v_41249 = v_41156 & v_41248;
assign v_41250 = v_41064 & v_41246;
assign v_41252 = v_41062 & v_41251;
assign v_41254 = v_41162 & v_41253;
assign v_41255 = v_41061 & v_41251;
assign v_41257 = v_41059 & v_41256;
assign v_41259 = v_41168 & v_41258;
assign v_41260 = v_41058 & v_41256;
assign v_41262 = v_41056 & v_41261;
assign v_41264 = v_41174 & v_41263;
assign v_41265 = v_41055 & v_41261;
assign v_41267 = v_41053 & v_41266;
assign v_41269 = v_41180 & v_41268;
assign v_41270 = v_41052 & v_41266;
assign v_41272 = v_41050 & v_41271;
assign v_41274 = v_41186 & v_41273;
assign v_41275 = v_41049 & v_41271;
assign v_41277 = v_41047 & v_41276;
assign v_41279 = v_41192 & v_41278;
assign v_41280 = v_41046 & v_41276;
assign v_41282 = v_41281;
assign v_41284 = v_41196 & v_41283;
assign v_41285 = v_41284;
assign v_41287 = v_41286;
assign v_41289 = ~v_3923;
assign v_41290 = ~v_37628;
assign v_41291 = v_37628;
assign v_41292 = ~v_3927;
assign v_41293 = ~v_37632;
assign v_41294 = v_37632;
assign v_41295 = ~v_3931;
assign v_41296 = ~v_37636;
assign v_41297 = v_37636;
assign v_41298 = ~v_3935;
assign v_41299 = ~v_37640;
assign v_41300 = v_37640;
assign v_41301 = ~v_37643;
assign v_41302 = ~v_3940;
assign v_41303 = v_3940;
assign v_41304 = ~v_37647;
assign v_41305 = ~v_3944;
assign v_41306 = v_3944;
assign v_41307 = ~v_37651;
assign v_41308 = ~v_3948;
assign v_41309 = v_3948;
assign v_41310 = ~v_37655;
assign v_41311 = ~v_3952;
assign v_41312 = v_3952;
assign v_41313 = ~v_37659;
assign v_41314 = ~v_3956;
assign v_41315 = v_3956;
assign v_41316 = ~v_37663;
assign v_41317 = ~v_3960;
assign v_41318 = v_3960;
assign v_41319 = ~v_37667;
assign v_41320 = ~v_3964;
assign v_41321 = v_3964;
assign v_41322 = ~v_37671;
assign v_41323 = ~v_3968;
assign v_41324 = v_3968;
assign v_41325 = ~v_37675;
assign v_41326 = ~v_3972;
assign v_41327 = v_3972;
assign v_41328 = ~v_37679;
assign v_41329 = ~v_3976;
assign v_41330 = v_3976;
assign v_41331 = ~v_37683;
assign v_41332 = ~v_3980;
assign v_41333 = v_3980;
assign v_41334 = ~v_37687;
assign v_41335 = ~v_3984;
assign v_41336 = v_3984;
assign v_41337 = ~v_37691;
assign v_41338 = ~v_3988;
assign v_41339 = v_41338;
assign v_41341 = v_41340;
assign v_41343 = v_41335 & v_41342;
assign v_41345 = v_37687;
assign v_41347 = v_41344 & v_41346;
assign v_41349 = v_41332 & v_41348;
assign v_41351 = v_37683;
assign v_41353 = v_41350 & v_41352;
assign v_41355 = v_41329 & v_41354;
assign v_41357 = v_37679;
assign v_41359 = v_41356 & v_41358;
assign v_41361 = v_41326 & v_41360;
assign v_41363 = v_37675;
assign v_41365 = v_41362 & v_41364;
assign v_41367 = v_41323 & v_41366;
assign v_41369 = v_37671;
assign v_41371 = v_41368 & v_41370;
assign v_41373 = v_41320 & v_41372;
assign v_41375 = v_37667;
assign v_41377 = v_41374 & v_41376;
assign v_41379 = v_41317 & v_41378;
assign v_41381 = v_37663;
assign v_41383 = v_41380 & v_41382;
assign v_41385 = v_41314 & v_41384;
assign v_41387 = v_37659;
assign v_41389 = v_41386 & v_41388;
assign v_41391 = v_41311 & v_41390;
assign v_41393 = v_37655;
assign v_41395 = v_41392 & v_41394;
assign v_41397 = v_41308 & v_41396;
assign v_41399 = v_37651;
assign v_41401 = v_41398 & v_41400;
assign v_41403 = v_41305 & v_41402;
assign v_41405 = v_37647;
assign v_41407 = v_41404 & v_41406;
assign v_41409 = v_41302 & v_41408;
assign v_41411 = v_37643;
assign v_41413 = v_41410 & v_41412;
assign v_41415 = v_41299 & v_41414;
assign v_41417 = v_3935;
assign v_41419 = v_41416 & v_41418;
assign v_41421 = v_41296 & v_41420;
assign v_41423 = v_3931;
assign v_41425 = v_41422 & v_41424;
assign v_41427 = v_41293 & v_41426;
assign v_41429 = v_3927;
assign v_41431 = v_41428 & v_41430;
assign v_41433 = v_41290 & v_41432;
assign v_41435 = v_3923;
assign v_41437 = v_41434 & v_41436;
assign v_41438 = v_41437;
assign v_41440 = v_37691;
assign v_41441 = v_3988;
assign v_41442 = v_41441;
assign v_41443 = v_41440 & v_41442;
assign v_41444 = v_41443;
assign v_41445 = v_41335 & v_41444;
assign v_41447 = v_41345 & v_41446;
assign v_41448 = v_41334 & v_41444;
assign v_41450 = v_41332 & v_41449;
assign v_41452 = v_41351 & v_41451;
assign v_41453 = v_41331 & v_41449;
assign v_41455 = v_41329 & v_41454;
assign v_41457 = v_41357 & v_41456;
assign v_41458 = v_41328 & v_41454;
assign v_41460 = v_41326 & v_41459;
assign v_41462 = v_41363 & v_41461;
assign v_41463 = v_41325 & v_41459;
assign v_41465 = v_41323 & v_41464;
assign v_41467 = v_41369 & v_41466;
assign v_41468 = v_41322 & v_41464;
assign v_41470 = v_41320 & v_41469;
assign v_41472 = v_41375 & v_41471;
assign v_41473 = v_41319 & v_41469;
assign v_41475 = v_41317 & v_41474;
assign v_41477 = v_41381 & v_41476;
assign v_41478 = v_41316 & v_41474;
assign v_41480 = v_41314 & v_41479;
assign v_41482 = v_41387 & v_41481;
assign v_41483 = v_41313 & v_41479;
assign v_41485 = v_41311 & v_41484;
assign v_41487 = v_41393 & v_41486;
assign v_41488 = v_41310 & v_41484;
assign v_41490 = v_41308 & v_41489;
assign v_41492 = v_41399 & v_41491;
assign v_41493 = v_41307 & v_41489;
assign v_41495 = v_41305 & v_41494;
assign v_41497 = v_41405 & v_41496;
assign v_41498 = v_41304 & v_41494;
assign v_41500 = v_41302 & v_41499;
assign v_41502 = v_41411 & v_41501;
assign v_41503 = v_41301 & v_41499;
assign v_41505 = v_41299 & v_41504;
assign v_41507 = v_41417 & v_41506;
assign v_41508 = v_41298 & v_41504;
assign v_41510 = v_41296 & v_41509;
assign v_41512 = v_41423 & v_41511;
assign v_41513 = v_41295 & v_41509;
assign v_41515 = v_41293 & v_41514;
assign v_41517 = v_41429 & v_41516;
assign v_41518 = v_41292 & v_41514;
assign v_41520 = v_41290 & v_41519;
assign v_41522 = v_41435 & v_41521;
assign v_41523 = v_41289 & v_41519;
assign v_41525 = v_41524;
assign v_41527 = v_41439 & v_41526;
assign v_41528 = v_41527;
assign v_41530 = v_41529;
assign v_41531 = ~v_4182;
assign v_41532 = ~v_37628;
assign v_41533 = v_37628;
assign v_41534 = ~v_4186;
assign v_41535 = ~v_37632;
assign v_41536 = v_37632;
assign v_41537 = ~v_4190;
assign v_41538 = ~v_37636;
assign v_41539 = v_37636;
assign v_41540 = ~v_4194;
assign v_41541 = ~v_37640;
assign v_41542 = v_37640;
assign v_41543 = ~v_37643;
assign v_41544 = ~v_4199;
assign v_41545 = v_4199;
assign v_41546 = ~v_37647;
assign v_41547 = ~v_4203;
assign v_41548 = v_4203;
assign v_41549 = ~v_37651;
assign v_41550 = ~v_4207;
assign v_41551 = v_4207;
assign v_41552 = ~v_37655;
assign v_41553 = ~v_4211;
assign v_41554 = v_4211;
assign v_41555 = ~v_37659;
assign v_41556 = ~v_4215;
assign v_41557 = v_4215;
assign v_41558 = ~v_37663;
assign v_41559 = ~v_4219;
assign v_41560 = v_4219;
assign v_41561 = ~v_37667;
assign v_41562 = ~v_4223;
assign v_41563 = v_4223;
assign v_41564 = ~v_37671;
assign v_41565 = ~v_4227;
assign v_41566 = v_4227;
assign v_41567 = ~v_37675;
assign v_41568 = ~v_4231;
assign v_41569 = v_4231;
assign v_41570 = ~v_37679;
assign v_41571 = ~v_4235;
assign v_41572 = v_4235;
assign v_41573 = ~v_37683;
assign v_41574 = ~v_4239;
assign v_41575 = v_4239;
assign v_41576 = ~v_37687;
assign v_41577 = ~v_4243;
assign v_41578 = v_4243;
assign v_41579 = ~v_37691;
assign v_41580 = ~v_4247;
assign v_41581 = v_41580;
assign v_41583 = v_41582;
assign v_41585 = v_41577 & v_41584;
assign v_41587 = v_37687;
assign v_41589 = v_41586 & v_41588;
assign v_41591 = v_41574 & v_41590;
assign v_41593 = v_37683;
assign v_41595 = v_41592 & v_41594;
assign v_41597 = v_41571 & v_41596;
assign v_41599 = v_37679;
assign v_41601 = v_41598 & v_41600;
assign v_41603 = v_41568 & v_41602;
assign v_41605 = v_37675;
assign v_41607 = v_41604 & v_41606;
assign v_41609 = v_41565 & v_41608;
assign v_41611 = v_37671;
assign v_41613 = v_41610 & v_41612;
assign v_41615 = v_41562 & v_41614;
assign v_41617 = v_37667;
assign v_41619 = v_41616 & v_41618;
assign v_41621 = v_41559 & v_41620;
assign v_41623 = v_37663;
assign v_41625 = v_41622 & v_41624;
assign v_41627 = v_41556 & v_41626;
assign v_41629 = v_37659;
assign v_41631 = v_41628 & v_41630;
assign v_41633 = v_41553 & v_41632;
assign v_41635 = v_37655;
assign v_41637 = v_41634 & v_41636;
assign v_41639 = v_41550 & v_41638;
assign v_41641 = v_37651;
assign v_41643 = v_41640 & v_41642;
assign v_41645 = v_41547 & v_41644;
assign v_41647 = v_37647;
assign v_41649 = v_41646 & v_41648;
assign v_41651 = v_41544 & v_41650;
assign v_41653 = v_37643;
assign v_41655 = v_41652 & v_41654;
assign v_41657 = v_41541 & v_41656;
assign v_41659 = v_4194;
assign v_41661 = v_41658 & v_41660;
assign v_41663 = v_41538 & v_41662;
assign v_41665 = v_4190;
assign v_41667 = v_41664 & v_41666;
assign v_41669 = v_41535 & v_41668;
assign v_41671 = v_4186;
assign v_41673 = v_41670 & v_41672;
assign v_41675 = v_41532 & v_41674;
assign v_41677 = v_4182;
assign v_41679 = v_41676 & v_41678;
assign v_41681 = ~v_41680;
assign v_41683 = v_37691;
assign v_41684 = v_4247;
assign v_41685 = v_41684;
assign v_41686 = v_41683 & v_41685;
assign v_41687 = v_41686;
assign v_41688 = v_41577 & v_41687;
assign v_41690 = v_41587 & v_41689;
assign v_41691 = v_41576 & v_41687;
assign v_41693 = v_41574 & v_41692;
assign v_41695 = v_41593 & v_41694;
assign v_41696 = v_41573 & v_41692;
assign v_41698 = v_41571 & v_41697;
assign v_41700 = v_41599 & v_41699;
assign v_41701 = v_41570 & v_41697;
assign v_41703 = v_41568 & v_41702;
assign v_41705 = v_41605 & v_41704;
assign v_41706 = v_41567 & v_41702;
assign v_41708 = v_41565 & v_41707;
assign v_41710 = v_41611 & v_41709;
assign v_41711 = v_41564 & v_41707;
assign v_41713 = v_41562 & v_41712;
assign v_41715 = v_41617 & v_41714;
assign v_41716 = v_41561 & v_41712;
assign v_41718 = v_41559 & v_41717;
assign v_41720 = v_41623 & v_41719;
assign v_41721 = v_41558 & v_41717;
assign v_41723 = v_41556 & v_41722;
assign v_41725 = v_41629 & v_41724;
assign v_41726 = v_41555 & v_41722;
assign v_41728 = v_41553 & v_41727;
assign v_41730 = v_41635 & v_41729;
assign v_41731 = v_41552 & v_41727;
assign v_41733 = v_41550 & v_41732;
assign v_41735 = v_41641 & v_41734;
assign v_41736 = v_41549 & v_41732;
assign v_41738 = v_41547 & v_41737;
assign v_41740 = v_41647 & v_41739;
assign v_41741 = v_41546 & v_41737;
assign v_41743 = v_41544 & v_41742;
assign v_41745 = v_41653 & v_41744;
assign v_41746 = v_41543 & v_41742;
assign v_41748 = v_41541 & v_41747;
assign v_41750 = v_41659 & v_41749;
assign v_41751 = v_41540 & v_41747;
assign v_41753 = v_41538 & v_41752;
assign v_41755 = v_41665 & v_41754;
assign v_41756 = v_41537 & v_41752;
assign v_41758 = v_41535 & v_41757;
assign v_41760 = v_41671 & v_41759;
assign v_41761 = v_41534 & v_41757;
assign v_41763 = v_41532 & v_41762;
assign v_41765 = v_41677 & v_41764;
assign v_41766 = v_41531 & v_41762;
assign v_41768 = v_41680;
assign v_41770 = v_41682 & v_41769;
assign v_41771 = v_41770;
assign v_41773 = v_41772;
assign v_41775 = ~v_6;
assign v_41777 = ~v_41776;
assign v_41778 = v_41776;
assign v_41779 = ~v_13;
assign v_41781 = ~v_41780;
assign v_41782 = v_41780;
assign v_41783 = ~v_18;
assign v_41785 = ~v_41784;
assign v_41786 = v_41784;
assign v_41787 = ~v_23;
assign v_41789 = ~v_41788;
assign v_41790 = v_41788;
assign v_41792 = ~v_41791;
assign v_41793 = ~v_30;
assign v_41794 = v_30;
assign v_41796 = ~v_41795;
assign v_41797 = ~v_35;
assign v_41798 = v_35;
assign v_41800 = ~v_41799;
assign v_41801 = ~v_40;
assign v_41802 = v_40;
assign v_41804 = ~v_41803;
assign v_41805 = ~v_45;
assign v_41806 = v_45;
assign v_41808 = ~v_41807;
assign v_41809 = ~v_50;
assign v_41810 = v_50;
assign v_41812 = ~v_41811;
assign v_41813 = ~v_55;
assign v_41814 = v_55;
assign v_41816 = ~v_41815;
assign v_41817 = ~v_60;
assign v_41818 = v_60;
assign v_41820 = ~v_41819;
assign v_41821 = ~v_65;
assign v_41822 = v_65;
assign v_41824 = ~v_41823;
assign v_41825 = ~v_70;
assign v_41826 = v_70;
assign v_41828 = ~v_41827;
assign v_41829 = ~v_75;
assign v_41830 = v_75;
assign v_41832 = ~v_41831;
assign v_41833 = ~v_80;
assign v_41834 = v_80;
assign v_41836 = ~v_41835;
assign v_41837 = ~v_85;
assign v_41838 = v_85;
assign v_41840 = ~v_41839;
assign v_41841 = ~v_90;
assign v_41842 = v_41841;
assign v_41844 = v_41843;
assign v_41846 = v_41837 & v_41845;
assign v_41848 = v_41835;
assign v_41850 = v_41847 & v_41849;
assign v_41852 = v_41833 & v_41851;
assign v_41854 = v_41831;
assign v_41856 = v_41853 & v_41855;
assign v_41858 = v_41829 & v_41857;
assign v_41860 = v_41827;
assign v_41862 = v_41859 & v_41861;
assign v_41864 = v_41825 & v_41863;
assign v_41866 = v_41823;
assign v_41868 = v_41865 & v_41867;
assign v_41870 = v_41821 & v_41869;
assign v_41872 = v_41819;
assign v_41874 = v_41871 & v_41873;
assign v_41876 = v_41817 & v_41875;
assign v_41878 = v_41815;
assign v_41880 = v_41877 & v_41879;
assign v_41882 = v_41813 & v_41881;
assign v_41884 = v_41811;
assign v_41886 = v_41883 & v_41885;
assign v_41888 = v_41809 & v_41887;
assign v_41890 = v_41807;
assign v_41892 = v_41889 & v_41891;
assign v_41894 = v_41805 & v_41893;
assign v_41896 = v_41803;
assign v_41898 = v_41895 & v_41897;
assign v_41900 = v_41801 & v_41899;
assign v_41902 = v_41799;
assign v_41904 = v_41901 & v_41903;
assign v_41906 = v_41797 & v_41905;
assign v_41908 = v_41795;
assign v_41910 = v_41907 & v_41909;
assign v_41912 = v_41793 & v_41911;
assign v_41914 = v_41791;
assign v_41916 = v_41913 & v_41915;
assign v_41918 = v_41789 & v_41917;
assign v_41920 = v_23;
assign v_41922 = v_41919 & v_41921;
assign v_41924 = v_41785 & v_41923;
assign v_41926 = v_18;
assign v_41928 = v_41925 & v_41927;
assign v_41930 = v_41781 & v_41929;
assign v_41932 = v_13;
assign v_41934 = v_41931 & v_41933;
assign v_41936 = v_41777 & v_41935;
assign v_41938 = v_6;
assign v_41940 = v_41937 & v_41939;
assign v_41941 = v_41940;
assign v_41943 = v_41839;
assign v_41944 = v_90;
assign v_41945 = v_41944;
assign v_41946 = v_41943 & v_41945;
assign v_41947 = v_41946;
assign v_41948 = v_41837 & v_41947;
assign v_41950 = v_41848 & v_41949;
assign v_41951 = v_41836 & v_41947;
assign v_41953 = v_41833 & v_41952;
assign v_41955 = v_41854 & v_41954;
assign v_41956 = v_41832 & v_41952;
assign v_41958 = v_41829 & v_41957;
assign v_41960 = v_41860 & v_41959;
assign v_41961 = v_41828 & v_41957;
assign v_41963 = v_41825 & v_41962;
assign v_41965 = v_41866 & v_41964;
assign v_41966 = v_41824 & v_41962;
assign v_41968 = v_41821 & v_41967;
assign v_41970 = v_41872 & v_41969;
assign v_41971 = v_41820 & v_41967;
assign v_41973 = v_41817 & v_41972;
assign v_41975 = v_41878 & v_41974;
assign v_41976 = v_41816 & v_41972;
assign v_41978 = v_41813 & v_41977;
assign v_41980 = v_41884 & v_41979;
assign v_41981 = v_41812 & v_41977;
assign v_41983 = v_41809 & v_41982;
assign v_41985 = v_41890 & v_41984;
assign v_41986 = v_41808 & v_41982;
assign v_41988 = v_41805 & v_41987;
assign v_41990 = v_41896 & v_41989;
assign v_41991 = v_41804 & v_41987;
assign v_41993 = v_41801 & v_41992;
assign v_41995 = v_41902 & v_41994;
assign v_41996 = v_41800 & v_41992;
assign v_41998 = v_41797 & v_41997;
assign v_42000 = v_41908 & v_41999;
assign v_42001 = v_41796 & v_41997;
assign v_42003 = v_41793 & v_42002;
assign v_42005 = v_41914 & v_42004;
assign v_42006 = v_41792 & v_42002;
assign v_42008 = v_41789 & v_42007;
assign v_42010 = v_41920 & v_42009;
assign v_42011 = v_41787 & v_42007;
assign v_42013 = v_41785 & v_42012;
assign v_42015 = v_41926 & v_42014;
assign v_42016 = v_41783 & v_42012;
assign v_42018 = v_41781 & v_42017;
assign v_42020 = v_41932 & v_42019;
assign v_42021 = v_41779 & v_42017;
assign v_42023 = v_41777 & v_42022;
assign v_42025 = v_41938 & v_42024;
assign v_42026 = v_41775 & v_42022;
assign v_42028 = v_42027;
assign v_42030 = v_41942 & v_42029;
assign v_42031 = v_42030;
assign v_42033 = v_42032;
assign v_42035 = ~v_283;
assign v_42036 = ~v_41776;
assign v_42037 = v_41776;
assign v_42038 = ~v_287;
assign v_42039 = ~v_41780;
assign v_42040 = v_41780;
assign v_42041 = ~v_291;
assign v_42042 = ~v_41784;
assign v_42043 = v_41784;
assign v_42044 = ~v_295;
assign v_42045 = ~v_41788;
assign v_42046 = v_41788;
assign v_42047 = ~v_41791;
assign v_42048 = ~v_300;
assign v_42049 = v_300;
assign v_42050 = ~v_41795;
assign v_42051 = ~v_304;
assign v_42052 = v_304;
assign v_42053 = ~v_41799;
assign v_42054 = ~v_308;
assign v_42055 = v_308;
assign v_42056 = ~v_41803;
assign v_42057 = ~v_312;
assign v_42058 = v_312;
assign v_42059 = ~v_41807;
assign v_42060 = ~v_316;
assign v_42061 = v_316;
assign v_42062 = ~v_41811;
assign v_42063 = ~v_320;
assign v_42064 = v_320;
assign v_42065 = ~v_41815;
assign v_42066 = ~v_324;
assign v_42067 = v_324;
assign v_42068 = ~v_41819;
assign v_42069 = ~v_328;
assign v_42070 = v_328;
assign v_42071 = ~v_41823;
assign v_42072 = ~v_332;
assign v_42073 = v_332;
assign v_42074 = ~v_41827;
assign v_42075 = ~v_336;
assign v_42076 = v_336;
assign v_42077 = ~v_41831;
assign v_42078 = ~v_340;
assign v_42079 = v_340;
assign v_42080 = ~v_41835;
assign v_42081 = ~v_344;
assign v_42082 = v_344;
assign v_42083 = ~v_41839;
assign v_42084 = ~v_348;
assign v_42085 = v_42084;
assign v_42087 = v_42086;
assign v_42089 = v_42081 & v_42088;
assign v_42091 = v_41835;
assign v_42093 = v_42090 & v_42092;
assign v_42095 = v_42078 & v_42094;
assign v_42097 = v_41831;
assign v_42099 = v_42096 & v_42098;
assign v_42101 = v_42075 & v_42100;
assign v_42103 = v_41827;
assign v_42105 = v_42102 & v_42104;
assign v_42107 = v_42072 & v_42106;
assign v_42109 = v_41823;
assign v_42111 = v_42108 & v_42110;
assign v_42113 = v_42069 & v_42112;
assign v_42115 = v_41819;
assign v_42117 = v_42114 & v_42116;
assign v_42119 = v_42066 & v_42118;
assign v_42121 = v_41815;
assign v_42123 = v_42120 & v_42122;
assign v_42125 = v_42063 & v_42124;
assign v_42127 = v_41811;
assign v_42129 = v_42126 & v_42128;
assign v_42131 = v_42060 & v_42130;
assign v_42133 = v_41807;
assign v_42135 = v_42132 & v_42134;
assign v_42137 = v_42057 & v_42136;
assign v_42139 = v_41803;
assign v_42141 = v_42138 & v_42140;
assign v_42143 = v_42054 & v_42142;
assign v_42145 = v_41799;
assign v_42147 = v_42144 & v_42146;
assign v_42149 = v_42051 & v_42148;
assign v_42151 = v_41795;
assign v_42153 = v_42150 & v_42152;
assign v_42155 = v_42048 & v_42154;
assign v_42157 = v_41791;
assign v_42159 = v_42156 & v_42158;
assign v_42161 = v_42045 & v_42160;
assign v_42163 = v_295;
assign v_42165 = v_42162 & v_42164;
assign v_42167 = v_42042 & v_42166;
assign v_42169 = v_291;
assign v_42171 = v_42168 & v_42170;
assign v_42173 = v_42039 & v_42172;
assign v_42175 = v_287;
assign v_42177 = v_42174 & v_42176;
assign v_42179 = v_42036 & v_42178;
assign v_42181 = v_283;
assign v_42183 = v_42180 & v_42182;
assign v_42184 = v_42183;
assign v_42186 = v_41839;
assign v_42187 = v_348;
assign v_42188 = v_42187;
assign v_42189 = v_42186 & v_42188;
assign v_42190 = v_42189;
assign v_42191 = v_42081 & v_42190;
assign v_42193 = v_42091 & v_42192;
assign v_42194 = v_42080 & v_42190;
assign v_42196 = v_42078 & v_42195;
assign v_42198 = v_42097 & v_42197;
assign v_42199 = v_42077 & v_42195;
assign v_42201 = v_42075 & v_42200;
assign v_42203 = v_42103 & v_42202;
assign v_42204 = v_42074 & v_42200;
assign v_42206 = v_42072 & v_42205;
assign v_42208 = v_42109 & v_42207;
assign v_42209 = v_42071 & v_42205;
assign v_42211 = v_42069 & v_42210;
assign v_42213 = v_42115 & v_42212;
assign v_42214 = v_42068 & v_42210;
assign v_42216 = v_42066 & v_42215;
assign v_42218 = v_42121 & v_42217;
assign v_42219 = v_42065 & v_42215;
assign v_42221 = v_42063 & v_42220;
assign v_42223 = v_42127 & v_42222;
assign v_42224 = v_42062 & v_42220;
assign v_42226 = v_42060 & v_42225;
assign v_42228 = v_42133 & v_42227;
assign v_42229 = v_42059 & v_42225;
assign v_42231 = v_42057 & v_42230;
assign v_42233 = v_42139 & v_42232;
assign v_42234 = v_42056 & v_42230;
assign v_42236 = v_42054 & v_42235;
assign v_42238 = v_42145 & v_42237;
assign v_42239 = v_42053 & v_42235;
assign v_42241 = v_42051 & v_42240;
assign v_42243 = v_42151 & v_42242;
assign v_42244 = v_42050 & v_42240;
assign v_42246 = v_42048 & v_42245;
assign v_42248 = v_42157 & v_42247;
assign v_42249 = v_42047 & v_42245;
assign v_42251 = v_42045 & v_42250;
assign v_42253 = v_42163 & v_42252;
assign v_42254 = v_42044 & v_42250;
assign v_42256 = v_42042 & v_42255;
assign v_42258 = v_42169 & v_42257;
assign v_42259 = v_42041 & v_42255;
assign v_42261 = v_42039 & v_42260;
assign v_42263 = v_42175 & v_42262;
assign v_42264 = v_42038 & v_42260;
assign v_42266 = v_42036 & v_42265;
assign v_42268 = v_42181 & v_42267;
assign v_42269 = v_42035 & v_42265;
assign v_42271 = v_42270;
assign v_42273 = v_42185 & v_42272;
assign v_42274 = v_42273;
assign v_42276 = v_42275;
assign v_42278 = ~v_543;
assign v_42279 = ~v_41776;
assign v_42280 = v_41776;
assign v_42281 = ~v_547;
assign v_42282 = ~v_41780;
assign v_42283 = v_41780;
assign v_42284 = ~v_551;
assign v_42285 = ~v_41784;
assign v_42286 = v_41784;
assign v_42287 = ~v_555;
assign v_42288 = ~v_41788;
assign v_42289 = v_41788;
assign v_42290 = ~v_41791;
assign v_42291 = ~v_560;
assign v_42292 = v_560;
assign v_42293 = ~v_41795;
assign v_42294 = ~v_564;
assign v_42295 = v_564;
assign v_42296 = ~v_41799;
assign v_42297 = ~v_568;
assign v_42298 = v_568;
assign v_42299 = ~v_41803;
assign v_42300 = ~v_572;
assign v_42301 = v_572;
assign v_42302 = ~v_41807;
assign v_42303 = ~v_576;
assign v_42304 = v_576;
assign v_42305 = ~v_41811;
assign v_42306 = ~v_580;
assign v_42307 = v_580;
assign v_42308 = ~v_41815;
assign v_42309 = ~v_584;
assign v_42310 = v_584;
assign v_42311 = ~v_41819;
assign v_42312 = ~v_588;
assign v_42313 = v_588;
assign v_42314 = ~v_41823;
assign v_42315 = ~v_592;
assign v_42316 = v_592;
assign v_42317 = ~v_41827;
assign v_42318 = ~v_596;
assign v_42319 = v_596;
assign v_42320 = ~v_41831;
assign v_42321 = ~v_600;
assign v_42322 = v_600;
assign v_42323 = ~v_41835;
assign v_42324 = ~v_604;
assign v_42325 = v_604;
assign v_42326 = ~v_41839;
assign v_42327 = ~v_608;
assign v_42328 = v_42327;
assign v_42330 = v_42329;
assign v_42332 = v_42324 & v_42331;
assign v_42334 = v_41835;
assign v_42336 = v_42333 & v_42335;
assign v_42338 = v_42321 & v_42337;
assign v_42340 = v_41831;
assign v_42342 = v_42339 & v_42341;
assign v_42344 = v_42318 & v_42343;
assign v_42346 = v_41827;
assign v_42348 = v_42345 & v_42347;
assign v_42350 = v_42315 & v_42349;
assign v_42352 = v_41823;
assign v_42354 = v_42351 & v_42353;
assign v_42356 = v_42312 & v_42355;
assign v_42358 = v_41819;
assign v_42360 = v_42357 & v_42359;
assign v_42362 = v_42309 & v_42361;
assign v_42364 = v_41815;
assign v_42366 = v_42363 & v_42365;
assign v_42368 = v_42306 & v_42367;
assign v_42370 = v_41811;
assign v_42372 = v_42369 & v_42371;
assign v_42374 = v_42303 & v_42373;
assign v_42376 = v_41807;
assign v_42378 = v_42375 & v_42377;
assign v_42380 = v_42300 & v_42379;
assign v_42382 = v_41803;
assign v_42384 = v_42381 & v_42383;
assign v_42386 = v_42297 & v_42385;
assign v_42388 = v_41799;
assign v_42390 = v_42387 & v_42389;
assign v_42392 = v_42294 & v_42391;
assign v_42394 = v_41795;
assign v_42396 = v_42393 & v_42395;
assign v_42398 = v_42291 & v_42397;
assign v_42400 = v_41791;
assign v_42402 = v_42399 & v_42401;
assign v_42404 = v_42288 & v_42403;
assign v_42406 = v_555;
assign v_42408 = v_42405 & v_42407;
assign v_42410 = v_42285 & v_42409;
assign v_42412 = v_551;
assign v_42414 = v_42411 & v_42413;
assign v_42416 = v_42282 & v_42415;
assign v_42418 = v_547;
assign v_42420 = v_42417 & v_42419;
assign v_42422 = v_42279 & v_42421;
assign v_42424 = v_543;
assign v_42426 = v_42423 & v_42425;
assign v_42427 = v_42426;
assign v_42429 = v_41839;
assign v_42430 = v_608;
assign v_42431 = v_42430;
assign v_42432 = v_42429 & v_42431;
assign v_42433 = v_42432;
assign v_42434 = v_42324 & v_42433;
assign v_42436 = v_42334 & v_42435;
assign v_42437 = v_42323 & v_42433;
assign v_42439 = v_42321 & v_42438;
assign v_42441 = v_42340 & v_42440;
assign v_42442 = v_42320 & v_42438;
assign v_42444 = v_42318 & v_42443;
assign v_42446 = v_42346 & v_42445;
assign v_42447 = v_42317 & v_42443;
assign v_42449 = v_42315 & v_42448;
assign v_42451 = v_42352 & v_42450;
assign v_42452 = v_42314 & v_42448;
assign v_42454 = v_42312 & v_42453;
assign v_42456 = v_42358 & v_42455;
assign v_42457 = v_42311 & v_42453;
assign v_42459 = v_42309 & v_42458;
assign v_42461 = v_42364 & v_42460;
assign v_42462 = v_42308 & v_42458;
assign v_42464 = v_42306 & v_42463;
assign v_42466 = v_42370 & v_42465;
assign v_42467 = v_42305 & v_42463;
assign v_42469 = v_42303 & v_42468;
assign v_42471 = v_42376 & v_42470;
assign v_42472 = v_42302 & v_42468;
assign v_42474 = v_42300 & v_42473;
assign v_42476 = v_42382 & v_42475;
assign v_42477 = v_42299 & v_42473;
assign v_42479 = v_42297 & v_42478;
assign v_42481 = v_42388 & v_42480;
assign v_42482 = v_42296 & v_42478;
assign v_42484 = v_42294 & v_42483;
assign v_42486 = v_42394 & v_42485;
assign v_42487 = v_42293 & v_42483;
assign v_42489 = v_42291 & v_42488;
assign v_42491 = v_42400 & v_42490;
assign v_42492 = v_42290 & v_42488;
assign v_42494 = v_42288 & v_42493;
assign v_42496 = v_42406 & v_42495;
assign v_42497 = v_42287 & v_42493;
assign v_42499 = v_42285 & v_42498;
assign v_42501 = v_42412 & v_42500;
assign v_42502 = v_42284 & v_42498;
assign v_42504 = v_42282 & v_42503;
assign v_42506 = v_42418 & v_42505;
assign v_42507 = v_42281 & v_42503;
assign v_42509 = v_42279 & v_42508;
assign v_42511 = v_42424 & v_42510;
assign v_42512 = v_42278 & v_42508;
assign v_42514 = v_42513;
assign v_42516 = v_42428 & v_42515;
assign v_42517 = v_42516;
assign v_42519 = v_42518;
assign v_42521 = ~v_803;
assign v_42522 = ~v_41776;
assign v_42523 = v_41776;
assign v_42524 = ~v_807;
assign v_42525 = ~v_41780;
assign v_42526 = v_41780;
assign v_42527 = ~v_811;
assign v_42528 = ~v_41784;
assign v_42529 = v_41784;
assign v_42530 = ~v_815;
assign v_42531 = ~v_41788;
assign v_42532 = v_41788;
assign v_42533 = ~v_41791;
assign v_42534 = ~v_820;
assign v_42535 = v_820;
assign v_42536 = ~v_41795;
assign v_42537 = ~v_824;
assign v_42538 = v_824;
assign v_42539 = ~v_41799;
assign v_42540 = ~v_828;
assign v_42541 = v_828;
assign v_42542 = ~v_41803;
assign v_42543 = ~v_832;
assign v_42544 = v_832;
assign v_42545 = ~v_41807;
assign v_42546 = ~v_836;
assign v_42547 = v_836;
assign v_42548 = ~v_41811;
assign v_42549 = ~v_840;
assign v_42550 = v_840;
assign v_42551 = ~v_41815;
assign v_42552 = ~v_844;
assign v_42553 = v_844;
assign v_42554 = ~v_41819;
assign v_42555 = ~v_848;
assign v_42556 = v_848;
assign v_42557 = ~v_41823;
assign v_42558 = ~v_852;
assign v_42559 = v_852;
assign v_42560 = ~v_41827;
assign v_42561 = ~v_856;
assign v_42562 = v_856;
assign v_42563 = ~v_41831;
assign v_42564 = ~v_860;
assign v_42565 = v_860;
assign v_42566 = ~v_41835;
assign v_42567 = ~v_864;
assign v_42568 = v_864;
assign v_42569 = ~v_41839;
assign v_42570 = ~v_868;
assign v_42571 = v_42570;
assign v_42573 = v_42572;
assign v_42575 = v_42567 & v_42574;
assign v_42577 = v_41835;
assign v_42579 = v_42576 & v_42578;
assign v_42581 = v_42564 & v_42580;
assign v_42583 = v_41831;
assign v_42585 = v_42582 & v_42584;
assign v_42587 = v_42561 & v_42586;
assign v_42589 = v_41827;
assign v_42591 = v_42588 & v_42590;
assign v_42593 = v_42558 & v_42592;
assign v_42595 = v_41823;
assign v_42597 = v_42594 & v_42596;
assign v_42599 = v_42555 & v_42598;
assign v_42601 = v_41819;
assign v_42603 = v_42600 & v_42602;
assign v_42605 = v_42552 & v_42604;
assign v_42607 = v_41815;
assign v_42609 = v_42606 & v_42608;
assign v_42611 = v_42549 & v_42610;
assign v_42613 = v_41811;
assign v_42615 = v_42612 & v_42614;
assign v_42617 = v_42546 & v_42616;
assign v_42619 = v_41807;
assign v_42621 = v_42618 & v_42620;
assign v_42623 = v_42543 & v_42622;
assign v_42625 = v_41803;
assign v_42627 = v_42624 & v_42626;
assign v_42629 = v_42540 & v_42628;
assign v_42631 = v_41799;
assign v_42633 = v_42630 & v_42632;
assign v_42635 = v_42537 & v_42634;
assign v_42637 = v_41795;
assign v_42639 = v_42636 & v_42638;
assign v_42641 = v_42534 & v_42640;
assign v_42643 = v_41791;
assign v_42645 = v_42642 & v_42644;
assign v_42647 = v_42531 & v_42646;
assign v_42649 = v_815;
assign v_42651 = v_42648 & v_42650;
assign v_42653 = v_42528 & v_42652;
assign v_42655 = v_811;
assign v_42657 = v_42654 & v_42656;
assign v_42659 = v_42525 & v_42658;
assign v_42661 = v_807;
assign v_42663 = v_42660 & v_42662;
assign v_42665 = v_42522 & v_42664;
assign v_42667 = v_803;
assign v_42669 = v_42666 & v_42668;
assign v_42670 = v_42669;
assign v_42672 = v_41839;
assign v_42673 = v_868;
assign v_42674 = v_42673;
assign v_42675 = v_42672 & v_42674;
assign v_42676 = v_42675;
assign v_42677 = v_42567 & v_42676;
assign v_42679 = v_42577 & v_42678;
assign v_42680 = v_42566 & v_42676;
assign v_42682 = v_42564 & v_42681;
assign v_42684 = v_42583 & v_42683;
assign v_42685 = v_42563 & v_42681;
assign v_42687 = v_42561 & v_42686;
assign v_42689 = v_42589 & v_42688;
assign v_42690 = v_42560 & v_42686;
assign v_42692 = v_42558 & v_42691;
assign v_42694 = v_42595 & v_42693;
assign v_42695 = v_42557 & v_42691;
assign v_42697 = v_42555 & v_42696;
assign v_42699 = v_42601 & v_42698;
assign v_42700 = v_42554 & v_42696;
assign v_42702 = v_42552 & v_42701;
assign v_42704 = v_42607 & v_42703;
assign v_42705 = v_42551 & v_42701;
assign v_42707 = v_42549 & v_42706;
assign v_42709 = v_42613 & v_42708;
assign v_42710 = v_42548 & v_42706;
assign v_42712 = v_42546 & v_42711;
assign v_42714 = v_42619 & v_42713;
assign v_42715 = v_42545 & v_42711;
assign v_42717 = v_42543 & v_42716;
assign v_42719 = v_42625 & v_42718;
assign v_42720 = v_42542 & v_42716;
assign v_42722 = v_42540 & v_42721;
assign v_42724 = v_42631 & v_42723;
assign v_42725 = v_42539 & v_42721;
assign v_42727 = v_42537 & v_42726;
assign v_42729 = v_42637 & v_42728;
assign v_42730 = v_42536 & v_42726;
assign v_42732 = v_42534 & v_42731;
assign v_42734 = v_42643 & v_42733;
assign v_42735 = v_42533 & v_42731;
assign v_42737 = v_42531 & v_42736;
assign v_42739 = v_42649 & v_42738;
assign v_42740 = v_42530 & v_42736;
assign v_42742 = v_42528 & v_42741;
assign v_42744 = v_42655 & v_42743;
assign v_42745 = v_42527 & v_42741;
assign v_42747 = v_42525 & v_42746;
assign v_42749 = v_42661 & v_42748;
assign v_42750 = v_42524 & v_42746;
assign v_42752 = v_42522 & v_42751;
assign v_42754 = v_42667 & v_42753;
assign v_42755 = v_42521 & v_42751;
assign v_42757 = v_42756;
assign v_42759 = v_42671 & v_42758;
assign v_42760 = v_42759;
assign v_42762 = v_42761;
assign v_42764 = ~v_1063;
assign v_42765 = ~v_41776;
assign v_42766 = v_41776;
assign v_42767 = ~v_1067;
assign v_42768 = ~v_41780;
assign v_42769 = v_41780;
assign v_42770 = ~v_1071;
assign v_42771 = ~v_41784;
assign v_42772 = v_41784;
assign v_42773 = ~v_1075;
assign v_42774 = ~v_41788;
assign v_42775 = v_41788;
assign v_42776 = ~v_41791;
assign v_42777 = ~v_1080;
assign v_42778 = v_1080;
assign v_42779 = ~v_41795;
assign v_42780 = ~v_1084;
assign v_42781 = v_1084;
assign v_42782 = ~v_41799;
assign v_42783 = ~v_1088;
assign v_42784 = v_1088;
assign v_42785 = ~v_41803;
assign v_42786 = ~v_1092;
assign v_42787 = v_1092;
assign v_42788 = ~v_41807;
assign v_42789 = ~v_1096;
assign v_42790 = v_1096;
assign v_42791 = ~v_41811;
assign v_42792 = ~v_1100;
assign v_42793 = v_1100;
assign v_42794 = ~v_41815;
assign v_42795 = ~v_1104;
assign v_42796 = v_1104;
assign v_42797 = ~v_41819;
assign v_42798 = ~v_1108;
assign v_42799 = v_1108;
assign v_42800 = ~v_41823;
assign v_42801 = ~v_1112;
assign v_42802 = v_1112;
assign v_42803 = ~v_41827;
assign v_42804 = ~v_1116;
assign v_42805 = v_1116;
assign v_42806 = ~v_41831;
assign v_42807 = ~v_1120;
assign v_42808 = v_1120;
assign v_42809 = ~v_41835;
assign v_42810 = ~v_1124;
assign v_42811 = v_1124;
assign v_42812 = ~v_41839;
assign v_42813 = ~v_1128;
assign v_42814 = v_42813;
assign v_42816 = v_42815;
assign v_42818 = v_42810 & v_42817;
assign v_42820 = v_41835;
assign v_42822 = v_42819 & v_42821;
assign v_42824 = v_42807 & v_42823;
assign v_42826 = v_41831;
assign v_42828 = v_42825 & v_42827;
assign v_42830 = v_42804 & v_42829;
assign v_42832 = v_41827;
assign v_42834 = v_42831 & v_42833;
assign v_42836 = v_42801 & v_42835;
assign v_42838 = v_41823;
assign v_42840 = v_42837 & v_42839;
assign v_42842 = v_42798 & v_42841;
assign v_42844 = v_41819;
assign v_42846 = v_42843 & v_42845;
assign v_42848 = v_42795 & v_42847;
assign v_42850 = v_41815;
assign v_42852 = v_42849 & v_42851;
assign v_42854 = v_42792 & v_42853;
assign v_42856 = v_41811;
assign v_42858 = v_42855 & v_42857;
assign v_42860 = v_42789 & v_42859;
assign v_42862 = v_41807;
assign v_42864 = v_42861 & v_42863;
assign v_42866 = v_42786 & v_42865;
assign v_42868 = v_41803;
assign v_42870 = v_42867 & v_42869;
assign v_42872 = v_42783 & v_42871;
assign v_42874 = v_41799;
assign v_42876 = v_42873 & v_42875;
assign v_42878 = v_42780 & v_42877;
assign v_42880 = v_41795;
assign v_42882 = v_42879 & v_42881;
assign v_42884 = v_42777 & v_42883;
assign v_42886 = v_41791;
assign v_42888 = v_42885 & v_42887;
assign v_42890 = v_42774 & v_42889;
assign v_42892 = v_1075;
assign v_42894 = v_42891 & v_42893;
assign v_42896 = v_42771 & v_42895;
assign v_42898 = v_1071;
assign v_42900 = v_42897 & v_42899;
assign v_42902 = v_42768 & v_42901;
assign v_42904 = v_1067;
assign v_42906 = v_42903 & v_42905;
assign v_42908 = v_42765 & v_42907;
assign v_42910 = v_1063;
assign v_42912 = v_42909 & v_42911;
assign v_42913 = v_42912;
assign v_42915 = v_41839;
assign v_42916 = v_1128;
assign v_42917 = v_42916;
assign v_42918 = v_42915 & v_42917;
assign v_42919 = v_42918;
assign v_42920 = v_42810 & v_42919;
assign v_42922 = v_42820 & v_42921;
assign v_42923 = v_42809 & v_42919;
assign v_42925 = v_42807 & v_42924;
assign v_42927 = v_42826 & v_42926;
assign v_42928 = v_42806 & v_42924;
assign v_42930 = v_42804 & v_42929;
assign v_42932 = v_42832 & v_42931;
assign v_42933 = v_42803 & v_42929;
assign v_42935 = v_42801 & v_42934;
assign v_42937 = v_42838 & v_42936;
assign v_42938 = v_42800 & v_42934;
assign v_42940 = v_42798 & v_42939;
assign v_42942 = v_42844 & v_42941;
assign v_42943 = v_42797 & v_42939;
assign v_42945 = v_42795 & v_42944;
assign v_42947 = v_42850 & v_42946;
assign v_42948 = v_42794 & v_42944;
assign v_42950 = v_42792 & v_42949;
assign v_42952 = v_42856 & v_42951;
assign v_42953 = v_42791 & v_42949;
assign v_42955 = v_42789 & v_42954;
assign v_42957 = v_42862 & v_42956;
assign v_42958 = v_42788 & v_42954;
assign v_42960 = v_42786 & v_42959;
assign v_42962 = v_42868 & v_42961;
assign v_42963 = v_42785 & v_42959;
assign v_42965 = v_42783 & v_42964;
assign v_42967 = v_42874 & v_42966;
assign v_42968 = v_42782 & v_42964;
assign v_42970 = v_42780 & v_42969;
assign v_42972 = v_42880 & v_42971;
assign v_42973 = v_42779 & v_42969;
assign v_42975 = v_42777 & v_42974;
assign v_42977 = v_42886 & v_42976;
assign v_42978 = v_42776 & v_42974;
assign v_42980 = v_42774 & v_42979;
assign v_42982 = v_42892 & v_42981;
assign v_42983 = v_42773 & v_42979;
assign v_42985 = v_42771 & v_42984;
assign v_42987 = v_42898 & v_42986;
assign v_42988 = v_42770 & v_42984;
assign v_42990 = v_42768 & v_42989;
assign v_42992 = v_42904 & v_42991;
assign v_42993 = v_42767 & v_42989;
assign v_42995 = v_42765 & v_42994;
assign v_42997 = v_42910 & v_42996;
assign v_42998 = v_42764 & v_42994;
assign v_43000 = v_42999;
assign v_43002 = v_42914 & v_43001;
assign v_43003 = v_43002;
assign v_43005 = v_43004;
assign v_43007 = ~v_1323;
assign v_43008 = ~v_41776;
assign v_43009 = v_41776;
assign v_43010 = ~v_1327;
assign v_43011 = ~v_41780;
assign v_43012 = v_41780;
assign v_43013 = ~v_1331;
assign v_43014 = ~v_41784;
assign v_43015 = v_41784;
assign v_43016 = ~v_1335;
assign v_43017 = ~v_41788;
assign v_43018 = v_41788;
assign v_43019 = ~v_41791;
assign v_43020 = ~v_1340;
assign v_43021 = v_1340;
assign v_43022 = ~v_41795;
assign v_43023 = ~v_1344;
assign v_43024 = v_1344;
assign v_43025 = ~v_41799;
assign v_43026 = ~v_1348;
assign v_43027 = v_1348;
assign v_43028 = ~v_41803;
assign v_43029 = ~v_1352;
assign v_43030 = v_1352;
assign v_43031 = ~v_41807;
assign v_43032 = ~v_1356;
assign v_43033 = v_1356;
assign v_43034 = ~v_41811;
assign v_43035 = ~v_1360;
assign v_43036 = v_1360;
assign v_43037 = ~v_41815;
assign v_43038 = ~v_1364;
assign v_43039 = v_1364;
assign v_43040 = ~v_41819;
assign v_43041 = ~v_1368;
assign v_43042 = v_1368;
assign v_43043 = ~v_41823;
assign v_43044 = ~v_1372;
assign v_43045 = v_1372;
assign v_43046 = ~v_41827;
assign v_43047 = ~v_1376;
assign v_43048 = v_1376;
assign v_43049 = ~v_41831;
assign v_43050 = ~v_1380;
assign v_43051 = v_1380;
assign v_43052 = ~v_41835;
assign v_43053 = ~v_1384;
assign v_43054 = v_1384;
assign v_43055 = ~v_41839;
assign v_43056 = ~v_1388;
assign v_43057 = v_43056;
assign v_43059 = v_43058;
assign v_43061 = v_43053 & v_43060;
assign v_43063 = v_41835;
assign v_43065 = v_43062 & v_43064;
assign v_43067 = v_43050 & v_43066;
assign v_43069 = v_41831;
assign v_43071 = v_43068 & v_43070;
assign v_43073 = v_43047 & v_43072;
assign v_43075 = v_41827;
assign v_43077 = v_43074 & v_43076;
assign v_43079 = v_43044 & v_43078;
assign v_43081 = v_41823;
assign v_43083 = v_43080 & v_43082;
assign v_43085 = v_43041 & v_43084;
assign v_43087 = v_41819;
assign v_43089 = v_43086 & v_43088;
assign v_43091 = v_43038 & v_43090;
assign v_43093 = v_41815;
assign v_43095 = v_43092 & v_43094;
assign v_43097 = v_43035 & v_43096;
assign v_43099 = v_41811;
assign v_43101 = v_43098 & v_43100;
assign v_43103 = v_43032 & v_43102;
assign v_43105 = v_41807;
assign v_43107 = v_43104 & v_43106;
assign v_43109 = v_43029 & v_43108;
assign v_43111 = v_41803;
assign v_43113 = v_43110 & v_43112;
assign v_43115 = v_43026 & v_43114;
assign v_43117 = v_41799;
assign v_43119 = v_43116 & v_43118;
assign v_43121 = v_43023 & v_43120;
assign v_43123 = v_41795;
assign v_43125 = v_43122 & v_43124;
assign v_43127 = v_43020 & v_43126;
assign v_43129 = v_41791;
assign v_43131 = v_43128 & v_43130;
assign v_43133 = v_43017 & v_43132;
assign v_43135 = v_1335;
assign v_43137 = v_43134 & v_43136;
assign v_43139 = v_43014 & v_43138;
assign v_43141 = v_1331;
assign v_43143 = v_43140 & v_43142;
assign v_43145 = v_43011 & v_43144;
assign v_43147 = v_1327;
assign v_43149 = v_43146 & v_43148;
assign v_43151 = v_43008 & v_43150;
assign v_43153 = v_1323;
assign v_43155 = v_43152 & v_43154;
assign v_43156 = v_43155;
assign v_43158 = v_41839;
assign v_43159 = v_1388;
assign v_43160 = v_43159;
assign v_43161 = v_43158 & v_43160;
assign v_43162 = v_43161;
assign v_43163 = v_43053 & v_43162;
assign v_43165 = v_43063 & v_43164;
assign v_43166 = v_43052 & v_43162;
assign v_43168 = v_43050 & v_43167;
assign v_43170 = v_43069 & v_43169;
assign v_43171 = v_43049 & v_43167;
assign v_43173 = v_43047 & v_43172;
assign v_43175 = v_43075 & v_43174;
assign v_43176 = v_43046 & v_43172;
assign v_43178 = v_43044 & v_43177;
assign v_43180 = v_43081 & v_43179;
assign v_43181 = v_43043 & v_43177;
assign v_43183 = v_43041 & v_43182;
assign v_43185 = v_43087 & v_43184;
assign v_43186 = v_43040 & v_43182;
assign v_43188 = v_43038 & v_43187;
assign v_43190 = v_43093 & v_43189;
assign v_43191 = v_43037 & v_43187;
assign v_43193 = v_43035 & v_43192;
assign v_43195 = v_43099 & v_43194;
assign v_43196 = v_43034 & v_43192;
assign v_43198 = v_43032 & v_43197;
assign v_43200 = v_43105 & v_43199;
assign v_43201 = v_43031 & v_43197;
assign v_43203 = v_43029 & v_43202;
assign v_43205 = v_43111 & v_43204;
assign v_43206 = v_43028 & v_43202;
assign v_43208 = v_43026 & v_43207;
assign v_43210 = v_43117 & v_43209;
assign v_43211 = v_43025 & v_43207;
assign v_43213 = v_43023 & v_43212;
assign v_43215 = v_43123 & v_43214;
assign v_43216 = v_43022 & v_43212;
assign v_43218 = v_43020 & v_43217;
assign v_43220 = v_43129 & v_43219;
assign v_43221 = v_43019 & v_43217;
assign v_43223 = v_43017 & v_43222;
assign v_43225 = v_43135 & v_43224;
assign v_43226 = v_43016 & v_43222;
assign v_43228 = v_43014 & v_43227;
assign v_43230 = v_43141 & v_43229;
assign v_43231 = v_43013 & v_43227;
assign v_43233 = v_43011 & v_43232;
assign v_43235 = v_43147 & v_43234;
assign v_43236 = v_43010 & v_43232;
assign v_43238 = v_43008 & v_43237;
assign v_43240 = v_43153 & v_43239;
assign v_43241 = v_43007 & v_43237;
assign v_43243 = v_43242;
assign v_43245 = v_43157 & v_43244;
assign v_43246 = v_43245;
assign v_43248 = v_43247;
assign v_43250 = ~v_1583;
assign v_43251 = ~v_41776;
assign v_43252 = v_41776;
assign v_43253 = ~v_1587;
assign v_43254 = ~v_41780;
assign v_43255 = v_41780;
assign v_43256 = ~v_1591;
assign v_43257 = ~v_41784;
assign v_43258 = v_41784;
assign v_43259 = ~v_1595;
assign v_43260 = ~v_41788;
assign v_43261 = v_41788;
assign v_43262 = ~v_41791;
assign v_43263 = ~v_1600;
assign v_43264 = v_1600;
assign v_43265 = ~v_41795;
assign v_43266 = ~v_1604;
assign v_43267 = v_1604;
assign v_43268 = ~v_41799;
assign v_43269 = ~v_1608;
assign v_43270 = v_1608;
assign v_43271 = ~v_41803;
assign v_43272 = ~v_1612;
assign v_43273 = v_1612;
assign v_43274 = ~v_41807;
assign v_43275 = ~v_1616;
assign v_43276 = v_1616;
assign v_43277 = ~v_41811;
assign v_43278 = ~v_1620;
assign v_43279 = v_1620;
assign v_43280 = ~v_41815;
assign v_43281 = ~v_1624;
assign v_43282 = v_1624;
assign v_43283 = ~v_41819;
assign v_43284 = ~v_1628;
assign v_43285 = v_1628;
assign v_43286 = ~v_41823;
assign v_43287 = ~v_1632;
assign v_43288 = v_1632;
assign v_43289 = ~v_41827;
assign v_43290 = ~v_1636;
assign v_43291 = v_1636;
assign v_43292 = ~v_41831;
assign v_43293 = ~v_1640;
assign v_43294 = v_1640;
assign v_43295 = ~v_41835;
assign v_43296 = ~v_1644;
assign v_43297 = v_1644;
assign v_43298 = ~v_41839;
assign v_43299 = ~v_1648;
assign v_43300 = v_43299;
assign v_43302 = v_43301;
assign v_43304 = v_43296 & v_43303;
assign v_43306 = v_41835;
assign v_43308 = v_43305 & v_43307;
assign v_43310 = v_43293 & v_43309;
assign v_43312 = v_41831;
assign v_43314 = v_43311 & v_43313;
assign v_43316 = v_43290 & v_43315;
assign v_43318 = v_41827;
assign v_43320 = v_43317 & v_43319;
assign v_43322 = v_43287 & v_43321;
assign v_43324 = v_41823;
assign v_43326 = v_43323 & v_43325;
assign v_43328 = v_43284 & v_43327;
assign v_43330 = v_41819;
assign v_43332 = v_43329 & v_43331;
assign v_43334 = v_43281 & v_43333;
assign v_43336 = v_41815;
assign v_43338 = v_43335 & v_43337;
assign v_43340 = v_43278 & v_43339;
assign v_43342 = v_41811;
assign v_43344 = v_43341 & v_43343;
assign v_43346 = v_43275 & v_43345;
assign v_43348 = v_41807;
assign v_43350 = v_43347 & v_43349;
assign v_43352 = v_43272 & v_43351;
assign v_43354 = v_41803;
assign v_43356 = v_43353 & v_43355;
assign v_43358 = v_43269 & v_43357;
assign v_43360 = v_41799;
assign v_43362 = v_43359 & v_43361;
assign v_43364 = v_43266 & v_43363;
assign v_43366 = v_41795;
assign v_43368 = v_43365 & v_43367;
assign v_43370 = v_43263 & v_43369;
assign v_43372 = v_41791;
assign v_43374 = v_43371 & v_43373;
assign v_43376 = v_43260 & v_43375;
assign v_43378 = v_1595;
assign v_43380 = v_43377 & v_43379;
assign v_43382 = v_43257 & v_43381;
assign v_43384 = v_1591;
assign v_43386 = v_43383 & v_43385;
assign v_43388 = v_43254 & v_43387;
assign v_43390 = v_1587;
assign v_43392 = v_43389 & v_43391;
assign v_43394 = v_43251 & v_43393;
assign v_43396 = v_1583;
assign v_43398 = v_43395 & v_43397;
assign v_43399 = v_43398;
assign v_43401 = v_41839;
assign v_43402 = v_1648;
assign v_43403 = v_43402;
assign v_43404 = v_43401 & v_43403;
assign v_43405 = v_43404;
assign v_43406 = v_43296 & v_43405;
assign v_43408 = v_43306 & v_43407;
assign v_43409 = v_43295 & v_43405;
assign v_43411 = v_43293 & v_43410;
assign v_43413 = v_43312 & v_43412;
assign v_43414 = v_43292 & v_43410;
assign v_43416 = v_43290 & v_43415;
assign v_43418 = v_43318 & v_43417;
assign v_43419 = v_43289 & v_43415;
assign v_43421 = v_43287 & v_43420;
assign v_43423 = v_43324 & v_43422;
assign v_43424 = v_43286 & v_43420;
assign v_43426 = v_43284 & v_43425;
assign v_43428 = v_43330 & v_43427;
assign v_43429 = v_43283 & v_43425;
assign v_43431 = v_43281 & v_43430;
assign v_43433 = v_43336 & v_43432;
assign v_43434 = v_43280 & v_43430;
assign v_43436 = v_43278 & v_43435;
assign v_43438 = v_43342 & v_43437;
assign v_43439 = v_43277 & v_43435;
assign v_43441 = v_43275 & v_43440;
assign v_43443 = v_43348 & v_43442;
assign v_43444 = v_43274 & v_43440;
assign v_43446 = v_43272 & v_43445;
assign v_43448 = v_43354 & v_43447;
assign v_43449 = v_43271 & v_43445;
assign v_43451 = v_43269 & v_43450;
assign v_43453 = v_43360 & v_43452;
assign v_43454 = v_43268 & v_43450;
assign v_43456 = v_43266 & v_43455;
assign v_43458 = v_43366 & v_43457;
assign v_43459 = v_43265 & v_43455;
assign v_43461 = v_43263 & v_43460;
assign v_43463 = v_43372 & v_43462;
assign v_43464 = v_43262 & v_43460;
assign v_43466 = v_43260 & v_43465;
assign v_43468 = v_43378 & v_43467;
assign v_43469 = v_43259 & v_43465;
assign v_43471 = v_43257 & v_43470;
assign v_43473 = v_43384 & v_43472;
assign v_43474 = v_43256 & v_43470;
assign v_43476 = v_43254 & v_43475;
assign v_43478 = v_43390 & v_43477;
assign v_43479 = v_43253 & v_43475;
assign v_43481 = v_43251 & v_43480;
assign v_43483 = v_43396 & v_43482;
assign v_43484 = v_43250 & v_43480;
assign v_43486 = v_43485;
assign v_43488 = v_43400 & v_43487;
assign v_43489 = v_43488;
assign v_43491 = v_43490;
assign v_43493 = ~v_1843;
assign v_43494 = ~v_41776;
assign v_43495 = v_41776;
assign v_43496 = ~v_1847;
assign v_43497 = ~v_41780;
assign v_43498 = v_41780;
assign v_43499 = ~v_1851;
assign v_43500 = ~v_41784;
assign v_43501 = v_41784;
assign v_43502 = ~v_1855;
assign v_43503 = ~v_41788;
assign v_43504 = v_41788;
assign v_43505 = ~v_41791;
assign v_43506 = ~v_1860;
assign v_43507 = v_1860;
assign v_43508 = ~v_41795;
assign v_43509 = ~v_1864;
assign v_43510 = v_1864;
assign v_43511 = ~v_41799;
assign v_43512 = ~v_1868;
assign v_43513 = v_1868;
assign v_43514 = ~v_41803;
assign v_43515 = ~v_1872;
assign v_43516 = v_1872;
assign v_43517 = ~v_41807;
assign v_43518 = ~v_1876;
assign v_43519 = v_1876;
assign v_43520 = ~v_41811;
assign v_43521 = ~v_1880;
assign v_43522 = v_1880;
assign v_43523 = ~v_41815;
assign v_43524 = ~v_1884;
assign v_43525 = v_1884;
assign v_43526 = ~v_41819;
assign v_43527 = ~v_1888;
assign v_43528 = v_1888;
assign v_43529 = ~v_41823;
assign v_43530 = ~v_1892;
assign v_43531 = v_1892;
assign v_43532 = ~v_41827;
assign v_43533 = ~v_1896;
assign v_43534 = v_1896;
assign v_43535 = ~v_41831;
assign v_43536 = ~v_1900;
assign v_43537 = v_1900;
assign v_43538 = ~v_41835;
assign v_43539 = ~v_1904;
assign v_43540 = v_1904;
assign v_43541 = ~v_41839;
assign v_43542 = ~v_1908;
assign v_43543 = v_43542;
assign v_43545 = v_43544;
assign v_43547 = v_43539 & v_43546;
assign v_43549 = v_41835;
assign v_43551 = v_43548 & v_43550;
assign v_43553 = v_43536 & v_43552;
assign v_43555 = v_41831;
assign v_43557 = v_43554 & v_43556;
assign v_43559 = v_43533 & v_43558;
assign v_43561 = v_41827;
assign v_43563 = v_43560 & v_43562;
assign v_43565 = v_43530 & v_43564;
assign v_43567 = v_41823;
assign v_43569 = v_43566 & v_43568;
assign v_43571 = v_43527 & v_43570;
assign v_43573 = v_41819;
assign v_43575 = v_43572 & v_43574;
assign v_43577 = v_43524 & v_43576;
assign v_43579 = v_41815;
assign v_43581 = v_43578 & v_43580;
assign v_43583 = v_43521 & v_43582;
assign v_43585 = v_41811;
assign v_43587 = v_43584 & v_43586;
assign v_43589 = v_43518 & v_43588;
assign v_43591 = v_41807;
assign v_43593 = v_43590 & v_43592;
assign v_43595 = v_43515 & v_43594;
assign v_43597 = v_41803;
assign v_43599 = v_43596 & v_43598;
assign v_43601 = v_43512 & v_43600;
assign v_43603 = v_41799;
assign v_43605 = v_43602 & v_43604;
assign v_43607 = v_43509 & v_43606;
assign v_43609 = v_41795;
assign v_43611 = v_43608 & v_43610;
assign v_43613 = v_43506 & v_43612;
assign v_43615 = v_41791;
assign v_43617 = v_43614 & v_43616;
assign v_43619 = v_43503 & v_43618;
assign v_43621 = v_1855;
assign v_43623 = v_43620 & v_43622;
assign v_43625 = v_43500 & v_43624;
assign v_43627 = v_1851;
assign v_43629 = v_43626 & v_43628;
assign v_43631 = v_43497 & v_43630;
assign v_43633 = v_1847;
assign v_43635 = v_43632 & v_43634;
assign v_43637 = v_43494 & v_43636;
assign v_43639 = v_1843;
assign v_43641 = v_43638 & v_43640;
assign v_43642 = v_43641;
assign v_43644 = v_41839;
assign v_43645 = v_1908;
assign v_43646 = v_43645;
assign v_43647 = v_43644 & v_43646;
assign v_43648 = v_43647;
assign v_43649 = v_43539 & v_43648;
assign v_43651 = v_43549 & v_43650;
assign v_43652 = v_43538 & v_43648;
assign v_43654 = v_43536 & v_43653;
assign v_43656 = v_43555 & v_43655;
assign v_43657 = v_43535 & v_43653;
assign v_43659 = v_43533 & v_43658;
assign v_43661 = v_43561 & v_43660;
assign v_43662 = v_43532 & v_43658;
assign v_43664 = v_43530 & v_43663;
assign v_43666 = v_43567 & v_43665;
assign v_43667 = v_43529 & v_43663;
assign v_43669 = v_43527 & v_43668;
assign v_43671 = v_43573 & v_43670;
assign v_43672 = v_43526 & v_43668;
assign v_43674 = v_43524 & v_43673;
assign v_43676 = v_43579 & v_43675;
assign v_43677 = v_43523 & v_43673;
assign v_43679 = v_43521 & v_43678;
assign v_43681 = v_43585 & v_43680;
assign v_43682 = v_43520 & v_43678;
assign v_43684 = v_43518 & v_43683;
assign v_43686 = v_43591 & v_43685;
assign v_43687 = v_43517 & v_43683;
assign v_43689 = v_43515 & v_43688;
assign v_43691 = v_43597 & v_43690;
assign v_43692 = v_43514 & v_43688;
assign v_43694 = v_43512 & v_43693;
assign v_43696 = v_43603 & v_43695;
assign v_43697 = v_43511 & v_43693;
assign v_43699 = v_43509 & v_43698;
assign v_43701 = v_43609 & v_43700;
assign v_43702 = v_43508 & v_43698;
assign v_43704 = v_43506 & v_43703;
assign v_43706 = v_43615 & v_43705;
assign v_43707 = v_43505 & v_43703;
assign v_43709 = v_43503 & v_43708;
assign v_43711 = v_43621 & v_43710;
assign v_43712 = v_43502 & v_43708;
assign v_43714 = v_43500 & v_43713;
assign v_43716 = v_43627 & v_43715;
assign v_43717 = v_43499 & v_43713;
assign v_43719 = v_43497 & v_43718;
assign v_43721 = v_43633 & v_43720;
assign v_43722 = v_43496 & v_43718;
assign v_43724 = v_43494 & v_43723;
assign v_43726 = v_43639 & v_43725;
assign v_43727 = v_43493 & v_43723;
assign v_43729 = v_43728;
assign v_43731 = v_43643 & v_43730;
assign v_43732 = v_43731;
assign v_43734 = v_43733;
assign v_43736 = ~v_2103;
assign v_43737 = ~v_41776;
assign v_43738 = v_41776;
assign v_43739 = ~v_2107;
assign v_43740 = ~v_41780;
assign v_43741 = v_41780;
assign v_43742 = ~v_2111;
assign v_43743 = ~v_41784;
assign v_43744 = v_41784;
assign v_43745 = ~v_2115;
assign v_43746 = ~v_41788;
assign v_43747 = v_41788;
assign v_43748 = ~v_41791;
assign v_43749 = ~v_2120;
assign v_43750 = v_2120;
assign v_43751 = ~v_41795;
assign v_43752 = ~v_2124;
assign v_43753 = v_2124;
assign v_43754 = ~v_41799;
assign v_43755 = ~v_2128;
assign v_43756 = v_2128;
assign v_43757 = ~v_41803;
assign v_43758 = ~v_2132;
assign v_43759 = v_2132;
assign v_43760 = ~v_41807;
assign v_43761 = ~v_2136;
assign v_43762 = v_2136;
assign v_43763 = ~v_41811;
assign v_43764 = ~v_2140;
assign v_43765 = v_2140;
assign v_43766 = ~v_41815;
assign v_43767 = ~v_2144;
assign v_43768 = v_2144;
assign v_43769 = ~v_41819;
assign v_43770 = ~v_2148;
assign v_43771 = v_2148;
assign v_43772 = ~v_41823;
assign v_43773 = ~v_2152;
assign v_43774 = v_2152;
assign v_43775 = ~v_41827;
assign v_43776 = ~v_2156;
assign v_43777 = v_2156;
assign v_43778 = ~v_41831;
assign v_43779 = ~v_2160;
assign v_43780 = v_2160;
assign v_43781 = ~v_41835;
assign v_43782 = ~v_2164;
assign v_43783 = v_2164;
assign v_43784 = ~v_41839;
assign v_43785 = ~v_2168;
assign v_43786 = v_43785;
assign v_43788 = v_43787;
assign v_43790 = v_43782 & v_43789;
assign v_43792 = v_41835;
assign v_43794 = v_43791 & v_43793;
assign v_43796 = v_43779 & v_43795;
assign v_43798 = v_41831;
assign v_43800 = v_43797 & v_43799;
assign v_43802 = v_43776 & v_43801;
assign v_43804 = v_41827;
assign v_43806 = v_43803 & v_43805;
assign v_43808 = v_43773 & v_43807;
assign v_43810 = v_41823;
assign v_43812 = v_43809 & v_43811;
assign v_43814 = v_43770 & v_43813;
assign v_43816 = v_41819;
assign v_43818 = v_43815 & v_43817;
assign v_43820 = v_43767 & v_43819;
assign v_43822 = v_41815;
assign v_43824 = v_43821 & v_43823;
assign v_43826 = v_43764 & v_43825;
assign v_43828 = v_41811;
assign v_43830 = v_43827 & v_43829;
assign v_43832 = v_43761 & v_43831;
assign v_43834 = v_41807;
assign v_43836 = v_43833 & v_43835;
assign v_43838 = v_43758 & v_43837;
assign v_43840 = v_41803;
assign v_43842 = v_43839 & v_43841;
assign v_43844 = v_43755 & v_43843;
assign v_43846 = v_41799;
assign v_43848 = v_43845 & v_43847;
assign v_43850 = v_43752 & v_43849;
assign v_43852 = v_41795;
assign v_43854 = v_43851 & v_43853;
assign v_43856 = v_43749 & v_43855;
assign v_43858 = v_41791;
assign v_43860 = v_43857 & v_43859;
assign v_43862 = v_43746 & v_43861;
assign v_43864 = v_2115;
assign v_43866 = v_43863 & v_43865;
assign v_43868 = v_43743 & v_43867;
assign v_43870 = v_2111;
assign v_43872 = v_43869 & v_43871;
assign v_43874 = v_43740 & v_43873;
assign v_43876 = v_2107;
assign v_43878 = v_43875 & v_43877;
assign v_43880 = v_43737 & v_43879;
assign v_43882 = v_2103;
assign v_43884 = v_43881 & v_43883;
assign v_43885 = v_43884;
assign v_43887 = v_41839;
assign v_43888 = v_2168;
assign v_43889 = v_43888;
assign v_43890 = v_43887 & v_43889;
assign v_43891 = v_43890;
assign v_43892 = v_43782 & v_43891;
assign v_43894 = v_43792 & v_43893;
assign v_43895 = v_43781 & v_43891;
assign v_43897 = v_43779 & v_43896;
assign v_43899 = v_43798 & v_43898;
assign v_43900 = v_43778 & v_43896;
assign v_43902 = v_43776 & v_43901;
assign v_43904 = v_43804 & v_43903;
assign v_43905 = v_43775 & v_43901;
assign v_43907 = v_43773 & v_43906;
assign v_43909 = v_43810 & v_43908;
assign v_43910 = v_43772 & v_43906;
assign v_43912 = v_43770 & v_43911;
assign v_43914 = v_43816 & v_43913;
assign v_43915 = v_43769 & v_43911;
assign v_43917 = v_43767 & v_43916;
assign v_43919 = v_43822 & v_43918;
assign v_43920 = v_43766 & v_43916;
assign v_43922 = v_43764 & v_43921;
assign v_43924 = v_43828 & v_43923;
assign v_43925 = v_43763 & v_43921;
assign v_43927 = v_43761 & v_43926;
assign v_43929 = v_43834 & v_43928;
assign v_43930 = v_43760 & v_43926;
assign v_43932 = v_43758 & v_43931;
assign v_43934 = v_43840 & v_43933;
assign v_43935 = v_43757 & v_43931;
assign v_43937 = v_43755 & v_43936;
assign v_43939 = v_43846 & v_43938;
assign v_43940 = v_43754 & v_43936;
assign v_43942 = v_43752 & v_43941;
assign v_43944 = v_43852 & v_43943;
assign v_43945 = v_43751 & v_43941;
assign v_43947 = v_43749 & v_43946;
assign v_43949 = v_43858 & v_43948;
assign v_43950 = v_43748 & v_43946;
assign v_43952 = v_43746 & v_43951;
assign v_43954 = v_43864 & v_43953;
assign v_43955 = v_43745 & v_43951;
assign v_43957 = v_43743 & v_43956;
assign v_43959 = v_43870 & v_43958;
assign v_43960 = v_43742 & v_43956;
assign v_43962 = v_43740 & v_43961;
assign v_43964 = v_43876 & v_43963;
assign v_43965 = v_43739 & v_43961;
assign v_43967 = v_43737 & v_43966;
assign v_43969 = v_43882 & v_43968;
assign v_43970 = v_43736 & v_43966;
assign v_43972 = v_43971;
assign v_43974 = v_43886 & v_43973;
assign v_43975 = v_43974;
assign v_43977 = v_43976;
assign v_43979 = ~v_2363;
assign v_43980 = ~v_41776;
assign v_43981 = v_41776;
assign v_43982 = ~v_2367;
assign v_43983 = ~v_41780;
assign v_43984 = v_41780;
assign v_43985 = ~v_2371;
assign v_43986 = ~v_41784;
assign v_43987 = v_41784;
assign v_43988 = ~v_2375;
assign v_43989 = ~v_41788;
assign v_43990 = v_41788;
assign v_43991 = ~v_41791;
assign v_43992 = ~v_2380;
assign v_43993 = v_2380;
assign v_43994 = ~v_41795;
assign v_43995 = ~v_2384;
assign v_43996 = v_2384;
assign v_43997 = ~v_41799;
assign v_43998 = ~v_2388;
assign v_43999 = v_2388;
assign v_44000 = ~v_41803;
assign v_44001 = ~v_2392;
assign v_44002 = v_2392;
assign v_44003 = ~v_41807;
assign v_44004 = ~v_2396;
assign v_44005 = v_2396;
assign v_44006 = ~v_41811;
assign v_44007 = ~v_2400;
assign v_44008 = v_2400;
assign v_44009 = ~v_41815;
assign v_44010 = ~v_2404;
assign v_44011 = v_2404;
assign v_44012 = ~v_41819;
assign v_44013 = ~v_2408;
assign v_44014 = v_2408;
assign v_44015 = ~v_41823;
assign v_44016 = ~v_2412;
assign v_44017 = v_2412;
assign v_44018 = ~v_41827;
assign v_44019 = ~v_2416;
assign v_44020 = v_2416;
assign v_44021 = ~v_41831;
assign v_44022 = ~v_2420;
assign v_44023 = v_2420;
assign v_44024 = ~v_41835;
assign v_44025 = ~v_2424;
assign v_44026 = v_2424;
assign v_44027 = ~v_41839;
assign v_44028 = ~v_2428;
assign v_44029 = v_44028;
assign v_44031 = v_44030;
assign v_44033 = v_44025 & v_44032;
assign v_44035 = v_41835;
assign v_44037 = v_44034 & v_44036;
assign v_44039 = v_44022 & v_44038;
assign v_44041 = v_41831;
assign v_44043 = v_44040 & v_44042;
assign v_44045 = v_44019 & v_44044;
assign v_44047 = v_41827;
assign v_44049 = v_44046 & v_44048;
assign v_44051 = v_44016 & v_44050;
assign v_44053 = v_41823;
assign v_44055 = v_44052 & v_44054;
assign v_44057 = v_44013 & v_44056;
assign v_44059 = v_41819;
assign v_44061 = v_44058 & v_44060;
assign v_44063 = v_44010 & v_44062;
assign v_44065 = v_41815;
assign v_44067 = v_44064 & v_44066;
assign v_44069 = v_44007 & v_44068;
assign v_44071 = v_41811;
assign v_44073 = v_44070 & v_44072;
assign v_44075 = v_44004 & v_44074;
assign v_44077 = v_41807;
assign v_44079 = v_44076 & v_44078;
assign v_44081 = v_44001 & v_44080;
assign v_44083 = v_41803;
assign v_44085 = v_44082 & v_44084;
assign v_44087 = v_43998 & v_44086;
assign v_44089 = v_41799;
assign v_44091 = v_44088 & v_44090;
assign v_44093 = v_43995 & v_44092;
assign v_44095 = v_41795;
assign v_44097 = v_44094 & v_44096;
assign v_44099 = v_43992 & v_44098;
assign v_44101 = v_41791;
assign v_44103 = v_44100 & v_44102;
assign v_44105 = v_43989 & v_44104;
assign v_44107 = v_2375;
assign v_44109 = v_44106 & v_44108;
assign v_44111 = v_43986 & v_44110;
assign v_44113 = v_2371;
assign v_44115 = v_44112 & v_44114;
assign v_44117 = v_43983 & v_44116;
assign v_44119 = v_2367;
assign v_44121 = v_44118 & v_44120;
assign v_44123 = v_43980 & v_44122;
assign v_44125 = v_2363;
assign v_44127 = v_44124 & v_44126;
assign v_44128 = v_44127;
assign v_44130 = v_41839;
assign v_44131 = v_2428;
assign v_44132 = v_44131;
assign v_44133 = v_44130 & v_44132;
assign v_44134 = v_44133;
assign v_44135 = v_44025 & v_44134;
assign v_44137 = v_44035 & v_44136;
assign v_44138 = v_44024 & v_44134;
assign v_44140 = v_44022 & v_44139;
assign v_44142 = v_44041 & v_44141;
assign v_44143 = v_44021 & v_44139;
assign v_44145 = v_44019 & v_44144;
assign v_44147 = v_44047 & v_44146;
assign v_44148 = v_44018 & v_44144;
assign v_44150 = v_44016 & v_44149;
assign v_44152 = v_44053 & v_44151;
assign v_44153 = v_44015 & v_44149;
assign v_44155 = v_44013 & v_44154;
assign v_44157 = v_44059 & v_44156;
assign v_44158 = v_44012 & v_44154;
assign v_44160 = v_44010 & v_44159;
assign v_44162 = v_44065 & v_44161;
assign v_44163 = v_44009 & v_44159;
assign v_44165 = v_44007 & v_44164;
assign v_44167 = v_44071 & v_44166;
assign v_44168 = v_44006 & v_44164;
assign v_44170 = v_44004 & v_44169;
assign v_44172 = v_44077 & v_44171;
assign v_44173 = v_44003 & v_44169;
assign v_44175 = v_44001 & v_44174;
assign v_44177 = v_44083 & v_44176;
assign v_44178 = v_44000 & v_44174;
assign v_44180 = v_43998 & v_44179;
assign v_44182 = v_44089 & v_44181;
assign v_44183 = v_43997 & v_44179;
assign v_44185 = v_43995 & v_44184;
assign v_44187 = v_44095 & v_44186;
assign v_44188 = v_43994 & v_44184;
assign v_44190 = v_43992 & v_44189;
assign v_44192 = v_44101 & v_44191;
assign v_44193 = v_43991 & v_44189;
assign v_44195 = v_43989 & v_44194;
assign v_44197 = v_44107 & v_44196;
assign v_44198 = v_43988 & v_44194;
assign v_44200 = v_43986 & v_44199;
assign v_44202 = v_44113 & v_44201;
assign v_44203 = v_43985 & v_44199;
assign v_44205 = v_43983 & v_44204;
assign v_44207 = v_44119 & v_44206;
assign v_44208 = v_43982 & v_44204;
assign v_44210 = v_43980 & v_44209;
assign v_44212 = v_44125 & v_44211;
assign v_44213 = v_43979 & v_44209;
assign v_44215 = v_44214;
assign v_44217 = v_44129 & v_44216;
assign v_44218 = v_44217;
assign v_44220 = v_44219;
assign v_44222 = ~v_2623;
assign v_44223 = ~v_41776;
assign v_44224 = v_41776;
assign v_44225 = ~v_2627;
assign v_44226 = ~v_41780;
assign v_44227 = v_41780;
assign v_44228 = ~v_2631;
assign v_44229 = ~v_41784;
assign v_44230 = v_41784;
assign v_44231 = ~v_2635;
assign v_44232 = ~v_41788;
assign v_44233 = v_41788;
assign v_44234 = ~v_41791;
assign v_44235 = ~v_2640;
assign v_44236 = v_2640;
assign v_44237 = ~v_41795;
assign v_44238 = ~v_2644;
assign v_44239 = v_2644;
assign v_44240 = ~v_41799;
assign v_44241 = ~v_2648;
assign v_44242 = v_2648;
assign v_44243 = ~v_41803;
assign v_44244 = ~v_2652;
assign v_44245 = v_2652;
assign v_44246 = ~v_41807;
assign v_44247 = ~v_2656;
assign v_44248 = v_2656;
assign v_44249 = ~v_41811;
assign v_44250 = ~v_2660;
assign v_44251 = v_2660;
assign v_44252 = ~v_41815;
assign v_44253 = ~v_2664;
assign v_44254 = v_2664;
assign v_44255 = ~v_41819;
assign v_44256 = ~v_2668;
assign v_44257 = v_2668;
assign v_44258 = ~v_41823;
assign v_44259 = ~v_2672;
assign v_44260 = v_2672;
assign v_44261 = ~v_41827;
assign v_44262 = ~v_2676;
assign v_44263 = v_2676;
assign v_44264 = ~v_41831;
assign v_44265 = ~v_2680;
assign v_44266 = v_2680;
assign v_44267 = ~v_41835;
assign v_44268 = ~v_2684;
assign v_44269 = v_2684;
assign v_44270 = ~v_41839;
assign v_44271 = ~v_2688;
assign v_44272 = v_44271;
assign v_44274 = v_44273;
assign v_44276 = v_44268 & v_44275;
assign v_44278 = v_41835;
assign v_44280 = v_44277 & v_44279;
assign v_44282 = v_44265 & v_44281;
assign v_44284 = v_41831;
assign v_44286 = v_44283 & v_44285;
assign v_44288 = v_44262 & v_44287;
assign v_44290 = v_41827;
assign v_44292 = v_44289 & v_44291;
assign v_44294 = v_44259 & v_44293;
assign v_44296 = v_41823;
assign v_44298 = v_44295 & v_44297;
assign v_44300 = v_44256 & v_44299;
assign v_44302 = v_41819;
assign v_44304 = v_44301 & v_44303;
assign v_44306 = v_44253 & v_44305;
assign v_44308 = v_41815;
assign v_44310 = v_44307 & v_44309;
assign v_44312 = v_44250 & v_44311;
assign v_44314 = v_41811;
assign v_44316 = v_44313 & v_44315;
assign v_44318 = v_44247 & v_44317;
assign v_44320 = v_41807;
assign v_44322 = v_44319 & v_44321;
assign v_44324 = v_44244 & v_44323;
assign v_44326 = v_41803;
assign v_44328 = v_44325 & v_44327;
assign v_44330 = v_44241 & v_44329;
assign v_44332 = v_41799;
assign v_44334 = v_44331 & v_44333;
assign v_44336 = v_44238 & v_44335;
assign v_44338 = v_41795;
assign v_44340 = v_44337 & v_44339;
assign v_44342 = v_44235 & v_44341;
assign v_44344 = v_41791;
assign v_44346 = v_44343 & v_44345;
assign v_44348 = v_44232 & v_44347;
assign v_44350 = v_2635;
assign v_44352 = v_44349 & v_44351;
assign v_44354 = v_44229 & v_44353;
assign v_44356 = v_2631;
assign v_44358 = v_44355 & v_44357;
assign v_44360 = v_44226 & v_44359;
assign v_44362 = v_2627;
assign v_44364 = v_44361 & v_44363;
assign v_44366 = v_44223 & v_44365;
assign v_44368 = v_2623;
assign v_44370 = v_44367 & v_44369;
assign v_44371 = v_44370;
assign v_44373 = v_41839;
assign v_44374 = v_2688;
assign v_44375 = v_44374;
assign v_44376 = v_44373 & v_44375;
assign v_44377 = v_44376;
assign v_44378 = v_44268 & v_44377;
assign v_44380 = v_44278 & v_44379;
assign v_44381 = v_44267 & v_44377;
assign v_44383 = v_44265 & v_44382;
assign v_44385 = v_44284 & v_44384;
assign v_44386 = v_44264 & v_44382;
assign v_44388 = v_44262 & v_44387;
assign v_44390 = v_44290 & v_44389;
assign v_44391 = v_44261 & v_44387;
assign v_44393 = v_44259 & v_44392;
assign v_44395 = v_44296 & v_44394;
assign v_44396 = v_44258 & v_44392;
assign v_44398 = v_44256 & v_44397;
assign v_44400 = v_44302 & v_44399;
assign v_44401 = v_44255 & v_44397;
assign v_44403 = v_44253 & v_44402;
assign v_44405 = v_44308 & v_44404;
assign v_44406 = v_44252 & v_44402;
assign v_44408 = v_44250 & v_44407;
assign v_44410 = v_44314 & v_44409;
assign v_44411 = v_44249 & v_44407;
assign v_44413 = v_44247 & v_44412;
assign v_44415 = v_44320 & v_44414;
assign v_44416 = v_44246 & v_44412;
assign v_44418 = v_44244 & v_44417;
assign v_44420 = v_44326 & v_44419;
assign v_44421 = v_44243 & v_44417;
assign v_44423 = v_44241 & v_44422;
assign v_44425 = v_44332 & v_44424;
assign v_44426 = v_44240 & v_44422;
assign v_44428 = v_44238 & v_44427;
assign v_44430 = v_44338 & v_44429;
assign v_44431 = v_44237 & v_44427;
assign v_44433 = v_44235 & v_44432;
assign v_44435 = v_44344 & v_44434;
assign v_44436 = v_44234 & v_44432;
assign v_44438 = v_44232 & v_44437;
assign v_44440 = v_44350 & v_44439;
assign v_44441 = v_44231 & v_44437;
assign v_44443 = v_44229 & v_44442;
assign v_44445 = v_44356 & v_44444;
assign v_44446 = v_44228 & v_44442;
assign v_44448 = v_44226 & v_44447;
assign v_44450 = v_44362 & v_44449;
assign v_44451 = v_44225 & v_44447;
assign v_44453 = v_44223 & v_44452;
assign v_44455 = v_44368 & v_44454;
assign v_44456 = v_44222 & v_44452;
assign v_44458 = v_44457;
assign v_44460 = v_44372 & v_44459;
assign v_44461 = v_44460;
assign v_44463 = v_44462;
assign v_44465 = ~v_2883;
assign v_44466 = ~v_41776;
assign v_44467 = v_41776;
assign v_44468 = ~v_2887;
assign v_44469 = ~v_41780;
assign v_44470 = v_41780;
assign v_44471 = ~v_2891;
assign v_44472 = ~v_41784;
assign v_44473 = v_41784;
assign v_44474 = ~v_2895;
assign v_44475 = ~v_41788;
assign v_44476 = v_41788;
assign v_44477 = ~v_41791;
assign v_44478 = ~v_2900;
assign v_44479 = v_2900;
assign v_44480 = ~v_41795;
assign v_44481 = ~v_2904;
assign v_44482 = v_2904;
assign v_44483 = ~v_41799;
assign v_44484 = ~v_2908;
assign v_44485 = v_2908;
assign v_44486 = ~v_41803;
assign v_44487 = ~v_2912;
assign v_44488 = v_2912;
assign v_44489 = ~v_41807;
assign v_44490 = ~v_2916;
assign v_44491 = v_2916;
assign v_44492 = ~v_41811;
assign v_44493 = ~v_2920;
assign v_44494 = v_2920;
assign v_44495 = ~v_41815;
assign v_44496 = ~v_2924;
assign v_44497 = v_2924;
assign v_44498 = ~v_41819;
assign v_44499 = ~v_2928;
assign v_44500 = v_2928;
assign v_44501 = ~v_41823;
assign v_44502 = ~v_2932;
assign v_44503 = v_2932;
assign v_44504 = ~v_41827;
assign v_44505 = ~v_2936;
assign v_44506 = v_2936;
assign v_44507 = ~v_41831;
assign v_44508 = ~v_2940;
assign v_44509 = v_2940;
assign v_44510 = ~v_41835;
assign v_44511 = ~v_2944;
assign v_44512 = v_2944;
assign v_44513 = ~v_41839;
assign v_44514 = ~v_2948;
assign v_44515 = v_44514;
assign v_44517 = v_44516;
assign v_44519 = v_44511 & v_44518;
assign v_44521 = v_41835;
assign v_44523 = v_44520 & v_44522;
assign v_44525 = v_44508 & v_44524;
assign v_44527 = v_41831;
assign v_44529 = v_44526 & v_44528;
assign v_44531 = v_44505 & v_44530;
assign v_44533 = v_41827;
assign v_44535 = v_44532 & v_44534;
assign v_44537 = v_44502 & v_44536;
assign v_44539 = v_41823;
assign v_44541 = v_44538 & v_44540;
assign v_44543 = v_44499 & v_44542;
assign v_44545 = v_41819;
assign v_44547 = v_44544 & v_44546;
assign v_44549 = v_44496 & v_44548;
assign v_44551 = v_41815;
assign v_44553 = v_44550 & v_44552;
assign v_44555 = v_44493 & v_44554;
assign v_44557 = v_41811;
assign v_44559 = v_44556 & v_44558;
assign v_44561 = v_44490 & v_44560;
assign v_44563 = v_41807;
assign v_44565 = v_44562 & v_44564;
assign v_44567 = v_44487 & v_44566;
assign v_44569 = v_41803;
assign v_44571 = v_44568 & v_44570;
assign v_44573 = v_44484 & v_44572;
assign v_44575 = v_41799;
assign v_44577 = v_44574 & v_44576;
assign v_44579 = v_44481 & v_44578;
assign v_44581 = v_41795;
assign v_44583 = v_44580 & v_44582;
assign v_44585 = v_44478 & v_44584;
assign v_44587 = v_41791;
assign v_44589 = v_44586 & v_44588;
assign v_44591 = v_44475 & v_44590;
assign v_44593 = v_2895;
assign v_44595 = v_44592 & v_44594;
assign v_44597 = v_44472 & v_44596;
assign v_44599 = v_2891;
assign v_44601 = v_44598 & v_44600;
assign v_44603 = v_44469 & v_44602;
assign v_44605 = v_2887;
assign v_44607 = v_44604 & v_44606;
assign v_44609 = v_44466 & v_44608;
assign v_44611 = v_2883;
assign v_44613 = v_44610 & v_44612;
assign v_44614 = v_44613;
assign v_44616 = v_41839;
assign v_44617 = v_2948;
assign v_44618 = v_44617;
assign v_44619 = v_44616 & v_44618;
assign v_44620 = v_44619;
assign v_44621 = v_44511 & v_44620;
assign v_44623 = v_44521 & v_44622;
assign v_44624 = v_44510 & v_44620;
assign v_44626 = v_44508 & v_44625;
assign v_44628 = v_44527 & v_44627;
assign v_44629 = v_44507 & v_44625;
assign v_44631 = v_44505 & v_44630;
assign v_44633 = v_44533 & v_44632;
assign v_44634 = v_44504 & v_44630;
assign v_44636 = v_44502 & v_44635;
assign v_44638 = v_44539 & v_44637;
assign v_44639 = v_44501 & v_44635;
assign v_44641 = v_44499 & v_44640;
assign v_44643 = v_44545 & v_44642;
assign v_44644 = v_44498 & v_44640;
assign v_44646 = v_44496 & v_44645;
assign v_44648 = v_44551 & v_44647;
assign v_44649 = v_44495 & v_44645;
assign v_44651 = v_44493 & v_44650;
assign v_44653 = v_44557 & v_44652;
assign v_44654 = v_44492 & v_44650;
assign v_44656 = v_44490 & v_44655;
assign v_44658 = v_44563 & v_44657;
assign v_44659 = v_44489 & v_44655;
assign v_44661 = v_44487 & v_44660;
assign v_44663 = v_44569 & v_44662;
assign v_44664 = v_44486 & v_44660;
assign v_44666 = v_44484 & v_44665;
assign v_44668 = v_44575 & v_44667;
assign v_44669 = v_44483 & v_44665;
assign v_44671 = v_44481 & v_44670;
assign v_44673 = v_44581 & v_44672;
assign v_44674 = v_44480 & v_44670;
assign v_44676 = v_44478 & v_44675;
assign v_44678 = v_44587 & v_44677;
assign v_44679 = v_44477 & v_44675;
assign v_44681 = v_44475 & v_44680;
assign v_44683 = v_44593 & v_44682;
assign v_44684 = v_44474 & v_44680;
assign v_44686 = v_44472 & v_44685;
assign v_44688 = v_44599 & v_44687;
assign v_44689 = v_44471 & v_44685;
assign v_44691 = v_44469 & v_44690;
assign v_44693 = v_44605 & v_44692;
assign v_44694 = v_44468 & v_44690;
assign v_44696 = v_44466 & v_44695;
assign v_44698 = v_44611 & v_44697;
assign v_44699 = v_44465 & v_44695;
assign v_44701 = v_44700;
assign v_44703 = v_44615 & v_44702;
assign v_44704 = v_44703;
assign v_44706 = v_44705;
assign v_44708 = ~v_3143;
assign v_44709 = ~v_41776;
assign v_44710 = v_41776;
assign v_44711 = ~v_3147;
assign v_44712 = ~v_41780;
assign v_44713 = v_41780;
assign v_44714 = ~v_3151;
assign v_44715 = ~v_41784;
assign v_44716 = v_41784;
assign v_44717 = ~v_3155;
assign v_44718 = ~v_41788;
assign v_44719 = v_41788;
assign v_44720 = ~v_41791;
assign v_44721 = ~v_3160;
assign v_44722 = v_3160;
assign v_44723 = ~v_41795;
assign v_44724 = ~v_3164;
assign v_44725 = v_3164;
assign v_44726 = ~v_41799;
assign v_44727 = ~v_3168;
assign v_44728 = v_3168;
assign v_44729 = ~v_41803;
assign v_44730 = ~v_3172;
assign v_44731 = v_3172;
assign v_44732 = ~v_41807;
assign v_44733 = ~v_3176;
assign v_44734 = v_3176;
assign v_44735 = ~v_41811;
assign v_44736 = ~v_3180;
assign v_44737 = v_3180;
assign v_44738 = ~v_41815;
assign v_44739 = ~v_3184;
assign v_44740 = v_3184;
assign v_44741 = ~v_41819;
assign v_44742 = ~v_3188;
assign v_44743 = v_3188;
assign v_44744 = ~v_41823;
assign v_44745 = ~v_3192;
assign v_44746 = v_3192;
assign v_44747 = ~v_41827;
assign v_44748 = ~v_3196;
assign v_44749 = v_3196;
assign v_44750 = ~v_41831;
assign v_44751 = ~v_3200;
assign v_44752 = v_3200;
assign v_44753 = ~v_41835;
assign v_44754 = ~v_3204;
assign v_44755 = v_3204;
assign v_44756 = ~v_41839;
assign v_44757 = ~v_3208;
assign v_44758 = v_44757;
assign v_44760 = v_44759;
assign v_44762 = v_44754 & v_44761;
assign v_44764 = v_41835;
assign v_44766 = v_44763 & v_44765;
assign v_44768 = v_44751 & v_44767;
assign v_44770 = v_41831;
assign v_44772 = v_44769 & v_44771;
assign v_44774 = v_44748 & v_44773;
assign v_44776 = v_41827;
assign v_44778 = v_44775 & v_44777;
assign v_44780 = v_44745 & v_44779;
assign v_44782 = v_41823;
assign v_44784 = v_44781 & v_44783;
assign v_44786 = v_44742 & v_44785;
assign v_44788 = v_41819;
assign v_44790 = v_44787 & v_44789;
assign v_44792 = v_44739 & v_44791;
assign v_44794 = v_41815;
assign v_44796 = v_44793 & v_44795;
assign v_44798 = v_44736 & v_44797;
assign v_44800 = v_41811;
assign v_44802 = v_44799 & v_44801;
assign v_44804 = v_44733 & v_44803;
assign v_44806 = v_41807;
assign v_44808 = v_44805 & v_44807;
assign v_44810 = v_44730 & v_44809;
assign v_44812 = v_41803;
assign v_44814 = v_44811 & v_44813;
assign v_44816 = v_44727 & v_44815;
assign v_44818 = v_41799;
assign v_44820 = v_44817 & v_44819;
assign v_44822 = v_44724 & v_44821;
assign v_44824 = v_41795;
assign v_44826 = v_44823 & v_44825;
assign v_44828 = v_44721 & v_44827;
assign v_44830 = v_41791;
assign v_44832 = v_44829 & v_44831;
assign v_44834 = v_44718 & v_44833;
assign v_44836 = v_3155;
assign v_44838 = v_44835 & v_44837;
assign v_44840 = v_44715 & v_44839;
assign v_44842 = v_3151;
assign v_44844 = v_44841 & v_44843;
assign v_44846 = v_44712 & v_44845;
assign v_44848 = v_3147;
assign v_44850 = v_44847 & v_44849;
assign v_44852 = v_44709 & v_44851;
assign v_44854 = v_3143;
assign v_44856 = v_44853 & v_44855;
assign v_44857 = v_44856;
assign v_44859 = v_41839;
assign v_44860 = v_3208;
assign v_44861 = v_44860;
assign v_44862 = v_44859 & v_44861;
assign v_44863 = v_44862;
assign v_44864 = v_44754 & v_44863;
assign v_44866 = v_44764 & v_44865;
assign v_44867 = v_44753 & v_44863;
assign v_44869 = v_44751 & v_44868;
assign v_44871 = v_44770 & v_44870;
assign v_44872 = v_44750 & v_44868;
assign v_44874 = v_44748 & v_44873;
assign v_44876 = v_44776 & v_44875;
assign v_44877 = v_44747 & v_44873;
assign v_44879 = v_44745 & v_44878;
assign v_44881 = v_44782 & v_44880;
assign v_44882 = v_44744 & v_44878;
assign v_44884 = v_44742 & v_44883;
assign v_44886 = v_44788 & v_44885;
assign v_44887 = v_44741 & v_44883;
assign v_44889 = v_44739 & v_44888;
assign v_44891 = v_44794 & v_44890;
assign v_44892 = v_44738 & v_44888;
assign v_44894 = v_44736 & v_44893;
assign v_44896 = v_44800 & v_44895;
assign v_44897 = v_44735 & v_44893;
assign v_44899 = v_44733 & v_44898;
assign v_44901 = v_44806 & v_44900;
assign v_44902 = v_44732 & v_44898;
assign v_44904 = v_44730 & v_44903;
assign v_44906 = v_44812 & v_44905;
assign v_44907 = v_44729 & v_44903;
assign v_44909 = v_44727 & v_44908;
assign v_44911 = v_44818 & v_44910;
assign v_44912 = v_44726 & v_44908;
assign v_44914 = v_44724 & v_44913;
assign v_44916 = v_44824 & v_44915;
assign v_44917 = v_44723 & v_44913;
assign v_44919 = v_44721 & v_44918;
assign v_44921 = v_44830 & v_44920;
assign v_44922 = v_44720 & v_44918;
assign v_44924 = v_44718 & v_44923;
assign v_44926 = v_44836 & v_44925;
assign v_44927 = v_44717 & v_44923;
assign v_44929 = v_44715 & v_44928;
assign v_44931 = v_44842 & v_44930;
assign v_44932 = v_44714 & v_44928;
assign v_44934 = v_44712 & v_44933;
assign v_44936 = v_44848 & v_44935;
assign v_44937 = v_44711 & v_44933;
assign v_44939 = v_44709 & v_44938;
assign v_44941 = v_44854 & v_44940;
assign v_44942 = v_44708 & v_44938;
assign v_44944 = v_44943;
assign v_44946 = v_44858 & v_44945;
assign v_44947 = v_44946;
assign v_44949 = v_44948;
assign v_44951 = ~v_3403;
assign v_44952 = ~v_41776;
assign v_44953 = v_41776;
assign v_44954 = ~v_3407;
assign v_44955 = ~v_41780;
assign v_44956 = v_41780;
assign v_44957 = ~v_3411;
assign v_44958 = ~v_41784;
assign v_44959 = v_41784;
assign v_44960 = ~v_3415;
assign v_44961 = ~v_41788;
assign v_44962 = v_41788;
assign v_44963 = ~v_41791;
assign v_44964 = ~v_3420;
assign v_44965 = v_3420;
assign v_44966 = ~v_41795;
assign v_44967 = ~v_3424;
assign v_44968 = v_3424;
assign v_44969 = ~v_41799;
assign v_44970 = ~v_3428;
assign v_44971 = v_3428;
assign v_44972 = ~v_41803;
assign v_44973 = ~v_3432;
assign v_44974 = v_3432;
assign v_44975 = ~v_41807;
assign v_44976 = ~v_3436;
assign v_44977 = v_3436;
assign v_44978 = ~v_41811;
assign v_44979 = ~v_3440;
assign v_44980 = v_3440;
assign v_44981 = ~v_41815;
assign v_44982 = ~v_3444;
assign v_44983 = v_3444;
assign v_44984 = ~v_41819;
assign v_44985 = ~v_3448;
assign v_44986 = v_3448;
assign v_44987 = ~v_41823;
assign v_44988 = ~v_3452;
assign v_44989 = v_3452;
assign v_44990 = ~v_41827;
assign v_44991 = ~v_3456;
assign v_44992 = v_3456;
assign v_44993 = ~v_41831;
assign v_44994 = ~v_3460;
assign v_44995 = v_3460;
assign v_44996 = ~v_41835;
assign v_44997 = ~v_3464;
assign v_44998 = v_3464;
assign v_44999 = ~v_41839;
assign v_45000 = ~v_3468;
assign v_45001 = v_45000;
assign v_45003 = v_45002;
assign v_45005 = v_44997 & v_45004;
assign v_45007 = v_41835;
assign v_45009 = v_45006 & v_45008;
assign v_45011 = v_44994 & v_45010;
assign v_45013 = v_41831;
assign v_45015 = v_45012 & v_45014;
assign v_45017 = v_44991 & v_45016;
assign v_45019 = v_41827;
assign v_45021 = v_45018 & v_45020;
assign v_45023 = v_44988 & v_45022;
assign v_45025 = v_41823;
assign v_45027 = v_45024 & v_45026;
assign v_45029 = v_44985 & v_45028;
assign v_45031 = v_41819;
assign v_45033 = v_45030 & v_45032;
assign v_45035 = v_44982 & v_45034;
assign v_45037 = v_41815;
assign v_45039 = v_45036 & v_45038;
assign v_45041 = v_44979 & v_45040;
assign v_45043 = v_41811;
assign v_45045 = v_45042 & v_45044;
assign v_45047 = v_44976 & v_45046;
assign v_45049 = v_41807;
assign v_45051 = v_45048 & v_45050;
assign v_45053 = v_44973 & v_45052;
assign v_45055 = v_41803;
assign v_45057 = v_45054 & v_45056;
assign v_45059 = v_44970 & v_45058;
assign v_45061 = v_41799;
assign v_45063 = v_45060 & v_45062;
assign v_45065 = v_44967 & v_45064;
assign v_45067 = v_41795;
assign v_45069 = v_45066 & v_45068;
assign v_45071 = v_44964 & v_45070;
assign v_45073 = v_41791;
assign v_45075 = v_45072 & v_45074;
assign v_45077 = v_44961 & v_45076;
assign v_45079 = v_3415;
assign v_45081 = v_45078 & v_45080;
assign v_45083 = v_44958 & v_45082;
assign v_45085 = v_3411;
assign v_45087 = v_45084 & v_45086;
assign v_45089 = v_44955 & v_45088;
assign v_45091 = v_3407;
assign v_45093 = v_45090 & v_45092;
assign v_45095 = v_44952 & v_45094;
assign v_45097 = v_3403;
assign v_45099 = v_45096 & v_45098;
assign v_45100 = v_45099;
assign v_45102 = v_41839;
assign v_45103 = v_3468;
assign v_45104 = v_45103;
assign v_45105 = v_45102 & v_45104;
assign v_45106 = v_45105;
assign v_45107 = v_44997 & v_45106;
assign v_45109 = v_45007 & v_45108;
assign v_45110 = v_44996 & v_45106;
assign v_45112 = v_44994 & v_45111;
assign v_45114 = v_45013 & v_45113;
assign v_45115 = v_44993 & v_45111;
assign v_45117 = v_44991 & v_45116;
assign v_45119 = v_45019 & v_45118;
assign v_45120 = v_44990 & v_45116;
assign v_45122 = v_44988 & v_45121;
assign v_45124 = v_45025 & v_45123;
assign v_45125 = v_44987 & v_45121;
assign v_45127 = v_44985 & v_45126;
assign v_45129 = v_45031 & v_45128;
assign v_45130 = v_44984 & v_45126;
assign v_45132 = v_44982 & v_45131;
assign v_45134 = v_45037 & v_45133;
assign v_45135 = v_44981 & v_45131;
assign v_45137 = v_44979 & v_45136;
assign v_45139 = v_45043 & v_45138;
assign v_45140 = v_44978 & v_45136;
assign v_45142 = v_44976 & v_45141;
assign v_45144 = v_45049 & v_45143;
assign v_45145 = v_44975 & v_45141;
assign v_45147 = v_44973 & v_45146;
assign v_45149 = v_45055 & v_45148;
assign v_45150 = v_44972 & v_45146;
assign v_45152 = v_44970 & v_45151;
assign v_45154 = v_45061 & v_45153;
assign v_45155 = v_44969 & v_45151;
assign v_45157 = v_44967 & v_45156;
assign v_45159 = v_45067 & v_45158;
assign v_45160 = v_44966 & v_45156;
assign v_45162 = v_44964 & v_45161;
assign v_45164 = v_45073 & v_45163;
assign v_45165 = v_44963 & v_45161;
assign v_45167 = v_44961 & v_45166;
assign v_45169 = v_45079 & v_45168;
assign v_45170 = v_44960 & v_45166;
assign v_45172 = v_44958 & v_45171;
assign v_45174 = v_45085 & v_45173;
assign v_45175 = v_44957 & v_45171;
assign v_45177 = v_44955 & v_45176;
assign v_45179 = v_45091 & v_45178;
assign v_45180 = v_44954 & v_45176;
assign v_45182 = v_44952 & v_45181;
assign v_45184 = v_45097 & v_45183;
assign v_45185 = v_44951 & v_45181;
assign v_45187 = v_45186;
assign v_45189 = v_45101 & v_45188;
assign v_45190 = v_45189;
assign v_45192 = v_45191;
assign v_45194 = ~v_3663;
assign v_45195 = ~v_41776;
assign v_45196 = v_41776;
assign v_45197 = ~v_3667;
assign v_45198 = ~v_41780;
assign v_45199 = v_41780;
assign v_45200 = ~v_3671;
assign v_45201 = ~v_41784;
assign v_45202 = v_41784;
assign v_45203 = ~v_3675;
assign v_45204 = ~v_41788;
assign v_45205 = v_41788;
assign v_45206 = ~v_41791;
assign v_45207 = ~v_3680;
assign v_45208 = v_3680;
assign v_45209 = ~v_41795;
assign v_45210 = ~v_3684;
assign v_45211 = v_3684;
assign v_45212 = ~v_41799;
assign v_45213 = ~v_3688;
assign v_45214 = v_3688;
assign v_45215 = ~v_41803;
assign v_45216 = ~v_3692;
assign v_45217 = v_3692;
assign v_45218 = ~v_41807;
assign v_45219 = ~v_3696;
assign v_45220 = v_3696;
assign v_45221 = ~v_41811;
assign v_45222 = ~v_3700;
assign v_45223 = v_3700;
assign v_45224 = ~v_41815;
assign v_45225 = ~v_3704;
assign v_45226 = v_3704;
assign v_45227 = ~v_41819;
assign v_45228 = ~v_3708;
assign v_45229 = v_3708;
assign v_45230 = ~v_41823;
assign v_45231 = ~v_3712;
assign v_45232 = v_3712;
assign v_45233 = ~v_41827;
assign v_45234 = ~v_3716;
assign v_45235 = v_3716;
assign v_45236 = ~v_41831;
assign v_45237 = ~v_3720;
assign v_45238 = v_3720;
assign v_45239 = ~v_41835;
assign v_45240 = ~v_3724;
assign v_45241 = v_3724;
assign v_45242 = ~v_41839;
assign v_45243 = ~v_3728;
assign v_45244 = v_45243;
assign v_45246 = v_45245;
assign v_45248 = v_45240 & v_45247;
assign v_45250 = v_41835;
assign v_45252 = v_45249 & v_45251;
assign v_45254 = v_45237 & v_45253;
assign v_45256 = v_41831;
assign v_45258 = v_45255 & v_45257;
assign v_45260 = v_45234 & v_45259;
assign v_45262 = v_41827;
assign v_45264 = v_45261 & v_45263;
assign v_45266 = v_45231 & v_45265;
assign v_45268 = v_41823;
assign v_45270 = v_45267 & v_45269;
assign v_45272 = v_45228 & v_45271;
assign v_45274 = v_41819;
assign v_45276 = v_45273 & v_45275;
assign v_45278 = v_45225 & v_45277;
assign v_45280 = v_41815;
assign v_45282 = v_45279 & v_45281;
assign v_45284 = v_45222 & v_45283;
assign v_45286 = v_41811;
assign v_45288 = v_45285 & v_45287;
assign v_45290 = v_45219 & v_45289;
assign v_45292 = v_41807;
assign v_45294 = v_45291 & v_45293;
assign v_45296 = v_45216 & v_45295;
assign v_45298 = v_41803;
assign v_45300 = v_45297 & v_45299;
assign v_45302 = v_45213 & v_45301;
assign v_45304 = v_41799;
assign v_45306 = v_45303 & v_45305;
assign v_45308 = v_45210 & v_45307;
assign v_45310 = v_41795;
assign v_45312 = v_45309 & v_45311;
assign v_45314 = v_45207 & v_45313;
assign v_45316 = v_41791;
assign v_45318 = v_45315 & v_45317;
assign v_45320 = v_45204 & v_45319;
assign v_45322 = v_3675;
assign v_45324 = v_45321 & v_45323;
assign v_45326 = v_45201 & v_45325;
assign v_45328 = v_3671;
assign v_45330 = v_45327 & v_45329;
assign v_45332 = v_45198 & v_45331;
assign v_45334 = v_3667;
assign v_45336 = v_45333 & v_45335;
assign v_45338 = v_45195 & v_45337;
assign v_45340 = v_3663;
assign v_45342 = v_45339 & v_45341;
assign v_45343 = v_45342;
assign v_45345 = v_41839;
assign v_45346 = v_3728;
assign v_45347 = v_45346;
assign v_45348 = v_45345 & v_45347;
assign v_45349 = v_45348;
assign v_45350 = v_45240 & v_45349;
assign v_45352 = v_45250 & v_45351;
assign v_45353 = v_45239 & v_45349;
assign v_45355 = v_45237 & v_45354;
assign v_45357 = v_45256 & v_45356;
assign v_45358 = v_45236 & v_45354;
assign v_45360 = v_45234 & v_45359;
assign v_45362 = v_45262 & v_45361;
assign v_45363 = v_45233 & v_45359;
assign v_45365 = v_45231 & v_45364;
assign v_45367 = v_45268 & v_45366;
assign v_45368 = v_45230 & v_45364;
assign v_45370 = v_45228 & v_45369;
assign v_45372 = v_45274 & v_45371;
assign v_45373 = v_45227 & v_45369;
assign v_45375 = v_45225 & v_45374;
assign v_45377 = v_45280 & v_45376;
assign v_45378 = v_45224 & v_45374;
assign v_45380 = v_45222 & v_45379;
assign v_45382 = v_45286 & v_45381;
assign v_45383 = v_45221 & v_45379;
assign v_45385 = v_45219 & v_45384;
assign v_45387 = v_45292 & v_45386;
assign v_45388 = v_45218 & v_45384;
assign v_45390 = v_45216 & v_45389;
assign v_45392 = v_45298 & v_45391;
assign v_45393 = v_45215 & v_45389;
assign v_45395 = v_45213 & v_45394;
assign v_45397 = v_45304 & v_45396;
assign v_45398 = v_45212 & v_45394;
assign v_45400 = v_45210 & v_45399;
assign v_45402 = v_45310 & v_45401;
assign v_45403 = v_45209 & v_45399;
assign v_45405 = v_45207 & v_45404;
assign v_45407 = v_45316 & v_45406;
assign v_45408 = v_45206 & v_45404;
assign v_45410 = v_45204 & v_45409;
assign v_45412 = v_45322 & v_45411;
assign v_45413 = v_45203 & v_45409;
assign v_45415 = v_45201 & v_45414;
assign v_45417 = v_45328 & v_45416;
assign v_45418 = v_45200 & v_45414;
assign v_45420 = v_45198 & v_45419;
assign v_45422 = v_45334 & v_45421;
assign v_45423 = v_45197 & v_45419;
assign v_45425 = v_45195 & v_45424;
assign v_45427 = v_45340 & v_45426;
assign v_45428 = v_45194 & v_45424;
assign v_45430 = v_45429;
assign v_45432 = v_45344 & v_45431;
assign v_45433 = v_45432;
assign v_45435 = v_45434;
assign v_45437 = ~v_3923;
assign v_45438 = ~v_41776;
assign v_45439 = v_41776;
assign v_45440 = ~v_3927;
assign v_45441 = ~v_41780;
assign v_45442 = v_41780;
assign v_45443 = ~v_3931;
assign v_45444 = ~v_41784;
assign v_45445 = v_41784;
assign v_45446 = ~v_3935;
assign v_45447 = ~v_41788;
assign v_45448 = v_41788;
assign v_45449 = ~v_41791;
assign v_45450 = ~v_3940;
assign v_45451 = v_3940;
assign v_45452 = ~v_41795;
assign v_45453 = ~v_3944;
assign v_45454 = v_3944;
assign v_45455 = ~v_41799;
assign v_45456 = ~v_3948;
assign v_45457 = v_3948;
assign v_45458 = ~v_41803;
assign v_45459 = ~v_3952;
assign v_45460 = v_3952;
assign v_45461 = ~v_41807;
assign v_45462 = ~v_3956;
assign v_45463 = v_3956;
assign v_45464 = ~v_41811;
assign v_45465 = ~v_3960;
assign v_45466 = v_3960;
assign v_45467 = ~v_41815;
assign v_45468 = ~v_3964;
assign v_45469 = v_3964;
assign v_45470 = ~v_41819;
assign v_45471 = ~v_3968;
assign v_45472 = v_3968;
assign v_45473 = ~v_41823;
assign v_45474 = ~v_3972;
assign v_45475 = v_3972;
assign v_45476 = ~v_41827;
assign v_45477 = ~v_3976;
assign v_45478 = v_3976;
assign v_45479 = ~v_41831;
assign v_45480 = ~v_3980;
assign v_45481 = v_3980;
assign v_45482 = ~v_41835;
assign v_45483 = ~v_3984;
assign v_45484 = v_3984;
assign v_45485 = ~v_41839;
assign v_45486 = ~v_3988;
assign v_45487 = v_45486;
assign v_45489 = v_45488;
assign v_45491 = v_45483 & v_45490;
assign v_45493 = v_41835;
assign v_45495 = v_45492 & v_45494;
assign v_45497 = v_45480 & v_45496;
assign v_45499 = v_41831;
assign v_45501 = v_45498 & v_45500;
assign v_45503 = v_45477 & v_45502;
assign v_45505 = v_41827;
assign v_45507 = v_45504 & v_45506;
assign v_45509 = v_45474 & v_45508;
assign v_45511 = v_41823;
assign v_45513 = v_45510 & v_45512;
assign v_45515 = v_45471 & v_45514;
assign v_45517 = v_41819;
assign v_45519 = v_45516 & v_45518;
assign v_45521 = v_45468 & v_45520;
assign v_45523 = v_41815;
assign v_45525 = v_45522 & v_45524;
assign v_45527 = v_45465 & v_45526;
assign v_45529 = v_41811;
assign v_45531 = v_45528 & v_45530;
assign v_45533 = v_45462 & v_45532;
assign v_45535 = v_41807;
assign v_45537 = v_45534 & v_45536;
assign v_45539 = v_45459 & v_45538;
assign v_45541 = v_41803;
assign v_45543 = v_45540 & v_45542;
assign v_45545 = v_45456 & v_45544;
assign v_45547 = v_41799;
assign v_45549 = v_45546 & v_45548;
assign v_45551 = v_45453 & v_45550;
assign v_45553 = v_41795;
assign v_45555 = v_45552 & v_45554;
assign v_45557 = v_45450 & v_45556;
assign v_45559 = v_41791;
assign v_45561 = v_45558 & v_45560;
assign v_45563 = v_45447 & v_45562;
assign v_45565 = v_3935;
assign v_45567 = v_45564 & v_45566;
assign v_45569 = v_45444 & v_45568;
assign v_45571 = v_3931;
assign v_45573 = v_45570 & v_45572;
assign v_45575 = v_45441 & v_45574;
assign v_45577 = v_3927;
assign v_45579 = v_45576 & v_45578;
assign v_45581 = v_45438 & v_45580;
assign v_45583 = v_3923;
assign v_45585 = v_45582 & v_45584;
assign v_45586 = v_45585;
assign v_45588 = v_41839;
assign v_45589 = v_3988;
assign v_45590 = v_45589;
assign v_45591 = v_45588 & v_45590;
assign v_45592 = v_45591;
assign v_45593 = v_45483 & v_45592;
assign v_45595 = v_45493 & v_45594;
assign v_45596 = v_45482 & v_45592;
assign v_45598 = v_45480 & v_45597;
assign v_45600 = v_45499 & v_45599;
assign v_45601 = v_45479 & v_45597;
assign v_45603 = v_45477 & v_45602;
assign v_45605 = v_45505 & v_45604;
assign v_45606 = v_45476 & v_45602;
assign v_45608 = v_45474 & v_45607;
assign v_45610 = v_45511 & v_45609;
assign v_45611 = v_45473 & v_45607;
assign v_45613 = v_45471 & v_45612;
assign v_45615 = v_45517 & v_45614;
assign v_45616 = v_45470 & v_45612;
assign v_45618 = v_45468 & v_45617;
assign v_45620 = v_45523 & v_45619;
assign v_45621 = v_45467 & v_45617;
assign v_45623 = v_45465 & v_45622;
assign v_45625 = v_45529 & v_45624;
assign v_45626 = v_45464 & v_45622;
assign v_45628 = v_45462 & v_45627;
assign v_45630 = v_45535 & v_45629;
assign v_45631 = v_45461 & v_45627;
assign v_45633 = v_45459 & v_45632;
assign v_45635 = v_45541 & v_45634;
assign v_45636 = v_45458 & v_45632;
assign v_45638 = v_45456 & v_45637;
assign v_45640 = v_45547 & v_45639;
assign v_45641 = v_45455 & v_45637;
assign v_45643 = v_45453 & v_45642;
assign v_45645 = v_45553 & v_45644;
assign v_45646 = v_45452 & v_45642;
assign v_45648 = v_45450 & v_45647;
assign v_45650 = v_45559 & v_45649;
assign v_45651 = v_45449 & v_45647;
assign v_45653 = v_45447 & v_45652;
assign v_45655 = v_45565 & v_45654;
assign v_45656 = v_45446 & v_45652;
assign v_45658 = v_45444 & v_45657;
assign v_45660 = v_45571 & v_45659;
assign v_45661 = v_45443 & v_45657;
assign v_45663 = v_45441 & v_45662;
assign v_45665 = v_45577 & v_45664;
assign v_45666 = v_45440 & v_45662;
assign v_45668 = v_45438 & v_45667;
assign v_45670 = v_45583 & v_45669;
assign v_45671 = v_45437 & v_45667;
assign v_45673 = v_45672;
assign v_45675 = v_45587 & v_45674;
assign v_45676 = v_45675;
assign v_45678 = v_45677;
assign v_45679 = ~v_4182;
assign v_45680 = ~v_41776;
assign v_45681 = v_41776;
assign v_45682 = ~v_4186;
assign v_45683 = ~v_41780;
assign v_45684 = v_41780;
assign v_45685 = ~v_4190;
assign v_45686 = ~v_41784;
assign v_45687 = v_41784;
assign v_45688 = ~v_4194;
assign v_45689 = ~v_41788;
assign v_45690 = v_41788;
assign v_45691 = ~v_41791;
assign v_45692 = ~v_4199;
assign v_45693 = v_4199;
assign v_45694 = ~v_41795;
assign v_45695 = ~v_4203;
assign v_45696 = v_4203;
assign v_45697 = ~v_41799;
assign v_45698 = ~v_4207;
assign v_45699 = v_4207;
assign v_45700 = ~v_41803;
assign v_45701 = ~v_4211;
assign v_45702 = v_4211;
assign v_45703 = ~v_41807;
assign v_45704 = ~v_4215;
assign v_45705 = v_4215;
assign v_45706 = ~v_41811;
assign v_45707 = ~v_4219;
assign v_45708 = v_4219;
assign v_45709 = ~v_41815;
assign v_45710 = ~v_4223;
assign v_45711 = v_4223;
assign v_45712 = ~v_41819;
assign v_45713 = ~v_4227;
assign v_45714 = v_4227;
assign v_45715 = ~v_41823;
assign v_45716 = ~v_4231;
assign v_45717 = v_4231;
assign v_45718 = ~v_41827;
assign v_45719 = ~v_4235;
assign v_45720 = v_4235;
assign v_45721 = ~v_41831;
assign v_45722 = ~v_4239;
assign v_45723 = v_4239;
assign v_45724 = ~v_41835;
assign v_45725 = ~v_4243;
assign v_45726 = v_4243;
assign v_45727 = ~v_41839;
assign v_45728 = ~v_4247;
assign v_45729 = v_45728;
assign v_45731 = v_45730;
assign v_45733 = v_45725 & v_45732;
assign v_45735 = v_41835;
assign v_45737 = v_45734 & v_45736;
assign v_45739 = v_45722 & v_45738;
assign v_45741 = v_41831;
assign v_45743 = v_45740 & v_45742;
assign v_45745 = v_45719 & v_45744;
assign v_45747 = v_41827;
assign v_45749 = v_45746 & v_45748;
assign v_45751 = v_45716 & v_45750;
assign v_45753 = v_41823;
assign v_45755 = v_45752 & v_45754;
assign v_45757 = v_45713 & v_45756;
assign v_45759 = v_41819;
assign v_45761 = v_45758 & v_45760;
assign v_45763 = v_45710 & v_45762;
assign v_45765 = v_41815;
assign v_45767 = v_45764 & v_45766;
assign v_45769 = v_45707 & v_45768;
assign v_45771 = v_41811;
assign v_45773 = v_45770 & v_45772;
assign v_45775 = v_45704 & v_45774;
assign v_45777 = v_41807;
assign v_45779 = v_45776 & v_45778;
assign v_45781 = v_45701 & v_45780;
assign v_45783 = v_41803;
assign v_45785 = v_45782 & v_45784;
assign v_45787 = v_45698 & v_45786;
assign v_45789 = v_41799;
assign v_45791 = v_45788 & v_45790;
assign v_45793 = v_45695 & v_45792;
assign v_45795 = v_41795;
assign v_45797 = v_45794 & v_45796;
assign v_45799 = v_45692 & v_45798;
assign v_45801 = v_41791;
assign v_45803 = v_45800 & v_45802;
assign v_45805 = v_45689 & v_45804;
assign v_45807 = v_4194;
assign v_45809 = v_45806 & v_45808;
assign v_45811 = v_45686 & v_45810;
assign v_45813 = v_4190;
assign v_45815 = v_45812 & v_45814;
assign v_45817 = v_45683 & v_45816;
assign v_45819 = v_4186;
assign v_45821 = v_45818 & v_45820;
assign v_45823 = v_45680 & v_45822;
assign v_45825 = v_4182;
assign v_45827 = v_45824 & v_45826;
assign v_45829 = ~v_45828;
assign v_45831 = v_41839;
assign v_45832 = v_4247;
assign v_45833 = v_45832;
assign v_45834 = v_45831 & v_45833;
assign v_45835 = v_45834;
assign v_45836 = v_45725 & v_45835;
assign v_45838 = v_45735 & v_45837;
assign v_45839 = v_45724 & v_45835;
assign v_45841 = v_45722 & v_45840;
assign v_45843 = v_45741 & v_45842;
assign v_45844 = v_45721 & v_45840;
assign v_45846 = v_45719 & v_45845;
assign v_45848 = v_45747 & v_45847;
assign v_45849 = v_45718 & v_45845;
assign v_45851 = v_45716 & v_45850;
assign v_45853 = v_45753 & v_45852;
assign v_45854 = v_45715 & v_45850;
assign v_45856 = v_45713 & v_45855;
assign v_45858 = v_45759 & v_45857;
assign v_45859 = v_45712 & v_45855;
assign v_45861 = v_45710 & v_45860;
assign v_45863 = v_45765 & v_45862;
assign v_45864 = v_45709 & v_45860;
assign v_45866 = v_45707 & v_45865;
assign v_45868 = v_45771 & v_45867;
assign v_45869 = v_45706 & v_45865;
assign v_45871 = v_45704 & v_45870;
assign v_45873 = v_45777 & v_45872;
assign v_45874 = v_45703 & v_45870;
assign v_45876 = v_45701 & v_45875;
assign v_45878 = v_45783 & v_45877;
assign v_45879 = v_45700 & v_45875;
assign v_45881 = v_45698 & v_45880;
assign v_45883 = v_45789 & v_45882;
assign v_45884 = v_45697 & v_45880;
assign v_45886 = v_45695 & v_45885;
assign v_45888 = v_45795 & v_45887;
assign v_45889 = v_45694 & v_45885;
assign v_45891 = v_45692 & v_45890;
assign v_45893 = v_45801 & v_45892;
assign v_45894 = v_45691 & v_45890;
assign v_45896 = v_45689 & v_45895;
assign v_45898 = v_45807 & v_45897;
assign v_45899 = v_45688 & v_45895;
assign v_45901 = v_45686 & v_45900;
assign v_45903 = v_45813 & v_45902;
assign v_45904 = v_45685 & v_45900;
assign v_45906 = v_45683 & v_45905;
assign v_45908 = v_45819 & v_45907;
assign v_45909 = v_45682 & v_45905;
assign v_45911 = v_45680 & v_45910;
assign v_45913 = v_45825 & v_45912;
assign v_45914 = v_45679 & v_45910;
assign v_45916 = v_45828;
assign v_45918 = v_45830 & v_45917;
assign v_45919 = v_45918;
assign v_45921 = v_45920;
assign v_45923 = ~v_6;
assign v_45925 = ~v_45924;
assign v_45926 = v_45924;
assign v_45927 = ~v_13;
assign v_45929 = ~v_45928;
assign v_45930 = v_45928;
assign v_45931 = ~v_18;
assign v_45933 = ~v_45932;
assign v_45934 = v_45932;
assign v_45935 = ~v_23;
assign v_45937 = ~v_45936;
assign v_45938 = v_45936;
assign v_45940 = ~v_45939;
assign v_45941 = ~v_30;
assign v_45942 = v_30;
assign v_45944 = ~v_45943;
assign v_45945 = ~v_35;
assign v_45946 = v_35;
assign v_45948 = ~v_45947;
assign v_45949 = ~v_40;
assign v_45950 = v_40;
assign v_45952 = ~v_45951;
assign v_45953 = ~v_45;
assign v_45954 = v_45;
assign v_45956 = ~v_45955;
assign v_45957 = ~v_50;
assign v_45958 = v_50;
assign v_45960 = ~v_45959;
assign v_45961 = ~v_55;
assign v_45962 = v_55;
assign v_45964 = ~v_45963;
assign v_45965 = ~v_60;
assign v_45966 = v_60;
assign v_45968 = ~v_45967;
assign v_45969 = ~v_65;
assign v_45970 = v_65;
assign v_45972 = ~v_45971;
assign v_45973 = ~v_70;
assign v_45974 = v_70;
assign v_45976 = ~v_45975;
assign v_45977 = ~v_75;
assign v_45978 = v_75;
assign v_45980 = ~v_45979;
assign v_45981 = ~v_80;
assign v_45982 = v_80;
assign v_45984 = ~v_45983;
assign v_45985 = ~v_85;
assign v_45986 = v_85;
assign v_45988 = ~v_45987;
assign v_45989 = ~v_90;
assign v_45990 = v_45989;
assign v_45992 = v_45991;
assign v_45994 = v_45985 & v_45993;
assign v_45996 = v_45983;
assign v_45998 = v_45995 & v_45997;
assign v_46000 = v_45981 & v_45999;
assign v_46002 = v_45979;
assign v_46004 = v_46001 & v_46003;
assign v_46006 = v_45977 & v_46005;
assign v_46008 = v_45975;
assign v_46010 = v_46007 & v_46009;
assign v_46012 = v_45973 & v_46011;
assign v_46014 = v_45971;
assign v_46016 = v_46013 & v_46015;
assign v_46018 = v_45969 & v_46017;
assign v_46020 = v_45967;
assign v_46022 = v_46019 & v_46021;
assign v_46024 = v_45965 & v_46023;
assign v_46026 = v_45963;
assign v_46028 = v_46025 & v_46027;
assign v_46030 = v_45961 & v_46029;
assign v_46032 = v_45959;
assign v_46034 = v_46031 & v_46033;
assign v_46036 = v_45957 & v_46035;
assign v_46038 = v_45955;
assign v_46040 = v_46037 & v_46039;
assign v_46042 = v_45953 & v_46041;
assign v_46044 = v_45951;
assign v_46046 = v_46043 & v_46045;
assign v_46048 = v_45949 & v_46047;
assign v_46050 = v_45947;
assign v_46052 = v_46049 & v_46051;
assign v_46054 = v_45945 & v_46053;
assign v_46056 = v_45943;
assign v_46058 = v_46055 & v_46057;
assign v_46060 = v_45941 & v_46059;
assign v_46062 = v_45939;
assign v_46064 = v_46061 & v_46063;
assign v_46066 = v_45937 & v_46065;
assign v_46068 = v_23;
assign v_46070 = v_46067 & v_46069;
assign v_46072 = v_45933 & v_46071;
assign v_46074 = v_18;
assign v_46076 = v_46073 & v_46075;
assign v_46078 = v_45929 & v_46077;
assign v_46080 = v_13;
assign v_46082 = v_46079 & v_46081;
assign v_46084 = v_45925 & v_46083;
assign v_46086 = v_6;
assign v_46088 = v_46085 & v_46087;
assign v_46089 = v_46088;
assign v_46091 = v_45987;
assign v_46092 = v_90;
assign v_46093 = v_46092;
assign v_46094 = v_46091 & v_46093;
assign v_46095 = v_46094;
assign v_46096 = v_45985 & v_46095;
assign v_46098 = v_45996 & v_46097;
assign v_46099 = v_45984 & v_46095;
assign v_46101 = v_45981 & v_46100;
assign v_46103 = v_46002 & v_46102;
assign v_46104 = v_45980 & v_46100;
assign v_46106 = v_45977 & v_46105;
assign v_46108 = v_46008 & v_46107;
assign v_46109 = v_45976 & v_46105;
assign v_46111 = v_45973 & v_46110;
assign v_46113 = v_46014 & v_46112;
assign v_46114 = v_45972 & v_46110;
assign v_46116 = v_45969 & v_46115;
assign v_46118 = v_46020 & v_46117;
assign v_46119 = v_45968 & v_46115;
assign v_46121 = v_45965 & v_46120;
assign v_46123 = v_46026 & v_46122;
assign v_46124 = v_45964 & v_46120;
assign v_46126 = v_45961 & v_46125;
assign v_46128 = v_46032 & v_46127;
assign v_46129 = v_45960 & v_46125;
assign v_46131 = v_45957 & v_46130;
assign v_46133 = v_46038 & v_46132;
assign v_46134 = v_45956 & v_46130;
assign v_46136 = v_45953 & v_46135;
assign v_46138 = v_46044 & v_46137;
assign v_46139 = v_45952 & v_46135;
assign v_46141 = v_45949 & v_46140;
assign v_46143 = v_46050 & v_46142;
assign v_46144 = v_45948 & v_46140;
assign v_46146 = v_45945 & v_46145;
assign v_46148 = v_46056 & v_46147;
assign v_46149 = v_45944 & v_46145;
assign v_46151 = v_45941 & v_46150;
assign v_46153 = v_46062 & v_46152;
assign v_46154 = v_45940 & v_46150;
assign v_46156 = v_45937 & v_46155;
assign v_46158 = v_46068 & v_46157;
assign v_46159 = v_45935 & v_46155;
assign v_46161 = v_45933 & v_46160;
assign v_46163 = v_46074 & v_46162;
assign v_46164 = v_45931 & v_46160;
assign v_46166 = v_45929 & v_46165;
assign v_46168 = v_46080 & v_46167;
assign v_46169 = v_45927 & v_46165;
assign v_46171 = v_45925 & v_46170;
assign v_46173 = v_46086 & v_46172;
assign v_46174 = v_45923 & v_46170;
assign v_46176 = v_46175;
assign v_46178 = v_46090 & v_46177;
assign v_46179 = v_46178;
assign v_46181 = v_46180;
assign v_46183 = ~v_283;
assign v_46184 = ~v_45924;
assign v_46185 = v_45924;
assign v_46186 = ~v_287;
assign v_46187 = ~v_45928;
assign v_46188 = v_45928;
assign v_46189 = ~v_291;
assign v_46190 = ~v_45932;
assign v_46191 = v_45932;
assign v_46192 = ~v_295;
assign v_46193 = ~v_45936;
assign v_46194 = v_45936;
assign v_46195 = ~v_45939;
assign v_46196 = ~v_300;
assign v_46197 = v_300;
assign v_46198 = ~v_45943;
assign v_46199 = ~v_304;
assign v_46200 = v_304;
assign v_46201 = ~v_45947;
assign v_46202 = ~v_308;
assign v_46203 = v_308;
assign v_46204 = ~v_45951;
assign v_46205 = ~v_312;
assign v_46206 = v_312;
assign v_46207 = ~v_45955;
assign v_46208 = ~v_316;
assign v_46209 = v_316;
assign v_46210 = ~v_45959;
assign v_46211 = ~v_320;
assign v_46212 = v_320;
assign v_46213 = ~v_45963;
assign v_46214 = ~v_324;
assign v_46215 = v_324;
assign v_46216 = ~v_45967;
assign v_46217 = ~v_328;
assign v_46218 = v_328;
assign v_46219 = ~v_45971;
assign v_46220 = ~v_332;
assign v_46221 = v_332;
assign v_46222 = ~v_45975;
assign v_46223 = ~v_336;
assign v_46224 = v_336;
assign v_46225 = ~v_45979;
assign v_46226 = ~v_340;
assign v_46227 = v_340;
assign v_46228 = ~v_45983;
assign v_46229 = ~v_344;
assign v_46230 = v_344;
assign v_46231 = ~v_45987;
assign v_46232 = ~v_348;
assign v_46233 = v_46232;
assign v_46235 = v_46234;
assign v_46237 = v_46229 & v_46236;
assign v_46239 = v_45983;
assign v_46241 = v_46238 & v_46240;
assign v_46243 = v_46226 & v_46242;
assign v_46245 = v_45979;
assign v_46247 = v_46244 & v_46246;
assign v_46249 = v_46223 & v_46248;
assign v_46251 = v_45975;
assign v_46253 = v_46250 & v_46252;
assign v_46255 = v_46220 & v_46254;
assign v_46257 = v_45971;
assign v_46259 = v_46256 & v_46258;
assign v_46261 = v_46217 & v_46260;
assign v_46263 = v_45967;
assign v_46265 = v_46262 & v_46264;
assign v_46267 = v_46214 & v_46266;
assign v_46269 = v_45963;
assign v_46271 = v_46268 & v_46270;
assign v_46273 = v_46211 & v_46272;
assign v_46275 = v_45959;
assign v_46277 = v_46274 & v_46276;
assign v_46279 = v_46208 & v_46278;
assign v_46281 = v_45955;
assign v_46283 = v_46280 & v_46282;
assign v_46285 = v_46205 & v_46284;
assign v_46287 = v_45951;
assign v_46289 = v_46286 & v_46288;
assign v_46291 = v_46202 & v_46290;
assign v_46293 = v_45947;
assign v_46295 = v_46292 & v_46294;
assign v_46297 = v_46199 & v_46296;
assign v_46299 = v_45943;
assign v_46301 = v_46298 & v_46300;
assign v_46303 = v_46196 & v_46302;
assign v_46305 = v_45939;
assign v_46307 = v_46304 & v_46306;
assign v_46309 = v_46193 & v_46308;
assign v_46311 = v_295;
assign v_46313 = v_46310 & v_46312;
assign v_46315 = v_46190 & v_46314;
assign v_46317 = v_291;
assign v_46319 = v_46316 & v_46318;
assign v_46321 = v_46187 & v_46320;
assign v_46323 = v_287;
assign v_46325 = v_46322 & v_46324;
assign v_46327 = v_46184 & v_46326;
assign v_46329 = v_283;
assign v_46331 = v_46328 & v_46330;
assign v_46332 = v_46331;
assign v_46334 = v_45987;
assign v_46335 = v_348;
assign v_46336 = v_46335;
assign v_46337 = v_46334 & v_46336;
assign v_46338 = v_46337;
assign v_46339 = v_46229 & v_46338;
assign v_46341 = v_46239 & v_46340;
assign v_46342 = v_46228 & v_46338;
assign v_46344 = v_46226 & v_46343;
assign v_46346 = v_46245 & v_46345;
assign v_46347 = v_46225 & v_46343;
assign v_46349 = v_46223 & v_46348;
assign v_46351 = v_46251 & v_46350;
assign v_46352 = v_46222 & v_46348;
assign v_46354 = v_46220 & v_46353;
assign v_46356 = v_46257 & v_46355;
assign v_46357 = v_46219 & v_46353;
assign v_46359 = v_46217 & v_46358;
assign v_46361 = v_46263 & v_46360;
assign v_46362 = v_46216 & v_46358;
assign v_46364 = v_46214 & v_46363;
assign v_46366 = v_46269 & v_46365;
assign v_46367 = v_46213 & v_46363;
assign v_46369 = v_46211 & v_46368;
assign v_46371 = v_46275 & v_46370;
assign v_46372 = v_46210 & v_46368;
assign v_46374 = v_46208 & v_46373;
assign v_46376 = v_46281 & v_46375;
assign v_46377 = v_46207 & v_46373;
assign v_46379 = v_46205 & v_46378;
assign v_46381 = v_46287 & v_46380;
assign v_46382 = v_46204 & v_46378;
assign v_46384 = v_46202 & v_46383;
assign v_46386 = v_46293 & v_46385;
assign v_46387 = v_46201 & v_46383;
assign v_46389 = v_46199 & v_46388;
assign v_46391 = v_46299 & v_46390;
assign v_46392 = v_46198 & v_46388;
assign v_46394 = v_46196 & v_46393;
assign v_46396 = v_46305 & v_46395;
assign v_46397 = v_46195 & v_46393;
assign v_46399 = v_46193 & v_46398;
assign v_46401 = v_46311 & v_46400;
assign v_46402 = v_46192 & v_46398;
assign v_46404 = v_46190 & v_46403;
assign v_46406 = v_46317 & v_46405;
assign v_46407 = v_46189 & v_46403;
assign v_46409 = v_46187 & v_46408;
assign v_46411 = v_46323 & v_46410;
assign v_46412 = v_46186 & v_46408;
assign v_46414 = v_46184 & v_46413;
assign v_46416 = v_46329 & v_46415;
assign v_46417 = v_46183 & v_46413;
assign v_46419 = v_46418;
assign v_46421 = v_46333 & v_46420;
assign v_46422 = v_46421;
assign v_46424 = v_46423;
assign v_46426 = ~v_543;
assign v_46427 = ~v_45924;
assign v_46428 = v_45924;
assign v_46429 = ~v_547;
assign v_46430 = ~v_45928;
assign v_46431 = v_45928;
assign v_46432 = ~v_551;
assign v_46433 = ~v_45932;
assign v_46434 = v_45932;
assign v_46435 = ~v_555;
assign v_46436 = ~v_45936;
assign v_46437 = v_45936;
assign v_46438 = ~v_45939;
assign v_46439 = ~v_560;
assign v_46440 = v_560;
assign v_46441 = ~v_45943;
assign v_46442 = ~v_564;
assign v_46443 = v_564;
assign v_46444 = ~v_45947;
assign v_46445 = ~v_568;
assign v_46446 = v_568;
assign v_46447 = ~v_45951;
assign v_46448 = ~v_572;
assign v_46449 = v_572;
assign v_46450 = ~v_45955;
assign v_46451 = ~v_576;
assign v_46452 = v_576;
assign v_46453 = ~v_45959;
assign v_46454 = ~v_580;
assign v_46455 = v_580;
assign v_46456 = ~v_45963;
assign v_46457 = ~v_584;
assign v_46458 = v_584;
assign v_46459 = ~v_45967;
assign v_46460 = ~v_588;
assign v_46461 = v_588;
assign v_46462 = ~v_45971;
assign v_46463 = ~v_592;
assign v_46464 = v_592;
assign v_46465 = ~v_45975;
assign v_46466 = ~v_596;
assign v_46467 = v_596;
assign v_46468 = ~v_45979;
assign v_46469 = ~v_600;
assign v_46470 = v_600;
assign v_46471 = ~v_45983;
assign v_46472 = ~v_604;
assign v_46473 = v_604;
assign v_46474 = ~v_45987;
assign v_46475 = ~v_608;
assign v_46476 = v_46475;
assign v_46478 = v_46477;
assign v_46480 = v_46472 & v_46479;
assign v_46482 = v_45983;
assign v_46484 = v_46481 & v_46483;
assign v_46486 = v_46469 & v_46485;
assign v_46488 = v_45979;
assign v_46490 = v_46487 & v_46489;
assign v_46492 = v_46466 & v_46491;
assign v_46494 = v_45975;
assign v_46496 = v_46493 & v_46495;
assign v_46498 = v_46463 & v_46497;
assign v_46500 = v_45971;
assign v_46502 = v_46499 & v_46501;
assign v_46504 = v_46460 & v_46503;
assign v_46506 = v_45967;
assign v_46508 = v_46505 & v_46507;
assign v_46510 = v_46457 & v_46509;
assign v_46512 = v_45963;
assign v_46514 = v_46511 & v_46513;
assign v_46516 = v_46454 & v_46515;
assign v_46518 = v_45959;
assign v_46520 = v_46517 & v_46519;
assign v_46522 = v_46451 & v_46521;
assign v_46524 = v_45955;
assign v_46526 = v_46523 & v_46525;
assign v_46528 = v_46448 & v_46527;
assign v_46530 = v_45951;
assign v_46532 = v_46529 & v_46531;
assign v_46534 = v_46445 & v_46533;
assign v_46536 = v_45947;
assign v_46538 = v_46535 & v_46537;
assign v_46540 = v_46442 & v_46539;
assign v_46542 = v_45943;
assign v_46544 = v_46541 & v_46543;
assign v_46546 = v_46439 & v_46545;
assign v_46548 = v_45939;
assign v_46550 = v_46547 & v_46549;
assign v_46552 = v_46436 & v_46551;
assign v_46554 = v_555;
assign v_46556 = v_46553 & v_46555;
assign v_46558 = v_46433 & v_46557;
assign v_46560 = v_551;
assign v_46562 = v_46559 & v_46561;
assign v_46564 = v_46430 & v_46563;
assign v_46566 = v_547;
assign v_46568 = v_46565 & v_46567;
assign v_46570 = v_46427 & v_46569;
assign v_46572 = v_543;
assign v_46574 = v_46571 & v_46573;
assign v_46575 = v_46574;
assign v_46577 = v_45987;
assign v_46578 = v_608;
assign v_46579 = v_46578;
assign v_46580 = v_46577 & v_46579;
assign v_46581 = v_46580;
assign v_46582 = v_46472 & v_46581;
assign v_46584 = v_46482 & v_46583;
assign v_46585 = v_46471 & v_46581;
assign v_46587 = v_46469 & v_46586;
assign v_46589 = v_46488 & v_46588;
assign v_46590 = v_46468 & v_46586;
assign v_46592 = v_46466 & v_46591;
assign v_46594 = v_46494 & v_46593;
assign v_46595 = v_46465 & v_46591;
assign v_46597 = v_46463 & v_46596;
assign v_46599 = v_46500 & v_46598;
assign v_46600 = v_46462 & v_46596;
assign v_46602 = v_46460 & v_46601;
assign v_46604 = v_46506 & v_46603;
assign v_46605 = v_46459 & v_46601;
assign v_46607 = v_46457 & v_46606;
assign v_46609 = v_46512 & v_46608;
assign v_46610 = v_46456 & v_46606;
assign v_46612 = v_46454 & v_46611;
assign v_46614 = v_46518 & v_46613;
assign v_46615 = v_46453 & v_46611;
assign v_46617 = v_46451 & v_46616;
assign v_46619 = v_46524 & v_46618;
assign v_46620 = v_46450 & v_46616;
assign v_46622 = v_46448 & v_46621;
assign v_46624 = v_46530 & v_46623;
assign v_46625 = v_46447 & v_46621;
assign v_46627 = v_46445 & v_46626;
assign v_46629 = v_46536 & v_46628;
assign v_46630 = v_46444 & v_46626;
assign v_46632 = v_46442 & v_46631;
assign v_46634 = v_46542 & v_46633;
assign v_46635 = v_46441 & v_46631;
assign v_46637 = v_46439 & v_46636;
assign v_46639 = v_46548 & v_46638;
assign v_46640 = v_46438 & v_46636;
assign v_46642 = v_46436 & v_46641;
assign v_46644 = v_46554 & v_46643;
assign v_46645 = v_46435 & v_46641;
assign v_46647 = v_46433 & v_46646;
assign v_46649 = v_46560 & v_46648;
assign v_46650 = v_46432 & v_46646;
assign v_46652 = v_46430 & v_46651;
assign v_46654 = v_46566 & v_46653;
assign v_46655 = v_46429 & v_46651;
assign v_46657 = v_46427 & v_46656;
assign v_46659 = v_46572 & v_46658;
assign v_46660 = v_46426 & v_46656;
assign v_46662 = v_46661;
assign v_46664 = v_46576 & v_46663;
assign v_46665 = v_46664;
assign v_46667 = v_46666;
assign v_46669 = ~v_803;
assign v_46670 = ~v_45924;
assign v_46671 = v_45924;
assign v_46672 = ~v_807;
assign v_46673 = ~v_45928;
assign v_46674 = v_45928;
assign v_46675 = ~v_811;
assign v_46676 = ~v_45932;
assign v_46677 = v_45932;
assign v_46678 = ~v_815;
assign v_46679 = ~v_45936;
assign v_46680 = v_45936;
assign v_46681 = ~v_45939;
assign v_46682 = ~v_820;
assign v_46683 = v_820;
assign v_46684 = ~v_45943;
assign v_46685 = ~v_824;
assign v_46686 = v_824;
assign v_46687 = ~v_45947;
assign v_46688 = ~v_828;
assign v_46689 = v_828;
assign v_46690 = ~v_45951;
assign v_46691 = ~v_832;
assign v_46692 = v_832;
assign v_46693 = ~v_45955;
assign v_46694 = ~v_836;
assign v_46695 = v_836;
assign v_46696 = ~v_45959;
assign v_46697 = ~v_840;
assign v_46698 = v_840;
assign v_46699 = ~v_45963;
assign v_46700 = ~v_844;
assign v_46701 = v_844;
assign v_46702 = ~v_45967;
assign v_46703 = ~v_848;
assign v_46704 = v_848;
assign v_46705 = ~v_45971;
assign v_46706 = ~v_852;
assign v_46707 = v_852;
assign v_46708 = ~v_45975;
assign v_46709 = ~v_856;
assign v_46710 = v_856;
assign v_46711 = ~v_45979;
assign v_46712 = ~v_860;
assign v_46713 = v_860;
assign v_46714 = ~v_45983;
assign v_46715 = ~v_864;
assign v_46716 = v_864;
assign v_46717 = ~v_45987;
assign v_46718 = ~v_868;
assign v_46719 = v_46718;
assign v_46721 = v_46720;
assign v_46723 = v_46715 & v_46722;
assign v_46725 = v_45983;
assign v_46727 = v_46724 & v_46726;
assign v_46729 = v_46712 & v_46728;
assign v_46731 = v_45979;
assign v_46733 = v_46730 & v_46732;
assign v_46735 = v_46709 & v_46734;
assign v_46737 = v_45975;
assign v_46739 = v_46736 & v_46738;
assign v_46741 = v_46706 & v_46740;
assign v_46743 = v_45971;
assign v_46745 = v_46742 & v_46744;
assign v_46747 = v_46703 & v_46746;
assign v_46749 = v_45967;
assign v_46751 = v_46748 & v_46750;
assign v_46753 = v_46700 & v_46752;
assign v_46755 = v_45963;
assign v_46757 = v_46754 & v_46756;
assign v_46759 = v_46697 & v_46758;
assign v_46761 = v_45959;
assign v_46763 = v_46760 & v_46762;
assign v_46765 = v_46694 & v_46764;
assign v_46767 = v_45955;
assign v_46769 = v_46766 & v_46768;
assign v_46771 = v_46691 & v_46770;
assign v_46773 = v_45951;
assign v_46775 = v_46772 & v_46774;
assign v_46777 = v_46688 & v_46776;
assign v_46779 = v_45947;
assign v_46781 = v_46778 & v_46780;
assign v_46783 = v_46685 & v_46782;
assign v_46785 = v_45943;
assign v_46787 = v_46784 & v_46786;
assign v_46789 = v_46682 & v_46788;
assign v_46791 = v_45939;
assign v_46793 = v_46790 & v_46792;
assign v_46795 = v_46679 & v_46794;
assign v_46797 = v_815;
assign v_46799 = v_46796 & v_46798;
assign v_46801 = v_46676 & v_46800;
assign v_46803 = v_811;
assign v_46805 = v_46802 & v_46804;
assign v_46807 = v_46673 & v_46806;
assign v_46809 = v_807;
assign v_46811 = v_46808 & v_46810;
assign v_46813 = v_46670 & v_46812;
assign v_46815 = v_803;
assign v_46817 = v_46814 & v_46816;
assign v_46818 = v_46817;
assign v_46820 = v_45987;
assign v_46821 = v_868;
assign v_46822 = v_46821;
assign v_46823 = v_46820 & v_46822;
assign v_46824 = v_46823;
assign v_46825 = v_46715 & v_46824;
assign v_46827 = v_46725 & v_46826;
assign v_46828 = v_46714 & v_46824;
assign v_46830 = v_46712 & v_46829;
assign v_46832 = v_46731 & v_46831;
assign v_46833 = v_46711 & v_46829;
assign v_46835 = v_46709 & v_46834;
assign v_46837 = v_46737 & v_46836;
assign v_46838 = v_46708 & v_46834;
assign v_46840 = v_46706 & v_46839;
assign v_46842 = v_46743 & v_46841;
assign v_46843 = v_46705 & v_46839;
assign v_46845 = v_46703 & v_46844;
assign v_46847 = v_46749 & v_46846;
assign v_46848 = v_46702 & v_46844;
assign v_46850 = v_46700 & v_46849;
assign v_46852 = v_46755 & v_46851;
assign v_46853 = v_46699 & v_46849;
assign v_46855 = v_46697 & v_46854;
assign v_46857 = v_46761 & v_46856;
assign v_46858 = v_46696 & v_46854;
assign v_46860 = v_46694 & v_46859;
assign v_46862 = v_46767 & v_46861;
assign v_46863 = v_46693 & v_46859;
assign v_46865 = v_46691 & v_46864;
assign v_46867 = v_46773 & v_46866;
assign v_46868 = v_46690 & v_46864;
assign v_46870 = v_46688 & v_46869;
assign v_46872 = v_46779 & v_46871;
assign v_46873 = v_46687 & v_46869;
assign v_46875 = v_46685 & v_46874;
assign v_46877 = v_46785 & v_46876;
assign v_46878 = v_46684 & v_46874;
assign v_46880 = v_46682 & v_46879;
assign v_46882 = v_46791 & v_46881;
assign v_46883 = v_46681 & v_46879;
assign v_46885 = v_46679 & v_46884;
assign v_46887 = v_46797 & v_46886;
assign v_46888 = v_46678 & v_46884;
assign v_46890 = v_46676 & v_46889;
assign v_46892 = v_46803 & v_46891;
assign v_46893 = v_46675 & v_46889;
assign v_46895 = v_46673 & v_46894;
assign v_46897 = v_46809 & v_46896;
assign v_46898 = v_46672 & v_46894;
assign v_46900 = v_46670 & v_46899;
assign v_46902 = v_46815 & v_46901;
assign v_46903 = v_46669 & v_46899;
assign v_46905 = v_46904;
assign v_46907 = v_46819 & v_46906;
assign v_46908 = v_46907;
assign v_46910 = v_46909;
assign v_46912 = ~v_1063;
assign v_46913 = ~v_45924;
assign v_46914 = v_45924;
assign v_46915 = ~v_1067;
assign v_46916 = ~v_45928;
assign v_46917 = v_45928;
assign v_46918 = ~v_1071;
assign v_46919 = ~v_45932;
assign v_46920 = v_45932;
assign v_46921 = ~v_1075;
assign v_46922 = ~v_45936;
assign v_46923 = v_45936;
assign v_46924 = ~v_45939;
assign v_46925 = ~v_1080;
assign v_46926 = v_1080;
assign v_46927 = ~v_45943;
assign v_46928 = ~v_1084;
assign v_46929 = v_1084;
assign v_46930 = ~v_45947;
assign v_46931 = ~v_1088;
assign v_46932 = v_1088;
assign v_46933 = ~v_45951;
assign v_46934 = ~v_1092;
assign v_46935 = v_1092;
assign v_46936 = ~v_45955;
assign v_46937 = ~v_1096;
assign v_46938 = v_1096;
assign v_46939 = ~v_45959;
assign v_46940 = ~v_1100;
assign v_46941 = v_1100;
assign v_46942 = ~v_45963;
assign v_46943 = ~v_1104;
assign v_46944 = v_1104;
assign v_46945 = ~v_45967;
assign v_46946 = ~v_1108;
assign v_46947 = v_1108;
assign v_46948 = ~v_45971;
assign v_46949 = ~v_1112;
assign v_46950 = v_1112;
assign v_46951 = ~v_45975;
assign v_46952 = ~v_1116;
assign v_46953 = v_1116;
assign v_46954 = ~v_45979;
assign v_46955 = ~v_1120;
assign v_46956 = v_1120;
assign v_46957 = ~v_45983;
assign v_46958 = ~v_1124;
assign v_46959 = v_1124;
assign v_46960 = ~v_45987;
assign v_46961 = ~v_1128;
assign v_46962 = v_46961;
assign v_46964 = v_46963;
assign v_46966 = v_46958 & v_46965;
assign v_46968 = v_45983;
assign v_46970 = v_46967 & v_46969;
assign v_46972 = v_46955 & v_46971;
assign v_46974 = v_45979;
assign v_46976 = v_46973 & v_46975;
assign v_46978 = v_46952 & v_46977;
assign v_46980 = v_45975;
assign v_46982 = v_46979 & v_46981;
assign v_46984 = v_46949 & v_46983;
assign v_46986 = v_45971;
assign v_46988 = v_46985 & v_46987;
assign v_46990 = v_46946 & v_46989;
assign v_46992 = v_45967;
assign v_46994 = v_46991 & v_46993;
assign v_46996 = v_46943 & v_46995;
assign v_46998 = v_45963;
assign v_47000 = v_46997 & v_46999;
assign v_47002 = v_46940 & v_47001;
assign v_47004 = v_45959;
assign v_47006 = v_47003 & v_47005;
assign v_47008 = v_46937 & v_47007;
assign v_47010 = v_45955;
assign v_47012 = v_47009 & v_47011;
assign v_47014 = v_46934 & v_47013;
assign v_47016 = v_45951;
assign v_47018 = v_47015 & v_47017;
assign v_47020 = v_46931 & v_47019;
assign v_47022 = v_45947;
assign v_47024 = v_47021 & v_47023;
assign v_47026 = v_46928 & v_47025;
assign v_47028 = v_45943;
assign v_47030 = v_47027 & v_47029;
assign v_47032 = v_46925 & v_47031;
assign v_47034 = v_45939;
assign v_47036 = v_47033 & v_47035;
assign v_47038 = v_46922 & v_47037;
assign v_47040 = v_1075;
assign v_47042 = v_47039 & v_47041;
assign v_47044 = v_46919 & v_47043;
assign v_47046 = v_1071;
assign v_47048 = v_47045 & v_47047;
assign v_47050 = v_46916 & v_47049;
assign v_47052 = v_1067;
assign v_47054 = v_47051 & v_47053;
assign v_47056 = v_46913 & v_47055;
assign v_47058 = v_1063;
assign v_47060 = v_47057 & v_47059;
assign v_47061 = v_47060;
assign v_47063 = v_45987;
assign v_47064 = v_1128;
assign v_47065 = v_47064;
assign v_47066 = v_47063 & v_47065;
assign v_47067 = v_47066;
assign v_47068 = v_46958 & v_47067;
assign v_47070 = v_46968 & v_47069;
assign v_47071 = v_46957 & v_47067;
assign v_47073 = v_46955 & v_47072;
assign v_47075 = v_46974 & v_47074;
assign v_47076 = v_46954 & v_47072;
assign v_47078 = v_46952 & v_47077;
assign v_47080 = v_46980 & v_47079;
assign v_47081 = v_46951 & v_47077;
assign v_47083 = v_46949 & v_47082;
assign v_47085 = v_46986 & v_47084;
assign v_47086 = v_46948 & v_47082;
assign v_47088 = v_46946 & v_47087;
assign v_47090 = v_46992 & v_47089;
assign v_47091 = v_46945 & v_47087;
assign v_47093 = v_46943 & v_47092;
assign v_47095 = v_46998 & v_47094;
assign v_47096 = v_46942 & v_47092;
assign v_47098 = v_46940 & v_47097;
assign v_47100 = v_47004 & v_47099;
assign v_47101 = v_46939 & v_47097;
assign v_47103 = v_46937 & v_47102;
assign v_47105 = v_47010 & v_47104;
assign v_47106 = v_46936 & v_47102;
assign v_47108 = v_46934 & v_47107;
assign v_47110 = v_47016 & v_47109;
assign v_47111 = v_46933 & v_47107;
assign v_47113 = v_46931 & v_47112;
assign v_47115 = v_47022 & v_47114;
assign v_47116 = v_46930 & v_47112;
assign v_47118 = v_46928 & v_47117;
assign v_47120 = v_47028 & v_47119;
assign v_47121 = v_46927 & v_47117;
assign v_47123 = v_46925 & v_47122;
assign v_47125 = v_47034 & v_47124;
assign v_47126 = v_46924 & v_47122;
assign v_47128 = v_46922 & v_47127;
assign v_47130 = v_47040 & v_47129;
assign v_47131 = v_46921 & v_47127;
assign v_47133 = v_46919 & v_47132;
assign v_47135 = v_47046 & v_47134;
assign v_47136 = v_46918 & v_47132;
assign v_47138 = v_46916 & v_47137;
assign v_47140 = v_47052 & v_47139;
assign v_47141 = v_46915 & v_47137;
assign v_47143 = v_46913 & v_47142;
assign v_47145 = v_47058 & v_47144;
assign v_47146 = v_46912 & v_47142;
assign v_47148 = v_47147;
assign v_47150 = v_47062 & v_47149;
assign v_47151 = v_47150;
assign v_47153 = v_47152;
assign v_47155 = ~v_1323;
assign v_47156 = ~v_45924;
assign v_47157 = v_45924;
assign v_47158 = ~v_1327;
assign v_47159 = ~v_45928;
assign v_47160 = v_45928;
assign v_47161 = ~v_1331;
assign v_47162 = ~v_45932;
assign v_47163 = v_45932;
assign v_47164 = ~v_1335;
assign v_47165 = ~v_45936;
assign v_47166 = v_45936;
assign v_47167 = ~v_45939;
assign v_47168 = ~v_1340;
assign v_47169 = v_1340;
assign v_47170 = ~v_45943;
assign v_47171 = ~v_1344;
assign v_47172 = v_1344;
assign v_47173 = ~v_45947;
assign v_47174 = ~v_1348;
assign v_47175 = v_1348;
assign v_47176 = ~v_45951;
assign v_47177 = ~v_1352;
assign v_47178 = v_1352;
assign v_47179 = ~v_45955;
assign v_47180 = ~v_1356;
assign v_47181 = v_1356;
assign v_47182 = ~v_45959;
assign v_47183 = ~v_1360;
assign v_47184 = v_1360;
assign v_47185 = ~v_45963;
assign v_47186 = ~v_1364;
assign v_47187 = v_1364;
assign v_47188 = ~v_45967;
assign v_47189 = ~v_1368;
assign v_47190 = v_1368;
assign v_47191 = ~v_45971;
assign v_47192 = ~v_1372;
assign v_47193 = v_1372;
assign v_47194 = ~v_45975;
assign v_47195 = ~v_1376;
assign v_47196 = v_1376;
assign v_47197 = ~v_45979;
assign v_47198 = ~v_1380;
assign v_47199 = v_1380;
assign v_47200 = ~v_45983;
assign v_47201 = ~v_1384;
assign v_47202 = v_1384;
assign v_47203 = ~v_45987;
assign v_47204 = ~v_1388;
assign v_47205 = v_47204;
assign v_47207 = v_47206;
assign v_47209 = v_47201 & v_47208;
assign v_47211 = v_45983;
assign v_47213 = v_47210 & v_47212;
assign v_47215 = v_47198 & v_47214;
assign v_47217 = v_45979;
assign v_47219 = v_47216 & v_47218;
assign v_47221 = v_47195 & v_47220;
assign v_47223 = v_45975;
assign v_47225 = v_47222 & v_47224;
assign v_47227 = v_47192 & v_47226;
assign v_47229 = v_45971;
assign v_47231 = v_47228 & v_47230;
assign v_47233 = v_47189 & v_47232;
assign v_47235 = v_45967;
assign v_47237 = v_47234 & v_47236;
assign v_47239 = v_47186 & v_47238;
assign v_47241 = v_45963;
assign v_47243 = v_47240 & v_47242;
assign v_47245 = v_47183 & v_47244;
assign v_47247 = v_45959;
assign v_47249 = v_47246 & v_47248;
assign v_47251 = v_47180 & v_47250;
assign v_47253 = v_45955;
assign v_47255 = v_47252 & v_47254;
assign v_47257 = v_47177 & v_47256;
assign v_47259 = v_45951;
assign v_47261 = v_47258 & v_47260;
assign v_47263 = v_47174 & v_47262;
assign v_47265 = v_45947;
assign v_47267 = v_47264 & v_47266;
assign v_47269 = v_47171 & v_47268;
assign v_47271 = v_45943;
assign v_47273 = v_47270 & v_47272;
assign v_47275 = v_47168 & v_47274;
assign v_47277 = v_45939;
assign v_47279 = v_47276 & v_47278;
assign v_47281 = v_47165 & v_47280;
assign v_47283 = v_1335;
assign v_47285 = v_47282 & v_47284;
assign v_47287 = v_47162 & v_47286;
assign v_47289 = v_1331;
assign v_47291 = v_47288 & v_47290;
assign v_47293 = v_47159 & v_47292;
assign v_47295 = v_1327;
assign v_47297 = v_47294 & v_47296;
assign v_47299 = v_47156 & v_47298;
assign v_47301 = v_1323;
assign v_47303 = v_47300 & v_47302;
assign v_47304 = v_47303;
assign v_47306 = v_45987;
assign v_47307 = v_1388;
assign v_47308 = v_47307;
assign v_47309 = v_47306 & v_47308;
assign v_47310 = v_47309;
assign v_47311 = v_47201 & v_47310;
assign v_47313 = v_47211 & v_47312;
assign v_47314 = v_47200 & v_47310;
assign v_47316 = v_47198 & v_47315;
assign v_47318 = v_47217 & v_47317;
assign v_47319 = v_47197 & v_47315;
assign v_47321 = v_47195 & v_47320;
assign v_47323 = v_47223 & v_47322;
assign v_47324 = v_47194 & v_47320;
assign v_47326 = v_47192 & v_47325;
assign v_47328 = v_47229 & v_47327;
assign v_47329 = v_47191 & v_47325;
assign v_47331 = v_47189 & v_47330;
assign v_47333 = v_47235 & v_47332;
assign v_47334 = v_47188 & v_47330;
assign v_47336 = v_47186 & v_47335;
assign v_47338 = v_47241 & v_47337;
assign v_47339 = v_47185 & v_47335;
assign v_47341 = v_47183 & v_47340;
assign v_47343 = v_47247 & v_47342;
assign v_47344 = v_47182 & v_47340;
assign v_47346 = v_47180 & v_47345;
assign v_47348 = v_47253 & v_47347;
assign v_47349 = v_47179 & v_47345;
assign v_47351 = v_47177 & v_47350;
assign v_47353 = v_47259 & v_47352;
assign v_47354 = v_47176 & v_47350;
assign v_47356 = v_47174 & v_47355;
assign v_47358 = v_47265 & v_47357;
assign v_47359 = v_47173 & v_47355;
assign v_47361 = v_47171 & v_47360;
assign v_47363 = v_47271 & v_47362;
assign v_47364 = v_47170 & v_47360;
assign v_47366 = v_47168 & v_47365;
assign v_47368 = v_47277 & v_47367;
assign v_47369 = v_47167 & v_47365;
assign v_47371 = v_47165 & v_47370;
assign v_47373 = v_47283 & v_47372;
assign v_47374 = v_47164 & v_47370;
assign v_47376 = v_47162 & v_47375;
assign v_47378 = v_47289 & v_47377;
assign v_47379 = v_47161 & v_47375;
assign v_47381 = v_47159 & v_47380;
assign v_47383 = v_47295 & v_47382;
assign v_47384 = v_47158 & v_47380;
assign v_47386 = v_47156 & v_47385;
assign v_47388 = v_47301 & v_47387;
assign v_47389 = v_47155 & v_47385;
assign v_47391 = v_47390;
assign v_47393 = v_47305 & v_47392;
assign v_47394 = v_47393;
assign v_47396 = v_47395;
assign v_47398 = ~v_1583;
assign v_47399 = ~v_45924;
assign v_47400 = v_45924;
assign v_47401 = ~v_1587;
assign v_47402 = ~v_45928;
assign v_47403 = v_45928;
assign v_47404 = ~v_1591;
assign v_47405 = ~v_45932;
assign v_47406 = v_45932;
assign v_47407 = ~v_1595;
assign v_47408 = ~v_45936;
assign v_47409 = v_45936;
assign v_47410 = ~v_45939;
assign v_47411 = ~v_1600;
assign v_47412 = v_1600;
assign v_47413 = ~v_45943;
assign v_47414 = ~v_1604;
assign v_47415 = v_1604;
assign v_47416 = ~v_45947;
assign v_47417 = ~v_1608;
assign v_47418 = v_1608;
assign v_47419 = ~v_45951;
assign v_47420 = ~v_1612;
assign v_47421 = v_1612;
assign v_47422 = ~v_45955;
assign v_47423 = ~v_1616;
assign v_47424 = v_1616;
assign v_47425 = ~v_45959;
assign v_47426 = ~v_1620;
assign v_47427 = v_1620;
assign v_47428 = ~v_45963;
assign v_47429 = ~v_1624;
assign v_47430 = v_1624;
assign v_47431 = ~v_45967;
assign v_47432 = ~v_1628;
assign v_47433 = v_1628;
assign v_47434 = ~v_45971;
assign v_47435 = ~v_1632;
assign v_47436 = v_1632;
assign v_47437 = ~v_45975;
assign v_47438 = ~v_1636;
assign v_47439 = v_1636;
assign v_47440 = ~v_45979;
assign v_47441 = ~v_1640;
assign v_47442 = v_1640;
assign v_47443 = ~v_45983;
assign v_47444 = ~v_1644;
assign v_47445 = v_1644;
assign v_47446 = ~v_45987;
assign v_47447 = ~v_1648;
assign v_47448 = v_47447;
assign v_47450 = v_47449;
assign v_47452 = v_47444 & v_47451;
assign v_47454 = v_45983;
assign v_47456 = v_47453 & v_47455;
assign v_47458 = v_47441 & v_47457;
assign v_47460 = v_45979;
assign v_47462 = v_47459 & v_47461;
assign v_47464 = v_47438 & v_47463;
assign v_47466 = v_45975;
assign v_47468 = v_47465 & v_47467;
assign v_47470 = v_47435 & v_47469;
assign v_47472 = v_45971;
assign v_47474 = v_47471 & v_47473;
assign v_47476 = v_47432 & v_47475;
assign v_47478 = v_45967;
assign v_47480 = v_47477 & v_47479;
assign v_47482 = v_47429 & v_47481;
assign v_47484 = v_45963;
assign v_47486 = v_47483 & v_47485;
assign v_47488 = v_47426 & v_47487;
assign v_47490 = v_45959;
assign v_47492 = v_47489 & v_47491;
assign v_47494 = v_47423 & v_47493;
assign v_47496 = v_45955;
assign v_47498 = v_47495 & v_47497;
assign v_47500 = v_47420 & v_47499;
assign v_47502 = v_45951;
assign v_47504 = v_47501 & v_47503;
assign v_47506 = v_47417 & v_47505;
assign v_47508 = v_45947;
assign v_47510 = v_47507 & v_47509;
assign v_47512 = v_47414 & v_47511;
assign v_47514 = v_45943;
assign v_47516 = v_47513 & v_47515;
assign v_47518 = v_47411 & v_47517;
assign v_47520 = v_45939;
assign v_47522 = v_47519 & v_47521;
assign v_47524 = v_47408 & v_47523;
assign v_47526 = v_1595;
assign v_47528 = v_47525 & v_47527;
assign v_47530 = v_47405 & v_47529;
assign v_47532 = v_1591;
assign v_47534 = v_47531 & v_47533;
assign v_47536 = v_47402 & v_47535;
assign v_47538 = v_1587;
assign v_47540 = v_47537 & v_47539;
assign v_47542 = v_47399 & v_47541;
assign v_47544 = v_1583;
assign v_47546 = v_47543 & v_47545;
assign v_47547 = v_47546;
assign v_47549 = v_45987;
assign v_47550 = v_1648;
assign v_47551 = v_47550;
assign v_47552 = v_47549 & v_47551;
assign v_47553 = v_47552;
assign v_47554 = v_47444 & v_47553;
assign v_47556 = v_47454 & v_47555;
assign v_47557 = v_47443 & v_47553;
assign v_47559 = v_47441 & v_47558;
assign v_47561 = v_47460 & v_47560;
assign v_47562 = v_47440 & v_47558;
assign v_47564 = v_47438 & v_47563;
assign v_47566 = v_47466 & v_47565;
assign v_47567 = v_47437 & v_47563;
assign v_47569 = v_47435 & v_47568;
assign v_47571 = v_47472 & v_47570;
assign v_47572 = v_47434 & v_47568;
assign v_47574 = v_47432 & v_47573;
assign v_47576 = v_47478 & v_47575;
assign v_47577 = v_47431 & v_47573;
assign v_47579 = v_47429 & v_47578;
assign v_47581 = v_47484 & v_47580;
assign v_47582 = v_47428 & v_47578;
assign v_47584 = v_47426 & v_47583;
assign v_47586 = v_47490 & v_47585;
assign v_47587 = v_47425 & v_47583;
assign v_47589 = v_47423 & v_47588;
assign v_47591 = v_47496 & v_47590;
assign v_47592 = v_47422 & v_47588;
assign v_47594 = v_47420 & v_47593;
assign v_47596 = v_47502 & v_47595;
assign v_47597 = v_47419 & v_47593;
assign v_47599 = v_47417 & v_47598;
assign v_47601 = v_47508 & v_47600;
assign v_47602 = v_47416 & v_47598;
assign v_47604 = v_47414 & v_47603;
assign v_47606 = v_47514 & v_47605;
assign v_47607 = v_47413 & v_47603;
assign v_47609 = v_47411 & v_47608;
assign v_47611 = v_47520 & v_47610;
assign v_47612 = v_47410 & v_47608;
assign v_47614 = v_47408 & v_47613;
assign v_47616 = v_47526 & v_47615;
assign v_47617 = v_47407 & v_47613;
assign v_47619 = v_47405 & v_47618;
assign v_47621 = v_47532 & v_47620;
assign v_47622 = v_47404 & v_47618;
assign v_47624 = v_47402 & v_47623;
assign v_47626 = v_47538 & v_47625;
assign v_47627 = v_47401 & v_47623;
assign v_47629 = v_47399 & v_47628;
assign v_47631 = v_47544 & v_47630;
assign v_47632 = v_47398 & v_47628;
assign v_47634 = v_47633;
assign v_47636 = v_47548 & v_47635;
assign v_47637 = v_47636;
assign v_47639 = v_47638;
assign v_47641 = ~v_1843;
assign v_47642 = ~v_45924;
assign v_47643 = v_45924;
assign v_47644 = ~v_1847;
assign v_47645 = ~v_45928;
assign v_47646 = v_45928;
assign v_47647 = ~v_1851;
assign v_47648 = ~v_45932;
assign v_47649 = v_45932;
assign v_47650 = ~v_1855;
assign v_47651 = ~v_45936;
assign v_47652 = v_45936;
assign v_47653 = ~v_45939;
assign v_47654 = ~v_1860;
assign v_47655 = v_1860;
assign v_47656 = ~v_45943;
assign v_47657 = ~v_1864;
assign v_47658 = v_1864;
assign v_47659 = ~v_45947;
assign v_47660 = ~v_1868;
assign v_47661 = v_1868;
assign v_47662 = ~v_45951;
assign v_47663 = ~v_1872;
assign v_47664 = v_1872;
assign v_47665 = ~v_45955;
assign v_47666 = ~v_1876;
assign v_47667 = v_1876;
assign v_47668 = ~v_45959;
assign v_47669 = ~v_1880;
assign v_47670 = v_1880;
assign v_47671 = ~v_45963;
assign v_47672 = ~v_1884;
assign v_47673 = v_1884;
assign v_47674 = ~v_45967;
assign v_47675 = ~v_1888;
assign v_47676 = v_1888;
assign v_47677 = ~v_45971;
assign v_47678 = ~v_1892;
assign v_47679 = v_1892;
assign v_47680 = ~v_45975;
assign v_47681 = ~v_1896;
assign v_47682 = v_1896;
assign v_47683 = ~v_45979;
assign v_47684 = ~v_1900;
assign v_47685 = v_1900;
assign v_47686 = ~v_45983;
assign v_47687 = ~v_1904;
assign v_47688 = v_1904;
assign v_47689 = ~v_45987;
assign v_47690 = ~v_1908;
assign v_47691 = v_47690;
assign v_47693 = v_47692;
assign v_47695 = v_47687 & v_47694;
assign v_47697 = v_45983;
assign v_47699 = v_47696 & v_47698;
assign v_47701 = v_47684 & v_47700;
assign v_47703 = v_45979;
assign v_47705 = v_47702 & v_47704;
assign v_47707 = v_47681 & v_47706;
assign v_47709 = v_45975;
assign v_47711 = v_47708 & v_47710;
assign v_47713 = v_47678 & v_47712;
assign v_47715 = v_45971;
assign v_47717 = v_47714 & v_47716;
assign v_47719 = v_47675 & v_47718;
assign v_47721 = v_45967;
assign v_47723 = v_47720 & v_47722;
assign v_47725 = v_47672 & v_47724;
assign v_47727 = v_45963;
assign v_47729 = v_47726 & v_47728;
assign v_47731 = v_47669 & v_47730;
assign v_47733 = v_45959;
assign v_47735 = v_47732 & v_47734;
assign v_47737 = v_47666 & v_47736;
assign v_47739 = v_45955;
assign v_47741 = v_47738 & v_47740;
assign v_47743 = v_47663 & v_47742;
assign v_47745 = v_45951;
assign v_47747 = v_47744 & v_47746;
assign v_47749 = v_47660 & v_47748;
assign v_47751 = v_45947;
assign v_47753 = v_47750 & v_47752;
assign v_47755 = v_47657 & v_47754;
assign v_47757 = v_45943;
assign v_47759 = v_47756 & v_47758;
assign v_47761 = v_47654 & v_47760;
assign v_47763 = v_45939;
assign v_47765 = v_47762 & v_47764;
assign v_47767 = v_47651 & v_47766;
assign v_47769 = v_1855;
assign v_47771 = v_47768 & v_47770;
assign v_47773 = v_47648 & v_47772;
assign v_47775 = v_1851;
assign v_47777 = v_47774 & v_47776;
assign v_47779 = v_47645 & v_47778;
assign v_47781 = v_1847;
assign v_47783 = v_47780 & v_47782;
assign v_47785 = v_47642 & v_47784;
assign v_47787 = v_1843;
assign v_47789 = v_47786 & v_47788;
assign v_47790 = v_47789;
assign v_47792 = v_45987;
assign v_47793 = v_1908;
assign v_47794 = v_47793;
assign v_47795 = v_47792 & v_47794;
assign v_47796 = v_47795;
assign v_47797 = v_47687 & v_47796;
assign v_47799 = v_47697 & v_47798;
assign v_47800 = v_47686 & v_47796;
assign v_47802 = v_47684 & v_47801;
assign v_47804 = v_47703 & v_47803;
assign v_47805 = v_47683 & v_47801;
assign v_47807 = v_47681 & v_47806;
assign v_47809 = v_47709 & v_47808;
assign v_47810 = v_47680 & v_47806;
assign v_47812 = v_47678 & v_47811;
assign v_47814 = v_47715 & v_47813;
assign v_47815 = v_47677 & v_47811;
assign v_47817 = v_47675 & v_47816;
assign v_47819 = v_47721 & v_47818;
assign v_47820 = v_47674 & v_47816;
assign v_47822 = v_47672 & v_47821;
assign v_47824 = v_47727 & v_47823;
assign v_47825 = v_47671 & v_47821;
assign v_47827 = v_47669 & v_47826;
assign v_47829 = v_47733 & v_47828;
assign v_47830 = v_47668 & v_47826;
assign v_47832 = v_47666 & v_47831;
assign v_47834 = v_47739 & v_47833;
assign v_47835 = v_47665 & v_47831;
assign v_47837 = v_47663 & v_47836;
assign v_47839 = v_47745 & v_47838;
assign v_47840 = v_47662 & v_47836;
assign v_47842 = v_47660 & v_47841;
assign v_47844 = v_47751 & v_47843;
assign v_47845 = v_47659 & v_47841;
assign v_47847 = v_47657 & v_47846;
assign v_47849 = v_47757 & v_47848;
assign v_47850 = v_47656 & v_47846;
assign v_47852 = v_47654 & v_47851;
assign v_47854 = v_47763 & v_47853;
assign v_47855 = v_47653 & v_47851;
assign v_47857 = v_47651 & v_47856;
assign v_47859 = v_47769 & v_47858;
assign v_47860 = v_47650 & v_47856;
assign v_47862 = v_47648 & v_47861;
assign v_47864 = v_47775 & v_47863;
assign v_47865 = v_47647 & v_47861;
assign v_47867 = v_47645 & v_47866;
assign v_47869 = v_47781 & v_47868;
assign v_47870 = v_47644 & v_47866;
assign v_47872 = v_47642 & v_47871;
assign v_47874 = v_47787 & v_47873;
assign v_47875 = v_47641 & v_47871;
assign v_47877 = v_47876;
assign v_47879 = v_47791 & v_47878;
assign v_47880 = v_47879;
assign v_47882 = v_47881;
assign v_47884 = ~v_2103;
assign v_47885 = ~v_45924;
assign v_47886 = v_45924;
assign v_47887 = ~v_2107;
assign v_47888 = ~v_45928;
assign v_47889 = v_45928;
assign v_47890 = ~v_2111;
assign v_47891 = ~v_45932;
assign v_47892 = v_45932;
assign v_47893 = ~v_2115;
assign v_47894 = ~v_45936;
assign v_47895 = v_45936;
assign v_47896 = ~v_45939;
assign v_47897 = ~v_2120;
assign v_47898 = v_2120;
assign v_47899 = ~v_45943;
assign v_47900 = ~v_2124;
assign v_47901 = v_2124;
assign v_47902 = ~v_45947;
assign v_47903 = ~v_2128;
assign v_47904 = v_2128;
assign v_47905 = ~v_45951;
assign v_47906 = ~v_2132;
assign v_47907 = v_2132;
assign v_47908 = ~v_45955;
assign v_47909 = ~v_2136;
assign v_47910 = v_2136;
assign v_47911 = ~v_45959;
assign v_47912 = ~v_2140;
assign v_47913 = v_2140;
assign v_47914 = ~v_45963;
assign v_47915 = ~v_2144;
assign v_47916 = v_2144;
assign v_47917 = ~v_45967;
assign v_47918 = ~v_2148;
assign v_47919 = v_2148;
assign v_47920 = ~v_45971;
assign v_47921 = ~v_2152;
assign v_47922 = v_2152;
assign v_47923 = ~v_45975;
assign v_47924 = ~v_2156;
assign v_47925 = v_2156;
assign v_47926 = ~v_45979;
assign v_47927 = ~v_2160;
assign v_47928 = v_2160;
assign v_47929 = ~v_45983;
assign v_47930 = ~v_2164;
assign v_47931 = v_2164;
assign v_47932 = ~v_45987;
assign v_47933 = ~v_2168;
assign v_47934 = v_47933;
assign v_47936 = v_47935;
assign v_47938 = v_47930 & v_47937;
assign v_47940 = v_45983;
assign v_47942 = v_47939 & v_47941;
assign v_47944 = v_47927 & v_47943;
assign v_47946 = v_45979;
assign v_47948 = v_47945 & v_47947;
assign v_47950 = v_47924 & v_47949;
assign v_47952 = v_45975;
assign v_47954 = v_47951 & v_47953;
assign v_47956 = v_47921 & v_47955;
assign v_47958 = v_45971;
assign v_47960 = v_47957 & v_47959;
assign v_47962 = v_47918 & v_47961;
assign v_47964 = v_45967;
assign v_47966 = v_47963 & v_47965;
assign v_47968 = v_47915 & v_47967;
assign v_47970 = v_45963;
assign v_47972 = v_47969 & v_47971;
assign v_47974 = v_47912 & v_47973;
assign v_47976 = v_45959;
assign v_47978 = v_47975 & v_47977;
assign v_47980 = v_47909 & v_47979;
assign v_47982 = v_45955;
assign v_47984 = v_47981 & v_47983;
assign v_47986 = v_47906 & v_47985;
assign v_47988 = v_45951;
assign v_47990 = v_47987 & v_47989;
assign v_47992 = v_47903 & v_47991;
assign v_47994 = v_45947;
assign v_47996 = v_47993 & v_47995;
assign v_47998 = v_47900 & v_47997;
assign v_48000 = v_45943;
assign v_48002 = v_47999 & v_48001;
assign v_48004 = v_47897 & v_48003;
assign v_48006 = v_45939;
assign v_48008 = v_48005 & v_48007;
assign v_48010 = v_47894 & v_48009;
assign v_48012 = v_2115;
assign v_48014 = v_48011 & v_48013;
assign v_48016 = v_47891 & v_48015;
assign v_48018 = v_2111;
assign v_48020 = v_48017 & v_48019;
assign v_48022 = v_47888 & v_48021;
assign v_48024 = v_2107;
assign v_48026 = v_48023 & v_48025;
assign v_48028 = v_47885 & v_48027;
assign v_48030 = v_2103;
assign v_48032 = v_48029 & v_48031;
assign v_48033 = v_48032;
assign v_48035 = v_45987;
assign v_48036 = v_2168;
assign v_48037 = v_48036;
assign v_48038 = v_48035 & v_48037;
assign v_48039 = v_48038;
assign v_48040 = v_47930 & v_48039;
assign v_48042 = v_47940 & v_48041;
assign v_48043 = v_47929 & v_48039;
assign v_48045 = v_47927 & v_48044;
assign v_48047 = v_47946 & v_48046;
assign v_48048 = v_47926 & v_48044;
assign v_48050 = v_47924 & v_48049;
assign v_48052 = v_47952 & v_48051;
assign v_48053 = v_47923 & v_48049;
assign v_48055 = v_47921 & v_48054;
assign v_48057 = v_47958 & v_48056;
assign v_48058 = v_47920 & v_48054;
assign v_48060 = v_47918 & v_48059;
assign v_48062 = v_47964 & v_48061;
assign v_48063 = v_47917 & v_48059;
assign v_48065 = v_47915 & v_48064;
assign v_48067 = v_47970 & v_48066;
assign v_48068 = v_47914 & v_48064;
assign v_48070 = v_47912 & v_48069;
assign v_48072 = v_47976 & v_48071;
assign v_48073 = v_47911 & v_48069;
assign v_48075 = v_47909 & v_48074;
assign v_48077 = v_47982 & v_48076;
assign v_48078 = v_47908 & v_48074;
assign v_48080 = v_47906 & v_48079;
assign v_48082 = v_47988 & v_48081;
assign v_48083 = v_47905 & v_48079;
assign v_48085 = v_47903 & v_48084;
assign v_48087 = v_47994 & v_48086;
assign v_48088 = v_47902 & v_48084;
assign v_48090 = v_47900 & v_48089;
assign v_48092 = v_48000 & v_48091;
assign v_48093 = v_47899 & v_48089;
assign v_48095 = v_47897 & v_48094;
assign v_48097 = v_48006 & v_48096;
assign v_48098 = v_47896 & v_48094;
assign v_48100 = v_47894 & v_48099;
assign v_48102 = v_48012 & v_48101;
assign v_48103 = v_47893 & v_48099;
assign v_48105 = v_47891 & v_48104;
assign v_48107 = v_48018 & v_48106;
assign v_48108 = v_47890 & v_48104;
assign v_48110 = v_47888 & v_48109;
assign v_48112 = v_48024 & v_48111;
assign v_48113 = v_47887 & v_48109;
assign v_48115 = v_47885 & v_48114;
assign v_48117 = v_48030 & v_48116;
assign v_48118 = v_47884 & v_48114;
assign v_48120 = v_48119;
assign v_48122 = v_48034 & v_48121;
assign v_48123 = v_48122;
assign v_48125 = v_48124;
assign v_48127 = ~v_2363;
assign v_48128 = ~v_45924;
assign v_48129 = v_45924;
assign v_48130 = ~v_2367;
assign v_48131 = ~v_45928;
assign v_48132 = v_45928;
assign v_48133 = ~v_2371;
assign v_48134 = ~v_45932;
assign v_48135 = v_45932;
assign v_48136 = ~v_2375;
assign v_48137 = ~v_45936;
assign v_48138 = v_45936;
assign v_48139 = ~v_45939;
assign v_48140 = ~v_2380;
assign v_48141 = v_2380;
assign v_48142 = ~v_45943;
assign v_48143 = ~v_2384;
assign v_48144 = v_2384;
assign v_48145 = ~v_45947;
assign v_48146 = ~v_2388;
assign v_48147 = v_2388;
assign v_48148 = ~v_45951;
assign v_48149 = ~v_2392;
assign v_48150 = v_2392;
assign v_48151 = ~v_45955;
assign v_48152 = ~v_2396;
assign v_48153 = v_2396;
assign v_48154 = ~v_45959;
assign v_48155 = ~v_2400;
assign v_48156 = v_2400;
assign v_48157 = ~v_45963;
assign v_48158 = ~v_2404;
assign v_48159 = v_2404;
assign v_48160 = ~v_45967;
assign v_48161 = ~v_2408;
assign v_48162 = v_2408;
assign v_48163 = ~v_45971;
assign v_48164 = ~v_2412;
assign v_48165 = v_2412;
assign v_48166 = ~v_45975;
assign v_48167 = ~v_2416;
assign v_48168 = v_2416;
assign v_48169 = ~v_45979;
assign v_48170 = ~v_2420;
assign v_48171 = v_2420;
assign v_48172 = ~v_45983;
assign v_48173 = ~v_2424;
assign v_48174 = v_2424;
assign v_48175 = ~v_45987;
assign v_48176 = ~v_2428;
assign v_48177 = v_48176;
assign v_48179 = v_48178;
assign v_48181 = v_48173 & v_48180;
assign v_48183 = v_45983;
assign v_48185 = v_48182 & v_48184;
assign v_48187 = v_48170 & v_48186;
assign v_48189 = v_45979;
assign v_48191 = v_48188 & v_48190;
assign v_48193 = v_48167 & v_48192;
assign v_48195 = v_45975;
assign v_48197 = v_48194 & v_48196;
assign v_48199 = v_48164 & v_48198;
assign v_48201 = v_45971;
assign v_48203 = v_48200 & v_48202;
assign v_48205 = v_48161 & v_48204;
assign v_48207 = v_45967;
assign v_48209 = v_48206 & v_48208;
assign v_48211 = v_48158 & v_48210;
assign v_48213 = v_45963;
assign v_48215 = v_48212 & v_48214;
assign v_48217 = v_48155 & v_48216;
assign v_48219 = v_45959;
assign v_48221 = v_48218 & v_48220;
assign v_48223 = v_48152 & v_48222;
assign v_48225 = v_45955;
assign v_48227 = v_48224 & v_48226;
assign v_48229 = v_48149 & v_48228;
assign v_48231 = v_45951;
assign v_48233 = v_48230 & v_48232;
assign v_48235 = v_48146 & v_48234;
assign v_48237 = v_45947;
assign v_48239 = v_48236 & v_48238;
assign v_48241 = v_48143 & v_48240;
assign v_48243 = v_45943;
assign v_48245 = v_48242 & v_48244;
assign v_48247 = v_48140 & v_48246;
assign v_48249 = v_45939;
assign v_48251 = v_48248 & v_48250;
assign v_48253 = v_48137 & v_48252;
assign v_48255 = v_2375;
assign v_48257 = v_48254 & v_48256;
assign v_48259 = v_48134 & v_48258;
assign v_48261 = v_2371;
assign v_48263 = v_48260 & v_48262;
assign v_48265 = v_48131 & v_48264;
assign v_48267 = v_2367;
assign v_48269 = v_48266 & v_48268;
assign v_48271 = v_48128 & v_48270;
assign v_48273 = v_2363;
assign v_48275 = v_48272 & v_48274;
assign v_48276 = v_48275;
assign v_48278 = v_45987;
assign v_48279 = v_2428;
assign v_48280 = v_48279;
assign v_48281 = v_48278 & v_48280;
assign v_48282 = v_48281;
assign v_48283 = v_48173 & v_48282;
assign v_48285 = v_48183 & v_48284;
assign v_48286 = v_48172 & v_48282;
assign v_48288 = v_48170 & v_48287;
assign v_48290 = v_48189 & v_48289;
assign v_48291 = v_48169 & v_48287;
assign v_48293 = v_48167 & v_48292;
assign v_48295 = v_48195 & v_48294;
assign v_48296 = v_48166 & v_48292;
assign v_48298 = v_48164 & v_48297;
assign v_48300 = v_48201 & v_48299;
assign v_48301 = v_48163 & v_48297;
assign v_48303 = v_48161 & v_48302;
assign v_48305 = v_48207 & v_48304;
assign v_48306 = v_48160 & v_48302;
assign v_48308 = v_48158 & v_48307;
assign v_48310 = v_48213 & v_48309;
assign v_48311 = v_48157 & v_48307;
assign v_48313 = v_48155 & v_48312;
assign v_48315 = v_48219 & v_48314;
assign v_48316 = v_48154 & v_48312;
assign v_48318 = v_48152 & v_48317;
assign v_48320 = v_48225 & v_48319;
assign v_48321 = v_48151 & v_48317;
assign v_48323 = v_48149 & v_48322;
assign v_48325 = v_48231 & v_48324;
assign v_48326 = v_48148 & v_48322;
assign v_48328 = v_48146 & v_48327;
assign v_48330 = v_48237 & v_48329;
assign v_48331 = v_48145 & v_48327;
assign v_48333 = v_48143 & v_48332;
assign v_48335 = v_48243 & v_48334;
assign v_48336 = v_48142 & v_48332;
assign v_48338 = v_48140 & v_48337;
assign v_48340 = v_48249 & v_48339;
assign v_48341 = v_48139 & v_48337;
assign v_48343 = v_48137 & v_48342;
assign v_48345 = v_48255 & v_48344;
assign v_48346 = v_48136 & v_48342;
assign v_48348 = v_48134 & v_48347;
assign v_48350 = v_48261 & v_48349;
assign v_48351 = v_48133 & v_48347;
assign v_48353 = v_48131 & v_48352;
assign v_48355 = v_48267 & v_48354;
assign v_48356 = v_48130 & v_48352;
assign v_48358 = v_48128 & v_48357;
assign v_48360 = v_48273 & v_48359;
assign v_48361 = v_48127 & v_48357;
assign v_48363 = v_48362;
assign v_48365 = v_48277 & v_48364;
assign v_48366 = v_48365;
assign v_48368 = v_48367;
assign v_48370 = ~v_2623;
assign v_48371 = ~v_45924;
assign v_48372 = v_45924;
assign v_48373 = ~v_2627;
assign v_48374 = ~v_45928;
assign v_48375 = v_45928;
assign v_48376 = ~v_2631;
assign v_48377 = ~v_45932;
assign v_48378 = v_45932;
assign v_48379 = ~v_2635;
assign v_48380 = ~v_45936;
assign v_48381 = v_45936;
assign v_48382 = ~v_45939;
assign v_48383 = ~v_2640;
assign v_48384 = v_2640;
assign v_48385 = ~v_45943;
assign v_48386 = ~v_2644;
assign v_48387 = v_2644;
assign v_48388 = ~v_45947;
assign v_48389 = ~v_2648;
assign v_48390 = v_2648;
assign v_48391 = ~v_45951;
assign v_48392 = ~v_2652;
assign v_48393 = v_2652;
assign v_48394 = ~v_45955;
assign v_48395 = ~v_2656;
assign v_48396 = v_2656;
assign v_48397 = ~v_45959;
assign v_48398 = ~v_2660;
assign v_48399 = v_2660;
assign v_48400 = ~v_45963;
assign v_48401 = ~v_2664;
assign v_48402 = v_2664;
assign v_48403 = ~v_45967;
assign v_48404 = ~v_2668;
assign v_48405 = v_2668;
assign v_48406 = ~v_45971;
assign v_48407 = ~v_2672;
assign v_48408 = v_2672;
assign v_48409 = ~v_45975;
assign v_48410 = ~v_2676;
assign v_48411 = v_2676;
assign v_48412 = ~v_45979;
assign v_48413 = ~v_2680;
assign v_48414 = v_2680;
assign v_48415 = ~v_45983;
assign v_48416 = ~v_2684;
assign v_48417 = v_2684;
assign v_48418 = ~v_45987;
assign v_48419 = ~v_2688;
assign v_48420 = v_48419;
assign v_48422 = v_48421;
assign v_48424 = v_48416 & v_48423;
assign v_48426 = v_45983;
assign v_48428 = v_48425 & v_48427;
assign v_48430 = v_48413 & v_48429;
assign v_48432 = v_45979;
assign v_48434 = v_48431 & v_48433;
assign v_48436 = v_48410 & v_48435;
assign v_48438 = v_45975;
assign v_48440 = v_48437 & v_48439;
assign v_48442 = v_48407 & v_48441;
assign v_48444 = v_45971;
assign v_48446 = v_48443 & v_48445;
assign v_48448 = v_48404 & v_48447;
assign v_48450 = v_45967;
assign v_48452 = v_48449 & v_48451;
assign v_48454 = v_48401 & v_48453;
assign v_48456 = v_45963;
assign v_48458 = v_48455 & v_48457;
assign v_48460 = v_48398 & v_48459;
assign v_48462 = v_45959;
assign v_48464 = v_48461 & v_48463;
assign v_48466 = v_48395 & v_48465;
assign v_48468 = v_45955;
assign v_48470 = v_48467 & v_48469;
assign v_48472 = v_48392 & v_48471;
assign v_48474 = v_45951;
assign v_48476 = v_48473 & v_48475;
assign v_48478 = v_48389 & v_48477;
assign v_48480 = v_45947;
assign v_48482 = v_48479 & v_48481;
assign v_48484 = v_48386 & v_48483;
assign v_48486 = v_45943;
assign v_48488 = v_48485 & v_48487;
assign v_48490 = v_48383 & v_48489;
assign v_48492 = v_45939;
assign v_48494 = v_48491 & v_48493;
assign v_48496 = v_48380 & v_48495;
assign v_48498 = v_2635;
assign v_48500 = v_48497 & v_48499;
assign v_48502 = v_48377 & v_48501;
assign v_48504 = v_2631;
assign v_48506 = v_48503 & v_48505;
assign v_48508 = v_48374 & v_48507;
assign v_48510 = v_2627;
assign v_48512 = v_48509 & v_48511;
assign v_48514 = v_48371 & v_48513;
assign v_48516 = v_2623;
assign v_48518 = v_48515 & v_48517;
assign v_48519 = v_48518;
assign v_48521 = v_45987;
assign v_48522 = v_2688;
assign v_48523 = v_48522;
assign v_48524 = v_48521 & v_48523;
assign v_48525 = v_48524;
assign v_48526 = v_48416 & v_48525;
assign v_48528 = v_48426 & v_48527;
assign v_48529 = v_48415 & v_48525;
assign v_48531 = v_48413 & v_48530;
assign v_48533 = v_48432 & v_48532;
assign v_48534 = v_48412 & v_48530;
assign v_48536 = v_48410 & v_48535;
assign v_48538 = v_48438 & v_48537;
assign v_48539 = v_48409 & v_48535;
assign v_48541 = v_48407 & v_48540;
assign v_48543 = v_48444 & v_48542;
assign v_48544 = v_48406 & v_48540;
assign v_48546 = v_48404 & v_48545;
assign v_48548 = v_48450 & v_48547;
assign v_48549 = v_48403 & v_48545;
assign v_48551 = v_48401 & v_48550;
assign v_48553 = v_48456 & v_48552;
assign v_48554 = v_48400 & v_48550;
assign v_48556 = v_48398 & v_48555;
assign v_48558 = v_48462 & v_48557;
assign v_48559 = v_48397 & v_48555;
assign v_48561 = v_48395 & v_48560;
assign v_48563 = v_48468 & v_48562;
assign v_48564 = v_48394 & v_48560;
assign v_48566 = v_48392 & v_48565;
assign v_48568 = v_48474 & v_48567;
assign v_48569 = v_48391 & v_48565;
assign v_48571 = v_48389 & v_48570;
assign v_48573 = v_48480 & v_48572;
assign v_48574 = v_48388 & v_48570;
assign v_48576 = v_48386 & v_48575;
assign v_48578 = v_48486 & v_48577;
assign v_48579 = v_48385 & v_48575;
assign v_48581 = v_48383 & v_48580;
assign v_48583 = v_48492 & v_48582;
assign v_48584 = v_48382 & v_48580;
assign v_48586 = v_48380 & v_48585;
assign v_48588 = v_48498 & v_48587;
assign v_48589 = v_48379 & v_48585;
assign v_48591 = v_48377 & v_48590;
assign v_48593 = v_48504 & v_48592;
assign v_48594 = v_48376 & v_48590;
assign v_48596 = v_48374 & v_48595;
assign v_48598 = v_48510 & v_48597;
assign v_48599 = v_48373 & v_48595;
assign v_48601 = v_48371 & v_48600;
assign v_48603 = v_48516 & v_48602;
assign v_48604 = v_48370 & v_48600;
assign v_48606 = v_48605;
assign v_48608 = v_48520 & v_48607;
assign v_48609 = v_48608;
assign v_48611 = v_48610;
assign v_48613 = ~v_2883;
assign v_48614 = ~v_45924;
assign v_48615 = v_45924;
assign v_48616 = ~v_2887;
assign v_48617 = ~v_45928;
assign v_48618 = v_45928;
assign v_48619 = ~v_2891;
assign v_48620 = ~v_45932;
assign v_48621 = v_45932;
assign v_48622 = ~v_2895;
assign v_48623 = ~v_45936;
assign v_48624 = v_45936;
assign v_48625 = ~v_45939;
assign v_48626 = ~v_2900;
assign v_48627 = v_2900;
assign v_48628 = ~v_45943;
assign v_48629 = ~v_2904;
assign v_48630 = v_2904;
assign v_48631 = ~v_45947;
assign v_48632 = ~v_2908;
assign v_48633 = v_2908;
assign v_48634 = ~v_45951;
assign v_48635 = ~v_2912;
assign v_48636 = v_2912;
assign v_48637 = ~v_45955;
assign v_48638 = ~v_2916;
assign v_48639 = v_2916;
assign v_48640 = ~v_45959;
assign v_48641 = ~v_2920;
assign v_48642 = v_2920;
assign v_48643 = ~v_45963;
assign v_48644 = ~v_2924;
assign v_48645 = v_2924;
assign v_48646 = ~v_45967;
assign v_48647 = ~v_2928;
assign v_48648 = v_2928;
assign v_48649 = ~v_45971;
assign v_48650 = ~v_2932;
assign v_48651 = v_2932;
assign v_48652 = ~v_45975;
assign v_48653 = ~v_2936;
assign v_48654 = v_2936;
assign v_48655 = ~v_45979;
assign v_48656 = ~v_2940;
assign v_48657 = v_2940;
assign v_48658 = ~v_45983;
assign v_48659 = ~v_2944;
assign v_48660 = v_2944;
assign v_48661 = ~v_45987;
assign v_48662 = ~v_2948;
assign v_48663 = v_48662;
assign v_48665 = v_48664;
assign v_48667 = v_48659 & v_48666;
assign v_48669 = v_45983;
assign v_48671 = v_48668 & v_48670;
assign v_48673 = v_48656 & v_48672;
assign v_48675 = v_45979;
assign v_48677 = v_48674 & v_48676;
assign v_48679 = v_48653 & v_48678;
assign v_48681 = v_45975;
assign v_48683 = v_48680 & v_48682;
assign v_48685 = v_48650 & v_48684;
assign v_48687 = v_45971;
assign v_48689 = v_48686 & v_48688;
assign v_48691 = v_48647 & v_48690;
assign v_48693 = v_45967;
assign v_48695 = v_48692 & v_48694;
assign v_48697 = v_48644 & v_48696;
assign v_48699 = v_45963;
assign v_48701 = v_48698 & v_48700;
assign v_48703 = v_48641 & v_48702;
assign v_48705 = v_45959;
assign v_48707 = v_48704 & v_48706;
assign v_48709 = v_48638 & v_48708;
assign v_48711 = v_45955;
assign v_48713 = v_48710 & v_48712;
assign v_48715 = v_48635 & v_48714;
assign v_48717 = v_45951;
assign v_48719 = v_48716 & v_48718;
assign v_48721 = v_48632 & v_48720;
assign v_48723 = v_45947;
assign v_48725 = v_48722 & v_48724;
assign v_48727 = v_48629 & v_48726;
assign v_48729 = v_45943;
assign v_48731 = v_48728 & v_48730;
assign v_48733 = v_48626 & v_48732;
assign v_48735 = v_45939;
assign v_48737 = v_48734 & v_48736;
assign v_48739 = v_48623 & v_48738;
assign v_48741 = v_2895;
assign v_48743 = v_48740 & v_48742;
assign v_48745 = v_48620 & v_48744;
assign v_48747 = v_2891;
assign v_48749 = v_48746 & v_48748;
assign v_48751 = v_48617 & v_48750;
assign v_48753 = v_2887;
assign v_48755 = v_48752 & v_48754;
assign v_48757 = v_48614 & v_48756;
assign v_48759 = v_2883;
assign v_48761 = v_48758 & v_48760;
assign v_48762 = v_48761;
assign v_48764 = v_45987;
assign v_48765 = v_2948;
assign v_48766 = v_48765;
assign v_48767 = v_48764 & v_48766;
assign v_48768 = v_48767;
assign v_48769 = v_48659 & v_48768;
assign v_48771 = v_48669 & v_48770;
assign v_48772 = v_48658 & v_48768;
assign v_48774 = v_48656 & v_48773;
assign v_48776 = v_48675 & v_48775;
assign v_48777 = v_48655 & v_48773;
assign v_48779 = v_48653 & v_48778;
assign v_48781 = v_48681 & v_48780;
assign v_48782 = v_48652 & v_48778;
assign v_48784 = v_48650 & v_48783;
assign v_48786 = v_48687 & v_48785;
assign v_48787 = v_48649 & v_48783;
assign v_48789 = v_48647 & v_48788;
assign v_48791 = v_48693 & v_48790;
assign v_48792 = v_48646 & v_48788;
assign v_48794 = v_48644 & v_48793;
assign v_48796 = v_48699 & v_48795;
assign v_48797 = v_48643 & v_48793;
assign v_48799 = v_48641 & v_48798;
assign v_48801 = v_48705 & v_48800;
assign v_48802 = v_48640 & v_48798;
assign v_48804 = v_48638 & v_48803;
assign v_48806 = v_48711 & v_48805;
assign v_48807 = v_48637 & v_48803;
assign v_48809 = v_48635 & v_48808;
assign v_48811 = v_48717 & v_48810;
assign v_48812 = v_48634 & v_48808;
assign v_48814 = v_48632 & v_48813;
assign v_48816 = v_48723 & v_48815;
assign v_48817 = v_48631 & v_48813;
assign v_48819 = v_48629 & v_48818;
assign v_48821 = v_48729 & v_48820;
assign v_48822 = v_48628 & v_48818;
assign v_48824 = v_48626 & v_48823;
assign v_48826 = v_48735 & v_48825;
assign v_48827 = v_48625 & v_48823;
assign v_48829 = v_48623 & v_48828;
assign v_48831 = v_48741 & v_48830;
assign v_48832 = v_48622 & v_48828;
assign v_48834 = v_48620 & v_48833;
assign v_48836 = v_48747 & v_48835;
assign v_48837 = v_48619 & v_48833;
assign v_48839 = v_48617 & v_48838;
assign v_48841 = v_48753 & v_48840;
assign v_48842 = v_48616 & v_48838;
assign v_48844 = v_48614 & v_48843;
assign v_48846 = v_48759 & v_48845;
assign v_48847 = v_48613 & v_48843;
assign v_48849 = v_48848;
assign v_48851 = v_48763 & v_48850;
assign v_48852 = v_48851;
assign v_48854 = v_48853;
assign v_48856 = ~v_3143;
assign v_48857 = ~v_45924;
assign v_48858 = v_45924;
assign v_48859 = ~v_3147;
assign v_48860 = ~v_45928;
assign v_48861 = v_45928;
assign v_48862 = ~v_3151;
assign v_48863 = ~v_45932;
assign v_48864 = v_45932;
assign v_48865 = ~v_3155;
assign v_48866 = ~v_45936;
assign v_48867 = v_45936;
assign v_48868 = ~v_45939;
assign v_48869 = ~v_3160;
assign v_48870 = v_3160;
assign v_48871 = ~v_45943;
assign v_48872 = ~v_3164;
assign v_48873 = v_3164;
assign v_48874 = ~v_45947;
assign v_48875 = ~v_3168;
assign v_48876 = v_3168;
assign v_48877 = ~v_45951;
assign v_48878 = ~v_3172;
assign v_48879 = v_3172;
assign v_48880 = ~v_45955;
assign v_48881 = ~v_3176;
assign v_48882 = v_3176;
assign v_48883 = ~v_45959;
assign v_48884 = ~v_3180;
assign v_48885 = v_3180;
assign v_48886 = ~v_45963;
assign v_48887 = ~v_3184;
assign v_48888 = v_3184;
assign v_48889 = ~v_45967;
assign v_48890 = ~v_3188;
assign v_48891 = v_3188;
assign v_48892 = ~v_45971;
assign v_48893 = ~v_3192;
assign v_48894 = v_3192;
assign v_48895 = ~v_45975;
assign v_48896 = ~v_3196;
assign v_48897 = v_3196;
assign v_48898 = ~v_45979;
assign v_48899 = ~v_3200;
assign v_48900 = v_3200;
assign v_48901 = ~v_45983;
assign v_48902 = ~v_3204;
assign v_48903 = v_3204;
assign v_48904 = ~v_45987;
assign v_48905 = ~v_3208;
assign v_48906 = v_48905;
assign v_48908 = v_48907;
assign v_48910 = v_48902 & v_48909;
assign v_48912 = v_45983;
assign v_48914 = v_48911 & v_48913;
assign v_48916 = v_48899 & v_48915;
assign v_48918 = v_45979;
assign v_48920 = v_48917 & v_48919;
assign v_48922 = v_48896 & v_48921;
assign v_48924 = v_45975;
assign v_48926 = v_48923 & v_48925;
assign v_48928 = v_48893 & v_48927;
assign v_48930 = v_45971;
assign v_48932 = v_48929 & v_48931;
assign v_48934 = v_48890 & v_48933;
assign v_48936 = v_45967;
assign v_48938 = v_48935 & v_48937;
assign v_48940 = v_48887 & v_48939;
assign v_48942 = v_45963;
assign v_48944 = v_48941 & v_48943;
assign v_48946 = v_48884 & v_48945;
assign v_48948 = v_45959;
assign v_48950 = v_48947 & v_48949;
assign v_48952 = v_48881 & v_48951;
assign v_48954 = v_45955;
assign v_48956 = v_48953 & v_48955;
assign v_48958 = v_48878 & v_48957;
assign v_48960 = v_45951;
assign v_48962 = v_48959 & v_48961;
assign v_48964 = v_48875 & v_48963;
assign v_48966 = v_45947;
assign v_48968 = v_48965 & v_48967;
assign v_48970 = v_48872 & v_48969;
assign v_48972 = v_45943;
assign v_48974 = v_48971 & v_48973;
assign v_48976 = v_48869 & v_48975;
assign v_48978 = v_45939;
assign v_48980 = v_48977 & v_48979;
assign v_48982 = v_48866 & v_48981;
assign v_48984 = v_3155;
assign v_48986 = v_48983 & v_48985;
assign v_48988 = v_48863 & v_48987;
assign v_48990 = v_3151;
assign v_48992 = v_48989 & v_48991;
assign v_48994 = v_48860 & v_48993;
assign v_48996 = v_3147;
assign v_48998 = v_48995 & v_48997;
assign v_49000 = v_48857 & v_48999;
assign v_49002 = v_3143;
assign v_49004 = v_49001 & v_49003;
assign v_49005 = v_49004;
assign v_49007 = v_45987;
assign v_49008 = v_3208;
assign v_49009 = v_49008;
assign v_49010 = v_49007 & v_49009;
assign v_49011 = v_49010;
assign v_49012 = v_48902 & v_49011;
assign v_49014 = v_48912 & v_49013;
assign v_49015 = v_48901 & v_49011;
assign v_49017 = v_48899 & v_49016;
assign v_49019 = v_48918 & v_49018;
assign v_49020 = v_48898 & v_49016;
assign v_49022 = v_48896 & v_49021;
assign v_49024 = v_48924 & v_49023;
assign v_49025 = v_48895 & v_49021;
assign v_49027 = v_48893 & v_49026;
assign v_49029 = v_48930 & v_49028;
assign v_49030 = v_48892 & v_49026;
assign v_49032 = v_48890 & v_49031;
assign v_49034 = v_48936 & v_49033;
assign v_49035 = v_48889 & v_49031;
assign v_49037 = v_48887 & v_49036;
assign v_49039 = v_48942 & v_49038;
assign v_49040 = v_48886 & v_49036;
assign v_49042 = v_48884 & v_49041;
assign v_49044 = v_48948 & v_49043;
assign v_49045 = v_48883 & v_49041;
assign v_49047 = v_48881 & v_49046;
assign v_49049 = v_48954 & v_49048;
assign v_49050 = v_48880 & v_49046;
assign v_49052 = v_48878 & v_49051;
assign v_49054 = v_48960 & v_49053;
assign v_49055 = v_48877 & v_49051;
assign v_49057 = v_48875 & v_49056;
assign v_49059 = v_48966 & v_49058;
assign v_49060 = v_48874 & v_49056;
assign v_49062 = v_48872 & v_49061;
assign v_49064 = v_48972 & v_49063;
assign v_49065 = v_48871 & v_49061;
assign v_49067 = v_48869 & v_49066;
assign v_49069 = v_48978 & v_49068;
assign v_49070 = v_48868 & v_49066;
assign v_49072 = v_48866 & v_49071;
assign v_49074 = v_48984 & v_49073;
assign v_49075 = v_48865 & v_49071;
assign v_49077 = v_48863 & v_49076;
assign v_49079 = v_48990 & v_49078;
assign v_49080 = v_48862 & v_49076;
assign v_49082 = v_48860 & v_49081;
assign v_49084 = v_48996 & v_49083;
assign v_49085 = v_48859 & v_49081;
assign v_49087 = v_48857 & v_49086;
assign v_49089 = v_49002 & v_49088;
assign v_49090 = v_48856 & v_49086;
assign v_49092 = v_49091;
assign v_49094 = v_49006 & v_49093;
assign v_49095 = v_49094;
assign v_49097 = v_49096;
assign v_49099 = ~v_3403;
assign v_49100 = ~v_45924;
assign v_49101 = v_45924;
assign v_49102 = ~v_3407;
assign v_49103 = ~v_45928;
assign v_49104 = v_45928;
assign v_49105 = ~v_3411;
assign v_49106 = ~v_45932;
assign v_49107 = v_45932;
assign v_49108 = ~v_3415;
assign v_49109 = ~v_45936;
assign v_49110 = v_45936;
assign v_49111 = ~v_45939;
assign v_49112 = ~v_3420;
assign v_49113 = v_3420;
assign v_49114 = ~v_45943;
assign v_49115 = ~v_3424;
assign v_49116 = v_3424;
assign v_49117 = ~v_45947;
assign v_49118 = ~v_3428;
assign v_49119 = v_3428;
assign v_49120 = ~v_45951;
assign v_49121 = ~v_3432;
assign v_49122 = v_3432;
assign v_49123 = ~v_45955;
assign v_49124 = ~v_3436;
assign v_49125 = v_3436;
assign v_49126 = ~v_45959;
assign v_49127 = ~v_3440;
assign v_49128 = v_3440;
assign v_49129 = ~v_45963;
assign v_49130 = ~v_3444;
assign v_49131 = v_3444;
assign v_49132 = ~v_45967;
assign v_49133 = ~v_3448;
assign v_49134 = v_3448;
assign v_49135 = ~v_45971;
assign v_49136 = ~v_3452;
assign v_49137 = v_3452;
assign v_49138 = ~v_45975;
assign v_49139 = ~v_3456;
assign v_49140 = v_3456;
assign v_49141 = ~v_45979;
assign v_49142 = ~v_3460;
assign v_49143 = v_3460;
assign v_49144 = ~v_45983;
assign v_49145 = ~v_3464;
assign v_49146 = v_3464;
assign v_49147 = ~v_45987;
assign v_49148 = ~v_3468;
assign v_49149 = v_49148;
assign v_49151 = v_49150;
assign v_49153 = v_49145 & v_49152;
assign v_49155 = v_45983;
assign v_49157 = v_49154 & v_49156;
assign v_49159 = v_49142 & v_49158;
assign v_49161 = v_45979;
assign v_49163 = v_49160 & v_49162;
assign v_49165 = v_49139 & v_49164;
assign v_49167 = v_45975;
assign v_49169 = v_49166 & v_49168;
assign v_49171 = v_49136 & v_49170;
assign v_49173 = v_45971;
assign v_49175 = v_49172 & v_49174;
assign v_49177 = v_49133 & v_49176;
assign v_49179 = v_45967;
assign v_49181 = v_49178 & v_49180;
assign v_49183 = v_49130 & v_49182;
assign v_49185 = v_45963;
assign v_49187 = v_49184 & v_49186;
assign v_49189 = v_49127 & v_49188;
assign v_49191 = v_45959;
assign v_49193 = v_49190 & v_49192;
assign v_49195 = v_49124 & v_49194;
assign v_49197 = v_45955;
assign v_49199 = v_49196 & v_49198;
assign v_49201 = v_49121 & v_49200;
assign v_49203 = v_45951;
assign v_49205 = v_49202 & v_49204;
assign v_49207 = v_49118 & v_49206;
assign v_49209 = v_45947;
assign v_49211 = v_49208 & v_49210;
assign v_49213 = v_49115 & v_49212;
assign v_49215 = v_45943;
assign v_49217 = v_49214 & v_49216;
assign v_49219 = v_49112 & v_49218;
assign v_49221 = v_45939;
assign v_49223 = v_49220 & v_49222;
assign v_49225 = v_49109 & v_49224;
assign v_49227 = v_3415;
assign v_49229 = v_49226 & v_49228;
assign v_49231 = v_49106 & v_49230;
assign v_49233 = v_3411;
assign v_49235 = v_49232 & v_49234;
assign v_49237 = v_49103 & v_49236;
assign v_49239 = v_3407;
assign v_49241 = v_49238 & v_49240;
assign v_49243 = v_49100 & v_49242;
assign v_49245 = v_3403;
assign v_49247 = v_49244 & v_49246;
assign v_49248 = v_49247;
assign v_49250 = v_45987;
assign v_49251 = v_3468;
assign v_49252 = v_49251;
assign v_49253 = v_49250 & v_49252;
assign v_49254 = v_49253;
assign v_49255 = v_49145 & v_49254;
assign v_49257 = v_49155 & v_49256;
assign v_49258 = v_49144 & v_49254;
assign v_49260 = v_49142 & v_49259;
assign v_49262 = v_49161 & v_49261;
assign v_49263 = v_49141 & v_49259;
assign v_49265 = v_49139 & v_49264;
assign v_49267 = v_49167 & v_49266;
assign v_49268 = v_49138 & v_49264;
assign v_49270 = v_49136 & v_49269;
assign v_49272 = v_49173 & v_49271;
assign v_49273 = v_49135 & v_49269;
assign v_49275 = v_49133 & v_49274;
assign v_49277 = v_49179 & v_49276;
assign v_49278 = v_49132 & v_49274;
assign v_49280 = v_49130 & v_49279;
assign v_49282 = v_49185 & v_49281;
assign v_49283 = v_49129 & v_49279;
assign v_49285 = v_49127 & v_49284;
assign v_49287 = v_49191 & v_49286;
assign v_49288 = v_49126 & v_49284;
assign v_49290 = v_49124 & v_49289;
assign v_49292 = v_49197 & v_49291;
assign v_49293 = v_49123 & v_49289;
assign v_49295 = v_49121 & v_49294;
assign v_49297 = v_49203 & v_49296;
assign v_49298 = v_49120 & v_49294;
assign v_49300 = v_49118 & v_49299;
assign v_49302 = v_49209 & v_49301;
assign v_49303 = v_49117 & v_49299;
assign v_49305 = v_49115 & v_49304;
assign v_49307 = v_49215 & v_49306;
assign v_49308 = v_49114 & v_49304;
assign v_49310 = v_49112 & v_49309;
assign v_49312 = v_49221 & v_49311;
assign v_49313 = v_49111 & v_49309;
assign v_49315 = v_49109 & v_49314;
assign v_49317 = v_49227 & v_49316;
assign v_49318 = v_49108 & v_49314;
assign v_49320 = v_49106 & v_49319;
assign v_49322 = v_49233 & v_49321;
assign v_49323 = v_49105 & v_49319;
assign v_49325 = v_49103 & v_49324;
assign v_49327 = v_49239 & v_49326;
assign v_49328 = v_49102 & v_49324;
assign v_49330 = v_49100 & v_49329;
assign v_49332 = v_49245 & v_49331;
assign v_49333 = v_49099 & v_49329;
assign v_49335 = v_49334;
assign v_49337 = v_49249 & v_49336;
assign v_49338 = v_49337;
assign v_49340 = v_49339;
assign v_49342 = ~v_3663;
assign v_49343 = ~v_45924;
assign v_49344 = v_45924;
assign v_49345 = ~v_3667;
assign v_49346 = ~v_45928;
assign v_49347 = v_45928;
assign v_49348 = ~v_3671;
assign v_49349 = ~v_45932;
assign v_49350 = v_45932;
assign v_49351 = ~v_3675;
assign v_49352 = ~v_45936;
assign v_49353 = v_45936;
assign v_49354 = ~v_45939;
assign v_49355 = ~v_3680;
assign v_49356 = v_3680;
assign v_49357 = ~v_45943;
assign v_49358 = ~v_3684;
assign v_49359 = v_3684;
assign v_49360 = ~v_45947;
assign v_49361 = ~v_3688;
assign v_49362 = v_3688;
assign v_49363 = ~v_45951;
assign v_49364 = ~v_3692;
assign v_49365 = v_3692;
assign v_49366 = ~v_45955;
assign v_49367 = ~v_3696;
assign v_49368 = v_3696;
assign v_49369 = ~v_45959;
assign v_49370 = ~v_3700;
assign v_49371 = v_3700;
assign v_49372 = ~v_45963;
assign v_49373 = ~v_3704;
assign v_49374 = v_3704;
assign v_49375 = ~v_45967;
assign v_49376 = ~v_3708;
assign v_49377 = v_3708;
assign v_49378 = ~v_45971;
assign v_49379 = ~v_3712;
assign v_49380 = v_3712;
assign v_49381 = ~v_45975;
assign v_49382 = ~v_3716;
assign v_49383 = v_3716;
assign v_49384 = ~v_45979;
assign v_49385 = ~v_3720;
assign v_49386 = v_3720;
assign v_49387 = ~v_45983;
assign v_49388 = ~v_3724;
assign v_49389 = v_3724;
assign v_49390 = ~v_45987;
assign v_49391 = ~v_3728;
assign v_49392 = v_49391;
assign v_49394 = v_49393;
assign v_49396 = v_49388 & v_49395;
assign v_49398 = v_45983;
assign v_49400 = v_49397 & v_49399;
assign v_49402 = v_49385 & v_49401;
assign v_49404 = v_45979;
assign v_49406 = v_49403 & v_49405;
assign v_49408 = v_49382 & v_49407;
assign v_49410 = v_45975;
assign v_49412 = v_49409 & v_49411;
assign v_49414 = v_49379 & v_49413;
assign v_49416 = v_45971;
assign v_49418 = v_49415 & v_49417;
assign v_49420 = v_49376 & v_49419;
assign v_49422 = v_45967;
assign v_49424 = v_49421 & v_49423;
assign v_49426 = v_49373 & v_49425;
assign v_49428 = v_45963;
assign v_49430 = v_49427 & v_49429;
assign v_49432 = v_49370 & v_49431;
assign v_49434 = v_45959;
assign v_49436 = v_49433 & v_49435;
assign v_49438 = v_49367 & v_49437;
assign v_49440 = v_45955;
assign v_49442 = v_49439 & v_49441;
assign v_49444 = v_49364 & v_49443;
assign v_49446 = v_45951;
assign v_49448 = v_49445 & v_49447;
assign v_49450 = v_49361 & v_49449;
assign v_49452 = v_45947;
assign v_49454 = v_49451 & v_49453;
assign v_49456 = v_49358 & v_49455;
assign v_49458 = v_45943;
assign v_49460 = v_49457 & v_49459;
assign v_49462 = v_49355 & v_49461;
assign v_49464 = v_45939;
assign v_49466 = v_49463 & v_49465;
assign v_49468 = v_49352 & v_49467;
assign v_49470 = v_3675;
assign v_49472 = v_49469 & v_49471;
assign v_49474 = v_49349 & v_49473;
assign v_49476 = v_3671;
assign v_49478 = v_49475 & v_49477;
assign v_49480 = v_49346 & v_49479;
assign v_49482 = v_3667;
assign v_49484 = v_49481 & v_49483;
assign v_49486 = v_49343 & v_49485;
assign v_49488 = v_3663;
assign v_49490 = v_49487 & v_49489;
assign v_49491 = v_49490;
assign v_49493 = v_45987;
assign v_49494 = v_3728;
assign v_49495 = v_49494;
assign v_49496 = v_49493 & v_49495;
assign v_49497 = v_49496;
assign v_49498 = v_49388 & v_49497;
assign v_49500 = v_49398 & v_49499;
assign v_49501 = v_49387 & v_49497;
assign v_49503 = v_49385 & v_49502;
assign v_49505 = v_49404 & v_49504;
assign v_49506 = v_49384 & v_49502;
assign v_49508 = v_49382 & v_49507;
assign v_49510 = v_49410 & v_49509;
assign v_49511 = v_49381 & v_49507;
assign v_49513 = v_49379 & v_49512;
assign v_49515 = v_49416 & v_49514;
assign v_49516 = v_49378 & v_49512;
assign v_49518 = v_49376 & v_49517;
assign v_49520 = v_49422 & v_49519;
assign v_49521 = v_49375 & v_49517;
assign v_49523 = v_49373 & v_49522;
assign v_49525 = v_49428 & v_49524;
assign v_49526 = v_49372 & v_49522;
assign v_49528 = v_49370 & v_49527;
assign v_49530 = v_49434 & v_49529;
assign v_49531 = v_49369 & v_49527;
assign v_49533 = v_49367 & v_49532;
assign v_49535 = v_49440 & v_49534;
assign v_49536 = v_49366 & v_49532;
assign v_49538 = v_49364 & v_49537;
assign v_49540 = v_49446 & v_49539;
assign v_49541 = v_49363 & v_49537;
assign v_49543 = v_49361 & v_49542;
assign v_49545 = v_49452 & v_49544;
assign v_49546 = v_49360 & v_49542;
assign v_49548 = v_49358 & v_49547;
assign v_49550 = v_49458 & v_49549;
assign v_49551 = v_49357 & v_49547;
assign v_49553 = v_49355 & v_49552;
assign v_49555 = v_49464 & v_49554;
assign v_49556 = v_49354 & v_49552;
assign v_49558 = v_49352 & v_49557;
assign v_49560 = v_49470 & v_49559;
assign v_49561 = v_49351 & v_49557;
assign v_49563 = v_49349 & v_49562;
assign v_49565 = v_49476 & v_49564;
assign v_49566 = v_49348 & v_49562;
assign v_49568 = v_49346 & v_49567;
assign v_49570 = v_49482 & v_49569;
assign v_49571 = v_49345 & v_49567;
assign v_49573 = v_49343 & v_49572;
assign v_49575 = v_49488 & v_49574;
assign v_49576 = v_49342 & v_49572;
assign v_49578 = v_49577;
assign v_49580 = v_49492 & v_49579;
assign v_49581 = v_49580;
assign v_49583 = v_49582;
assign v_49585 = ~v_3923;
assign v_49586 = ~v_45924;
assign v_49587 = v_45924;
assign v_49588 = ~v_3927;
assign v_49589 = ~v_45928;
assign v_49590 = v_45928;
assign v_49591 = ~v_3931;
assign v_49592 = ~v_45932;
assign v_49593 = v_45932;
assign v_49594 = ~v_3935;
assign v_49595 = ~v_45936;
assign v_49596 = v_45936;
assign v_49597 = ~v_45939;
assign v_49598 = ~v_3940;
assign v_49599 = v_3940;
assign v_49600 = ~v_45943;
assign v_49601 = ~v_3944;
assign v_49602 = v_3944;
assign v_49603 = ~v_45947;
assign v_49604 = ~v_3948;
assign v_49605 = v_3948;
assign v_49606 = ~v_45951;
assign v_49607 = ~v_3952;
assign v_49608 = v_3952;
assign v_49609 = ~v_45955;
assign v_49610 = ~v_3956;
assign v_49611 = v_3956;
assign v_49612 = ~v_45959;
assign v_49613 = ~v_3960;
assign v_49614 = v_3960;
assign v_49615 = ~v_45963;
assign v_49616 = ~v_3964;
assign v_49617 = v_3964;
assign v_49618 = ~v_45967;
assign v_49619 = ~v_3968;
assign v_49620 = v_3968;
assign v_49621 = ~v_45971;
assign v_49622 = ~v_3972;
assign v_49623 = v_3972;
assign v_49624 = ~v_45975;
assign v_49625 = ~v_3976;
assign v_49626 = v_3976;
assign v_49627 = ~v_45979;
assign v_49628 = ~v_3980;
assign v_49629 = v_3980;
assign v_49630 = ~v_45983;
assign v_49631 = ~v_3984;
assign v_49632 = v_3984;
assign v_49633 = ~v_45987;
assign v_49634 = ~v_3988;
assign v_49635 = v_49634;
assign v_49637 = v_49636;
assign v_49639 = v_49631 & v_49638;
assign v_49641 = v_45983;
assign v_49643 = v_49640 & v_49642;
assign v_49645 = v_49628 & v_49644;
assign v_49647 = v_45979;
assign v_49649 = v_49646 & v_49648;
assign v_49651 = v_49625 & v_49650;
assign v_49653 = v_45975;
assign v_49655 = v_49652 & v_49654;
assign v_49657 = v_49622 & v_49656;
assign v_49659 = v_45971;
assign v_49661 = v_49658 & v_49660;
assign v_49663 = v_49619 & v_49662;
assign v_49665 = v_45967;
assign v_49667 = v_49664 & v_49666;
assign v_49669 = v_49616 & v_49668;
assign v_49671 = v_45963;
assign v_49673 = v_49670 & v_49672;
assign v_49675 = v_49613 & v_49674;
assign v_49677 = v_45959;
assign v_49679 = v_49676 & v_49678;
assign v_49681 = v_49610 & v_49680;
assign v_49683 = v_45955;
assign v_49685 = v_49682 & v_49684;
assign v_49687 = v_49607 & v_49686;
assign v_49689 = v_45951;
assign v_49691 = v_49688 & v_49690;
assign v_49693 = v_49604 & v_49692;
assign v_49695 = v_45947;
assign v_49697 = v_49694 & v_49696;
assign v_49699 = v_49601 & v_49698;
assign v_49701 = v_45943;
assign v_49703 = v_49700 & v_49702;
assign v_49705 = v_49598 & v_49704;
assign v_49707 = v_45939;
assign v_49709 = v_49706 & v_49708;
assign v_49711 = v_49595 & v_49710;
assign v_49713 = v_3935;
assign v_49715 = v_49712 & v_49714;
assign v_49717 = v_49592 & v_49716;
assign v_49719 = v_3931;
assign v_49721 = v_49718 & v_49720;
assign v_49723 = v_49589 & v_49722;
assign v_49725 = v_3927;
assign v_49727 = v_49724 & v_49726;
assign v_49729 = v_49586 & v_49728;
assign v_49731 = v_3923;
assign v_49733 = v_49730 & v_49732;
assign v_49734 = v_49733;
assign v_49736 = v_45987;
assign v_49737 = v_3988;
assign v_49738 = v_49737;
assign v_49739 = v_49736 & v_49738;
assign v_49740 = v_49739;
assign v_49741 = v_49631 & v_49740;
assign v_49743 = v_49641 & v_49742;
assign v_49744 = v_49630 & v_49740;
assign v_49746 = v_49628 & v_49745;
assign v_49748 = v_49647 & v_49747;
assign v_49749 = v_49627 & v_49745;
assign v_49751 = v_49625 & v_49750;
assign v_49753 = v_49653 & v_49752;
assign v_49754 = v_49624 & v_49750;
assign v_49756 = v_49622 & v_49755;
assign v_49758 = v_49659 & v_49757;
assign v_49759 = v_49621 & v_49755;
assign v_49761 = v_49619 & v_49760;
assign v_49763 = v_49665 & v_49762;
assign v_49764 = v_49618 & v_49760;
assign v_49766 = v_49616 & v_49765;
assign v_49768 = v_49671 & v_49767;
assign v_49769 = v_49615 & v_49765;
assign v_49771 = v_49613 & v_49770;
assign v_49773 = v_49677 & v_49772;
assign v_49774 = v_49612 & v_49770;
assign v_49776 = v_49610 & v_49775;
assign v_49778 = v_49683 & v_49777;
assign v_49779 = v_49609 & v_49775;
assign v_49781 = v_49607 & v_49780;
assign v_49783 = v_49689 & v_49782;
assign v_49784 = v_49606 & v_49780;
assign v_49786 = v_49604 & v_49785;
assign v_49788 = v_49695 & v_49787;
assign v_49789 = v_49603 & v_49785;
assign v_49791 = v_49601 & v_49790;
assign v_49793 = v_49701 & v_49792;
assign v_49794 = v_49600 & v_49790;
assign v_49796 = v_49598 & v_49795;
assign v_49798 = v_49707 & v_49797;
assign v_49799 = v_49597 & v_49795;
assign v_49801 = v_49595 & v_49800;
assign v_49803 = v_49713 & v_49802;
assign v_49804 = v_49594 & v_49800;
assign v_49806 = v_49592 & v_49805;
assign v_49808 = v_49719 & v_49807;
assign v_49809 = v_49591 & v_49805;
assign v_49811 = v_49589 & v_49810;
assign v_49813 = v_49725 & v_49812;
assign v_49814 = v_49588 & v_49810;
assign v_49816 = v_49586 & v_49815;
assign v_49818 = v_49731 & v_49817;
assign v_49819 = v_49585 & v_49815;
assign v_49821 = v_49820;
assign v_49823 = v_49735 & v_49822;
assign v_49824 = v_49823;
assign v_49826 = v_49825;
assign v_49827 = ~v_4182;
assign v_49828 = ~v_45924;
assign v_49829 = v_45924;
assign v_49830 = ~v_4186;
assign v_49831 = ~v_45928;
assign v_49832 = v_45928;
assign v_49833 = ~v_4190;
assign v_49834 = ~v_45932;
assign v_49835 = v_45932;
assign v_49836 = ~v_4194;
assign v_49837 = ~v_45936;
assign v_49838 = v_45936;
assign v_49839 = ~v_45939;
assign v_49840 = ~v_4199;
assign v_49841 = v_4199;
assign v_49842 = ~v_45943;
assign v_49843 = ~v_4203;
assign v_49844 = v_4203;
assign v_49845 = ~v_45947;
assign v_49846 = ~v_4207;
assign v_49847 = v_4207;
assign v_49848 = ~v_45951;
assign v_49849 = ~v_4211;
assign v_49850 = v_4211;
assign v_49851 = ~v_45955;
assign v_49852 = ~v_4215;
assign v_49853 = v_4215;
assign v_49854 = ~v_45959;
assign v_49855 = ~v_4219;
assign v_49856 = v_4219;
assign v_49857 = ~v_45963;
assign v_49858 = ~v_4223;
assign v_49859 = v_4223;
assign v_49860 = ~v_45967;
assign v_49861 = ~v_4227;
assign v_49862 = v_4227;
assign v_49863 = ~v_45971;
assign v_49864 = ~v_4231;
assign v_49865 = v_4231;
assign v_49866 = ~v_45975;
assign v_49867 = ~v_4235;
assign v_49868 = v_4235;
assign v_49869 = ~v_45979;
assign v_49870 = ~v_4239;
assign v_49871 = v_4239;
assign v_49872 = ~v_45983;
assign v_49873 = ~v_4243;
assign v_49874 = v_4243;
assign v_49875 = ~v_45987;
assign v_49876 = ~v_4247;
assign v_49877 = v_49876;
assign v_49879 = v_49878;
assign v_49881 = v_49873 & v_49880;
assign v_49883 = v_45983;
assign v_49885 = v_49882 & v_49884;
assign v_49887 = v_49870 & v_49886;
assign v_49889 = v_45979;
assign v_49891 = v_49888 & v_49890;
assign v_49893 = v_49867 & v_49892;
assign v_49895 = v_45975;
assign v_49897 = v_49894 & v_49896;
assign v_49899 = v_49864 & v_49898;
assign v_49901 = v_45971;
assign v_49903 = v_49900 & v_49902;
assign v_49905 = v_49861 & v_49904;
assign v_49907 = v_45967;
assign v_49909 = v_49906 & v_49908;
assign v_49911 = v_49858 & v_49910;
assign v_49913 = v_45963;
assign v_49915 = v_49912 & v_49914;
assign v_49917 = v_49855 & v_49916;
assign v_49919 = v_45959;
assign v_49921 = v_49918 & v_49920;
assign v_49923 = v_49852 & v_49922;
assign v_49925 = v_45955;
assign v_49927 = v_49924 & v_49926;
assign v_49929 = v_49849 & v_49928;
assign v_49931 = v_45951;
assign v_49933 = v_49930 & v_49932;
assign v_49935 = v_49846 & v_49934;
assign v_49937 = v_45947;
assign v_49939 = v_49936 & v_49938;
assign v_49941 = v_49843 & v_49940;
assign v_49943 = v_45943;
assign v_49945 = v_49942 & v_49944;
assign v_49947 = v_49840 & v_49946;
assign v_49949 = v_45939;
assign v_49951 = v_49948 & v_49950;
assign v_49953 = v_49837 & v_49952;
assign v_49955 = v_4194;
assign v_49957 = v_49954 & v_49956;
assign v_49959 = v_49834 & v_49958;
assign v_49961 = v_4190;
assign v_49963 = v_49960 & v_49962;
assign v_49965 = v_49831 & v_49964;
assign v_49967 = v_4186;
assign v_49969 = v_49966 & v_49968;
assign v_49971 = v_49828 & v_49970;
assign v_49973 = v_4182;
assign v_49975 = v_49972 & v_49974;
assign v_49977 = ~v_49976;
assign v_49979 = v_45987;
assign v_49980 = v_4247;
assign v_49981 = v_49980;
assign v_49982 = v_49979 & v_49981;
assign v_49983 = v_49982;
assign v_49984 = v_49873 & v_49983;
assign v_49986 = v_49883 & v_49985;
assign v_49987 = v_49872 & v_49983;
assign v_49989 = v_49870 & v_49988;
assign v_49991 = v_49889 & v_49990;
assign v_49992 = v_49869 & v_49988;
assign v_49994 = v_49867 & v_49993;
assign v_49996 = v_49895 & v_49995;
assign v_49997 = v_49866 & v_49993;
assign v_49999 = v_49864 & v_49998;
assign v_50001 = v_49901 & v_50000;
assign v_50002 = v_49863 & v_49998;
assign v_50004 = v_49861 & v_50003;
assign v_50006 = v_49907 & v_50005;
assign v_50007 = v_49860 & v_50003;
assign v_50009 = v_49858 & v_50008;
assign v_50011 = v_49913 & v_50010;
assign v_50012 = v_49857 & v_50008;
assign v_50014 = v_49855 & v_50013;
assign v_50016 = v_49919 & v_50015;
assign v_50017 = v_49854 & v_50013;
assign v_50019 = v_49852 & v_50018;
assign v_50021 = v_49925 & v_50020;
assign v_50022 = v_49851 & v_50018;
assign v_50024 = v_49849 & v_50023;
assign v_50026 = v_49931 & v_50025;
assign v_50027 = v_49848 & v_50023;
assign v_50029 = v_49846 & v_50028;
assign v_50031 = v_49937 & v_50030;
assign v_50032 = v_49845 & v_50028;
assign v_50034 = v_49843 & v_50033;
assign v_50036 = v_49943 & v_50035;
assign v_50037 = v_49842 & v_50033;
assign v_50039 = v_49840 & v_50038;
assign v_50041 = v_49949 & v_50040;
assign v_50042 = v_49839 & v_50038;
assign v_50044 = v_49837 & v_50043;
assign v_50046 = v_49955 & v_50045;
assign v_50047 = v_49836 & v_50043;
assign v_50049 = v_49834 & v_50048;
assign v_50051 = v_49961 & v_50050;
assign v_50052 = v_49833 & v_50048;
assign v_50054 = v_49831 & v_50053;
assign v_50056 = v_49967 & v_50055;
assign v_50057 = v_49830 & v_50053;
assign v_50059 = v_49828 & v_50058;
assign v_50061 = v_49973 & v_50060;
assign v_50062 = v_49827 & v_50058;
assign v_50064 = v_49976;
assign v_50066 = v_49978 & v_50065;
assign v_50067 = v_50066;
assign v_50069 = v_50068;
assign v_50071 = ~v_6;
assign v_50073 = ~v_50072;
assign v_50074 = v_50072;
assign v_50075 = ~v_13;
assign v_50077 = ~v_50076;
assign v_50078 = v_50076;
assign v_50079 = ~v_18;
assign v_50081 = ~v_50080;
assign v_50082 = v_50080;
assign v_50083 = ~v_23;
assign v_50085 = ~v_50084;
assign v_50086 = v_50084;
assign v_50088 = ~v_50087;
assign v_50089 = ~v_30;
assign v_50090 = v_30;
assign v_50092 = ~v_50091;
assign v_50093 = ~v_35;
assign v_50094 = v_35;
assign v_50096 = ~v_50095;
assign v_50097 = ~v_40;
assign v_50098 = v_40;
assign v_50100 = ~v_50099;
assign v_50101 = ~v_45;
assign v_50102 = v_45;
assign v_50104 = ~v_50103;
assign v_50105 = ~v_50;
assign v_50106 = v_50;
assign v_50108 = ~v_50107;
assign v_50109 = ~v_55;
assign v_50110 = v_55;
assign v_50112 = ~v_50111;
assign v_50113 = ~v_60;
assign v_50114 = v_60;
assign v_50116 = ~v_50115;
assign v_50117 = ~v_65;
assign v_50118 = v_65;
assign v_50120 = ~v_50119;
assign v_50121 = ~v_70;
assign v_50122 = v_70;
assign v_50124 = ~v_50123;
assign v_50125 = ~v_75;
assign v_50126 = v_75;
assign v_50128 = ~v_50127;
assign v_50129 = ~v_80;
assign v_50130 = v_80;
assign v_50132 = ~v_50131;
assign v_50133 = ~v_85;
assign v_50134 = v_85;
assign v_50136 = ~v_50135;
assign v_50137 = ~v_90;
assign v_50138 = v_50137;
assign v_50140 = v_50139;
assign v_50142 = v_50133 & v_50141;
assign v_50144 = v_50131;
assign v_50146 = v_50143 & v_50145;
assign v_50148 = v_50129 & v_50147;
assign v_50150 = v_50127;
assign v_50152 = v_50149 & v_50151;
assign v_50154 = v_50125 & v_50153;
assign v_50156 = v_50123;
assign v_50158 = v_50155 & v_50157;
assign v_50160 = v_50121 & v_50159;
assign v_50162 = v_50119;
assign v_50164 = v_50161 & v_50163;
assign v_50166 = v_50117 & v_50165;
assign v_50168 = v_50115;
assign v_50170 = v_50167 & v_50169;
assign v_50172 = v_50113 & v_50171;
assign v_50174 = v_50111;
assign v_50176 = v_50173 & v_50175;
assign v_50178 = v_50109 & v_50177;
assign v_50180 = v_50107;
assign v_50182 = v_50179 & v_50181;
assign v_50184 = v_50105 & v_50183;
assign v_50186 = v_50103;
assign v_50188 = v_50185 & v_50187;
assign v_50190 = v_50101 & v_50189;
assign v_50192 = v_50099;
assign v_50194 = v_50191 & v_50193;
assign v_50196 = v_50097 & v_50195;
assign v_50198 = v_50095;
assign v_50200 = v_50197 & v_50199;
assign v_50202 = v_50093 & v_50201;
assign v_50204 = v_50091;
assign v_50206 = v_50203 & v_50205;
assign v_50208 = v_50089 & v_50207;
assign v_50210 = v_50087;
assign v_50212 = v_50209 & v_50211;
assign v_50214 = v_50085 & v_50213;
assign v_50216 = v_23;
assign v_50218 = v_50215 & v_50217;
assign v_50220 = v_50081 & v_50219;
assign v_50222 = v_18;
assign v_50224 = v_50221 & v_50223;
assign v_50226 = v_50077 & v_50225;
assign v_50228 = v_13;
assign v_50230 = v_50227 & v_50229;
assign v_50232 = v_50073 & v_50231;
assign v_50234 = v_6;
assign v_50236 = v_50233 & v_50235;
assign v_50237 = v_50236;
assign v_50239 = v_50135;
assign v_50240 = v_90;
assign v_50241 = v_50240;
assign v_50242 = v_50239 & v_50241;
assign v_50243 = v_50242;
assign v_50244 = v_50133 & v_50243;
assign v_50246 = v_50144 & v_50245;
assign v_50247 = v_50132 & v_50243;
assign v_50249 = v_50129 & v_50248;
assign v_50251 = v_50150 & v_50250;
assign v_50252 = v_50128 & v_50248;
assign v_50254 = v_50125 & v_50253;
assign v_50256 = v_50156 & v_50255;
assign v_50257 = v_50124 & v_50253;
assign v_50259 = v_50121 & v_50258;
assign v_50261 = v_50162 & v_50260;
assign v_50262 = v_50120 & v_50258;
assign v_50264 = v_50117 & v_50263;
assign v_50266 = v_50168 & v_50265;
assign v_50267 = v_50116 & v_50263;
assign v_50269 = v_50113 & v_50268;
assign v_50271 = v_50174 & v_50270;
assign v_50272 = v_50112 & v_50268;
assign v_50274 = v_50109 & v_50273;
assign v_50276 = v_50180 & v_50275;
assign v_50277 = v_50108 & v_50273;
assign v_50279 = v_50105 & v_50278;
assign v_50281 = v_50186 & v_50280;
assign v_50282 = v_50104 & v_50278;
assign v_50284 = v_50101 & v_50283;
assign v_50286 = v_50192 & v_50285;
assign v_50287 = v_50100 & v_50283;
assign v_50289 = v_50097 & v_50288;
assign v_50291 = v_50198 & v_50290;
assign v_50292 = v_50096 & v_50288;
assign v_50294 = v_50093 & v_50293;
assign v_50296 = v_50204 & v_50295;
assign v_50297 = v_50092 & v_50293;
assign v_50299 = v_50089 & v_50298;
assign v_50301 = v_50210 & v_50300;
assign v_50302 = v_50088 & v_50298;
assign v_50304 = v_50085 & v_50303;
assign v_50306 = v_50216 & v_50305;
assign v_50307 = v_50083 & v_50303;
assign v_50309 = v_50081 & v_50308;
assign v_50311 = v_50222 & v_50310;
assign v_50312 = v_50079 & v_50308;
assign v_50314 = v_50077 & v_50313;
assign v_50316 = v_50228 & v_50315;
assign v_50317 = v_50075 & v_50313;
assign v_50319 = v_50073 & v_50318;
assign v_50321 = v_50234 & v_50320;
assign v_50322 = v_50071 & v_50318;
assign v_50324 = v_50323;
assign v_50326 = v_50238 & v_50325;
assign v_50327 = v_50326;
assign v_50329 = v_50328;
assign v_50331 = ~v_283;
assign v_50332 = ~v_50072;
assign v_50333 = v_50072;
assign v_50334 = ~v_287;
assign v_50335 = ~v_50076;
assign v_50336 = v_50076;
assign v_50337 = ~v_291;
assign v_50338 = ~v_50080;
assign v_50339 = v_50080;
assign v_50340 = ~v_295;
assign v_50341 = ~v_50084;
assign v_50342 = v_50084;
assign v_50343 = ~v_50087;
assign v_50344 = ~v_300;
assign v_50345 = v_300;
assign v_50346 = ~v_50091;
assign v_50347 = ~v_304;
assign v_50348 = v_304;
assign v_50349 = ~v_50095;
assign v_50350 = ~v_308;
assign v_50351 = v_308;
assign v_50352 = ~v_50099;
assign v_50353 = ~v_312;
assign v_50354 = v_312;
assign v_50355 = ~v_50103;
assign v_50356 = ~v_316;
assign v_50357 = v_316;
assign v_50358 = ~v_50107;
assign v_50359 = ~v_320;
assign v_50360 = v_320;
assign v_50361 = ~v_50111;
assign v_50362 = ~v_324;
assign v_50363 = v_324;
assign v_50364 = ~v_50115;
assign v_50365 = ~v_328;
assign v_50366 = v_328;
assign v_50367 = ~v_50119;
assign v_50368 = ~v_332;
assign v_50369 = v_332;
assign v_50370 = ~v_50123;
assign v_50371 = ~v_336;
assign v_50372 = v_336;
assign v_50373 = ~v_50127;
assign v_50374 = ~v_340;
assign v_50375 = v_340;
assign v_50376 = ~v_50131;
assign v_50377 = ~v_344;
assign v_50378 = v_344;
assign v_50379 = ~v_50135;
assign v_50380 = ~v_348;
assign v_50381 = v_50380;
assign v_50383 = v_50382;
assign v_50385 = v_50377 & v_50384;
assign v_50387 = v_50131;
assign v_50389 = v_50386 & v_50388;
assign v_50391 = v_50374 & v_50390;
assign v_50393 = v_50127;
assign v_50395 = v_50392 & v_50394;
assign v_50397 = v_50371 & v_50396;
assign v_50399 = v_50123;
assign v_50401 = v_50398 & v_50400;
assign v_50403 = v_50368 & v_50402;
assign v_50405 = v_50119;
assign v_50407 = v_50404 & v_50406;
assign v_50409 = v_50365 & v_50408;
assign v_50411 = v_50115;
assign v_50413 = v_50410 & v_50412;
assign v_50415 = v_50362 & v_50414;
assign v_50417 = v_50111;
assign v_50419 = v_50416 & v_50418;
assign v_50421 = v_50359 & v_50420;
assign v_50423 = v_50107;
assign v_50425 = v_50422 & v_50424;
assign v_50427 = v_50356 & v_50426;
assign v_50429 = v_50103;
assign v_50431 = v_50428 & v_50430;
assign v_50433 = v_50353 & v_50432;
assign v_50435 = v_50099;
assign v_50437 = v_50434 & v_50436;
assign v_50439 = v_50350 & v_50438;
assign v_50441 = v_50095;
assign v_50443 = v_50440 & v_50442;
assign v_50445 = v_50347 & v_50444;
assign v_50447 = v_50091;
assign v_50449 = v_50446 & v_50448;
assign v_50451 = v_50344 & v_50450;
assign v_50453 = v_50087;
assign v_50455 = v_50452 & v_50454;
assign v_50457 = v_50341 & v_50456;
assign v_50459 = v_295;
assign v_50461 = v_50458 & v_50460;
assign v_50463 = v_50338 & v_50462;
assign v_50465 = v_291;
assign v_50467 = v_50464 & v_50466;
assign v_50469 = v_50335 & v_50468;
assign v_50471 = v_287;
assign v_50473 = v_50470 & v_50472;
assign v_50475 = v_50332 & v_50474;
assign v_50477 = v_283;
assign v_50479 = v_50476 & v_50478;
assign v_50480 = v_50479;
assign v_50482 = v_50135;
assign v_50483 = v_348;
assign v_50484 = v_50483;
assign v_50485 = v_50482 & v_50484;
assign v_50486 = v_50485;
assign v_50487 = v_50377 & v_50486;
assign v_50489 = v_50387 & v_50488;
assign v_50490 = v_50376 & v_50486;
assign v_50492 = v_50374 & v_50491;
assign v_50494 = v_50393 & v_50493;
assign v_50495 = v_50373 & v_50491;
assign v_50497 = v_50371 & v_50496;
assign v_50499 = v_50399 & v_50498;
assign v_50500 = v_50370 & v_50496;
assign v_50502 = v_50368 & v_50501;
assign v_50504 = v_50405 & v_50503;
assign v_50505 = v_50367 & v_50501;
assign v_50507 = v_50365 & v_50506;
assign v_50509 = v_50411 & v_50508;
assign v_50510 = v_50364 & v_50506;
assign v_50512 = v_50362 & v_50511;
assign v_50514 = v_50417 & v_50513;
assign v_50515 = v_50361 & v_50511;
assign v_50517 = v_50359 & v_50516;
assign v_50519 = v_50423 & v_50518;
assign v_50520 = v_50358 & v_50516;
assign v_50522 = v_50356 & v_50521;
assign v_50524 = v_50429 & v_50523;
assign v_50525 = v_50355 & v_50521;
assign v_50527 = v_50353 & v_50526;
assign v_50529 = v_50435 & v_50528;
assign v_50530 = v_50352 & v_50526;
assign v_50532 = v_50350 & v_50531;
assign v_50534 = v_50441 & v_50533;
assign v_50535 = v_50349 & v_50531;
assign v_50537 = v_50347 & v_50536;
assign v_50539 = v_50447 & v_50538;
assign v_50540 = v_50346 & v_50536;
assign v_50542 = v_50344 & v_50541;
assign v_50544 = v_50453 & v_50543;
assign v_50545 = v_50343 & v_50541;
assign v_50547 = v_50341 & v_50546;
assign v_50549 = v_50459 & v_50548;
assign v_50550 = v_50340 & v_50546;
assign v_50552 = v_50338 & v_50551;
assign v_50554 = v_50465 & v_50553;
assign v_50555 = v_50337 & v_50551;
assign v_50557 = v_50335 & v_50556;
assign v_50559 = v_50471 & v_50558;
assign v_50560 = v_50334 & v_50556;
assign v_50562 = v_50332 & v_50561;
assign v_50564 = v_50477 & v_50563;
assign v_50565 = v_50331 & v_50561;
assign v_50567 = v_50566;
assign v_50569 = v_50481 & v_50568;
assign v_50570 = v_50569;
assign v_50572 = v_50571;
assign v_50574 = ~v_543;
assign v_50575 = ~v_50072;
assign v_50576 = v_50072;
assign v_50577 = ~v_547;
assign v_50578 = ~v_50076;
assign v_50579 = v_50076;
assign v_50580 = ~v_551;
assign v_50581 = ~v_50080;
assign v_50582 = v_50080;
assign v_50583 = ~v_555;
assign v_50584 = ~v_50084;
assign v_50585 = v_50084;
assign v_50586 = ~v_50087;
assign v_50587 = ~v_560;
assign v_50588 = v_560;
assign v_50589 = ~v_50091;
assign v_50590 = ~v_564;
assign v_50591 = v_564;
assign v_50592 = ~v_50095;
assign v_50593 = ~v_568;
assign v_50594 = v_568;
assign v_50595 = ~v_50099;
assign v_50596 = ~v_572;
assign v_50597 = v_572;
assign v_50598 = ~v_50103;
assign v_50599 = ~v_576;
assign v_50600 = v_576;
assign v_50601 = ~v_50107;
assign v_50602 = ~v_580;
assign v_50603 = v_580;
assign v_50604 = ~v_50111;
assign v_50605 = ~v_584;
assign v_50606 = v_584;
assign v_50607 = ~v_50115;
assign v_50608 = ~v_588;
assign v_50609 = v_588;
assign v_50610 = ~v_50119;
assign v_50611 = ~v_592;
assign v_50612 = v_592;
assign v_50613 = ~v_50123;
assign v_50614 = ~v_596;
assign v_50615 = v_596;
assign v_50616 = ~v_50127;
assign v_50617 = ~v_600;
assign v_50618 = v_600;
assign v_50619 = ~v_50131;
assign v_50620 = ~v_604;
assign v_50621 = v_604;
assign v_50622 = ~v_50135;
assign v_50623 = ~v_608;
assign v_50624 = v_50623;
assign v_50626 = v_50625;
assign v_50628 = v_50620 & v_50627;
assign v_50630 = v_50131;
assign v_50632 = v_50629 & v_50631;
assign v_50634 = v_50617 & v_50633;
assign v_50636 = v_50127;
assign v_50638 = v_50635 & v_50637;
assign v_50640 = v_50614 & v_50639;
assign v_50642 = v_50123;
assign v_50644 = v_50641 & v_50643;
assign v_50646 = v_50611 & v_50645;
assign v_50648 = v_50119;
assign v_50650 = v_50647 & v_50649;
assign v_50652 = v_50608 & v_50651;
assign v_50654 = v_50115;
assign v_50656 = v_50653 & v_50655;
assign v_50658 = v_50605 & v_50657;
assign v_50660 = v_50111;
assign v_50662 = v_50659 & v_50661;
assign v_50664 = v_50602 & v_50663;
assign v_50666 = v_50107;
assign v_50668 = v_50665 & v_50667;
assign v_50670 = v_50599 & v_50669;
assign v_50672 = v_50103;
assign v_50674 = v_50671 & v_50673;
assign v_50676 = v_50596 & v_50675;
assign v_50678 = v_50099;
assign v_50680 = v_50677 & v_50679;
assign v_50682 = v_50593 & v_50681;
assign v_50684 = v_50095;
assign v_50686 = v_50683 & v_50685;
assign v_50688 = v_50590 & v_50687;
assign v_50690 = v_50091;
assign v_50692 = v_50689 & v_50691;
assign v_50694 = v_50587 & v_50693;
assign v_50696 = v_50087;
assign v_50698 = v_50695 & v_50697;
assign v_50700 = v_50584 & v_50699;
assign v_50702 = v_555;
assign v_50704 = v_50701 & v_50703;
assign v_50706 = v_50581 & v_50705;
assign v_50708 = v_551;
assign v_50710 = v_50707 & v_50709;
assign v_50712 = v_50578 & v_50711;
assign v_50714 = v_547;
assign v_50716 = v_50713 & v_50715;
assign v_50718 = v_50575 & v_50717;
assign v_50720 = v_543;
assign v_50722 = v_50719 & v_50721;
assign v_50723 = v_50722;
assign v_50725 = v_50135;
assign v_50726 = v_608;
assign v_50727 = v_50726;
assign v_50728 = v_50725 & v_50727;
assign v_50729 = v_50728;
assign v_50730 = v_50620 & v_50729;
assign v_50732 = v_50630 & v_50731;
assign v_50733 = v_50619 & v_50729;
assign v_50735 = v_50617 & v_50734;
assign v_50737 = v_50636 & v_50736;
assign v_50738 = v_50616 & v_50734;
assign v_50740 = v_50614 & v_50739;
assign v_50742 = v_50642 & v_50741;
assign v_50743 = v_50613 & v_50739;
assign v_50745 = v_50611 & v_50744;
assign v_50747 = v_50648 & v_50746;
assign v_50748 = v_50610 & v_50744;
assign v_50750 = v_50608 & v_50749;
assign v_50752 = v_50654 & v_50751;
assign v_50753 = v_50607 & v_50749;
assign v_50755 = v_50605 & v_50754;
assign v_50757 = v_50660 & v_50756;
assign v_50758 = v_50604 & v_50754;
assign v_50760 = v_50602 & v_50759;
assign v_50762 = v_50666 & v_50761;
assign v_50763 = v_50601 & v_50759;
assign v_50765 = v_50599 & v_50764;
assign v_50767 = v_50672 & v_50766;
assign v_50768 = v_50598 & v_50764;
assign v_50770 = v_50596 & v_50769;
assign v_50772 = v_50678 & v_50771;
assign v_50773 = v_50595 & v_50769;
assign v_50775 = v_50593 & v_50774;
assign v_50777 = v_50684 & v_50776;
assign v_50778 = v_50592 & v_50774;
assign v_50780 = v_50590 & v_50779;
assign v_50782 = v_50690 & v_50781;
assign v_50783 = v_50589 & v_50779;
assign v_50785 = v_50587 & v_50784;
assign v_50787 = v_50696 & v_50786;
assign v_50788 = v_50586 & v_50784;
assign v_50790 = v_50584 & v_50789;
assign v_50792 = v_50702 & v_50791;
assign v_50793 = v_50583 & v_50789;
assign v_50795 = v_50581 & v_50794;
assign v_50797 = v_50708 & v_50796;
assign v_50798 = v_50580 & v_50794;
assign v_50800 = v_50578 & v_50799;
assign v_50802 = v_50714 & v_50801;
assign v_50803 = v_50577 & v_50799;
assign v_50805 = v_50575 & v_50804;
assign v_50807 = v_50720 & v_50806;
assign v_50808 = v_50574 & v_50804;
assign v_50810 = v_50809;
assign v_50812 = v_50724 & v_50811;
assign v_50813 = v_50812;
assign v_50815 = v_50814;
assign v_50817 = ~v_803;
assign v_50818 = ~v_50072;
assign v_50819 = v_50072;
assign v_50820 = ~v_807;
assign v_50821 = ~v_50076;
assign v_50822 = v_50076;
assign v_50823 = ~v_811;
assign v_50824 = ~v_50080;
assign v_50825 = v_50080;
assign v_50826 = ~v_815;
assign v_50827 = ~v_50084;
assign v_50828 = v_50084;
assign v_50829 = ~v_50087;
assign v_50830 = ~v_820;
assign v_50831 = v_820;
assign v_50832 = ~v_50091;
assign v_50833 = ~v_824;
assign v_50834 = v_824;
assign v_50835 = ~v_50095;
assign v_50836 = ~v_828;
assign v_50837 = v_828;
assign v_50838 = ~v_50099;
assign v_50839 = ~v_832;
assign v_50840 = v_832;
assign v_50841 = ~v_50103;
assign v_50842 = ~v_836;
assign v_50843 = v_836;
assign v_50844 = ~v_50107;
assign v_50845 = ~v_840;
assign v_50846 = v_840;
assign v_50847 = ~v_50111;
assign v_50848 = ~v_844;
assign v_50849 = v_844;
assign v_50850 = ~v_50115;
assign v_50851 = ~v_848;
assign v_50852 = v_848;
assign v_50853 = ~v_50119;
assign v_50854 = ~v_852;
assign v_50855 = v_852;
assign v_50856 = ~v_50123;
assign v_50857 = ~v_856;
assign v_50858 = v_856;
assign v_50859 = ~v_50127;
assign v_50860 = ~v_860;
assign v_50861 = v_860;
assign v_50862 = ~v_50131;
assign v_50863 = ~v_864;
assign v_50864 = v_864;
assign v_50865 = ~v_50135;
assign v_50866 = ~v_868;
assign v_50867 = v_50866;
assign v_50869 = v_50868;
assign v_50871 = v_50863 & v_50870;
assign v_50873 = v_50131;
assign v_50875 = v_50872 & v_50874;
assign v_50877 = v_50860 & v_50876;
assign v_50879 = v_50127;
assign v_50881 = v_50878 & v_50880;
assign v_50883 = v_50857 & v_50882;
assign v_50885 = v_50123;
assign v_50887 = v_50884 & v_50886;
assign v_50889 = v_50854 & v_50888;
assign v_50891 = v_50119;
assign v_50893 = v_50890 & v_50892;
assign v_50895 = v_50851 & v_50894;
assign v_50897 = v_50115;
assign v_50899 = v_50896 & v_50898;
assign v_50901 = v_50848 & v_50900;
assign v_50903 = v_50111;
assign v_50905 = v_50902 & v_50904;
assign v_50907 = v_50845 & v_50906;
assign v_50909 = v_50107;
assign v_50911 = v_50908 & v_50910;
assign v_50913 = v_50842 & v_50912;
assign v_50915 = v_50103;
assign v_50917 = v_50914 & v_50916;
assign v_50919 = v_50839 & v_50918;
assign v_50921 = v_50099;
assign v_50923 = v_50920 & v_50922;
assign v_50925 = v_50836 & v_50924;
assign v_50927 = v_50095;
assign v_50929 = v_50926 & v_50928;
assign v_50931 = v_50833 & v_50930;
assign v_50933 = v_50091;
assign v_50935 = v_50932 & v_50934;
assign v_50937 = v_50830 & v_50936;
assign v_50939 = v_50087;
assign v_50941 = v_50938 & v_50940;
assign v_50943 = v_50827 & v_50942;
assign v_50945 = v_815;
assign v_50947 = v_50944 & v_50946;
assign v_50949 = v_50824 & v_50948;
assign v_50951 = v_811;
assign v_50953 = v_50950 & v_50952;
assign v_50955 = v_50821 & v_50954;
assign v_50957 = v_807;
assign v_50959 = v_50956 & v_50958;
assign v_50961 = v_50818 & v_50960;
assign v_50963 = v_803;
assign v_50965 = v_50962 & v_50964;
assign v_50966 = v_50965;
assign v_50968 = v_50135;
assign v_50969 = v_868;
assign v_50970 = v_50969;
assign v_50971 = v_50968 & v_50970;
assign v_50972 = v_50971;
assign v_50973 = v_50863 & v_50972;
assign v_50975 = v_50873 & v_50974;
assign v_50976 = v_50862 & v_50972;
assign v_50978 = v_50860 & v_50977;
assign v_50980 = v_50879 & v_50979;
assign v_50981 = v_50859 & v_50977;
assign v_50983 = v_50857 & v_50982;
assign v_50985 = v_50885 & v_50984;
assign v_50986 = v_50856 & v_50982;
assign v_50988 = v_50854 & v_50987;
assign v_50990 = v_50891 & v_50989;
assign v_50991 = v_50853 & v_50987;
assign v_50993 = v_50851 & v_50992;
assign v_50995 = v_50897 & v_50994;
assign v_50996 = v_50850 & v_50992;
assign v_50998 = v_50848 & v_50997;
assign v_51000 = v_50903 & v_50999;
assign v_51001 = v_50847 & v_50997;
assign v_51003 = v_50845 & v_51002;
assign v_51005 = v_50909 & v_51004;
assign v_51006 = v_50844 & v_51002;
assign v_51008 = v_50842 & v_51007;
assign v_51010 = v_50915 & v_51009;
assign v_51011 = v_50841 & v_51007;
assign v_51013 = v_50839 & v_51012;
assign v_51015 = v_50921 & v_51014;
assign v_51016 = v_50838 & v_51012;
assign v_51018 = v_50836 & v_51017;
assign v_51020 = v_50927 & v_51019;
assign v_51021 = v_50835 & v_51017;
assign v_51023 = v_50833 & v_51022;
assign v_51025 = v_50933 & v_51024;
assign v_51026 = v_50832 & v_51022;
assign v_51028 = v_50830 & v_51027;
assign v_51030 = v_50939 & v_51029;
assign v_51031 = v_50829 & v_51027;
assign v_51033 = v_50827 & v_51032;
assign v_51035 = v_50945 & v_51034;
assign v_51036 = v_50826 & v_51032;
assign v_51038 = v_50824 & v_51037;
assign v_51040 = v_50951 & v_51039;
assign v_51041 = v_50823 & v_51037;
assign v_51043 = v_50821 & v_51042;
assign v_51045 = v_50957 & v_51044;
assign v_51046 = v_50820 & v_51042;
assign v_51048 = v_50818 & v_51047;
assign v_51050 = v_50963 & v_51049;
assign v_51051 = v_50817 & v_51047;
assign v_51053 = v_51052;
assign v_51055 = v_50967 & v_51054;
assign v_51056 = v_51055;
assign v_51058 = v_51057;
assign v_51060 = ~v_1063;
assign v_51061 = ~v_50072;
assign v_51062 = v_50072;
assign v_51063 = ~v_1067;
assign v_51064 = ~v_50076;
assign v_51065 = v_50076;
assign v_51066 = ~v_1071;
assign v_51067 = ~v_50080;
assign v_51068 = v_50080;
assign v_51069 = ~v_1075;
assign v_51070 = ~v_50084;
assign v_51071 = v_50084;
assign v_51072 = ~v_50087;
assign v_51073 = ~v_1080;
assign v_51074 = v_1080;
assign v_51075 = ~v_50091;
assign v_51076 = ~v_1084;
assign v_51077 = v_1084;
assign v_51078 = ~v_50095;
assign v_51079 = ~v_1088;
assign v_51080 = v_1088;
assign v_51081 = ~v_50099;
assign v_51082 = ~v_1092;
assign v_51083 = v_1092;
assign v_51084 = ~v_50103;
assign v_51085 = ~v_1096;
assign v_51086 = v_1096;
assign v_51087 = ~v_50107;
assign v_51088 = ~v_1100;
assign v_51089 = v_1100;
assign v_51090 = ~v_50111;
assign v_51091 = ~v_1104;
assign v_51092 = v_1104;
assign v_51093 = ~v_50115;
assign v_51094 = ~v_1108;
assign v_51095 = v_1108;
assign v_51096 = ~v_50119;
assign v_51097 = ~v_1112;
assign v_51098 = v_1112;
assign v_51099 = ~v_50123;
assign v_51100 = ~v_1116;
assign v_51101 = v_1116;
assign v_51102 = ~v_50127;
assign v_51103 = ~v_1120;
assign v_51104 = v_1120;
assign v_51105 = ~v_50131;
assign v_51106 = ~v_1124;
assign v_51107 = v_1124;
assign v_51108 = ~v_50135;
assign v_51109 = ~v_1128;
assign v_51110 = v_51109;
assign v_51112 = v_51111;
assign v_51114 = v_51106 & v_51113;
assign v_51116 = v_50131;
assign v_51118 = v_51115 & v_51117;
assign v_51120 = v_51103 & v_51119;
assign v_51122 = v_50127;
assign v_51124 = v_51121 & v_51123;
assign v_51126 = v_51100 & v_51125;
assign v_51128 = v_50123;
assign v_51130 = v_51127 & v_51129;
assign v_51132 = v_51097 & v_51131;
assign v_51134 = v_50119;
assign v_51136 = v_51133 & v_51135;
assign v_51138 = v_51094 & v_51137;
assign v_51140 = v_50115;
assign v_51142 = v_51139 & v_51141;
assign v_51144 = v_51091 & v_51143;
assign v_51146 = v_50111;
assign v_51148 = v_51145 & v_51147;
assign v_51150 = v_51088 & v_51149;
assign v_51152 = v_50107;
assign v_51154 = v_51151 & v_51153;
assign v_51156 = v_51085 & v_51155;
assign v_51158 = v_50103;
assign v_51160 = v_51157 & v_51159;
assign v_51162 = v_51082 & v_51161;
assign v_51164 = v_50099;
assign v_51166 = v_51163 & v_51165;
assign v_51168 = v_51079 & v_51167;
assign v_51170 = v_50095;
assign v_51172 = v_51169 & v_51171;
assign v_51174 = v_51076 & v_51173;
assign v_51176 = v_50091;
assign v_51178 = v_51175 & v_51177;
assign v_51180 = v_51073 & v_51179;
assign v_51182 = v_50087;
assign v_51184 = v_51181 & v_51183;
assign v_51186 = v_51070 & v_51185;
assign v_51188 = v_1075;
assign v_51190 = v_51187 & v_51189;
assign v_51192 = v_51067 & v_51191;
assign v_51194 = v_1071;
assign v_51196 = v_51193 & v_51195;
assign v_51198 = v_51064 & v_51197;
assign v_51200 = v_1067;
assign v_51202 = v_51199 & v_51201;
assign v_51204 = v_51061 & v_51203;
assign v_51206 = v_1063;
assign v_51208 = v_51205 & v_51207;
assign v_51209 = v_51208;
assign v_51211 = v_50135;
assign v_51212 = v_1128;
assign v_51213 = v_51212;
assign v_51214 = v_51211 & v_51213;
assign v_51215 = v_51214;
assign v_51216 = v_51106 & v_51215;
assign v_51218 = v_51116 & v_51217;
assign v_51219 = v_51105 & v_51215;
assign v_51221 = v_51103 & v_51220;
assign v_51223 = v_51122 & v_51222;
assign v_51224 = v_51102 & v_51220;
assign v_51226 = v_51100 & v_51225;
assign v_51228 = v_51128 & v_51227;
assign v_51229 = v_51099 & v_51225;
assign v_51231 = v_51097 & v_51230;
assign v_51233 = v_51134 & v_51232;
assign v_51234 = v_51096 & v_51230;
assign v_51236 = v_51094 & v_51235;
assign v_51238 = v_51140 & v_51237;
assign v_51239 = v_51093 & v_51235;
assign v_51241 = v_51091 & v_51240;
assign v_51243 = v_51146 & v_51242;
assign v_51244 = v_51090 & v_51240;
assign v_51246 = v_51088 & v_51245;
assign v_51248 = v_51152 & v_51247;
assign v_51249 = v_51087 & v_51245;
assign v_51251 = v_51085 & v_51250;
assign v_51253 = v_51158 & v_51252;
assign v_51254 = v_51084 & v_51250;
assign v_51256 = v_51082 & v_51255;
assign v_51258 = v_51164 & v_51257;
assign v_51259 = v_51081 & v_51255;
assign v_51261 = v_51079 & v_51260;
assign v_51263 = v_51170 & v_51262;
assign v_51264 = v_51078 & v_51260;
assign v_51266 = v_51076 & v_51265;
assign v_51268 = v_51176 & v_51267;
assign v_51269 = v_51075 & v_51265;
assign v_51271 = v_51073 & v_51270;
assign v_51273 = v_51182 & v_51272;
assign v_51274 = v_51072 & v_51270;
assign v_51276 = v_51070 & v_51275;
assign v_51278 = v_51188 & v_51277;
assign v_51279 = v_51069 & v_51275;
assign v_51281 = v_51067 & v_51280;
assign v_51283 = v_51194 & v_51282;
assign v_51284 = v_51066 & v_51280;
assign v_51286 = v_51064 & v_51285;
assign v_51288 = v_51200 & v_51287;
assign v_51289 = v_51063 & v_51285;
assign v_51291 = v_51061 & v_51290;
assign v_51293 = v_51206 & v_51292;
assign v_51294 = v_51060 & v_51290;
assign v_51296 = v_51295;
assign v_51298 = v_51210 & v_51297;
assign v_51299 = v_51298;
assign v_51301 = v_51300;
assign v_51303 = ~v_1323;
assign v_51304 = ~v_50072;
assign v_51305 = v_50072;
assign v_51306 = ~v_1327;
assign v_51307 = ~v_50076;
assign v_51308 = v_50076;
assign v_51309 = ~v_1331;
assign v_51310 = ~v_50080;
assign v_51311 = v_50080;
assign v_51312 = ~v_1335;
assign v_51313 = ~v_50084;
assign v_51314 = v_50084;
assign v_51315 = ~v_50087;
assign v_51316 = ~v_1340;
assign v_51317 = v_1340;
assign v_51318 = ~v_50091;
assign v_51319 = ~v_1344;
assign v_51320 = v_1344;
assign v_51321 = ~v_50095;
assign v_51322 = ~v_1348;
assign v_51323 = v_1348;
assign v_51324 = ~v_50099;
assign v_51325 = ~v_1352;
assign v_51326 = v_1352;
assign v_51327 = ~v_50103;
assign v_51328 = ~v_1356;
assign v_51329 = v_1356;
assign v_51330 = ~v_50107;
assign v_51331 = ~v_1360;
assign v_51332 = v_1360;
assign v_51333 = ~v_50111;
assign v_51334 = ~v_1364;
assign v_51335 = v_1364;
assign v_51336 = ~v_50115;
assign v_51337 = ~v_1368;
assign v_51338 = v_1368;
assign v_51339 = ~v_50119;
assign v_51340 = ~v_1372;
assign v_51341 = v_1372;
assign v_51342 = ~v_50123;
assign v_51343 = ~v_1376;
assign v_51344 = v_1376;
assign v_51345 = ~v_50127;
assign v_51346 = ~v_1380;
assign v_51347 = v_1380;
assign v_51348 = ~v_50131;
assign v_51349 = ~v_1384;
assign v_51350 = v_1384;
assign v_51351 = ~v_50135;
assign v_51352 = ~v_1388;
assign v_51353 = v_51352;
assign v_51355 = v_51354;
assign v_51357 = v_51349 & v_51356;
assign v_51359 = v_50131;
assign v_51361 = v_51358 & v_51360;
assign v_51363 = v_51346 & v_51362;
assign v_51365 = v_50127;
assign v_51367 = v_51364 & v_51366;
assign v_51369 = v_51343 & v_51368;
assign v_51371 = v_50123;
assign v_51373 = v_51370 & v_51372;
assign v_51375 = v_51340 & v_51374;
assign v_51377 = v_50119;
assign v_51379 = v_51376 & v_51378;
assign v_51381 = v_51337 & v_51380;
assign v_51383 = v_50115;
assign v_51385 = v_51382 & v_51384;
assign v_51387 = v_51334 & v_51386;
assign v_51389 = v_50111;
assign v_51391 = v_51388 & v_51390;
assign v_51393 = v_51331 & v_51392;
assign v_51395 = v_50107;
assign v_51397 = v_51394 & v_51396;
assign v_51399 = v_51328 & v_51398;
assign v_51401 = v_50103;
assign v_51403 = v_51400 & v_51402;
assign v_51405 = v_51325 & v_51404;
assign v_51407 = v_50099;
assign v_51409 = v_51406 & v_51408;
assign v_51411 = v_51322 & v_51410;
assign v_51413 = v_50095;
assign v_51415 = v_51412 & v_51414;
assign v_51417 = v_51319 & v_51416;
assign v_51419 = v_50091;
assign v_51421 = v_51418 & v_51420;
assign v_51423 = v_51316 & v_51422;
assign v_51425 = v_50087;
assign v_51427 = v_51424 & v_51426;
assign v_51429 = v_51313 & v_51428;
assign v_51431 = v_1335;
assign v_51433 = v_51430 & v_51432;
assign v_51435 = v_51310 & v_51434;
assign v_51437 = v_1331;
assign v_51439 = v_51436 & v_51438;
assign v_51441 = v_51307 & v_51440;
assign v_51443 = v_1327;
assign v_51445 = v_51442 & v_51444;
assign v_51447 = v_51304 & v_51446;
assign v_51449 = v_1323;
assign v_51451 = v_51448 & v_51450;
assign v_51452 = v_51451;
assign v_51454 = v_50135;
assign v_51455 = v_1388;
assign v_51456 = v_51455;
assign v_51457 = v_51454 & v_51456;
assign v_51458 = v_51457;
assign v_51459 = v_51349 & v_51458;
assign v_51461 = v_51359 & v_51460;
assign v_51462 = v_51348 & v_51458;
assign v_51464 = v_51346 & v_51463;
assign v_51466 = v_51365 & v_51465;
assign v_51467 = v_51345 & v_51463;
assign v_51469 = v_51343 & v_51468;
assign v_51471 = v_51371 & v_51470;
assign v_51472 = v_51342 & v_51468;
assign v_51474 = v_51340 & v_51473;
assign v_51476 = v_51377 & v_51475;
assign v_51477 = v_51339 & v_51473;
assign v_51479 = v_51337 & v_51478;
assign v_51481 = v_51383 & v_51480;
assign v_51482 = v_51336 & v_51478;
assign v_51484 = v_51334 & v_51483;
assign v_51486 = v_51389 & v_51485;
assign v_51487 = v_51333 & v_51483;
assign v_51489 = v_51331 & v_51488;
assign v_51491 = v_51395 & v_51490;
assign v_51492 = v_51330 & v_51488;
assign v_51494 = v_51328 & v_51493;
assign v_51496 = v_51401 & v_51495;
assign v_51497 = v_51327 & v_51493;
assign v_51499 = v_51325 & v_51498;
assign v_51501 = v_51407 & v_51500;
assign v_51502 = v_51324 & v_51498;
assign v_51504 = v_51322 & v_51503;
assign v_51506 = v_51413 & v_51505;
assign v_51507 = v_51321 & v_51503;
assign v_51509 = v_51319 & v_51508;
assign v_51511 = v_51419 & v_51510;
assign v_51512 = v_51318 & v_51508;
assign v_51514 = v_51316 & v_51513;
assign v_51516 = v_51425 & v_51515;
assign v_51517 = v_51315 & v_51513;
assign v_51519 = v_51313 & v_51518;
assign v_51521 = v_51431 & v_51520;
assign v_51522 = v_51312 & v_51518;
assign v_51524 = v_51310 & v_51523;
assign v_51526 = v_51437 & v_51525;
assign v_51527 = v_51309 & v_51523;
assign v_51529 = v_51307 & v_51528;
assign v_51531 = v_51443 & v_51530;
assign v_51532 = v_51306 & v_51528;
assign v_51534 = v_51304 & v_51533;
assign v_51536 = v_51449 & v_51535;
assign v_51537 = v_51303 & v_51533;
assign v_51539 = v_51538;
assign v_51541 = v_51453 & v_51540;
assign v_51542 = v_51541;
assign v_51544 = v_51543;
assign v_51546 = ~v_1583;
assign v_51547 = ~v_50072;
assign v_51548 = v_50072;
assign v_51549 = ~v_1587;
assign v_51550 = ~v_50076;
assign v_51551 = v_50076;
assign v_51552 = ~v_1591;
assign v_51553 = ~v_50080;
assign v_51554 = v_50080;
assign v_51555 = ~v_1595;
assign v_51556 = ~v_50084;
assign v_51557 = v_50084;
assign v_51558 = ~v_50087;
assign v_51559 = ~v_1600;
assign v_51560 = v_1600;
assign v_51561 = ~v_50091;
assign v_51562 = ~v_1604;
assign v_51563 = v_1604;
assign v_51564 = ~v_50095;
assign v_51565 = ~v_1608;
assign v_51566 = v_1608;
assign v_51567 = ~v_50099;
assign v_51568 = ~v_1612;
assign v_51569 = v_1612;
assign v_51570 = ~v_50103;
assign v_51571 = ~v_1616;
assign v_51572 = v_1616;
assign v_51573 = ~v_50107;
assign v_51574 = ~v_1620;
assign v_51575 = v_1620;
assign v_51576 = ~v_50111;
assign v_51577 = ~v_1624;
assign v_51578 = v_1624;
assign v_51579 = ~v_50115;
assign v_51580 = ~v_1628;
assign v_51581 = v_1628;
assign v_51582 = ~v_50119;
assign v_51583 = ~v_1632;
assign v_51584 = v_1632;
assign v_51585 = ~v_50123;
assign v_51586 = ~v_1636;
assign v_51587 = v_1636;
assign v_51588 = ~v_50127;
assign v_51589 = ~v_1640;
assign v_51590 = v_1640;
assign v_51591 = ~v_50131;
assign v_51592 = ~v_1644;
assign v_51593 = v_1644;
assign v_51594 = ~v_50135;
assign v_51595 = ~v_1648;
assign v_51596 = v_51595;
assign v_51598 = v_51597;
assign v_51600 = v_51592 & v_51599;
assign v_51602 = v_50131;
assign v_51604 = v_51601 & v_51603;
assign v_51606 = v_51589 & v_51605;
assign v_51608 = v_50127;
assign v_51610 = v_51607 & v_51609;
assign v_51612 = v_51586 & v_51611;
assign v_51614 = v_50123;
assign v_51616 = v_51613 & v_51615;
assign v_51618 = v_51583 & v_51617;
assign v_51620 = v_50119;
assign v_51622 = v_51619 & v_51621;
assign v_51624 = v_51580 & v_51623;
assign v_51626 = v_50115;
assign v_51628 = v_51625 & v_51627;
assign v_51630 = v_51577 & v_51629;
assign v_51632 = v_50111;
assign v_51634 = v_51631 & v_51633;
assign v_51636 = v_51574 & v_51635;
assign v_51638 = v_50107;
assign v_51640 = v_51637 & v_51639;
assign v_51642 = v_51571 & v_51641;
assign v_51644 = v_50103;
assign v_51646 = v_51643 & v_51645;
assign v_51648 = v_51568 & v_51647;
assign v_51650 = v_50099;
assign v_51652 = v_51649 & v_51651;
assign v_51654 = v_51565 & v_51653;
assign v_51656 = v_50095;
assign v_51658 = v_51655 & v_51657;
assign v_51660 = v_51562 & v_51659;
assign v_51662 = v_50091;
assign v_51664 = v_51661 & v_51663;
assign v_51666 = v_51559 & v_51665;
assign v_51668 = v_50087;
assign v_51670 = v_51667 & v_51669;
assign v_51672 = v_51556 & v_51671;
assign v_51674 = v_1595;
assign v_51676 = v_51673 & v_51675;
assign v_51678 = v_51553 & v_51677;
assign v_51680 = v_1591;
assign v_51682 = v_51679 & v_51681;
assign v_51684 = v_51550 & v_51683;
assign v_51686 = v_1587;
assign v_51688 = v_51685 & v_51687;
assign v_51690 = v_51547 & v_51689;
assign v_51692 = v_1583;
assign v_51694 = v_51691 & v_51693;
assign v_51695 = v_51694;
assign v_51697 = v_50135;
assign v_51698 = v_1648;
assign v_51699 = v_51698;
assign v_51700 = v_51697 & v_51699;
assign v_51701 = v_51700;
assign v_51702 = v_51592 & v_51701;
assign v_51704 = v_51602 & v_51703;
assign v_51705 = v_51591 & v_51701;
assign v_51707 = v_51589 & v_51706;
assign v_51709 = v_51608 & v_51708;
assign v_51710 = v_51588 & v_51706;
assign v_51712 = v_51586 & v_51711;
assign v_51714 = v_51614 & v_51713;
assign v_51715 = v_51585 & v_51711;
assign v_51717 = v_51583 & v_51716;
assign v_51719 = v_51620 & v_51718;
assign v_51720 = v_51582 & v_51716;
assign v_51722 = v_51580 & v_51721;
assign v_51724 = v_51626 & v_51723;
assign v_51725 = v_51579 & v_51721;
assign v_51727 = v_51577 & v_51726;
assign v_51729 = v_51632 & v_51728;
assign v_51730 = v_51576 & v_51726;
assign v_51732 = v_51574 & v_51731;
assign v_51734 = v_51638 & v_51733;
assign v_51735 = v_51573 & v_51731;
assign v_51737 = v_51571 & v_51736;
assign v_51739 = v_51644 & v_51738;
assign v_51740 = v_51570 & v_51736;
assign v_51742 = v_51568 & v_51741;
assign v_51744 = v_51650 & v_51743;
assign v_51745 = v_51567 & v_51741;
assign v_51747 = v_51565 & v_51746;
assign v_51749 = v_51656 & v_51748;
assign v_51750 = v_51564 & v_51746;
assign v_51752 = v_51562 & v_51751;
assign v_51754 = v_51662 & v_51753;
assign v_51755 = v_51561 & v_51751;
assign v_51757 = v_51559 & v_51756;
assign v_51759 = v_51668 & v_51758;
assign v_51760 = v_51558 & v_51756;
assign v_51762 = v_51556 & v_51761;
assign v_51764 = v_51674 & v_51763;
assign v_51765 = v_51555 & v_51761;
assign v_51767 = v_51553 & v_51766;
assign v_51769 = v_51680 & v_51768;
assign v_51770 = v_51552 & v_51766;
assign v_51772 = v_51550 & v_51771;
assign v_51774 = v_51686 & v_51773;
assign v_51775 = v_51549 & v_51771;
assign v_51777 = v_51547 & v_51776;
assign v_51779 = v_51692 & v_51778;
assign v_51780 = v_51546 & v_51776;
assign v_51782 = v_51781;
assign v_51784 = v_51696 & v_51783;
assign v_51785 = v_51784;
assign v_51787 = v_51786;
assign v_51789 = ~v_1843;
assign v_51790 = ~v_50072;
assign v_51791 = v_50072;
assign v_51792 = ~v_1847;
assign v_51793 = ~v_50076;
assign v_51794 = v_50076;
assign v_51795 = ~v_1851;
assign v_51796 = ~v_50080;
assign v_51797 = v_50080;
assign v_51798 = ~v_1855;
assign v_51799 = ~v_50084;
assign v_51800 = v_50084;
assign v_51801 = ~v_50087;
assign v_51802 = ~v_1860;
assign v_51803 = v_1860;
assign v_51804 = ~v_50091;
assign v_51805 = ~v_1864;
assign v_51806 = v_1864;
assign v_51807 = ~v_50095;
assign v_51808 = ~v_1868;
assign v_51809 = v_1868;
assign v_51810 = ~v_50099;
assign v_51811 = ~v_1872;
assign v_51812 = v_1872;
assign v_51813 = ~v_50103;
assign v_51814 = ~v_1876;
assign v_51815 = v_1876;
assign v_51816 = ~v_50107;
assign v_51817 = ~v_1880;
assign v_51818 = v_1880;
assign v_51819 = ~v_50111;
assign v_51820 = ~v_1884;
assign v_51821 = v_1884;
assign v_51822 = ~v_50115;
assign v_51823 = ~v_1888;
assign v_51824 = v_1888;
assign v_51825 = ~v_50119;
assign v_51826 = ~v_1892;
assign v_51827 = v_1892;
assign v_51828 = ~v_50123;
assign v_51829 = ~v_1896;
assign v_51830 = v_1896;
assign v_51831 = ~v_50127;
assign v_51832 = ~v_1900;
assign v_51833 = v_1900;
assign v_51834 = ~v_50131;
assign v_51835 = ~v_1904;
assign v_51836 = v_1904;
assign v_51837 = ~v_50135;
assign v_51838 = ~v_1908;
assign v_51839 = v_51838;
assign v_51841 = v_51840;
assign v_51843 = v_51835 & v_51842;
assign v_51845 = v_50131;
assign v_51847 = v_51844 & v_51846;
assign v_51849 = v_51832 & v_51848;
assign v_51851 = v_50127;
assign v_51853 = v_51850 & v_51852;
assign v_51855 = v_51829 & v_51854;
assign v_51857 = v_50123;
assign v_51859 = v_51856 & v_51858;
assign v_51861 = v_51826 & v_51860;
assign v_51863 = v_50119;
assign v_51865 = v_51862 & v_51864;
assign v_51867 = v_51823 & v_51866;
assign v_51869 = v_50115;
assign v_51871 = v_51868 & v_51870;
assign v_51873 = v_51820 & v_51872;
assign v_51875 = v_50111;
assign v_51877 = v_51874 & v_51876;
assign v_51879 = v_51817 & v_51878;
assign v_51881 = v_50107;
assign v_51883 = v_51880 & v_51882;
assign v_51885 = v_51814 & v_51884;
assign v_51887 = v_50103;
assign v_51889 = v_51886 & v_51888;
assign v_51891 = v_51811 & v_51890;
assign v_51893 = v_50099;
assign v_51895 = v_51892 & v_51894;
assign v_51897 = v_51808 & v_51896;
assign v_51899 = v_50095;
assign v_51901 = v_51898 & v_51900;
assign v_51903 = v_51805 & v_51902;
assign v_51905 = v_50091;
assign v_51907 = v_51904 & v_51906;
assign v_51909 = v_51802 & v_51908;
assign v_51911 = v_50087;
assign v_51913 = v_51910 & v_51912;
assign v_51915 = v_51799 & v_51914;
assign v_51917 = v_1855;
assign v_51919 = v_51916 & v_51918;
assign v_51921 = v_51796 & v_51920;
assign v_51923 = v_1851;
assign v_51925 = v_51922 & v_51924;
assign v_51927 = v_51793 & v_51926;
assign v_51929 = v_1847;
assign v_51931 = v_51928 & v_51930;
assign v_51933 = v_51790 & v_51932;
assign v_51935 = v_1843;
assign v_51937 = v_51934 & v_51936;
assign v_51938 = v_51937;
assign v_51940 = v_50135;
assign v_51941 = v_1908;
assign v_51942 = v_51941;
assign v_51943 = v_51940 & v_51942;
assign v_51944 = v_51943;
assign v_51945 = v_51835 & v_51944;
assign v_51947 = v_51845 & v_51946;
assign v_51948 = v_51834 & v_51944;
assign v_51950 = v_51832 & v_51949;
assign v_51952 = v_51851 & v_51951;
assign v_51953 = v_51831 & v_51949;
assign v_51955 = v_51829 & v_51954;
assign v_51957 = v_51857 & v_51956;
assign v_51958 = v_51828 & v_51954;
assign v_51960 = v_51826 & v_51959;
assign v_51962 = v_51863 & v_51961;
assign v_51963 = v_51825 & v_51959;
assign v_51965 = v_51823 & v_51964;
assign v_51967 = v_51869 & v_51966;
assign v_51968 = v_51822 & v_51964;
assign v_51970 = v_51820 & v_51969;
assign v_51972 = v_51875 & v_51971;
assign v_51973 = v_51819 & v_51969;
assign v_51975 = v_51817 & v_51974;
assign v_51977 = v_51881 & v_51976;
assign v_51978 = v_51816 & v_51974;
assign v_51980 = v_51814 & v_51979;
assign v_51982 = v_51887 & v_51981;
assign v_51983 = v_51813 & v_51979;
assign v_51985 = v_51811 & v_51984;
assign v_51987 = v_51893 & v_51986;
assign v_51988 = v_51810 & v_51984;
assign v_51990 = v_51808 & v_51989;
assign v_51992 = v_51899 & v_51991;
assign v_51993 = v_51807 & v_51989;
assign v_51995 = v_51805 & v_51994;
assign v_51997 = v_51905 & v_51996;
assign v_51998 = v_51804 & v_51994;
assign v_52000 = v_51802 & v_51999;
assign v_52002 = v_51911 & v_52001;
assign v_52003 = v_51801 & v_51999;
assign v_52005 = v_51799 & v_52004;
assign v_52007 = v_51917 & v_52006;
assign v_52008 = v_51798 & v_52004;
assign v_52010 = v_51796 & v_52009;
assign v_52012 = v_51923 & v_52011;
assign v_52013 = v_51795 & v_52009;
assign v_52015 = v_51793 & v_52014;
assign v_52017 = v_51929 & v_52016;
assign v_52018 = v_51792 & v_52014;
assign v_52020 = v_51790 & v_52019;
assign v_52022 = v_51935 & v_52021;
assign v_52023 = v_51789 & v_52019;
assign v_52025 = v_52024;
assign v_52027 = v_51939 & v_52026;
assign v_52028 = v_52027;
assign v_52030 = v_52029;
assign v_52032 = ~v_2103;
assign v_52033 = ~v_50072;
assign v_52034 = v_50072;
assign v_52035 = ~v_2107;
assign v_52036 = ~v_50076;
assign v_52037 = v_50076;
assign v_52038 = ~v_2111;
assign v_52039 = ~v_50080;
assign v_52040 = v_50080;
assign v_52041 = ~v_2115;
assign v_52042 = ~v_50084;
assign v_52043 = v_50084;
assign v_52044 = ~v_50087;
assign v_52045 = ~v_2120;
assign v_52046 = v_2120;
assign v_52047 = ~v_50091;
assign v_52048 = ~v_2124;
assign v_52049 = v_2124;
assign v_52050 = ~v_50095;
assign v_52051 = ~v_2128;
assign v_52052 = v_2128;
assign v_52053 = ~v_50099;
assign v_52054 = ~v_2132;
assign v_52055 = v_2132;
assign v_52056 = ~v_50103;
assign v_52057 = ~v_2136;
assign v_52058 = v_2136;
assign v_52059 = ~v_50107;
assign v_52060 = ~v_2140;
assign v_52061 = v_2140;
assign v_52062 = ~v_50111;
assign v_52063 = ~v_2144;
assign v_52064 = v_2144;
assign v_52065 = ~v_50115;
assign v_52066 = ~v_2148;
assign v_52067 = v_2148;
assign v_52068 = ~v_50119;
assign v_52069 = ~v_2152;
assign v_52070 = v_2152;
assign v_52071 = ~v_50123;
assign v_52072 = ~v_2156;
assign v_52073 = v_2156;
assign v_52074 = ~v_50127;
assign v_52075 = ~v_2160;
assign v_52076 = v_2160;
assign v_52077 = ~v_50131;
assign v_52078 = ~v_2164;
assign v_52079 = v_2164;
assign v_52080 = ~v_50135;
assign v_52081 = ~v_2168;
assign v_52082 = v_52081;
assign v_52084 = v_52083;
assign v_52086 = v_52078 & v_52085;
assign v_52088 = v_50131;
assign v_52090 = v_52087 & v_52089;
assign v_52092 = v_52075 & v_52091;
assign v_52094 = v_50127;
assign v_52096 = v_52093 & v_52095;
assign v_52098 = v_52072 & v_52097;
assign v_52100 = v_50123;
assign v_52102 = v_52099 & v_52101;
assign v_52104 = v_52069 & v_52103;
assign v_52106 = v_50119;
assign v_52108 = v_52105 & v_52107;
assign v_52110 = v_52066 & v_52109;
assign v_52112 = v_50115;
assign v_52114 = v_52111 & v_52113;
assign v_52116 = v_52063 & v_52115;
assign v_52118 = v_50111;
assign v_52120 = v_52117 & v_52119;
assign v_52122 = v_52060 & v_52121;
assign v_52124 = v_50107;
assign v_52126 = v_52123 & v_52125;
assign v_52128 = v_52057 & v_52127;
assign v_52130 = v_50103;
assign v_52132 = v_52129 & v_52131;
assign v_52134 = v_52054 & v_52133;
assign v_52136 = v_50099;
assign v_52138 = v_52135 & v_52137;
assign v_52140 = v_52051 & v_52139;
assign v_52142 = v_50095;
assign v_52144 = v_52141 & v_52143;
assign v_52146 = v_52048 & v_52145;
assign v_52148 = v_50091;
assign v_52150 = v_52147 & v_52149;
assign v_52152 = v_52045 & v_52151;
assign v_52154 = v_50087;
assign v_52156 = v_52153 & v_52155;
assign v_52158 = v_52042 & v_52157;
assign v_52160 = v_2115;
assign v_52162 = v_52159 & v_52161;
assign v_52164 = v_52039 & v_52163;
assign v_52166 = v_2111;
assign v_52168 = v_52165 & v_52167;
assign v_52170 = v_52036 & v_52169;
assign v_52172 = v_2107;
assign v_52174 = v_52171 & v_52173;
assign v_52176 = v_52033 & v_52175;
assign v_52178 = v_2103;
assign v_52180 = v_52177 & v_52179;
assign v_52181 = v_52180;
assign v_52183 = v_50135;
assign v_52184 = v_2168;
assign v_52185 = v_52184;
assign v_52186 = v_52183 & v_52185;
assign v_52187 = v_52186;
assign v_52188 = v_52078 & v_52187;
assign v_52190 = v_52088 & v_52189;
assign v_52191 = v_52077 & v_52187;
assign v_52193 = v_52075 & v_52192;
assign v_52195 = v_52094 & v_52194;
assign v_52196 = v_52074 & v_52192;
assign v_52198 = v_52072 & v_52197;
assign v_52200 = v_52100 & v_52199;
assign v_52201 = v_52071 & v_52197;
assign v_52203 = v_52069 & v_52202;
assign v_52205 = v_52106 & v_52204;
assign v_52206 = v_52068 & v_52202;
assign v_52208 = v_52066 & v_52207;
assign v_52210 = v_52112 & v_52209;
assign v_52211 = v_52065 & v_52207;
assign v_52213 = v_52063 & v_52212;
assign v_52215 = v_52118 & v_52214;
assign v_52216 = v_52062 & v_52212;
assign v_52218 = v_52060 & v_52217;
assign v_52220 = v_52124 & v_52219;
assign v_52221 = v_52059 & v_52217;
assign v_52223 = v_52057 & v_52222;
assign v_52225 = v_52130 & v_52224;
assign v_52226 = v_52056 & v_52222;
assign v_52228 = v_52054 & v_52227;
assign v_52230 = v_52136 & v_52229;
assign v_52231 = v_52053 & v_52227;
assign v_52233 = v_52051 & v_52232;
assign v_52235 = v_52142 & v_52234;
assign v_52236 = v_52050 & v_52232;
assign v_52238 = v_52048 & v_52237;
assign v_52240 = v_52148 & v_52239;
assign v_52241 = v_52047 & v_52237;
assign v_52243 = v_52045 & v_52242;
assign v_52245 = v_52154 & v_52244;
assign v_52246 = v_52044 & v_52242;
assign v_52248 = v_52042 & v_52247;
assign v_52250 = v_52160 & v_52249;
assign v_52251 = v_52041 & v_52247;
assign v_52253 = v_52039 & v_52252;
assign v_52255 = v_52166 & v_52254;
assign v_52256 = v_52038 & v_52252;
assign v_52258 = v_52036 & v_52257;
assign v_52260 = v_52172 & v_52259;
assign v_52261 = v_52035 & v_52257;
assign v_52263 = v_52033 & v_52262;
assign v_52265 = v_52178 & v_52264;
assign v_52266 = v_52032 & v_52262;
assign v_52268 = v_52267;
assign v_52270 = v_52182 & v_52269;
assign v_52271 = v_52270;
assign v_52273 = v_52272;
assign v_52275 = ~v_2363;
assign v_52276 = ~v_50072;
assign v_52277 = v_50072;
assign v_52278 = ~v_2367;
assign v_52279 = ~v_50076;
assign v_52280 = v_50076;
assign v_52281 = ~v_2371;
assign v_52282 = ~v_50080;
assign v_52283 = v_50080;
assign v_52284 = ~v_2375;
assign v_52285 = ~v_50084;
assign v_52286 = v_50084;
assign v_52287 = ~v_50087;
assign v_52288 = ~v_2380;
assign v_52289 = v_2380;
assign v_52290 = ~v_50091;
assign v_52291 = ~v_2384;
assign v_52292 = v_2384;
assign v_52293 = ~v_50095;
assign v_52294 = ~v_2388;
assign v_52295 = v_2388;
assign v_52296 = ~v_50099;
assign v_52297 = ~v_2392;
assign v_52298 = v_2392;
assign v_52299 = ~v_50103;
assign v_52300 = ~v_2396;
assign v_52301 = v_2396;
assign v_52302 = ~v_50107;
assign v_52303 = ~v_2400;
assign v_52304 = v_2400;
assign v_52305 = ~v_50111;
assign v_52306 = ~v_2404;
assign v_52307 = v_2404;
assign v_52308 = ~v_50115;
assign v_52309 = ~v_2408;
assign v_52310 = v_2408;
assign v_52311 = ~v_50119;
assign v_52312 = ~v_2412;
assign v_52313 = v_2412;
assign v_52314 = ~v_50123;
assign v_52315 = ~v_2416;
assign v_52316 = v_2416;
assign v_52317 = ~v_50127;
assign v_52318 = ~v_2420;
assign v_52319 = v_2420;
assign v_52320 = ~v_50131;
assign v_52321 = ~v_2424;
assign v_52322 = v_2424;
assign v_52323 = ~v_50135;
assign v_52324 = ~v_2428;
assign v_52325 = v_52324;
assign v_52327 = v_52326;
assign v_52329 = v_52321 & v_52328;
assign v_52331 = v_50131;
assign v_52333 = v_52330 & v_52332;
assign v_52335 = v_52318 & v_52334;
assign v_52337 = v_50127;
assign v_52339 = v_52336 & v_52338;
assign v_52341 = v_52315 & v_52340;
assign v_52343 = v_50123;
assign v_52345 = v_52342 & v_52344;
assign v_52347 = v_52312 & v_52346;
assign v_52349 = v_50119;
assign v_52351 = v_52348 & v_52350;
assign v_52353 = v_52309 & v_52352;
assign v_52355 = v_50115;
assign v_52357 = v_52354 & v_52356;
assign v_52359 = v_52306 & v_52358;
assign v_52361 = v_50111;
assign v_52363 = v_52360 & v_52362;
assign v_52365 = v_52303 & v_52364;
assign v_52367 = v_50107;
assign v_52369 = v_52366 & v_52368;
assign v_52371 = v_52300 & v_52370;
assign v_52373 = v_50103;
assign v_52375 = v_52372 & v_52374;
assign v_52377 = v_52297 & v_52376;
assign v_52379 = v_50099;
assign v_52381 = v_52378 & v_52380;
assign v_52383 = v_52294 & v_52382;
assign v_52385 = v_50095;
assign v_52387 = v_52384 & v_52386;
assign v_52389 = v_52291 & v_52388;
assign v_52391 = v_50091;
assign v_52393 = v_52390 & v_52392;
assign v_52395 = v_52288 & v_52394;
assign v_52397 = v_50087;
assign v_52399 = v_52396 & v_52398;
assign v_52401 = v_52285 & v_52400;
assign v_52403 = v_2375;
assign v_52405 = v_52402 & v_52404;
assign v_52407 = v_52282 & v_52406;
assign v_52409 = v_2371;
assign v_52411 = v_52408 & v_52410;
assign v_52413 = v_52279 & v_52412;
assign v_52415 = v_2367;
assign v_52417 = v_52414 & v_52416;
assign v_52419 = v_52276 & v_52418;
assign v_52421 = v_2363;
assign v_52423 = v_52420 & v_52422;
assign v_52424 = v_52423;
assign v_52426 = v_50135;
assign v_52427 = v_2428;
assign v_52428 = v_52427;
assign v_52429 = v_52426 & v_52428;
assign v_52430 = v_52429;
assign v_52431 = v_52321 & v_52430;
assign v_52433 = v_52331 & v_52432;
assign v_52434 = v_52320 & v_52430;
assign v_52436 = v_52318 & v_52435;
assign v_52438 = v_52337 & v_52437;
assign v_52439 = v_52317 & v_52435;
assign v_52441 = v_52315 & v_52440;
assign v_52443 = v_52343 & v_52442;
assign v_52444 = v_52314 & v_52440;
assign v_52446 = v_52312 & v_52445;
assign v_52448 = v_52349 & v_52447;
assign v_52449 = v_52311 & v_52445;
assign v_52451 = v_52309 & v_52450;
assign v_52453 = v_52355 & v_52452;
assign v_52454 = v_52308 & v_52450;
assign v_52456 = v_52306 & v_52455;
assign v_52458 = v_52361 & v_52457;
assign v_52459 = v_52305 & v_52455;
assign v_52461 = v_52303 & v_52460;
assign v_52463 = v_52367 & v_52462;
assign v_52464 = v_52302 & v_52460;
assign v_52466 = v_52300 & v_52465;
assign v_52468 = v_52373 & v_52467;
assign v_52469 = v_52299 & v_52465;
assign v_52471 = v_52297 & v_52470;
assign v_52473 = v_52379 & v_52472;
assign v_52474 = v_52296 & v_52470;
assign v_52476 = v_52294 & v_52475;
assign v_52478 = v_52385 & v_52477;
assign v_52479 = v_52293 & v_52475;
assign v_52481 = v_52291 & v_52480;
assign v_52483 = v_52391 & v_52482;
assign v_52484 = v_52290 & v_52480;
assign v_52486 = v_52288 & v_52485;
assign v_52488 = v_52397 & v_52487;
assign v_52489 = v_52287 & v_52485;
assign v_52491 = v_52285 & v_52490;
assign v_52493 = v_52403 & v_52492;
assign v_52494 = v_52284 & v_52490;
assign v_52496 = v_52282 & v_52495;
assign v_52498 = v_52409 & v_52497;
assign v_52499 = v_52281 & v_52495;
assign v_52501 = v_52279 & v_52500;
assign v_52503 = v_52415 & v_52502;
assign v_52504 = v_52278 & v_52500;
assign v_52506 = v_52276 & v_52505;
assign v_52508 = v_52421 & v_52507;
assign v_52509 = v_52275 & v_52505;
assign v_52511 = v_52510;
assign v_52513 = v_52425 & v_52512;
assign v_52514 = v_52513;
assign v_52516 = v_52515;
assign v_52518 = ~v_2623;
assign v_52519 = ~v_50072;
assign v_52520 = v_50072;
assign v_52521 = ~v_2627;
assign v_52522 = ~v_50076;
assign v_52523 = v_50076;
assign v_52524 = ~v_2631;
assign v_52525 = ~v_50080;
assign v_52526 = v_50080;
assign v_52527 = ~v_2635;
assign v_52528 = ~v_50084;
assign v_52529 = v_50084;
assign v_52530 = ~v_50087;
assign v_52531 = ~v_2640;
assign v_52532 = v_2640;
assign v_52533 = ~v_50091;
assign v_52534 = ~v_2644;
assign v_52535 = v_2644;
assign v_52536 = ~v_50095;
assign v_52537 = ~v_2648;
assign v_52538 = v_2648;
assign v_52539 = ~v_50099;
assign v_52540 = ~v_2652;
assign v_52541 = v_2652;
assign v_52542 = ~v_50103;
assign v_52543 = ~v_2656;
assign v_52544 = v_2656;
assign v_52545 = ~v_50107;
assign v_52546 = ~v_2660;
assign v_52547 = v_2660;
assign v_52548 = ~v_50111;
assign v_52549 = ~v_2664;
assign v_52550 = v_2664;
assign v_52551 = ~v_50115;
assign v_52552 = ~v_2668;
assign v_52553 = v_2668;
assign v_52554 = ~v_50119;
assign v_52555 = ~v_2672;
assign v_52556 = v_2672;
assign v_52557 = ~v_50123;
assign v_52558 = ~v_2676;
assign v_52559 = v_2676;
assign v_52560 = ~v_50127;
assign v_52561 = ~v_2680;
assign v_52562 = v_2680;
assign v_52563 = ~v_50131;
assign v_52564 = ~v_2684;
assign v_52565 = v_2684;
assign v_52566 = ~v_50135;
assign v_52567 = ~v_2688;
assign v_52568 = v_52567;
assign v_52570 = v_52569;
assign v_52572 = v_52564 & v_52571;
assign v_52574 = v_50131;
assign v_52576 = v_52573 & v_52575;
assign v_52578 = v_52561 & v_52577;
assign v_52580 = v_50127;
assign v_52582 = v_52579 & v_52581;
assign v_52584 = v_52558 & v_52583;
assign v_52586 = v_50123;
assign v_52588 = v_52585 & v_52587;
assign v_52590 = v_52555 & v_52589;
assign v_52592 = v_50119;
assign v_52594 = v_52591 & v_52593;
assign v_52596 = v_52552 & v_52595;
assign v_52598 = v_50115;
assign v_52600 = v_52597 & v_52599;
assign v_52602 = v_52549 & v_52601;
assign v_52604 = v_50111;
assign v_52606 = v_52603 & v_52605;
assign v_52608 = v_52546 & v_52607;
assign v_52610 = v_50107;
assign v_52612 = v_52609 & v_52611;
assign v_52614 = v_52543 & v_52613;
assign v_52616 = v_50103;
assign v_52618 = v_52615 & v_52617;
assign v_52620 = v_52540 & v_52619;
assign v_52622 = v_50099;
assign v_52624 = v_52621 & v_52623;
assign v_52626 = v_52537 & v_52625;
assign v_52628 = v_50095;
assign v_52630 = v_52627 & v_52629;
assign v_52632 = v_52534 & v_52631;
assign v_52634 = v_50091;
assign v_52636 = v_52633 & v_52635;
assign v_52638 = v_52531 & v_52637;
assign v_52640 = v_50087;
assign v_52642 = v_52639 & v_52641;
assign v_52644 = v_52528 & v_52643;
assign v_52646 = v_2635;
assign v_52648 = v_52645 & v_52647;
assign v_52650 = v_52525 & v_52649;
assign v_52652 = v_2631;
assign v_52654 = v_52651 & v_52653;
assign v_52656 = v_52522 & v_52655;
assign v_52658 = v_2627;
assign v_52660 = v_52657 & v_52659;
assign v_52662 = v_52519 & v_52661;
assign v_52664 = v_2623;
assign v_52666 = v_52663 & v_52665;
assign v_52667 = v_52666;
assign v_52669 = v_50135;
assign v_52670 = v_2688;
assign v_52671 = v_52670;
assign v_52672 = v_52669 & v_52671;
assign v_52673 = v_52672;
assign v_52674 = v_52564 & v_52673;
assign v_52676 = v_52574 & v_52675;
assign v_52677 = v_52563 & v_52673;
assign v_52679 = v_52561 & v_52678;
assign v_52681 = v_52580 & v_52680;
assign v_52682 = v_52560 & v_52678;
assign v_52684 = v_52558 & v_52683;
assign v_52686 = v_52586 & v_52685;
assign v_52687 = v_52557 & v_52683;
assign v_52689 = v_52555 & v_52688;
assign v_52691 = v_52592 & v_52690;
assign v_52692 = v_52554 & v_52688;
assign v_52694 = v_52552 & v_52693;
assign v_52696 = v_52598 & v_52695;
assign v_52697 = v_52551 & v_52693;
assign v_52699 = v_52549 & v_52698;
assign v_52701 = v_52604 & v_52700;
assign v_52702 = v_52548 & v_52698;
assign v_52704 = v_52546 & v_52703;
assign v_52706 = v_52610 & v_52705;
assign v_52707 = v_52545 & v_52703;
assign v_52709 = v_52543 & v_52708;
assign v_52711 = v_52616 & v_52710;
assign v_52712 = v_52542 & v_52708;
assign v_52714 = v_52540 & v_52713;
assign v_52716 = v_52622 & v_52715;
assign v_52717 = v_52539 & v_52713;
assign v_52719 = v_52537 & v_52718;
assign v_52721 = v_52628 & v_52720;
assign v_52722 = v_52536 & v_52718;
assign v_52724 = v_52534 & v_52723;
assign v_52726 = v_52634 & v_52725;
assign v_52727 = v_52533 & v_52723;
assign v_52729 = v_52531 & v_52728;
assign v_52731 = v_52640 & v_52730;
assign v_52732 = v_52530 & v_52728;
assign v_52734 = v_52528 & v_52733;
assign v_52736 = v_52646 & v_52735;
assign v_52737 = v_52527 & v_52733;
assign v_52739 = v_52525 & v_52738;
assign v_52741 = v_52652 & v_52740;
assign v_52742 = v_52524 & v_52738;
assign v_52744 = v_52522 & v_52743;
assign v_52746 = v_52658 & v_52745;
assign v_52747 = v_52521 & v_52743;
assign v_52749 = v_52519 & v_52748;
assign v_52751 = v_52664 & v_52750;
assign v_52752 = v_52518 & v_52748;
assign v_52754 = v_52753;
assign v_52756 = v_52668 & v_52755;
assign v_52757 = v_52756;
assign v_52759 = v_52758;
assign v_52761 = ~v_2883;
assign v_52762 = ~v_50072;
assign v_52763 = v_50072;
assign v_52764 = ~v_2887;
assign v_52765 = ~v_50076;
assign v_52766 = v_50076;
assign v_52767 = ~v_2891;
assign v_52768 = ~v_50080;
assign v_52769 = v_50080;
assign v_52770 = ~v_2895;
assign v_52771 = ~v_50084;
assign v_52772 = v_50084;
assign v_52773 = ~v_50087;
assign v_52774 = ~v_2900;
assign v_52775 = v_2900;
assign v_52776 = ~v_50091;
assign v_52777 = ~v_2904;
assign v_52778 = v_2904;
assign v_52779 = ~v_50095;
assign v_52780 = ~v_2908;
assign v_52781 = v_2908;
assign v_52782 = ~v_50099;
assign v_52783 = ~v_2912;
assign v_52784 = v_2912;
assign v_52785 = ~v_50103;
assign v_52786 = ~v_2916;
assign v_52787 = v_2916;
assign v_52788 = ~v_50107;
assign v_52789 = ~v_2920;
assign v_52790 = v_2920;
assign v_52791 = ~v_50111;
assign v_52792 = ~v_2924;
assign v_52793 = v_2924;
assign v_52794 = ~v_50115;
assign v_52795 = ~v_2928;
assign v_52796 = v_2928;
assign v_52797 = ~v_50119;
assign v_52798 = ~v_2932;
assign v_52799 = v_2932;
assign v_52800 = ~v_50123;
assign v_52801 = ~v_2936;
assign v_52802 = v_2936;
assign v_52803 = ~v_50127;
assign v_52804 = ~v_2940;
assign v_52805 = v_2940;
assign v_52806 = ~v_50131;
assign v_52807 = ~v_2944;
assign v_52808 = v_2944;
assign v_52809 = ~v_50135;
assign v_52810 = ~v_2948;
assign v_52811 = v_52810;
assign v_52813 = v_52812;
assign v_52815 = v_52807 & v_52814;
assign v_52817 = v_50131;
assign v_52819 = v_52816 & v_52818;
assign v_52821 = v_52804 & v_52820;
assign v_52823 = v_50127;
assign v_52825 = v_52822 & v_52824;
assign v_52827 = v_52801 & v_52826;
assign v_52829 = v_50123;
assign v_52831 = v_52828 & v_52830;
assign v_52833 = v_52798 & v_52832;
assign v_52835 = v_50119;
assign v_52837 = v_52834 & v_52836;
assign v_52839 = v_52795 & v_52838;
assign v_52841 = v_50115;
assign v_52843 = v_52840 & v_52842;
assign v_52845 = v_52792 & v_52844;
assign v_52847 = v_50111;
assign v_52849 = v_52846 & v_52848;
assign v_52851 = v_52789 & v_52850;
assign v_52853 = v_50107;
assign v_52855 = v_52852 & v_52854;
assign v_52857 = v_52786 & v_52856;
assign v_52859 = v_50103;
assign v_52861 = v_52858 & v_52860;
assign v_52863 = v_52783 & v_52862;
assign v_52865 = v_50099;
assign v_52867 = v_52864 & v_52866;
assign v_52869 = v_52780 & v_52868;
assign v_52871 = v_50095;
assign v_52873 = v_52870 & v_52872;
assign v_52875 = v_52777 & v_52874;
assign v_52877 = v_50091;
assign v_52879 = v_52876 & v_52878;
assign v_52881 = v_52774 & v_52880;
assign v_52883 = v_50087;
assign v_52885 = v_52882 & v_52884;
assign v_52887 = v_52771 & v_52886;
assign v_52889 = v_2895;
assign v_52891 = v_52888 & v_52890;
assign v_52893 = v_52768 & v_52892;
assign v_52895 = v_2891;
assign v_52897 = v_52894 & v_52896;
assign v_52899 = v_52765 & v_52898;
assign v_52901 = v_2887;
assign v_52903 = v_52900 & v_52902;
assign v_52905 = v_52762 & v_52904;
assign v_52907 = v_2883;
assign v_52909 = v_52906 & v_52908;
assign v_52910 = v_52909;
assign v_52912 = v_50135;
assign v_52913 = v_2948;
assign v_52914 = v_52913;
assign v_52915 = v_52912 & v_52914;
assign v_52916 = v_52915;
assign v_52917 = v_52807 & v_52916;
assign v_52919 = v_52817 & v_52918;
assign v_52920 = v_52806 & v_52916;
assign v_52922 = v_52804 & v_52921;
assign v_52924 = v_52823 & v_52923;
assign v_52925 = v_52803 & v_52921;
assign v_52927 = v_52801 & v_52926;
assign v_52929 = v_52829 & v_52928;
assign v_52930 = v_52800 & v_52926;
assign v_52932 = v_52798 & v_52931;
assign v_52934 = v_52835 & v_52933;
assign v_52935 = v_52797 & v_52931;
assign v_52937 = v_52795 & v_52936;
assign v_52939 = v_52841 & v_52938;
assign v_52940 = v_52794 & v_52936;
assign v_52942 = v_52792 & v_52941;
assign v_52944 = v_52847 & v_52943;
assign v_52945 = v_52791 & v_52941;
assign v_52947 = v_52789 & v_52946;
assign v_52949 = v_52853 & v_52948;
assign v_52950 = v_52788 & v_52946;
assign v_52952 = v_52786 & v_52951;
assign v_52954 = v_52859 & v_52953;
assign v_52955 = v_52785 & v_52951;
assign v_52957 = v_52783 & v_52956;
assign v_52959 = v_52865 & v_52958;
assign v_52960 = v_52782 & v_52956;
assign v_52962 = v_52780 & v_52961;
assign v_52964 = v_52871 & v_52963;
assign v_52965 = v_52779 & v_52961;
assign v_52967 = v_52777 & v_52966;
assign v_52969 = v_52877 & v_52968;
assign v_52970 = v_52776 & v_52966;
assign v_52972 = v_52774 & v_52971;
assign v_52974 = v_52883 & v_52973;
assign v_52975 = v_52773 & v_52971;
assign v_52977 = v_52771 & v_52976;
assign v_52979 = v_52889 & v_52978;
assign v_52980 = v_52770 & v_52976;
assign v_52982 = v_52768 & v_52981;
assign v_52984 = v_52895 & v_52983;
assign v_52985 = v_52767 & v_52981;
assign v_52987 = v_52765 & v_52986;
assign v_52989 = v_52901 & v_52988;
assign v_52990 = v_52764 & v_52986;
assign v_52992 = v_52762 & v_52991;
assign v_52994 = v_52907 & v_52993;
assign v_52995 = v_52761 & v_52991;
assign v_52997 = v_52996;
assign v_52999 = v_52911 & v_52998;
assign v_53000 = v_52999;
assign v_53002 = v_53001;
assign v_53004 = ~v_3143;
assign v_53005 = ~v_50072;
assign v_53006 = v_50072;
assign v_53007 = ~v_3147;
assign v_53008 = ~v_50076;
assign v_53009 = v_50076;
assign v_53010 = ~v_3151;
assign v_53011 = ~v_50080;
assign v_53012 = v_50080;
assign v_53013 = ~v_3155;
assign v_53014 = ~v_50084;
assign v_53015 = v_50084;
assign v_53016 = ~v_50087;
assign v_53017 = ~v_3160;
assign v_53018 = v_3160;
assign v_53019 = ~v_50091;
assign v_53020 = ~v_3164;
assign v_53021 = v_3164;
assign v_53022 = ~v_50095;
assign v_53023 = ~v_3168;
assign v_53024 = v_3168;
assign v_53025 = ~v_50099;
assign v_53026 = ~v_3172;
assign v_53027 = v_3172;
assign v_53028 = ~v_50103;
assign v_53029 = ~v_3176;
assign v_53030 = v_3176;
assign v_53031 = ~v_50107;
assign v_53032 = ~v_3180;
assign v_53033 = v_3180;
assign v_53034 = ~v_50111;
assign v_53035 = ~v_3184;
assign v_53036 = v_3184;
assign v_53037 = ~v_50115;
assign v_53038 = ~v_3188;
assign v_53039 = v_3188;
assign v_53040 = ~v_50119;
assign v_53041 = ~v_3192;
assign v_53042 = v_3192;
assign v_53043 = ~v_50123;
assign v_53044 = ~v_3196;
assign v_53045 = v_3196;
assign v_53046 = ~v_50127;
assign v_53047 = ~v_3200;
assign v_53048 = v_3200;
assign v_53049 = ~v_50131;
assign v_53050 = ~v_3204;
assign v_53051 = v_3204;
assign v_53052 = ~v_50135;
assign v_53053 = ~v_3208;
assign v_53054 = v_53053;
assign v_53056 = v_53055;
assign v_53058 = v_53050 & v_53057;
assign v_53060 = v_50131;
assign v_53062 = v_53059 & v_53061;
assign v_53064 = v_53047 & v_53063;
assign v_53066 = v_50127;
assign v_53068 = v_53065 & v_53067;
assign v_53070 = v_53044 & v_53069;
assign v_53072 = v_50123;
assign v_53074 = v_53071 & v_53073;
assign v_53076 = v_53041 & v_53075;
assign v_53078 = v_50119;
assign v_53080 = v_53077 & v_53079;
assign v_53082 = v_53038 & v_53081;
assign v_53084 = v_50115;
assign v_53086 = v_53083 & v_53085;
assign v_53088 = v_53035 & v_53087;
assign v_53090 = v_50111;
assign v_53092 = v_53089 & v_53091;
assign v_53094 = v_53032 & v_53093;
assign v_53096 = v_50107;
assign v_53098 = v_53095 & v_53097;
assign v_53100 = v_53029 & v_53099;
assign v_53102 = v_50103;
assign v_53104 = v_53101 & v_53103;
assign v_53106 = v_53026 & v_53105;
assign v_53108 = v_50099;
assign v_53110 = v_53107 & v_53109;
assign v_53112 = v_53023 & v_53111;
assign v_53114 = v_50095;
assign v_53116 = v_53113 & v_53115;
assign v_53118 = v_53020 & v_53117;
assign v_53120 = v_50091;
assign v_53122 = v_53119 & v_53121;
assign v_53124 = v_53017 & v_53123;
assign v_53126 = v_50087;
assign v_53128 = v_53125 & v_53127;
assign v_53130 = v_53014 & v_53129;
assign v_53132 = v_3155;
assign v_53134 = v_53131 & v_53133;
assign v_53136 = v_53011 & v_53135;
assign v_53138 = v_3151;
assign v_53140 = v_53137 & v_53139;
assign v_53142 = v_53008 & v_53141;
assign v_53144 = v_3147;
assign v_53146 = v_53143 & v_53145;
assign v_53148 = v_53005 & v_53147;
assign v_53150 = v_3143;
assign v_53152 = v_53149 & v_53151;
assign v_53153 = v_53152;
assign v_53155 = v_50135;
assign v_53156 = v_3208;
assign v_53157 = v_53156;
assign v_53158 = v_53155 & v_53157;
assign v_53159 = v_53158;
assign v_53160 = v_53050 & v_53159;
assign v_53162 = v_53060 & v_53161;
assign v_53163 = v_53049 & v_53159;
assign v_53165 = v_53047 & v_53164;
assign v_53167 = v_53066 & v_53166;
assign v_53168 = v_53046 & v_53164;
assign v_53170 = v_53044 & v_53169;
assign v_53172 = v_53072 & v_53171;
assign v_53173 = v_53043 & v_53169;
assign v_53175 = v_53041 & v_53174;
assign v_53177 = v_53078 & v_53176;
assign v_53178 = v_53040 & v_53174;
assign v_53180 = v_53038 & v_53179;
assign v_53182 = v_53084 & v_53181;
assign v_53183 = v_53037 & v_53179;
assign v_53185 = v_53035 & v_53184;
assign v_53187 = v_53090 & v_53186;
assign v_53188 = v_53034 & v_53184;
assign v_53190 = v_53032 & v_53189;
assign v_53192 = v_53096 & v_53191;
assign v_53193 = v_53031 & v_53189;
assign v_53195 = v_53029 & v_53194;
assign v_53197 = v_53102 & v_53196;
assign v_53198 = v_53028 & v_53194;
assign v_53200 = v_53026 & v_53199;
assign v_53202 = v_53108 & v_53201;
assign v_53203 = v_53025 & v_53199;
assign v_53205 = v_53023 & v_53204;
assign v_53207 = v_53114 & v_53206;
assign v_53208 = v_53022 & v_53204;
assign v_53210 = v_53020 & v_53209;
assign v_53212 = v_53120 & v_53211;
assign v_53213 = v_53019 & v_53209;
assign v_53215 = v_53017 & v_53214;
assign v_53217 = v_53126 & v_53216;
assign v_53218 = v_53016 & v_53214;
assign v_53220 = v_53014 & v_53219;
assign v_53222 = v_53132 & v_53221;
assign v_53223 = v_53013 & v_53219;
assign v_53225 = v_53011 & v_53224;
assign v_53227 = v_53138 & v_53226;
assign v_53228 = v_53010 & v_53224;
assign v_53230 = v_53008 & v_53229;
assign v_53232 = v_53144 & v_53231;
assign v_53233 = v_53007 & v_53229;
assign v_53235 = v_53005 & v_53234;
assign v_53237 = v_53150 & v_53236;
assign v_53238 = v_53004 & v_53234;
assign v_53240 = v_53239;
assign v_53242 = v_53154 & v_53241;
assign v_53243 = v_53242;
assign v_53245 = v_53244;
assign v_53247 = ~v_3403;
assign v_53248 = ~v_50072;
assign v_53249 = v_50072;
assign v_53250 = ~v_3407;
assign v_53251 = ~v_50076;
assign v_53252 = v_50076;
assign v_53253 = ~v_3411;
assign v_53254 = ~v_50080;
assign v_53255 = v_50080;
assign v_53256 = ~v_3415;
assign v_53257 = ~v_50084;
assign v_53258 = v_50084;
assign v_53259 = ~v_50087;
assign v_53260 = ~v_3420;
assign v_53261 = v_3420;
assign v_53262 = ~v_50091;
assign v_53263 = ~v_3424;
assign v_53264 = v_3424;
assign v_53265 = ~v_50095;
assign v_53266 = ~v_3428;
assign v_53267 = v_3428;
assign v_53268 = ~v_50099;
assign v_53269 = ~v_3432;
assign v_53270 = v_3432;
assign v_53271 = ~v_50103;
assign v_53272 = ~v_3436;
assign v_53273 = v_3436;
assign v_53274 = ~v_50107;
assign v_53275 = ~v_3440;
assign v_53276 = v_3440;
assign v_53277 = ~v_50111;
assign v_53278 = ~v_3444;
assign v_53279 = v_3444;
assign v_53280 = ~v_50115;
assign v_53281 = ~v_3448;
assign v_53282 = v_3448;
assign v_53283 = ~v_50119;
assign v_53284 = ~v_3452;
assign v_53285 = v_3452;
assign v_53286 = ~v_50123;
assign v_53287 = ~v_3456;
assign v_53288 = v_3456;
assign v_53289 = ~v_50127;
assign v_53290 = ~v_3460;
assign v_53291 = v_3460;
assign v_53292 = ~v_50131;
assign v_53293 = ~v_3464;
assign v_53294 = v_3464;
assign v_53295 = ~v_50135;
assign v_53296 = ~v_3468;
assign v_53297 = v_53296;
assign v_53299 = v_53298;
assign v_53301 = v_53293 & v_53300;
assign v_53303 = v_50131;
assign v_53305 = v_53302 & v_53304;
assign v_53307 = v_53290 & v_53306;
assign v_53309 = v_50127;
assign v_53311 = v_53308 & v_53310;
assign v_53313 = v_53287 & v_53312;
assign v_53315 = v_50123;
assign v_53317 = v_53314 & v_53316;
assign v_53319 = v_53284 & v_53318;
assign v_53321 = v_50119;
assign v_53323 = v_53320 & v_53322;
assign v_53325 = v_53281 & v_53324;
assign v_53327 = v_50115;
assign v_53329 = v_53326 & v_53328;
assign v_53331 = v_53278 & v_53330;
assign v_53333 = v_50111;
assign v_53335 = v_53332 & v_53334;
assign v_53337 = v_53275 & v_53336;
assign v_53339 = v_50107;
assign v_53341 = v_53338 & v_53340;
assign v_53343 = v_53272 & v_53342;
assign v_53345 = v_50103;
assign v_53347 = v_53344 & v_53346;
assign v_53349 = v_53269 & v_53348;
assign v_53351 = v_50099;
assign v_53353 = v_53350 & v_53352;
assign v_53355 = v_53266 & v_53354;
assign v_53357 = v_50095;
assign v_53359 = v_53356 & v_53358;
assign v_53361 = v_53263 & v_53360;
assign v_53363 = v_50091;
assign v_53365 = v_53362 & v_53364;
assign v_53367 = v_53260 & v_53366;
assign v_53369 = v_50087;
assign v_53371 = v_53368 & v_53370;
assign v_53373 = v_53257 & v_53372;
assign v_53375 = v_3415;
assign v_53377 = v_53374 & v_53376;
assign v_53379 = v_53254 & v_53378;
assign v_53381 = v_3411;
assign v_53383 = v_53380 & v_53382;
assign v_53385 = v_53251 & v_53384;
assign v_53387 = v_3407;
assign v_53389 = v_53386 & v_53388;
assign v_53391 = v_53248 & v_53390;
assign v_53393 = v_3403;
assign v_53395 = v_53392 & v_53394;
assign v_53396 = v_53395;
assign v_53398 = v_50135;
assign v_53399 = v_3468;
assign v_53400 = v_53399;
assign v_53401 = v_53398 & v_53400;
assign v_53402 = v_53401;
assign v_53403 = v_53293 & v_53402;
assign v_53405 = v_53303 & v_53404;
assign v_53406 = v_53292 & v_53402;
assign v_53408 = v_53290 & v_53407;
assign v_53410 = v_53309 & v_53409;
assign v_53411 = v_53289 & v_53407;
assign v_53413 = v_53287 & v_53412;
assign v_53415 = v_53315 & v_53414;
assign v_53416 = v_53286 & v_53412;
assign v_53418 = v_53284 & v_53417;
assign v_53420 = v_53321 & v_53419;
assign v_53421 = v_53283 & v_53417;
assign v_53423 = v_53281 & v_53422;
assign v_53425 = v_53327 & v_53424;
assign v_53426 = v_53280 & v_53422;
assign v_53428 = v_53278 & v_53427;
assign v_53430 = v_53333 & v_53429;
assign v_53431 = v_53277 & v_53427;
assign v_53433 = v_53275 & v_53432;
assign v_53435 = v_53339 & v_53434;
assign v_53436 = v_53274 & v_53432;
assign v_53438 = v_53272 & v_53437;
assign v_53440 = v_53345 & v_53439;
assign v_53441 = v_53271 & v_53437;
assign v_53443 = v_53269 & v_53442;
assign v_53445 = v_53351 & v_53444;
assign v_53446 = v_53268 & v_53442;
assign v_53448 = v_53266 & v_53447;
assign v_53450 = v_53357 & v_53449;
assign v_53451 = v_53265 & v_53447;
assign v_53453 = v_53263 & v_53452;
assign v_53455 = v_53363 & v_53454;
assign v_53456 = v_53262 & v_53452;
assign v_53458 = v_53260 & v_53457;
assign v_53460 = v_53369 & v_53459;
assign v_53461 = v_53259 & v_53457;
assign v_53463 = v_53257 & v_53462;
assign v_53465 = v_53375 & v_53464;
assign v_53466 = v_53256 & v_53462;
assign v_53468 = v_53254 & v_53467;
assign v_53470 = v_53381 & v_53469;
assign v_53471 = v_53253 & v_53467;
assign v_53473 = v_53251 & v_53472;
assign v_53475 = v_53387 & v_53474;
assign v_53476 = v_53250 & v_53472;
assign v_53478 = v_53248 & v_53477;
assign v_53480 = v_53393 & v_53479;
assign v_53481 = v_53247 & v_53477;
assign v_53483 = v_53482;
assign v_53485 = v_53397 & v_53484;
assign v_53486 = v_53485;
assign v_53488 = v_53487;
assign v_53490 = ~v_3663;
assign v_53491 = ~v_50072;
assign v_53492 = v_50072;
assign v_53493 = ~v_3667;
assign v_53494 = ~v_50076;
assign v_53495 = v_50076;
assign v_53496 = ~v_3671;
assign v_53497 = ~v_50080;
assign v_53498 = v_50080;
assign v_53499 = ~v_3675;
assign v_53500 = ~v_50084;
assign v_53501 = v_50084;
assign v_53502 = ~v_50087;
assign v_53503 = ~v_3680;
assign v_53504 = v_3680;
assign v_53505 = ~v_50091;
assign v_53506 = ~v_3684;
assign v_53507 = v_3684;
assign v_53508 = ~v_50095;
assign v_53509 = ~v_3688;
assign v_53510 = v_3688;
assign v_53511 = ~v_50099;
assign v_53512 = ~v_3692;
assign v_53513 = v_3692;
assign v_53514 = ~v_50103;
assign v_53515 = ~v_3696;
assign v_53516 = v_3696;
assign v_53517 = ~v_50107;
assign v_53518 = ~v_3700;
assign v_53519 = v_3700;
assign v_53520 = ~v_50111;
assign v_53521 = ~v_3704;
assign v_53522 = v_3704;
assign v_53523 = ~v_50115;
assign v_53524 = ~v_3708;
assign v_53525 = v_3708;
assign v_53526 = ~v_50119;
assign v_53527 = ~v_3712;
assign v_53528 = v_3712;
assign v_53529 = ~v_50123;
assign v_53530 = ~v_3716;
assign v_53531 = v_3716;
assign v_53532 = ~v_50127;
assign v_53533 = ~v_3720;
assign v_53534 = v_3720;
assign v_53535 = ~v_50131;
assign v_53536 = ~v_3724;
assign v_53537 = v_3724;
assign v_53538 = ~v_50135;
assign v_53539 = ~v_3728;
assign v_53540 = v_53539;
assign v_53542 = v_53541;
assign v_53544 = v_53536 & v_53543;
assign v_53546 = v_50131;
assign v_53548 = v_53545 & v_53547;
assign v_53550 = v_53533 & v_53549;
assign v_53552 = v_50127;
assign v_53554 = v_53551 & v_53553;
assign v_53556 = v_53530 & v_53555;
assign v_53558 = v_50123;
assign v_53560 = v_53557 & v_53559;
assign v_53562 = v_53527 & v_53561;
assign v_53564 = v_50119;
assign v_53566 = v_53563 & v_53565;
assign v_53568 = v_53524 & v_53567;
assign v_53570 = v_50115;
assign v_53572 = v_53569 & v_53571;
assign v_53574 = v_53521 & v_53573;
assign v_53576 = v_50111;
assign v_53578 = v_53575 & v_53577;
assign v_53580 = v_53518 & v_53579;
assign v_53582 = v_50107;
assign v_53584 = v_53581 & v_53583;
assign v_53586 = v_53515 & v_53585;
assign v_53588 = v_50103;
assign v_53590 = v_53587 & v_53589;
assign v_53592 = v_53512 & v_53591;
assign v_53594 = v_50099;
assign v_53596 = v_53593 & v_53595;
assign v_53598 = v_53509 & v_53597;
assign v_53600 = v_50095;
assign v_53602 = v_53599 & v_53601;
assign v_53604 = v_53506 & v_53603;
assign v_53606 = v_50091;
assign v_53608 = v_53605 & v_53607;
assign v_53610 = v_53503 & v_53609;
assign v_53612 = v_50087;
assign v_53614 = v_53611 & v_53613;
assign v_53616 = v_53500 & v_53615;
assign v_53618 = v_3675;
assign v_53620 = v_53617 & v_53619;
assign v_53622 = v_53497 & v_53621;
assign v_53624 = v_3671;
assign v_53626 = v_53623 & v_53625;
assign v_53628 = v_53494 & v_53627;
assign v_53630 = v_3667;
assign v_53632 = v_53629 & v_53631;
assign v_53634 = v_53491 & v_53633;
assign v_53636 = v_3663;
assign v_53638 = v_53635 & v_53637;
assign v_53639 = v_53638;
assign v_53641 = v_50135;
assign v_53642 = v_3728;
assign v_53643 = v_53642;
assign v_53644 = v_53641 & v_53643;
assign v_53645 = v_53644;
assign v_53646 = v_53536 & v_53645;
assign v_53648 = v_53546 & v_53647;
assign v_53649 = v_53535 & v_53645;
assign v_53651 = v_53533 & v_53650;
assign v_53653 = v_53552 & v_53652;
assign v_53654 = v_53532 & v_53650;
assign v_53656 = v_53530 & v_53655;
assign v_53658 = v_53558 & v_53657;
assign v_53659 = v_53529 & v_53655;
assign v_53661 = v_53527 & v_53660;
assign v_53663 = v_53564 & v_53662;
assign v_53664 = v_53526 & v_53660;
assign v_53666 = v_53524 & v_53665;
assign v_53668 = v_53570 & v_53667;
assign v_53669 = v_53523 & v_53665;
assign v_53671 = v_53521 & v_53670;
assign v_53673 = v_53576 & v_53672;
assign v_53674 = v_53520 & v_53670;
assign v_53676 = v_53518 & v_53675;
assign v_53678 = v_53582 & v_53677;
assign v_53679 = v_53517 & v_53675;
assign v_53681 = v_53515 & v_53680;
assign v_53683 = v_53588 & v_53682;
assign v_53684 = v_53514 & v_53680;
assign v_53686 = v_53512 & v_53685;
assign v_53688 = v_53594 & v_53687;
assign v_53689 = v_53511 & v_53685;
assign v_53691 = v_53509 & v_53690;
assign v_53693 = v_53600 & v_53692;
assign v_53694 = v_53508 & v_53690;
assign v_53696 = v_53506 & v_53695;
assign v_53698 = v_53606 & v_53697;
assign v_53699 = v_53505 & v_53695;
assign v_53701 = v_53503 & v_53700;
assign v_53703 = v_53612 & v_53702;
assign v_53704 = v_53502 & v_53700;
assign v_53706 = v_53500 & v_53705;
assign v_53708 = v_53618 & v_53707;
assign v_53709 = v_53499 & v_53705;
assign v_53711 = v_53497 & v_53710;
assign v_53713 = v_53624 & v_53712;
assign v_53714 = v_53496 & v_53710;
assign v_53716 = v_53494 & v_53715;
assign v_53718 = v_53630 & v_53717;
assign v_53719 = v_53493 & v_53715;
assign v_53721 = v_53491 & v_53720;
assign v_53723 = v_53636 & v_53722;
assign v_53724 = v_53490 & v_53720;
assign v_53726 = v_53725;
assign v_53728 = v_53640 & v_53727;
assign v_53729 = v_53728;
assign v_53731 = v_53730;
assign v_53733 = ~v_3923;
assign v_53734 = ~v_50072;
assign v_53735 = v_50072;
assign v_53736 = ~v_3927;
assign v_53737 = ~v_50076;
assign v_53738 = v_50076;
assign v_53739 = ~v_3931;
assign v_53740 = ~v_50080;
assign v_53741 = v_50080;
assign v_53742 = ~v_3935;
assign v_53743 = ~v_50084;
assign v_53744 = v_50084;
assign v_53745 = ~v_50087;
assign v_53746 = ~v_3940;
assign v_53747 = v_3940;
assign v_53748 = ~v_50091;
assign v_53749 = ~v_3944;
assign v_53750 = v_3944;
assign v_53751 = ~v_50095;
assign v_53752 = ~v_3948;
assign v_53753 = v_3948;
assign v_53754 = ~v_50099;
assign v_53755 = ~v_3952;
assign v_53756 = v_3952;
assign v_53757 = ~v_50103;
assign v_53758 = ~v_3956;
assign v_53759 = v_3956;
assign v_53760 = ~v_50107;
assign v_53761 = ~v_3960;
assign v_53762 = v_3960;
assign v_53763 = ~v_50111;
assign v_53764 = ~v_3964;
assign v_53765 = v_3964;
assign v_53766 = ~v_50115;
assign v_53767 = ~v_3968;
assign v_53768 = v_3968;
assign v_53769 = ~v_50119;
assign v_53770 = ~v_3972;
assign v_53771 = v_3972;
assign v_53772 = ~v_50123;
assign v_53773 = ~v_3976;
assign v_53774 = v_3976;
assign v_53775 = ~v_50127;
assign v_53776 = ~v_3980;
assign v_53777 = v_3980;
assign v_53778 = ~v_50131;
assign v_53779 = ~v_3984;
assign v_53780 = v_3984;
assign v_53781 = ~v_50135;
assign v_53782 = ~v_3988;
assign v_53783 = v_53782;
assign v_53785 = v_53784;
assign v_53787 = v_53779 & v_53786;
assign v_53789 = v_50131;
assign v_53791 = v_53788 & v_53790;
assign v_53793 = v_53776 & v_53792;
assign v_53795 = v_50127;
assign v_53797 = v_53794 & v_53796;
assign v_53799 = v_53773 & v_53798;
assign v_53801 = v_50123;
assign v_53803 = v_53800 & v_53802;
assign v_53805 = v_53770 & v_53804;
assign v_53807 = v_50119;
assign v_53809 = v_53806 & v_53808;
assign v_53811 = v_53767 & v_53810;
assign v_53813 = v_50115;
assign v_53815 = v_53812 & v_53814;
assign v_53817 = v_53764 & v_53816;
assign v_53819 = v_50111;
assign v_53821 = v_53818 & v_53820;
assign v_53823 = v_53761 & v_53822;
assign v_53825 = v_50107;
assign v_53827 = v_53824 & v_53826;
assign v_53829 = v_53758 & v_53828;
assign v_53831 = v_50103;
assign v_53833 = v_53830 & v_53832;
assign v_53835 = v_53755 & v_53834;
assign v_53837 = v_50099;
assign v_53839 = v_53836 & v_53838;
assign v_53841 = v_53752 & v_53840;
assign v_53843 = v_50095;
assign v_53845 = v_53842 & v_53844;
assign v_53847 = v_53749 & v_53846;
assign v_53849 = v_50091;
assign v_53851 = v_53848 & v_53850;
assign v_53853 = v_53746 & v_53852;
assign v_53855 = v_50087;
assign v_53857 = v_53854 & v_53856;
assign v_53859 = v_53743 & v_53858;
assign v_53861 = v_3935;
assign v_53863 = v_53860 & v_53862;
assign v_53865 = v_53740 & v_53864;
assign v_53867 = v_3931;
assign v_53869 = v_53866 & v_53868;
assign v_53871 = v_53737 & v_53870;
assign v_53873 = v_3927;
assign v_53875 = v_53872 & v_53874;
assign v_53877 = v_53734 & v_53876;
assign v_53879 = v_3923;
assign v_53881 = v_53878 & v_53880;
assign v_53882 = v_53881;
assign v_53884 = v_50135;
assign v_53885 = v_3988;
assign v_53886 = v_53885;
assign v_53887 = v_53884 & v_53886;
assign v_53888 = v_53887;
assign v_53889 = v_53779 & v_53888;
assign v_53891 = v_53789 & v_53890;
assign v_53892 = v_53778 & v_53888;
assign v_53894 = v_53776 & v_53893;
assign v_53896 = v_53795 & v_53895;
assign v_53897 = v_53775 & v_53893;
assign v_53899 = v_53773 & v_53898;
assign v_53901 = v_53801 & v_53900;
assign v_53902 = v_53772 & v_53898;
assign v_53904 = v_53770 & v_53903;
assign v_53906 = v_53807 & v_53905;
assign v_53907 = v_53769 & v_53903;
assign v_53909 = v_53767 & v_53908;
assign v_53911 = v_53813 & v_53910;
assign v_53912 = v_53766 & v_53908;
assign v_53914 = v_53764 & v_53913;
assign v_53916 = v_53819 & v_53915;
assign v_53917 = v_53763 & v_53913;
assign v_53919 = v_53761 & v_53918;
assign v_53921 = v_53825 & v_53920;
assign v_53922 = v_53760 & v_53918;
assign v_53924 = v_53758 & v_53923;
assign v_53926 = v_53831 & v_53925;
assign v_53927 = v_53757 & v_53923;
assign v_53929 = v_53755 & v_53928;
assign v_53931 = v_53837 & v_53930;
assign v_53932 = v_53754 & v_53928;
assign v_53934 = v_53752 & v_53933;
assign v_53936 = v_53843 & v_53935;
assign v_53937 = v_53751 & v_53933;
assign v_53939 = v_53749 & v_53938;
assign v_53941 = v_53849 & v_53940;
assign v_53942 = v_53748 & v_53938;
assign v_53944 = v_53746 & v_53943;
assign v_53946 = v_53855 & v_53945;
assign v_53947 = v_53745 & v_53943;
assign v_53949 = v_53743 & v_53948;
assign v_53951 = v_53861 & v_53950;
assign v_53952 = v_53742 & v_53948;
assign v_53954 = v_53740 & v_53953;
assign v_53956 = v_53867 & v_53955;
assign v_53957 = v_53739 & v_53953;
assign v_53959 = v_53737 & v_53958;
assign v_53961 = v_53873 & v_53960;
assign v_53962 = v_53736 & v_53958;
assign v_53964 = v_53734 & v_53963;
assign v_53966 = v_53879 & v_53965;
assign v_53967 = v_53733 & v_53963;
assign v_53969 = v_53968;
assign v_53971 = v_53883 & v_53970;
assign v_53972 = v_53971;
assign v_53974 = v_53973;
assign v_53975 = ~v_4182;
assign v_53976 = ~v_50072;
assign v_53977 = v_50072;
assign v_53978 = ~v_4186;
assign v_53979 = ~v_50076;
assign v_53980 = v_50076;
assign v_53981 = ~v_4190;
assign v_53982 = ~v_50080;
assign v_53983 = v_50080;
assign v_53984 = ~v_4194;
assign v_53985 = ~v_50084;
assign v_53986 = v_50084;
assign v_53987 = ~v_50087;
assign v_53988 = ~v_4199;
assign v_53989 = v_4199;
assign v_53990 = ~v_50091;
assign v_53991 = ~v_4203;
assign v_53992 = v_4203;
assign v_53993 = ~v_50095;
assign v_53994 = ~v_4207;
assign v_53995 = v_4207;
assign v_53996 = ~v_50099;
assign v_53997 = ~v_4211;
assign v_53998 = v_4211;
assign v_53999 = ~v_50103;
assign v_54000 = ~v_4215;
assign v_54001 = v_4215;
assign v_54002 = ~v_50107;
assign v_54003 = ~v_4219;
assign v_54004 = v_4219;
assign v_54005 = ~v_50111;
assign v_54006 = ~v_4223;
assign v_54007 = v_4223;
assign v_54008 = ~v_50115;
assign v_54009 = ~v_4227;
assign v_54010 = v_4227;
assign v_54011 = ~v_50119;
assign v_54012 = ~v_4231;
assign v_54013 = v_4231;
assign v_54014 = ~v_50123;
assign v_54015 = ~v_4235;
assign v_54016 = v_4235;
assign v_54017 = ~v_50127;
assign v_54018 = ~v_4239;
assign v_54019 = v_4239;
assign v_54020 = ~v_50131;
assign v_54021 = ~v_4243;
assign v_54022 = v_4243;
assign v_54023 = ~v_50135;
assign v_54024 = ~v_4247;
assign v_54025 = v_54024;
assign v_54027 = v_54026;
assign v_54029 = v_54021 & v_54028;
assign v_54031 = v_50131;
assign v_54033 = v_54030 & v_54032;
assign v_54035 = v_54018 & v_54034;
assign v_54037 = v_50127;
assign v_54039 = v_54036 & v_54038;
assign v_54041 = v_54015 & v_54040;
assign v_54043 = v_50123;
assign v_54045 = v_54042 & v_54044;
assign v_54047 = v_54012 & v_54046;
assign v_54049 = v_50119;
assign v_54051 = v_54048 & v_54050;
assign v_54053 = v_54009 & v_54052;
assign v_54055 = v_50115;
assign v_54057 = v_54054 & v_54056;
assign v_54059 = v_54006 & v_54058;
assign v_54061 = v_50111;
assign v_54063 = v_54060 & v_54062;
assign v_54065 = v_54003 & v_54064;
assign v_54067 = v_50107;
assign v_54069 = v_54066 & v_54068;
assign v_54071 = v_54000 & v_54070;
assign v_54073 = v_50103;
assign v_54075 = v_54072 & v_54074;
assign v_54077 = v_53997 & v_54076;
assign v_54079 = v_50099;
assign v_54081 = v_54078 & v_54080;
assign v_54083 = v_53994 & v_54082;
assign v_54085 = v_50095;
assign v_54087 = v_54084 & v_54086;
assign v_54089 = v_53991 & v_54088;
assign v_54091 = v_50091;
assign v_54093 = v_54090 & v_54092;
assign v_54095 = v_53988 & v_54094;
assign v_54097 = v_50087;
assign v_54099 = v_54096 & v_54098;
assign v_54101 = v_53985 & v_54100;
assign v_54103 = v_4194;
assign v_54105 = v_54102 & v_54104;
assign v_54107 = v_53982 & v_54106;
assign v_54109 = v_4190;
assign v_54111 = v_54108 & v_54110;
assign v_54113 = v_53979 & v_54112;
assign v_54115 = v_4186;
assign v_54117 = v_54114 & v_54116;
assign v_54119 = v_53976 & v_54118;
assign v_54121 = v_4182;
assign v_54123 = v_54120 & v_54122;
assign v_54125 = ~v_54124;
assign v_54127 = v_50135;
assign v_54128 = v_4247;
assign v_54129 = v_54128;
assign v_54130 = v_54127 & v_54129;
assign v_54131 = v_54130;
assign v_54132 = v_54021 & v_54131;
assign v_54134 = v_54031 & v_54133;
assign v_54135 = v_54020 & v_54131;
assign v_54137 = v_54018 & v_54136;
assign v_54139 = v_54037 & v_54138;
assign v_54140 = v_54017 & v_54136;
assign v_54142 = v_54015 & v_54141;
assign v_54144 = v_54043 & v_54143;
assign v_54145 = v_54014 & v_54141;
assign v_54147 = v_54012 & v_54146;
assign v_54149 = v_54049 & v_54148;
assign v_54150 = v_54011 & v_54146;
assign v_54152 = v_54009 & v_54151;
assign v_54154 = v_54055 & v_54153;
assign v_54155 = v_54008 & v_54151;
assign v_54157 = v_54006 & v_54156;
assign v_54159 = v_54061 & v_54158;
assign v_54160 = v_54005 & v_54156;
assign v_54162 = v_54003 & v_54161;
assign v_54164 = v_54067 & v_54163;
assign v_54165 = v_54002 & v_54161;
assign v_54167 = v_54000 & v_54166;
assign v_54169 = v_54073 & v_54168;
assign v_54170 = v_53999 & v_54166;
assign v_54172 = v_53997 & v_54171;
assign v_54174 = v_54079 & v_54173;
assign v_54175 = v_53996 & v_54171;
assign v_54177 = v_53994 & v_54176;
assign v_54179 = v_54085 & v_54178;
assign v_54180 = v_53993 & v_54176;
assign v_54182 = v_53991 & v_54181;
assign v_54184 = v_54091 & v_54183;
assign v_54185 = v_53990 & v_54181;
assign v_54187 = v_53988 & v_54186;
assign v_54189 = v_54097 & v_54188;
assign v_54190 = v_53987 & v_54186;
assign v_54192 = v_53985 & v_54191;
assign v_54194 = v_54103 & v_54193;
assign v_54195 = v_53984 & v_54191;
assign v_54197 = v_53982 & v_54196;
assign v_54199 = v_54109 & v_54198;
assign v_54200 = v_53981 & v_54196;
assign v_54202 = v_53979 & v_54201;
assign v_54204 = v_54115 & v_54203;
assign v_54205 = v_53978 & v_54201;
assign v_54207 = v_53976 & v_54206;
assign v_54209 = v_54121 & v_54208;
assign v_54210 = v_53975 & v_54206;
assign v_54212 = v_54124;
assign v_54214 = v_54126 & v_54213;
assign v_54215 = v_54214;
assign v_54217 = v_54216;
assign v_54219 = ~v_6;
assign v_54221 = ~v_54220;
assign v_54222 = v_54220;
assign v_54223 = ~v_13;
assign v_54225 = ~v_54224;
assign v_54226 = v_54224;
assign v_54227 = ~v_18;
assign v_54229 = ~v_54228;
assign v_54230 = v_54228;
assign v_54231 = ~v_23;
assign v_54233 = ~v_54232;
assign v_54234 = v_54232;
assign v_54236 = ~v_54235;
assign v_54237 = ~v_30;
assign v_54238 = v_30;
assign v_54240 = ~v_54239;
assign v_54241 = ~v_35;
assign v_54242 = v_35;
assign v_54244 = ~v_54243;
assign v_54245 = ~v_40;
assign v_54246 = v_40;
assign v_54248 = ~v_54247;
assign v_54249 = ~v_45;
assign v_54250 = v_45;
assign v_54252 = ~v_54251;
assign v_54253 = ~v_50;
assign v_54254 = v_50;
assign v_54256 = ~v_54255;
assign v_54257 = ~v_55;
assign v_54258 = v_55;
assign v_54260 = ~v_54259;
assign v_54261 = ~v_60;
assign v_54262 = v_60;
assign v_54264 = ~v_54263;
assign v_54265 = ~v_65;
assign v_54266 = v_65;
assign v_54268 = ~v_54267;
assign v_54269 = ~v_70;
assign v_54270 = v_70;
assign v_54272 = ~v_54271;
assign v_54273 = ~v_75;
assign v_54274 = v_75;
assign v_54276 = ~v_54275;
assign v_54277 = ~v_80;
assign v_54278 = v_80;
assign v_54280 = ~v_54279;
assign v_54281 = ~v_85;
assign v_54282 = v_85;
assign v_54284 = ~v_54283;
assign v_54285 = ~v_90;
assign v_54286 = v_54285;
assign v_54288 = v_54287;
assign v_54290 = v_54281 & v_54289;
assign v_54292 = v_54279;
assign v_54294 = v_54291 & v_54293;
assign v_54296 = v_54277 & v_54295;
assign v_54298 = v_54275;
assign v_54300 = v_54297 & v_54299;
assign v_54302 = v_54273 & v_54301;
assign v_54304 = v_54271;
assign v_54306 = v_54303 & v_54305;
assign v_54308 = v_54269 & v_54307;
assign v_54310 = v_54267;
assign v_54312 = v_54309 & v_54311;
assign v_54314 = v_54265 & v_54313;
assign v_54316 = v_54263;
assign v_54318 = v_54315 & v_54317;
assign v_54320 = v_54261 & v_54319;
assign v_54322 = v_54259;
assign v_54324 = v_54321 & v_54323;
assign v_54326 = v_54257 & v_54325;
assign v_54328 = v_54255;
assign v_54330 = v_54327 & v_54329;
assign v_54332 = v_54253 & v_54331;
assign v_54334 = v_54251;
assign v_54336 = v_54333 & v_54335;
assign v_54338 = v_54249 & v_54337;
assign v_54340 = v_54247;
assign v_54342 = v_54339 & v_54341;
assign v_54344 = v_54245 & v_54343;
assign v_54346 = v_54243;
assign v_54348 = v_54345 & v_54347;
assign v_54350 = v_54241 & v_54349;
assign v_54352 = v_54239;
assign v_54354 = v_54351 & v_54353;
assign v_54356 = v_54237 & v_54355;
assign v_54358 = v_54235;
assign v_54360 = v_54357 & v_54359;
assign v_54362 = v_54233 & v_54361;
assign v_54364 = v_23;
assign v_54366 = v_54363 & v_54365;
assign v_54368 = v_54229 & v_54367;
assign v_54370 = v_18;
assign v_54372 = v_54369 & v_54371;
assign v_54374 = v_54225 & v_54373;
assign v_54376 = v_13;
assign v_54378 = v_54375 & v_54377;
assign v_54380 = v_54221 & v_54379;
assign v_54382 = v_6;
assign v_54384 = v_54381 & v_54383;
assign v_54385 = v_54384;
assign v_54387 = v_54283;
assign v_54388 = v_90;
assign v_54389 = v_54388;
assign v_54390 = v_54387 & v_54389;
assign v_54391 = v_54390;
assign v_54392 = v_54281 & v_54391;
assign v_54394 = v_54292 & v_54393;
assign v_54395 = v_54280 & v_54391;
assign v_54397 = v_54277 & v_54396;
assign v_54399 = v_54298 & v_54398;
assign v_54400 = v_54276 & v_54396;
assign v_54402 = v_54273 & v_54401;
assign v_54404 = v_54304 & v_54403;
assign v_54405 = v_54272 & v_54401;
assign v_54407 = v_54269 & v_54406;
assign v_54409 = v_54310 & v_54408;
assign v_54410 = v_54268 & v_54406;
assign v_54412 = v_54265 & v_54411;
assign v_54414 = v_54316 & v_54413;
assign v_54415 = v_54264 & v_54411;
assign v_54417 = v_54261 & v_54416;
assign v_54419 = v_54322 & v_54418;
assign v_54420 = v_54260 & v_54416;
assign v_54422 = v_54257 & v_54421;
assign v_54424 = v_54328 & v_54423;
assign v_54425 = v_54256 & v_54421;
assign v_54427 = v_54253 & v_54426;
assign v_54429 = v_54334 & v_54428;
assign v_54430 = v_54252 & v_54426;
assign v_54432 = v_54249 & v_54431;
assign v_54434 = v_54340 & v_54433;
assign v_54435 = v_54248 & v_54431;
assign v_54437 = v_54245 & v_54436;
assign v_54439 = v_54346 & v_54438;
assign v_54440 = v_54244 & v_54436;
assign v_54442 = v_54241 & v_54441;
assign v_54444 = v_54352 & v_54443;
assign v_54445 = v_54240 & v_54441;
assign v_54447 = v_54237 & v_54446;
assign v_54449 = v_54358 & v_54448;
assign v_54450 = v_54236 & v_54446;
assign v_54452 = v_54233 & v_54451;
assign v_54454 = v_54364 & v_54453;
assign v_54455 = v_54231 & v_54451;
assign v_54457 = v_54229 & v_54456;
assign v_54459 = v_54370 & v_54458;
assign v_54460 = v_54227 & v_54456;
assign v_54462 = v_54225 & v_54461;
assign v_54464 = v_54376 & v_54463;
assign v_54465 = v_54223 & v_54461;
assign v_54467 = v_54221 & v_54466;
assign v_54469 = v_54382 & v_54468;
assign v_54470 = v_54219 & v_54466;
assign v_54472 = v_54471;
assign v_54474 = v_54386 & v_54473;
assign v_54475 = v_54474;
assign v_54477 = v_54476;
assign v_54479 = ~v_283;
assign v_54480 = ~v_54220;
assign v_54481 = v_54220;
assign v_54482 = ~v_287;
assign v_54483 = ~v_54224;
assign v_54484 = v_54224;
assign v_54485 = ~v_291;
assign v_54486 = ~v_54228;
assign v_54487 = v_54228;
assign v_54488 = ~v_295;
assign v_54489 = ~v_54232;
assign v_54490 = v_54232;
assign v_54491 = ~v_54235;
assign v_54492 = ~v_300;
assign v_54493 = v_300;
assign v_54494 = ~v_54239;
assign v_54495 = ~v_304;
assign v_54496 = v_304;
assign v_54497 = ~v_54243;
assign v_54498 = ~v_308;
assign v_54499 = v_308;
assign v_54500 = ~v_54247;
assign v_54501 = ~v_312;
assign v_54502 = v_312;
assign v_54503 = ~v_54251;
assign v_54504 = ~v_316;
assign v_54505 = v_316;
assign v_54506 = ~v_54255;
assign v_54507 = ~v_320;
assign v_54508 = v_320;
assign v_54509 = ~v_54259;
assign v_54510 = ~v_324;
assign v_54511 = v_324;
assign v_54512 = ~v_54263;
assign v_54513 = ~v_328;
assign v_54514 = v_328;
assign v_54515 = ~v_54267;
assign v_54516 = ~v_332;
assign v_54517 = v_332;
assign v_54518 = ~v_54271;
assign v_54519 = ~v_336;
assign v_54520 = v_336;
assign v_54521 = ~v_54275;
assign v_54522 = ~v_340;
assign v_54523 = v_340;
assign v_54524 = ~v_54279;
assign v_54525 = ~v_344;
assign v_54526 = v_344;
assign v_54527 = ~v_54283;
assign v_54528 = ~v_348;
assign v_54529 = v_54528;
assign v_54531 = v_54530;
assign v_54533 = v_54525 & v_54532;
assign v_54535 = v_54279;
assign v_54537 = v_54534 & v_54536;
assign v_54539 = v_54522 & v_54538;
assign v_54541 = v_54275;
assign v_54543 = v_54540 & v_54542;
assign v_54545 = v_54519 & v_54544;
assign v_54547 = v_54271;
assign v_54549 = v_54546 & v_54548;
assign v_54551 = v_54516 & v_54550;
assign v_54553 = v_54267;
assign v_54555 = v_54552 & v_54554;
assign v_54557 = v_54513 & v_54556;
assign v_54559 = v_54263;
assign v_54561 = v_54558 & v_54560;
assign v_54563 = v_54510 & v_54562;
assign v_54565 = v_54259;
assign v_54567 = v_54564 & v_54566;
assign v_54569 = v_54507 & v_54568;
assign v_54571 = v_54255;
assign v_54573 = v_54570 & v_54572;
assign v_54575 = v_54504 & v_54574;
assign v_54577 = v_54251;
assign v_54579 = v_54576 & v_54578;
assign v_54581 = v_54501 & v_54580;
assign v_54583 = v_54247;
assign v_54585 = v_54582 & v_54584;
assign v_54587 = v_54498 & v_54586;
assign v_54589 = v_54243;
assign v_54591 = v_54588 & v_54590;
assign v_54593 = v_54495 & v_54592;
assign v_54595 = v_54239;
assign v_54597 = v_54594 & v_54596;
assign v_54599 = v_54492 & v_54598;
assign v_54601 = v_54235;
assign v_54603 = v_54600 & v_54602;
assign v_54605 = v_54489 & v_54604;
assign v_54607 = v_295;
assign v_54609 = v_54606 & v_54608;
assign v_54611 = v_54486 & v_54610;
assign v_54613 = v_291;
assign v_54615 = v_54612 & v_54614;
assign v_54617 = v_54483 & v_54616;
assign v_54619 = v_287;
assign v_54621 = v_54618 & v_54620;
assign v_54623 = v_54480 & v_54622;
assign v_54625 = v_283;
assign v_54627 = v_54624 & v_54626;
assign v_54628 = v_54627;
assign v_54630 = v_54283;
assign v_54631 = v_348;
assign v_54632 = v_54631;
assign v_54633 = v_54630 & v_54632;
assign v_54634 = v_54633;
assign v_54635 = v_54525 & v_54634;
assign v_54637 = v_54535 & v_54636;
assign v_54638 = v_54524 & v_54634;
assign v_54640 = v_54522 & v_54639;
assign v_54642 = v_54541 & v_54641;
assign v_54643 = v_54521 & v_54639;
assign v_54645 = v_54519 & v_54644;
assign v_54647 = v_54547 & v_54646;
assign v_54648 = v_54518 & v_54644;
assign v_54650 = v_54516 & v_54649;
assign v_54652 = v_54553 & v_54651;
assign v_54653 = v_54515 & v_54649;
assign v_54655 = v_54513 & v_54654;
assign v_54657 = v_54559 & v_54656;
assign v_54658 = v_54512 & v_54654;
assign v_54660 = v_54510 & v_54659;
assign v_54662 = v_54565 & v_54661;
assign v_54663 = v_54509 & v_54659;
assign v_54665 = v_54507 & v_54664;
assign v_54667 = v_54571 & v_54666;
assign v_54668 = v_54506 & v_54664;
assign v_54670 = v_54504 & v_54669;
assign v_54672 = v_54577 & v_54671;
assign v_54673 = v_54503 & v_54669;
assign v_54675 = v_54501 & v_54674;
assign v_54677 = v_54583 & v_54676;
assign v_54678 = v_54500 & v_54674;
assign v_54680 = v_54498 & v_54679;
assign v_54682 = v_54589 & v_54681;
assign v_54683 = v_54497 & v_54679;
assign v_54685 = v_54495 & v_54684;
assign v_54687 = v_54595 & v_54686;
assign v_54688 = v_54494 & v_54684;
assign v_54690 = v_54492 & v_54689;
assign v_54692 = v_54601 & v_54691;
assign v_54693 = v_54491 & v_54689;
assign v_54695 = v_54489 & v_54694;
assign v_54697 = v_54607 & v_54696;
assign v_54698 = v_54488 & v_54694;
assign v_54700 = v_54486 & v_54699;
assign v_54702 = v_54613 & v_54701;
assign v_54703 = v_54485 & v_54699;
assign v_54705 = v_54483 & v_54704;
assign v_54707 = v_54619 & v_54706;
assign v_54708 = v_54482 & v_54704;
assign v_54710 = v_54480 & v_54709;
assign v_54712 = v_54625 & v_54711;
assign v_54713 = v_54479 & v_54709;
assign v_54715 = v_54714;
assign v_54717 = v_54629 & v_54716;
assign v_54718 = v_54717;
assign v_54720 = v_54719;
assign v_54722 = ~v_543;
assign v_54723 = ~v_54220;
assign v_54724 = v_54220;
assign v_54725 = ~v_547;
assign v_54726 = ~v_54224;
assign v_54727 = v_54224;
assign v_54728 = ~v_551;
assign v_54729 = ~v_54228;
assign v_54730 = v_54228;
assign v_54731 = ~v_555;
assign v_54732 = ~v_54232;
assign v_54733 = v_54232;
assign v_54734 = ~v_54235;
assign v_54735 = ~v_560;
assign v_54736 = v_560;
assign v_54737 = ~v_54239;
assign v_54738 = ~v_564;
assign v_54739 = v_564;
assign v_54740 = ~v_54243;
assign v_54741 = ~v_568;
assign v_54742 = v_568;
assign v_54743 = ~v_54247;
assign v_54744 = ~v_572;
assign v_54745 = v_572;
assign v_54746 = ~v_54251;
assign v_54747 = ~v_576;
assign v_54748 = v_576;
assign v_54749 = ~v_54255;
assign v_54750 = ~v_580;
assign v_54751 = v_580;
assign v_54752 = ~v_54259;
assign v_54753 = ~v_584;
assign v_54754 = v_584;
assign v_54755 = ~v_54263;
assign v_54756 = ~v_588;
assign v_54757 = v_588;
assign v_54758 = ~v_54267;
assign v_54759 = ~v_592;
assign v_54760 = v_592;
assign v_54761 = ~v_54271;
assign v_54762 = ~v_596;
assign v_54763 = v_596;
assign v_54764 = ~v_54275;
assign v_54765 = ~v_600;
assign v_54766 = v_600;
assign v_54767 = ~v_54279;
assign v_54768 = ~v_604;
assign v_54769 = v_604;
assign v_54770 = ~v_54283;
assign v_54771 = ~v_608;
assign v_54772 = v_54771;
assign v_54774 = v_54773;
assign v_54776 = v_54768 & v_54775;
assign v_54778 = v_54279;
assign v_54780 = v_54777 & v_54779;
assign v_54782 = v_54765 & v_54781;
assign v_54784 = v_54275;
assign v_54786 = v_54783 & v_54785;
assign v_54788 = v_54762 & v_54787;
assign v_54790 = v_54271;
assign v_54792 = v_54789 & v_54791;
assign v_54794 = v_54759 & v_54793;
assign v_54796 = v_54267;
assign v_54798 = v_54795 & v_54797;
assign v_54800 = v_54756 & v_54799;
assign v_54802 = v_54263;
assign v_54804 = v_54801 & v_54803;
assign v_54806 = v_54753 & v_54805;
assign v_54808 = v_54259;
assign v_54810 = v_54807 & v_54809;
assign v_54812 = v_54750 & v_54811;
assign v_54814 = v_54255;
assign v_54816 = v_54813 & v_54815;
assign v_54818 = v_54747 & v_54817;
assign v_54820 = v_54251;
assign v_54822 = v_54819 & v_54821;
assign v_54824 = v_54744 & v_54823;
assign v_54826 = v_54247;
assign v_54828 = v_54825 & v_54827;
assign v_54830 = v_54741 & v_54829;
assign v_54832 = v_54243;
assign v_54834 = v_54831 & v_54833;
assign v_54836 = v_54738 & v_54835;
assign v_54838 = v_54239;
assign v_54840 = v_54837 & v_54839;
assign v_54842 = v_54735 & v_54841;
assign v_54844 = v_54235;
assign v_54846 = v_54843 & v_54845;
assign v_54848 = v_54732 & v_54847;
assign v_54850 = v_555;
assign v_54852 = v_54849 & v_54851;
assign v_54854 = v_54729 & v_54853;
assign v_54856 = v_551;
assign v_54858 = v_54855 & v_54857;
assign v_54860 = v_54726 & v_54859;
assign v_54862 = v_547;
assign v_54864 = v_54861 & v_54863;
assign v_54866 = v_54723 & v_54865;
assign v_54868 = v_543;
assign v_54870 = v_54867 & v_54869;
assign v_54871 = v_54870;
assign v_54873 = v_54283;
assign v_54874 = v_608;
assign v_54875 = v_54874;
assign v_54876 = v_54873 & v_54875;
assign v_54877 = v_54876;
assign v_54878 = v_54768 & v_54877;
assign v_54880 = v_54778 & v_54879;
assign v_54881 = v_54767 & v_54877;
assign v_54883 = v_54765 & v_54882;
assign v_54885 = v_54784 & v_54884;
assign v_54886 = v_54764 & v_54882;
assign v_54888 = v_54762 & v_54887;
assign v_54890 = v_54790 & v_54889;
assign v_54891 = v_54761 & v_54887;
assign v_54893 = v_54759 & v_54892;
assign v_54895 = v_54796 & v_54894;
assign v_54896 = v_54758 & v_54892;
assign v_54898 = v_54756 & v_54897;
assign v_54900 = v_54802 & v_54899;
assign v_54901 = v_54755 & v_54897;
assign v_54903 = v_54753 & v_54902;
assign v_54905 = v_54808 & v_54904;
assign v_54906 = v_54752 & v_54902;
assign v_54908 = v_54750 & v_54907;
assign v_54910 = v_54814 & v_54909;
assign v_54911 = v_54749 & v_54907;
assign v_54913 = v_54747 & v_54912;
assign v_54915 = v_54820 & v_54914;
assign v_54916 = v_54746 & v_54912;
assign v_54918 = v_54744 & v_54917;
assign v_54920 = v_54826 & v_54919;
assign v_54921 = v_54743 & v_54917;
assign v_54923 = v_54741 & v_54922;
assign v_54925 = v_54832 & v_54924;
assign v_54926 = v_54740 & v_54922;
assign v_54928 = v_54738 & v_54927;
assign v_54930 = v_54838 & v_54929;
assign v_54931 = v_54737 & v_54927;
assign v_54933 = v_54735 & v_54932;
assign v_54935 = v_54844 & v_54934;
assign v_54936 = v_54734 & v_54932;
assign v_54938 = v_54732 & v_54937;
assign v_54940 = v_54850 & v_54939;
assign v_54941 = v_54731 & v_54937;
assign v_54943 = v_54729 & v_54942;
assign v_54945 = v_54856 & v_54944;
assign v_54946 = v_54728 & v_54942;
assign v_54948 = v_54726 & v_54947;
assign v_54950 = v_54862 & v_54949;
assign v_54951 = v_54725 & v_54947;
assign v_54953 = v_54723 & v_54952;
assign v_54955 = v_54868 & v_54954;
assign v_54956 = v_54722 & v_54952;
assign v_54958 = v_54957;
assign v_54960 = v_54872 & v_54959;
assign v_54961 = v_54960;
assign v_54963 = v_54962;
assign v_54965 = ~v_803;
assign v_54966 = ~v_54220;
assign v_54967 = v_54220;
assign v_54968 = ~v_807;
assign v_54969 = ~v_54224;
assign v_54970 = v_54224;
assign v_54971 = ~v_811;
assign v_54972 = ~v_54228;
assign v_54973 = v_54228;
assign v_54974 = ~v_815;
assign v_54975 = ~v_54232;
assign v_54976 = v_54232;
assign v_54977 = ~v_54235;
assign v_54978 = ~v_820;
assign v_54979 = v_820;
assign v_54980 = ~v_54239;
assign v_54981 = ~v_824;
assign v_54982 = v_824;
assign v_54983 = ~v_54243;
assign v_54984 = ~v_828;
assign v_54985 = v_828;
assign v_54986 = ~v_54247;
assign v_54987 = ~v_832;
assign v_54988 = v_832;
assign v_54989 = ~v_54251;
assign v_54990 = ~v_836;
assign v_54991 = v_836;
assign v_54992 = ~v_54255;
assign v_54993 = ~v_840;
assign v_54994 = v_840;
assign v_54995 = ~v_54259;
assign v_54996 = ~v_844;
assign v_54997 = v_844;
assign v_54998 = ~v_54263;
assign v_54999 = ~v_848;
assign v_55000 = v_848;
assign v_55001 = ~v_54267;
assign v_55002 = ~v_852;
assign v_55003 = v_852;
assign v_55004 = ~v_54271;
assign v_55005 = ~v_856;
assign v_55006 = v_856;
assign v_55007 = ~v_54275;
assign v_55008 = ~v_860;
assign v_55009 = v_860;
assign v_55010 = ~v_54279;
assign v_55011 = ~v_864;
assign v_55012 = v_864;
assign v_55013 = ~v_54283;
assign v_55014 = ~v_868;
assign v_55015 = v_55014;
assign v_55017 = v_55016;
assign v_55019 = v_55011 & v_55018;
assign v_55021 = v_54279;
assign v_55023 = v_55020 & v_55022;
assign v_55025 = v_55008 & v_55024;
assign v_55027 = v_54275;
assign v_55029 = v_55026 & v_55028;
assign v_55031 = v_55005 & v_55030;
assign v_55033 = v_54271;
assign v_55035 = v_55032 & v_55034;
assign v_55037 = v_55002 & v_55036;
assign v_55039 = v_54267;
assign v_55041 = v_55038 & v_55040;
assign v_55043 = v_54999 & v_55042;
assign v_55045 = v_54263;
assign v_55047 = v_55044 & v_55046;
assign v_55049 = v_54996 & v_55048;
assign v_55051 = v_54259;
assign v_55053 = v_55050 & v_55052;
assign v_55055 = v_54993 & v_55054;
assign v_55057 = v_54255;
assign v_55059 = v_55056 & v_55058;
assign v_55061 = v_54990 & v_55060;
assign v_55063 = v_54251;
assign v_55065 = v_55062 & v_55064;
assign v_55067 = v_54987 & v_55066;
assign v_55069 = v_54247;
assign v_55071 = v_55068 & v_55070;
assign v_55073 = v_54984 & v_55072;
assign v_55075 = v_54243;
assign v_55077 = v_55074 & v_55076;
assign v_55079 = v_54981 & v_55078;
assign v_55081 = v_54239;
assign v_55083 = v_55080 & v_55082;
assign v_55085 = v_54978 & v_55084;
assign v_55087 = v_54235;
assign v_55089 = v_55086 & v_55088;
assign v_55091 = v_54975 & v_55090;
assign v_55093 = v_815;
assign v_55095 = v_55092 & v_55094;
assign v_55097 = v_54972 & v_55096;
assign v_55099 = v_811;
assign v_55101 = v_55098 & v_55100;
assign v_55103 = v_54969 & v_55102;
assign v_55105 = v_807;
assign v_55107 = v_55104 & v_55106;
assign v_55109 = v_54966 & v_55108;
assign v_55111 = v_803;
assign v_55113 = v_55110 & v_55112;
assign v_55114 = v_55113;
assign v_55116 = v_54283;
assign v_55117 = v_868;
assign v_55118 = v_55117;
assign v_55119 = v_55116 & v_55118;
assign v_55120 = v_55119;
assign v_55121 = v_55011 & v_55120;
assign v_55123 = v_55021 & v_55122;
assign v_55124 = v_55010 & v_55120;
assign v_55126 = v_55008 & v_55125;
assign v_55128 = v_55027 & v_55127;
assign v_55129 = v_55007 & v_55125;
assign v_55131 = v_55005 & v_55130;
assign v_55133 = v_55033 & v_55132;
assign v_55134 = v_55004 & v_55130;
assign v_55136 = v_55002 & v_55135;
assign v_55138 = v_55039 & v_55137;
assign v_55139 = v_55001 & v_55135;
assign v_55141 = v_54999 & v_55140;
assign v_55143 = v_55045 & v_55142;
assign v_55144 = v_54998 & v_55140;
assign v_55146 = v_54996 & v_55145;
assign v_55148 = v_55051 & v_55147;
assign v_55149 = v_54995 & v_55145;
assign v_55151 = v_54993 & v_55150;
assign v_55153 = v_55057 & v_55152;
assign v_55154 = v_54992 & v_55150;
assign v_55156 = v_54990 & v_55155;
assign v_55158 = v_55063 & v_55157;
assign v_55159 = v_54989 & v_55155;
assign v_55161 = v_54987 & v_55160;
assign v_55163 = v_55069 & v_55162;
assign v_55164 = v_54986 & v_55160;
assign v_55166 = v_54984 & v_55165;
assign v_55168 = v_55075 & v_55167;
assign v_55169 = v_54983 & v_55165;
assign v_55171 = v_54981 & v_55170;
assign v_55173 = v_55081 & v_55172;
assign v_55174 = v_54980 & v_55170;
assign v_55176 = v_54978 & v_55175;
assign v_55178 = v_55087 & v_55177;
assign v_55179 = v_54977 & v_55175;
assign v_55181 = v_54975 & v_55180;
assign v_55183 = v_55093 & v_55182;
assign v_55184 = v_54974 & v_55180;
assign v_55186 = v_54972 & v_55185;
assign v_55188 = v_55099 & v_55187;
assign v_55189 = v_54971 & v_55185;
assign v_55191 = v_54969 & v_55190;
assign v_55193 = v_55105 & v_55192;
assign v_55194 = v_54968 & v_55190;
assign v_55196 = v_54966 & v_55195;
assign v_55198 = v_55111 & v_55197;
assign v_55199 = v_54965 & v_55195;
assign v_55201 = v_55200;
assign v_55203 = v_55115 & v_55202;
assign v_55204 = v_55203;
assign v_55206 = v_55205;
assign v_55208 = ~v_1063;
assign v_55209 = ~v_54220;
assign v_55210 = v_54220;
assign v_55211 = ~v_1067;
assign v_55212 = ~v_54224;
assign v_55213 = v_54224;
assign v_55214 = ~v_1071;
assign v_55215 = ~v_54228;
assign v_55216 = v_54228;
assign v_55217 = ~v_1075;
assign v_55218 = ~v_54232;
assign v_55219 = v_54232;
assign v_55220 = ~v_54235;
assign v_55221 = ~v_1080;
assign v_55222 = v_1080;
assign v_55223 = ~v_54239;
assign v_55224 = ~v_1084;
assign v_55225 = v_1084;
assign v_55226 = ~v_54243;
assign v_55227 = ~v_1088;
assign v_55228 = v_1088;
assign v_55229 = ~v_54247;
assign v_55230 = ~v_1092;
assign v_55231 = v_1092;
assign v_55232 = ~v_54251;
assign v_55233 = ~v_1096;
assign v_55234 = v_1096;
assign v_55235 = ~v_54255;
assign v_55236 = ~v_1100;
assign v_55237 = v_1100;
assign v_55238 = ~v_54259;
assign v_55239 = ~v_1104;
assign v_55240 = v_1104;
assign v_55241 = ~v_54263;
assign v_55242 = ~v_1108;
assign v_55243 = v_1108;
assign v_55244 = ~v_54267;
assign v_55245 = ~v_1112;
assign v_55246 = v_1112;
assign v_55247 = ~v_54271;
assign v_55248 = ~v_1116;
assign v_55249 = v_1116;
assign v_55250 = ~v_54275;
assign v_55251 = ~v_1120;
assign v_55252 = v_1120;
assign v_55253 = ~v_54279;
assign v_55254 = ~v_1124;
assign v_55255 = v_1124;
assign v_55256 = ~v_54283;
assign v_55257 = ~v_1128;
assign v_55258 = v_55257;
assign v_55260 = v_55259;
assign v_55262 = v_55254 & v_55261;
assign v_55264 = v_54279;
assign v_55266 = v_55263 & v_55265;
assign v_55268 = v_55251 & v_55267;
assign v_55270 = v_54275;
assign v_55272 = v_55269 & v_55271;
assign v_55274 = v_55248 & v_55273;
assign v_55276 = v_54271;
assign v_55278 = v_55275 & v_55277;
assign v_55280 = v_55245 & v_55279;
assign v_55282 = v_54267;
assign v_55284 = v_55281 & v_55283;
assign v_55286 = v_55242 & v_55285;
assign v_55288 = v_54263;
assign v_55290 = v_55287 & v_55289;
assign v_55292 = v_55239 & v_55291;
assign v_55294 = v_54259;
assign v_55296 = v_55293 & v_55295;
assign v_55298 = v_55236 & v_55297;
assign v_55300 = v_54255;
assign v_55302 = v_55299 & v_55301;
assign v_55304 = v_55233 & v_55303;
assign v_55306 = v_54251;
assign v_55308 = v_55305 & v_55307;
assign v_55310 = v_55230 & v_55309;
assign v_55312 = v_54247;
assign v_55314 = v_55311 & v_55313;
assign v_55316 = v_55227 & v_55315;
assign v_55318 = v_54243;
assign v_55320 = v_55317 & v_55319;
assign v_55322 = v_55224 & v_55321;
assign v_55324 = v_54239;
assign v_55326 = v_55323 & v_55325;
assign v_55328 = v_55221 & v_55327;
assign v_55330 = v_54235;
assign v_55332 = v_55329 & v_55331;
assign v_55334 = v_55218 & v_55333;
assign v_55336 = v_1075;
assign v_55338 = v_55335 & v_55337;
assign v_55340 = v_55215 & v_55339;
assign v_55342 = v_1071;
assign v_55344 = v_55341 & v_55343;
assign v_55346 = v_55212 & v_55345;
assign v_55348 = v_1067;
assign v_55350 = v_55347 & v_55349;
assign v_55352 = v_55209 & v_55351;
assign v_55354 = v_1063;
assign v_55356 = v_55353 & v_55355;
assign v_55357 = v_55356;
assign v_55359 = v_54283;
assign v_55360 = v_1128;
assign v_55361 = v_55360;
assign v_55362 = v_55359 & v_55361;
assign v_55363 = v_55362;
assign v_55364 = v_55254 & v_55363;
assign v_55366 = v_55264 & v_55365;
assign v_55367 = v_55253 & v_55363;
assign v_55369 = v_55251 & v_55368;
assign v_55371 = v_55270 & v_55370;
assign v_55372 = v_55250 & v_55368;
assign v_55374 = v_55248 & v_55373;
assign v_55376 = v_55276 & v_55375;
assign v_55377 = v_55247 & v_55373;
assign v_55379 = v_55245 & v_55378;
assign v_55381 = v_55282 & v_55380;
assign v_55382 = v_55244 & v_55378;
assign v_55384 = v_55242 & v_55383;
assign v_55386 = v_55288 & v_55385;
assign v_55387 = v_55241 & v_55383;
assign v_55389 = v_55239 & v_55388;
assign v_55391 = v_55294 & v_55390;
assign v_55392 = v_55238 & v_55388;
assign v_55394 = v_55236 & v_55393;
assign v_55396 = v_55300 & v_55395;
assign v_55397 = v_55235 & v_55393;
assign v_55399 = v_55233 & v_55398;
assign v_55401 = v_55306 & v_55400;
assign v_55402 = v_55232 & v_55398;
assign v_55404 = v_55230 & v_55403;
assign v_55406 = v_55312 & v_55405;
assign v_55407 = v_55229 & v_55403;
assign v_55409 = v_55227 & v_55408;
assign v_55411 = v_55318 & v_55410;
assign v_55412 = v_55226 & v_55408;
assign v_55414 = v_55224 & v_55413;
assign v_55416 = v_55324 & v_55415;
assign v_55417 = v_55223 & v_55413;
assign v_55419 = v_55221 & v_55418;
assign v_55421 = v_55330 & v_55420;
assign v_55422 = v_55220 & v_55418;
assign v_55424 = v_55218 & v_55423;
assign v_55426 = v_55336 & v_55425;
assign v_55427 = v_55217 & v_55423;
assign v_55429 = v_55215 & v_55428;
assign v_55431 = v_55342 & v_55430;
assign v_55432 = v_55214 & v_55428;
assign v_55434 = v_55212 & v_55433;
assign v_55436 = v_55348 & v_55435;
assign v_55437 = v_55211 & v_55433;
assign v_55439 = v_55209 & v_55438;
assign v_55441 = v_55354 & v_55440;
assign v_55442 = v_55208 & v_55438;
assign v_55444 = v_55443;
assign v_55446 = v_55358 & v_55445;
assign v_55447 = v_55446;
assign v_55449 = v_55448;
assign v_55451 = ~v_1323;
assign v_55452 = ~v_54220;
assign v_55453 = v_54220;
assign v_55454 = ~v_1327;
assign v_55455 = ~v_54224;
assign v_55456 = v_54224;
assign v_55457 = ~v_1331;
assign v_55458 = ~v_54228;
assign v_55459 = v_54228;
assign v_55460 = ~v_1335;
assign v_55461 = ~v_54232;
assign v_55462 = v_54232;
assign v_55463 = ~v_54235;
assign v_55464 = ~v_1340;
assign v_55465 = v_1340;
assign v_55466 = ~v_54239;
assign v_55467 = ~v_1344;
assign v_55468 = v_1344;
assign v_55469 = ~v_54243;
assign v_55470 = ~v_1348;
assign v_55471 = v_1348;
assign v_55472 = ~v_54247;
assign v_55473 = ~v_1352;
assign v_55474 = v_1352;
assign v_55475 = ~v_54251;
assign v_55476 = ~v_1356;
assign v_55477 = v_1356;
assign v_55478 = ~v_54255;
assign v_55479 = ~v_1360;
assign v_55480 = v_1360;
assign v_55481 = ~v_54259;
assign v_55482 = ~v_1364;
assign v_55483 = v_1364;
assign v_55484 = ~v_54263;
assign v_55485 = ~v_1368;
assign v_55486 = v_1368;
assign v_55487 = ~v_54267;
assign v_55488 = ~v_1372;
assign v_55489 = v_1372;
assign v_55490 = ~v_54271;
assign v_55491 = ~v_1376;
assign v_55492 = v_1376;
assign v_55493 = ~v_54275;
assign v_55494 = ~v_1380;
assign v_55495 = v_1380;
assign v_55496 = ~v_54279;
assign v_55497 = ~v_1384;
assign v_55498 = v_1384;
assign v_55499 = ~v_54283;
assign v_55500 = ~v_1388;
assign v_55501 = v_55500;
assign v_55503 = v_55502;
assign v_55505 = v_55497 & v_55504;
assign v_55507 = v_54279;
assign v_55509 = v_55506 & v_55508;
assign v_55511 = v_55494 & v_55510;
assign v_55513 = v_54275;
assign v_55515 = v_55512 & v_55514;
assign v_55517 = v_55491 & v_55516;
assign v_55519 = v_54271;
assign v_55521 = v_55518 & v_55520;
assign v_55523 = v_55488 & v_55522;
assign v_55525 = v_54267;
assign v_55527 = v_55524 & v_55526;
assign v_55529 = v_55485 & v_55528;
assign v_55531 = v_54263;
assign v_55533 = v_55530 & v_55532;
assign v_55535 = v_55482 & v_55534;
assign v_55537 = v_54259;
assign v_55539 = v_55536 & v_55538;
assign v_55541 = v_55479 & v_55540;
assign v_55543 = v_54255;
assign v_55545 = v_55542 & v_55544;
assign v_55547 = v_55476 & v_55546;
assign v_55549 = v_54251;
assign v_55551 = v_55548 & v_55550;
assign v_55553 = v_55473 & v_55552;
assign v_55555 = v_54247;
assign v_55557 = v_55554 & v_55556;
assign v_55559 = v_55470 & v_55558;
assign v_55561 = v_54243;
assign v_55563 = v_55560 & v_55562;
assign v_55565 = v_55467 & v_55564;
assign v_55567 = v_54239;
assign v_55569 = v_55566 & v_55568;
assign v_55571 = v_55464 & v_55570;
assign v_55573 = v_54235;
assign v_55575 = v_55572 & v_55574;
assign v_55577 = v_55461 & v_55576;
assign v_55579 = v_1335;
assign v_55581 = v_55578 & v_55580;
assign v_55583 = v_55458 & v_55582;
assign v_55585 = v_1331;
assign v_55587 = v_55584 & v_55586;
assign v_55589 = v_55455 & v_55588;
assign v_55591 = v_1327;
assign v_55593 = v_55590 & v_55592;
assign v_55595 = v_55452 & v_55594;
assign v_55597 = v_1323;
assign v_55599 = v_55596 & v_55598;
assign v_55600 = v_55599;
assign v_55602 = v_54283;
assign v_55603 = v_1388;
assign v_55604 = v_55603;
assign v_55605 = v_55602 & v_55604;
assign v_55606 = v_55605;
assign v_55607 = v_55497 & v_55606;
assign v_55609 = v_55507 & v_55608;
assign v_55610 = v_55496 & v_55606;
assign v_55612 = v_55494 & v_55611;
assign v_55614 = v_55513 & v_55613;
assign v_55615 = v_55493 & v_55611;
assign v_55617 = v_55491 & v_55616;
assign v_55619 = v_55519 & v_55618;
assign v_55620 = v_55490 & v_55616;
assign v_55622 = v_55488 & v_55621;
assign v_55624 = v_55525 & v_55623;
assign v_55625 = v_55487 & v_55621;
assign v_55627 = v_55485 & v_55626;
assign v_55629 = v_55531 & v_55628;
assign v_55630 = v_55484 & v_55626;
assign v_55632 = v_55482 & v_55631;
assign v_55634 = v_55537 & v_55633;
assign v_55635 = v_55481 & v_55631;
assign v_55637 = v_55479 & v_55636;
assign v_55639 = v_55543 & v_55638;
assign v_55640 = v_55478 & v_55636;
assign v_55642 = v_55476 & v_55641;
assign v_55644 = v_55549 & v_55643;
assign v_55645 = v_55475 & v_55641;
assign v_55647 = v_55473 & v_55646;
assign v_55649 = v_55555 & v_55648;
assign v_55650 = v_55472 & v_55646;
assign v_55652 = v_55470 & v_55651;
assign v_55654 = v_55561 & v_55653;
assign v_55655 = v_55469 & v_55651;
assign v_55657 = v_55467 & v_55656;
assign v_55659 = v_55567 & v_55658;
assign v_55660 = v_55466 & v_55656;
assign v_55662 = v_55464 & v_55661;
assign v_55664 = v_55573 & v_55663;
assign v_55665 = v_55463 & v_55661;
assign v_55667 = v_55461 & v_55666;
assign v_55669 = v_55579 & v_55668;
assign v_55670 = v_55460 & v_55666;
assign v_55672 = v_55458 & v_55671;
assign v_55674 = v_55585 & v_55673;
assign v_55675 = v_55457 & v_55671;
assign v_55677 = v_55455 & v_55676;
assign v_55679 = v_55591 & v_55678;
assign v_55680 = v_55454 & v_55676;
assign v_55682 = v_55452 & v_55681;
assign v_55684 = v_55597 & v_55683;
assign v_55685 = v_55451 & v_55681;
assign v_55687 = v_55686;
assign v_55689 = v_55601 & v_55688;
assign v_55690 = v_55689;
assign v_55692 = v_55691;
assign v_55694 = ~v_1583;
assign v_55695 = ~v_54220;
assign v_55696 = v_54220;
assign v_55697 = ~v_1587;
assign v_55698 = ~v_54224;
assign v_55699 = v_54224;
assign v_55700 = ~v_1591;
assign v_55701 = ~v_54228;
assign v_55702 = v_54228;
assign v_55703 = ~v_1595;
assign v_55704 = ~v_54232;
assign v_55705 = v_54232;
assign v_55706 = ~v_54235;
assign v_55707 = ~v_1600;
assign v_55708 = v_1600;
assign v_55709 = ~v_54239;
assign v_55710 = ~v_1604;
assign v_55711 = v_1604;
assign v_55712 = ~v_54243;
assign v_55713 = ~v_1608;
assign v_55714 = v_1608;
assign v_55715 = ~v_54247;
assign v_55716 = ~v_1612;
assign v_55717 = v_1612;
assign v_55718 = ~v_54251;
assign v_55719 = ~v_1616;
assign v_55720 = v_1616;
assign v_55721 = ~v_54255;
assign v_55722 = ~v_1620;
assign v_55723 = v_1620;
assign v_55724 = ~v_54259;
assign v_55725 = ~v_1624;
assign v_55726 = v_1624;
assign v_55727 = ~v_54263;
assign v_55728 = ~v_1628;
assign v_55729 = v_1628;
assign v_55730 = ~v_54267;
assign v_55731 = ~v_1632;
assign v_55732 = v_1632;
assign v_55733 = ~v_54271;
assign v_55734 = ~v_1636;
assign v_55735 = v_1636;
assign v_55736 = ~v_54275;
assign v_55737 = ~v_1640;
assign v_55738 = v_1640;
assign v_55739 = ~v_54279;
assign v_55740 = ~v_1644;
assign v_55741 = v_1644;
assign v_55742 = ~v_54283;
assign v_55743 = ~v_1648;
assign v_55744 = v_55743;
assign v_55746 = v_55745;
assign v_55748 = v_55740 & v_55747;
assign v_55750 = v_54279;
assign v_55752 = v_55749 & v_55751;
assign v_55754 = v_55737 & v_55753;
assign v_55756 = v_54275;
assign v_55758 = v_55755 & v_55757;
assign v_55760 = v_55734 & v_55759;
assign v_55762 = v_54271;
assign v_55764 = v_55761 & v_55763;
assign v_55766 = v_55731 & v_55765;
assign v_55768 = v_54267;
assign v_55770 = v_55767 & v_55769;
assign v_55772 = v_55728 & v_55771;
assign v_55774 = v_54263;
assign v_55776 = v_55773 & v_55775;
assign v_55778 = v_55725 & v_55777;
assign v_55780 = v_54259;
assign v_55782 = v_55779 & v_55781;
assign v_55784 = v_55722 & v_55783;
assign v_55786 = v_54255;
assign v_55788 = v_55785 & v_55787;
assign v_55790 = v_55719 & v_55789;
assign v_55792 = v_54251;
assign v_55794 = v_55791 & v_55793;
assign v_55796 = v_55716 & v_55795;
assign v_55798 = v_54247;
assign v_55800 = v_55797 & v_55799;
assign v_55802 = v_55713 & v_55801;
assign v_55804 = v_54243;
assign v_55806 = v_55803 & v_55805;
assign v_55808 = v_55710 & v_55807;
assign v_55810 = v_54239;
assign v_55812 = v_55809 & v_55811;
assign v_55814 = v_55707 & v_55813;
assign v_55816 = v_54235;
assign v_55818 = v_55815 & v_55817;
assign v_55820 = v_55704 & v_55819;
assign v_55822 = v_1595;
assign v_55824 = v_55821 & v_55823;
assign v_55826 = v_55701 & v_55825;
assign v_55828 = v_1591;
assign v_55830 = v_55827 & v_55829;
assign v_55832 = v_55698 & v_55831;
assign v_55834 = v_1587;
assign v_55836 = v_55833 & v_55835;
assign v_55838 = v_55695 & v_55837;
assign v_55840 = v_1583;
assign v_55842 = v_55839 & v_55841;
assign v_55843 = v_55842;
assign v_55845 = v_54283;
assign v_55846 = v_1648;
assign v_55847 = v_55846;
assign v_55848 = v_55845 & v_55847;
assign v_55849 = v_55848;
assign v_55850 = v_55740 & v_55849;
assign v_55852 = v_55750 & v_55851;
assign v_55853 = v_55739 & v_55849;
assign v_55855 = v_55737 & v_55854;
assign v_55857 = v_55756 & v_55856;
assign v_55858 = v_55736 & v_55854;
assign v_55860 = v_55734 & v_55859;
assign v_55862 = v_55762 & v_55861;
assign v_55863 = v_55733 & v_55859;
assign v_55865 = v_55731 & v_55864;
assign v_55867 = v_55768 & v_55866;
assign v_55868 = v_55730 & v_55864;
assign v_55870 = v_55728 & v_55869;
assign v_55872 = v_55774 & v_55871;
assign v_55873 = v_55727 & v_55869;
assign v_55875 = v_55725 & v_55874;
assign v_55877 = v_55780 & v_55876;
assign v_55878 = v_55724 & v_55874;
assign v_55880 = v_55722 & v_55879;
assign v_55882 = v_55786 & v_55881;
assign v_55883 = v_55721 & v_55879;
assign v_55885 = v_55719 & v_55884;
assign v_55887 = v_55792 & v_55886;
assign v_55888 = v_55718 & v_55884;
assign v_55890 = v_55716 & v_55889;
assign v_55892 = v_55798 & v_55891;
assign v_55893 = v_55715 & v_55889;
assign v_55895 = v_55713 & v_55894;
assign v_55897 = v_55804 & v_55896;
assign v_55898 = v_55712 & v_55894;
assign v_55900 = v_55710 & v_55899;
assign v_55902 = v_55810 & v_55901;
assign v_55903 = v_55709 & v_55899;
assign v_55905 = v_55707 & v_55904;
assign v_55907 = v_55816 & v_55906;
assign v_55908 = v_55706 & v_55904;
assign v_55910 = v_55704 & v_55909;
assign v_55912 = v_55822 & v_55911;
assign v_55913 = v_55703 & v_55909;
assign v_55915 = v_55701 & v_55914;
assign v_55917 = v_55828 & v_55916;
assign v_55918 = v_55700 & v_55914;
assign v_55920 = v_55698 & v_55919;
assign v_55922 = v_55834 & v_55921;
assign v_55923 = v_55697 & v_55919;
assign v_55925 = v_55695 & v_55924;
assign v_55927 = v_55840 & v_55926;
assign v_55928 = v_55694 & v_55924;
assign v_55930 = v_55929;
assign v_55932 = v_55844 & v_55931;
assign v_55933 = v_55932;
assign v_55935 = v_55934;
assign v_55937 = ~v_1843;
assign v_55938 = ~v_54220;
assign v_55939 = v_54220;
assign v_55940 = ~v_1847;
assign v_55941 = ~v_54224;
assign v_55942 = v_54224;
assign v_55943 = ~v_1851;
assign v_55944 = ~v_54228;
assign v_55945 = v_54228;
assign v_55946 = ~v_1855;
assign v_55947 = ~v_54232;
assign v_55948 = v_54232;
assign v_55949 = ~v_54235;
assign v_55950 = ~v_1860;
assign v_55951 = v_1860;
assign v_55952 = ~v_54239;
assign v_55953 = ~v_1864;
assign v_55954 = v_1864;
assign v_55955 = ~v_54243;
assign v_55956 = ~v_1868;
assign v_55957 = v_1868;
assign v_55958 = ~v_54247;
assign v_55959 = ~v_1872;
assign v_55960 = v_1872;
assign v_55961 = ~v_54251;
assign v_55962 = ~v_1876;
assign v_55963 = v_1876;
assign v_55964 = ~v_54255;
assign v_55965 = ~v_1880;
assign v_55966 = v_1880;
assign v_55967 = ~v_54259;
assign v_55968 = ~v_1884;
assign v_55969 = v_1884;
assign v_55970 = ~v_54263;
assign v_55971 = ~v_1888;
assign v_55972 = v_1888;
assign v_55973 = ~v_54267;
assign v_55974 = ~v_1892;
assign v_55975 = v_1892;
assign v_55976 = ~v_54271;
assign v_55977 = ~v_1896;
assign v_55978 = v_1896;
assign v_55979 = ~v_54275;
assign v_55980 = ~v_1900;
assign v_55981 = v_1900;
assign v_55982 = ~v_54279;
assign v_55983 = ~v_1904;
assign v_55984 = v_1904;
assign v_55985 = ~v_54283;
assign v_55986 = ~v_1908;
assign v_55987 = v_55986;
assign v_55989 = v_55988;
assign v_55991 = v_55983 & v_55990;
assign v_55993 = v_54279;
assign v_55995 = v_55992 & v_55994;
assign v_55997 = v_55980 & v_55996;
assign v_55999 = v_54275;
assign v_56001 = v_55998 & v_56000;
assign v_56003 = v_55977 & v_56002;
assign v_56005 = v_54271;
assign v_56007 = v_56004 & v_56006;
assign v_56009 = v_55974 & v_56008;
assign v_56011 = v_54267;
assign v_56013 = v_56010 & v_56012;
assign v_56015 = v_55971 & v_56014;
assign v_56017 = v_54263;
assign v_56019 = v_56016 & v_56018;
assign v_56021 = v_55968 & v_56020;
assign v_56023 = v_54259;
assign v_56025 = v_56022 & v_56024;
assign v_56027 = v_55965 & v_56026;
assign v_56029 = v_54255;
assign v_56031 = v_56028 & v_56030;
assign v_56033 = v_55962 & v_56032;
assign v_56035 = v_54251;
assign v_56037 = v_56034 & v_56036;
assign v_56039 = v_55959 & v_56038;
assign v_56041 = v_54247;
assign v_56043 = v_56040 & v_56042;
assign v_56045 = v_55956 & v_56044;
assign v_56047 = v_54243;
assign v_56049 = v_56046 & v_56048;
assign v_56051 = v_55953 & v_56050;
assign v_56053 = v_54239;
assign v_56055 = v_56052 & v_56054;
assign v_56057 = v_55950 & v_56056;
assign v_56059 = v_54235;
assign v_56061 = v_56058 & v_56060;
assign v_56063 = v_55947 & v_56062;
assign v_56065 = v_1855;
assign v_56067 = v_56064 & v_56066;
assign v_56069 = v_55944 & v_56068;
assign v_56071 = v_1851;
assign v_56073 = v_56070 & v_56072;
assign v_56075 = v_55941 & v_56074;
assign v_56077 = v_1847;
assign v_56079 = v_56076 & v_56078;
assign v_56081 = v_55938 & v_56080;
assign v_56083 = v_1843;
assign v_56085 = v_56082 & v_56084;
assign v_56086 = v_56085;
assign v_56088 = v_54283;
assign v_56089 = v_1908;
assign v_56090 = v_56089;
assign v_56091 = v_56088 & v_56090;
assign v_56092 = v_56091;
assign v_56093 = v_55983 & v_56092;
assign v_56095 = v_55993 & v_56094;
assign v_56096 = v_55982 & v_56092;
assign v_56098 = v_55980 & v_56097;
assign v_56100 = v_55999 & v_56099;
assign v_56101 = v_55979 & v_56097;
assign v_56103 = v_55977 & v_56102;
assign v_56105 = v_56005 & v_56104;
assign v_56106 = v_55976 & v_56102;
assign v_56108 = v_55974 & v_56107;
assign v_56110 = v_56011 & v_56109;
assign v_56111 = v_55973 & v_56107;
assign v_56113 = v_55971 & v_56112;
assign v_56115 = v_56017 & v_56114;
assign v_56116 = v_55970 & v_56112;
assign v_56118 = v_55968 & v_56117;
assign v_56120 = v_56023 & v_56119;
assign v_56121 = v_55967 & v_56117;
assign v_56123 = v_55965 & v_56122;
assign v_56125 = v_56029 & v_56124;
assign v_56126 = v_55964 & v_56122;
assign v_56128 = v_55962 & v_56127;
assign v_56130 = v_56035 & v_56129;
assign v_56131 = v_55961 & v_56127;
assign v_56133 = v_55959 & v_56132;
assign v_56135 = v_56041 & v_56134;
assign v_56136 = v_55958 & v_56132;
assign v_56138 = v_55956 & v_56137;
assign v_56140 = v_56047 & v_56139;
assign v_56141 = v_55955 & v_56137;
assign v_56143 = v_55953 & v_56142;
assign v_56145 = v_56053 & v_56144;
assign v_56146 = v_55952 & v_56142;
assign v_56148 = v_55950 & v_56147;
assign v_56150 = v_56059 & v_56149;
assign v_56151 = v_55949 & v_56147;
assign v_56153 = v_55947 & v_56152;
assign v_56155 = v_56065 & v_56154;
assign v_56156 = v_55946 & v_56152;
assign v_56158 = v_55944 & v_56157;
assign v_56160 = v_56071 & v_56159;
assign v_56161 = v_55943 & v_56157;
assign v_56163 = v_55941 & v_56162;
assign v_56165 = v_56077 & v_56164;
assign v_56166 = v_55940 & v_56162;
assign v_56168 = v_55938 & v_56167;
assign v_56170 = v_56083 & v_56169;
assign v_56171 = v_55937 & v_56167;
assign v_56173 = v_56172;
assign v_56175 = v_56087 & v_56174;
assign v_56176 = v_56175;
assign v_56178 = v_56177;
assign v_56180 = ~v_2103;
assign v_56181 = ~v_54220;
assign v_56182 = v_54220;
assign v_56183 = ~v_2107;
assign v_56184 = ~v_54224;
assign v_56185 = v_54224;
assign v_56186 = ~v_2111;
assign v_56187 = ~v_54228;
assign v_56188 = v_54228;
assign v_56189 = ~v_2115;
assign v_56190 = ~v_54232;
assign v_56191 = v_54232;
assign v_56192 = ~v_54235;
assign v_56193 = ~v_2120;
assign v_56194 = v_2120;
assign v_56195 = ~v_54239;
assign v_56196 = ~v_2124;
assign v_56197 = v_2124;
assign v_56198 = ~v_54243;
assign v_56199 = ~v_2128;
assign v_56200 = v_2128;
assign v_56201 = ~v_54247;
assign v_56202 = ~v_2132;
assign v_56203 = v_2132;
assign v_56204 = ~v_54251;
assign v_56205 = ~v_2136;
assign v_56206 = v_2136;
assign v_56207 = ~v_54255;
assign v_56208 = ~v_2140;
assign v_56209 = v_2140;
assign v_56210 = ~v_54259;
assign v_56211 = ~v_2144;
assign v_56212 = v_2144;
assign v_56213 = ~v_54263;
assign v_56214 = ~v_2148;
assign v_56215 = v_2148;
assign v_56216 = ~v_54267;
assign v_56217 = ~v_2152;
assign v_56218 = v_2152;
assign v_56219 = ~v_54271;
assign v_56220 = ~v_2156;
assign v_56221 = v_2156;
assign v_56222 = ~v_54275;
assign v_56223 = ~v_2160;
assign v_56224 = v_2160;
assign v_56225 = ~v_54279;
assign v_56226 = ~v_2164;
assign v_56227 = v_2164;
assign v_56228 = ~v_54283;
assign v_56229 = ~v_2168;
assign v_56230 = v_56229;
assign v_56232 = v_56231;
assign v_56234 = v_56226 & v_56233;
assign v_56236 = v_54279;
assign v_56238 = v_56235 & v_56237;
assign v_56240 = v_56223 & v_56239;
assign v_56242 = v_54275;
assign v_56244 = v_56241 & v_56243;
assign v_56246 = v_56220 & v_56245;
assign v_56248 = v_54271;
assign v_56250 = v_56247 & v_56249;
assign v_56252 = v_56217 & v_56251;
assign v_56254 = v_54267;
assign v_56256 = v_56253 & v_56255;
assign v_56258 = v_56214 & v_56257;
assign v_56260 = v_54263;
assign v_56262 = v_56259 & v_56261;
assign v_56264 = v_56211 & v_56263;
assign v_56266 = v_54259;
assign v_56268 = v_56265 & v_56267;
assign v_56270 = v_56208 & v_56269;
assign v_56272 = v_54255;
assign v_56274 = v_56271 & v_56273;
assign v_56276 = v_56205 & v_56275;
assign v_56278 = v_54251;
assign v_56280 = v_56277 & v_56279;
assign v_56282 = v_56202 & v_56281;
assign v_56284 = v_54247;
assign v_56286 = v_56283 & v_56285;
assign v_56288 = v_56199 & v_56287;
assign v_56290 = v_54243;
assign v_56292 = v_56289 & v_56291;
assign v_56294 = v_56196 & v_56293;
assign v_56296 = v_54239;
assign v_56298 = v_56295 & v_56297;
assign v_56300 = v_56193 & v_56299;
assign v_56302 = v_54235;
assign v_56304 = v_56301 & v_56303;
assign v_56306 = v_56190 & v_56305;
assign v_56308 = v_2115;
assign v_56310 = v_56307 & v_56309;
assign v_56312 = v_56187 & v_56311;
assign v_56314 = v_2111;
assign v_56316 = v_56313 & v_56315;
assign v_56318 = v_56184 & v_56317;
assign v_56320 = v_2107;
assign v_56322 = v_56319 & v_56321;
assign v_56324 = v_56181 & v_56323;
assign v_56326 = v_2103;
assign v_56328 = v_56325 & v_56327;
assign v_56329 = v_56328;
assign v_56331 = v_54283;
assign v_56332 = v_2168;
assign v_56333 = v_56332;
assign v_56334 = v_56331 & v_56333;
assign v_56335 = v_56334;
assign v_56336 = v_56226 & v_56335;
assign v_56338 = v_56236 & v_56337;
assign v_56339 = v_56225 & v_56335;
assign v_56341 = v_56223 & v_56340;
assign v_56343 = v_56242 & v_56342;
assign v_56344 = v_56222 & v_56340;
assign v_56346 = v_56220 & v_56345;
assign v_56348 = v_56248 & v_56347;
assign v_56349 = v_56219 & v_56345;
assign v_56351 = v_56217 & v_56350;
assign v_56353 = v_56254 & v_56352;
assign v_56354 = v_56216 & v_56350;
assign v_56356 = v_56214 & v_56355;
assign v_56358 = v_56260 & v_56357;
assign v_56359 = v_56213 & v_56355;
assign v_56361 = v_56211 & v_56360;
assign v_56363 = v_56266 & v_56362;
assign v_56364 = v_56210 & v_56360;
assign v_56366 = v_56208 & v_56365;
assign v_56368 = v_56272 & v_56367;
assign v_56369 = v_56207 & v_56365;
assign v_56371 = v_56205 & v_56370;
assign v_56373 = v_56278 & v_56372;
assign v_56374 = v_56204 & v_56370;
assign v_56376 = v_56202 & v_56375;
assign v_56378 = v_56284 & v_56377;
assign v_56379 = v_56201 & v_56375;
assign v_56381 = v_56199 & v_56380;
assign v_56383 = v_56290 & v_56382;
assign v_56384 = v_56198 & v_56380;
assign v_56386 = v_56196 & v_56385;
assign v_56388 = v_56296 & v_56387;
assign v_56389 = v_56195 & v_56385;
assign v_56391 = v_56193 & v_56390;
assign v_56393 = v_56302 & v_56392;
assign v_56394 = v_56192 & v_56390;
assign v_56396 = v_56190 & v_56395;
assign v_56398 = v_56308 & v_56397;
assign v_56399 = v_56189 & v_56395;
assign v_56401 = v_56187 & v_56400;
assign v_56403 = v_56314 & v_56402;
assign v_56404 = v_56186 & v_56400;
assign v_56406 = v_56184 & v_56405;
assign v_56408 = v_56320 & v_56407;
assign v_56409 = v_56183 & v_56405;
assign v_56411 = v_56181 & v_56410;
assign v_56413 = v_56326 & v_56412;
assign v_56414 = v_56180 & v_56410;
assign v_56416 = v_56415;
assign v_56418 = v_56330 & v_56417;
assign v_56419 = v_56418;
assign v_56421 = v_56420;
assign v_56423 = ~v_2363;
assign v_56424 = ~v_54220;
assign v_56425 = v_54220;
assign v_56426 = ~v_2367;
assign v_56427 = ~v_54224;
assign v_56428 = v_54224;
assign v_56429 = ~v_2371;
assign v_56430 = ~v_54228;
assign v_56431 = v_54228;
assign v_56432 = ~v_2375;
assign v_56433 = ~v_54232;
assign v_56434 = v_54232;
assign v_56435 = ~v_54235;
assign v_56436 = ~v_2380;
assign v_56437 = v_2380;
assign v_56438 = ~v_54239;
assign v_56439 = ~v_2384;
assign v_56440 = v_2384;
assign v_56441 = ~v_54243;
assign v_56442 = ~v_2388;
assign v_56443 = v_2388;
assign v_56444 = ~v_54247;
assign v_56445 = ~v_2392;
assign v_56446 = v_2392;
assign v_56447 = ~v_54251;
assign v_56448 = ~v_2396;
assign v_56449 = v_2396;
assign v_56450 = ~v_54255;
assign v_56451 = ~v_2400;
assign v_56452 = v_2400;
assign v_56453 = ~v_54259;
assign v_56454 = ~v_2404;
assign v_56455 = v_2404;
assign v_56456 = ~v_54263;
assign v_56457 = ~v_2408;
assign v_56458 = v_2408;
assign v_56459 = ~v_54267;
assign v_56460 = ~v_2412;
assign v_56461 = v_2412;
assign v_56462 = ~v_54271;
assign v_56463 = ~v_2416;
assign v_56464 = v_2416;
assign v_56465 = ~v_54275;
assign v_56466 = ~v_2420;
assign v_56467 = v_2420;
assign v_56468 = ~v_54279;
assign v_56469 = ~v_2424;
assign v_56470 = v_2424;
assign v_56471 = ~v_54283;
assign v_56472 = ~v_2428;
assign v_56473 = v_56472;
assign v_56475 = v_56474;
assign v_56477 = v_56469 & v_56476;
assign v_56479 = v_54279;
assign v_56481 = v_56478 & v_56480;
assign v_56483 = v_56466 & v_56482;
assign v_56485 = v_54275;
assign v_56487 = v_56484 & v_56486;
assign v_56489 = v_56463 & v_56488;
assign v_56491 = v_54271;
assign v_56493 = v_56490 & v_56492;
assign v_56495 = v_56460 & v_56494;
assign v_56497 = v_54267;
assign v_56499 = v_56496 & v_56498;
assign v_56501 = v_56457 & v_56500;
assign v_56503 = v_54263;
assign v_56505 = v_56502 & v_56504;
assign v_56507 = v_56454 & v_56506;
assign v_56509 = v_54259;
assign v_56511 = v_56508 & v_56510;
assign v_56513 = v_56451 & v_56512;
assign v_56515 = v_54255;
assign v_56517 = v_56514 & v_56516;
assign v_56519 = v_56448 & v_56518;
assign v_56521 = v_54251;
assign v_56523 = v_56520 & v_56522;
assign v_56525 = v_56445 & v_56524;
assign v_56527 = v_54247;
assign v_56529 = v_56526 & v_56528;
assign v_56531 = v_56442 & v_56530;
assign v_56533 = v_54243;
assign v_56535 = v_56532 & v_56534;
assign v_56537 = v_56439 & v_56536;
assign v_56539 = v_54239;
assign v_56541 = v_56538 & v_56540;
assign v_56543 = v_56436 & v_56542;
assign v_56545 = v_54235;
assign v_56547 = v_56544 & v_56546;
assign v_56549 = v_56433 & v_56548;
assign v_56551 = v_2375;
assign v_56553 = v_56550 & v_56552;
assign v_56555 = v_56430 & v_56554;
assign v_56557 = v_2371;
assign v_56559 = v_56556 & v_56558;
assign v_56561 = v_56427 & v_56560;
assign v_56563 = v_2367;
assign v_56565 = v_56562 & v_56564;
assign v_56567 = v_56424 & v_56566;
assign v_56569 = v_2363;
assign v_56571 = v_56568 & v_56570;
assign v_56572 = v_56571;
assign v_56574 = v_54283;
assign v_56575 = v_2428;
assign v_56576 = v_56575;
assign v_56577 = v_56574 & v_56576;
assign v_56578 = v_56577;
assign v_56579 = v_56469 & v_56578;
assign v_56581 = v_56479 & v_56580;
assign v_56582 = v_56468 & v_56578;
assign v_56584 = v_56466 & v_56583;
assign v_56586 = v_56485 & v_56585;
assign v_56587 = v_56465 & v_56583;
assign v_56589 = v_56463 & v_56588;
assign v_56591 = v_56491 & v_56590;
assign v_56592 = v_56462 & v_56588;
assign v_56594 = v_56460 & v_56593;
assign v_56596 = v_56497 & v_56595;
assign v_56597 = v_56459 & v_56593;
assign v_56599 = v_56457 & v_56598;
assign v_56601 = v_56503 & v_56600;
assign v_56602 = v_56456 & v_56598;
assign v_56604 = v_56454 & v_56603;
assign v_56606 = v_56509 & v_56605;
assign v_56607 = v_56453 & v_56603;
assign v_56609 = v_56451 & v_56608;
assign v_56611 = v_56515 & v_56610;
assign v_56612 = v_56450 & v_56608;
assign v_56614 = v_56448 & v_56613;
assign v_56616 = v_56521 & v_56615;
assign v_56617 = v_56447 & v_56613;
assign v_56619 = v_56445 & v_56618;
assign v_56621 = v_56527 & v_56620;
assign v_56622 = v_56444 & v_56618;
assign v_56624 = v_56442 & v_56623;
assign v_56626 = v_56533 & v_56625;
assign v_56627 = v_56441 & v_56623;
assign v_56629 = v_56439 & v_56628;
assign v_56631 = v_56539 & v_56630;
assign v_56632 = v_56438 & v_56628;
assign v_56634 = v_56436 & v_56633;
assign v_56636 = v_56545 & v_56635;
assign v_56637 = v_56435 & v_56633;
assign v_56639 = v_56433 & v_56638;
assign v_56641 = v_56551 & v_56640;
assign v_56642 = v_56432 & v_56638;
assign v_56644 = v_56430 & v_56643;
assign v_56646 = v_56557 & v_56645;
assign v_56647 = v_56429 & v_56643;
assign v_56649 = v_56427 & v_56648;
assign v_56651 = v_56563 & v_56650;
assign v_56652 = v_56426 & v_56648;
assign v_56654 = v_56424 & v_56653;
assign v_56656 = v_56569 & v_56655;
assign v_56657 = v_56423 & v_56653;
assign v_56659 = v_56658;
assign v_56661 = v_56573 & v_56660;
assign v_56662 = v_56661;
assign v_56664 = v_56663;
assign v_56666 = ~v_2623;
assign v_56667 = ~v_54220;
assign v_56668 = v_54220;
assign v_56669 = ~v_2627;
assign v_56670 = ~v_54224;
assign v_56671 = v_54224;
assign v_56672 = ~v_2631;
assign v_56673 = ~v_54228;
assign v_56674 = v_54228;
assign v_56675 = ~v_2635;
assign v_56676 = ~v_54232;
assign v_56677 = v_54232;
assign v_56678 = ~v_54235;
assign v_56679 = ~v_2640;
assign v_56680 = v_2640;
assign v_56681 = ~v_54239;
assign v_56682 = ~v_2644;
assign v_56683 = v_2644;
assign v_56684 = ~v_54243;
assign v_56685 = ~v_2648;
assign v_56686 = v_2648;
assign v_56687 = ~v_54247;
assign v_56688 = ~v_2652;
assign v_56689 = v_2652;
assign v_56690 = ~v_54251;
assign v_56691 = ~v_2656;
assign v_56692 = v_2656;
assign v_56693 = ~v_54255;
assign v_56694 = ~v_2660;
assign v_56695 = v_2660;
assign v_56696 = ~v_54259;
assign v_56697 = ~v_2664;
assign v_56698 = v_2664;
assign v_56699 = ~v_54263;
assign v_56700 = ~v_2668;
assign v_56701 = v_2668;
assign v_56702 = ~v_54267;
assign v_56703 = ~v_2672;
assign v_56704 = v_2672;
assign v_56705 = ~v_54271;
assign v_56706 = ~v_2676;
assign v_56707 = v_2676;
assign v_56708 = ~v_54275;
assign v_56709 = ~v_2680;
assign v_56710 = v_2680;
assign v_56711 = ~v_54279;
assign v_56712 = ~v_2684;
assign v_56713 = v_2684;
assign v_56714 = ~v_54283;
assign v_56715 = ~v_2688;
assign v_56716 = v_56715;
assign v_56718 = v_56717;
assign v_56720 = v_56712 & v_56719;
assign v_56722 = v_54279;
assign v_56724 = v_56721 & v_56723;
assign v_56726 = v_56709 & v_56725;
assign v_56728 = v_54275;
assign v_56730 = v_56727 & v_56729;
assign v_56732 = v_56706 & v_56731;
assign v_56734 = v_54271;
assign v_56736 = v_56733 & v_56735;
assign v_56738 = v_56703 & v_56737;
assign v_56740 = v_54267;
assign v_56742 = v_56739 & v_56741;
assign v_56744 = v_56700 & v_56743;
assign v_56746 = v_54263;
assign v_56748 = v_56745 & v_56747;
assign v_56750 = v_56697 & v_56749;
assign v_56752 = v_54259;
assign v_56754 = v_56751 & v_56753;
assign v_56756 = v_56694 & v_56755;
assign v_56758 = v_54255;
assign v_56760 = v_56757 & v_56759;
assign v_56762 = v_56691 & v_56761;
assign v_56764 = v_54251;
assign v_56766 = v_56763 & v_56765;
assign v_56768 = v_56688 & v_56767;
assign v_56770 = v_54247;
assign v_56772 = v_56769 & v_56771;
assign v_56774 = v_56685 & v_56773;
assign v_56776 = v_54243;
assign v_56778 = v_56775 & v_56777;
assign v_56780 = v_56682 & v_56779;
assign v_56782 = v_54239;
assign v_56784 = v_56781 & v_56783;
assign v_56786 = v_56679 & v_56785;
assign v_56788 = v_54235;
assign v_56790 = v_56787 & v_56789;
assign v_56792 = v_56676 & v_56791;
assign v_56794 = v_2635;
assign v_56796 = v_56793 & v_56795;
assign v_56798 = v_56673 & v_56797;
assign v_56800 = v_2631;
assign v_56802 = v_56799 & v_56801;
assign v_56804 = v_56670 & v_56803;
assign v_56806 = v_2627;
assign v_56808 = v_56805 & v_56807;
assign v_56810 = v_56667 & v_56809;
assign v_56812 = v_2623;
assign v_56814 = v_56811 & v_56813;
assign v_56815 = v_56814;
assign v_56817 = v_54283;
assign v_56818 = v_2688;
assign v_56819 = v_56818;
assign v_56820 = v_56817 & v_56819;
assign v_56821 = v_56820;
assign v_56822 = v_56712 & v_56821;
assign v_56824 = v_56722 & v_56823;
assign v_56825 = v_56711 & v_56821;
assign v_56827 = v_56709 & v_56826;
assign v_56829 = v_56728 & v_56828;
assign v_56830 = v_56708 & v_56826;
assign v_56832 = v_56706 & v_56831;
assign v_56834 = v_56734 & v_56833;
assign v_56835 = v_56705 & v_56831;
assign v_56837 = v_56703 & v_56836;
assign v_56839 = v_56740 & v_56838;
assign v_56840 = v_56702 & v_56836;
assign v_56842 = v_56700 & v_56841;
assign v_56844 = v_56746 & v_56843;
assign v_56845 = v_56699 & v_56841;
assign v_56847 = v_56697 & v_56846;
assign v_56849 = v_56752 & v_56848;
assign v_56850 = v_56696 & v_56846;
assign v_56852 = v_56694 & v_56851;
assign v_56854 = v_56758 & v_56853;
assign v_56855 = v_56693 & v_56851;
assign v_56857 = v_56691 & v_56856;
assign v_56859 = v_56764 & v_56858;
assign v_56860 = v_56690 & v_56856;
assign v_56862 = v_56688 & v_56861;
assign v_56864 = v_56770 & v_56863;
assign v_56865 = v_56687 & v_56861;
assign v_56867 = v_56685 & v_56866;
assign v_56869 = v_56776 & v_56868;
assign v_56870 = v_56684 & v_56866;
assign v_56872 = v_56682 & v_56871;
assign v_56874 = v_56782 & v_56873;
assign v_56875 = v_56681 & v_56871;
assign v_56877 = v_56679 & v_56876;
assign v_56879 = v_56788 & v_56878;
assign v_56880 = v_56678 & v_56876;
assign v_56882 = v_56676 & v_56881;
assign v_56884 = v_56794 & v_56883;
assign v_56885 = v_56675 & v_56881;
assign v_56887 = v_56673 & v_56886;
assign v_56889 = v_56800 & v_56888;
assign v_56890 = v_56672 & v_56886;
assign v_56892 = v_56670 & v_56891;
assign v_56894 = v_56806 & v_56893;
assign v_56895 = v_56669 & v_56891;
assign v_56897 = v_56667 & v_56896;
assign v_56899 = v_56812 & v_56898;
assign v_56900 = v_56666 & v_56896;
assign v_56902 = v_56901;
assign v_56904 = v_56816 & v_56903;
assign v_56905 = v_56904;
assign v_56907 = v_56906;
assign v_56909 = ~v_2883;
assign v_56910 = ~v_54220;
assign v_56911 = v_54220;
assign v_56912 = ~v_2887;
assign v_56913 = ~v_54224;
assign v_56914 = v_54224;
assign v_56915 = ~v_2891;
assign v_56916 = ~v_54228;
assign v_56917 = v_54228;
assign v_56918 = ~v_2895;
assign v_56919 = ~v_54232;
assign v_56920 = v_54232;
assign v_56921 = ~v_54235;
assign v_56922 = ~v_2900;
assign v_56923 = v_2900;
assign v_56924 = ~v_54239;
assign v_56925 = ~v_2904;
assign v_56926 = v_2904;
assign v_56927 = ~v_54243;
assign v_56928 = ~v_2908;
assign v_56929 = v_2908;
assign v_56930 = ~v_54247;
assign v_56931 = ~v_2912;
assign v_56932 = v_2912;
assign v_56933 = ~v_54251;
assign v_56934 = ~v_2916;
assign v_56935 = v_2916;
assign v_56936 = ~v_54255;
assign v_56937 = ~v_2920;
assign v_56938 = v_2920;
assign v_56939 = ~v_54259;
assign v_56940 = ~v_2924;
assign v_56941 = v_2924;
assign v_56942 = ~v_54263;
assign v_56943 = ~v_2928;
assign v_56944 = v_2928;
assign v_56945 = ~v_54267;
assign v_56946 = ~v_2932;
assign v_56947 = v_2932;
assign v_56948 = ~v_54271;
assign v_56949 = ~v_2936;
assign v_56950 = v_2936;
assign v_56951 = ~v_54275;
assign v_56952 = ~v_2940;
assign v_56953 = v_2940;
assign v_56954 = ~v_54279;
assign v_56955 = ~v_2944;
assign v_56956 = v_2944;
assign v_56957 = ~v_54283;
assign v_56958 = ~v_2948;
assign v_56959 = v_56958;
assign v_56961 = v_56960;
assign v_56963 = v_56955 & v_56962;
assign v_56965 = v_54279;
assign v_56967 = v_56964 & v_56966;
assign v_56969 = v_56952 & v_56968;
assign v_56971 = v_54275;
assign v_56973 = v_56970 & v_56972;
assign v_56975 = v_56949 & v_56974;
assign v_56977 = v_54271;
assign v_56979 = v_56976 & v_56978;
assign v_56981 = v_56946 & v_56980;
assign v_56983 = v_54267;
assign v_56985 = v_56982 & v_56984;
assign v_56987 = v_56943 & v_56986;
assign v_56989 = v_54263;
assign v_56991 = v_56988 & v_56990;
assign v_56993 = v_56940 & v_56992;
assign v_56995 = v_54259;
assign v_56997 = v_56994 & v_56996;
assign v_56999 = v_56937 & v_56998;
assign v_57001 = v_54255;
assign v_57003 = v_57000 & v_57002;
assign v_57005 = v_56934 & v_57004;
assign v_57007 = v_54251;
assign v_57009 = v_57006 & v_57008;
assign v_57011 = v_56931 & v_57010;
assign v_57013 = v_54247;
assign v_57015 = v_57012 & v_57014;
assign v_57017 = v_56928 & v_57016;
assign v_57019 = v_54243;
assign v_57021 = v_57018 & v_57020;
assign v_57023 = v_56925 & v_57022;
assign v_57025 = v_54239;
assign v_57027 = v_57024 & v_57026;
assign v_57029 = v_56922 & v_57028;
assign v_57031 = v_54235;
assign v_57033 = v_57030 & v_57032;
assign v_57035 = v_56919 & v_57034;
assign v_57037 = v_2895;
assign v_57039 = v_57036 & v_57038;
assign v_57041 = v_56916 & v_57040;
assign v_57043 = v_2891;
assign v_57045 = v_57042 & v_57044;
assign v_57047 = v_56913 & v_57046;
assign v_57049 = v_2887;
assign v_57051 = v_57048 & v_57050;
assign v_57053 = v_56910 & v_57052;
assign v_57055 = v_2883;
assign v_57057 = v_57054 & v_57056;
assign v_57058 = v_57057;
assign v_57060 = v_54283;
assign v_57061 = v_2948;
assign v_57062 = v_57061;
assign v_57063 = v_57060 & v_57062;
assign v_57064 = v_57063;
assign v_57065 = v_56955 & v_57064;
assign v_57067 = v_56965 & v_57066;
assign v_57068 = v_56954 & v_57064;
assign v_57070 = v_56952 & v_57069;
assign v_57072 = v_56971 & v_57071;
assign v_57073 = v_56951 & v_57069;
assign v_57075 = v_56949 & v_57074;
assign v_57077 = v_56977 & v_57076;
assign v_57078 = v_56948 & v_57074;
assign v_57080 = v_56946 & v_57079;
assign v_57082 = v_56983 & v_57081;
assign v_57083 = v_56945 & v_57079;
assign v_57085 = v_56943 & v_57084;
assign v_57087 = v_56989 & v_57086;
assign v_57088 = v_56942 & v_57084;
assign v_57090 = v_56940 & v_57089;
assign v_57092 = v_56995 & v_57091;
assign v_57093 = v_56939 & v_57089;
assign v_57095 = v_56937 & v_57094;
assign v_57097 = v_57001 & v_57096;
assign v_57098 = v_56936 & v_57094;
assign v_57100 = v_56934 & v_57099;
assign v_57102 = v_57007 & v_57101;
assign v_57103 = v_56933 & v_57099;
assign v_57105 = v_56931 & v_57104;
assign v_57107 = v_57013 & v_57106;
assign v_57108 = v_56930 & v_57104;
assign v_57110 = v_56928 & v_57109;
assign v_57112 = v_57019 & v_57111;
assign v_57113 = v_56927 & v_57109;
assign v_57115 = v_56925 & v_57114;
assign v_57117 = v_57025 & v_57116;
assign v_57118 = v_56924 & v_57114;
assign v_57120 = v_56922 & v_57119;
assign v_57122 = v_57031 & v_57121;
assign v_57123 = v_56921 & v_57119;
assign v_57125 = v_56919 & v_57124;
assign v_57127 = v_57037 & v_57126;
assign v_57128 = v_56918 & v_57124;
assign v_57130 = v_56916 & v_57129;
assign v_57132 = v_57043 & v_57131;
assign v_57133 = v_56915 & v_57129;
assign v_57135 = v_56913 & v_57134;
assign v_57137 = v_57049 & v_57136;
assign v_57138 = v_56912 & v_57134;
assign v_57140 = v_56910 & v_57139;
assign v_57142 = v_57055 & v_57141;
assign v_57143 = v_56909 & v_57139;
assign v_57145 = v_57144;
assign v_57147 = v_57059 & v_57146;
assign v_57148 = v_57147;
assign v_57150 = v_57149;
assign v_57152 = ~v_3143;
assign v_57153 = ~v_54220;
assign v_57154 = v_54220;
assign v_57155 = ~v_3147;
assign v_57156 = ~v_54224;
assign v_57157 = v_54224;
assign v_57158 = ~v_3151;
assign v_57159 = ~v_54228;
assign v_57160 = v_54228;
assign v_57161 = ~v_3155;
assign v_57162 = ~v_54232;
assign v_57163 = v_54232;
assign v_57164 = ~v_54235;
assign v_57165 = ~v_3160;
assign v_57166 = v_3160;
assign v_57167 = ~v_54239;
assign v_57168 = ~v_3164;
assign v_57169 = v_3164;
assign v_57170 = ~v_54243;
assign v_57171 = ~v_3168;
assign v_57172 = v_3168;
assign v_57173 = ~v_54247;
assign v_57174 = ~v_3172;
assign v_57175 = v_3172;
assign v_57176 = ~v_54251;
assign v_57177 = ~v_3176;
assign v_57178 = v_3176;
assign v_57179 = ~v_54255;
assign v_57180 = ~v_3180;
assign v_57181 = v_3180;
assign v_57182 = ~v_54259;
assign v_57183 = ~v_3184;
assign v_57184 = v_3184;
assign v_57185 = ~v_54263;
assign v_57186 = ~v_3188;
assign v_57187 = v_3188;
assign v_57188 = ~v_54267;
assign v_57189 = ~v_3192;
assign v_57190 = v_3192;
assign v_57191 = ~v_54271;
assign v_57192 = ~v_3196;
assign v_57193 = v_3196;
assign v_57194 = ~v_54275;
assign v_57195 = ~v_3200;
assign v_57196 = v_3200;
assign v_57197 = ~v_54279;
assign v_57198 = ~v_3204;
assign v_57199 = v_3204;
assign v_57200 = ~v_54283;
assign v_57201 = ~v_3208;
assign v_57202 = v_57201;
assign v_57204 = v_57203;
assign v_57206 = v_57198 & v_57205;
assign v_57208 = v_54279;
assign v_57210 = v_57207 & v_57209;
assign v_57212 = v_57195 & v_57211;
assign v_57214 = v_54275;
assign v_57216 = v_57213 & v_57215;
assign v_57218 = v_57192 & v_57217;
assign v_57220 = v_54271;
assign v_57222 = v_57219 & v_57221;
assign v_57224 = v_57189 & v_57223;
assign v_57226 = v_54267;
assign v_57228 = v_57225 & v_57227;
assign v_57230 = v_57186 & v_57229;
assign v_57232 = v_54263;
assign v_57234 = v_57231 & v_57233;
assign v_57236 = v_57183 & v_57235;
assign v_57238 = v_54259;
assign v_57240 = v_57237 & v_57239;
assign v_57242 = v_57180 & v_57241;
assign v_57244 = v_54255;
assign v_57246 = v_57243 & v_57245;
assign v_57248 = v_57177 & v_57247;
assign v_57250 = v_54251;
assign v_57252 = v_57249 & v_57251;
assign v_57254 = v_57174 & v_57253;
assign v_57256 = v_54247;
assign v_57258 = v_57255 & v_57257;
assign v_57260 = v_57171 & v_57259;
assign v_57262 = v_54243;
assign v_57264 = v_57261 & v_57263;
assign v_57266 = v_57168 & v_57265;
assign v_57268 = v_54239;
assign v_57270 = v_57267 & v_57269;
assign v_57272 = v_57165 & v_57271;
assign v_57274 = v_54235;
assign v_57276 = v_57273 & v_57275;
assign v_57278 = v_57162 & v_57277;
assign v_57280 = v_3155;
assign v_57282 = v_57279 & v_57281;
assign v_57284 = v_57159 & v_57283;
assign v_57286 = v_3151;
assign v_57288 = v_57285 & v_57287;
assign v_57290 = v_57156 & v_57289;
assign v_57292 = v_3147;
assign v_57294 = v_57291 & v_57293;
assign v_57296 = v_57153 & v_57295;
assign v_57298 = v_3143;
assign v_57300 = v_57297 & v_57299;
assign v_57301 = v_57300;
assign v_57303 = v_54283;
assign v_57304 = v_3208;
assign v_57305 = v_57304;
assign v_57306 = v_57303 & v_57305;
assign v_57307 = v_57306;
assign v_57308 = v_57198 & v_57307;
assign v_57310 = v_57208 & v_57309;
assign v_57311 = v_57197 & v_57307;
assign v_57313 = v_57195 & v_57312;
assign v_57315 = v_57214 & v_57314;
assign v_57316 = v_57194 & v_57312;
assign v_57318 = v_57192 & v_57317;
assign v_57320 = v_57220 & v_57319;
assign v_57321 = v_57191 & v_57317;
assign v_57323 = v_57189 & v_57322;
assign v_57325 = v_57226 & v_57324;
assign v_57326 = v_57188 & v_57322;
assign v_57328 = v_57186 & v_57327;
assign v_57330 = v_57232 & v_57329;
assign v_57331 = v_57185 & v_57327;
assign v_57333 = v_57183 & v_57332;
assign v_57335 = v_57238 & v_57334;
assign v_57336 = v_57182 & v_57332;
assign v_57338 = v_57180 & v_57337;
assign v_57340 = v_57244 & v_57339;
assign v_57341 = v_57179 & v_57337;
assign v_57343 = v_57177 & v_57342;
assign v_57345 = v_57250 & v_57344;
assign v_57346 = v_57176 & v_57342;
assign v_57348 = v_57174 & v_57347;
assign v_57350 = v_57256 & v_57349;
assign v_57351 = v_57173 & v_57347;
assign v_57353 = v_57171 & v_57352;
assign v_57355 = v_57262 & v_57354;
assign v_57356 = v_57170 & v_57352;
assign v_57358 = v_57168 & v_57357;
assign v_57360 = v_57268 & v_57359;
assign v_57361 = v_57167 & v_57357;
assign v_57363 = v_57165 & v_57362;
assign v_57365 = v_57274 & v_57364;
assign v_57366 = v_57164 & v_57362;
assign v_57368 = v_57162 & v_57367;
assign v_57370 = v_57280 & v_57369;
assign v_57371 = v_57161 & v_57367;
assign v_57373 = v_57159 & v_57372;
assign v_57375 = v_57286 & v_57374;
assign v_57376 = v_57158 & v_57372;
assign v_57378 = v_57156 & v_57377;
assign v_57380 = v_57292 & v_57379;
assign v_57381 = v_57155 & v_57377;
assign v_57383 = v_57153 & v_57382;
assign v_57385 = v_57298 & v_57384;
assign v_57386 = v_57152 & v_57382;
assign v_57388 = v_57387;
assign v_57390 = v_57302 & v_57389;
assign v_57391 = v_57390;
assign v_57393 = v_57392;
assign v_57395 = ~v_3403;
assign v_57396 = ~v_54220;
assign v_57397 = v_54220;
assign v_57398 = ~v_3407;
assign v_57399 = ~v_54224;
assign v_57400 = v_54224;
assign v_57401 = ~v_3411;
assign v_57402 = ~v_54228;
assign v_57403 = v_54228;
assign v_57404 = ~v_3415;
assign v_57405 = ~v_54232;
assign v_57406 = v_54232;
assign v_57407 = ~v_54235;
assign v_57408 = ~v_3420;
assign v_57409 = v_3420;
assign v_57410 = ~v_54239;
assign v_57411 = ~v_3424;
assign v_57412 = v_3424;
assign v_57413 = ~v_54243;
assign v_57414 = ~v_3428;
assign v_57415 = v_3428;
assign v_57416 = ~v_54247;
assign v_57417 = ~v_3432;
assign v_57418 = v_3432;
assign v_57419 = ~v_54251;
assign v_57420 = ~v_3436;
assign v_57421 = v_3436;
assign v_57422 = ~v_54255;
assign v_57423 = ~v_3440;
assign v_57424 = v_3440;
assign v_57425 = ~v_54259;
assign v_57426 = ~v_3444;
assign v_57427 = v_3444;
assign v_57428 = ~v_54263;
assign v_57429 = ~v_3448;
assign v_57430 = v_3448;
assign v_57431 = ~v_54267;
assign v_57432 = ~v_3452;
assign v_57433 = v_3452;
assign v_57434 = ~v_54271;
assign v_57435 = ~v_3456;
assign v_57436 = v_3456;
assign v_57437 = ~v_54275;
assign v_57438 = ~v_3460;
assign v_57439 = v_3460;
assign v_57440 = ~v_54279;
assign v_57441 = ~v_3464;
assign v_57442 = v_3464;
assign v_57443 = ~v_54283;
assign v_57444 = ~v_3468;
assign v_57445 = v_57444;
assign v_57447 = v_57446;
assign v_57449 = v_57441 & v_57448;
assign v_57451 = v_54279;
assign v_57453 = v_57450 & v_57452;
assign v_57455 = v_57438 & v_57454;
assign v_57457 = v_54275;
assign v_57459 = v_57456 & v_57458;
assign v_57461 = v_57435 & v_57460;
assign v_57463 = v_54271;
assign v_57465 = v_57462 & v_57464;
assign v_57467 = v_57432 & v_57466;
assign v_57469 = v_54267;
assign v_57471 = v_57468 & v_57470;
assign v_57473 = v_57429 & v_57472;
assign v_57475 = v_54263;
assign v_57477 = v_57474 & v_57476;
assign v_57479 = v_57426 & v_57478;
assign v_57481 = v_54259;
assign v_57483 = v_57480 & v_57482;
assign v_57485 = v_57423 & v_57484;
assign v_57487 = v_54255;
assign v_57489 = v_57486 & v_57488;
assign v_57491 = v_57420 & v_57490;
assign v_57493 = v_54251;
assign v_57495 = v_57492 & v_57494;
assign v_57497 = v_57417 & v_57496;
assign v_57499 = v_54247;
assign v_57501 = v_57498 & v_57500;
assign v_57503 = v_57414 & v_57502;
assign v_57505 = v_54243;
assign v_57507 = v_57504 & v_57506;
assign v_57509 = v_57411 & v_57508;
assign v_57511 = v_54239;
assign v_57513 = v_57510 & v_57512;
assign v_57515 = v_57408 & v_57514;
assign v_57517 = v_54235;
assign v_57519 = v_57516 & v_57518;
assign v_57521 = v_57405 & v_57520;
assign v_57523 = v_3415;
assign v_57525 = v_57522 & v_57524;
assign v_57527 = v_57402 & v_57526;
assign v_57529 = v_3411;
assign v_57531 = v_57528 & v_57530;
assign v_57533 = v_57399 & v_57532;
assign v_57535 = v_3407;
assign v_57537 = v_57534 & v_57536;
assign v_57539 = v_57396 & v_57538;
assign v_57541 = v_3403;
assign v_57543 = v_57540 & v_57542;
assign v_57544 = v_57543;
assign v_57546 = v_54283;
assign v_57547 = v_3468;
assign v_57548 = v_57547;
assign v_57549 = v_57546 & v_57548;
assign v_57550 = v_57549;
assign v_57551 = v_57441 & v_57550;
assign v_57553 = v_57451 & v_57552;
assign v_57554 = v_57440 & v_57550;
assign v_57556 = v_57438 & v_57555;
assign v_57558 = v_57457 & v_57557;
assign v_57559 = v_57437 & v_57555;
assign v_57561 = v_57435 & v_57560;
assign v_57563 = v_57463 & v_57562;
assign v_57564 = v_57434 & v_57560;
assign v_57566 = v_57432 & v_57565;
assign v_57568 = v_57469 & v_57567;
assign v_57569 = v_57431 & v_57565;
assign v_57571 = v_57429 & v_57570;
assign v_57573 = v_57475 & v_57572;
assign v_57574 = v_57428 & v_57570;
assign v_57576 = v_57426 & v_57575;
assign v_57578 = v_57481 & v_57577;
assign v_57579 = v_57425 & v_57575;
assign v_57581 = v_57423 & v_57580;
assign v_57583 = v_57487 & v_57582;
assign v_57584 = v_57422 & v_57580;
assign v_57586 = v_57420 & v_57585;
assign v_57588 = v_57493 & v_57587;
assign v_57589 = v_57419 & v_57585;
assign v_57591 = v_57417 & v_57590;
assign v_57593 = v_57499 & v_57592;
assign v_57594 = v_57416 & v_57590;
assign v_57596 = v_57414 & v_57595;
assign v_57598 = v_57505 & v_57597;
assign v_57599 = v_57413 & v_57595;
assign v_57601 = v_57411 & v_57600;
assign v_57603 = v_57511 & v_57602;
assign v_57604 = v_57410 & v_57600;
assign v_57606 = v_57408 & v_57605;
assign v_57608 = v_57517 & v_57607;
assign v_57609 = v_57407 & v_57605;
assign v_57611 = v_57405 & v_57610;
assign v_57613 = v_57523 & v_57612;
assign v_57614 = v_57404 & v_57610;
assign v_57616 = v_57402 & v_57615;
assign v_57618 = v_57529 & v_57617;
assign v_57619 = v_57401 & v_57615;
assign v_57621 = v_57399 & v_57620;
assign v_57623 = v_57535 & v_57622;
assign v_57624 = v_57398 & v_57620;
assign v_57626 = v_57396 & v_57625;
assign v_57628 = v_57541 & v_57627;
assign v_57629 = v_57395 & v_57625;
assign v_57631 = v_57630;
assign v_57633 = v_57545 & v_57632;
assign v_57634 = v_57633;
assign v_57636 = v_57635;
assign v_57638 = ~v_3663;
assign v_57639 = ~v_54220;
assign v_57640 = v_54220;
assign v_57641 = ~v_3667;
assign v_57642 = ~v_54224;
assign v_57643 = v_54224;
assign v_57644 = ~v_3671;
assign v_57645 = ~v_54228;
assign v_57646 = v_54228;
assign v_57647 = ~v_3675;
assign v_57648 = ~v_54232;
assign v_57649 = v_54232;
assign v_57650 = ~v_54235;
assign v_57651 = ~v_3680;
assign v_57652 = v_3680;
assign v_57653 = ~v_54239;
assign v_57654 = ~v_3684;
assign v_57655 = v_3684;
assign v_57656 = ~v_54243;
assign v_57657 = ~v_3688;
assign v_57658 = v_3688;
assign v_57659 = ~v_54247;
assign v_57660 = ~v_3692;
assign v_57661 = v_3692;
assign v_57662 = ~v_54251;
assign v_57663 = ~v_3696;
assign v_57664 = v_3696;
assign v_57665 = ~v_54255;
assign v_57666 = ~v_3700;
assign v_57667 = v_3700;
assign v_57668 = ~v_54259;
assign v_57669 = ~v_3704;
assign v_57670 = v_3704;
assign v_57671 = ~v_54263;
assign v_57672 = ~v_3708;
assign v_57673 = v_3708;
assign v_57674 = ~v_54267;
assign v_57675 = ~v_3712;
assign v_57676 = v_3712;
assign v_57677 = ~v_54271;
assign v_57678 = ~v_3716;
assign v_57679 = v_3716;
assign v_57680 = ~v_54275;
assign v_57681 = ~v_3720;
assign v_57682 = v_3720;
assign v_57683 = ~v_54279;
assign v_57684 = ~v_3724;
assign v_57685 = v_3724;
assign v_57686 = ~v_54283;
assign v_57687 = ~v_3728;
assign v_57688 = v_57687;
assign v_57690 = v_57689;
assign v_57692 = v_57684 & v_57691;
assign v_57694 = v_54279;
assign v_57696 = v_57693 & v_57695;
assign v_57698 = v_57681 & v_57697;
assign v_57700 = v_54275;
assign v_57702 = v_57699 & v_57701;
assign v_57704 = v_57678 & v_57703;
assign v_57706 = v_54271;
assign v_57708 = v_57705 & v_57707;
assign v_57710 = v_57675 & v_57709;
assign v_57712 = v_54267;
assign v_57714 = v_57711 & v_57713;
assign v_57716 = v_57672 & v_57715;
assign v_57718 = v_54263;
assign v_57720 = v_57717 & v_57719;
assign v_57722 = v_57669 & v_57721;
assign v_57724 = v_54259;
assign v_57726 = v_57723 & v_57725;
assign v_57728 = v_57666 & v_57727;
assign v_57730 = v_54255;
assign v_57732 = v_57729 & v_57731;
assign v_57734 = v_57663 & v_57733;
assign v_57736 = v_54251;
assign v_57738 = v_57735 & v_57737;
assign v_57740 = v_57660 & v_57739;
assign v_57742 = v_54247;
assign v_57744 = v_57741 & v_57743;
assign v_57746 = v_57657 & v_57745;
assign v_57748 = v_54243;
assign v_57750 = v_57747 & v_57749;
assign v_57752 = v_57654 & v_57751;
assign v_57754 = v_54239;
assign v_57756 = v_57753 & v_57755;
assign v_57758 = v_57651 & v_57757;
assign v_57760 = v_54235;
assign v_57762 = v_57759 & v_57761;
assign v_57764 = v_57648 & v_57763;
assign v_57766 = v_3675;
assign v_57768 = v_57765 & v_57767;
assign v_57770 = v_57645 & v_57769;
assign v_57772 = v_3671;
assign v_57774 = v_57771 & v_57773;
assign v_57776 = v_57642 & v_57775;
assign v_57778 = v_3667;
assign v_57780 = v_57777 & v_57779;
assign v_57782 = v_57639 & v_57781;
assign v_57784 = v_3663;
assign v_57786 = v_57783 & v_57785;
assign v_57787 = v_57786;
assign v_57789 = v_54283;
assign v_57790 = v_3728;
assign v_57791 = v_57790;
assign v_57792 = v_57789 & v_57791;
assign v_57793 = v_57792;
assign v_57794 = v_57684 & v_57793;
assign v_57796 = v_57694 & v_57795;
assign v_57797 = v_57683 & v_57793;
assign v_57799 = v_57681 & v_57798;
assign v_57801 = v_57700 & v_57800;
assign v_57802 = v_57680 & v_57798;
assign v_57804 = v_57678 & v_57803;
assign v_57806 = v_57706 & v_57805;
assign v_57807 = v_57677 & v_57803;
assign v_57809 = v_57675 & v_57808;
assign v_57811 = v_57712 & v_57810;
assign v_57812 = v_57674 & v_57808;
assign v_57814 = v_57672 & v_57813;
assign v_57816 = v_57718 & v_57815;
assign v_57817 = v_57671 & v_57813;
assign v_57819 = v_57669 & v_57818;
assign v_57821 = v_57724 & v_57820;
assign v_57822 = v_57668 & v_57818;
assign v_57824 = v_57666 & v_57823;
assign v_57826 = v_57730 & v_57825;
assign v_57827 = v_57665 & v_57823;
assign v_57829 = v_57663 & v_57828;
assign v_57831 = v_57736 & v_57830;
assign v_57832 = v_57662 & v_57828;
assign v_57834 = v_57660 & v_57833;
assign v_57836 = v_57742 & v_57835;
assign v_57837 = v_57659 & v_57833;
assign v_57839 = v_57657 & v_57838;
assign v_57841 = v_57748 & v_57840;
assign v_57842 = v_57656 & v_57838;
assign v_57844 = v_57654 & v_57843;
assign v_57846 = v_57754 & v_57845;
assign v_57847 = v_57653 & v_57843;
assign v_57849 = v_57651 & v_57848;
assign v_57851 = v_57760 & v_57850;
assign v_57852 = v_57650 & v_57848;
assign v_57854 = v_57648 & v_57853;
assign v_57856 = v_57766 & v_57855;
assign v_57857 = v_57647 & v_57853;
assign v_57859 = v_57645 & v_57858;
assign v_57861 = v_57772 & v_57860;
assign v_57862 = v_57644 & v_57858;
assign v_57864 = v_57642 & v_57863;
assign v_57866 = v_57778 & v_57865;
assign v_57867 = v_57641 & v_57863;
assign v_57869 = v_57639 & v_57868;
assign v_57871 = v_57784 & v_57870;
assign v_57872 = v_57638 & v_57868;
assign v_57874 = v_57873;
assign v_57876 = v_57788 & v_57875;
assign v_57877 = v_57876;
assign v_57879 = v_57878;
assign v_57881 = ~v_3923;
assign v_57882 = ~v_54220;
assign v_57883 = v_54220;
assign v_57884 = ~v_3927;
assign v_57885 = ~v_54224;
assign v_57886 = v_54224;
assign v_57887 = ~v_3931;
assign v_57888 = ~v_54228;
assign v_57889 = v_54228;
assign v_57890 = ~v_3935;
assign v_57891 = ~v_54232;
assign v_57892 = v_54232;
assign v_57893 = ~v_54235;
assign v_57894 = ~v_3940;
assign v_57895 = v_3940;
assign v_57896 = ~v_54239;
assign v_57897 = ~v_3944;
assign v_57898 = v_3944;
assign v_57899 = ~v_54243;
assign v_57900 = ~v_3948;
assign v_57901 = v_3948;
assign v_57902 = ~v_54247;
assign v_57903 = ~v_3952;
assign v_57904 = v_3952;
assign v_57905 = ~v_54251;
assign v_57906 = ~v_3956;
assign v_57907 = v_3956;
assign v_57908 = ~v_54255;
assign v_57909 = ~v_3960;
assign v_57910 = v_3960;
assign v_57911 = ~v_54259;
assign v_57912 = ~v_3964;
assign v_57913 = v_3964;
assign v_57914 = ~v_54263;
assign v_57915 = ~v_3968;
assign v_57916 = v_3968;
assign v_57917 = ~v_54267;
assign v_57918 = ~v_3972;
assign v_57919 = v_3972;
assign v_57920 = ~v_54271;
assign v_57921 = ~v_3976;
assign v_57922 = v_3976;
assign v_57923 = ~v_54275;
assign v_57924 = ~v_3980;
assign v_57925 = v_3980;
assign v_57926 = ~v_54279;
assign v_57927 = ~v_3984;
assign v_57928 = v_3984;
assign v_57929 = ~v_54283;
assign v_57930 = ~v_3988;
assign v_57931 = v_57930;
assign v_57933 = v_57932;
assign v_57935 = v_57927 & v_57934;
assign v_57937 = v_54279;
assign v_57939 = v_57936 & v_57938;
assign v_57941 = v_57924 & v_57940;
assign v_57943 = v_54275;
assign v_57945 = v_57942 & v_57944;
assign v_57947 = v_57921 & v_57946;
assign v_57949 = v_54271;
assign v_57951 = v_57948 & v_57950;
assign v_57953 = v_57918 & v_57952;
assign v_57955 = v_54267;
assign v_57957 = v_57954 & v_57956;
assign v_57959 = v_57915 & v_57958;
assign v_57961 = v_54263;
assign v_57963 = v_57960 & v_57962;
assign v_57965 = v_57912 & v_57964;
assign v_57967 = v_54259;
assign v_57969 = v_57966 & v_57968;
assign v_57971 = v_57909 & v_57970;
assign v_57973 = v_54255;
assign v_57975 = v_57972 & v_57974;
assign v_57977 = v_57906 & v_57976;
assign v_57979 = v_54251;
assign v_57981 = v_57978 & v_57980;
assign v_57983 = v_57903 & v_57982;
assign v_57985 = v_54247;
assign v_57987 = v_57984 & v_57986;
assign v_57989 = v_57900 & v_57988;
assign v_57991 = v_54243;
assign v_57993 = v_57990 & v_57992;
assign v_57995 = v_57897 & v_57994;
assign v_57997 = v_54239;
assign v_57999 = v_57996 & v_57998;
assign v_58001 = v_57894 & v_58000;
assign v_58003 = v_54235;
assign v_58005 = v_58002 & v_58004;
assign v_58007 = v_57891 & v_58006;
assign v_58009 = v_3935;
assign v_58011 = v_58008 & v_58010;
assign v_58013 = v_57888 & v_58012;
assign v_58015 = v_3931;
assign v_58017 = v_58014 & v_58016;
assign v_58019 = v_57885 & v_58018;
assign v_58021 = v_3927;
assign v_58023 = v_58020 & v_58022;
assign v_58025 = v_57882 & v_58024;
assign v_58027 = v_3923;
assign v_58029 = v_58026 & v_58028;
assign v_58030 = v_58029;
assign v_58032 = v_54283;
assign v_58033 = v_3988;
assign v_58034 = v_58033;
assign v_58035 = v_58032 & v_58034;
assign v_58036 = v_58035;
assign v_58037 = v_57927 & v_58036;
assign v_58039 = v_57937 & v_58038;
assign v_58040 = v_57926 & v_58036;
assign v_58042 = v_57924 & v_58041;
assign v_58044 = v_57943 & v_58043;
assign v_58045 = v_57923 & v_58041;
assign v_58047 = v_57921 & v_58046;
assign v_58049 = v_57949 & v_58048;
assign v_58050 = v_57920 & v_58046;
assign v_58052 = v_57918 & v_58051;
assign v_58054 = v_57955 & v_58053;
assign v_58055 = v_57917 & v_58051;
assign v_58057 = v_57915 & v_58056;
assign v_58059 = v_57961 & v_58058;
assign v_58060 = v_57914 & v_58056;
assign v_58062 = v_57912 & v_58061;
assign v_58064 = v_57967 & v_58063;
assign v_58065 = v_57911 & v_58061;
assign v_58067 = v_57909 & v_58066;
assign v_58069 = v_57973 & v_58068;
assign v_58070 = v_57908 & v_58066;
assign v_58072 = v_57906 & v_58071;
assign v_58074 = v_57979 & v_58073;
assign v_58075 = v_57905 & v_58071;
assign v_58077 = v_57903 & v_58076;
assign v_58079 = v_57985 & v_58078;
assign v_58080 = v_57902 & v_58076;
assign v_58082 = v_57900 & v_58081;
assign v_58084 = v_57991 & v_58083;
assign v_58085 = v_57899 & v_58081;
assign v_58087 = v_57897 & v_58086;
assign v_58089 = v_57997 & v_58088;
assign v_58090 = v_57896 & v_58086;
assign v_58092 = v_57894 & v_58091;
assign v_58094 = v_58003 & v_58093;
assign v_58095 = v_57893 & v_58091;
assign v_58097 = v_57891 & v_58096;
assign v_58099 = v_58009 & v_58098;
assign v_58100 = v_57890 & v_58096;
assign v_58102 = v_57888 & v_58101;
assign v_58104 = v_58015 & v_58103;
assign v_58105 = v_57887 & v_58101;
assign v_58107 = v_57885 & v_58106;
assign v_58109 = v_58021 & v_58108;
assign v_58110 = v_57884 & v_58106;
assign v_58112 = v_57882 & v_58111;
assign v_58114 = v_58027 & v_58113;
assign v_58115 = v_57881 & v_58111;
assign v_58117 = v_58116;
assign v_58119 = v_58031 & v_58118;
assign v_58120 = v_58119;
assign v_58122 = v_58121;
assign v_58123 = ~v_4182;
assign v_58124 = ~v_54220;
assign v_58125 = v_54220;
assign v_58126 = ~v_4186;
assign v_58127 = ~v_54224;
assign v_58128 = v_54224;
assign v_58129 = ~v_4190;
assign v_58130 = ~v_54228;
assign v_58131 = v_54228;
assign v_58132 = ~v_4194;
assign v_58133 = ~v_54232;
assign v_58134 = v_54232;
assign v_58135 = ~v_54235;
assign v_58136 = ~v_4199;
assign v_58137 = v_4199;
assign v_58138 = ~v_54239;
assign v_58139 = ~v_4203;
assign v_58140 = v_4203;
assign v_58141 = ~v_54243;
assign v_58142 = ~v_4207;
assign v_58143 = v_4207;
assign v_58144 = ~v_54247;
assign v_58145 = ~v_4211;
assign v_58146 = v_4211;
assign v_58147 = ~v_54251;
assign v_58148 = ~v_4215;
assign v_58149 = v_4215;
assign v_58150 = ~v_54255;
assign v_58151 = ~v_4219;
assign v_58152 = v_4219;
assign v_58153 = ~v_54259;
assign v_58154 = ~v_4223;
assign v_58155 = v_4223;
assign v_58156 = ~v_54263;
assign v_58157 = ~v_4227;
assign v_58158 = v_4227;
assign v_58159 = ~v_54267;
assign v_58160 = ~v_4231;
assign v_58161 = v_4231;
assign v_58162 = ~v_54271;
assign v_58163 = ~v_4235;
assign v_58164 = v_4235;
assign v_58165 = ~v_54275;
assign v_58166 = ~v_4239;
assign v_58167 = v_4239;
assign v_58168 = ~v_54279;
assign v_58169 = ~v_4243;
assign v_58170 = v_4243;
assign v_58171 = ~v_54283;
assign v_58172 = ~v_4247;
assign v_58173 = v_58172;
assign v_58175 = v_58174;
assign v_58177 = v_58169 & v_58176;
assign v_58179 = v_54279;
assign v_58181 = v_58178 & v_58180;
assign v_58183 = v_58166 & v_58182;
assign v_58185 = v_54275;
assign v_58187 = v_58184 & v_58186;
assign v_58189 = v_58163 & v_58188;
assign v_58191 = v_54271;
assign v_58193 = v_58190 & v_58192;
assign v_58195 = v_58160 & v_58194;
assign v_58197 = v_54267;
assign v_58199 = v_58196 & v_58198;
assign v_58201 = v_58157 & v_58200;
assign v_58203 = v_54263;
assign v_58205 = v_58202 & v_58204;
assign v_58207 = v_58154 & v_58206;
assign v_58209 = v_54259;
assign v_58211 = v_58208 & v_58210;
assign v_58213 = v_58151 & v_58212;
assign v_58215 = v_54255;
assign v_58217 = v_58214 & v_58216;
assign v_58219 = v_58148 & v_58218;
assign v_58221 = v_54251;
assign v_58223 = v_58220 & v_58222;
assign v_58225 = v_58145 & v_58224;
assign v_58227 = v_54247;
assign v_58229 = v_58226 & v_58228;
assign v_58231 = v_58142 & v_58230;
assign v_58233 = v_54243;
assign v_58235 = v_58232 & v_58234;
assign v_58237 = v_58139 & v_58236;
assign v_58239 = v_54239;
assign v_58241 = v_58238 & v_58240;
assign v_58243 = v_58136 & v_58242;
assign v_58245 = v_54235;
assign v_58247 = v_58244 & v_58246;
assign v_58249 = v_58133 & v_58248;
assign v_58251 = v_4194;
assign v_58253 = v_58250 & v_58252;
assign v_58255 = v_58130 & v_58254;
assign v_58257 = v_4190;
assign v_58259 = v_58256 & v_58258;
assign v_58261 = v_58127 & v_58260;
assign v_58263 = v_4186;
assign v_58265 = v_58262 & v_58264;
assign v_58267 = v_58124 & v_58266;
assign v_58269 = v_4182;
assign v_58271 = v_58268 & v_58270;
assign v_58273 = ~v_58272;
assign v_58275 = v_54283;
assign v_58276 = v_4247;
assign v_58277 = v_58276;
assign v_58278 = v_58275 & v_58277;
assign v_58279 = v_58278;
assign v_58280 = v_58169 & v_58279;
assign v_58282 = v_58179 & v_58281;
assign v_58283 = v_58168 & v_58279;
assign v_58285 = v_58166 & v_58284;
assign v_58287 = v_58185 & v_58286;
assign v_58288 = v_58165 & v_58284;
assign v_58290 = v_58163 & v_58289;
assign v_58292 = v_58191 & v_58291;
assign v_58293 = v_58162 & v_58289;
assign v_58295 = v_58160 & v_58294;
assign v_58297 = v_58197 & v_58296;
assign v_58298 = v_58159 & v_58294;
assign v_58300 = v_58157 & v_58299;
assign v_58302 = v_58203 & v_58301;
assign v_58303 = v_58156 & v_58299;
assign v_58305 = v_58154 & v_58304;
assign v_58307 = v_58209 & v_58306;
assign v_58308 = v_58153 & v_58304;
assign v_58310 = v_58151 & v_58309;
assign v_58312 = v_58215 & v_58311;
assign v_58313 = v_58150 & v_58309;
assign v_58315 = v_58148 & v_58314;
assign v_58317 = v_58221 & v_58316;
assign v_58318 = v_58147 & v_58314;
assign v_58320 = v_58145 & v_58319;
assign v_58322 = v_58227 & v_58321;
assign v_58323 = v_58144 & v_58319;
assign v_58325 = v_58142 & v_58324;
assign v_58327 = v_58233 & v_58326;
assign v_58328 = v_58141 & v_58324;
assign v_58330 = v_58139 & v_58329;
assign v_58332 = v_58239 & v_58331;
assign v_58333 = v_58138 & v_58329;
assign v_58335 = v_58136 & v_58334;
assign v_58337 = v_58245 & v_58336;
assign v_58338 = v_58135 & v_58334;
assign v_58340 = v_58133 & v_58339;
assign v_58342 = v_58251 & v_58341;
assign v_58343 = v_58132 & v_58339;
assign v_58345 = v_58130 & v_58344;
assign v_58347 = v_58257 & v_58346;
assign v_58348 = v_58129 & v_58344;
assign v_58350 = v_58127 & v_58349;
assign v_58352 = v_58263 & v_58351;
assign v_58353 = v_58126 & v_58349;
assign v_58355 = v_58124 & v_58354;
assign v_58357 = v_58269 & v_58356;
assign v_58358 = v_58123 & v_58354;
assign v_58360 = v_58272;
assign v_58362 = v_58274 & v_58361;
assign v_58363 = v_58362;
assign v_58365 = v_58364;
assign v_58367 = ~v_6;
assign v_58369 = ~v_58368;
assign v_58370 = v_58368;
assign v_58371 = ~v_13;
assign v_58373 = ~v_58372;
assign v_58374 = v_58372;
assign v_58375 = ~v_18;
assign v_58377 = ~v_58376;
assign v_58378 = v_58376;
assign v_58379 = ~v_23;
assign v_58381 = ~v_58380;
assign v_58382 = v_58380;
assign v_58384 = ~v_58383;
assign v_58385 = ~v_30;
assign v_58386 = v_30;
assign v_58388 = ~v_58387;
assign v_58389 = ~v_35;
assign v_58390 = v_35;
assign v_58392 = ~v_58391;
assign v_58393 = ~v_40;
assign v_58394 = v_40;
assign v_58396 = ~v_58395;
assign v_58397 = ~v_45;
assign v_58398 = v_45;
assign v_58400 = ~v_58399;
assign v_58401 = ~v_50;
assign v_58402 = v_50;
assign v_58404 = ~v_58403;
assign v_58405 = ~v_55;
assign v_58406 = v_55;
assign v_58408 = ~v_58407;
assign v_58409 = ~v_60;
assign v_58410 = v_60;
assign v_58412 = ~v_58411;
assign v_58413 = ~v_65;
assign v_58414 = v_65;
assign v_58416 = ~v_58415;
assign v_58417 = ~v_70;
assign v_58418 = v_70;
assign v_58420 = ~v_58419;
assign v_58421 = ~v_75;
assign v_58422 = v_75;
assign v_58424 = ~v_58423;
assign v_58425 = ~v_80;
assign v_58426 = v_80;
assign v_58428 = ~v_58427;
assign v_58429 = ~v_85;
assign v_58430 = v_85;
assign v_58432 = ~v_58431;
assign v_58433 = ~v_90;
assign v_58434 = v_58433;
assign v_58436 = v_58435;
assign v_58438 = v_58429 & v_58437;
assign v_58440 = v_58427;
assign v_58442 = v_58439 & v_58441;
assign v_58444 = v_58425 & v_58443;
assign v_58446 = v_58423;
assign v_58448 = v_58445 & v_58447;
assign v_58450 = v_58421 & v_58449;
assign v_58452 = v_58419;
assign v_58454 = v_58451 & v_58453;
assign v_58456 = v_58417 & v_58455;
assign v_58458 = v_58415;
assign v_58460 = v_58457 & v_58459;
assign v_58462 = v_58413 & v_58461;
assign v_58464 = v_58411;
assign v_58466 = v_58463 & v_58465;
assign v_58468 = v_58409 & v_58467;
assign v_58470 = v_58407;
assign v_58472 = v_58469 & v_58471;
assign v_58474 = v_58405 & v_58473;
assign v_58476 = v_58403;
assign v_58478 = v_58475 & v_58477;
assign v_58480 = v_58401 & v_58479;
assign v_58482 = v_58399;
assign v_58484 = v_58481 & v_58483;
assign v_58486 = v_58397 & v_58485;
assign v_58488 = v_58395;
assign v_58490 = v_58487 & v_58489;
assign v_58492 = v_58393 & v_58491;
assign v_58494 = v_58391;
assign v_58496 = v_58493 & v_58495;
assign v_58498 = v_58389 & v_58497;
assign v_58500 = v_58387;
assign v_58502 = v_58499 & v_58501;
assign v_58504 = v_58385 & v_58503;
assign v_58506 = v_58383;
assign v_58508 = v_58505 & v_58507;
assign v_58510 = v_58381 & v_58509;
assign v_58512 = v_23;
assign v_58514 = v_58511 & v_58513;
assign v_58516 = v_58377 & v_58515;
assign v_58518 = v_18;
assign v_58520 = v_58517 & v_58519;
assign v_58522 = v_58373 & v_58521;
assign v_58524 = v_13;
assign v_58526 = v_58523 & v_58525;
assign v_58528 = v_58369 & v_58527;
assign v_58530 = v_6;
assign v_58532 = v_58529 & v_58531;
assign v_58533 = v_58532;
assign v_58535 = v_58431;
assign v_58536 = v_90;
assign v_58537 = v_58536;
assign v_58538 = v_58535 & v_58537;
assign v_58539 = v_58538;
assign v_58540 = v_58429 & v_58539;
assign v_58542 = v_58440 & v_58541;
assign v_58543 = v_58428 & v_58539;
assign v_58545 = v_58425 & v_58544;
assign v_58547 = v_58446 & v_58546;
assign v_58548 = v_58424 & v_58544;
assign v_58550 = v_58421 & v_58549;
assign v_58552 = v_58452 & v_58551;
assign v_58553 = v_58420 & v_58549;
assign v_58555 = v_58417 & v_58554;
assign v_58557 = v_58458 & v_58556;
assign v_58558 = v_58416 & v_58554;
assign v_58560 = v_58413 & v_58559;
assign v_58562 = v_58464 & v_58561;
assign v_58563 = v_58412 & v_58559;
assign v_58565 = v_58409 & v_58564;
assign v_58567 = v_58470 & v_58566;
assign v_58568 = v_58408 & v_58564;
assign v_58570 = v_58405 & v_58569;
assign v_58572 = v_58476 & v_58571;
assign v_58573 = v_58404 & v_58569;
assign v_58575 = v_58401 & v_58574;
assign v_58577 = v_58482 & v_58576;
assign v_58578 = v_58400 & v_58574;
assign v_58580 = v_58397 & v_58579;
assign v_58582 = v_58488 & v_58581;
assign v_58583 = v_58396 & v_58579;
assign v_58585 = v_58393 & v_58584;
assign v_58587 = v_58494 & v_58586;
assign v_58588 = v_58392 & v_58584;
assign v_58590 = v_58389 & v_58589;
assign v_58592 = v_58500 & v_58591;
assign v_58593 = v_58388 & v_58589;
assign v_58595 = v_58385 & v_58594;
assign v_58597 = v_58506 & v_58596;
assign v_58598 = v_58384 & v_58594;
assign v_58600 = v_58381 & v_58599;
assign v_58602 = v_58512 & v_58601;
assign v_58603 = v_58379 & v_58599;
assign v_58605 = v_58377 & v_58604;
assign v_58607 = v_58518 & v_58606;
assign v_58608 = v_58375 & v_58604;
assign v_58610 = v_58373 & v_58609;
assign v_58612 = v_58524 & v_58611;
assign v_58613 = v_58371 & v_58609;
assign v_58615 = v_58369 & v_58614;
assign v_58617 = v_58530 & v_58616;
assign v_58618 = v_58367 & v_58614;
assign v_58620 = v_58619;
assign v_58622 = v_58534 & v_58621;
assign v_58623 = v_58622;
assign v_58625 = v_58624;
assign v_58627 = ~v_283;
assign v_58628 = ~v_58368;
assign v_58629 = v_58368;
assign v_58630 = ~v_287;
assign v_58631 = ~v_58372;
assign v_58632 = v_58372;
assign v_58633 = ~v_291;
assign v_58634 = ~v_58376;
assign v_58635 = v_58376;
assign v_58636 = ~v_295;
assign v_58637 = ~v_58380;
assign v_58638 = v_58380;
assign v_58639 = ~v_58383;
assign v_58640 = ~v_300;
assign v_58641 = v_300;
assign v_58642 = ~v_58387;
assign v_58643 = ~v_304;
assign v_58644 = v_304;
assign v_58645 = ~v_58391;
assign v_58646 = ~v_308;
assign v_58647 = v_308;
assign v_58648 = ~v_58395;
assign v_58649 = ~v_312;
assign v_58650 = v_312;
assign v_58651 = ~v_58399;
assign v_58652 = ~v_316;
assign v_58653 = v_316;
assign v_58654 = ~v_58403;
assign v_58655 = ~v_320;
assign v_58656 = v_320;
assign v_58657 = ~v_58407;
assign v_58658 = ~v_324;
assign v_58659 = v_324;
assign v_58660 = ~v_58411;
assign v_58661 = ~v_328;
assign v_58662 = v_328;
assign v_58663 = ~v_58415;
assign v_58664 = ~v_332;
assign v_58665 = v_332;
assign v_58666 = ~v_58419;
assign v_58667 = ~v_336;
assign v_58668 = v_336;
assign v_58669 = ~v_58423;
assign v_58670 = ~v_340;
assign v_58671 = v_340;
assign v_58672 = ~v_58427;
assign v_58673 = ~v_344;
assign v_58674 = v_344;
assign v_58675 = ~v_58431;
assign v_58676 = ~v_348;
assign v_58677 = v_58676;
assign v_58679 = v_58678;
assign v_58681 = v_58673 & v_58680;
assign v_58683 = v_58427;
assign v_58685 = v_58682 & v_58684;
assign v_58687 = v_58670 & v_58686;
assign v_58689 = v_58423;
assign v_58691 = v_58688 & v_58690;
assign v_58693 = v_58667 & v_58692;
assign v_58695 = v_58419;
assign v_58697 = v_58694 & v_58696;
assign v_58699 = v_58664 & v_58698;
assign v_58701 = v_58415;
assign v_58703 = v_58700 & v_58702;
assign v_58705 = v_58661 & v_58704;
assign v_58707 = v_58411;
assign v_58709 = v_58706 & v_58708;
assign v_58711 = v_58658 & v_58710;
assign v_58713 = v_58407;
assign v_58715 = v_58712 & v_58714;
assign v_58717 = v_58655 & v_58716;
assign v_58719 = v_58403;
assign v_58721 = v_58718 & v_58720;
assign v_58723 = v_58652 & v_58722;
assign v_58725 = v_58399;
assign v_58727 = v_58724 & v_58726;
assign v_58729 = v_58649 & v_58728;
assign v_58731 = v_58395;
assign v_58733 = v_58730 & v_58732;
assign v_58735 = v_58646 & v_58734;
assign v_58737 = v_58391;
assign v_58739 = v_58736 & v_58738;
assign v_58741 = v_58643 & v_58740;
assign v_58743 = v_58387;
assign v_58745 = v_58742 & v_58744;
assign v_58747 = v_58640 & v_58746;
assign v_58749 = v_58383;
assign v_58751 = v_58748 & v_58750;
assign v_58753 = v_58637 & v_58752;
assign v_58755 = v_295;
assign v_58757 = v_58754 & v_58756;
assign v_58759 = v_58634 & v_58758;
assign v_58761 = v_291;
assign v_58763 = v_58760 & v_58762;
assign v_58765 = v_58631 & v_58764;
assign v_58767 = v_287;
assign v_58769 = v_58766 & v_58768;
assign v_58771 = v_58628 & v_58770;
assign v_58773 = v_283;
assign v_58775 = v_58772 & v_58774;
assign v_58776 = v_58775;
assign v_58778 = v_58431;
assign v_58779 = v_348;
assign v_58780 = v_58779;
assign v_58781 = v_58778 & v_58780;
assign v_58782 = v_58781;
assign v_58783 = v_58673 & v_58782;
assign v_58785 = v_58683 & v_58784;
assign v_58786 = v_58672 & v_58782;
assign v_58788 = v_58670 & v_58787;
assign v_58790 = v_58689 & v_58789;
assign v_58791 = v_58669 & v_58787;
assign v_58793 = v_58667 & v_58792;
assign v_58795 = v_58695 & v_58794;
assign v_58796 = v_58666 & v_58792;
assign v_58798 = v_58664 & v_58797;
assign v_58800 = v_58701 & v_58799;
assign v_58801 = v_58663 & v_58797;
assign v_58803 = v_58661 & v_58802;
assign v_58805 = v_58707 & v_58804;
assign v_58806 = v_58660 & v_58802;
assign v_58808 = v_58658 & v_58807;
assign v_58810 = v_58713 & v_58809;
assign v_58811 = v_58657 & v_58807;
assign v_58813 = v_58655 & v_58812;
assign v_58815 = v_58719 & v_58814;
assign v_58816 = v_58654 & v_58812;
assign v_58818 = v_58652 & v_58817;
assign v_58820 = v_58725 & v_58819;
assign v_58821 = v_58651 & v_58817;
assign v_58823 = v_58649 & v_58822;
assign v_58825 = v_58731 & v_58824;
assign v_58826 = v_58648 & v_58822;
assign v_58828 = v_58646 & v_58827;
assign v_58830 = v_58737 & v_58829;
assign v_58831 = v_58645 & v_58827;
assign v_58833 = v_58643 & v_58832;
assign v_58835 = v_58743 & v_58834;
assign v_58836 = v_58642 & v_58832;
assign v_58838 = v_58640 & v_58837;
assign v_58840 = v_58749 & v_58839;
assign v_58841 = v_58639 & v_58837;
assign v_58843 = v_58637 & v_58842;
assign v_58845 = v_58755 & v_58844;
assign v_58846 = v_58636 & v_58842;
assign v_58848 = v_58634 & v_58847;
assign v_58850 = v_58761 & v_58849;
assign v_58851 = v_58633 & v_58847;
assign v_58853 = v_58631 & v_58852;
assign v_58855 = v_58767 & v_58854;
assign v_58856 = v_58630 & v_58852;
assign v_58858 = v_58628 & v_58857;
assign v_58860 = v_58773 & v_58859;
assign v_58861 = v_58627 & v_58857;
assign v_58863 = v_58862;
assign v_58865 = v_58777 & v_58864;
assign v_58866 = v_58865;
assign v_58868 = v_58867;
assign v_58870 = ~v_543;
assign v_58871 = ~v_58368;
assign v_58872 = v_58368;
assign v_58873 = ~v_547;
assign v_58874 = ~v_58372;
assign v_58875 = v_58372;
assign v_58876 = ~v_551;
assign v_58877 = ~v_58376;
assign v_58878 = v_58376;
assign v_58879 = ~v_555;
assign v_58880 = ~v_58380;
assign v_58881 = v_58380;
assign v_58882 = ~v_58383;
assign v_58883 = ~v_560;
assign v_58884 = v_560;
assign v_58885 = ~v_58387;
assign v_58886 = ~v_564;
assign v_58887 = v_564;
assign v_58888 = ~v_58391;
assign v_58889 = ~v_568;
assign v_58890 = v_568;
assign v_58891 = ~v_58395;
assign v_58892 = ~v_572;
assign v_58893 = v_572;
assign v_58894 = ~v_58399;
assign v_58895 = ~v_576;
assign v_58896 = v_576;
assign v_58897 = ~v_58403;
assign v_58898 = ~v_580;
assign v_58899 = v_580;
assign v_58900 = ~v_58407;
assign v_58901 = ~v_584;
assign v_58902 = v_584;
assign v_58903 = ~v_58411;
assign v_58904 = ~v_588;
assign v_58905 = v_588;
assign v_58906 = ~v_58415;
assign v_58907 = ~v_592;
assign v_58908 = v_592;
assign v_58909 = ~v_58419;
assign v_58910 = ~v_596;
assign v_58911 = v_596;
assign v_58912 = ~v_58423;
assign v_58913 = ~v_600;
assign v_58914 = v_600;
assign v_58915 = ~v_58427;
assign v_58916 = ~v_604;
assign v_58917 = v_604;
assign v_58918 = ~v_58431;
assign v_58919 = ~v_608;
assign v_58920 = v_58919;
assign v_58922 = v_58921;
assign v_58924 = v_58916 & v_58923;
assign v_58926 = v_58427;
assign v_58928 = v_58925 & v_58927;
assign v_58930 = v_58913 & v_58929;
assign v_58932 = v_58423;
assign v_58934 = v_58931 & v_58933;
assign v_58936 = v_58910 & v_58935;
assign v_58938 = v_58419;
assign v_58940 = v_58937 & v_58939;
assign v_58942 = v_58907 & v_58941;
assign v_58944 = v_58415;
assign v_58946 = v_58943 & v_58945;
assign v_58948 = v_58904 & v_58947;
assign v_58950 = v_58411;
assign v_58952 = v_58949 & v_58951;
assign v_58954 = v_58901 & v_58953;
assign v_58956 = v_58407;
assign v_58958 = v_58955 & v_58957;
assign v_58960 = v_58898 & v_58959;
assign v_58962 = v_58403;
assign v_58964 = v_58961 & v_58963;
assign v_58966 = v_58895 & v_58965;
assign v_58968 = v_58399;
assign v_58970 = v_58967 & v_58969;
assign v_58972 = v_58892 & v_58971;
assign v_58974 = v_58395;
assign v_58976 = v_58973 & v_58975;
assign v_58978 = v_58889 & v_58977;
assign v_58980 = v_58391;
assign v_58982 = v_58979 & v_58981;
assign v_58984 = v_58886 & v_58983;
assign v_58986 = v_58387;
assign v_58988 = v_58985 & v_58987;
assign v_58990 = v_58883 & v_58989;
assign v_58992 = v_58383;
assign v_58994 = v_58991 & v_58993;
assign v_58996 = v_58880 & v_58995;
assign v_58998 = v_555;
assign v_59000 = v_58997 & v_58999;
assign v_59002 = v_58877 & v_59001;
assign v_59004 = v_551;
assign v_59006 = v_59003 & v_59005;
assign v_59008 = v_58874 & v_59007;
assign v_59010 = v_547;
assign v_59012 = v_59009 & v_59011;
assign v_59014 = v_58871 & v_59013;
assign v_59016 = v_543;
assign v_59018 = v_59015 & v_59017;
assign v_59019 = v_59018;
assign v_59021 = v_58431;
assign v_59022 = v_608;
assign v_59023 = v_59022;
assign v_59024 = v_59021 & v_59023;
assign v_59025 = v_59024;
assign v_59026 = v_58916 & v_59025;
assign v_59028 = v_58926 & v_59027;
assign v_59029 = v_58915 & v_59025;
assign v_59031 = v_58913 & v_59030;
assign v_59033 = v_58932 & v_59032;
assign v_59034 = v_58912 & v_59030;
assign v_59036 = v_58910 & v_59035;
assign v_59038 = v_58938 & v_59037;
assign v_59039 = v_58909 & v_59035;
assign v_59041 = v_58907 & v_59040;
assign v_59043 = v_58944 & v_59042;
assign v_59044 = v_58906 & v_59040;
assign v_59046 = v_58904 & v_59045;
assign v_59048 = v_58950 & v_59047;
assign v_59049 = v_58903 & v_59045;
assign v_59051 = v_58901 & v_59050;
assign v_59053 = v_58956 & v_59052;
assign v_59054 = v_58900 & v_59050;
assign v_59056 = v_58898 & v_59055;
assign v_59058 = v_58962 & v_59057;
assign v_59059 = v_58897 & v_59055;
assign v_59061 = v_58895 & v_59060;
assign v_59063 = v_58968 & v_59062;
assign v_59064 = v_58894 & v_59060;
assign v_59066 = v_58892 & v_59065;
assign v_59068 = v_58974 & v_59067;
assign v_59069 = v_58891 & v_59065;
assign v_59071 = v_58889 & v_59070;
assign v_59073 = v_58980 & v_59072;
assign v_59074 = v_58888 & v_59070;
assign v_59076 = v_58886 & v_59075;
assign v_59078 = v_58986 & v_59077;
assign v_59079 = v_58885 & v_59075;
assign v_59081 = v_58883 & v_59080;
assign v_59083 = v_58992 & v_59082;
assign v_59084 = v_58882 & v_59080;
assign v_59086 = v_58880 & v_59085;
assign v_59088 = v_58998 & v_59087;
assign v_59089 = v_58879 & v_59085;
assign v_59091 = v_58877 & v_59090;
assign v_59093 = v_59004 & v_59092;
assign v_59094 = v_58876 & v_59090;
assign v_59096 = v_58874 & v_59095;
assign v_59098 = v_59010 & v_59097;
assign v_59099 = v_58873 & v_59095;
assign v_59101 = v_58871 & v_59100;
assign v_59103 = v_59016 & v_59102;
assign v_59104 = v_58870 & v_59100;
assign v_59106 = v_59105;
assign v_59108 = v_59020 & v_59107;
assign v_59109 = v_59108;
assign v_59111 = v_59110;
assign v_59113 = ~v_803;
assign v_59114 = ~v_58368;
assign v_59115 = v_58368;
assign v_59116 = ~v_807;
assign v_59117 = ~v_58372;
assign v_59118 = v_58372;
assign v_59119 = ~v_811;
assign v_59120 = ~v_58376;
assign v_59121 = v_58376;
assign v_59122 = ~v_815;
assign v_59123 = ~v_58380;
assign v_59124 = v_58380;
assign v_59125 = ~v_58383;
assign v_59126 = ~v_820;
assign v_59127 = v_820;
assign v_59128 = ~v_58387;
assign v_59129 = ~v_824;
assign v_59130 = v_824;
assign v_59131 = ~v_58391;
assign v_59132 = ~v_828;
assign v_59133 = v_828;
assign v_59134 = ~v_58395;
assign v_59135 = ~v_832;
assign v_59136 = v_832;
assign v_59137 = ~v_58399;
assign v_59138 = ~v_836;
assign v_59139 = v_836;
assign v_59140 = ~v_58403;
assign v_59141 = ~v_840;
assign v_59142 = v_840;
assign v_59143 = ~v_58407;
assign v_59144 = ~v_844;
assign v_59145 = v_844;
assign v_59146 = ~v_58411;
assign v_59147 = ~v_848;
assign v_59148 = v_848;
assign v_59149 = ~v_58415;
assign v_59150 = ~v_852;
assign v_59151 = v_852;
assign v_59152 = ~v_58419;
assign v_59153 = ~v_856;
assign v_59154 = v_856;
assign v_59155 = ~v_58423;
assign v_59156 = ~v_860;
assign v_59157 = v_860;
assign v_59158 = ~v_58427;
assign v_59159 = ~v_864;
assign v_59160 = v_864;
assign v_59161 = ~v_58431;
assign v_59162 = ~v_868;
assign v_59163 = v_59162;
assign v_59165 = v_59164;
assign v_59167 = v_59159 & v_59166;
assign v_59169 = v_58427;
assign v_59171 = v_59168 & v_59170;
assign v_59173 = v_59156 & v_59172;
assign v_59175 = v_58423;
assign v_59177 = v_59174 & v_59176;
assign v_59179 = v_59153 & v_59178;
assign v_59181 = v_58419;
assign v_59183 = v_59180 & v_59182;
assign v_59185 = v_59150 & v_59184;
assign v_59187 = v_58415;
assign v_59189 = v_59186 & v_59188;
assign v_59191 = v_59147 & v_59190;
assign v_59193 = v_58411;
assign v_59195 = v_59192 & v_59194;
assign v_59197 = v_59144 & v_59196;
assign v_59199 = v_58407;
assign v_59201 = v_59198 & v_59200;
assign v_59203 = v_59141 & v_59202;
assign v_59205 = v_58403;
assign v_59207 = v_59204 & v_59206;
assign v_59209 = v_59138 & v_59208;
assign v_59211 = v_58399;
assign v_59213 = v_59210 & v_59212;
assign v_59215 = v_59135 & v_59214;
assign v_59217 = v_58395;
assign v_59219 = v_59216 & v_59218;
assign v_59221 = v_59132 & v_59220;
assign v_59223 = v_58391;
assign v_59225 = v_59222 & v_59224;
assign v_59227 = v_59129 & v_59226;
assign v_59229 = v_58387;
assign v_59231 = v_59228 & v_59230;
assign v_59233 = v_59126 & v_59232;
assign v_59235 = v_58383;
assign v_59237 = v_59234 & v_59236;
assign v_59239 = v_59123 & v_59238;
assign v_59241 = v_815;
assign v_59243 = v_59240 & v_59242;
assign v_59245 = v_59120 & v_59244;
assign v_59247 = v_811;
assign v_59249 = v_59246 & v_59248;
assign v_59251 = v_59117 & v_59250;
assign v_59253 = v_807;
assign v_59255 = v_59252 & v_59254;
assign v_59257 = v_59114 & v_59256;
assign v_59259 = v_803;
assign v_59261 = v_59258 & v_59260;
assign v_59262 = v_59261;
assign v_59264 = v_58431;
assign v_59265 = v_868;
assign v_59266 = v_59265;
assign v_59267 = v_59264 & v_59266;
assign v_59268 = v_59267;
assign v_59269 = v_59159 & v_59268;
assign v_59271 = v_59169 & v_59270;
assign v_59272 = v_59158 & v_59268;
assign v_59274 = v_59156 & v_59273;
assign v_59276 = v_59175 & v_59275;
assign v_59277 = v_59155 & v_59273;
assign v_59279 = v_59153 & v_59278;
assign v_59281 = v_59181 & v_59280;
assign v_59282 = v_59152 & v_59278;
assign v_59284 = v_59150 & v_59283;
assign v_59286 = v_59187 & v_59285;
assign v_59287 = v_59149 & v_59283;
assign v_59289 = v_59147 & v_59288;
assign v_59291 = v_59193 & v_59290;
assign v_59292 = v_59146 & v_59288;
assign v_59294 = v_59144 & v_59293;
assign v_59296 = v_59199 & v_59295;
assign v_59297 = v_59143 & v_59293;
assign v_59299 = v_59141 & v_59298;
assign v_59301 = v_59205 & v_59300;
assign v_59302 = v_59140 & v_59298;
assign v_59304 = v_59138 & v_59303;
assign v_59306 = v_59211 & v_59305;
assign v_59307 = v_59137 & v_59303;
assign v_59309 = v_59135 & v_59308;
assign v_59311 = v_59217 & v_59310;
assign v_59312 = v_59134 & v_59308;
assign v_59314 = v_59132 & v_59313;
assign v_59316 = v_59223 & v_59315;
assign v_59317 = v_59131 & v_59313;
assign v_59319 = v_59129 & v_59318;
assign v_59321 = v_59229 & v_59320;
assign v_59322 = v_59128 & v_59318;
assign v_59324 = v_59126 & v_59323;
assign v_59326 = v_59235 & v_59325;
assign v_59327 = v_59125 & v_59323;
assign v_59329 = v_59123 & v_59328;
assign v_59331 = v_59241 & v_59330;
assign v_59332 = v_59122 & v_59328;
assign v_59334 = v_59120 & v_59333;
assign v_59336 = v_59247 & v_59335;
assign v_59337 = v_59119 & v_59333;
assign v_59339 = v_59117 & v_59338;
assign v_59341 = v_59253 & v_59340;
assign v_59342 = v_59116 & v_59338;
assign v_59344 = v_59114 & v_59343;
assign v_59346 = v_59259 & v_59345;
assign v_59347 = v_59113 & v_59343;
assign v_59349 = v_59348;
assign v_59351 = v_59263 & v_59350;
assign v_59352 = v_59351;
assign v_59354 = v_59353;
assign v_59356 = ~v_1063;
assign v_59357 = ~v_58368;
assign v_59358 = v_58368;
assign v_59359 = ~v_1067;
assign v_59360 = ~v_58372;
assign v_59361 = v_58372;
assign v_59362 = ~v_1071;
assign v_59363 = ~v_58376;
assign v_59364 = v_58376;
assign v_59365 = ~v_1075;
assign v_59366 = ~v_58380;
assign v_59367 = v_58380;
assign v_59368 = ~v_58383;
assign v_59369 = ~v_1080;
assign v_59370 = v_1080;
assign v_59371 = ~v_58387;
assign v_59372 = ~v_1084;
assign v_59373 = v_1084;
assign v_59374 = ~v_58391;
assign v_59375 = ~v_1088;
assign v_59376 = v_1088;
assign v_59377 = ~v_58395;
assign v_59378 = ~v_1092;
assign v_59379 = v_1092;
assign v_59380 = ~v_58399;
assign v_59381 = ~v_1096;
assign v_59382 = v_1096;
assign v_59383 = ~v_58403;
assign v_59384 = ~v_1100;
assign v_59385 = v_1100;
assign v_59386 = ~v_58407;
assign v_59387 = ~v_1104;
assign v_59388 = v_1104;
assign v_59389 = ~v_58411;
assign v_59390 = ~v_1108;
assign v_59391 = v_1108;
assign v_59392 = ~v_58415;
assign v_59393 = ~v_1112;
assign v_59394 = v_1112;
assign v_59395 = ~v_58419;
assign v_59396 = ~v_1116;
assign v_59397 = v_1116;
assign v_59398 = ~v_58423;
assign v_59399 = ~v_1120;
assign v_59400 = v_1120;
assign v_59401 = ~v_58427;
assign v_59402 = ~v_1124;
assign v_59403 = v_1124;
assign v_59404 = ~v_58431;
assign v_59405 = ~v_1128;
assign v_59406 = v_59405;
assign v_59408 = v_59407;
assign v_59410 = v_59402 & v_59409;
assign v_59412 = v_58427;
assign v_59414 = v_59411 & v_59413;
assign v_59416 = v_59399 & v_59415;
assign v_59418 = v_58423;
assign v_59420 = v_59417 & v_59419;
assign v_59422 = v_59396 & v_59421;
assign v_59424 = v_58419;
assign v_59426 = v_59423 & v_59425;
assign v_59428 = v_59393 & v_59427;
assign v_59430 = v_58415;
assign v_59432 = v_59429 & v_59431;
assign v_59434 = v_59390 & v_59433;
assign v_59436 = v_58411;
assign v_59438 = v_59435 & v_59437;
assign v_59440 = v_59387 & v_59439;
assign v_59442 = v_58407;
assign v_59444 = v_59441 & v_59443;
assign v_59446 = v_59384 & v_59445;
assign v_59448 = v_58403;
assign v_59450 = v_59447 & v_59449;
assign v_59452 = v_59381 & v_59451;
assign v_59454 = v_58399;
assign v_59456 = v_59453 & v_59455;
assign v_59458 = v_59378 & v_59457;
assign v_59460 = v_58395;
assign v_59462 = v_59459 & v_59461;
assign v_59464 = v_59375 & v_59463;
assign v_59466 = v_58391;
assign v_59468 = v_59465 & v_59467;
assign v_59470 = v_59372 & v_59469;
assign v_59472 = v_58387;
assign v_59474 = v_59471 & v_59473;
assign v_59476 = v_59369 & v_59475;
assign v_59478 = v_58383;
assign v_59480 = v_59477 & v_59479;
assign v_59482 = v_59366 & v_59481;
assign v_59484 = v_1075;
assign v_59486 = v_59483 & v_59485;
assign v_59488 = v_59363 & v_59487;
assign v_59490 = v_1071;
assign v_59492 = v_59489 & v_59491;
assign v_59494 = v_59360 & v_59493;
assign v_59496 = v_1067;
assign v_59498 = v_59495 & v_59497;
assign v_59500 = v_59357 & v_59499;
assign v_59502 = v_1063;
assign v_59504 = v_59501 & v_59503;
assign v_59505 = v_59504;
assign v_59507 = v_58431;
assign v_59508 = v_1128;
assign v_59509 = v_59508;
assign v_59510 = v_59507 & v_59509;
assign v_59511 = v_59510;
assign v_59512 = v_59402 & v_59511;
assign v_59514 = v_59412 & v_59513;
assign v_59515 = v_59401 & v_59511;
assign v_59517 = v_59399 & v_59516;
assign v_59519 = v_59418 & v_59518;
assign v_59520 = v_59398 & v_59516;
assign v_59522 = v_59396 & v_59521;
assign v_59524 = v_59424 & v_59523;
assign v_59525 = v_59395 & v_59521;
assign v_59527 = v_59393 & v_59526;
assign v_59529 = v_59430 & v_59528;
assign v_59530 = v_59392 & v_59526;
assign v_59532 = v_59390 & v_59531;
assign v_59534 = v_59436 & v_59533;
assign v_59535 = v_59389 & v_59531;
assign v_59537 = v_59387 & v_59536;
assign v_59539 = v_59442 & v_59538;
assign v_59540 = v_59386 & v_59536;
assign v_59542 = v_59384 & v_59541;
assign v_59544 = v_59448 & v_59543;
assign v_59545 = v_59383 & v_59541;
assign v_59547 = v_59381 & v_59546;
assign v_59549 = v_59454 & v_59548;
assign v_59550 = v_59380 & v_59546;
assign v_59552 = v_59378 & v_59551;
assign v_59554 = v_59460 & v_59553;
assign v_59555 = v_59377 & v_59551;
assign v_59557 = v_59375 & v_59556;
assign v_59559 = v_59466 & v_59558;
assign v_59560 = v_59374 & v_59556;
assign v_59562 = v_59372 & v_59561;
assign v_59564 = v_59472 & v_59563;
assign v_59565 = v_59371 & v_59561;
assign v_59567 = v_59369 & v_59566;
assign v_59569 = v_59478 & v_59568;
assign v_59570 = v_59368 & v_59566;
assign v_59572 = v_59366 & v_59571;
assign v_59574 = v_59484 & v_59573;
assign v_59575 = v_59365 & v_59571;
assign v_59577 = v_59363 & v_59576;
assign v_59579 = v_59490 & v_59578;
assign v_59580 = v_59362 & v_59576;
assign v_59582 = v_59360 & v_59581;
assign v_59584 = v_59496 & v_59583;
assign v_59585 = v_59359 & v_59581;
assign v_59587 = v_59357 & v_59586;
assign v_59589 = v_59502 & v_59588;
assign v_59590 = v_59356 & v_59586;
assign v_59592 = v_59591;
assign v_59594 = v_59506 & v_59593;
assign v_59595 = v_59594;
assign v_59597 = v_59596;
assign v_59599 = ~v_1323;
assign v_59600 = ~v_58368;
assign v_59601 = v_58368;
assign v_59602 = ~v_1327;
assign v_59603 = ~v_58372;
assign v_59604 = v_58372;
assign v_59605 = ~v_1331;
assign v_59606 = ~v_58376;
assign v_59607 = v_58376;
assign v_59608 = ~v_1335;
assign v_59609 = ~v_58380;
assign v_59610 = v_58380;
assign v_59611 = ~v_58383;
assign v_59612 = ~v_1340;
assign v_59613 = v_1340;
assign v_59614 = ~v_58387;
assign v_59615 = ~v_1344;
assign v_59616 = v_1344;
assign v_59617 = ~v_58391;
assign v_59618 = ~v_1348;
assign v_59619 = v_1348;
assign v_59620 = ~v_58395;
assign v_59621 = ~v_1352;
assign v_59622 = v_1352;
assign v_59623 = ~v_58399;
assign v_59624 = ~v_1356;
assign v_59625 = v_1356;
assign v_59626 = ~v_58403;
assign v_59627 = ~v_1360;
assign v_59628 = v_1360;
assign v_59629 = ~v_58407;
assign v_59630 = ~v_1364;
assign v_59631 = v_1364;
assign v_59632 = ~v_58411;
assign v_59633 = ~v_1368;
assign v_59634 = v_1368;
assign v_59635 = ~v_58415;
assign v_59636 = ~v_1372;
assign v_59637 = v_1372;
assign v_59638 = ~v_58419;
assign v_59639 = ~v_1376;
assign v_59640 = v_1376;
assign v_59641 = ~v_58423;
assign v_59642 = ~v_1380;
assign v_59643 = v_1380;
assign v_59644 = ~v_58427;
assign v_59645 = ~v_1384;
assign v_59646 = v_1384;
assign v_59647 = ~v_58431;
assign v_59648 = ~v_1388;
assign v_59649 = v_59648;
assign v_59651 = v_59650;
assign v_59653 = v_59645 & v_59652;
assign v_59655 = v_58427;
assign v_59657 = v_59654 & v_59656;
assign v_59659 = v_59642 & v_59658;
assign v_59661 = v_58423;
assign v_59663 = v_59660 & v_59662;
assign v_59665 = v_59639 & v_59664;
assign v_59667 = v_58419;
assign v_59669 = v_59666 & v_59668;
assign v_59671 = v_59636 & v_59670;
assign v_59673 = v_58415;
assign v_59675 = v_59672 & v_59674;
assign v_59677 = v_59633 & v_59676;
assign v_59679 = v_58411;
assign v_59681 = v_59678 & v_59680;
assign v_59683 = v_59630 & v_59682;
assign v_59685 = v_58407;
assign v_59687 = v_59684 & v_59686;
assign v_59689 = v_59627 & v_59688;
assign v_59691 = v_58403;
assign v_59693 = v_59690 & v_59692;
assign v_59695 = v_59624 & v_59694;
assign v_59697 = v_58399;
assign v_59699 = v_59696 & v_59698;
assign v_59701 = v_59621 & v_59700;
assign v_59703 = v_58395;
assign v_59705 = v_59702 & v_59704;
assign v_59707 = v_59618 & v_59706;
assign v_59709 = v_58391;
assign v_59711 = v_59708 & v_59710;
assign v_59713 = v_59615 & v_59712;
assign v_59715 = v_58387;
assign v_59717 = v_59714 & v_59716;
assign v_59719 = v_59612 & v_59718;
assign v_59721 = v_58383;
assign v_59723 = v_59720 & v_59722;
assign v_59725 = v_59609 & v_59724;
assign v_59727 = v_1335;
assign v_59729 = v_59726 & v_59728;
assign v_59731 = v_59606 & v_59730;
assign v_59733 = v_1331;
assign v_59735 = v_59732 & v_59734;
assign v_59737 = v_59603 & v_59736;
assign v_59739 = v_1327;
assign v_59741 = v_59738 & v_59740;
assign v_59743 = v_59600 & v_59742;
assign v_59745 = v_1323;
assign v_59747 = v_59744 & v_59746;
assign v_59748 = v_59747;
assign v_59750 = v_58431;
assign v_59751 = v_1388;
assign v_59752 = v_59751;
assign v_59753 = v_59750 & v_59752;
assign v_59754 = v_59753;
assign v_59755 = v_59645 & v_59754;
assign v_59757 = v_59655 & v_59756;
assign v_59758 = v_59644 & v_59754;
assign v_59760 = v_59642 & v_59759;
assign v_59762 = v_59661 & v_59761;
assign v_59763 = v_59641 & v_59759;
assign v_59765 = v_59639 & v_59764;
assign v_59767 = v_59667 & v_59766;
assign v_59768 = v_59638 & v_59764;
assign v_59770 = v_59636 & v_59769;
assign v_59772 = v_59673 & v_59771;
assign v_59773 = v_59635 & v_59769;
assign v_59775 = v_59633 & v_59774;
assign v_59777 = v_59679 & v_59776;
assign v_59778 = v_59632 & v_59774;
assign v_59780 = v_59630 & v_59779;
assign v_59782 = v_59685 & v_59781;
assign v_59783 = v_59629 & v_59779;
assign v_59785 = v_59627 & v_59784;
assign v_59787 = v_59691 & v_59786;
assign v_59788 = v_59626 & v_59784;
assign v_59790 = v_59624 & v_59789;
assign v_59792 = v_59697 & v_59791;
assign v_59793 = v_59623 & v_59789;
assign v_59795 = v_59621 & v_59794;
assign v_59797 = v_59703 & v_59796;
assign v_59798 = v_59620 & v_59794;
assign v_59800 = v_59618 & v_59799;
assign v_59802 = v_59709 & v_59801;
assign v_59803 = v_59617 & v_59799;
assign v_59805 = v_59615 & v_59804;
assign v_59807 = v_59715 & v_59806;
assign v_59808 = v_59614 & v_59804;
assign v_59810 = v_59612 & v_59809;
assign v_59812 = v_59721 & v_59811;
assign v_59813 = v_59611 & v_59809;
assign v_59815 = v_59609 & v_59814;
assign v_59817 = v_59727 & v_59816;
assign v_59818 = v_59608 & v_59814;
assign v_59820 = v_59606 & v_59819;
assign v_59822 = v_59733 & v_59821;
assign v_59823 = v_59605 & v_59819;
assign v_59825 = v_59603 & v_59824;
assign v_59827 = v_59739 & v_59826;
assign v_59828 = v_59602 & v_59824;
assign v_59830 = v_59600 & v_59829;
assign v_59832 = v_59745 & v_59831;
assign v_59833 = v_59599 & v_59829;
assign v_59835 = v_59834;
assign v_59837 = v_59749 & v_59836;
assign v_59838 = v_59837;
assign v_59840 = v_59839;
assign v_59842 = ~v_1583;
assign v_59843 = ~v_58368;
assign v_59844 = v_58368;
assign v_59845 = ~v_1587;
assign v_59846 = ~v_58372;
assign v_59847 = v_58372;
assign v_59848 = ~v_1591;
assign v_59849 = ~v_58376;
assign v_59850 = v_58376;
assign v_59851 = ~v_1595;
assign v_59852 = ~v_58380;
assign v_59853 = v_58380;
assign v_59854 = ~v_58383;
assign v_59855 = ~v_1600;
assign v_59856 = v_1600;
assign v_59857 = ~v_58387;
assign v_59858 = ~v_1604;
assign v_59859 = v_1604;
assign v_59860 = ~v_58391;
assign v_59861 = ~v_1608;
assign v_59862 = v_1608;
assign v_59863 = ~v_58395;
assign v_59864 = ~v_1612;
assign v_59865 = v_1612;
assign v_59866 = ~v_58399;
assign v_59867 = ~v_1616;
assign v_59868 = v_1616;
assign v_59869 = ~v_58403;
assign v_59870 = ~v_1620;
assign v_59871 = v_1620;
assign v_59872 = ~v_58407;
assign v_59873 = ~v_1624;
assign v_59874 = v_1624;
assign v_59875 = ~v_58411;
assign v_59876 = ~v_1628;
assign v_59877 = v_1628;
assign v_59878 = ~v_58415;
assign v_59879 = ~v_1632;
assign v_59880 = v_1632;
assign v_59881 = ~v_58419;
assign v_59882 = ~v_1636;
assign v_59883 = v_1636;
assign v_59884 = ~v_58423;
assign v_59885 = ~v_1640;
assign v_59886 = v_1640;
assign v_59887 = ~v_58427;
assign v_59888 = ~v_1644;
assign v_59889 = v_1644;
assign v_59890 = ~v_58431;
assign v_59891 = ~v_1648;
assign v_59892 = v_59891;
assign v_59894 = v_59893;
assign v_59896 = v_59888 & v_59895;
assign v_59898 = v_58427;
assign v_59900 = v_59897 & v_59899;
assign v_59902 = v_59885 & v_59901;
assign v_59904 = v_58423;
assign v_59906 = v_59903 & v_59905;
assign v_59908 = v_59882 & v_59907;
assign v_59910 = v_58419;
assign v_59912 = v_59909 & v_59911;
assign v_59914 = v_59879 & v_59913;
assign v_59916 = v_58415;
assign v_59918 = v_59915 & v_59917;
assign v_59920 = v_59876 & v_59919;
assign v_59922 = v_58411;
assign v_59924 = v_59921 & v_59923;
assign v_59926 = v_59873 & v_59925;
assign v_59928 = v_58407;
assign v_59930 = v_59927 & v_59929;
assign v_59932 = v_59870 & v_59931;
assign v_59934 = v_58403;
assign v_59936 = v_59933 & v_59935;
assign v_59938 = v_59867 & v_59937;
assign v_59940 = v_58399;
assign v_59942 = v_59939 & v_59941;
assign v_59944 = v_59864 & v_59943;
assign v_59946 = v_58395;
assign v_59948 = v_59945 & v_59947;
assign v_59950 = v_59861 & v_59949;
assign v_59952 = v_58391;
assign v_59954 = v_59951 & v_59953;
assign v_59956 = v_59858 & v_59955;
assign v_59958 = v_58387;
assign v_59960 = v_59957 & v_59959;
assign v_59962 = v_59855 & v_59961;
assign v_59964 = v_58383;
assign v_59966 = v_59963 & v_59965;
assign v_59968 = v_59852 & v_59967;
assign v_59970 = v_1595;
assign v_59972 = v_59969 & v_59971;
assign v_59974 = v_59849 & v_59973;
assign v_59976 = v_1591;
assign v_59978 = v_59975 & v_59977;
assign v_59980 = v_59846 & v_59979;
assign v_59982 = v_1587;
assign v_59984 = v_59981 & v_59983;
assign v_59986 = v_59843 & v_59985;
assign v_59988 = v_1583;
assign v_59990 = v_59987 & v_59989;
assign v_59991 = v_59990;
assign v_59993 = v_58431;
assign v_59994 = v_1648;
assign v_59995 = v_59994;
assign v_59996 = v_59993 & v_59995;
assign v_59997 = v_59996;
assign v_59998 = v_59888 & v_59997;
assign v_60000 = v_59898 & v_59999;
assign v_60001 = v_59887 & v_59997;
assign v_60003 = v_59885 & v_60002;
assign v_60005 = v_59904 & v_60004;
assign v_60006 = v_59884 & v_60002;
assign v_60008 = v_59882 & v_60007;
assign v_60010 = v_59910 & v_60009;
assign v_60011 = v_59881 & v_60007;
assign v_60013 = v_59879 & v_60012;
assign v_60015 = v_59916 & v_60014;
assign v_60016 = v_59878 & v_60012;
assign v_60018 = v_59876 & v_60017;
assign v_60020 = v_59922 & v_60019;
assign v_60021 = v_59875 & v_60017;
assign v_60023 = v_59873 & v_60022;
assign v_60025 = v_59928 & v_60024;
assign v_60026 = v_59872 & v_60022;
assign v_60028 = v_59870 & v_60027;
assign v_60030 = v_59934 & v_60029;
assign v_60031 = v_59869 & v_60027;
assign v_60033 = v_59867 & v_60032;
assign v_60035 = v_59940 & v_60034;
assign v_60036 = v_59866 & v_60032;
assign v_60038 = v_59864 & v_60037;
assign v_60040 = v_59946 & v_60039;
assign v_60041 = v_59863 & v_60037;
assign v_60043 = v_59861 & v_60042;
assign v_60045 = v_59952 & v_60044;
assign v_60046 = v_59860 & v_60042;
assign v_60048 = v_59858 & v_60047;
assign v_60050 = v_59958 & v_60049;
assign v_60051 = v_59857 & v_60047;
assign v_60053 = v_59855 & v_60052;
assign v_60055 = v_59964 & v_60054;
assign v_60056 = v_59854 & v_60052;
assign v_60058 = v_59852 & v_60057;
assign v_60060 = v_59970 & v_60059;
assign v_60061 = v_59851 & v_60057;
assign v_60063 = v_59849 & v_60062;
assign v_60065 = v_59976 & v_60064;
assign v_60066 = v_59848 & v_60062;
assign v_60068 = v_59846 & v_60067;
assign v_60070 = v_59982 & v_60069;
assign v_60071 = v_59845 & v_60067;
assign v_60073 = v_59843 & v_60072;
assign v_60075 = v_59988 & v_60074;
assign v_60076 = v_59842 & v_60072;
assign v_60078 = v_60077;
assign v_60080 = v_59992 & v_60079;
assign v_60081 = v_60080;
assign v_60083 = v_60082;
assign v_60085 = ~v_1843;
assign v_60086 = ~v_58368;
assign v_60087 = v_58368;
assign v_60088 = ~v_1847;
assign v_60089 = ~v_58372;
assign v_60090 = v_58372;
assign v_60091 = ~v_1851;
assign v_60092 = ~v_58376;
assign v_60093 = v_58376;
assign v_60094 = ~v_1855;
assign v_60095 = ~v_58380;
assign v_60096 = v_58380;
assign v_60097 = ~v_58383;
assign v_60098 = ~v_1860;
assign v_60099 = v_1860;
assign v_60100 = ~v_58387;
assign v_60101 = ~v_1864;
assign v_60102 = v_1864;
assign v_60103 = ~v_58391;
assign v_60104 = ~v_1868;
assign v_60105 = v_1868;
assign v_60106 = ~v_58395;
assign v_60107 = ~v_1872;
assign v_60108 = v_1872;
assign v_60109 = ~v_58399;
assign v_60110 = ~v_1876;
assign v_60111 = v_1876;
assign v_60112 = ~v_58403;
assign v_60113 = ~v_1880;
assign v_60114 = v_1880;
assign v_60115 = ~v_58407;
assign v_60116 = ~v_1884;
assign v_60117 = v_1884;
assign v_60118 = ~v_58411;
assign v_60119 = ~v_1888;
assign v_60120 = v_1888;
assign v_60121 = ~v_58415;
assign v_60122 = ~v_1892;
assign v_60123 = v_1892;
assign v_60124 = ~v_58419;
assign v_60125 = ~v_1896;
assign v_60126 = v_1896;
assign v_60127 = ~v_58423;
assign v_60128 = ~v_1900;
assign v_60129 = v_1900;
assign v_60130 = ~v_58427;
assign v_60131 = ~v_1904;
assign v_60132 = v_1904;
assign v_60133 = ~v_58431;
assign v_60134 = ~v_1908;
assign v_60135 = v_60134;
assign v_60137 = v_60136;
assign v_60139 = v_60131 & v_60138;
assign v_60141 = v_58427;
assign v_60143 = v_60140 & v_60142;
assign v_60145 = v_60128 & v_60144;
assign v_60147 = v_58423;
assign v_60149 = v_60146 & v_60148;
assign v_60151 = v_60125 & v_60150;
assign v_60153 = v_58419;
assign v_60155 = v_60152 & v_60154;
assign v_60157 = v_60122 & v_60156;
assign v_60159 = v_58415;
assign v_60161 = v_60158 & v_60160;
assign v_60163 = v_60119 & v_60162;
assign v_60165 = v_58411;
assign v_60167 = v_60164 & v_60166;
assign v_60169 = v_60116 & v_60168;
assign v_60171 = v_58407;
assign v_60173 = v_60170 & v_60172;
assign v_60175 = v_60113 & v_60174;
assign v_60177 = v_58403;
assign v_60179 = v_60176 & v_60178;
assign v_60181 = v_60110 & v_60180;
assign v_60183 = v_58399;
assign v_60185 = v_60182 & v_60184;
assign v_60187 = v_60107 & v_60186;
assign v_60189 = v_58395;
assign v_60191 = v_60188 & v_60190;
assign v_60193 = v_60104 & v_60192;
assign v_60195 = v_58391;
assign v_60197 = v_60194 & v_60196;
assign v_60199 = v_60101 & v_60198;
assign v_60201 = v_58387;
assign v_60203 = v_60200 & v_60202;
assign v_60205 = v_60098 & v_60204;
assign v_60207 = v_58383;
assign v_60209 = v_60206 & v_60208;
assign v_60211 = v_60095 & v_60210;
assign v_60213 = v_1855;
assign v_60215 = v_60212 & v_60214;
assign v_60217 = v_60092 & v_60216;
assign v_60219 = v_1851;
assign v_60221 = v_60218 & v_60220;
assign v_60223 = v_60089 & v_60222;
assign v_60225 = v_1847;
assign v_60227 = v_60224 & v_60226;
assign v_60229 = v_60086 & v_60228;
assign v_60231 = v_1843;
assign v_60233 = v_60230 & v_60232;
assign v_60234 = v_60233;
assign v_60236 = v_58431;
assign v_60237 = v_1908;
assign v_60238 = v_60237;
assign v_60239 = v_60236 & v_60238;
assign v_60240 = v_60239;
assign v_60241 = v_60131 & v_60240;
assign v_60243 = v_60141 & v_60242;
assign v_60244 = v_60130 & v_60240;
assign v_60246 = v_60128 & v_60245;
assign v_60248 = v_60147 & v_60247;
assign v_60249 = v_60127 & v_60245;
assign v_60251 = v_60125 & v_60250;
assign v_60253 = v_60153 & v_60252;
assign v_60254 = v_60124 & v_60250;
assign v_60256 = v_60122 & v_60255;
assign v_60258 = v_60159 & v_60257;
assign v_60259 = v_60121 & v_60255;
assign v_60261 = v_60119 & v_60260;
assign v_60263 = v_60165 & v_60262;
assign v_60264 = v_60118 & v_60260;
assign v_60266 = v_60116 & v_60265;
assign v_60268 = v_60171 & v_60267;
assign v_60269 = v_60115 & v_60265;
assign v_60271 = v_60113 & v_60270;
assign v_60273 = v_60177 & v_60272;
assign v_60274 = v_60112 & v_60270;
assign v_60276 = v_60110 & v_60275;
assign v_60278 = v_60183 & v_60277;
assign v_60279 = v_60109 & v_60275;
assign v_60281 = v_60107 & v_60280;
assign v_60283 = v_60189 & v_60282;
assign v_60284 = v_60106 & v_60280;
assign v_60286 = v_60104 & v_60285;
assign v_60288 = v_60195 & v_60287;
assign v_60289 = v_60103 & v_60285;
assign v_60291 = v_60101 & v_60290;
assign v_60293 = v_60201 & v_60292;
assign v_60294 = v_60100 & v_60290;
assign v_60296 = v_60098 & v_60295;
assign v_60298 = v_60207 & v_60297;
assign v_60299 = v_60097 & v_60295;
assign v_60301 = v_60095 & v_60300;
assign v_60303 = v_60213 & v_60302;
assign v_60304 = v_60094 & v_60300;
assign v_60306 = v_60092 & v_60305;
assign v_60308 = v_60219 & v_60307;
assign v_60309 = v_60091 & v_60305;
assign v_60311 = v_60089 & v_60310;
assign v_60313 = v_60225 & v_60312;
assign v_60314 = v_60088 & v_60310;
assign v_60316 = v_60086 & v_60315;
assign v_60318 = v_60231 & v_60317;
assign v_60319 = v_60085 & v_60315;
assign v_60321 = v_60320;
assign v_60323 = v_60235 & v_60322;
assign v_60324 = v_60323;
assign v_60326 = v_60325;
assign v_60328 = ~v_2103;
assign v_60329 = ~v_58368;
assign v_60330 = v_58368;
assign v_60331 = ~v_2107;
assign v_60332 = ~v_58372;
assign v_60333 = v_58372;
assign v_60334 = ~v_2111;
assign v_60335 = ~v_58376;
assign v_60336 = v_58376;
assign v_60337 = ~v_2115;
assign v_60338 = ~v_58380;
assign v_60339 = v_58380;
assign v_60340 = ~v_58383;
assign v_60341 = ~v_2120;
assign v_60342 = v_2120;
assign v_60343 = ~v_58387;
assign v_60344 = ~v_2124;
assign v_60345 = v_2124;
assign v_60346 = ~v_58391;
assign v_60347 = ~v_2128;
assign v_60348 = v_2128;
assign v_60349 = ~v_58395;
assign v_60350 = ~v_2132;
assign v_60351 = v_2132;
assign v_60352 = ~v_58399;
assign v_60353 = ~v_2136;
assign v_60354 = v_2136;
assign v_60355 = ~v_58403;
assign v_60356 = ~v_2140;
assign v_60357 = v_2140;
assign v_60358 = ~v_58407;
assign v_60359 = ~v_2144;
assign v_60360 = v_2144;
assign v_60361 = ~v_58411;
assign v_60362 = ~v_2148;
assign v_60363 = v_2148;
assign v_60364 = ~v_58415;
assign v_60365 = ~v_2152;
assign v_60366 = v_2152;
assign v_60367 = ~v_58419;
assign v_60368 = ~v_2156;
assign v_60369 = v_2156;
assign v_60370 = ~v_58423;
assign v_60371 = ~v_2160;
assign v_60372 = v_2160;
assign v_60373 = ~v_58427;
assign v_60374 = ~v_2164;
assign v_60375 = v_2164;
assign v_60376 = ~v_58431;
assign v_60377 = ~v_2168;
assign v_60378 = v_60377;
assign v_60380 = v_60379;
assign v_60382 = v_60374 & v_60381;
assign v_60384 = v_58427;
assign v_60386 = v_60383 & v_60385;
assign v_60388 = v_60371 & v_60387;
assign v_60390 = v_58423;
assign v_60392 = v_60389 & v_60391;
assign v_60394 = v_60368 & v_60393;
assign v_60396 = v_58419;
assign v_60398 = v_60395 & v_60397;
assign v_60400 = v_60365 & v_60399;
assign v_60402 = v_58415;
assign v_60404 = v_60401 & v_60403;
assign v_60406 = v_60362 & v_60405;
assign v_60408 = v_58411;
assign v_60410 = v_60407 & v_60409;
assign v_60412 = v_60359 & v_60411;
assign v_60414 = v_58407;
assign v_60416 = v_60413 & v_60415;
assign v_60418 = v_60356 & v_60417;
assign v_60420 = v_58403;
assign v_60422 = v_60419 & v_60421;
assign v_60424 = v_60353 & v_60423;
assign v_60426 = v_58399;
assign v_60428 = v_60425 & v_60427;
assign v_60430 = v_60350 & v_60429;
assign v_60432 = v_58395;
assign v_60434 = v_60431 & v_60433;
assign v_60436 = v_60347 & v_60435;
assign v_60438 = v_58391;
assign v_60440 = v_60437 & v_60439;
assign v_60442 = v_60344 & v_60441;
assign v_60444 = v_58387;
assign v_60446 = v_60443 & v_60445;
assign v_60448 = v_60341 & v_60447;
assign v_60450 = v_58383;
assign v_60452 = v_60449 & v_60451;
assign v_60454 = v_60338 & v_60453;
assign v_60456 = v_2115;
assign v_60458 = v_60455 & v_60457;
assign v_60460 = v_60335 & v_60459;
assign v_60462 = v_2111;
assign v_60464 = v_60461 & v_60463;
assign v_60466 = v_60332 & v_60465;
assign v_60468 = v_2107;
assign v_60470 = v_60467 & v_60469;
assign v_60472 = v_60329 & v_60471;
assign v_60474 = v_2103;
assign v_60476 = v_60473 & v_60475;
assign v_60477 = v_60476;
assign v_60479 = v_58431;
assign v_60480 = v_2168;
assign v_60481 = v_60480;
assign v_60482 = v_60479 & v_60481;
assign v_60483 = v_60482;
assign v_60484 = v_60374 & v_60483;
assign v_60486 = v_60384 & v_60485;
assign v_60487 = v_60373 & v_60483;
assign v_60489 = v_60371 & v_60488;
assign v_60491 = v_60390 & v_60490;
assign v_60492 = v_60370 & v_60488;
assign v_60494 = v_60368 & v_60493;
assign v_60496 = v_60396 & v_60495;
assign v_60497 = v_60367 & v_60493;
assign v_60499 = v_60365 & v_60498;
assign v_60501 = v_60402 & v_60500;
assign v_60502 = v_60364 & v_60498;
assign v_60504 = v_60362 & v_60503;
assign v_60506 = v_60408 & v_60505;
assign v_60507 = v_60361 & v_60503;
assign v_60509 = v_60359 & v_60508;
assign v_60511 = v_60414 & v_60510;
assign v_60512 = v_60358 & v_60508;
assign v_60514 = v_60356 & v_60513;
assign v_60516 = v_60420 & v_60515;
assign v_60517 = v_60355 & v_60513;
assign v_60519 = v_60353 & v_60518;
assign v_60521 = v_60426 & v_60520;
assign v_60522 = v_60352 & v_60518;
assign v_60524 = v_60350 & v_60523;
assign v_60526 = v_60432 & v_60525;
assign v_60527 = v_60349 & v_60523;
assign v_60529 = v_60347 & v_60528;
assign v_60531 = v_60438 & v_60530;
assign v_60532 = v_60346 & v_60528;
assign v_60534 = v_60344 & v_60533;
assign v_60536 = v_60444 & v_60535;
assign v_60537 = v_60343 & v_60533;
assign v_60539 = v_60341 & v_60538;
assign v_60541 = v_60450 & v_60540;
assign v_60542 = v_60340 & v_60538;
assign v_60544 = v_60338 & v_60543;
assign v_60546 = v_60456 & v_60545;
assign v_60547 = v_60337 & v_60543;
assign v_60549 = v_60335 & v_60548;
assign v_60551 = v_60462 & v_60550;
assign v_60552 = v_60334 & v_60548;
assign v_60554 = v_60332 & v_60553;
assign v_60556 = v_60468 & v_60555;
assign v_60557 = v_60331 & v_60553;
assign v_60559 = v_60329 & v_60558;
assign v_60561 = v_60474 & v_60560;
assign v_60562 = v_60328 & v_60558;
assign v_60564 = v_60563;
assign v_60566 = v_60478 & v_60565;
assign v_60567 = v_60566;
assign v_60569 = v_60568;
assign v_60571 = ~v_2363;
assign v_60572 = ~v_58368;
assign v_60573 = v_58368;
assign v_60574 = ~v_2367;
assign v_60575 = ~v_58372;
assign v_60576 = v_58372;
assign v_60577 = ~v_2371;
assign v_60578 = ~v_58376;
assign v_60579 = v_58376;
assign v_60580 = ~v_2375;
assign v_60581 = ~v_58380;
assign v_60582 = v_58380;
assign v_60583 = ~v_58383;
assign v_60584 = ~v_2380;
assign v_60585 = v_2380;
assign v_60586 = ~v_58387;
assign v_60587 = ~v_2384;
assign v_60588 = v_2384;
assign v_60589 = ~v_58391;
assign v_60590 = ~v_2388;
assign v_60591 = v_2388;
assign v_60592 = ~v_58395;
assign v_60593 = ~v_2392;
assign v_60594 = v_2392;
assign v_60595 = ~v_58399;
assign v_60596 = ~v_2396;
assign v_60597 = v_2396;
assign v_60598 = ~v_58403;
assign v_60599 = ~v_2400;
assign v_60600 = v_2400;
assign v_60601 = ~v_58407;
assign v_60602 = ~v_2404;
assign v_60603 = v_2404;
assign v_60604 = ~v_58411;
assign v_60605 = ~v_2408;
assign v_60606 = v_2408;
assign v_60607 = ~v_58415;
assign v_60608 = ~v_2412;
assign v_60609 = v_2412;
assign v_60610 = ~v_58419;
assign v_60611 = ~v_2416;
assign v_60612 = v_2416;
assign v_60613 = ~v_58423;
assign v_60614 = ~v_2420;
assign v_60615 = v_2420;
assign v_60616 = ~v_58427;
assign v_60617 = ~v_2424;
assign v_60618 = v_2424;
assign v_60619 = ~v_58431;
assign v_60620 = ~v_2428;
assign v_60621 = v_60620;
assign v_60623 = v_60622;
assign v_60625 = v_60617 & v_60624;
assign v_60627 = v_58427;
assign v_60629 = v_60626 & v_60628;
assign v_60631 = v_60614 & v_60630;
assign v_60633 = v_58423;
assign v_60635 = v_60632 & v_60634;
assign v_60637 = v_60611 & v_60636;
assign v_60639 = v_58419;
assign v_60641 = v_60638 & v_60640;
assign v_60643 = v_60608 & v_60642;
assign v_60645 = v_58415;
assign v_60647 = v_60644 & v_60646;
assign v_60649 = v_60605 & v_60648;
assign v_60651 = v_58411;
assign v_60653 = v_60650 & v_60652;
assign v_60655 = v_60602 & v_60654;
assign v_60657 = v_58407;
assign v_60659 = v_60656 & v_60658;
assign v_60661 = v_60599 & v_60660;
assign v_60663 = v_58403;
assign v_60665 = v_60662 & v_60664;
assign v_60667 = v_60596 & v_60666;
assign v_60669 = v_58399;
assign v_60671 = v_60668 & v_60670;
assign v_60673 = v_60593 & v_60672;
assign v_60675 = v_58395;
assign v_60677 = v_60674 & v_60676;
assign v_60679 = v_60590 & v_60678;
assign v_60681 = v_58391;
assign v_60683 = v_60680 & v_60682;
assign v_60685 = v_60587 & v_60684;
assign v_60687 = v_58387;
assign v_60689 = v_60686 & v_60688;
assign v_60691 = v_60584 & v_60690;
assign v_60693 = v_58383;
assign v_60695 = v_60692 & v_60694;
assign v_60697 = v_60581 & v_60696;
assign v_60699 = v_2375;
assign v_60701 = v_60698 & v_60700;
assign v_60703 = v_60578 & v_60702;
assign v_60705 = v_2371;
assign v_60707 = v_60704 & v_60706;
assign v_60709 = v_60575 & v_60708;
assign v_60711 = v_2367;
assign v_60713 = v_60710 & v_60712;
assign v_60715 = v_60572 & v_60714;
assign v_60717 = v_2363;
assign v_60719 = v_60716 & v_60718;
assign v_60720 = v_60719;
assign v_60722 = v_58431;
assign v_60723 = v_2428;
assign v_60724 = v_60723;
assign v_60725 = v_60722 & v_60724;
assign v_60726 = v_60725;
assign v_60727 = v_60617 & v_60726;
assign v_60729 = v_60627 & v_60728;
assign v_60730 = v_60616 & v_60726;
assign v_60732 = v_60614 & v_60731;
assign v_60734 = v_60633 & v_60733;
assign v_60735 = v_60613 & v_60731;
assign v_60737 = v_60611 & v_60736;
assign v_60739 = v_60639 & v_60738;
assign v_60740 = v_60610 & v_60736;
assign v_60742 = v_60608 & v_60741;
assign v_60744 = v_60645 & v_60743;
assign v_60745 = v_60607 & v_60741;
assign v_60747 = v_60605 & v_60746;
assign v_60749 = v_60651 & v_60748;
assign v_60750 = v_60604 & v_60746;
assign v_60752 = v_60602 & v_60751;
assign v_60754 = v_60657 & v_60753;
assign v_60755 = v_60601 & v_60751;
assign v_60757 = v_60599 & v_60756;
assign v_60759 = v_60663 & v_60758;
assign v_60760 = v_60598 & v_60756;
assign v_60762 = v_60596 & v_60761;
assign v_60764 = v_60669 & v_60763;
assign v_60765 = v_60595 & v_60761;
assign v_60767 = v_60593 & v_60766;
assign v_60769 = v_60675 & v_60768;
assign v_60770 = v_60592 & v_60766;
assign v_60772 = v_60590 & v_60771;
assign v_60774 = v_60681 & v_60773;
assign v_60775 = v_60589 & v_60771;
assign v_60777 = v_60587 & v_60776;
assign v_60779 = v_60687 & v_60778;
assign v_60780 = v_60586 & v_60776;
assign v_60782 = v_60584 & v_60781;
assign v_60784 = v_60693 & v_60783;
assign v_60785 = v_60583 & v_60781;
assign v_60787 = v_60581 & v_60786;
assign v_60789 = v_60699 & v_60788;
assign v_60790 = v_60580 & v_60786;
assign v_60792 = v_60578 & v_60791;
assign v_60794 = v_60705 & v_60793;
assign v_60795 = v_60577 & v_60791;
assign v_60797 = v_60575 & v_60796;
assign v_60799 = v_60711 & v_60798;
assign v_60800 = v_60574 & v_60796;
assign v_60802 = v_60572 & v_60801;
assign v_60804 = v_60717 & v_60803;
assign v_60805 = v_60571 & v_60801;
assign v_60807 = v_60806;
assign v_60809 = v_60721 & v_60808;
assign v_60810 = v_60809;
assign v_60812 = v_60811;
assign v_60814 = ~v_2623;
assign v_60815 = ~v_58368;
assign v_60816 = v_58368;
assign v_60817 = ~v_2627;
assign v_60818 = ~v_58372;
assign v_60819 = v_58372;
assign v_60820 = ~v_2631;
assign v_60821 = ~v_58376;
assign v_60822 = v_58376;
assign v_60823 = ~v_2635;
assign v_60824 = ~v_58380;
assign v_60825 = v_58380;
assign v_60826 = ~v_58383;
assign v_60827 = ~v_2640;
assign v_60828 = v_2640;
assign v_60829 = ~v_58387;
assign v_60830 = ~v_2644;
assign v_60831 = v_2644;
assign v_60832 = ~v_58391;
assign v_60833 = ~v_2648;
assign v_60834 = v_2648;
assign v_60835 = ~v_58395;
assign v_60836 = ~v_2652;
assign v_60837 = v_2652;
assign v_60838 = ~v_58399;
assign v_60839 = ~v_2656;
assign v_60840 = v_2656;
assign v_60841 = ~v_58403;
assign v_60842 = ~v_2660;
assign v_60843 = v_2660;
assign v_60844 = ~v_58407;
assign v_60845 = ~v_2664;
assign v_60846 = v_2664;
assign v_60847 = ~v_58411;
assign v_60848 = ~v_2668;
assign v_60849 = v_2668;
assign v_60850 = ~v_58415;
assign v_60851 = ~v_2672;
assign v_60852 = v_2672;
assign v_60853 = ~v_58419;
assign v_60854 = ~v_2676;
assign v_60855 = v_2676;
assign v_60856 = ~v_58423;
assign v_60857 = ~v_2680;
assign v_60858 = v_2680;
assign v_60859 = ~v_58427;
assign v_60860 = ~v_2684;
assign v_60861 = v_2684;
assign v_60862 = ~v_58431;
assign v_60863 = ~v_2688;
assign v_60864 = v_60863;
assign v_60866 = v_60865;
assign v_60868 = v_60860 & v_60867;
assign v_60870 = v_58427;
assign v_60872 = v_60869 & v_60871;
assign v_60874 = v_60857 & v_60873;
assign v_60876 = v_58423;
assign v_60878 = v_60875 & v_60877;
assign v_60880 = v_60854 & v_60879;
assign v_60882 = v_58419;
assign v_60884 = v_60881 & v_60883;
assign v_60886 = v_60851 & v_60885;
assign v_60888 = v_58415;
assign v_60890 = v_60887 & v_60889;
assign v_60892 = v_60848 & v_60891;
assign v_60894 = v_58411;
assign v_60896 = v_60893 & v_60895;
assign v_60898 = v_60845 & v_60897;
assign v_60900 = v_58407;
assign v_60902 = v_60899 & v_60901;
assign v_60904 = v_60842 & v_60903;
assign v_60906 = v_58403;
assign v_60908 = v_60905 & v_60907;
assign v_60910 = v_60839 & v_60909;
assign v_60912 = v_58399;
assign v_60914 = v_60911 & v_60913;
assign v_60916 = v_60836 & v_60915;
assign v_60918 = v_58395;
assign v_60920 = v_60917 & v_60919;
assign v_60922 = v_60833 & v_60921;
assign v_60924 = v_58391;
assign v_60926 = v_60923 & v_60925;
assign v_60928 = v_60830 & v_60927;
assign v_60930 = v_58387;
assign v_60932 = v_60929 & v_60931;
assign v_60934 = v_60827 & v_60933;
assign v_60936 = v_58383;
assign v_60938 = v_60935 & v_60937;
assign v_60940 = v_60824 & v_60939;
assign v_60942 = v_2635;
assign v_60944 = v_60941 & v_60943;
assign v_60946 = v_60821 & v_60945;
assign v_60948 = v_2631;
assign v_60950 = v_60947 & v_60949;
assign v_60952 = v_60818 & v_60951;
assign v_60954 = v_2627;
assign v_60956 = v_60953 & v_60955;
assign v_60958 = v_60815 & v_60957;
assign v_60960 = v_2623;
assign v_60962 = v_60959 & v_60961;
assign v_60963 = v_60962;
assign v_60965 = v_58431;
assign v_60966 = v_2688;
assign v_60967 = v_60966;
assign v_60968 = v_60965 & v_60967;
assign v_60969 = v_60968;
assign v_60970 = v_60860 & v_60969;
assign v_60972 = v_60870 & v_60971;
assign v_60973 = v_60859 & v_60969;
assign v_60975 = v_60857 & v_60974;
assign v_60977 = v_60876 & v_60976;
assign v_60978 = v_60856 & v_60974;
assign v_60980 = v_60854 & v_60979;
assign v_60982 = v_60882 & v_60981;
assign v_60983 = v_60853 & v_60979;
assign v_60985 = v_60851 & v_60984;
assign v_60987 = v_60888 & v_60986;
assign v_60988 = v_60850 & v_60984;
assign v_60990 = v_60848 & v_60989;
assign v_60992 = v_60894 & v_60991;
assign v_60993 = v_60847 & v_60989;
assign v_60995 = v_60845 & v_60994;
assign v_60997 = v_60900 & v_60996;
assign v_60998 = v_60844 & v_60994;
assign v_61000 = v_60842 & v_60999;
assign v_61002 = v_60906 & v_61001;
assign v_61003 = v_60841 & v_60999;
assign v_61005 = v_60839 & v_61004;
assign v_61007 = v_60912 & v_61006;
assign v_61008 = v_60838 & v_61004;
assign v_61010 = v_60836 & v_61009;
assign v_61012 = v_60918 & v_61011;
assign v_61013 = v_60835 & v_61009;
assign v_61015 = v_60833 & v_61014;
assign v_61017 = v_60924 & v_61016;
assign v_61018 = v_60832 & v_61014;
assign v_61020 = v_60830 & v_61019;
assign v_61022 = v_60930 & v_61021;
assign v_61023 = v_60829 & v_61019;
assign v_61025 = v_60827 & v_61024;
assign v_61027 = v_60936 & v_61026;
assign v_61028 = v_60826 & v_61024;
assign v_61030 = v_60824 & v_61029;
assign v_61032 = v_60942 & v_61031;
assign v_61033 = v_60823 & v_61029;
assign v_61035 = v_60821 & v_61034;
assign v_61037 = v_60948 & v_61036;
assign v_61038 = v_60820 & v_61034;
assign v_61040 = v_60818 & v_61039;
assign v_61042 = v_60954 & v_61041;
assign v_61043 = v_60817 & v_61039;
assign v_61045 = v_60815 & v_61044;
assign v_61047 = v_60960 & v_61046;
assign v_61048 = v_60814 & v_61044;
assign v_61050 = v_61049;
assign v_61052 = v_60964 & v_61051;
assign v_61053 = v_61052;
assign v_61055 = v_61054;
assign v_61057 = ~v_2883;
assign v_61058 = ~v_58368;
assign v_61059 = v_58368;
assign v_61060 = ~v_2887;
assign v_61061 = ~v_58372;
assign v_61062 = v_58372;
assign v_61063 = ~v_2891;
assign v_61064 = ~v_58376;
assign v_61065 = v_58376;
assign v_61066 = ~v_2895;
assign v_61067 = ~v_58380;
assign v_61068 = v_58380;
assign v_61069 = ~v_58383;
assign v_61070 = ~v_2900;
assign v_61071 = v_2900;
assign v_61072 = ~v_58387;
assign v_61073 = ~v_2904;
assign v_61074 = v_2904;
assign v_61075 = ~v_58391;
assign v_61076 = ~v_2908;
assign v_61077 = v_2908;
assign v_61078 = ~v_58395;
assign v_61079 = ~v_2912;
assign v_61080 = v_2912;
assign v_61081 = ~v_58399;
assign v_61082 = ~v_2916;
assign v_61083 = v_2916;
assign v_61084 = ~v_58403;
assign v_61085 = ~v_2920;
assign v_61086 = v_2920;
assign v_61087 = ~v_58407;
assign v_61088 = ~v_2924;
assign v_61089 = v_2924;
assign v_61090 = ~v_58411;
assign v_61091 = ~v_2928;
assign v_61092 = v_2928;
assign v_61093 = ~v_58415;
assign v_61094 = ~v_2932;
assign v_61095 = v_2932;
assign v_61096 = ~v_58419;
assign v_61097 = ~v_2936;
assign v_61098 = v_2936;
assign v_61099 = ~v_58423;
assign v_61100 = ~v_2940;
assign v_61101 = v_2940;
assign v_61102 = ~v_58427;
assign v_61103 = ~v_2944;
assign v_61104 = v_2944;
assign v_61105 = ~v_58431;
assign v_61106 = ~v_2948;
assign v_61107 = v_61106;
assign v_61109 = v_61108;
assign v_61111 = v_61103 & v_61110;
assign v_61113 = v_58427;
assign v_61115 = v_61112 & v_61114;
assign v_61117 = v_61100 & v_61116;
assign v_61119 = v_58423;
assign v_61121 = v_61118 & v_61120;
assign v_61123 = v_61097 & v_61122;
assign v_61125 = v_58419;
assign v_61127 = v_61124 & v_61126;
assign v_61129 = v_61094 & v_61128;
assign v_61131 = v_58415;
assign v_61133 = v_61130 & v_61132;
assign v_61135 = v_61091 & v_61134;
assign v_61137 = v_58411;
assign v_61139 = v_61136 & v_61138;
assign v_61141 = v_61088 & v_61140;
assign v_61143 = v_58407;
assign v_61145 = v_61142 & v_61144;
assign v_61147 = v_61085 & v_61146;
assign v_61149 = v_58403;
assign v_61151 = v_61148 & v_61150;
assign v_61153 = v_61082 & v_61152;
assign v_61155 = v_58399;
assign v_61157 = v_61154 & v_61156;
assign v_61159 = v_61079 & v_61158;
assign v_61161 = v_58395;
assign v_61163 = v_61160 & v_61162;
assign v_61165 = v_61076 & v_61164;
assign v_61167 = v_58391;
assign v_61169 = v_61166 & v_61168;
assign v_61171 = v_61073 & v_61170;
assign v_61173 = v_58387;
assign v_61175 = v_61172 & v_61174;
assign v_61177 = v_61070 & v_61176;
assign v_61179 = v_58383;
assign v_61181 = v_61178 & v_61180;
assign v_61183 = v_61067 & v_61182;
assign v_61185 = v_2895;
assign v_61187 = v_61184 & v_61186;
assign v_61189 = v_61064 & v_61188;
assign v_61191 = v_2891;
assign v_61193 = v_61190 & v_61192;
assign v_61195 = v_61061 & v_61194;
assign v_61197 = v_2887;
assign v_61199 = v_61196 & v_61198;
assign v_61201 = v_61058 & v_61200;
assign v_61203 = v_2883;
assign v_61205 = v_61202 & v_61204;
assign v_61206 = v_61205;
assign v_61208 = v_58431;
assign v_61209 = v_2948;
assign v_61210 = v_61209;
assign v_61211 = v_61208 & v_61210;
assign v_61212 = v_61211;
assign v_61213 = v_61103 & v_61212;
assign v_61215 = v_61113 & v_61214;
assign v_61216 = v_61102 & v_61212;
assign v_61218 = v_61100 & v_61217;
assign v_61220 = v_61119 & v_61219;
assign v_61221 = v_61099 & v_61217;
assign v_61223 = v_61097 & v_61222;
assign v_61225 = v_61125 & v_61224;
assign v_61226 = v_61096 & v_61222;
assign v_61228 = v_61094 & v_61227;
assign v_61230 = v_61131 & v_61229;
assign v_61231 = v_61093 & v_61227;
assign v_61233 = v_61091 & v_61232;
assign v_61235 = v_61137 & v_61234;
assign v_61236 = v_61090 & v_61232;
assign v_61238 = v_61088 & v_61237;
assign v_61240 = v_61143 & v_61239;
assign v_61241 = v_61087 & v_61237;
assign v_61243 = v_61085 & v_61242;
assign v_61245 = v_61149 & v_61244;
assign v_61246 = v_61084 & v_61242;
assign v_61248 = v_61082 & v_61247;
assign v_61250 = v_61155 & v_61249;
assign v_61251 = v_61081 & v_61247;
assign v_61253 = v_61079 & v_61252;
assign v_61255 = v_61161 & v_61254;
assign v_61256 = v_61078 & v_61252;
assign v_61258 = v_61076 & v_61257;
assign v_61260 = v_61167 & v_61259;
assign v_61261 = v_61075 & v_61257;
assign v_61263 = v_61073 & v_61262;
assign v_61265 = v_61173 & v_61264;
assign v_61266 = v_61072 & v_61262;
assign v_61268 = v_61070 & v_61267;
assign v_61270 = v_61179 & v_61269;
assign v_61271 = v_61069 & v_61267;
assign v_61273 = v_61067 & v_61272;
assign v_61275 = v_61185 & v_61274;
assign v_61276 = v_61066 & v_61272;
assign v_61278 = v_61064 & v_61277;
assign v_61280 = v_61191 & v_61279;
assign v_61281 = v_61063 & v_61277;
assign v_61283 = v_61061 & v_61282;
assign v_61285 = v_61197 & v_61284;
assign v_61286 = v_61060 & v_61282;
assign v_61288 = v_61058 & v_61287;
assign v_61290 = v_61203 & v_61289;
assign v_61291 = v_61057 & v_61287;
assign v_61293 = v_61292;
assign v_61295 = v_61207 & v_61294;
assign v_61296 = v_61295;
assign v_61298 = v_61297;
assign v_61300 = ~v_3143;
assign v_61301 = ~v_58368;
assign v_61302 = v_58368;
assign v_61303 = ~v_3147;
assign v_61304 = ~v_58372;
assign v_61305 = v_58372;
assign v_61306 = ~v_3151;
assign v_61307 = ~v_58376;
assign v_61308 = v_58376;
assign v_61309 = ~v_3155;
assign v_61310 = ~v_58380;
assign v_61311 = v_58380;
assign v_61312 = ~v_58383;
assign v_61313 = ~v_3160;
assign v_61314 = v_3160;
assign v_61315 = ~v_58387;
assign v_61316 = ~v_3164;
assign v_61317 = v_3164;
assign v_61318 = ~v_58391;
assign v_61319 = ~v_3168;
assign v_61320 = v_3168;
assign v_61321 = ~v_58395;
assign v_61322 = ~v_3172;
assign v_61323 = v_3172;
assign v_61324 = ~v_58399;
assign v_61325 = ~v_3176;
assign v_61326 = v_3176;
assign v_61327 = ~v_58403;
assign v_61328 = ~v_3180;
assign v_61329 = v_3180;
assign v_61330 = ~v_58407;
assign v_61331 = ~v_3184;
assign v_61332 = v_3184;
assign v_61333 = ~v_58411;
assign v_61334 = ~v_3188;
assign v_61335 = v_3188;
assign v_61336 = ~v_58415;
assign v_61337 = ~v_3192;
assign v_61338 = v_3192;
assign v_61339 = ~v_58419;
assign v_61340 = ~v_3196;
assign v_61341 = v_3196;
assign v_61342 = ~v_58423;
assign v_61343 = ~v_3200;
assign v_61344 = v_3200;
assign v_61345 = ~v_58427;
assign v_61346 = ~v_3204;
assign v_61347 = v_3204;
assign v_61348 = ~v_58431;
assign v_61349 = ~v_3208;
assign v_61350 = v_61349;
assign v_61352 = v_61351;
assign v_61354 = v_61346 & v_61353;
assign v_61356 = v_58427;
assign v_61358 = v_61355 & v_61357;
assign v_61360 = v_61343 & v_61359;
assign v_61362 = v_58423;
assign v_61364 = v_61361 & v_61363;
assign v_61366 = v_61340 & v_61365;
assign v_61368 = v_58419;
assign v_61370 = v_61367 & v_61369;
assign v_61372 = v_61337 & v_61371;
assign v_61374 = v_58415;
assign v_61376 = v_61373 & v_61375;
assign v_61378 = v_61334 & v_61377;
assign v_61380 = v_58411;
assign v_61382 = v_61379 & v_61381;
assign v_61384 = v_61331 & v_61383;
assign v_61386 = v_58407;
assign v_61388 = v_61385 & v_61387;
assign v_61390 = v_61328 & v_61389;
assign v_61392 = v_58403;
assign v_61394 = v_61391 & v_61393;
assign v_61396 = v_61325 & v_61395;
assign v_61398 = v_58399;
assign v_61400 = v_61397 & v_61399;
assign v_61402 = v_61322 & v_61401;
assign v_61404 = v_58395;
assign v_61406 = v_61403 & v_61405;
assign v_61408 = v_61319 & v_61407;
assign v_61410 = v_58391;
assign v_61412 = v_61409 & v_61411;
assign v_61414 = v_61316 & v_61413;
assign v_61416 = v_58387;
assign v_61418 = v_61415 & v_61417;
assign v_61420 = v_61313 & v_61419;
assign v_61422 = v_58383;
assign v_61424 = v_61421 & v_61423;
assign v_61426 = v_61310 & v_61425;
assign v_61428 = v_3155;
assign v_61430 = v_61427 & v_61429;
assign v_61432 = v_61307 & v_61431;
assign v_61434 = v_3151;
assign v_61436 = v_61433 & v_61435;
assign v_61438 = v_61304 & v_61437;
assign v_61440 = v_3147;
assign v_61442 = v_61439 & v_61441;
assign v_61444 = v_61301 & v_61443;
assign v_61446 = v_3143;
assign v_61448 = v_61445 & v_61447;
assign v_61449 = v_61448;
assign v_61451 = v_58431;
assign v_61452 = v_3208;
assign v_61453 = v_61452;
assign v_61454 = v_61451 & v_61453;
assign v_61455 = v_61454;
assign v_61456 = v_61346 & v_61455;
assign v_61458 = v_61356 & v_61457;
assign v_61459 = v_61345 & v_61455;
assign v_61461 = v_61343 & v_61460;
assign v_61463 = v_61362 & v_61462;
assign v_61464 = v_61342 & v_61460;
assign v_61466 = v_61340 & v_61465;
assign v_61468 = v_61368 & v_61467;
assign v_61469 = v_61339 & v_61465;
assign v_61471 = v_61337 & v_61470;
assign v_61473 = v_61374 & v_61472;
assign v_61474 = v_61336 & v_61470;
assign v_61476 = v_61334 & v_61475;
assign v_61478 = v_61380 & v_61477;
assign v_61479 = v_61333 & v_61475;
assign v_61481 = v_61331 & v_61480;
assign v_61483 = v_61386 & v_61482;
assign v_61484 = v_61330 & v_61480;
assign v_61486 = v_61328 & v_61485;
assign v_61488 = v_61392 & v_61487;
assign v_61489 = v_61327 & v_61485;
assign v_61491 = v_61325 & v_61490;
assign v_61493 = v_61398 & v_61492;
assign v_61494 = v_61324 & v_61490;
assign v_61496 = v_61322 & v_61495;
assign v_61498 = v_61404 & v_61497;
assign v_61499 = v_61321 & v_61495;
assign v_61501 = v_61319 & v_61500;
assign v_61503 = v_61410 & v_61502;
assign v_61504 = v_61318 & v_61500;
assign v_61506 = v_61316 & v_61505;
assign v_61508 = v_61416 & v_61507;
assign v_61509 = v_61315 & v_61505;
assign v_61511 = v_61313 & v_61510;
assign v_61513 = v_61422 & v_61512;
assign v_61514 = v_61312 & v_61510;
assign v_61516 = v_61310 & v_61515;
assign v_61518 = v_61428 & v_61517;
assign v_61519 = v_61309 & v_61515;
assign v_61521 = v_61307 & v_61520;
assign v_61523 = v_61434 & v_61522;
assign v_61524 = v_61306 & v_61520;
assign v_61526 = v_61304 & v_61525;
assign v_61528 = v_61440 & v_61527;
assign v_61529 = v_61303 & v_61525;
assign v_61531 = v_61301 & v_61530;
assign v_61533 = v_61446 & v_61532;
assign v_61534 = v_61300 & v_61530;
assign v_61536 = v_61535;
assign v_61538 = v_61450 & v_61537;
assign v_61539 = v_61538;
assign v_61541 = v_61540;
assign v_61543 = ~v_3403;
assign v_61544 = ~v_58368;
assign v_61545 = v_58368;
assign v_61546 = ~v_3407;
assign v_61547 = ~v_58372;
assign v_61548 = v_58372;
assign v_61549 = ~v_3411;
assign v_61550 = ~v_58376;
assign v_61551 = v_58376;
assign v_61552 = ~v_3415;
assign v_61553 = ~v_58380;
assign v_61554 = v_58380;
assign v_61555 = ~v_58383;
assign v_61556 = ~v_3420;
assign v_61557 = v_3420;
assign v_61558 = ~v_58387;
assign v_61559 = ~v_3424;
assign v_61560 = v_3424;
assign v_61561 = ~v_58391;
assign v_61562 = ~v_3428;
assign v_61563 = v_3428;
assign v_61564 = ~v_58395;
assign v_61565 = ~v_3432;
assign v_61566 = v_3432;
assign v_61567 = ~v_58399;
assign v_61568 = ~v_3436;
assign v_61569 = v_3436;
assign v_61570 = ~v_58403;
assign v_61571 = ~v_3440;
assign v_61572 = v_3440;
assign v_61573 = ~v_58407;
assign v_61574 = ~v_3444;
assign v_61575 = v_3444;
assign v_61576 = ~v_58411;
assign v_61577 = ~v_3448;
assign v_61578 = v_3448;
assign v_61579 = ~v_58415;
assign v_61580 = ~v_3452;
assign v_61581 = v_3452;
assign v_61582 = ~v_58419;
assign v_61583 = ~v_3456;
assign v_61584 = v_3456;
assign v_61585 = ~v_58423;
assign v_61586 = ~v_3460;
assign v_61587 = v_3460;
assign v_61588 = ~v_58427;
assign v_61589 = ~v_3464;
assign v_61590 = v_3464;
assign v_61591 = ~v_58431;
assign v_61592 = ~v_3468;
assign v_61593 = v_61592;
assign v_61595 = v_61594;
assign v_61597 = v_61589 & v_61596;
assign v_61599 = v_58427;
assign v_61601 = v_61598 & v_61600;
assign v_61603 = v_61586 & v_61602;
assign v_61605 = v_58423;
assign v_61607 = v_61604 & v_61606;
assign v_61609 = v_61583 & v_61608;
assign v_61611 = v_58419;
assign v_61613 = v_61610 & v_61612;
assign v_61615 = v_61580 & v_61614;
assign v_61617 = v_58415;
assign v_61619 = v_61616 & v_61618;
assign v_61621 = v_61577 & v_61620;
assign v_61623 = v_58411;
assign v_61625 = v_61622 & v_61624;
assign v_61627 = v_61574 & v_61626;
assign v_61629 = v_58407;
assign v_61631 = v_61628 & v_61630;
assign v_61633 = v_61571 & v_61632;
assign v_61635 = v_58403;
assign v_61637 = v_61634 & v_61636;
assign v_61639 = v_61568 & v_61638;
assign v_61641 = v_58399;
assign v_61643 = v_61640 & v_61642;
assign v_61645 = v_61565 & v_61644;
assign v_61647 = v_58395;
assign v_61649 = v_61646 & v_61648;
assign v_61651 = v_61562 & v_61650;
assign v_61653 = v_58391;
assign v_61655 = v_61652 & v_61654;
assign v_61657 = v_61559 & v_61656;
assign v_61659 = v_58387;
assign v_61661 = v_61658 & v_61660;
assign v_61663 = v_61556 & v_61662;
assign v_61665 = v_58383;
assign v_61667 = v_61664 & v_61666;
assign v_61669 = v_61553 & v_61668;
assign v_61671 = v_3415;
assign v_61673 = v_61670 & v_61672;
assign v_61675 = v_61550 & v_61674;
assign v_61677 = v_3411;
assign v_61679 = v_61676 & v_61678;
assign v_61681 = v_61547 & v_61680;
assign v_61683 = v_3407;
assign v_61685 = v_61682 & v_61684;
assign v_61687 = v_61544 & v_61686;
assign v_61689 = v_3403;
assign v_61691 = v_61688 & v_61690;
assign v_61692 = v_61691;
assign v_61694 = v_58431;
assign v_61695 = v_3468;
assign v_61696 = v_61695;
assign v_61697 = v_61694 & v_61696;
assign v_61698 = v_61697;
assign v_61699 = v_61589 & v_61698;
assign v_61701 = v_61599 & v_61700;
assign v_61702 = v_61588 & v_61698;
assign v_61704 = v_61586 & v_61703;
assign v_61706 = v_61605 & v_61705;
assign v_61707 = v_61585 & v_61703;
assign v_61709 = v_61583 & v_61708;
assign v_61711 = v_61611 & v_61710;
assign v_61712 = v_61582 & v_61708;
assign v_61714 = v_61580 & v_61713;
assign v_61716 = v_61617 & v_61715;
assign v_61717 = v_61579 & v_61713;
assign v_61719 = v_61577 & v_61718;
assign v_61721 = v_61623 & v_61720;
assign v_61722 = v_61576 & v_61718;
assign v_61724 = v_61574 & v_61723;
assign v_61726 = v_61629 & v_61725;
assign v_61727 = v_61573 & v_61723;
assign v_61729 = v_61571 & v_61728;
assign v_61731 = v_61635 & v_61730;
assign v_61732 = v_61570 & v_61728;
assign v_61734 = v_61568 & v_61733;
assign v_61736 = v_61641 & v_61735;
assign v_61737 = v_61567 & v_61733;
assign v_61739 = v_61565 & v_61738;
assign v_61741 = v_61647 & v_61740;
assign v_61742 = v_61564 & v_61738;
assign v_61744 = v_61562 & v_61743;
assign v_61746 = v_61653 & v_61745;
assign v_61747 = v_61561 & v_61743;
assign v_61749 = v_61559 & v_61748;
assign v_61751 = v_61659 & v_61750;
assign v_61752 = v_61558 & v_61748;
assign v_61754 = v_61556 & v_61753;
assign v_61756 = v_61665 & v_61755;
assign v_61757 = v_61555 & v_61753;
assign v_61759 = v_61553 & v_61758;
assign v_61761 = v_61671 & v_61760;
assign v_61762 = v_61552 & v_61758;
assign v_61764 = v_61550 & v_61763;
assign v_61766 = v_61677 & v_61765;
assign v_61767 = v_61549 & v_61763;
assign v_61769 = v_61547 & v_61768;
assign v_61771 = v_61683 & v_61770;
assign v_61772 = v_61546 & v_61768;
assign v_61774 = v_61544 & v_61773;
assign v_61776 = v_61689 & v_61775;
assign v_61777 = v_61543 & v_61773;
assign v_61779 = v_61778;
assign v_61781 = v_61693 & v_61780;
assign v_61782 = v_61781;
assign v_61784 = v_61783;
assign v_61786 = ~v_3663;
assign v_61787 = ~v_58368;
assign v_61788 = v_58368;
assign v_61789 = ~v_3667;
assign v_61790 = ~v_58372;
assign v_61791 = v_58372;
assign v_61792 = ~v_3671;
assign v_61793 = ~v_58376;
assign v_61794 = v_58376;
assign v_61795 = ~v_3675;
assign v_61796 = ~v_58380;
assign v_61797 = v_58380;
assign v_61798 = ~v_58383;
assign v_61799 = ~v_3680;
assign v_61800 = v_3680;
assign v_61801 = ~v_58387;
assign v_61802 = ~v_3684;
assign v_61803 = v_3684;
assign v_61804 = ~v_58391;
assign v_61805 = ~v_3688;
assign v_61806 = v_3688;
assign v_61807 = ~v_58395;
assign v_61808 = ~v_3692;
assign v_61809 = v_3692;
assign v_61810 = ~v_58399;
assign v_61811 = ~v_3696;
assign v_61812 = v_3696;
assign v_61813 = ~v_58403;
assign v_61814 = ~v_3700;
assign v_61815 = v_3700;
assign v_61816 = ~v_58407;
assign v_61817 = ~v_3704;
assign v_61818 = v_3704;
assign v_61819 = ~v_58411;
assign v_61820 = ~v_3708;
assign v_61821 = v_3708;
assign v_61822 = ~v_58415;
assign v_61823 = ~v_3712;
assign v_61824 = v_3712;
assign v_61825 = ~v_58419;
assign v_61826 = ~v_3716;
assign v_61827 = v_3716;
assign v_61828 = ~v_58423;
assign v_61829 = ~v_3720;
assign v_61830 = v_3720;
assign v_61831 = ~v_58427;
assign v_61832 = ~v_3724;
assign v_61833 = v_3724;
assign v_61834 = ~v_58431;
assign v_61835 = ~v_3728;
assign v_61836 = v_61835;
assign v_61838 = v_61837;
assign v_61840 = v_61832 & v_61839;
assign v_61842 = v_58427;
assign v_61844 = v_61841 & v_61843;
assign v_61846 = v_61829 & v_61845;
assign v_61848 = v_58423;
assign v_61850 = v_61847 & v_61849;
assign v_61852 = v_61826 & v_61851;
assign v_61854 = v_58419;
assign v_61856 = v_61853 & v_61855;
assign v_61858 = v_61823 & v_61857;
assign v_61860 = v_58415;
assign v_61862 = v_61859 & v_61861;
assign v_61864 = v_61820 & v_61863;
assign v_61866 = v_58411;
assign v_61868 = v_61865 & v_61867;
assign v_61870 = v_61817 & v_61869;
assign v_61872 = v_58407;
assign v_61874 = v_61871 & v_61873;
assign v_61876 = v_61814 & v_61875;
assign v_61878 = v_58403;
assign v_61880 = v_61877 & v_61879;
assign v_61882 = v_61811 & v_61881;
assign v_61884 = v_58399;
assign v_61886 = v_61883 & v_61885;
assign v_61888 = v_61808 & v_61887;
assign v_61890 = v_58395;
assign v_61892 = v_61889 & v_61891;
assign v_61894 = v_61805 & v_61893;
assign v_61896 = v_58391;
assign v_61898 = v_61895 & v_61897;
assign v_61900 = v_61802 & v_61899;
assign v_61902 = v_58387;
assign v_61904 = v_61901 & v_61903;
assign v_61906 = v_61799 & v_61905;
assign v_61908 = v_58383;
assign v_61910 = v_61907 & v_61909;
assign v_61912 = v_61796 & v_61911;
assign v_61914 = v_3675;
assign v_61916 = v_61913 & v_61915;
assign v_61918 = v_61793 & v_61917;
assign v_61920 = v_3671;
assign v_61922 = v_61919 & v_61921;
assign v_61924 = v_61790 & v_61923;
assign v_61926 = v_3667;
assign v_61928 = v_61925 & v_61927;
assign v_61930 = v_61787 & v_61929;
assign v_61932 = v_3663;
assign v_61934 = v_61931 & v_61933;
assign v_61935 = v_61934;
assign v_61937 = v_58431;
assign v_61938 = v_3728;
assign v_61939 = v_61938;
assign v_61940 = v_61937 & v_61939;
assign v_61941 = v_61940;
assign v_61942 = v_61832 & v_61941;
assign v_61944 = v_61842 & v_61943;
assign v_61945 = v_61831 & v_61941;
assign v_61947 = v_61829 & v_61946;
assign v_61949 = v_61848 & v_61948;
assign v_61950 = v_61828 & v_61946;
assign v_61952 = v_61826 & v_61951;
assign v_61954 = v_61854 & v_61953;
assign v_61955 = v_61825 & v_61951;
assign v_61957 = v_61823 & v_61956;
assign v_61959 = v_61860 & v_61958;
assign v_61960 = v_61822 & v_61956;
assign v_61962 = v_61820 & v_61961;
assign v_61964 = v_61866 & v_61963;
assign v_61965 = v_61819 & v_61961;
assign v_61967 = v_61817 & v_61966;
assign v_61969 = v_61872 & v_61968;
assign v_61970 = v_61816 & v_61966;
assign v_61972 = v_61814 & v_61971;
assign v_61974 = v_61878 & v_61973;
assign v_61975 = v_61813 & v_61971;
assign v_61977 = v_61811 & v_61976;
assign v_61979 = v_61884 & v_61978;
assign v_61980 = v_61810 & v_61976;
assign v_61982 = v_61808 & v_61981;
assign v_61984 = v_61890 & v_61983;
assign v_61985 = v_61807 & v_61981;
assign v_61987 = v_61805 & v_61986;
assign v_61989 = v_61896 & v_61988;
assign v_61990 = v_61804 & v_61986;
assign v_61992 = v_61802 & v_61991;
assign v_61994 = v_61902 & v_61993;
assign v_61995 = v_61801 & v_61991;
assign v_61997 = v_61799 & v_61996;
assign v_61999 = v_61908 & v_61998;
assign v_62000 = v_61798 & v_61996;
assign v_62002 = v_61796 & v_62001;
assign v_62004 = v_61914 & v_62003;
assign v_62005 = v_61795 & v_62001;
assign v_62007 = v_61793 & v_62006;
assign v_62009 = v_61920 & v_62008;
assign v_62010 = v_61792 & v_62006;
assign v_62012 = v_61790 & v_62011;
assign v_62014 = v_61926 & v_62013;
assign v_62015 = v_61789 & v_62011;
assign v_62017 = v_61787 & v_62016;
assign v_62019 = v_61932 & v_62018;
assign v_62020 = v_61786 & v_62016;
assign v_62022 = v_62021;
assign v_62024 = v_61936 & v_62023;
assign v_62025 = v_62024;
assign v_62027 = v_62026;
assign v_62029 = ~v_3923;
assign v_62030 = ~v_58368;
assign v_62031 = v_58368;
assign v_62032 = ~v_3927;
assign v_62033 = ~v_58372;
assign v_62034 = v_58372;
assign v_62035 = ~v_3931;
assign v_62036 = ~v_58376;
assign v_62037 = v_58376;
assign v_62038 = ~v_3935;
assign v_62039 = ~v_58380;
assign v_62040 = v_58380;
assign v_62041 = ~v_58383;
assign v_62042 = ~v_3940;
assign v_62043 = v_3940;
assign v_62044 = ~v_58387;
assign v_62045 = ~v_3944;
assign v_62046 = v_3944;
assign v_62047 = ~v_58391;
assign v_62048 = ~v_3948;
assign v_62049 = v_3948;
assign v_62050 = ~v_58395;
assign v_62051 = ~v_3952;
assign v_62052 = v_3952;
assign v_62053 = ~v_58399;
assign v_62054 = ~v_3956;
assign v_62055 = v_3956;
assign v_62056 = ~v_58403;
assign v_62057 = ~v_3960;
assign v_62058 = v_3960;
assign v_62059 = ~v_58407;
assign v_62060 = ~v_3964;
assign v_62061 = v_3964;
assign v_62062 = ~v_58411;
assign v_62063 = ~v_3968;
assign v_62064 = v_3968;
assign v_62065 = ~v_58415;
assign v_62066 = ~v_3972;
assign v_62067 = v_3972;
assign v_62068 = ~v_58419;
assign v_62069 = ~v_3976;
assign v_62070 = v_3976;
assign v_62071 = ~v_58423;
assign v_62072 = ~v_3980;
assign v_62073 = v_3980;
assign v_62074 = ~v_58427;
assign v_62075 = ~v_3984;
assign v_62076 = v_3984;
assign v_62077 = ~v_58431;
assign v_62078 = ~v_3988;
assign v_62079 = v_62078;
assign v_62081 = v_62080;
assign v_62083 = v_62075 & v_62082;
assign v_62085 = v_58427;
assign v_62087 = v_62084 & v_62086;
assign v_62089 = v_62072 & v_62088;
assign v_62091 = v_58423;
assign v_62093 = v_62090 & v_62092;
assign v_62095 = v_62069 & v_62094;
assign v_62097 = v_58419;
assign v_62099 = v_62096 & v_62098;
assign v_62101 = v_62066 & v_62100;
assign v_62103 = v_58415;
assign v_62105 = v_62102 & v_62104;
assign v_62107 = v_62063 & v_62106;
assign v_62109 = v_58411;
assign v_62111 = v_62108 & v_62110;
assign v_62113 = v_62060 & v_62112;
assign v_62115 = v_58407;
assign v_62117 = v_62114 & v_62116;
assign v_62119 = v_62057 & v_62118;
assign v_62121 = v_58403;
assign v_62123 = v_62120 & v_62122;
assign v_62125 = v_62054 & v_62124;
assign v_62127 = v_58399;
assign v_62129 = v_62126 & v_62128;
assign v_62131 = v_62051 & v_62130;
assign v_62133 = v_58395;
assign v_62135 = v_62132 & v_62134;
assign v_62137 = v_62048 & v_62136;
assign v_62139 = v_58391;
assign v_62141 = v_62138 & v_62140;
assign v_62143 = v_62045 & v_62142;
assign v_62145 = v_58387;
assign v_62147 = v_62144 & v_62146;
assign v_62149 = v_62042 & v_62148;
assign v_62151 = v_58383;
assign v_62153 = v_62150 & v_62152;
assign v_62155 = v_62039 & v_62154;
assign v_62157 = v_3935;
assign v_62159 = v_62156 & v_62158;
assign v_62161 = v_62036 & v_62160;
assign v_62163 = v_3931;
assign v_62165 = v_62162 & v_62164;
assign v_62167 = v_62033 & v_62166;
assign v_62169 = v_3927;
assign v_62171 = v_62168 & v_62170;
assign v_62173 = v_62030 & v_62172;
assign v_62175 = v_3923;
assign v_62177 = v_62174 & v_62176;
assign v_62178 = v_62177;
assign v_62180 = v_58431;
assign v_62181 = v_3988;
assign v_62182 = v_62181;
assign v_62183 = v_62180 & v_62182;
assign v_62184 = v_62183;
assign v_62185 = v_62075 & v_62184;
assign v_62187 = v_62085 & v_62186;
assign v_62188 = v_62074 & v_62184;
assign v_62190 = v_62072 & v_62189;
assign v_62192 = v_62091 & v_62191;
assign v_62193 = v_62071 & v_62189;
assign v_62195 = v_62069 & v_62194;
assign v_62197 = v_62097 & v_62196;
assign v_62198 = v_62068 & v_62194;
assign v_62200 = v_62066 & v_62199;
assign v_62202 = v_62103 & v_62201;
assign v_62203 = v_62065 & v_62199;
assign v_62205 = v_62063 & v_62204;
assign v_62207 = v_62109 & v_62206;
assign v_62208 = v_62062 & v_62204;
assign v_62210 = v_62060 & v_62209;
assign v_62212 = v_62115 & v_62211;
assign v_62213 = v_62059 & v_62209;
assign v_62215 = v_62057 & v_62214;
assign v_62217 = v_62121 & v_62216;
assign v_62218 = v_62056 & v_62214;
assign v_62220 = v_62054 & v_62219;
assign v_62222 = v_62127 & v_62221;
assign v_62223 = v_62053 & v_62219;
assign v_62225 = v_62051 & v_62224;
assign v_62227 = v_62133 & v_62226;
assign v_62228 = v_62050 & v_62224;
assign v_62230 = v_62048 & v_62229;
assign v_62232 = v_62139 & v_62231;
assign v_62233 = v_62047 & v_62229;
assign v_62235 = v_62045 & v_62234;
assign v_62237 = v_62145 & v_62236;
assign v_62238 = v_62044 & v_62234;
assign v_62240 = v_62042 & v_62239;
assign v_62242 = v_62151 & v_62241;
assign v_62243 = v_62041 & v_62239;
assign v_62245 = v_62039 & v_62244;
assign v_62247 = v_62157 & v_62246;
assign v_62248 = v_62038 & v_62244;
assign v_62250 = v_62036 & v_62249;
assign v_62252 = v_62163 & v_62251;
assign v_62253 = v_62035 & v_62249;
assign v_62255 = v_62033 & v_62254;
assign v_62257 = v_62169 & v_62256;
assign v_62258 = v_62032 & v_62254;
assign v_62260 = v_62030 & v_62259;
assign v_62262 = v_62175 & v_62261;
assign v_62263 = v_62029 & v_62259;
assign v_62265 = v_62264;
assign v_62267 = v_62179 & v_62266;
assign v_62268 = v_62267;
assign v_62270 = v_62269;
assign v_62271 = ~v_4182;
assign v_62272 = ~v_58368;
assign v_62273 = v_58368;
assign v_62274 = ~v_4186;
assign v_62275 = ~v_58372;
assign v_62276 = v_58372;
assign v_62277 = ~v_4190;
assign v_62278 = ~v_58376;
assign v_62279 = v_58376;
assign v_62280 = ~v_4194;
assign v_62281 = ~v_58380;
assign v_62282 = v_58380;
assign v_62283 = ~v_58383;
assign v_62284 = ~v_4199;
assign v_62285 = v_4199;
assign v_62286 = ~v_58387;
assign v_62287 = ~v_4203;
assign v_62288 = v_4203;
assign v_62289 = ~v_58391;
assign v_62290 = ~v_4207;
assign v_62291 = v_4207;
assign v_62292 = ~v_58395;
assign v_62293 = ~v_4211;
assign v_62294 = v_4211;
assign v_62295 = ~v_58399;
assign v_62296 = ~v_4215;
assign v_62297 = v_4215;
assign v_62298 = ~v_58403;
assign v_62299 = ~v_4219;
assign v_62300 = v_4219;
assign v_62301 = ~v_58407;
assign v_62302 = ~v_4223;
assign v_62303 = v_4223;
assign v_62304 = ~v_58411;
assign v_62305 = ~v_4227;
assign v_62306 = v_4227;
assign v_62307 = ~v_58415;
assign v_62308 = ~v_4231;
assign v_62309 = v_4231;
assign v_62310 = ~v_58419;
assign v_62311 = ~v_4235;
assign v_62312 = v_4235;
assign v_62313 = ~v_58423;
assign v_62314 = ~v_4239;
assign v_62315 = v_4239;
assign v_62316 = ~v_58427;
assign v_62317 = ~v_4243;
assign v_62318 = v_4243;
assign v_62319 = ~v_58431;
assign v_62320 = ~v_4247;
assign v_62321 = v_62320;
assign v_62323 = v_62322;
assign v_62325 = v_62317 & v_62324;
assign v_62327 = v_58427;
assign v_62329 = v_62326 & v_62328;
assign v_62331 = v_62314 & v_62330;
assign v_62333 = v_58423;
assign v_62335 = v_62332 & v_62334;
assign v_62337 = v_62311 & v_62336;
assign v_62339 = v_58419;
assign v_62341 = v_62338 & v_62340;
assign v_62343 = v_62308 & v_62342;
assign v_62345 = v_58415;
assign v_62347 = v_62344 & v_62346;
assign v_62349 = v_62305 & v_62348;
assign v_62351 = v_58411;
assign v_62353 = v_62350 & v_62352;
assign v_62355 = v_62302 & v_62354;
assign v_62357 = v_58407;
assign v_62359 = v_62356 & v_62358;
assign v_62361 = v_62299 & v_62360;
assign v_62363 = v_58403;
assign v_62365 = v_62362 & v_62364;
assign v_62367 = v_62296 & v_62366;
assign v_62369 = v_58399;
assign v_62371 = v_62368 & v_62370;
assign v_62373 = v_62293 & v_62372;
assign v_62375 = v_58395;
assign v_62377 = v_62374 & v_62376;
assign v_62379 = v_62290 & v_62378;
assign v_62381 = v_58391;
assign v_62383 = v_62380 & v_62382;
assign v_62385 = v_62287 & v_62384;
assign v_62387 = v_58387;
assign v_62389 = v_62386 & v_62388;
assign v_62391 = v_62284 & v_62390;
assign v_62393 = v_58383;
assign v_62395 = v_62392 & v_62394;
assign v_62397 = v_62281 & v_62396;
assign v_62399 = v_4194;
assign v_62401 = v_62398 & v_62400;
assign v_62403 = v_62278 & v_62402;
assign v_62405 = v_4190;
assign v_62407 = v_62404 & v_62406;
assign v_62409 = v_62275 & v_62408;
assign v_62411 = v_4186;
assign v_62413 = v_62410 & v_62412;
assign v_62415 = v_62272 & v_62414;
assign v_62417 = v_4182;
assign v_62419 = v_62416 & v_62418;
assign v_62421 = ~v_62420;
assign v_62423 = v_58431;
assign v_62424 = v_4247;
assign v_62425 = v_62424;
assign v_62426 = v_62423 & v_62425;
assign v_62427 = v_62426;
assign v_62428 = v_62317 & v_62427;
assign v_62430 = v_62327 & v_62429;
assign v_62431 = v_62316 & v_62427;
assign v_62433 = v_62314 & v_62432;
assign v_62435 = v_62333 & v_62434;
assign v_62436 = v_62313 & v_62432;
assign v_62438 = v_62311 & v_62437;
assign v_62440 = v_62339 & v_62439;
assign v_62441 = v_62310 & v_62437;
assign v_62443 = v_62308 & v_62442;
assign v_62445 = v_62345 & v_62444;
assign v_62446 = v_62307 & v_62442;
assign v_62448 = v_62305 & v_62447;
assign v_62450 = v_62351 & v_62449;
assign v_62451 = v_62304 & v_62447;
assign v_62453 = v_62302 & v_62452;
assign v_62455 = v_62357 & v_62454;
assign v_62456 = v_62301 & v_62452;
assign v_62458 = v_62299 & v_62457;
assign v_62460 = v_62363 & v_62459;
assign v_62461 = v_62298 & v_62457;
assign v_62463 = v_62296 & v_62462;
assign v_62465 = v_62369 & v_62464;
assign v_62466 = v_62295 & v_62462;
assign v_62468 = v_62293 & v_62467;
assign v_62470 = v_62375 & v_62469;
assign v_62471 = v_62292 & v_62467;
assign v_62473 = v_62290 & v_62472;
assign v_62475 = v_62381 & v_62474;
assign v_62476 = v_62289 & v_62472;
assign v_62478 = v_62287 & v_62477;
assign v_62480 = v_62387 & v_62479;
assign v_62481 = v_62286 & v_62477;
assign v_62483 = v_62284 & v_62482;
assign v_62485 = v_62393 & v_62484;
assign v_62486 = v_62283 & v_62482;
assign v_62488 = v_62281 & v_62487;
assign v_62490 = v_62399 & v_62489;
assign v_62491 = v_62280 & v_62487;
assign v_62493 = v_62278 & v_62492;
assign v_62495 = v_62405 & v_62494;
assign v_62496 = v_62277 & v_62492;
assign v_62498 = v_62275 & v_62497;
assign v_62500 = v_62411 & v_62499;
assign v_62501 = v_62274 & v_62497;
assign v_62503 = v_62272 & v_62502;
assign v_62505 = v_62417 & v_62504;
assign v_62506 = v_62271 & v_62502;
assign v_62508 = v_62420;
assign v_62510 = v_62422 & v_62509;
assign v_62511 = v_62510;
assign v_62513 = v_62512;
assign v_62515 = ~v_6;
assign v_62517 = ~v_62516;
assign v_62518 = v_62516;
assign v_62519 = ~v_13;
assign v_62521 = ~v_62520;
assign v_62522 = v_62520;
assign v_62523 = ~v_18;
assign v_62525 = ~v_62524;
assign v_62526 = v_62524;
assign v_62527 = ~v_23;
assign v_62529 = ~v_62528;
assign v_62530 = v_62528;
assign v_62532 = ~v_62531;
assign v_62533 = ~v_30;
assign v_62534 = v_30;
assign v_62536 = ~v_62535;
assign v_62537 = ~v_35;
assign v_62538 = v_35;
assign v_62540 = ~v_62539;
assign v_62541 = ~v_40;
assign v_62542 = v_40;
assign v_62544 = ~v_62543;
assign v_62545 = ~v_45;
assign v_62546 = v_45;
assign v_62548 = ~v_62547;
assign v_62549 = ~v_50;
assign v_62550 = v_50;
assign v_62552 = ~v_62551;
assign v_62553 = ~v_55;
assign v_62554 = v_55;
assign v_62556 = ~v_62555;
assign v_62557 = ~v_60;
assign v_62558 = v_60;
assign v_62560 = ~v_62559;
assign v_62561 = ~v_65;
assign v_62562 = v_65;
assign v_62564 = ~v_62563;
assign v_62565 = ~v_70;
assign v_62566 = v_70;
assign v_62568 = ~v_62567;
assign v_62569 = ~v_75;
assign v_62570 = v_75;
assign v_62572 = ~v_62571;
assign v_62573 = ~v_80;
assign v_62574 = v_80;
assign v_62576 = ~v_62575;
assign v_62577 = ~v_85;
assign v_62578 = v_85;
assign v_62580 = ~v_62579;
assign v_62581 = ~v_90;
assign v_62582 = v_62581;
assign v_62584 = v_62583;
assign v_62586 = v_62577 & v_62585;
assign v_62588 = v_62575;
assign v_62590 = v_62587 & v_62589;
assign v_62592 = v_62573 & v_62591;
assign v_62594 = v_62571;
assign v_62596 = v_62593 & v_62595;
assign v_62598 = v_62569 & v_62597;
assign v_62600 = v_62567;
assign v_62602 = v_62599 & v_62601;
assign v_62604 = v_62565 & v_62603;
assign v_62606 = v_62563;
assign v_62608 = v_62605 & v_62607;
assign v_62610 = v_62561 & v_62609;
assign v_62612 = v_62559;
assign v_62614 = v_62611 & v_62613;
assign v_62616 = v_62557 & v_62615;
assign v_62618 = v_62555;
assign v_62620 = v_62617 & v_62619;
assign v_62622 = v_62553 & v_62621;
assign v_62624 = v_62551;
assign v_62626 = v_62623 & v_62625;
assign v_62628 = v_62549 & v_62627;
assign v_62630 = v_62547;
assign v_62632 = v_62629 & v_62631;
assign v_62634 = v_62545 & v_62633;
assign v_62636 = v_62543;
assign v_62638 = v_62635 & v_62637;
assign v_62640 = v_62541 & v_62639;
assign v_62642 = v_62539;
assign v_62644 = v_62641 & v_62643;
assign v_62646 = v_62537 & v_62645;
assign v_62648 = v_62535;
assign v_62650 = v_62647 & v_62649;
assign v_62652 = v_62533 & v_62651;
assign v_62654 = v_62531;
assign v_62656 = v_62653 & v_62655;
assign v_62658 = v_62529 & v_62657;
assign v_62660 = v_23;
assign v_62662 = v_62659 & v_62661;
assign v_62664 = v_62525 & v_62663;
assign v_62666 = v_18;
assign v_62668 = v_62665 & v_62667;
assign v_62670 = v_62521 & v_62669;
assign v_62672 = v_13;
assign v_62674 = v_62671 & v_62673;
assign v_62676 = v_62517 & v_62675;
assign v_62678 = v_6;
assign v_62680 = v_62677 & v_62679;
assign v_62681 = v_62680;
assign v_62683 = v_62579;
assign v_62684 = v_90;
assign v_62685 = v_62684;
assign v_62686 = v_62683 & v_62685;
assign v_62687 = v_62686;
assign v_62688 = v_62577 & v_62687;
assign v_62690 = v_62588 & v_62689;
assign v_62691 = v_62576 & v_62687;
assign v_62693 = v_62573 & v_62692;
assign v_62695 = v_62594 & v_62694;
assign v_62696 = v_62572 & v_62692;
assign v_62698 = v_62569 & v_62697;
assign v_62700 = v_62600 & v_62699;
assign v_62701 = v_62568 & v_62697;
assign v_62703 = v_62565 & v_62702;
assign v_62705 = v_62606 & v_62704;
assign v_62706 = v_62564 & v_62702;
assign v_62708 = v_62561 & v_62707;
assign v_62710 = v_62612 & v_62709;
assign v_62711 = v_62560 & v_62707;
assign v_62713 = v_62557 & v_62712;
assign v_62715 = v_62618 & v_62714;
assign v_62716 = v_62556 & v_62712;
assign v_62718 = v_62553 & v_62717;
assign v_62720 = v_62624 & v_62719;
assign v_62721 = v_62552 & v_62717;
assign v_62723 = v_62549 & v_62722;
assign v_62725 = v_62630 & v_62724;
assign v_62726 = v_62548 & v_62722;
assign v_62728 = v_62545 & v_62727;
assign v_62730 = v_62636 & v_62729;
assign v_62731 = v_62544 & v_62727;
assign v_62733 = v_62541 & v_62732;
assign v_62735 = v_62642 & v_62734;
assign v_62736 = v_62540 & v_62732;
assign v_62738 = v_62537 & v_62737;
assign v_62740 = v_62648 & v_62739;
assign v_62741 = v_62536 & v_62737;
assign v_62743 = v_62533 & v_62742;
assign v_62745 = v_62654 & v_62744;
assign v_62746 = v_62532 & v_62742;
assign v_62748 = v_62529 & v_62747;
assign v_62750 = v_62660 & v_62749;
assign v_62751 = v_62527 & v_62747;
assign v_62753 = v_62525 & v_62752;
assign v_62755 = v_62666 & v_62754;
assign v_62756 = v_62523 & v_62752;
assign v_62758 = v_62521 & v_62757;
assign v_62760 = v_62672 & v_62759;
assign v_62761 = v_62519 & v_62757;
assign v_62763 = v_62517 & v_62762;
assign v_62765 = v_62678 & v_62764;
assign v_62766 = v_62515 & v_62762;
assign v_62768 = v_62767;
assign v_62770 = v_62682 & v_62769;
assign v_62771 = v_62770;
assign v_62773 = v_62772;
assign v_62775 = ~v_283;
assign v_62776 = ~v_62516;
assign v_62777 = v_62516;
assign v_62778 = ~v_287;
assign v_62779 = ~v_62520;
assign v_62780 = v_62520;
assign v_62781 = ~v_291;
assign v_62782 = ~v_62524;
assign v_62783 = v_62524;
assign v_62784 = ~v_295;
assign v_62785 = ~v_62528;
assign v_62786 = v_62528;
assign v_62787 = ~v_62531;
assign v_62788 = ~v_300;
assign v_62789 = v_300;
assign v_62790 = ~v_62535;
assign v_62791 = ~v_304;
assign v_62792 = v_304;
assign v_62793 = ~v_62539;
assign v_62794 = ~v_308;
assign v_62795 = v_308;
assign v_62796 = ~v_62543;
assign v_62797 = ~v_312;
assign v_62798 = v_312;
assign v_62799 = ~v_62547;
assign v_62800 = ~v_316;
assign v_62801 = v_316;
assign v_62802 = ~v_62551;
assign v_62803 = ~v_320;
assign v_62804 = v_320;
assign v_62805 = ~v_62555;
assign v_62806 = ~v_324;
assign v_62807 = v_324;
assign v_62808 = ~v_62559;
assign v_62809 = ~v_328;
assign v_62810 = v_328;
assign v_62811 = ~v_62563;
assign v_62812 = ~v_332;
assign v_62813 = v_332;
assign v_62814 = ~v_62567;
assign v_62815 = ~v_336;
assign v_62816 = v_336;
assign v_62817 = ~v_62571;
assign v_62818 = ~v_340;
assign v_62819 = v_340;
assign v_62820 = ~v_62575;
assign v_62821 = ~v_344;
assign v_62822 = v_344;
assign v_62823 = ~v_62579;
assign v_62824 = ~v_348;
assign v_62825 = v_62824;
assign v_62827 = v_62826;
assign v_62829 = v_62821 & v_62828;
assign v_62831 = v_62575;
assign v_62833 = v_62830 & v_62832;
assign v_62835 = v_62818 & v_62834;
assign v_62837 = v_62571;
assign v_62839 = v_62836 & v_62838;
assign v_62841 = v_62815 & v_62840;
assign v_62843 = v_62567;
assign v_62845 = v_62842 & v_62844;
assign v_62847 = v_62812 & v_62846;
assign v_62849 = v_62563;
assign v_62851 = v_62848 & v_62850;
assign v_62853 = v_62809 & v_62852;
assign v_62855 = v_62559;
assign v_62857 = v_62854 & v_62856;
assign v_62859 = v_62806 & v_62858;
assign v_62861 = v_62555;
assign v_62863 = v_62860 & v_62862;
assign v_62865 = v_62803 & v_62864;
assign v_62867 = v_62551;
assign v_62869 = v_62866 & v_62868;
assign v_62871 = v_62800 & v_62870;
assign v_62873 = v_62547;
assign v_62875 = v_62872 & v_62874;
assign v_62877 = v_62797 & v_62876;
assign v_62879 = v_62543;
assign v_62881 = v_62878 & v_62880;
assign v_62883 = v_62794 & v_62882;
assign v_62885 = v_62539;
assign v_62887 = v_62884 & v_62886;
assign v_62889 = v_62791 & v_62888;
assign v_62891 = v_62535;
assign v_62893 = v_62890 & v_62892;
assign v_62895 = v_62788 & v_62894;
assign v_62897 = v_62531;
assign v_62899 = v_62896 & v_62898;
assign v_62901 = v_62785 & v_62900;
assign v_62903 = v_295;
assign v_62905 = v_62902 & v_62904;
assign v_62907 = v_62782 & v_62906;
assign v_62909 = v_291;
assign v_62911 = v_62908 & v_62910;
assign v_62913 = v_62779 & v_62912;
assign v_62915 = v_287;
assign v_62917 = v_62914 & v_62916;
assign v_62919 = v_62776 & v_62918;
assign v_62921 = v_283;
assign v_62923 = v_62920 & v_62922;
assign v_62924 = v_62923;
assign v_62926 = v_62579;
assign v_62927 = v_348;
assign v_62928 = v_62927;
assign v_62929 = v_62926 & v_62928;
assign v_62930 = v_62929;
assign v_62931 = v_62821 & v_62930;
assign v_62933 = v_62831 & v_62932;
assign v_62934 = v_62820 & v_62930;
assign v_62936 = v_62818 & v_62935;
assign v_62938 = v_62837 & v_62937;
assign v_62939 = v_62817 & v_62935;
assign v_62941 = v_62815 & v_62940;
assign v_62943 = v_62843 & v_62942;
assign v_62944 = v_62814 & v_62940;
assign v_62946 = v_62812 & v_62945;
assign v_62948 = v_62849 & v_62947;
assign v_62949 = v_62811 & v_62945;
assign v_62951 = v_62809 & v_62950;
assign v_62953 = v_62855 & v_62952;
assign v_62954 = v_62808 & v_62950;
assign v_62956 = v_62806 & v_62955;
assign v_62958 = v_62861 & v_62957;
assign v_62959 = v_62805 & v_62955;
assign v_62961 = v_62803 & v_62960;
assign v_62963 = v_62867 & v_62962;
assign v_62964 = v_62802 & v_62960;
assign v_62966 = v_62800 & v_62965;
assign v_62968 = v_62873 & v_62967;
assign v_62969 = v_62799 & v_62965;
assign v_62971 = v_62797 & v_62970;
assign v_62973 = v_62879 & v_62972;
assign v_62974 = v_62796 & v_62970;
assign v_62976 = v_62794 & v_62975;
assign v_62978 = v_62885 & v_62977;
assign v_62979 = v_62793 & v_62975;
assign v_62981 = v_62791 & v_62980;
assign v_62983 = v_62891 & v_62982;
assign v_62984 = v_62790 & v_62980;
assign v_62986 = v_62788 & v_62985;
assign v_62988 = v_62897 & v_62987;
assign v_62989 = v_62787 & v_62985;
assign v_62991 = v_62785 & v_62990;
assign v_62993 = v_62903 & v_62992;
assign v_62994 = v_62784 & v_62990;
assign v_62996 = v_62782 & v_62995;
assign v_62998 = v_62909 & v_62997;
assign v_62999 = v_62781 & v_62995;
assign v_63001 = v_62779 & v_63000;
assign v_63003 = v_62915 & v_63002;
assign v_63004 = v_62778 & v_63000;
assign v_63006 = v_62776 & v_63005;
assign v_63008 = v_62921 & v_63007;
assign v_63009 = v_62775 & v_63005;
assign v_63011 = v_63010;
assign v_63013 = v_62925 & v_63012;
assign v_63014 = v_63013;
assign v_63016 = v_63015;
assign v_63018 = ~v_543;
assign v_63019 = ~v_62516;
assign v_63020 = v_62516;
assign v_63021 = ~v_547;
assign v_63022 = ~v_62520;
assign v_63023 = v_62520;
assign v_63024 = ~v_551;
assign v_63025 = ~v_62524;
assign v_63026 = v_62524;
assign v_63027 = ~v_555;
assign v_63028 = ~v_62528;
assign v_63029 = v_62528;
assign v_63030 = ~v_62531;
assign v_63031 = ~v_560;
assign v_63032 = v_560;
assign v_63033 = ~v_62535;
assign v_63034 = ~v_564;
assign v_63035 = v_564;
assign v_63036 = ~v_62539;
assign v_63037 = ~v_568;
assign v_63038 = v_568;
assign v_63039 = ~v_62543;
assign v_63040 = ~v_572;
assign v_63041 = v_572;
assign v_63042 = ~v_62547;
assign v_63043 = ~v_576;
assign v_63044 = v_576;
assign v_63045 = ~v_62551;
assign v_63046 = ~v_580;
assign v_63047 = v_580;
assign v_63048 = ~v_62555;
assign v_63049 = ~v_584;
assign v_63050 = v_584;
assign v_63051 = ~v_62559;
assign v_63052 = ~v_588;
assign v_63053 = v_588;
assign v_63054 = ~v_62563;
assign v_63055 = ~v_592;
assign v_63056 = v_592;
assign v_63057 = ~v_62567;
assign v_63058 = ~v_596;
assign v_63059 = v_596;
assign v_63060 = ~v_62571;
assign v_63061 = ~v_600;
assign v_63062 = v_600;
assign v_63063 = ~v_62575;
assign v_63064 = ~v_604;
assign v_63065 = v_604;
assign v_63066 = ~v_62579;
assign v_63067 = ~v_608;
assign v_63068 = v_63067;
assign v_63070 = v_63069;
assign v_63072 = v_63064 & v_63071;
assign v_63074 = v_62575;
assign v_63076 = v_63073 & v_63075;
assign v_63078 = v_63061 & v_63077;
assign v_63080 = v_62571;
assign v_63082 = v_63079 & v_63081;
assign v_63084 = v_63058 & v_63083;
assign v_63086 = v_62567;
assign v_63088 = v_63085 & v_63087;
assign v_63090 = v_63055 & v_63089;
assign v_63092 = v_62563;
assign v_63094 = v_63091 & v_63093;
assign v_63096 = v_63052 & v_63095;
assign v_63098 = v_62559;
assign v_63100 = v_63097 & v_63099;
assign v_63102 = v_63049 & v_63101;
assign v_63104 = v_62555;
assign v_63106 = v_63103 & v_63105;
assign v_63108 = v_63046 & v_63107;
assign v_63110 = v_62551;
assign v_63112 = v_63109 & v_63111;
assign v_63114 = v_63043 & v_63113;
assign v_63116 = v_62547;
assign v_63118 = v_63115 & v_63117;
assign v_63120 = v_63040 & v_63119;
assign v_63122 = v_62543;
assign v_63124 = v_63121 & v_63123;
assign v_63126 = v_63037 & v_63125;
assign v_63128 = v_62539;
assign v_63130 = v_63127 & v_63129;
assign v_63132 = v_63034 & v_63131;
assign v_63134 = v_62535;
assign v_63136 = v_63133 & v_63135;
assign v_63138 = v_63031 & v_63137;
assign v_63140 = v_62531;
assign v_63142 = v_63139 & v_63141;
assign v_63144 = v_63028 & v_63143;
assign v_63146 = v_555;
assign v_63148 = v_63145 & v_63147;
assign v_63150 = v_63025 & v_63149;
assign v_63152 = v_551;
assign v_63154 = v_63151 & v_63153;
assign v_63156 = v_63022 & v_63155;
assign v_63158 = v_547;
assign v_63160 = v_63157 & v_63159;
assign v_63162 = v_63019 & v_63161;
assign v_63164 = v_543;
assign v_63166 = v_63163 & v_63165;
assign v_63167 = v_63166;
assign v_63169 = v_62579;
assign v_63170 = v_608;
assign v_63171 = v_63170;
assign v_63172 = v_63169 & v_63171;
assign v_63173 = v_63172;
assign v_63174 = v_63064 & v_63173;
assign v_63176 = v_63074 & v_63175;
assign v_63177 = v_63063 & v_63173;
assign v_63179 = v_63061 & v_63178;
assign v_63181 = v_63080 & v_63180;
assign v_63182 = v_63060 & v_63178;
assign v_63184 = v_63058 & v_63183;
assign v_63186 = v_63086 & v_63185;
assign v_63187 = v_63057 & v_63183;
assign v_63189 = v_63055 & v_63188;
assign v_63191 = v_63092 & v_63190;
assign v_63192 = v_63054 & v_63188;
assign v_63194 = v_63052 & v_63193;
assign v_63196 = v_63098 & v_63195;
assign v_63197 = v_63051 & v_63193;
assign v_63199 = v_63049 & v_63198;
assign v_63201 = v_63104 & v_63200;
assign v_63202 = v_63048 & v_63198;
assign v_63204 = v_63046 & v_63203;
assign v_63206 = v_63110 & v_63205;
assign v_63207 = v_63045 & v_63203;
assign v_63209 = v_63043 & v_63208;
assign v_63211 = v_63116 & v_63210;
assign v_63212 = v_63042 & v_63208;
assign v_63214 = v_63040 & v_63213;
assign v_63216 = v_63122 & v_63215;
assign v_63217 = v_63039 & v_63213;
assign v_63219 = v_63037 & v_63218;
assign v_63221 = v_63128 & v_63220;
assign v_63222 = v_63036 & v_63218;
assign v_63224 = v_63034 & v_63223;
assign v_63226 = v_63134 & v_63225;
assign v_63227 = v_63033 & v_63223;
assign v_63229 = v_63031 & v_63228;
assign v_63231 = v_63140 & v_63230;
assign v_63232 = v_63030 & v_63228;
assign v_63234 = v_63028 & v_63233;
assign v_63236 = v_63146 & v_63235;
assign v_63237 = v_63027 & v_63233;
assign v_63239 = v_63025 & v_63238;
assign v_63241 = v_63152 & v_63240;
assign v_63242 = v_63024 & v_63238;
assign v_63244 = v_63022 & v_63243;
assign v_63246 = v_63158 & v_63245;
assign v_63247 = v_63021 & v_63243;
assign v_63249 = v_63019 & v_63248;
assign v_63251 = v_63164 & v_63250;
assign v_63252 = v_63018 & v_63248;
assign v_63254 = v_63253;
assign v_63256 = v_63168 & v_63255;
assign v_63257 = v_63256;
assign v_63259 = v_63258;
assign v_63261 = ~v_803;
assign v_63262 = ~v_62516;
assign v_63263 = v_62516;
assign v_63264 = ~v_807;
assign v_63265 = ~v_62520;
assign v_63266 = v_62520;
assign v_63267 = ~v_811;
assign v_63268 = ~v_62524;
assign v_63269 = v_62524;
assign v_63270 = ~v_815;
assign v_63271 = ~v_62528;
assign v_63272 = v_62528;
assign v_63273 = ~v_62531;
assign v_63274 = ~v_820;
assign v_63275 = v_820;
assign v_63276 = ~v_62535;
assign v_63277 = ~v_824;
assign v_63278 = v_824;
assign v_63279 = ~v_62539;
assign v_63280 = ~v_828;
assign v_63281 = v_828;
assign v_63282 = ~v_62543;
assign v_63283 = ~v_832;
assign v_63284 = v_832;
assign v_63285 = ~v_62547;
assign v_63286 = ~v_836;
assign v_63287 = v_836;
assign v_63288 = ~v_62551;
assign v_63289 = ~v_840;
assign v_63290 = v_840;
assign v_63291 = ~v_62555;
assign v_63292 = ~v_844;
assign v_63293 = v_844;
assign v_63294 = ~v_62559;
assign v_63295 = ~v_848;
assign v_63296 = v_848;
assign v_63297 = ~v_62563;
assign v_63298 = ~v_852;
assign v_63299 = v_852;
assign v_63300 = ~v_62567;
assign v_63301 = ~v_856;
assign v_63302 = v_856;
assign v_63303 = ~v_62571;
assign v_63304 = ~v_860;
assign v_63305 = v_860;
assign v_63306 = ~v_62575;
assign v_63307 = ~v_864;
assign v_63308 = v_864;
assign v_63309 = ~v_62579;
assign v_63310 = ~v_868;
assign v_63311 = v_63310;
assign v_63313 = v_63312;
assign v_63315 = v_63307 & v_63314;
assign v_63317 = v_62575;
assign v_63319 = v_63316 & v_63318;
assign v_63321 = v_63304 & v_63320;
assign v_63323 = v_62571;
assign v_63325 = v_63322 & v_63324;
assign v_63327 = v_63301 & v_63326;
assign v_63329 = v_62567;
assign v_63331 = v_63328 & v_63330;
assign v_63333 = v_63298 & v_63332;
assign v_63335 = v_62563;
assign v_63337 = v_63334 & v_63336;
assign v_63339 = v_63295 & v_63338;
assign v_63341 = v_62559;
assign v_63343 = v_63340 & v_63342;
assign v_63345 = v_63292 & v_63344;
assign v_63347 = v_62555;
assign v_63349 = v_63346 & v_63348;
assign v_63351 = v_63289 & v_63350;
assign v_63353 = v_62551;
assign v_63355 = v_63352 & v_63354;
assign v_63357 = v_63286 & v_63356;
assign v_63359 = v_62547;
assign v_63361 = v_63358 & v_63360;
assign v_63363 = v_63283 & v_63362;
assign v_63365 = v_62543;
assign v_63367 = v_63364 & v_63366;
assign v_63369 = v_63280 & v_63368;
assign v_63371 = v_62539;
assign v_63373 = v_63370 & v_63372;
assign v_63375 = v_63277 & v_63374;
assign v_63377 = v_62535;
assign v_63379 = v_63376 & v_63378;
assign v_63381 = v_63274 & v_63380;
assign v_63383 = v_62531;
assign v_63385 = v_63382 & v_63384;
assign v_63387 = v_63271 & v_63386;
assign v_63389 = v_815;
assign v_63391 = v_63388 & v_63390;
assign v_63393 = v_63268 & v_63392;
assign v_63395 = v_811;
assign v_63397 = v_63394 & v_63396;
assign v_63399 = v_63265 & v_63398;
assign v_63401 = v_807;
assign v_63403 = v_63400 & v_63402;
assign v_63405 = v_63262 & v_63404;
assign v_63407 = v_803;
assign v_63409 = v_63406 & v_63408;
assign v_63410 = v_63409;
assign v_63412 = v_62579;
assign v_63413 = v_868;
assign v_63414 = v_63413;
assign v_63415 = v_63412 & v_63414;
assign v_63416 = v_63415;
assign v_63417 = v_63307 & v_63416;
assign v_63419 = v_63317 & v_63418;
assign v_63420 = v_63306 & v_63416;
assign v_63422 = v_63304 & v_63421;
assign v_63424 = v_63323 & v_63423;
assign v_63425 = v_63303 & v_63421;
assign v_63427 = v_63301 & v_63426;
assign v_63429 = v_63329 & v_63428;
assign v_63430 = v_63300 & v_63426;
assign v_63432 = v_63298 & v_63431;
assign v_63434 = v_63335 & v_63433;
assign v_63435 = v_63297 & v_63431;
assign v_63437 = v_63295 & v_63436;
assign v_63439 = v_63341 & v_63438;
assign v_63440 = v_63294 & v_63436;
assign v_63442 = v_63292 & v_63441;
assign v_63444 = v_63347 & v_63443;
assign v_63445 = v_63291 & v_63441;
assign v_63447 = v_63289 & v_63446;
assign v_63449 = v_63353 & v_63448;
assign v_63450 = v_63288 & v_63446;
assign v_63452 = v_63286 & v_63451;
assign v_63454 = v_63359 & v_63453;
assign v_63455 = v_63285 & v_63451;
assign v_63457 = v_63283 & v_63456;
assign v_63459 = v_63365 & v_63458;
assign v_63460 = v_63282 & v_63456;
assign v_63462 = v_63280 & v_63461;
assign v_63464 = v_63371 & v_63463;
assign v_63465 = v_63279 & v_63461;
assign v_63467 = v_63277 & v_63466;
assign v_63469 = v_63377 & v_63468;
assign v_63470 = v_63276 & v_63466;
assign v_63472 = v_63274 & v_63471;
assign v_63474 = v_63383 & v_63473;
assign v_63475 = v_63273 & v_63471;
assign v_63477 = v_63271 & v_63476;
assign v_63479 = v_63389 & v_63478;
assign v_63480 = v_63270 & v_63476;
assign v_63482 = v_63268 & v_63481;
assign v_63484 = v_63395 & v_63483;
assign v_63485 = v_63267 & v_63481;
assign v_63487 = v_63265 & v_63486;
assign v_63489 = v_63401 & v_63488;
assign v_63490 = v_63264 & v_63486;
assign v_63492 = v_63262 & v_63491;
assign v_63494 = v_63407 & v_63493;
assign v_63495 = v_63261 & v_63491;
assign v_63497 = v_63496;
assign v_63499 = v_63411 & v_63498;
assign v_63500 = v_63499;
assign v_63502 = v_63501;
assign v_63504 = ~v_1063;
assign v_63505 = ~v_62516;
assign v_63506 = v_62516;
assign v_63507 = ~v_1067;
assign v_63508 = ~v_62520;
assign v_63509 = v_62520;
assign v_63510 = ~v_1071;
assign v_63511 = ~v_62524;
assign v_63512 = v_62524;
assign v_63513 = ~v_1075;
assign v_63514 = ~v_62528;
assign v_63515 = v_62528;
assign v_63516 = ~v_62531;
assign v_63517 = ~v_1080;
assign v_63518 = v_1080;
assign v_63519 = ~v_62535;
assign v_63520 = ~v_1084;
assign v_63521 = v_1084;
assign v_63522 = ~v_62539;
assign v_63523 = ~v_1088;
assign v_63524 = v_1088;
assign v_63525 = ~v_62543;
assign v_63526 = ~v_1092;
assign v_63527 = v_1092;
assign v_63528 = ~v_62547;
assign v_63529 = ~v_1096;
assign v_63530 = v_1096;
assign v_63531 = ~v_62551;
assign v_63532 = ~v_1100;
assign v_63533 = v_1100;
assign v_63534 = ~v_62555;
assign v_63535 = ~v_1104;
assign v_63536 = v_1104;
assign v_63537 = ~v_62559;
assign v_63538 = ~v_1108;
assign v_63539 = v_1108;
assign v_63540 = ~v_62563;
assign v_63541 = ~v_1112;
assign v_63542 = v_1112;
assign v_63543 = ~v_62567;
assign v_63544 = ~v_1116;
assign v_63545 = v_1116;
assign v_63546 = ~v_62571;
assign v_63547 = ~v_1120;
assign v_63548 = v_1120;
assign v_63549 = ~v_62575;
assign v_63550 = ~v_1124;
assign v_63551 = v_1124;
assign v_63552 = ~v_62579;
assign v_63553 = ~v_1128;
assign v_63554 = v_63553;
assign v_63556 = v_63555;
assign v_63558 = v_63550 & v_63557;
assign v_63560 = v_62575;
assign v_63562 = v_63559 & v_63561;
assign v_63564 = v_63547 & v_63563;
assign v_63566 = v_62571;
assign v_63568 = v_63565 & v_63567;
assign v_63570 = v_63544 & v_63569;
assign v_63572 = v_62567;
assign v_63574 = v_63571 & v_63573;
assign v_63576 = v_63541 & v_63575;
assign v_63578 = v_62563;
assign v_63580 = v_63577 & v_63579;
assign v_63582 = v_63538 & v_63581;
assign v_63584 = v_62559;
assign v_63586 = v_63583 & v_63585;
assign v_63588 = v_63535 & v_63587;
assign v_63590 = v_62555;
assign v_63592 = v_63589 & v_63591;
assign v_63594 = v_63532 & v_63593;
assign v_63596 = v_62551;
assign v_63598 = v_63595 & v_63597;
assign v_63600 = v_63529 & v_63599;
assign v_63602 = v_62547;
assign v_63604 = v_63601 & v_63603;
assign v_63606 = v_63526 & v_63605;
assign v_63608 = v_62543;
assign v_63610 = v_63607 & v_63609;
assign v_63612 = v_63523 & v_63611;
assign v_63614 = v_62539;
assign v_63616 = v_63613 & v_63615;
assign v_63618 = v_63520 & v_63617;
assign v_63620 = v_62535;
assign v_63622 = v_63619 & v_63621;
assign v_63624 = v_63517 & v_63623;
assign v_63626 = v_62531;
assign v_63628 = v_63625 & v_63627;
assign v_63630 = v_63514 & v_63629;
assign v_63632 = v_1075;
assign v_63634 = v_63631 & v_63633;
assign v_63636 = v_63511 & v_63635;
assign v_63638 = v_1071;
assign v_63640 = v_63637 & v_63639;
assign v_63642 = v_63508 & v_63641;
assign v_63644 = v_1067;
assign v_63646 = v_63643 & v_63645;
assign v_63648 = v_63505 & v_63647;
assign v_63650 = v_1063;
assign v_63652 = v_63649 & v_63651;
assign v_63653 = v_63652;
assign v_63655 = v_62579;
assign v_63656 = v_1128;
assign v_63657 = v_63656;
assign v_63658 = v_63655 & v_63657;
assign v_63659 = v_63658;
assign v_63660 = v_63550 & v_63659;
assign v_63662 = v_63560 & v_63661;
assign v_63663 = v_63549 & v_63659;
assign v_63665 = v_63547 & v_63664;
assign v_63667 = v_63566 & v_63666;
assign v_63668 = v_63546 & v_63664;
assign v_63670 = v_63544 & v_63669;
assign v_63672 = v_63572 & v_63671;
assign v_63673 = v_63543 & v_63669;
assign v_63675 = v_63541 & v_63674;
assign v_63677 = v_63578 & v_63676;
assign v_63678 = v_63540 & v_63674;
assign v_63680 = v_63538 & v_63679;
assign v_63682 = v_63584 & v_63681;
assign v_63683 = v_63537 & v_63679;
assign v_63685 = v_63535 & v_63684;
assign v_63687 = v_63590 & v_63686;
assign v_63688 = v_63534 & v_63684;
assign v_63690 = v_63532 & v_63689;
assign v_63692 = v_63596 & v_63691;
assign v_63693 = v_63531 & v_63689;
assign v_63695 = v_63529 & v_63694;
assign v_63697 = v_63602 & v_63696;
assign v_63698 = v_63528 & v_63694;
assign v_63700 = v_63526 & v_63699;
assign v_63702 = v_63608 & v_63701;
assign v_63703 = v_63525 & v_63699;
assign v_63705 = v_63523 & v_63704;
assign v_63707 = v_63614 & v_63706;
assign v_63708 = v_63522 & v_63704;
assign v_63710 = v_63520 & v_63709;
assign v_63712 = v_63620 & v_63711;
assign v_63713 = v_63519 & v_63709;
assign v_63715 = v_63517 & v_63714;
assign v_63717 = v_63626 & v_63716;
assign v_63718 = v_63516 & v_63714;
assign v_63720 = v_63514 & v_63719;
assign v_63722 = v_63632 & v_63721;
assign v_63723 = v_63513 & v_63719;
assign v_63725 = v_63511 & v_63724;
assign v_63727 = v_63638 & v_63726;
assign v_63728 = v_63510 & v_63724;
assign v_63730 = v_63508 & v_63729;
assign v_63732 = v_63644 & v_63731;
assign v_63733 = v_63507 & v_63729;
assign v_63735 = v_63505 & v_63734;
assign v_63737 = v_63650 & v_63736;
assign v_63738 = v_63504 & v_63734;
assign v_63740 = v_63739;
assign v_63742 = v_63654 & v_63741;
assign v_63743 = v_63742;
assign v_63745 = v_63744;
assign v_63747 = ~v_1323;
assign v_63748 = ~v_62516;
assign v_63749 = v_62516;
assign v_63750 = ~v_1327;
assign v_63751 = ~v_62520;
assign v_63752 = v_62520;
assign v_63753 = ~v_1331;
assign v_63754 = ~v_62524;
assign v_63755 = v_62524;
assign v_63756 = ~v_1335;
assign v_63757 = ~v_62528;
assign v_63758 = v_62528;
assign v_63759 = ~v_62531;
assign v_63760 = ~v_1340;
assign v_63761 = v_1340;
assign v_63762 = ~v_62535;
assign v_63763 = ~v_1344;
assign v_63764 = v_1344;
assign v_63765 = ~v_62539;
assign v_63766 = ~v_1348;
assign v_63767 = v_1348;
assign v_63768 = ~v_62543;
assign v_63769 = ~v_1352;
assign v_63770 = v_1352;
assign v_63771 = ~v_62547;
assign v_63772 = ~v_1356;
assign v_63773 = v_1356;
assign v_63774 = ~v_62551;
assign v_63775 = ~v_1360;
assign v_63776 = v_1360;
assign v_63777 = ~v_62555;
assign v_63778 = ~v_1364;
assign v_63779 = v_1364;
assign v_63780 = ~v_62559;
assign v_63781 = ~v_1368;
assign v_63782 = v_1368;
assign v_63783 = ~v_62563;
assign v_63784 = ~v_1372;
assign v_63785 = v_1372;
assign v_63786 = ~v_62567;
assign v_63787 = ~v_1376;
assign v_63788 = v_1376;
assign v_63789 = ~v_62571;
assign v_63790 = ~v_1380;
assign v_63791 = v_1380;
assign v_63792 = ~v_62575;
assign v_63793 = ~v_1384;
assign v_63794 = v_1384;
assign v_63795 = ~v_62579;
assign v_63796 = ~v_1388;
assign v_63797 = v_63796;
assign v_63799 = v_63798;
assign v_63801 = v_63793 & v_63800;
assign v_63803 = v_62575;
assign v_63805 = v_63802 & v_63804;
assign v_63807 = v_63790 & v_63806;
assign v_63809 = v_62571;
assign v_63811 = v_63808 & v_63810;
assign v_63813 = v_63787 & v_63812;
assign v_63815 = v_62567;
assign v_63817 = v_63814 & v_63816;
assign v_63819 = v_63784 & v_63818;
assign v_63821 = v_62563;
assign v_63823 = v_63820 & v_63822;
assign v_63825 = v_63781 & v_63824;
assign v_63827 = v_62559;
assign v_63829 = v_63826 & v_63828;
assign v_63831 = v_63778 & v_63830;
assign v_63833 = v_62555;
assign v_63835 = v_63832 & v_63834;
assign v_63837 = v_63775 & v_63836;
assign v_63839 = v_62551;
assign v_63841 = v_63838 & v_63840;
assign v_63843 = v_63772 & v_63842;
assign v_63845 = v_62547;
assign v_63847 = v_63844 & v_63846;
assign v_63849 = v_63769 & v_63848;
assign v_63851 = v_62543;
assign v_63853 = v_63850 & v_63852;
assign v_63855 = v_63766 & v_63854;
assign v_63857 = v_62539;
assign v_63859 = v_63856 & v_63858;
assign v_63861 = v_63763 & v_63860;
assign v_63863 = v_62535;
assign v_63865 = v_63862 & v_63864;
assign v_63867 = v_63760 & v_63866;
assign v_63869 = v_62531;
assign v_63871 = v_63868 & v_63870;
assign v_63873 = v_63757 & v_63872;
assign v_63875 = v_1335;
assign v_63877 = v_63874 & v_63876;
assign v_63879 = v_63754 & v_63878;
assign v_63881 = v_1331;
assign v_63883 = v_63880 & v_63882;
assign v_63885 = v_63751 & v_63884;
assign v_63887 = v_1327;
assign v_63889 = v_63886 & v_63888;
assign v_63891 = v_63748 & v_63890;
assign v_63893 = v_1323;
assign v_63895 = v_63892 & v_63894;
assign v_63896 = v_63895;
assign v_63898 = v_62579;
assign v_63899 = v_1388;
assign v_63900 = v_63899;
assign v_63901 = v_63898 & v_63900;
assign v_63902 = v_63901;
assign v_63903 = v_63793 & v_63902;
assign v_63905 = v_63803 & v_63904;
assign v_63906 = v_63792 & v_63902;
assign v_63908 = v_63790 & v_63907;
assign v_63910 = v_63809 & v_63909;
assign v_63911 = v_63789 & v_63907;
assign v_63913 = v_63787 & v_63912;
assign v_63915 = v_63815 & v_63914;
assign v_63916 = v_63786 & v_63912;
assign v_63918 = v_63784 & v_63917;
assign v_63920 = v_63821 & v_63919;
assign v_63921 = v_63783 & v_63917;
assign v_63923 = v_63781 & v_63922;
assign v_63925 = v_63827 & v_63924;
assign v_63926 = v_63780 & v_63922;
assign v_63928 = v_63778 & v_63927;
assign v_63930 = v_63833 & v_63929;
assign v_63931 = v_63777 & v_63927;
assign v_63933 = v_63775 & v_63932;
assign v_63935 = v_63839 & v_63934;
assign v_63936 = v_63774 & v_63932;
assign v_63938 = v_63772 & v_63937;
assign v_63940 = v_63845 & v_63939;
assign v_63941 = v_63771 & v_63937;
assign v_63943 = v_63769 & v_63942;
assign v_63945 = v_63851 & v_63944;
assign v_63946 = v_63768 & v_63942;
assign v_63948 = v_63766 & v_63947;
assign v_63950 = v_63857 & v_63949;
assign v_63951 = v_63765 & v_63947;
assign v_63953 = v_63763 & v_63952;
assign v_63955 = v_63863 & v_63954;
assign v_63956 = v_63762 & v_63952;
assign v_63958 = v_63760 & v_63957;
assign v_63960 = v_63869 & v_63959;
assign v_63961 = v_63759 & v_63957;
assign v_63963 = v_63757 & v_63962;
assign v_63965 = v_63875 & v_63964;
assign v_63966 = v_63756 & v_63962;
assign v_63968 = v_63754 & v_63967;
assign v_63970 = v_63881 & v_63969;
assign v_63971 = v_63753 & v_63967;
assign v_63973 = v_63751 & v_63972;
assign v_63975 = v_63887 & v_63974;
assign v_63976 = v_63750 & v_63972;
assign v_63978 = v_63748 & v_63977;
assign v_63980 = v_63893 & v_63979;
assign v_63981 = v_63747 & v_63977;
assign v_63983 = v_63982;
assign v_63985 = v_63897 & v_63984;
assign v_63986 = v_63985;
assign v_63988 = v_63987;
assign v_63990 = ~v_1583;
assign v_63991 = ~v_62516;
assign v_63992 = v_62516;
assign v_63993 = ~v_1587;
assign v_63994 = ~v_62520;
assign v_63995 = v_62520;
assign v_63996 = ~v_1591;
assign v_63997 = ~v_62524;
assign v_63998 = v_62524;
assign v_63999 = ~v_1595;
assign v_64000 = ~v_62528;
assign v_64001 = v_62528;
assign v_64002 = ~v_62531;
assign v_64003 = ~v_1600;
assign v_64004 = v_1600;
assign v_64005 = ~v_62535;
assign v_64006 = ~v_1604;
assign v_64007 = v_1604;
assign v_64008 = ~v_62539;
assign v_64009 = ~v_1608;
assign v_64010 = v_1608;
assign v_64011 = ~v_62543;
assign v_64012 = ~v_1612;
assign v_64013 = v_1612;
assign v_64014 = ~v_62547;
assign v_64015 = ~v_1616;
assign v_64016 = v_1616;
assign v_64017 = ~v_62551;
assign v_64018 = ~v_1620;
assign v_64019 = v_1620;
assign v_64020 = ~v_62555;
assign v_64021 = ~v_1624;
assign v_64022 = v_1624;
assign v_64023 = ~v_62559;
assign v_64024 = ~v_1628;
assign v_64025 = v_1628;
assign v_64026 = ~v_62563;
assign v_64027 = ~v_1632;
assign v_64028 = v_1632;
assign v_64029 = ~v_62567;
assign v_64030 = ~v_1636;
assign v_64031 = v_1636;
assign v_64032 = ~v_62571;
assign v_64033 = ~v_1640;
assign v_64034 = v_1640;
assign v_64035 = ~v_62575;
assign v_64036 = ~v_1644;
assign v_64037 = v_1644;
assign v_64038 = ~v_62579;
assign v_64039 = ~v_1648;
assign v_64040 = v_64039;
assign v_64042 = v_64041;
assign v_64044 = v_64036 & v_64043;
assign v_64046 = v_62575;
assign v_64048 = v_64045 & v_64047;
assign v_64050 = v_64033 & v_64049;
assign v_64052 = v_62571;
assign v_64054 = v_64051 & v_64053;
assign v_64056 = v_64030 & v_64055;
assign v_64058 = v_62567;
assign v_64060 = v_64057 & v_64059;
assign v_64062 = v_64027 & v_64061;
assign v_64064 = v_62563;
assign v_64066 = v_64063 & v_64065;
assign v_64068 = v_64024 & v_64067;
assign v_64070 = v_62559;
assign v_64072 = v_64069 & v_64071;
assign v_64074 = v_64021 & v_64073;
assign v_64076 = v_62555;
assign v_64078 = v_64075 & v_64077;
assign v_64080 = v_64018 & v_64079;
assign v_64082 = v_62551;
assign v_64084 = v_64081 & v_64083;
assign v_64086 = v_64015 & v_64085;
assign v_64088 = v_62547;
assign v_64090 = v_64087 & v_64089;
assign v_64092 = v_64012 & v_64091;
assign v_64094 = v_62543;
assign v_64096 = v_64093 & v_64095;
assign v_64098 = v_64009 & v_64097;
assign v_64100 = v_62539;
assign v_64102 = v_64099 & v_64101;
assign v_64104 = v_64006 & v_64103;
assign v_64106 = v_62535;
assign v_64108 = v_64105 & v_64107;
assign v_64110 = v_64003 & v_64109;
assign v_64112 = v_62531;
assign v_64114 = v_64111 & v_64113;
assign v_64116 = v_64000 & v_64115;
assign v_64118 = v_1595;
assign v_64120 = v_64117 & v_64119;
assign v_64122 = v_63997 & v_64121;
assign v_64124 = v_1591;
assign v_64126 = v_64123 & v_64125;
assign v_64128 = v_63994 & v_64127;
assign v_64130 = v_1587;
assign v_64132 = v_64129 & v_64131;
assign v_64134 = v_63991 & v_64133;
assign v_64136 = v_1583;
assign v_64138 = v_64135 & v_64137;
assign v_64139 = v_64138;
assign v_64141 = v_62579;
assign v_64142 = v_1648;
assign v_64143 = v_64142;
assign v_64144 = v_64141 & v_64143;
assign v_64145 = v_64144;
assign v_64146 = v_64036 & v_64145;
assign v_64148 = v_64046 & v_64147;
assign v_64149 = v_64035 & v_64145;
assign v_64151 = v_64033 & v_64150;
assign v_64153 = v_64052 & v_64152;
assign v_64154 = v_64032 & v_64150;
assign v_64156 = v_64030 & v_64155;
assign v_64158 = v_64058 & v_64157;
assign v_64159 = v_64029 & v_64155;
assign v_64161 = v_64027 & v_64160;
assign v_64163 = v_64064 & v_64162;
assign v_64164 = v_64026 & v_64160;
assign v_64166 = v_64024 & v_64165;
assign v_64168 = v_64070 & v_64167;
assign v_64169 = v_64023 & v_64165;
assign v_64171 = v_64021 & v_64170;
assign v_64173 = v_64076 & v_64172;
assign v_64174 = v_64020 & v_64170;
assign v_64176 = v_64018 & v_64175;
assign v_64178 = v_64082 & v_64177;
assign v_64179 = v_64017 & v_64175;
assign v_64181 = v_64015 & v_64180;
assign v_64183 = v_64088 & v_64182;
assign v_64184 = v_64014 & v_64180;
assign v_64186 = v_64012 & v_64185;
assign v_64188 = v_64094 & v_64187;
assign v_64189 = v_64011 & v_64185;
assign v_64191 = v_64009 & v_64190;
assign v_64193 = v_64100 & v_64192;
assign v_64194 = v_64008 & v_64190;
assign v_64196 = v_64006 & v_64195;
assign v_64198 = v_64106 & v_64197;
assign v_64199 = v_64005 & v_64195;
assign v_64201 = v_64003 & v_64200;
assign v_64203 = v_64112 & v_64202;
assign v_64204 = v_64002 & v_64200;
assign v_64206 = v_64000 & v_64205;
assign v_64208 = v_64118 & v_64207;
assign v_64209 = v_63999 & v_64205;
assign v_64211 = v_63997 & v_64210;
assign v_64213 = v_64124 & v_64212;
assign v_64214 = v_63996 & v_64210;
assign v_64216 = v_63994 & v_64215;
assign v_64218 = v_64130 & v_64217;
assign v_64219 = v_63993 & v_64215;
assign v_64221 = v_63991 & v_64220;
assign v_64223 = v_64136 & v_64222;
assign v_64224 = v_63990 & v_64220;
assign v_64226 = v_64225;
assign v_64228 = v_64140 & v_64227;
assign v_64229 = v_64228;
assign v_64231 = v_64230;
assign v_64233 = ~v_1843;
assign v_64234 = ~v_62516;
assign v_64235 = v_62516;
assign v_64236 = ~v_1847;
assign v_64237 = ~v_62520;
assign v_64238 = v_62520;
assign v_64239 = ~v_1851;
assign v_64240 = ~v_62524;
assign v_64241 = v_62524;
assign v_64242 = ~v_1855;
assign v_64243 = ~v_62528;
assign v_64244 = v_62528;
assign v_64245 = ~v_62531;
assign v_64246 = ~v_1860;
assign v_64247 = v_1860;
assign v_64248 = ~v_62535;
assign v_64249 = ~v_1864;
assign v_64250 = v_1864;
assign v_64251 = ~v_62539;
assign v_64252 = ~v_1868;
assign v_64253 = v_1868;
assign v_64254 = ~v_62543;
assign v_64255 = ~v_1872;
assign v_64256 = v_1872;
assign v_64257 = ~v_62547;
assign v_64258 = ~v_1876;
assign v_64259 = v_1876;
assign v_64260 = ~v_62551;
assign v_64261 = ~v_1880;
assign v_64262 = v_1880;
assign v_64263 = ~v_62555;
assign v_64264 = ~v_1884;
assign v_64265 = v_1884;
assign v_64266 = ~v_62559;
assign v_64267 = ~v_1888;
assign v_64268 = v_1888;
assign v_64269 = ~v_62563;
assign v_64270 = ~v_1892;
assign v_64271 = v_1892;
assign v_64272 = ~v_62567;
assign v_64273 = ~v_1896;
assign v_64274 = v_1896;
assign v_64275 = ~v_62571;
assign v_64276 = ~v_1900;
assign v_64277 = v_1900;
assign v_64278 = ~v_62575;
assign v_64279 = ~v_1904;
assign v_64280 = v_1904;
assign v_64281 = ~v_62579;
assign v_64282 = ~v_1908;
assign v_64283 = v_64282;
assign v_64285 = v_64284;
assign v_64287 = v_64279 & v_64286;
assign v_64289 = v_62575;
assign v_64291 = v_64288 & v_64290;
assign v_64293 = v_64276 & v_64292;
assign v_64295 = v_62571;
assign v_64297 = v_64294 & v_64296;
assign v_64299 = v_64273 & v_64298;
assign v_64301 = v_62567;
assign v_64303 = v_64300 & v_64302;
assign v_64305 = v_64270 & v_64304;
assign v_64307 = v_62563;
assign v_64309 = v_64306 & v_64308;
assign v_64311 = v_64267 & v_64310;
assign v_64313 = v_62559;
assign v_64315 = v_64312 & v_64314;
assign v_64317 = v_64264 & v_64316;
assign v_64319 = v_62555;
assign v_64321 = v_64318 & v_64320;
assign v_64323 = v_64261 & v_64322;
assign v_64325 = v_62551;
assign v_64327 = v_64324 & v_64326;
assign v_64329 = v_64258 & v_64328;
assign v_64331 = v_62547;
assign v_64333 = v_64330 & v_64332;
assign v_64335 = v_64255 & v_64334;
assign v_64337 = v_62543;
assign v_64339 = v_64336 & v_64338;
assign v_64341 = v_64252 & v_64340;
assign v_64343 = v_62539;
assign v_64345 = v_64342 & v_64344;
assign v_64347 = v_64249 & v_64346;
assign v_64349 = v_62535;
assign v_64351 = v_64348 & v_64350;
assign v_64353 = v_64246 & v_64352;
assign v_64355 = v_62531;
assign v_64357 = v_64354 & v_64356;
assign v_64359 = v_64243 & v_64358;
assign v_64361 = v_1855;
assign v_64363 = v_64360 & v_64362;
assign v_64365 = v_64240 & v_64364;
assign v_64367 = v_1851;
assign v_64369 = v_64366 & v_64368;
assign v_64371 = v_64237 & v_64370;
assign v_64373 = v_1847;
assign v_64375 = v_64372 & v_64374;
assign v_64377 = v_64234 & v_64376;
assign v_64379 = v_1843;
assign v_64381 = v_64378 & v_64380;
assign v_64382 = v_64381;
assign v_64384 = v_62579;
assign v_64385 = v_1908;
assign v_64386 = v_64385;
assign v_64387 = v_64384 & v_64386;
assign v_64388 = v_64387;
assign v_64389 = v_64279 & v_64388;
assign v_64391 = v_64289 & v_64390;
assign v_64392 = v_64278 & v_64388;
assign v_64394 = v_64276 & v_64393;
assign v_64396 = v_64295 & v_64395;
assign v_64397 = v_64275 & v_64393;
assign v_64399 = v_64273 & v_64398;
assign v_64401 = v_64301 & v_64400;
assign v_64402 = v_64272 & v_64398;
assign v_64404 = v_64270 & v_64403;
assign v_64406 = v_64307 & v_64405;
assign v_64407 = v_64269 & v_64403;
assign v_64409 = v_64267 & v_64408;
assign v_64411 = v_64313 & v_64410;
assign v_64412 = v_64266 & v_64408;
assign v_64414 = v_64264 & v_64413;
assign v_64416 = v_64319 & v_64415;
assign v_64417 = v_64263 & v_64413;
assign v_64419 = v_64261 & v_64418;
assign v_64421 = v_64325 & v_64420;
assign v_64422 = v_64260 & v_64418;
assign v_64424 = v_64258 & v_64423;
assign v_64426 = v_64331 & v_64425;
assign v_64427 = v_64257 & v_64423;
assign v_64429 = v_64255 & v_64428;
assign v_64431 = v_64337 & v_64430;
assign v_64432 = v_64254 & v_64428;
assign v_64434 = v_64252 & v_64433;
assign v_64436 = v_64343 & v_64435;
assign v_64437 = v_64251 & v_64433;
assign v_64439 = v_64249 & v_64438;
assign v_64441 = v_64349 & v_64440;
assign v_64442 = v_64248 & v_64438;
assign v_64444 = v_64246 & v_64443;
assign v_64446 = v_64355 & v_64445;
assign v_64447 = v_64245 & v_64443;
assign v_64449 = v_64243 & v_64448;
assign v_64451 = v_64361 & v_64450;
assign v_64452 = v_64242 & v_64448;
assign v_64454 = v_64240 & v_64453;
assign v_64456 = v_64367 & v_64455;
assign v_64457 = v_64239 & v_64453;
assign v_64459 = v_64237 & v_64458;
assign v_64461 = v_64373 & v_64460;
assign v_64462 = v_64236 & v_64458;
assign v_64464 = v_64234 & v_64463;
assign v_64466 = v_64379 & v_64465;
assign v_64467 = v_64233 & v_64463;
assign v_64469 = v_64468;
assign v_64471 = v_64383 & v_64470;
assign v_64472 = v_64471;
assign v_64474 = v_64473;
assign v_64476 = ~v_2103;
assign v_64477 = ~v_62516;
assign v_64478 = v_62516;
assign v_64479 = ~v_2107;
assign v_64480 = ~v_62520;
assign v_64481 = v_62520;
assign v_64482 = ~v_2111;
assign v_64483 = ~v_62524;
assign v_64484 = v_62524;
assign v_64485 = ~v_2115;
assign v_64486 = ~v_62528;
assign v_64487 = v_62528;
assign v_64488 = ~v_62531;
assign v_64489 = ~v_2120;
assign v_64490 = v_2120;
assign v_64491 = ~v_62535;
assign v_64492 = ~v_2124;
assign v_64493 = v_2124;
assign v_64494 = ~v_62539;
assign v_64495 = ~v_2128;
assign v_64496 = v_2128;
assign v_64497 = ~v_62543;
assign v_64498 = ~v_2132;
assign v_64499 = v_2132;
assign v_64500 = ~v_62547;
assign v_64501 = ~v_2136;
assign v_64502 = v_2136;
assign v_64503 = ~v_62551;
assign v_64504 = ~v_2140;
assign v_64505 = v_2140;
assign v_64506 = ~v_62555;
assign v_64507 = ~v_2144;
assign v_64508 = v_2144;
assign v_64509 = ~v_62559;
assign v_64510 = ~v_2148;
assign v_64511 = v_2148;
assign v_64512 = ~v_62563;
assign v_64513 = ~v_2152;
assign v_64514 = v_2152;
assign v_64515 = ~v_62567;
assign v_64516 = ~v_2156;
assign v_64517 = v_2156;
assign v_64518 = ~v_62571;
assign v_64519 = ~v_2160;
assign v_64520 = v_2160;
assign v_64521 = ~v_62575;
assign v_64522 = ~v_2164;
assign v_64523 = v_2164;
assign v_64524 = ~v_62579;
assign v_64525 = ~v_2168;
assign v_64526 = v_64525;
assign v_64528 = v_64527;
assign v_64530 = v_64522 & v_64529;
assign v_64532 = v_62575;
assign v_64534 = v_64531 & v_64533;
assign v_64536 = v_64519 & v_64535;
assign v_64538 = v_62571;
assign v_64540 = v_64537 & v_64539;
assign v_64542 = v_64516 & v_64541;
assign v_64544 = v_62567;
assign v_64546 = v_64543 & v_64545;
assign v_64548 = v_64513 & v_64547;
assign v_64550 = v_62563;
assign v_64552 = v_64549 & v_64551;
assign v_64554 = v_64510 & v_64553;
assign v_64556 = v_62559;
assign v_64558 = v_64555 & v_64557;
assign v_64560 = v_64507 & v_64559;
assign v_64562 = v_62555;
assign v_64564 = v_64561 & v_64563;
assign v_64566 = v_64504 & v_64565;
assign v_64568 = v_62551;
assign v_64570 = v_64567 & v_64569;
assign v_64572 = v_64501 & v_64571;
assign v_64574 = v_62547;
assign v_64576 = v_64573 & v_64575;
assign v_64578 = v_64498 & v_64577;
assign v_64580 = v_62543;
assign v_64582 = v_64579 & v_64581;
assign v_64584 = v_64495 & v_64583;
assign v_64586 = v_62539;
assign v_64588 = v_64585 & v_64587;
assign v_64590 = v_64492 & v_64589;
assign v_64592 = v_62535;
assign v_64594 = v_64591 & v_64593;
assign v_64596 = v_64489 & v_64595;
assign v_64598 = v_62531;
assign v_64600 = v_64597 & v_64599;
assign v_64602 = v_64486 & v_64601;
assign v_64604 = v_2115;
assign v_64606 = v_64603 & v_64605;
assign v_64608 = v_64483 & v_64607;
assign v_64610 = v_2111;
assign v_64612 = v_64609 & v_64611;
assign v_64614 = v_64480 & v_64613;
assign v_64616 = v_2107;
assign v_64618 = v_64615 & v_64617;
assign v_64620 = v_64477 & v_64619;
assign v_64622 = v_2103;
assign v_64624 = v_64621 & v_64623;
assign v_64625 = v_64624;
assign v_64627 = v_62579;
assign v_64628 = v_2168;
assign v_64629 = v_64628;
assign v_64630 = v_64627 & v_64629;
assign v_64631 = v_64630;
assign v_64632 = v_64522 & v_64631;
assign v_64634 = v_64532 & v_64633;
assign v_64635 = v_64521 & v_64631;
assign v_64637 = v_64519 & v_64636;
assign v_64639 = v_64538 & v_64638;
assign v_64640 = v_64518 & v_64636;
assign v_64642 = v_64516 & v_64641;
assign v_64644 = v_64544 & v_64643;
assign v_64645 = v_64515 & v_64641;
assign v_64647 = v_64513 & v_64646;
assign v_64649 = v_64550 & v_64648;
assign v_64650 = v_64512 & v_64646;
assign v_64652 = v_64510 & v_64651;
assign v_64654 = v_64556 & v_64653;
assign v_64655 = v_64509 & v_64651;
assign v_64657 = v_64507 & v_64656;
assign v_64659 = v_64562 & v_64658;
assign v_64660 = v_64506 & v_64656;
assign v_64662 = v_64504 & v_64661;
assign v_64664 = v_64568 & v_64663;
assign v_64665 = v_64503 & v_64661;
assign v_64667 = v_64501 & v_64666;
assign v_64669 = v_64574 & v_64668;
assign v_64670 = v_64500 & v_64666;
assign v_64672 = v_64498 & v_64671;
assign v_64674 = v_64580 & v_64673;
assign v_64675 = v_64497 & v_64671;
assign v_64677 = v_64495 & v_64676;
assign v_64679 = v_64586 & v_64678;
assign v_64680 = v_64494 & v_64676;
assign v_64682 = v_64492 & v_64681;
assign v_64684 = v_64592 & v_64683;
assign v_64685 = v_64491 & v_64681;
assign v_64687 = v_64489 & v_64686;
assign v_64689 = v_64598 & v_64688;
assign v_64690 = v_64488 & v_64686;
assign v_64692 = v_64486 & v_64691;
assign v_64694 = v_64604 & v_64693;
assign v_64695 = v_64485 & v_64691;
assign v_64697 = v_64483 & v_64696;
assign v_64699 = v_64610 & v_64698;
assign v_64700 = v_64482 & v_64696;
assign v_64702 = v_64480 & v_64701;
assign v_64704 = v_64616 & v_64703;
assign v_64705 = v_64479 & v_64701;
assign v_64707 = v_64477 & v_64706;
assign v_64709 = v_64622 & v_64708;
assign v_64710 = v_64476 & v_64706;
assign v_64712 = v_64711;
assign v_64714 = v_64626 & v_64713;
assign v_64715 = v_64714;
assign v_64717 = v_64716;
assign v_64719 = ~v_2363;
assign v_64720 = ~v_62516;
assign v_64721 = v_62516;
assign v_64722 = ~v_2367;
assign v_64723 = ~v_62520;
assign v_64724 = v_62520;
assign v_64725 = ~v_2371;
assign v_64726 = ~v_62524;
assign v_64727 = v_62524;
assign v_64728 = ~v_2375;
assign v_64729 = ~v_62528;
assign v_64730 = v_62528;
assign v_64731 = ~v_62531;
assign v_64732 = ~v_2380;
assign v_64733 = v_2380;
assign v_64734 = ~v_62535;
assign v_64735 = ~v_2384;
assign v_64736 = v_2384;
assign v_64737 = ~v_62539;
assign v_64738 = ~v_2388;
assign v_64739 = v_2388;
assign v_64740 = ~v_62543;
assign v_64741 = ~v_2392;
assign v_64742 = v_2392;
assign v_64743 = ~v_62547;
assign v_64744 = ~v_2396;
assign v_64745 = v_2396;
assign v_64746 = ~v_62551;
assign v_64747 = ~v_2400;
assign v_64748 = v_2400;
assign v_64749 = ~v_62555;
assign v_64750 = ~v_2404;
assign v_64751 = v_2404;
assign v_64752 = ~v_62559;
assign v_64753 = ~v_2408;
assign v_64754 = v_2408;
assign v_64755 = ~v_62563;
assign v_64756 = ~v_2412;
assign v_64757 = v_2412;
assign v_64758 = ~v_62567;
assign v_64759 = ~v_2416;
assign v_64760 = v_2416;
assign v_64761 = ~v_62571;
assign v_64762 = ~v_2420;
assign v_64763 = v_2420;
assign v_64764 = ~v_62575;
assign v_64765 = ~v_2424;
assign v_64766 = v_2424;
assign v_64767 = ~v_62579;
assign v_64768 = ~v_2428;
assign v_64769 = v_64768;
assign v_64771 = v_64770;
assign v_64773 = v_64765 & v_64772;
assign v_64775 = v_62575;
assign v_64777 = v_64774 & v_64776;
assign v_64779 = v_64762 & v_64778;
assign v_64781 = v_62571;
assign v_64783 = v_64780 & v_64782;
assign v_64785 = v_64759 & v_64784;
assign v_64787 = v_62567;
assign v_64789 = v_64786 & v_64788;
assign v_64791 = v_64756 & v_64790;
assign v_64793 = v_62563;
assign v_64795 = v_64792 & v_64794;
assign v_64797 = v_64753 & v_64796;
assign v_64799 = v_62559;
assign v_64801 = v_64798 & v_64800;
assign v_64803 = v_64750 & v_64802;
assign v_64805 = v_62555;
assign v_64807 = v_64804 & v_64806;
assign v_64809 = v_64747 & v_64808;
assign v_64811 = v_62551;
assign v_64813 = v_64810 & v_64812;
assign v_64815 = v_64744 & v_64814;
assign v_64817 = v_62547;
assign v_64819 = v_64816 & v_64818;
assign v_64821 = v_64741 & v_64820;
assign v_64823 = v_62543;
assign v_64825 = v_64822 & v_64824;
assign v_64827 = v_64738 & v_64826;
assign v_64829 = v_62539;
assign v_64831 = v_64828 & v_64830;
assign v_64833 = v_64735 & v_64832;
assign v_64835 = v_62535;
assign v_64837 = v_64834 & v_64836;
assign v_64839 = v_64732 & v_64838;
assign v_64841 = v_62531;
assign v_64843 = v_64840 & v_64842;
assign v_64845 = v_64729 & v_64844;
assign v_64847 = v_2375;
assign v_64849 = v_64846 & v_64848;
assign v_64851 = v_64726 & v_64850;
assign v_64853 = v_2371;
assign v_64855 = v_64852 & v_64854;
assign v_64857 = v_64723 & v_64856;
assign v_64859 = v_2367;
assign v_64861 = v_64858 & v_64860;
assign v_64863 = v_64720 & v_64862;
assign v_64865 = v_2363;
assign v_64867 = v_64864 & v_64866;
assign v_64868 = v_64867;
assign v_64870 = v_62579;
assign v_64871 = v_2428;
assign v_64872 = v_64871;
assign v_64873 = v_64870 & v_64872;
assign v_64874 = v_64873;
assign v_64875 = v_64765 & v_64874;
assign v_64877 = v_64775 & v_64876;
assign v_64878 = v_64764 & v_64874;
assign v_64880 = v_64762 & v_64879;
assign v_64882 = v_64781 & v_64881;
assign v_64883 = v_64761 & v_64879;
assign v_64885 = v_64759 & v_64884;
assign v_64887 = v_64787 & v_64886;
assign v_64888 = v_64758 & v_64884;
assign v_64890 = v_64756 & v_64889;
assign v_64892 = v_64793 & v_64891;
assign v_64893 = v_64755 & v_64889;
assign v_64895 = v_64753 & v_64894;
assign v_64897 = v_64799 & v_64896;
assign v_64898 = v_64752 & v_64894;
assign v_64900 = v_64750 & v_64899;
assign v_64902 = v_64805 & v_64901;
assign v_64903 = v_64749 & v_64899;
assign v_64905 = v_64747 & v_64904;
assign v_64907 = v_64811 & v_64906;
assign v_64908 = v_64746 & v_64904;
assign v_64910 = v_64744 & v_64909;
assign v_64912 = v_64817 & v_64911;
assign v_64913 = v_64743 & v_64909;
assign v_64915 = v_64741 & v_64914;
assign v_64917 = v_64823 & v_64916;
assign v_64918 = v_64740 & v_64914;
assign v_64920 = v_64738 & v_64919;
assign v_64922 = v_64829 & v_64921;
assign v_64923 = v_64737 & v_64919;
assign v_64925 = v_64735 & v_64924;
assign v_64927 = v_64835 & v_64926;
assign v_64928 = v_64734 & v_64924;
assign v_64930 = v_64732 & v_64929;
assign v_64932 = v_64841 & v_64931;
assign v_64933 = v_64731 & v_64929;
assign v_64935 = v_64729 & v_64934;
assign v_64937 = v_64847 & v_64936;
assign v_64938 = v_64728 & v_64934;
assign v_64940 = v_64726 & v_64939;
assign v_64942 = v_64853 & v_64941;
assign v_64943 = v_64725 & v_64939;
assign v_64945 = v_64723 & v_64944;
assign v_64947 = v_64859 & v_64946;
assign v_64948 = v_64722 & v_64944;
assign v_64950 = v_64720 & v_64949;
assign v_64952 = v_64865 & v_64951;
assign v_64953 = v_64719 & v_64949;
assign v_64955 = v_64954;
assign v_64957 = v_64869 & v_64956;
assign v_64958 = v_64957;
assign v_64960 = v_64959;
assign v_64962 = ~v_2623;
assign v_64963 = ~v_62516;
assign v_64964 = v_62516;
assign v_64965 = ~v_2627;
assign v_64966 = ~v_62520;
assign v_64967 = v_62520;
assign v_64968 = ~v_2631;
assign v_64969 = ~v_62524;
assign v_64970 = v_62524;
assign v_64971 = ~v_2635;
assign v_64972 = ~v_62528;
assign v_64973 = v_62528;
assign v_64974 = ~v_62531;
assign v_64975 = ~v_2640;
assign v_64976 = v_2640;
assign v_64977 = ~v_62535;
assign v_64978 = ~v_2644;
assign v_64979 = v_2644;
assign v_64980 = ~v_62539;
assign v_64981 = ~v_2648;
assign v_64982 = v_2648;
assign v_64983 = ~v_62543;
assign v_64984 = ~v_2652;
assign v_64985 = v_2652;
assign v_64986 = ~v_62547;
assign v_64987 = ~v_2656;
assign v_64988 = v_2656;
assign v_64989 = ~v_62551;
assign v_64990 = ~v_2660;
assign v_64991 = v_2660;
assign v_64992 = ~v_62555;
assign v_64993 = ~v_2664;
assign v_64994 = v_2664;
assign v_64995 = ~v_62559;
assign v_64996 = ~v_2668;
assign v_64997 = v_2668;
assign v_64998 = ~v_62563;
assign v_64999 = ~v_2672;
assign v_65000 = v_2672;
assign v_65001 = ~v_62567;
assign v_65002 = ~v_2676;
assign v_65003 = v_2676;
assign v_65004 = ~v_62571;
assign v_65005 = ~v_2680;
assign v_65006 = v_2680;
assign v_65007 = ~v_62575;
assign v_65008 = ~v_2684;
assign v_65009 = v_2684;
assign v_65010 = ~v_62579;
assign v_65011 = ~v_2688;
assign v_65012 = v_65011;
assign v_65014 = v_65013;
assign v_65016 = v_65008 & v_65015;
assign v_65018 = v_62575;
assign v_65020 = v_65017 & v_65019;
assign v_65022 = v_65005 & v_65021;
assign v_65024 = v_62571;
assign v_65026 = v_65023 & v_65025;
assign v_65028 = v_65002 & v_65027;
assign v_65030 = v_62567;
assign v_65032 = v_65029 & v_65031;
assign v_65034 = v_64999 & v_65033;
assign v_65036 = v_62563;
assign v_65038 = v_65035 & v_65037;
assign v_65040 = v_64996 & v_65039;
assign v_65042 = v_62559;
assign v_65044 = v_65041 & v_65043;
assign v_65046 = v_64993 & v_65045;
assign v_65048 = v_62555;
assign v_65050 = v_65047 & v_65049;
assign v_65052 = v_64990 & v_65051;
assign v_65054 = v_62551;
assign v_65056 = v_65053 & v_65055;
assign v_65058 = v_64987 & v_65057;
assign v_65060 = v_62547;
assign v_65062 = v_65059 & v_65061;
assign v_65064 = v_64984 & v_65063;
assign v_65066 = v_62543;
assign v_65068 = v_65065 & v_65067;
assign v_65070 = v_64981 & v_65069;
assign v_65072 = v_62539;
assign v_65074 = v_65071 & v_65073;
assign v_65076 = v_64978 & v_65075;
assign v_65078 = v_62535;
assign v_65080 = v_65077 & v_65079;
assign v_65082 = v_64975 & v_65081;
assign v_65084 = v_62531;
assign v_65086 = v_65083 & v_65085;
assign v_65088 = v_64972 & v_65087;
assign v_65090 = v_2635;
assign v_65092 = v_65089 & v_65091;
assign v_65094 = v_64969 & v_65093;
assign v_65096 = v_2631;
assign v_65098 = v_65095 & v_65097;
assign v_65100 = v_64966 & v_65099;
assign v_65102 = v_2627;
assign v_65104 = v_65101 & v_65103;
assign v_65106 = v_64963 & v_65105;
assign v_65108 = v_2623;
assign v_65110 = v_65107 & v_65109;
assign v_65111 = v_65110;
assign v_65113 = v_62579;
assign v_65114 = v_2688;
assign v_65115 = v_65114;
assign v_65116 = v_65113 & v_65115;
assign v_65117 = v_65116;
assign v_65118 = v_65008 & v_65117;
assign v_65120 = v_65018 & v_65119;
assign v_65121 = v_65007 & v_65117;
assign v_65123 = v_65005 & v_65122;
assign v_65125 = v_65024 & v_65124;
assign v_65126 = v_65004 & v_65122;
assign v_65128 = v_65002 & v_65127;
assign v_65130 = v_65030 & v_65129;
assign v_65131 = v_65001 & v_65127;
assign v_65133 = v_64999 & v_65132;
assign v_65135 = v_65036 & v_65134;
assign v_65136 = v_64998 & v_65132;
assign v_65138 = v_64996 & v_65137;
assign v_65140 = v_65042 & v_65139;
assign v_65141 = v_64995 & v_65137;
assign v_65143 = v_64993 & v_65142;
assign v_65145 = v_65048 & v_65144;
assign v_65146 = v_64992 & v_65142;
assign v_65148 = v_64990 & v_65147;
assign v_65150 = v_65054 & v_65149;
assign v_65151 = v_64989 & v_65147;
assign v_65153 = v_64987 & v_65152;
assign v_65155 = v_65060 & v_65154;
assign v_65156 = v_64986 & v_65152;
assign v_65158 = v_64984 & v_65157;
assign v_65160 = v_65066 & v_65159;
assign v_65161 = v_64983 & v_65157;
assign v_65163 = v_64981 & v_65162;
assign v_65165 = v_65072 & v_65164;
assign v_65166 = v_64980 & v_65162;
assign v_65168 = v_64978 & v_65167;
assign v_65170 = v_65078 & v_65169;
assign v_65171 = v_64977 & v_65167;
assign v_65173 = v_64975 & v_65172;
assign v_65175 = v_65084 & v_65174;
assign v_65176 = v_64974 & v_65172;
assign v_65178 = v_64972 & v_65177;
assign v_65180 = v_65090 & v_65179;
assign v_65181 = v_64971 & v_65177;
assign v_65183 = v_64969 & v_65182;
assign v_65185 = v_65096 & v_65184;
assign v_65186 = v_64968 & v_65182;
assign v_65188 = v_64966 & v_65187;
assign v_65190 = v_65102 & v_65189;
assign v_65191 = v_64965 & v_65187;
assign v_65193 = v_64963 & v_65192;
assign v_65195 = v_65108 & v_65194;
assign v_65196 = v_64962 & v_65192;
assign v_65198 = v_65197;
assign v_65200 = v_65112 & v_65199;
assign v_65201 = v_65200;
assign v_65203 = v_65202;
assign v_65205 = ~v_2883;
assign v_65206 = ~v_62516;
assign v_65207 = v_62516;
assign v_65208 = ~v_2887;
assign v_65209 = ~v_62520;
assign v_65210 = v_62520;
assign v_65211 = ~v_2891;
assign v_65212 = ~v_62524;
assign v_65213 = v_62524;
assign v_65214 = ~v_2895;
assign v_65215 = ~v_62528;
assign v_65216 = v_62528;
assign v_65217 = ~v_62531;
assign v_65218 = ~v_2900;
assign v_65219 = v_2900;
assign v_65220 = ~v_62535;
assign v_65221 = ~v_2904;
assign v_65222 = v_2904;
assign v_65223 = ~v_62539;
assign v_65224 = ~v_2908;
assign v_65225 = v_2908;
assign v_65226 = ~v_62543;
assign v_65227 = ~v_2912;
assign v_65228 = v_2912;
assign v_65229 = ~v_62547;
assign v_65230 = ~v_2916;
assign v_65231 = v_2916;
assign v_65232 = ~v_62551;
assign v_65233 = ~v_2920;
assign v_65234 = v_2920;
assign v_65235 = ~v_62555;
assign v_65236 = ~v_2924;
assign v_65237 = v_2924;
assign v_65238 = ~v_62559;
assign v_65239 = ~v_2928;
assign v_65240 = v_2928;
assign v_65241 = ~v_62563;
assign v_65242 = ~v_2932;
assign v_65243 = v_2932;
assign v_65244 = ~v_62567;
assign v_65245 = ~v_2936;
assign v_65246 = v_2936;
assign v_65247 = ~v_62571;
assign v_65248 = ~v_2940;
assign v_65249 = v_2940;
assign v_65250 = ~v_62575;
assign v_65251 = ~v_2944;
assign v_65252 = v_2944;
assign v_65253 = ~v_62579;
assign v_65254 = ~v_2948;
assign v_65255 = v_65254;
assign v_65257 = v_65256;
assign v_65259 = v_65251 & v_65258;
assign v_65261 = v_62575;
assign v_65263 = v_65260 & v_65262;
assign v_65265 = v_65248 & v_65264;
assign v_65267 = v_62571;
assign v_65269 = v_65266 & v_65268;
assign v_65271 = v_65245 & v_65270;
assign v_65273 = v_62567;
assign v_65275 = v_65272 & v_65274;
assign v_65277 = v_65242 & v_65276;
assign v_65279 = v_62563;
assign v_65281 = v_65278 & v_65280;
assign v_65283 = v_65239 & v_65282;
assign v_65285 = v_62559;
assign v_65287 = v_65284 & v_65286;
assign v_65289 = v_65236 & v_65288;
assign v_65291 = v_62555;
assign v_65293 = v_65290 & v_65292;
assign v_65295 = v_65233 & v_65294;
assign v_65297 = v_62551;
assign v_65299 = v_65296 & v_65298;
assign v_65301 = v_65230 & v_65300;
assign v_65303 = v_62547;
assign v_65305 = v_65302 & v_65304;
assign v_65307 = v_65227 & v_65306;
assign v_65309 = v_62543;
assign v_65311 = v_65308 & v_65310;
assign v_65313 = v_65224 & v_65312;
assign v_65315 = v_62539;
assign v_65317 = v_65314 & v_65316;
assign v_65319 = v_65221 & v_65318;
assign v_65321 = v_62535;
assign v_65323 = v_65320 & v_65322;
assign v_65325 = v_65218 & v_65324;
assign v_65327 = v_62531;
assign v_65329 = v_65326 & v_65328;
assign v_65331 = v_65215 & v_65330;
assign v_65333 = v_2895;
assign v_65335 = v_65332 & v_65334;
assign v_65337 = v_65212 & v_65336;
assign v_65339 = v_2891;
assign v_65341 = v_65338 & v_65340;
assign v_65343 = v_65209 & v_65342;
assign v_65345 = v_2887;
assign v_65347 = v_65344 & v_65346;
assign v_65349 = v_65206 & v_65348;
assign v_65351 = v_2883;
assign v_65353 = v_65350 & v_65352;
assign v_65354 = v_65353;
assign v_65356 = v_62579;
assign v_65357 = v_2948;
assign v_65358 = v_65357;
assign v_65359 = v_65356 & v_65358;
assign v_65360 = v_65359;
assign v_65361 = v_65251 & v_65360;
assign v_65363 = v_65261 & v_65362;
assign v_65364 = v_65250 & v_65360;
assign v_65366 = v_65248 & v_65365;
assign v_65368 = v_65267 & v_65367;
assign v_65369 = v_65247 & v_65365;
assign v_65371 = v_65245 & v_65370;
assign v_65373 = v_65273 & v_65372;
assign v_65374 = v_65244 & v_65370;
assign v_65376 = v_65242 & v_65375;
assign v_65378 = v_65279 & v_65377;
assign v_65379 = v_65241 & v_65375;
assign v_65381 = v_65239 & v_65380;
assign v_65383 = v_65285 & v_65382;
assign v_65384 = v_65238 & v_65380;
assign v_65386 = v_65236 & v_65385;
assign v_65388 = v_65291 & v_65387;
assign v_65389 = v_65235 & v_65385;
assign v_65391 = v_65233 & v_65390;
assign v_65393 = v_65297 & v_65392;
assign v_65394 = v_65232 & v_65390;
assign v_65396 = v_65230 & v_65395;
assign v_65398 = v_65303 & v_65397;
assign v_65399 = v_65229 & v_65395;
assign v_65401 = v_65227 & v_65400;
assign v_65403 = v_65309 & v_65402;
assign v_65404 = v_65226 & v_65400;
assign v_65406 = v_65224 & v_65405;
assign v_65408 = v_65315 & v_65407;
assign v_65409 = v_65223 & v_65405;
assign v_65411 = v_65221 & v_65410;
assign v_65413 = v_65321 & v_65412;
assign v_65414 = v_65220 & v_65410;
assign v_65416 = v_65218 & v_65415;
assign v_65418 = v_65327 & v_65417;
assign v_65419 = v_65217 & v_65415;
assign v_65421 = v_65215 & v_65420;
assign v_65423 = v_65333 & v_65422;
assign v_65424 = v_65214 & v_65420;
assign v_65426 = v_65212 & v_65425;
assign v_65428 = v_65339 & v_65427;
assign v_65429 = v_65211 & v_65425;
assign v_65431 = v_65209 & v_65430;
assign v_65433 = v_65345 & v_65432;
assign v_65434 = v_65208 & v_65430;
assign v_65436 = v_65206 & v_65435;
assign v_65438 = v_65351 & v_65437;
assign v_65439 = v_65205 & v_65435;
assign v_65441 = v_65440;
assign v_65443 = v_65355 & v_65442;
assign v_65444 = v_65443;
assign v_65446 = v_65445;
assign v_65448 = ~v_3143;
assign v_65449 = ~v_62516;
assign v_65450 = v_62516;
assign v_65451 = ~v_3147;
assign v_65452 = ~v_62520;
assign v_65453 = v_62520;
assign v_65454 = ~v_3151;
assign v_65455 = ~v_62524;
assign v_65456 = v_62524;
assign v_65457 = ~v_3155;
assign v_65458 = ~v_62528;
assign v_65459 = v_62528;
assign v_65460 = ~v_62531;
assign v_65461 = ~v_3160;
assign v_65462 = v_3160;
assign v_65463 = ~v_62535;
assign v_65464 = ~v_3164;
assign v_65465 = v_3164;
assign v_65466 = ~v_62539;
assign v_65467 = ~v_3168;
assign v_65468 = v_3168;
assign v_65469 = ~v_62543;
assign v_65470 = ~v_3172;
assign v_65471 = v_3172;
assign v_65472 = ~v_62547;
assign v_65473 = ~v_3176;
assign v_65474 = v_3176;
assign v_65475 = ~v_62551;
assign v_65476 = ~v_3180;
assign v_65477 = v_3180;
assign v_65478 = ~v_62555;
assign v_65479 = ~v_3184;
assign v_65480 = v_3184;
assign v_65481 = ~v_62559;
assign v_65482 = ~v_3188;
assign v_65483 = v_3188;
assign v_65484 = ~v_62563;
assign v_65485 = ~v_3192;
assign v_65486 = v_3192;
assign v_65487 = ~v_62567;
assign v_65488 = ~v_3196;
assign v_65489 = v_3196;
assign v_65490 = ~v_62571;
assign v_65491 = ~v_3200;
assign v_65492 = v_3200;
assign v_65493 = ~v_62575;
assign v_65494 = ~v_3204;
assign v_65495 = v_3204;
assign v_65496 = ~v_62579;
assign v_65497 = ~v_3208;
assign v_65498 = v_65497;
assign v_65500 = v_65499;
assign v_65502 = v_65494 & v_65501;
assign v_65504 = v_62575;
assign v_65506 = v_65503 & v_65505;
assign v_65508 = v_65491 & v_65507;
assign v_65510 = v_62571;
assign v_65512 = v_65509 & v_65511;
assign v_65514 = v_65488 & v_65513;
assign v_65516 = v_62567;
assign v_65518 = v_65515 & v_65517;
assign v_65520 = v_65485 & v_65519;
assign v_65522 = v_62563;
assign v_65524 = v_65521 & v_65523;
assign v_65526 = v_65482 & v_65525;
assign v_65528 = v_62559;
assign v_65530 = v_65527 & v_65529;
assign v_65532 = v_65479 & v_65531;
assign v_65534 = v_62555;
assign v_65536 = v_65533 & v_65535;
assign v_65538 = v_65476 & v_65537;
assign v_65540 = v_62551;
assign v_65542 = v_65539 & v_65541;
assign v_65544 = v_65473 & v_65543;
assign v_65546 = v_62547;
assign v_65548 = v_65545 & v_65547;
assign v_65550 = v_65470 & v_65549;
assign v_65552 = v_62543;
assign v_65554 = v_65551 & v_65553;
assign v_65556 = v_65467 & v_65555;
assign v_65558 = v_62539;
assign v_65560 = v_65557 & v_65559;
assign v_65562 = v_65464 & v_65561;
assign v_65564 = v_62535;
assign v_65566 = v_65563 & v_65565;
assign v_65568 = v_65461 & v_65567;
assign v_65570 = v_62531;
assign v_65572 = v_65569 & v_65571;
assign v_65574 = v_65458 & v_65573;
assign v_65576 = v_3155;
assign v_65578 = v_65575 & v_65577;
assign v_65580 = v_65455 & v_65579;
assign v_65582 = v_3151;
assign v_65584 = v_65581 & v_65583;
assign v_65586 = v_65452 & v_65585;
assign v_65588 = v_3147;
assign v_65590 = v_65587 & v_65589;
assign v_65592 = v_65449 & v_65591;
assign v_65594 = v_3143;
assign v_65596 = v_65593 & v_65595;
assign v_65597 = v_65596;
assign v_65599 = v_62579;
assign v_65600 = v_3208;
assign v_65601 = v_65600;
assign v_65602 = v_65599 & v_65601;
assign v_65603 = v_65602;
assign v_65604 = v_65494 & v_65603;
assign v_65606 = v_65504 & v_65605;
assign v_65607 = v_65493 & v_65603;
assign v_65609 = v_65491 & v_65608;
assign v_65611 = v_65510 & v_65610;
assign v_65612 = v_65490 & v_65608;
assign v_65614 = v_65488 & v_65613;
assign v_65616 = v_65516 & v_65615;
assign v_65617 = v_65487 & v_65613;
assign v_65619 = v_65485 & v_65618;
assign v_65621 = v_65522 & v_65620;
assign v_65622 = v_65484 & v_65618;
assign v_65624 = v_65482 & v_65623;
assign v_65626 = v_65528 & v_65625;
assign v_65627 = v_65481 & v_65623;
assign v_65629 = v_65479 & v_65628;
assign v_65631 = v_65534 & v_65630;
assign v_65632 = v_65478 & v_65628;
assign v_65634 = v_65476 & v_65633;
assign v_65636 = v_65540 & v_65635;
assign v_65637 = v_65475 & v_65633;
assign v_65639 = v_65473 & v_65638;
assign v_65641 = v_65546 & v_65640;
assign v_65642 = v_65472 & v_65638;
assign v_65644 = v_65470 & v_65643;
assign v_65646 = v_65552 & v_65645;
assign v_65647 = v_65469 & v_65643;
assign v_65649 = v_65467 & v_65648;
assign v_65651 = v_65558 & v_65650;
assign v_65652 = v_65466 & v_65648;
assign v_65654 = v_65464 & v_65653;
assign v_65656 = v_65564 & v_65655;
assign v_65657 = v_65463 & v_65653;
assign v_65659 = v_65461 & v_65658;
assign v_65661 = v_65570 & v_65660;
assign v_65662 = v_65460 & v_65658;
assign v_65664 = v_65458 & v_65663;
assign v_65666 = v_65576 & v_65665;
assign v_65667 = v_65457 & v_65663;
assign v_65669 = v_65455 & v_65668;
assign v_65671 = v_65582 & v_65670;
assign v_65672 = v_65454 & v_65668;
assign v_65674 = v_65452 & v_65673;
assign v_65676 = v_65588 & v_65675;
assign v_65677 = v_65451 & v_65673;
assign v_65679 = v_65449 & v_65678;
assign v_65681 = v_65594 & v_65680;
assign v_65682 = v_65448 & v_65678;
assign v_65684 = v_65683;
assign v_65686 = v_65598 & v_65685;
assign v_65687 = v_65686;
assign v_65689 = v_65688;
assign v_65691 = ~v_3403;
assign v_65692 = ~v_62516;
assign v_65693 = v_62516;
assign v_65694 = ~v_3407;
assign v_65695 = ~v_62520;
assign v_65696 = v_62520;
assign v_65697 = ~v_3411;
assign v_65698 = ~v_62524;
assign v_65699 = v_62524;
assign v_65700 = ~v_3415;
assign v_65701 = ~v_62528;
assign v_65702 = v_62528;
assign v_65703 = ~v_62531;
assign v_65704 = ~v_3420;
assign v_65705 = v_3420;
assign v_65706 = ~v_62535;
assign v_65707 = ~v_3424;
assign v_65708 = v_3424;
assign v_65709 = ~v_62539;
assign v_65710 = ~v_3428;
assign v_65711 = v_3428;
assign v_65712 = ~v_62543;
assign v_65713 = ~v_3432;
assign v_65714 = v_3432;
assign v_65715 = ~v_62547;
assign v_65716 = ~v_3436;
assign v_65717 = v_3436;
assign v_65718 = ~v_62551;
assign v_65719 = ~v_3440;
assign v_65720 = v_3440;
assign v_65721 = ~v_62555;
assign v_65722 = ~v_3444;
assign v_65723 = v_3444;
assign v_65724 = ~v_62559;
assign v_65725 = ~v_3448;
assign v_65726 = v_3448;
assign v_65727 = ~v_62563;
assign v_65728 = ~v_3452;
assign v_65729 = v_3452;
assign v_65730 = ~v_62567;
assign v_65731 = ~v_3456;
assign v_65732 = v_3456;
assign v_65733 = ~v_62571;
assign v_65734 = ~v_3460;
assign v_65735 = v_3460;
assign v_65736 = ~v_62575;
assign v_65737 = ~v_3464;
assign v_65738 = v_3464;
assign v_65739 = ~v_62579;
assign v_65740 = ~v_3468;
assign v_65741 = v_65740;
assign v_65743 = v_65742;
assign v_65745 = v_65737 & v_65744;
assign v_65747 = v_62575;
assign v_65749 = v_65746 & v_65748;
assign v_65751 = v_65734 & v_65750;
assign v_65753 = v_62571;
assign v_65755 = v_65752 & v_65754;
assign v_65757 = v_65731 & v_65756;
assign v_65759 = v_62567;
assign v_65761 = v_65758 & v_65760;
assign v_65763 = v_65728 & v_65762;
assign v_65765 = v_62563;
assign v_65767 = v_65764 & v_65766;
assign v_65769 = v_65725 & v_65768;
assign v_65771 = v_62559;
assign v_65773 = v_65770 & v_65772;
assign v_65775 = v_65722 & v_65774;
assign v_65777 = v_62555;
assign v_65779 = v_65776 & v_65778;
assign v_65781 = v_65719 & v_65780;
assign v_65783 = v_62551;
assign v_65785 = v_65782 & v_65784;
assign v_65787 = v_65716 & v_65786;
assign v_65789 = v_62547;
assign v_65791 = v_65788 & v_65790;
assign v_65793 = v_65713 & v_65792;
assign v_65795 = v_62543;
assign v_65797 = v_65794 & v_65796;
assign v_65799 = v_65710 & v_65798;
assign v_65801 = v_62539;
assign v_65803 = v_65800 & v_65802;
assign v_65805 = v_65707 & v_65804;
assign v_65807 = v_62535;
assign v_65809 = v_65806 & v_65808;
assign v_65811 = v_65704 & v_65810;
assign v_65813 = v_62531;
assign v_65815 = v_65812 & v_65814;
assign v_65817 = v_65701 & v_65816;
assign v_65819 = v_3415;
assign v_65821 = v_65818 & v_65820;
assign v_65823 = v_65698 & v_65822;
assign v_65825 = v_3411;
assign v_65827 = v_65824 & v_65826;
assign v_65829 = v_65695 & v_65828;
assign v_65831 = v_3407;
assign v_65833 = v_65830 & v_65832;
assign v_65835 = v_65692 & v_65834;
assign v_65837 = v_3403;
assign v_65839 = v_65836 & v_65838;
assign v_65840 = v_65839;
assign v_65842 = v_62579;
assign v_65843 = v_3468;
assign v_65844 = v_65843;
assign v_65845 = v_65842 & v_65844;
assign v_65846 = v_65845;
assign v_65847 = v_65737 & v_65846;
assign v_65849 = v_65747 & v_65848;
assign v_65850 = v_65736 & v_65846;
assign v_65852 = v_65734 & v_65851;
assign v_65854 = v_65753 & v_65853;
assign v_65855 = v_65733 & v_65851;
assign v_65857 = v_65731 & v_65856;
assign v_65859 = v_65759 & v_65858;
assign v_65860 = v_65730 & v_65856;
assign v_65862 = v_65728 & v_65861;
assign v_65864 = v_65765 & v_65863;
assign v_65865 = v_65727 & v_65861;
assign v_65867 = v_65725 & v_65866;
assign v_65869 = v_65771 & v_65868;
assign v_65870 = v_65724 & v_65866;
assign v_65872 = v_65722 & v_65871;
assign v_65874 = v_65777 & v_65873;
assign v_65875 = v_65721 & v_65871;
assign v_65877 = v_65719 & v_65876;
assign v_65879 = v_65783 & v_65878;
assign v_65880 = v_65718 & v_65876;
assign v_65882 = v_65716 & v_65881;
assign v_65884 = v_65789 & v_65883;
assign v_65885 = v_65715 & v_65881;
assign v_65887 = v_65713 & v_65886;
assign v_65889 = v_65795 & v_65888;
assign v_65890 = v_65712 & v_65886;
assign v_65892 = v_65710 & v_65891;
assign v_65894 = v_65801 & v_65893;
assign v_65895 = v_65709 & v_65891;
assign v_65897 = v_65707 & v_65896;
assign v_65899 = v_65807 & v_65898;
assign v_65900 = v_65706 & v_65896;
assign v_65902 = v_65704 & v_65901;
assign v_65904 = v_65813 & v_65903;
assign v_65905 = v_65703 & v_65901;
assign v_65907 = v_65701 & v_65906;
assign v_65909 = v_65819 & v_65908;
assign v_65910 = v_65700 & v_65906;
assign v_65912 = v_65698 & v_65911;
assign v_65914 = v_65825 & v_65913;
assign v_65915 = v_65697 & v_65911;
assign v_65917 = v_65695 & v_65916;
assign v_65919 = v_65831 & v_65918;
assign v_65920 = v_65694 & v_65916;
assign v_65922 = v_65692 & v_65921;
assign v_65924 = v_65837 & v_65923;
assign v_65925 = v_65691 & v_65921;
assign v_65927 = v_65926;
assign v_65929 = v_65841 & v_65928;
assign v_65930 = v_65929;
assign v_65932 = v_65931;
assign v_65934 = ~v_3663;
assign v_65935 = ~v_62516;
assign v_65936 = v_62516;
assign v_65937 = ~v_3667;
assign v_65938 = ~v_62520;
assign v_65939 = v_62520;
assign v_65940 = ~v_3671;
assign v_65941 = ~v_62524;
assign v_65942 = v_62524;
assign v_65943 = ~v_3675;
assign v_65944 = ~v_62528;
assign v_65945 = v_62528;
assign v_65946 = ~v_62531;
assign v_65947 = ~v_3680;
assign v_65948 = v_3680;
assign v_65949 = ~v_62535;
assign v_65950 = ~v_3684;
assign v_65951 = v_3684;
assign v_65952 = ~v_62539;
assign v_65953 = ~v_3688;
assign v_65954 = v_3688;
assign v_65955 = ~v_62543;
assign v_65956 = ~v_3692;
assign v_65957 = v_3692;
assign v_65958 = ~v_62547;
assign v_65959 = ~v_3696;
assign v_65960 = v_3696;
assign v_65961 = ~v_62551;
assign v_65962 = ~v_3700;
assign v_65963 = v_3700;
assign v_65964 = ~v_62555;
assign v_65965 = ~v_3704;
assign v_65966 = v_3704;
assign v_65967 = ~v_62559;
assign v_65968 = ~v_3708;
assign v_65969 = v_3708;
assign v_65970 = ~v_62563;
assign v_65971 = ~v_3712;
assign v_65972 = v_3712;
assign v_65973 = ~v_62567;
assign v_65974 = ~v_3716;
assign v_65975 = v_3716;
assign v_65976 = ~v_62571;
assign v_65977 = ~v_3720;
assign v_65978 = v_3720;
assign v_65979 = ~v_62575;
assign v_65980 = ~v_3724;
assign v_65981 = v_3724;
assign v_65982 = ~v_62579;
assign v_65983 = ~v_3728;
assign v_65984 = v_65983;
assign v_65986 = v_65985;
assign v_65988 = v_65980 & v_65987;
assign v_65990 = v_62575;
assign v_65992 = v_65989 & v_65991;
assign v_65994 = v_65977 & v_65993;
assign v_65996 = v_62571;
assign v_65998 = v_65995 & v_65997;
assign v_66000 = v_65974 & v_65999;
assign v_66002 = v_62567;
assign v_66004 = v_66001 & v_66003;
assign v_66006 = v_65971 & v_66005;
assign v_66008 = v_62563;
assign v_66010 = v_66007 & v_66009;
assign v_66012 = v_65968 & v_66011;
assign v_66014 = v_62559;
assign v_66016 = v_66013 & v_66015;
assign v_66018 = v_65965 & v_66017;
assign v_66020 = v_62555;
assign v_66022 = v_66019 & v_66021;
assign v_66024 = v_65962 & v_66023;
assign v_66026 = v_62551;
assign v_66028 = v_66025 & v_66027;
assign v_66030 = v_65959 & v_66029;
assign v_66032 = v_62547;
assign v_66034 = v_66031 & v_66033;
assign v_66036 = v_65956 & v_66035;
assign v_66038 = v_62543;
assign v_66040 = v_66037 & v_66039;
assign v_66042 = v_65953 & v_66041;
assign v_66044 = v_62539;
assign v_66046 = v_66043 & v_66045;
assign v_66048 = v_65950 & v_66047;
assign v_66050 = v_62535;
assign v_66052 = v_66049 & v_66051;
assign v_66054 = v_65947 & v_66053;
assign v_66056 = v_62531;
assign v_66058 = v_66055 & v_66057;
assign v_66060 = v_65944 & v_66059;
assign v_66062 = v_3675;
assign v_66064 = v_66061 & v_66063;
assign v_66066 = v_65941 & v_66065;
assign v_66068 = v_3671;
assign v_66070 = v_66067 & v_66069;
assign v_66072 = v_65938 & v_66071;
assign v_66074 = v_3667;
assign v_66076 = v_66073 & v_66075;
assign v_66078 = v_65935 & v_66077;
assign v_66080 = v_3663;
assign v_66082 = v_66079 & v_66081;
assign v_66083 = v_66082;
assign v_66085 = v_62579;
assign v_66086 = v_3728;
assign v_66087 = v_66086;
assign v_66088 = v_66085 & v_66087;
assign v_66089 = v_66088;
assign v_66090 = v_65980 & v_66089;
assign v_66092 = v_65990 & v_66091;
assign v_66093 = v_65979 & v_66089;
assign v_66095 = v_65977 & v_66094;
assign v_66097 = v_65996 & v_66096;
assign v_66098 = v_65976 & v_66094;
assign v_66100 = v_65974 & v_66099;
assign v_66102 = v_66002 & v_66101;
assign v_66103 = v_65973 & v_66099;
assign v_66105 = v_65971 & v_66104;
assign v_66107 = v_66008 & v_66106;
assign v_66108 = v_65970 & v_66104;
assign v_66110 = v_65968 & v_66109;
assign v_66112 = v_66014 & v_66111;
assign v_66113 = v_65967 & v_66109;
assign v_66115 = v_65965 & v_66114;
assign v_66117 = v_66020 & v_66116;
assign v_66118 = v_65964 & v_66114;
assign v_66120 = v_65962 & v_66119;
assign v_66122 = v_66026 & v_66121;
assign v_66123 = v_65961 & v_66119;
assign v_66125 = v_65959 & v_66124;
assign v_66127 = v_66032 & v_66126;
assign v_66128 = v_65958 & v_66124;
assign v_66130 = v_65956 & v_66129;
assign v_66132 = v_66038 & v_66131;
assign v_66133 = v_65955 & v_66129;
assign v_66135 = v_65953 & v_66134;
assign v_66137 = v_66044 & v_66136;
assign v_66138 = v_65952 & v_66134;
assign v_66140 = v_65950 & v_66139;
assign v_66142 = v_66050 & v_66141;
assign v_66143 = v_65949 & v_66139;
assign v_66145 = v_65947 & v_66144;
assign v_66147 = v_66056 & v_66146;
assign v_66148 = v_65946 & v_66144;
assign v_66150 = v_65944 & v_66149;
assign v_66152 = v_66062 & v_66151;
assign v_66153 = v_65943 & v_66149;
assign v_66155 = v_65941 & v_66154;
assign v_66157 = v_66068 & v_66156;
assign v_66158 = v_65940 & v_66154;
assign v_66160 = v_65938 & v_66159;
assign v_66162 = v_66074 & v_66161;
assign v_66163 = v_65937 & v_66159;
assign v_66165 = v_65935 & v_66164;
assign v_66167 = v_66080 & v_66166;
assign v_66168 = v_65934 & v_66164;
assign v_66170 = v_66169;
assign v_66172 = v_66084 & v_66171;
assign v_66173 = v_66172;
assign v_66175 = v_66174;
assign v_66177 = ~v_3923;
assign v_66178 = ~v_62516;
assign v_66179 = v_62516;
assign v_66180 = ~v_3927;
assign v_66181 = ~v_62520;
assign v_66182 = v_62520;
assign v_66183 = ~v_3931;
assign v_66184 = ~v_62524;
assign v_66185 = v_62524;
assign v_66186 = ~v_3935;
assign v_66187 = ~v_62528;
assign v_66188 = v_62528;
assign v_66189 = ~v_62531;
assign v_66190 = ~v_3940;
assign v_66191 = v_3940;
assign v_66192 = ~v_62535;
assign v_66193 = ~v_3944;
assign v_66194 = v_3944;
assign v_66195 = ~v_62539;
assign v_66196 = ~v_3948;
assign v_66197 = v_3948;
assign v_66198 = ~v_62543;
assign v_66199 = ~v_3952;
assign v_66200 = v_3952;
assign v_66201 = ~v_62547;
assign v_66202 = ~v_3956;
assign v_66203 = v_3956;
assign v_66204 = ~v_62551;
assign v_66205 = ~v_3960;
assign v_66206 = v_3960;
assign v_66207 = ~v_62555;
assign v_66208 = ~v_3964;
assign v_66209 = v_3964;
assign v_66210 = ~v_62559;
assign v_66211 = ~v_3968;
assign v_66212 = v_3968;
assign v_66213 = ~v_62563;
assign v_66214 = ~v_3972;
assign v_66215 = v_3972;
assign v_66216 = ~v_62567;
assign v_66217 = ~v_3976;
assign v_66218 = v_3976;
assign v_66219 = ~v_62571;
assign v_66220 = ~v_3980;
assign v_66221 = v_3980;
assign v_66222 = ~v_62575;
assign v_66223 = ~v_3984;
assign v_66224 = v_3984;
assign v_66225 = ~v_62579;
assign v_66226 = ~v_3988;
assign v_66227 = v_66226;
assign v_66229 = v_66228;
assign v_66231 = v_66223 & v_66230;
assign v_66233 = v_62575;
assign v_66235 = v_66232 & v_66234;
assign v_66237 = v_66220 & v_66236;
assign v_66239 = v_62571;
assign v_66241 = v_66238 & v_66240;
assign v_66243 = v_66217 & v_66242;
assign v_66245 = v_62567;
assign v_66247 = v_66244 & v_66246;
assign v_66249 = v_66214 & v_66248;
assign v_66251 = v_62563;
assign v_66253 = v_66250 & v_66252;
assign v_66255 = v_66211 & v_66254;
assign v_66257 = v_62559;
assign v_66259 = v_66256 & v_66258;
assign v_66261 = v_66208 & v_66260;
assign v_66263 = v_62555;
assign v_66265 = v_66262 & v_66264;
assign v_66267 = v_66205 & v_66266;
assign v_66269 = v_62551;
assign v_66271 = v_66268 & v_66270;
assign v_66273 = v_66202 & v_66272;
assign v_66275 = v_62547;
assign v_66277 = v_66274 & v_66276;
assign v_66279 = v_66199 & v_66278;
assign v_66281 = v_62543;
assign v_66283 = v_66280 & v_66282;
assign v_66285 = v_66196 & v_66284;
assign v_66287 = v_62539;
assign v_66289 = v_66286 & v_66288;
assign v_66291 = v_66193 & v_66290;
assign v_66293 = v_62535;
assign v_66295 = v_66292 & v_66294;
assign v_66297 = v_66190 & v_66296;
assign v_66299 = v_62531;
assign v_66301 = v_66298 & v_66300;
assign v_66303 = v_66187 & v_66302;
assign v_66305 = v_3935;
assign v_66307 = v_66304 & v_66306;
assign v_66309 = v_66184 & v_66308;
assign v_66311 = v_3931;
assign v_66313 = v_66310 & v_66312;
assign v_66315 = v_66181 & v_66314;
assign v_66317 = v_3927;
assign v_66319 = v_66316 & v_66318;
assign v_66321 = v_66178 & v_66320;
assign v_66323 = v_3923;
assign v_66325 = v_66322 & v_66324;
assign v_66326 = v_66325;
assign v_66328 = v_62579;
assign v_66329 = v_3988;
assign v_66330 = v_66329;
assign v_66331 = v_66328 & v_66330;
assign v_66332 = v_66331;
assign v_66333 = v_66223 & v_66332;
assign v_66335 = v_66233 & v_66334;
assign v_66336 = v_66222 & v_66332;
assign v_66338 = v_66220 & v_66337;
assign v_66340 = v_66239 & v_66339;
assign v_66341 = v_66219 & v_66337;
assign v_66343 = v_66217 & v_66342;
assign v_66345 = v_66245 & v_66344;
assign v_66346 = v_66216 & v_66342;
assign v_66348 = v_66214 & v_66347;
assign v_66350 = v_66251 & v_66349;
assign v_66351 = v_66213 & v_66347;
assign v_66353 = v_66211 & v_66352;
assign v_66355 = v_66257 & v_66354;
assign v_66356 = v_66210 & v_66352;
assign v_66358 = v_66208 & v_66357;
assign v_66360 = v_66263 & v_66359;
assign v_66361 = v_66207 & v_66357;
assign v_66363 = v_66205 & v_66362;
assign v_66365 = v_66269 & v_66364;
assign v_66366 = v_66204 & v_66362;
assign v_66368 = v_66202 & v_66367;
assign v_66370 = v_66275 & v_66369;
assign v_66371 = v_66201 & v_66367;
assign v_66373 = v_66199 & v_66372;
assign v_66375 = v_66281 & v_66374;
assign v_66376 = v_66198 & v_66372;
assign v_66378 = v_66196 & v_66377;
assign v_66380 = v_66287 & v_66379;
assign v_66381 = v_66195 & v_66377;
assign v_66383 = v_66193 & v_66382;
assign v_66385 = v_66293 & v_66384;
assign v_66386 = v_66192 & v_66382;
assign v_66388 = v_66190 & v_66387;
assign v_66390 = v_66299 & v_66389;
assign v_66391 = v_66189 & v_66387;
assign v_66393 = v_66187 & v_66392;
assign v_66395 = v_66305 & v_66394;
assign v_66396 = v_66186 & v_66392;
assign v_66398 = v_66184 & v_66397;
assign v_66400 = v_66311 & v_66399;
assign v_66401 = v_66183 & v_66397;
assign v_66403 = v_66181 & v_66402;
assign v_66405 = v_66317 & v_66404;
assign v_66406 = v_66180 & v_66402;
assign v_66408 = v_66178 & v_66407;
assign v_66410 = v_66323 & v_66409;
assign v_66411 = v_66177 & v_66407;
assign v_66413 = v_66412;
assign v_66415 = v_66327 & v_66414;
assign v_66416 = v_66415;
assign v_66418 = v_66417;
assign v_66419 = ~v_4182;
assign v_66420 = ~v_62516;
assign v_66421 = v_62516;
assign v_66422 = ~v_4186;
assign v_66423 = ~v_62520;
assign v_66424 = v_62520;
assign v_66425 = ~v_4190;
assign v_66426 = ~v_62524;
assign v_66427 = v_62524;
assign v_66428 = ~v_4194;
assign v_66429 = ~v_62528;
assign v_66430 = v_62528;
assign v_66431 = ~v_62531;
assign v_66432 = ~v_4199;
assign v_66433 = v_4199;
assign v_66434 = ~v_62535;
assign v_66435 = ~v_4203;
assign v_66436 = v_4203;
assign v_66437 = ~v_62539;
assign v_66438 = ~v_4207;
assign v_66439 = v_4207;
assign v_66440 = ~v_62543;
assign v_66441 = ~v_4211;
assign v_66442 = v_4211;
assign v_66443 = ~v_62547;
assign v_66444 = ~v_4215;
assign v_66445 = v_4215;
assign v_66446 = ~v_62551;
assign v_66447 = ~v_4219;
assign v_66448 = v_4219;
assign v_66449 = ~v_62555;
assign v_66450 = ~v_4223;
assign v_66451 = v_4223;
assign v_66452 = ~v_62559;
assign v_66453 = ~v_4227;
assign v_66454 = v_4227;
assign v_66455 = ~v_62563;
assign v_66456 = ~v_4231;
assign v_66457 = v_4231;
assign v_66458 = ~v_62567;
assign v_66459 = ~v_4235;
assign v_66460 = v_4235;
assign v_66461 = ~v_62571;
assign v_66462 = ~v_4239;
assign v_66463 = v_4239;
assign v_66464 = ~v_62575;
assign v_66465 = ~v_4243;
assign v_66466 = v_4243;
assign v_66467 = ~v_62579;
assign v_66468 = ~v_4247;
assign v_66469 = v_66468;
assign v_66471 = v_66470;
assign v_66473 = v_66465 & v_66472;
assign v_66475 = v_62575;
assign v_66477 = v_66474 & v_66476;
assign v_66479 = v_66462 & v_66478;
assign v_66481 = v_62571;
assign v_66483 = v_66480 & v_66482;
assign v_66485 = v_66459 & v_66484;
assign v_66487 = v_62567;
assign v_66489 = v_66486 & v_66488;
assign v_66491 = v_66456 & v_66490;
assign v_66493 = v_62563;
assign v_66495 = v_66492 & v_66494;
assign v_66497 = v_66453 & v_66496;
assign v_66499 = v_62559;
assign v_66501 = v_66498 & v_66500;
assign v_66503 = v_66450 & v_66502;
assign v_66505 = v_62555;
assign v_66507 = v_66504 & v_66506;
assign v_66509 = v_66447 & v_66508;
assign v_66511 = v_62551;
assign v_66513 = v_66510 & v_66512;
assign v_66515 = v_66444 & v_66514;
assign v_66517 = v_62547;
assign v_66519 = v_66516 & v_66518;
assign v_66521 = v_66441 & v_66520;
assign v_66523 = v_62543;
assign v_66525 = v_66522 & v_66524;
assign v_66527 = v_66438 & v_66526;
assign v_66529 = v_62539;
assign v_66531 = v_66528 & v_66530;
assign v_66533 = v_66435 & v_66532;
assign v_66535 = v_62535;
assign v_66537 = v_66534 & v_66536;
assign v_66539 = v_66432 & v_66538;
assign v_66541 = v_62531;
assign v_66543 = v_66540 & v_66542;
assign v_66545 = v_66429 & v_66544;
assign v_66547 = v_4194;
assign v_66549 = v_66546 & v_66548;
assign v_66551 = v_66426 & v_66550;
assign v_66553 = v_4190;
assign v_66555 = v_66552 & v_66554;
assign v_66557 = v_66423 & v_66556;
assign v_66559 = v_4186;
assign v_66561 = v_66558 & v_66560;
assign v_66563 = v_66420 & v_66562;
assign v_66565 = v_4182;
assign v_66567 = v_66564 & v_66566;
assign v_66569 = ~v_66568;
assign v_66571 = v_62579;
assign v_66572 = v_4247;
assign v_66573 = v_66572;
assign v_66574 = v_66571 & v_66573;
assign v_66575 = v_66574;
assign v_66576 = v_66465 & v_66575;
assign v_66578 = v_66475 & v_66577;
assign v_66579 = v_66464 & v_66575;
assign v_66581 = v_66462 & v_66580;
assign v_66583 = v_66481 & v_66582;
assign v_66584 = v_66461 & v_66580;
assign v_66586 = v_66459 & v_66585;
assign v_66588 = v_66487 & v_66587;
assign v_66589 = v_66458 & v_66585;
assign v_66591 = v_66456 & v_66590;
assign v_66593 = v_66493 & v_66592;
assign v_66594 = v_66455 & v_66590;
assign v_66596 = v_66453 & v_66595;
assign v_66598 = v_66499 & v_66597;
assign v_66599 = v_66452 & v_66595;
assign v_66601 = v_66450 & v_66600;
assign v_66603 = v_66505 & v_66602;
assign v_66604 = v_66449 & v_66600;
assign v_66606 = v_66447 & v_66605;
assign v_66608 = v_66511 & v_66607;
assign v_66609 = v_66446 & v_66605;
assign v_66611 = v_66444 & v_66610;
assign v_66613 = v_66517 & v_66612;
assign v_66614 = v_66443 & v_66610;
assign v_66616 = v_66441 & v_66615;
assign v_66618 = v_66523 & v_66617;
assign v_66619 = v_66440 & v_66615;
assign v_66621 = v_66438 & v_66620;
assign v_66623 = v_66529 & v_66622;
assign v_66624 = v_66437 & v_66620;
assign v_66626 = v_66435 & v_66625;
assign v_66628 = v_66535 & v_66627;
assign v_66629 = v_66434 & v_66625;
assign v_66631 = v_66432 & v_66630;
assign v_66633 = v_66541 & v_66632;
assign v_66634 = v_66431 & v_66630;
assign v_66636 = v_66429 & v_66635;
assign v_66638 = v_66547 & v_66637;
assign v_66639 = v_66428 & v_66635;
assign v_66641 = v_66426 & v_66640;
assign v_66643 = v_66553 & v_66642;
assign v_66644 = v_66425 & v_66640;
assign v_66646 = v_66423 & v_66645;
assign v_66648 = v_66559 & v_66647;
assign v_66649 = v_66422 & v_66645;
assign v_66651 = v_66420 & v_66650;
assign v_66653 = v_66565 & v_66652;
assign v_66654 = v_66419 & v_66650;
assign v_66656 = v_66568;
assign v_66658 = v_66570 & v_66657;
assign v_66659 = v_66658;
assign v_66661 = v_66660;
assign v_66662 = ~v_6;
assign v_66664 = ~v_66663;
assign v_66665 = v_66663;
assign v_66666 = ~v_13;
assign v_66668 = ~v_66667;
assign v_66669 = v_66667;
assign v_66670 = ~v_18;
assign v_66672 = ~v_66671;
assign v_66673 = v_66671;
assign v_66674 = ~v_23;
assign v_66676 = ~v_66675;
assign v_66677 = v_66675;
assign v_66679 = ~v_66678;
assign v_66680 = ~v_30;
assign v_66681 = v_30;
assign v_66683 = ~v_66682;
assign v_66684 = ~v_35;
assign v_66685 = v_35;
assign v_66687 = ~v_66686;
assign v_66688 = ~v_40;
assign v_66689 = v_40;
assign v_66691 = ~v_66690;
assign v_66692 = ~v_45;
assign v_66693 = v_45;
assign v_66695 = ~v_66694;
assign v_66696 = ~v_50;
assign v_66697 = v_50;
assign v_66699 = ~v_66698;
assign v_66700 = ~v_55;
assign v_66701 = v_55;
assign v_66703 = ~v_66702;
assign v_66704 = ~v_60;
assign v_66705 = v_60;
assign v_66707 = ~v_66706;
assign v_66708 = ~v_65;
assign v_66709 = v_65;
assign v_66711 = ~v_66710;
assign v_66712 = ~v_70;
assign v_66713 = v_70;
assign v_66715 = ~v_66714;
assign v_66716 = ~v_75;
assign v_66717 = v_75;
assign v_66719 = ~v_66718;
assign v_66720 = ~v_80;
assign v_66721 = v_80;
assign v_66723 = ~v_66722;
assign v_66724 = ~v_85;
assign v_66725 = v_85;
assign v_66727 = ~v_66726;
assign v_66728 = ~v_90;
assign v_66729 = v_66728;
assign v_66731 = v_66730;
assign v_66733 = v_66724 & v_66732;
assign v_66735 = v_66722;
assign v_66737 = v_66734 & v_66736;
assign v_66739 = v_66720 & v_66738;
assign v_66741 = v_66718;
assign v_66743 = v_66740 & v_66742;
assign v_66745 = v_66716 & v_66744;
assign v_66747 = v_66714;
assign v_66749 = v_66746 & v_66748;
assign v_66751 = v_66712 & v_66750;
assign v_66753 = v_66710;
assign v_66755 = v_66752 & v_66754;
assign v_66757 = v_66708 & v_66756;
assign v_66759 = v_66706;
assign v_66761 = v_66758 & v_66760;
assign v_66763 = v_66704 & v_66762;
assign v_66765 = v_66702;
assign v_66767 = v_66764 & v_66766;
assign v_66769 = v_66700 & v_66768;
assign v_66771 = v_66698;
assign v_66773 = v_66770 & v_66772;
assign v_66775 = v_66696 & v_66774;
assign v_66777 = v_66694;
assign v_66779 = v_66776 & v_66778;
assign v_66781 = v_66692 & v_66780;
assign v_66783 = v_66690;
assign v_66785 = v_66782 & v_66784;
assign v_66787 = v_66688 & v_66786;
assign v_66789 = v_66686;
assign v_66791 = v_66788 & v_66790;
assign v_66793 = v_66684 & v_66792;
assign v_66795 = v_66682;
assign v_66797 = v_66794 & v_66796;
assign v_66799 = v_66680 & v_66798;
assign v_66801 = v_66678;
assign v_66803 = v_66800 & v_66802;
assign v_66805 = v_66676 & v_66804;
assign v_66807 = v_23;
assign v_66809 = v_66806 & v_66808;
assign v_66811 = v_66672 & v_66810;
assign v_66813 = v_18;
assign v_66815 = v_66812 & v_66814;
assign v_66817 = v_66668 & v_66816;
assign v_66819 = v_13;
assign v_66821 = v_66818 & v_66820;
assign v_66823 = v_66664 & v_66822;
assign v_66825 = v_6;
assign v_66827 = v_66824 & v_66826;
assign v_66829 = ~v_66828;
assign v_66831 = v_66726;
assign v_66832 = v_90;
assign v_66833 = v_66832;
assign v_66834 = v_66831 & v_66833;
assign v_66835 = v_66834;
assign v_66836 = v_66724 & v_66835;
assign v_66838 = v_66735 & v_66837;
assign v_66839 = v_66723 & v_66835;
assign v_66841 = v_66720 & v_66840;
assign v_66843 = v_66741 & v_66842;
assign v_66844 = v_66719 & v_66840;
assign v_66846 = v_66716 & v_66845;
assign v_66848 = v_66747 & v_66847;
assign v_66849 = v_66715 & v_66845;
assign v_66851 = v_66712 & v_66850;
assign v_66853 = v_66753 & v_66852;
assign v_66854 = v_66711 & v_66850;
assign v_66856 = v_66708 & v_66855;
assign v_66858 = v_66759 & v_66857;
assign v_66859 = v_66707 & v_66855;
assign v_66861 = v_66704 & v_66860;
assign v_66863 = v_66765 & v_66862;
assign v_66864 = v_66703 & v_66860;
assign v_66866 = v_66700 & v_66865;
assign v_66868 = v_66771 & v_66867;
assign v_66869 = v_66699 & v_66865;
assign v_66871 = v_66696 & v_66870;
assign v_66873 = v_66777 & v_66872;
assign v_66874 = v_66695 & v_66870;
assign v_66876 = v_66692 & v_66875;
assign v_66878 = v_66783 & v_66877;
assign v_66879 = v_66691 & v_66875;
assign v_66881 = v_66688 & v_66880;
assign v_66883 = v_66789 & v_66882;
assign v_66884 = v_66687 & v_66880;
assign v_66886 = v_66684 & v_66885;
assign v_66888 = v_66795 & v_66887;
assign v_66889 = v_66683 & v_66885;
assign v_66891 = v_66680 & v_66890;
assign v_66893 = v_66801 & v_66892;
assign v_66894 = v_66679 & v_66890;
assign v_66896 = v_66676 & v_66895;
assign v_66898 = v_66807 & v_66897;
assign v_66899 = v_66674 & v_66895;
assign v_66901 = v_66672 & v_66900;
assign v_66903 = v_66813 & v_66902;
assign v_66904 = v_66670 & v_66900;
assign v_66906 = v_66668 & v_66905;
assign v_66908 = v_66819 & v_66907;
assign v_66909 = v_66666 & v_66905;
assign v_66911 = v_66664 & v_66910;
assign v_66913 = v_66825 & v_66912;
assign v_66914 = v_66662 & v_66910;
assign v_66916 = v_66828;
assign v_66918 = v_66830 & v_66917;
assign v_66919 = v_66918;
assign v_66921 = v_66920;
assign v_66922 = ~v_283;
assign v_66923 = ~v_66663;
assign v_66924 = v_66663;
assign v_66925 = ~v_287;
assign v_66926 = ~v_66667;
assign v_66927 = v_66667;
assign v_66928 = ~v_291;
assign v_66929 = ~v_66671;
assign v_66930 = v_66671;
assign v_66931 = ~v_295;
assign v_66932 = ~v_66675;
assign v_66933 = v_66675;
assign v_66934 = ~v_66678;
assign v_66935 = ~v_300;
assign v_66936 = v_300;
assign v_66937 = ~v_66682;
assign v_66938 = ~v_304;
assign v_66939 = v_304;
assign v_66940 = ~v_66686;
assign v_66941 = ~v_308;
assign v_66942 = v_308;
assign v_66943 = ~v_66690;
assign v_66944 = ~v_312;
assign v_66945 = v_312;
assign v_66946 = ~v_66694;
assign v_66947 = ~v_316;
assign v_66948 = v_316;
assign v_66949 = ~v_66698;
assign v_66950 = ~v_320;
assign v_66951 = v_320;
assign v_66952 = ~v_66702;
assign v_66953 = ~v_324;
assign v_66954 = v_324;
assign v_66955 = ~v_66706;
assign v_66956 = ~v_328;
assign v_66957 = v_328;
assign v_66958 = ~v_66710;
assign v_66959 = ~v_332;
assign v_66960 = v_332;
assign v_66961 = ~v_66714;
assign v_66962 = ~v_336;
assign v_66963 = v_336;
assign v_66964 = ~v_66718;
assign v_66965 = ~v_340;
assign v_66966 = v_340;
assign v_66967 = ~v_66722;
assign v_66968 = ~v_344;
assign v_66969 = v_344;
assign v_66970 = ~v_66726;
assign v_66971 = ~v_348;
assign v_66972 = v_66971;
assign v_66974 = v_66973;
assign v_66976 = v_66968 & v_66975;
assign v_66978 = v_66722;
assign v_66980 = v_66977 & v_66979;
assign v_66982 = v_66965 & v_66981;
assign v_66984 = v_66718;
assign v_66986 = v_66983 & v_66985;
assign v_66988 = v_66962 & v_66987;
assign v_66990 = v_66714;
assign v_66992 = v_66989 & v_66991;
assign v_66994 = v_66959 & v_66993;
assign v_66996 = v_66710;
assign v_66998 = v_66995 & v_66997;
assign v_67000 = v_66956 & v_66999;
assign v_67002 = v_66706;
assign v_67004 = v_67001 & v_67003;
assign v_67006 = v_66953 & v_67005;
assign v_67008 = v_66702;
assign v_67010 = v_67007 & v_67009;
assign v_67012 = v_66950 & v_67011;
assign v_67014 = v_66698;
assign v_67016 = v_67013 & v_67015;
assign v_67018 = v_66947 & v_67017;
assign v_67020 = v_66694;
assign v_67022 = v_67019 & v_67021;
assign v_67024 = v_66944 & v_67023;
assign v_67026 = v_66690;
assign v_67028 = v_67025 & v_67027;
assign v_67030 = v_66941 & v_67029;
assign v_67032 = v_66686;
assign v_67034 = v_67031 & v_67033;
assign v_67036 = v_66938 & v_67035;
assign v_67038 = v_66682;
assign v_67040 = v_67037 & v_67039;
assign v_67042 = v_66935 & v_67041;
assign v_67044 = v_66678;
assign v_67046 = v_67043 & v_67045;
assign v_67048 = v_66932 & v_67047;
assign v_67050 = v_295;
assign v_67052 = v_67049 & v_67051;
assign v_67054 = v_66929 & v_67053;
assign v_67056 = v_291;
assign v_67058 = v_67055 & v_67057;
assign v_67060 = v_66926 & v_67059;
assign v_67062 = v_287;
assign v_67064 = v_67061 & v_67063;
assign v_67066 = v_66923 & v_67065;
assign v_67068 = v_283;
assign v_67070 = v_67067 & v_67069;
assign v_67072 = ~v_67071;
assign v_67074 = v_66726;
assign v_67075 = v_348;
assign v_67076 = v_67075;
assign v_67077 = v_67074 & v_67076;
assign v_67078 = v_67077;
assign v_67079 = v_66968 & v_67078;
assign v_67081 = v_66978 & v_67080;
assign v_67082 = v_66967 & v_67078;
assign v_67084 = v_66965 & v_67083;
assign v_67086 = v_66984 & v_67085;
assign v_67087 = v_66964 & v_67083;
assign v_67089 = v_66962 & v_67088;
assign v_67091 = v_66990 & v_67090;
assign v_67092 = v_66961 & v_67088;
assign v_67094 = v_66959 & v_67093;
assign v_67096 = v_66996 & v_67095;
assign v_67097 = v_66958 & v_67093;
assign v_67099 = v_66956 & v_67098;
assign v_67101 = v_67002 & v_67100;
assign v_67102 = v_66955 & v_67098;
assign v_67104 = v_66953 & v_67103;
assign v_67106 = v_67008 & v_67105;
assign v_67107 = v_66952 & v_67103;
assign v_67109 = v_66950 & v_67108;
assign v_67111 = v_67014 & v_67110;
assign v_67112 = v_66949 & v_67108;
assign v_67114 = v_66947 & v_67113;
assign v_67116 = v_67020 & v_67115;
assign v_67117 = v_66946 & v_67113;
assign v_67119 = v_66944 & v_67118;
assign v_67121 = v_67026 & v_67120;
assign v_67122 = v_66943 & v_67118;
assign v_67124 = v_66941 & v_67123;
assign v_67126 = v_67032 & v_67125;
assign v_67127 = v_66940 & v_67123;
assign v_67129 = v_66938 & v_67128;
assign v_67131 = v_67038 & v_67130;
assign v_67132 = v_66937 & v_67128;
assign v_67134 = v_66935 & v_67133;
assign v_67136 = v_67044 & v_67135;
assign v_67137 = v_66934 & v_67133;
assign v_67139 = v_66932 & v_67138;
assign v_67141 = v_67050 & v_67140;
assign v_67142 = v_66931 & v_67138;
assign v_67144 = v_66929 & v_67143;
assign v_67146 = v_67056 & v_67145;
assign v_67147 = v_66928 & v_67143;
assign v_67149 = v_66926 & v_67148;
assign v_67151 = v_67062 & v_67150;
assign v_67152 = v_66925 & v_67148;
assign v_67154 = v_66923 & v_67153;
assign v_67156 = v_67068 & v_67155;
assign v_67157 = v_66922 & v_67153;
assign v_67159 = v_67071;
assign v_67161 = v_67073 & v_67160;
assign v_67162 = v_67161;
assign v_67164 = v_67163;
assign v_67165 = ~v_543;
assign v_67166 = ~v_66663;
assign v_67167 = v_66663;
assign v_67168 = ~v_547;
assign v_67169 = ~v_66667;
assign v_67170 = v_66667;
assign v_67171 = ~v_551;
assign v_67172 = ~v_66671;
assign v_67173 = v_66671;
assign v_67174 = ~v_555;
assign v_67175 = ~v_66675;
assign v_67176 = v_66675;
assign v_67177 = ~v_66678;
assign v_67178 = ~v_560;
assign v_67179 = v_560;
assign v_67180 = ~v_66682;
assign v_67181 = ~v_564;
assign v_67182 = v_564;
assign v_67183 = ~v_66686;
assign v_67184 = ~v_568;
assign v_67185 = v_568;
assign v_67186 = ~v_66690;
assign v_67187 = ~v_572;
assign v_67188 = v_572;
assign v_67189 = ~v_66694;
assign v_67190 = ~v_576;
assign v_67191 = v_576;
assign v_67192 = ~v_66698;
assign v_67193 = ~v_580;
assign v_67194 = v_580;
assign v_67195 = ~v_66702;
assign v_67196 = ~v_584;
assign v_67197 = v_584;
assign v_67198 = ~v_66706;
assign v_67199 = ~v_588;
assign v_67200 = v_588;
assign v_67201 = ~v_66710;
assign v_67202 = ~v_592;
assign v_67203 = v_592;
assign v_67204 = ~v_66714;
assign v_67205 = ~v_596;
assign v_67206 = v_596;
assign v_67207 = ~v_66718;
assign v_67208 = ~v_600;
assign v_67209 = v_600;
assign v_67210 = ~v_66722;
assign v_67211 = ~v_604;
assign v_67212 = v_604;
assign v_67213 = ~v_66726;
assign v_67214 = ~v_608;
assign v_67215 = v_67214;
assign v_67217 = v_67216;
assign v_67219 = v_67211 & v_67218;
assign v_67221 = v_66722;
assign v_67223 = v_67220 & v_67222;
assign v_67225 = v_67208 & v_67224;
assign v_67227 = v_66718;
assign v_67229 = v_67226 & v_67228;
assign v_67231 = v_67205 & v_67230;
assign v_67233 = v_66714;
assign v_67235 = v_67232 & v_67234;
assign v_67237 = v_67202 & v_67236;
assign v_67239 = v_66710;
assign v_67241 = v_67238 & v_67240;
assign v_67243 = v_67199 & v_67242;
assign v_67245 = v_66706;
assign v_67247 = v_67244 & v_67246;
assign v_67249 = v_67196 & v_67248;
assign v_67251 = v_66702;
assign v_67253 = v_67250 & v_67252;
assign v_67255 = v_67193 & v_67254;
assign v_67257 = v_66698;
assign v_67259 = v_67256 & v_67258;
assign v_67261 = v_67190 & v_67260;
assign v_67263 = v_66694;
assign v_67265 = v_67262 & v_67264;
assign v_67267 = v_67187 & v_67266;
assign v_67269 = v_66690;
assign v_67271 = v_67268 & v_67270;
assign v_67273 = v_67184 & v_67272;
assign v_67275 = v_66686;
assign v_67277 = v_67274 & v_67276;
assign v_67279 = v_67181 & v_67278;
assign v_67281 = v_66682;
assign v_67283 = v_67280 & v_67282;
assign v_67285 = v_67178 & v_67284;
assign v_67287 = v_66678;
assign v_67289 = v_67286 & v_67288;
assign v_67291 = v_67175 & v_67290;
assign v_67293 = v_555;
assign v_67295 = v_67292 & v_67294;
assign v_67297 = v_67172 & v_67296;
assign v_67299 = v_551;
assign v_67301 = v_67298 & v_67300;
assign v_67303 = v_67169 & v_67302;
assign v_67305 = v_547;
assign v_67307 = v_67304 & v_67306;
assign v_67309 = v_67166 & v_67308;
assign v_67311 = v_543;
assign v_67313 = v_67310 & v_67312;
assign v_67315 = ~v_67314;
assign v_67317 = v_66726;
assign v_67318 = v_608;
assign v_67319 = v_67318;
assign v_67320 = v_67317 & v_67319;
assign v_67321 = v_67320;
assign v_67322 = v_67211 & v_67321;
assign v_67324 = v_67221 & v_67323;
assign v_67325 = v_67210 & v_67321;
assign v_67327 = v_67208 & v_67326;
assign v_67329 = v_67227 & v_67328;
assign v_67330 = v_67207 & v_67326;
assign v_67332 = v_67205 & v_67331;
assign v_67334 = v_67233 & v_67333;
assign v_67335 = v_67204 & v_67331;
assign v_67337 = v_67202 & v_67336;
assign v_67339 = v_67239 & v_67338;
assign v_67340 = v_67201 & v_67336;
assign v_67342 = v_67199 & v_67341;
assign v_67344 = v_67245 & v_67343;
assign v_67345 = v_67198 & v_67341;
assign v_67347 = v_67196 & v_67346;
assign v_67349 = v_67251 & v_67348;
assign v_67350 = v_67195 & v_67346;
assign v_67352 = v_67193 & v_67351;
assign v_67354 = v_67257 & v_67353;
assign v_67355 = v_67192 & v_67351;
assign v_67357 = v_67190 & v_67356;
assign v_67359 = v_67263 & v_67358;
assign v_67360 = v_67189 & v_67356;
assign v_67362 = v_67187 & v_67361;
assign v_67364 = v_67269 & v_67363;
assign v_67365 = v_67186 & v_67361;
assign v_67367 = v_67184 & v_67366;
assign v_67369 = v_67275 & v_67368;
assign v_67370 = v_67183 & v_67366;
assign v_67372 = v_67181 & v_67371;
assign v_67374 = v_67281 & v_67373;
assign v_67375 = v_67180 & v_67371;
assign v_67377 = v_67178 & v_67376;
assign v_67379 = v_67287 & v_67378;
assign v_67380 = v_67177 & v_67376;
assign v_67382 = v_67175 & v_67381;
assign v_67384 = v_67293 & v_67383;
assign v_67385 = v_67174 & v_67381;
assign v_67387 = v_67172 & v_67386;
assign v_67389 = v_67299 & v_67388;
assign v_67390 = v_67171 & v_67386;
assign v_67392 = v_67169 & v_67391;
assign v_67394 = v_67305 & v_67393;
assign v_67395 = v_67168 & v_67391;
assign v_67397 = v_67166 & v_67396;
assign v_67399 = v_67311 & v_67398;
assign v_67400 = v_67165 & v_67396;
assign v_67402 = v_67314;
assign v_67404 = v_67316 & v_67403;
assign v_67405 = v_67404;
assign v_67407 = v_67406;
assign v_67408 = ~v_803;
assign v_67409 = ~v_66663;
assign v_67410 = v_66663;
assign v_67411 = ~v_807;
assign v_67412 = ~v_66667;
assign v_67413 = v_66667;
assign v_67414 = ~v_811;
assign v_67415 = ~v_66671;
assign v_67416 = v_66671;
assign v_67417 = ~v_815;
assign v_67418 = ~v_66675;
assign v_67419 = v_66675;
assign v_67420 = ~v_66678;
assign v_67421 = ~v_820;
assign v_67422 = v_820;
assign v_67423 = ~v_66682;
assign v_67424 = ~v_824;
assign v_67425 = v_824;
assign v_67426 = ~v_66686;
assign v_67427 = ~v_828;
assign v_67428 = v_828;
assign v_67429 = ~v_66690;
assign v_67430 = ~v_832;
assign v_67431 = v_832;
assign v_67432 = ~v_66694;
assign v_67433 = ~v_836;
assign v_67434 = v_836;
assign v_67435 = ~v_66698;
assign v_67436 = ~v_840;
assign v_67437 = v_840;
assign v_67438 = ~v_66702;
assign v_67439 = ~v_844;
assign v_67440 = v_844;
assign v_67441 = ~v_66706;
assign v_67442 = ~v_848;
assign v_67443 = v_848;
assign v_67444 = ~v_66710;
assign v_67445 = ~v_852;
assign v_67446 = v_852;
assign v_67447 = ~v_66714;
assign v_67448 = ~v_856;
assign v_67449 = v_856;
assign v_67450 = ~v_66718;
assign v_67451 = ~v_860;
assign v_67452 = v_860;
assign v_67453 = ~v_66722;
assign v_67454 = ~v_864;
assign v_67455 = v_864;
assign v_67456 = ~v_66726;
assign v_67457 = ~v_868;
assign v_67458 = v_67457;
assign v_67460 = v_67459;
assign v_67462 = v_67454 & v_67461;
assign v_67464 = v_66722;
assign v_67466 = v_67463 & v_67465;
assign v_67468 = v_67451 & v_67467;
assign v_67470 = v_66718;
assign v_67472 = v_67469 & v_67471;
assign v_67474 = v_67448 & v_67473;
assign v_67476 = v_66714;
assign v_67478 = v_67475 & v_67477;
assign v_67480 = v_67445 & v_67479;
assign v_67482 = v_66710;
assign v_67484 = v_67481 & v_67483;
assign v_67486 = v_67442 & v_67485;
assign v_67488 = v_66706;
assign v_67490 = v_67487 & v_67489;
assign v_67492 = v_67439 & v_67491;
assign v_67494 = v_66702;
assign v_67496 = v_67493 & v_67495;
assign v_67498 = v_67436 & v_67497;
assign v_67500 = v_66698;
assign v_67502 = v_67499 & v_67501;
assign v_67504 = v_67433 & v_67503;
assign v_67506 = v_66694;
assign v_67508 = v_67505 & v_67507;
assign v_67510 = v_67430 & v_67509;
assign v_67512 = v_66690;
assign v_67514 = v_67511 & v_67513;
assign v_67516 = v_67427 & v_67515;
assign v_67518 = v_66686;
assign v_67520 = v_67517 & v_67519;
assign v_67522 = v_67424 & v_67521;
assign v_67524 = v_66682;
assign v_67526 = v_67523 & v_67525;
assign v_67528 = v_67421 & v_67527;
assign v_67530 = v_66678;
assign v_67532 = v_67529 & v_67531;
assign v_67534 = v_67418 & v_67533;
assign v_67536 = v_815;
assign v_67538 = v_67535 & v_67537;
assign v_67540 = v_67415 & v_67539;
assign v_67542 = v_811;
assign v_67544 = v_67541 & v_67543;
assign v_67546 = v_67412 & v_67545;
assign v_67548 = v_807;
assign v_67550 = v_67547 & v_67549;
assign v_67552 = v_67409 & v_67551;
assign v_67554 = v_803;
assign v_67556 = v_67553 & v_67555;
assign v_67558 = ~v_67557;
assign v_67560 = v_66726;
assign v_67561 = v_868;
assign v_67562 = v_67561;
assign v_67563 = v_67560 & v_67562;
assign v_67564 = v_67563;
assign v_67565 = v_67454 & v_67564;
assign v_67567 = v_67464 & v_67566;
assign v_67568 = v_67453 & v_67564;
assign v_67570 = v_67451 & v_67569;
assign v_67572 = v_67470 & v_67571;
assign v_67573 = v_67450 & v_67569;
assign v_67575 = v_67448 & v_67574;
assign v_67577 = v_67476 & v_67576;
assign v_67578 = v_67447 & v_67574;
assign v_67580 = v_67445 & v_67579;
assign v_67582 = v_67482 & v_67581;
assign v_67583 = v_67444 & v_67579;
assign v_67585 = v_67442 & v_67584;
assign v_67587 = v_67488 & v_67586;
assign v_67588 = v_67441 & v_67584;
assign v_67590 = v_67439 & v_67589;
assign v_67592 = v_67494 & v_67591;
assign v_67593 = v_67438 & v_67589;
assign v_67595 = v_67436 & v_67594;
assign v_67597 = v_67500 & v_67596;
assign v_67598 = v_67435 & v_67594;
assign v_67600 = v_67433 & v_67599;
assign v_67602 = v_67506 & v_67601;
assign v_67603 = v_67432 & v_67599;
assign v_67605 = v_67430 & v_67604;
assign v_67607 = v_67512 & v_67606;
assign v_67608 = v_67429 & v_67604;
assign v_67610 = v_67427 & v_67609;
assign v_67612 = v_67518 & v_67611;
assign v_67613 = v_67426 & v_67609;
assign v_67615 = v_67424 & v_67614;
assign v_67617 = v_67524 & v_67616;
assign v_67618 = v_67423 & v_67614;
assign v_67620 = v_67421 & v_67619;
assign v_67622 = v_67530 & v_67621;
assign v_67623 = v_67420 & v_67619;
assign v_67625 = v_67418 & v_67624;
assign v_67627 = v_67536 & v_67626;
assign v_67628 = v_67417 & v_67624;
assign v_67630 = v_67415 & v_67629;
assign v_67632 = v_67542 & v_67631;
assign v_67633 = v_67414 & v_67629;
assign v_67635 = v_67412 & v_67634;
assign v_67637 = v_67548 & v_67636;
assign v_67638 = v_67411 & v_67634;
assign v_67640 = v_67409 & v_67639;
assign v_67642 = v_67554 & v_67641;
assign v_67643 = v_67408 & v_67639;
assign v_67645 = v_67557;
assign v_67647 = v_67559 & v_67646;
assign v_67648 = v_67647;
assign v_67650 = v_67649;
assign v_67651 = ~v_1063;
assign v_67652 = ~v_66663;
assign v_67653 = v_66663;
assign v_67654 = ~v_1067;
assign v_67655 = ~v_66667;
assign v_67656 = v_66667;
assign v_67657 = ~v_1071;
assign v_67658 = ~v_66671;
assign v_67659 = v_66671;
assign v_67660 = ~v_1075;
assign v_67661 = ~v_66675;
assign v_67662 = v_66675;
assign v_67663 = ~v_66678;
assign v_67664 = ~v_1080;
assign v_67665 = v_1080;
assign v_67666 = ~v_66682;
assign v_67667 = ~v_1084;
assign v_67668 = v_1084;
assign v_67669 = ~v_66686;
assign v_67670 = ~v_1088;
assign v_67671 = v_1088;
assign v_67672 = ~v_66690;
assign v_67673 = ~v_1092;
assign v_67674 = v_1092;
assign v_67675 = ~v_66694;
assign v_67676 = ~v_1096;
assign v_67677 = v_1096;
assign v_67678 = ~v_66698;
assign v_67679 = ~v_1100;
assign v_67680 = v_1100;
assign v_67681 = ~v_66702;
assign v_67682 = ~v_1104;
assign v_67683 = v_1104;
assign v_67684 = ~v_66706;
assign v_67685 = ~v_1108;
assign v_67686 = v_1108;
assign v_67687 = ~v_66710;
assign v_67688 = ~v_1112;
assign v_67689 = v_1112;
assign v_67690 = ~v_66714;
assign v_67691 = ~v_1116;
assign v_67692 = v_1116;
assign v_67693 = ~v_66718;
assign v_67694 = ~v_1120;
assign v_67695 = v_1120;
assign v_67696 = ~v_66722;
assign v_67697 = ~v_1124;
assign v_67698 = v_1124;
assign v_67699 = ~v_66726;
assign v_67700 = ~v_1128;
assign v_67701 = v_67700;
assign v_67703 = v_67702;
assign v_67705 = v_67697 & v_67704;
assign v_67707 = v_66722;
assign v_67709 = v_67706 & v_67708;
assign v_67711 = v_67694 & v_67710;
assign v_67713 = v_66718;
assign v_67715 = v_67712 & v_67714;
assign v_67717 = v_67691 & v_67716;
assign v_67719 = v_66714;
assign v_67721 = v_67718 & v_67720;
assign v_67723 = v_67688 & v_67722;
assign v_67725 = v_66710;
assign v_67727 = v_67724 & v_67726;
assign v_67729 = v_67685 & v_67728;
assign v_67731 = v_66706;
assign v_67733 = v_67730 & v_67732;
assign v_67735 = v_67682 & v_67734;
assign v_67737 = v_66702;
assign v_67739 = v_67736 & v_67738;
assign v_67741 = v_67679 & v_67740;
assign v_67743 = v_66698;
assign v_67745 = v_67742 & v_67744;
assign v_67747 = v_67676 & v_67746;
assign v_67749 = v_66694;
assign v_67751 = v_67748 & v_67750;
assign v_67753 = v_67673 & v_67752;
assign v_67755 = v_66690;
assign v_67757 = v_67754 & v_67756;
assign v_67759 = v_67670 & v_67758;
assign v_67761 = v_66686;
assign v_67763 = v_67760 & v_67762;
assign v_67765 = v_67667 & v_67764;
assign v_67767 = v_66682;
assign v_67769 = v_67766 & v_67768;
assign v_67771 = v_67664 & v_67770;
assign v_67773 = v_66678;
assign v_67775 = v_67772 & v_67774;
assign v_67777 = v_67661 & v_67776;
assign v_67779 = v_1075;
assign v_67781 = v_67778 & v_67780;
assign v_67783 = v_67658 & v_67782;
assign v_67785 = v_1071;
assign v_67787 = v_67784 & v_67786;
assign v_67789 = v_67655 & v_67788;
assign v_67791 = v_1067;
assign v_67793 = v_67790 & v_67792;
assign v_67795 = v_67652 & v_67794;
assign v_67797 = v_1063;
assign v_67799 = v_67796 & v_67798;
assign v_67801 = ~v_67800;
assign v_67803 = v_66726;
assign v_67804 = v_1128;
assign v_67805 = v_67804;
assign v_67806 = v_67803 & v_67805;
assign v_67807 = v_67806;
assign v_67808 = v_67697 & v_67807;
assign v_67810 = v_67707 & v_67809;
assign v_67811 = v_67696 & v_67807;
assign v_67813 = v_67694 & v_67812;
assign v_67815 = v_67713 & v_67814;
assign v_67816 = v_67693 & v_67812;
assign v_67818 = v_67691 & v_67817;
assign v_67820 = v_67719 & v_67819;
assign v_67821 = v_67690 & v_67817;
assign v_67823 = v_67688 & v_67822;
assign v_67825 = v_67725 & v_67824;
assign v_67826 = v_67687 & v_67822;
assign v_67828 = v_67685 & v_67827;
assign v_67830 = v_67731 & v_67829;
assign v_67831 = v_67684 & v_67827;
assign v_67833 = v_67682 & v_67832;
assign v_67835 = v_67737 & v_67834;
assign v_67836 = v_67681 & v_67832;
assign v_67838 = v_67679 & v_67837;
assign v_67840 = v_67743 & v_67839;
assign v_67841 = v_67678 & v_67837;
assign v_67843 = v_67676 & v_67842;
assign v_67845 = v_67749 & v_67844;
assign v_67846 = v_67675 & v_67842;
assign v_67848 = v_67673 & v_67847;
assign v_67850 = v_67755 & v_67849;
assign v_67851 = v_67672 & v_67847;
assign v_67853 = v_67670 & v_67852;
assign v_67855 = v_67761 & v_67854;
assign v_67856 = v_67669 & v_67852;
assign v_67858 = v_67667 & v_67857;
assign v_67860 = v_67767 & v_67859;
assign v_67861 = v_67666 & v_67857;
assign v_67863 = v_67664 & v_67862;
assign v_67865 = v_67773 & v_67864;
assign v_67866 = v_67663 & v_67862;
assign v_67868 = v_67661 & v_67867;
assign v_67870 = v_67779 & v_67869;
assign v_67871 = v_67660 & v_67867;
assign v_67873 = v_67658 & v_67872;
assign v_67875 = v_67785 & v_67874;
assign v_67876 = v_67657 & v_67872;
assign v_67878 = v_67655 & v_67877;
assign v_67880 = v_67791 & v_67879;
assign v_67881 = v_67654 & v_67877;
assign v_67883 = v_67652 & v_67882;
assign v_67885 = v_67797 & v_67884;
assign v_67886 = v_67651 & v_67882;
assign v_67888 = v_67800;
assign v_67890 = v_67802 & v_67889;
assign v_67891 = v_67890;
assign v_67893 = v_67892;
assign v_67894 = ~v_1323;
assign v_67895 = ~v_66663;
assign v_67896 = v_66663;
assign v_67897 = ~v_1327;
assign v_67898 = ~v_66667;
assign v_67899 = v_66667;
assign v_67900 = ~v_1331;
assign v_67901 = ~v_66671;
assign v_67902 = v_66671;
assign v_67903 = ~v_1335;
assign v_67904 = ~v_66675;
assign v_67905 = v_66675;
assign v_67906 = ~v_66678;
assign v_67907 = ~v_1340;
assign v_67908 = v_1340;
assign v_67909 = ~v_66682;
assign v_67910 = ~v_1344;
assign v_67911 = v_1344;
assign v_67912 = ~v_66686;
assign v_67913 = ~v_1348;
assign v_67914 = v_1348;
assign v_67915 = ~v_66690;
assign v_67916 = ~v_1352;
assign v_67917 = v_1352;
assign v_67918 = ~v_66694;
assign v_67919 = ~v_1356;
assign v_67920 = v_1356;
assign v_67921 = ~v_66698;
assign v_67922 = ~v_1360;
assign v_67923 = v_1360;
assign v_67924 = ~v_66702;
assign v_67925 = ~v_1364;
assign v_67926 = v_1364;
assign v_67927 = ~v_66706;
assign v_67928 = ~v_1368;
assign v_67929 = v_1368;
assign v_67930 = ~v_66710;
assign v_67931 = ~v_1372;
assign v_67932 = v_1372;
assign v_67933 = ~v_66714;
assign v_67934 = ~v_1376;
assign v_67935 = v_1376;
assign v_67936 = ~v_66718;
assign v_67937 = ~v_1380;
assign v_67938 = v_1380;
assign v_67939 = ~v_66722;
assign v_67940 = ~v_1384;
assign v_67941 = v_1384;
assign v_67942 = ~v_66726;
assign v_67943 = ~v_1388;
assign v_67944 = v_67943;
assign v_67946 = v_67945;
assign v_67948 = v_67940 & v_67947;
assign v_67950 = v_66722;
assign v_67952 = v_67949 & v_67951;
assign v_67954 = v_67937 & v_67953;
assign v_67956 = v_66718;
assign v_67958 = v_67955 & v_67957;
assign v_67960 = v_67934 & v_67959;
assign v_67962 = v_66714;
assign v_67964 = v_67961 & v_67963;
assign v_67966 = v_67931 & v_67965;
assign v_67968 = v_66710;
assign v_67970 = v_67967 & v_67969;
assign v_67972 = v_67928 & v_67971;
assign v_67974 = v_66706;
assign v_67976 = v_67973 & v_67975;
assign v_67978 = v_67925 & v_67977;
assign v_67980 = v_66702;
assign v_67982 = v_67979 & v_67981;
assign v_67984 = v_67922 & v_67983;
assign v_67986 = v_66698;
assign v_67988 = v_67985 & v_67987;
assign v_67990 = v_67919 & v_67989;
assign v_67992 = v_66694;
assign v_67994 = v_67991 & v_67993;
assign v_67996 = v_67916 & v_67995;
assign v_67998 = v_66690;
assign v_68000 = v_67997 & v_67999;
assign v_68002 = v_67913 & v_68001;
assign v_68004 = v_66686;
assign v_68006 = v_68003 & v_68005;
assign v_68008 = v_67910 & v_68007;
assign v_68010 = v_66682;
assign v_68012 = v_68009 & v_68011;
assign v_68014 = v_67907 & v_68013;
assign v_68016 = v_66678;
assign v_68018 = v_68015 & v_68017;
assign v_68020 = v_67904 & v_68019;
assign v_68022 = v_1335;
assign v_68024 = v_68021 & v_68023;
assign v_68026 = v_67901 & v_68025;
assign v_68028 = v_1331;
assign v_68030 = v_68027 & v_68029;
assign v_68032 = v_67898 & v_68031;
assign v_68034 = v_1327;
assign v_68036 = v_68033 & v_68035;
assign v_68038 = v_67895 & v_68037;
assign v_68040 = v_1323;
assign v_68042 = v_68039 & v_68041;
assign v_68044 = ~v_68043;
assign v_68046 = v_66726;
assign v_68047 = v_1388;
assign v_68048 = v_68047;
assign v_68049 = v_68046 & v_68048;
assign v_68050 = v_68049;
assign v_68051 = v_67940 & v_68050;
assign v_68053 = v_67950 & v_68052;
assign v_68054 = v_67939 & v_68050;
assign v_68056 = v_67937 & v_68055;
assign v_68058 = v_67956 & v_68057;
assign v_68059 = v_67936 & v_68055;
assign v_68061 = v_67934 & v_68060;
assign v_68063 = v_67962 & v_68062;
assign v_68064 = v_67933 & v_68060;
assign v_68066 = v_67931 & v_68065;
assign v_68068 = v_67968 & v_68067;
assign v_68069 = v_67930 & v_68065;
assign v_68071 = v_67928 & v_68070;
assign v_68073 = v_67974 & v_68072;
assign v_68074 = v_67927 & v_68070;
assign v_68076 = v_67925 & v_68075;
assign v_68078 = v_67980 & v_68077;
assign v_68079 = v_67924 & v_68075;
assign v_68081 = v_67922 & v_68080;
assign v_68083 = v_67986 & v_68082;
assign v_68084 = v_67921 & v_68080;
assign v_68086 = v_67919 & v_68085;
assign v_68088 = v_67992 & v_68087;
assign v_68089 = v_67918 & v_68085;
assign v_68091 = v_67916 & v_68090;
assign v_68093 = v_67998 & v_68092;
assign v_68094 = v_67915 & v_68090;
assign v_68096 = v_67913 & v_68095;
assign v_68098 = v_68004 & v_68097;
assign v_68099 = v_67912 & v_68095;
assign v_68101 = v_67910 & v_68100;
assign v_68103 = v_68010 & v_68102;
assign v_68104 = v_67909 & v_68100;
assign v_68106 = v_67907 & v_68105;
assign v_68108 = v_68016 & v_68107;
assign v_68109 = v_67906 & v_68105;
assign v_68111 = v_67904 & v_68110;
assign v_68113 = v_68022 & v_68112;
assign v_68114 = v_67903 & v_68110;
assign v_68116 = v_67901 & v_68115;
assign v_68118 = v_68028 & v_68117;
assign v_68119 = v_67900 & v_68115;
assign v_68121 = v_67898 & v_68120;
assign v_68123 = v_68034 & v_68122;
assign v_68124 = v_67897 & v_68120;
assign v_68126 = v_67895 & v_68125;
assign v_68128 = v_68040 & v_68127;
assign v_68129 = v_67894 & v_68125;
assign v_68131 = v_68043;
assign v_68133 = v_68045 & v_68132;
assign v_68134 = v_68133;
assign v_68136 = v_68135;
assign v_68137 = ~v_1583;
assign v_68138 = ~v_66663;
assign v_68139 = v_66663;
assign v_68140 = ~v_1587;
assign v_68141 = ~v_66667;
assign v_68142 = v_66667;
assign v_68143 = ~v_1591;
assign v_68144 = ~v_66671;
assign v_68145 = v_66671;
assign v_68146 = ~v_1595;
assign v_68147 = ~v_66675;
assign v_68148 = v_66675;
assign v_68149 = ~v_66678;
assign v_68150 = ~v_1600;
assign v_68151 = v_1600;
assign v_68152 = ~v_66682;
assign v_68153 = ~v_1604;
assign v_68154 = v_1604;
assign v_68155 = ~v_66686;
assign v_68156 = ~v_1608;
assign v_68157 = v_1608;
assign v_68158 = ~v_66690;
assign v_68159 = ~v_1612;
assign v_68160 = v_1612;
assign v_68161 = ~v_66694;
assign v_68162 = ~v_1616;
assign v_68163 = v_1616;
assign v_68164 = ~v_66698;
assign v_68165 = ~v_1620;
assign v_68166 = v_1620;
assign v_68167 = ~v_66702;
assign v_68168 = ~v_1624;
assign v_68169 = v_1624;
assign v_68170 = ~v_66706;
assign v_68171 = ~v_1628;
assign v_68172 = v_1628;
assign v_68173 = ~v_66710;
assign v_68174 = ~v_1632;
assign v_68175 = v_1632;
assign v_68176 = ~v_66714;
assign v_68177 = ~v_1636;
assign v_68178 = v_1636;
assign v_68179 = ~v_66718;
assign v_68180 = ~v_1640;
assign v_68181 = v_1640;
assign v_68182 = ~v_66722;
assign v_68183 = ~v_1644;
assign v_68184 = v_1644;
assign v_68185 = ~v_66726;
assign v_68186 = ~v_1648;
assign v_68187 = v_68186;
assign v_68189 = v_68188;
assign v_68191 = v_68183 & v_68190;
assign v_68193 = v_66722;
assign v_68195 = v_68192 & v_68194;
assign v_68197 = v_68180 & v_68196;
assign v_68199 = v_66718;
assign v_68201 = v_68198 & v_68200;
assign v_68203 = v_68177 & v_68202;
assign v_68205 = v_66714;
assign v_68207 = v_68204 & v_68206;
assign v_68209 = v_68174 & v_68208;
assign v_68211 = v_66710;
assign v_68213 = v_68210 & v_68212;
assign v_68215 = v_68171 & v_68214;
assign v_68217 = v_66706;
assign v_68219 = v_68216 & v_68218;
assign v_68221 = v_68168 & v_68220;
assign v_68223 = v_66702;
assign v_68225 = v_68222 & v_68224;
assign v_68227 = v_68165 & v_68226;
assign v_68229 = v_66698;
assign v_68231 = v_68228 & v_68230;
assign v_68233 = v_68162 & v_68232;
assign v_68235 = v_66694;
assign v_68237 = v_68234 & v_68236;
assign v_68239 = v_68159 & v_68238;
assign v_68241 = v_66690;
assign v_68243 = v_68240 & v_68242;
assign v_68245 = v_68156 & v_68244;
assign v_68247 = v_66686;
assign v_68249 = v_68246 & v_68248;
assign v_68251 = v_68153 & v_68250;
assign v_68253 = v_66682;
assign v_68255 = v_68252 & v_68254;
assign v_68257 = v_68150 & v_68256;
assign v_68259 = v_66678;
assign v_68261 = v_68258 & v_68260;
assign v_68263 = v_68147 & v_68262;
assign v_68265 = v_1595;
assign v_68267 = v_68264 & v_68266;
assign v_68269 = v_68144 & v_68268;
assign v_68271 = v_1591;
assign v_68273 = v_68270 & v_68272;
assign v_68275 = v_68141 & v_68274;
assign v_68277 = v_1587;
assign v_68279 = v_68276 & v_68278;
assign v_68281 = v_68138 & v_68280;
assign v_68283 = v_1583;
assign v_68285 = v_68282 & v_68284;
assign v_68287 = ~v_68286;
assign v_68289 = v_66726;
assign v_68290 = v_1648;
assign v_68291 = v_68290;
assign v_68292 = v_68289 & v_68291;
assign v_68293 = v_68292;
assign v_68294 = v_68183 & v_68293;
assign v_68296 = v_68193 & v_68295;
assign v_68297 = v_68182 & v_68293;
assign v_68299 = v_68180 & v_68298;
assign v_68301 = v_68199 & v_68300;
assign v_68302 = v_68179 & v_68298;
assign v_68304 = v_68177 & v_68303;
assign v_68306 = v_68205 & v_68305;
assign v_68307 = v_68176 & v_68303;
assign v_68309 = v_68174 & v_68308;
assign v_68311 = v_68211 & v_68310;
assign v_68312 = v_68173 & v_68308;
assign v_68314 = v_68171 & v_68313;
assign v_68316 = v_68217 & v_68315;
assign v_68317 = v_68170 & v_68313;
assign v_68319 = v_68168 & v_68318;
assign v_68321 = v_68223 & v_68320;
assign v_68322 = v_68167 & v_68318;
assign v_68324 = v_68165 & v_68323;
assign v_68326 = v_68229 & v_68325;
assign v_68327 = v_68164 & v_68323;
assign v_68329 = v_68162 & v_68328;
assign v_68331 = v_68235 & v_68330;
assign v_68332 = v_68161 & v_68328;
assign v_68334 = v_68159 & v_68333;
assign v_68336 = v_68241 & v_68335;
assign v_68337 = v_68158 & v_68333;
assign v_68339 = v_68156 & v_68338;
assign v_68341 = v_68247 & v_68340;
assign v_68342 = v_68155 & v_68338;
assign v_68344 = v_68153 & v_68343;
assign v_68346 = v_68253 & v_68345;
assign v_68347 = v_68152 & v_68343;
assign v_68349 = v_68150 & v_68348;
assign v_68351 = v_68259 & v_68350;
assign v_68352 = v_68149 & v_68348;
assign v_68354 = v_68147 & v_68353;
assign v_68356 = v_68265 & v_68355;
assign v_68357 = v_68146 & v_68353;
assign v_68359 = v_68144 & v_68358;
assign v_68361 = v_68271 & v_68360;
assign v_68362 = v_68143 & v_68358;
assign v_68364 = v_68141 & v_68363;
assign v_68366 = v_68277 & v_68365;
assign v_68367 = v_68140 & v_68363;
assign v_68369 = v_68138 & v_68368;
assign v_68371 = v_68283 & v_68370;
assign v_68372 = v_68137 & v_68368;
assign v_68374 = v_68286;
assign v_68376 = v_68288 & v_68375;
assign v_68377 = v_68376;
assign v_68379 = v_68378;
assign v_68380 = ~v_1843;
assign v_68381 = ~v_66663;
assign v_68382 = v_66663;
assign v_68383 = ~v_1847;
assign v_68384 = ~v_66667;
assign v_68385 = v_66667;
assign v_68386 = ~v_1851;
assign v_68387 = ~v_66671;
assign v_68388 = v_66671;
assign v_68389 = ~v_1855;
assign v_68390 = ~v_66675;
assign v_68391 = v_66675;
assign v_68392 = ~v_66678;
assign v_68393 = ~v_1860;
assign v_68394 = v_1860;
assign v_68395 = ~v_66682;
assign v_68396 = ~v_1864;
assign v_68397 = v_1864;
assign v_68398 = ~v_66686;
assign v_68399 = ~v_1868;
assign v_68400 = v_1868;
assign v_68401 = ~v_66690;
assign v_68402 = ~v_1872;
assign v_68403 = v_1872;
assign v_68404 = ~v_66694;
assign v_68405 = ~v_1876;
assign v_68406 = v_1876;
assign v_68407 = ~v_66698;
assign v_68408 = ~v_1880;
assign v_68409 = v_1880;
assign v_68410 = ~v_66702;
assign v_68411 = ~v_1884;
assign v_68412 = v_1884;
assign v_68413 = ~v_66706;
assign v_68414 = ~v_1888;
assign v_68415 = v_1888;
assign v_68416 = ~v_66710;
assign v_68417 = ~v_1892;
assign v_68418 = v_1892;
assign v_68419 = ~v_66714;
assign v_68420 = ~v_1896;
assign v_68421 = v_1896;
assign v_68422 = ~v_66718;
assign v_68423 = ~v_1900;
assign v_68424 = v_1900;
assign v_68425 = ~v_66722;
assign v_68426 = ~v_1904;
assign v_68427 = v_1904;
assign v_68428 = ~v_66726;
assign v_68429 = ~v_1908;
assign v_68430 = v_68429;
assign v_68432 = v_68431;
assign v_68434 = v_68426 & v_68433;
assign v_68436 = v_66722;
assign v_68438 = v_68435 & v_68437;
assign v_68440 = v_68423 & v_68439;
assign v_68442 = v_66718;
assign v_68444 = v_68441 & v_68443;
assign v_68446 = v_68420 & v_68445;
assign v_68448 = v_66714;
assign v_68450 = v_68447 & v_68449;
assign v_68452 = v_68417 & v_68451;
assign v_68454 = v_66710;
assign v_68456 = v_68453 & v_68455;
assign v_68458 = v_68414 & v_68457;
assign v_68460 = v_66706;
assign v_68462 = v_68459 & v_68461;
assign v_68464 = v_68411 & v_68463;
assign v_68466 = v_66702;
assign v_68468 = v_68465 & v_68467;
assign v_68470 = v_68408 & v_68469;
assign v_68472 = v_66698;
assign v_68474 = v_68471 & v_68473;
assign v_68476 = v_68405 & v_68475;
assign v_68478 = v_66694;
assign v_68480 = v_68477 & v_68479;
assign v_68482 = v_68402 & v_68481;
assign v_68484 = v_66690;
assign v_68486 = v_68483 & v_68485;
assign v_68488 = v_68399 & v_68487;
assign v_68490 = v_66686;
assign v_68492 = v_68489 & v_68491;
assign v_68494 = v_68396 & v_68493;
assign v_68496 = v_66682;
assign v_68498 = v_68495 & v_68497;
assign v_68500 = v_68393 & v_68499;
assign v_68502 = v_66678;
assign v_68504 = v_68501 & v_68503;
assign v_68506 = v_68390 & v_68505;
assign v_68508 = v_1855;
assign v_68510 = v_68507 & v_68509;
assign v_68512 = v_68387 & v_68511;
assign v_68514 = v_1851;
assign v_68516 = v_68513 & v_68515;
assign v_68518 = v_68384 & v_68517;
assign v_68520 = v_1847;
assign v_68522 = v_68519 & v_68521;
assign v_68524 = v_68381 & v_68523;
assign v_68526 = v_1843;
assign v_68528 = v_68525 & v_68527;
assign v_68530 = ~v_68529;
assign v_68532 = v_66726;
assign v_68533 = v_1908;
assign v_68534 = v_68533;
assign v_68535 = v_68532 & v_68534;
assign v_68536 = v_68535;
assign v_68537 = v_68426 & v_68536;
assign v_68539 = v_68436 & v_68538;
assign v_68540 = v_68425 & v_68536;
assign v_68542 = v_68423 & v_68541;
assign v_68544 = v_68442 & v_68543;
assign v_68545 = v_68422 & v_68541;
assign v_68547 = v_68420 & v_68546;
assign v_68549 = v_68448 & v_68548;
assign v_68550 = v_68419 & v_68546;
assign v_68552 = v_68417 & v_68551;
assign v_68554 = v_68454 & v_68553;
assign v_68555 = v_68416 & v_68551;
assign v_68557 = v_68414 & v_68556;
assign v_68559 = v_68460 & v_68558;
assign v_68560 = v_68413 & v_68556;
assign v_68562 = v_68411 & v_68561;
assign v_68564 = v_68466 & v_68563;
assign v_68565 = v_68410 & v_68561;
assign v_68567 = v_68408 & v_68566;
assign v_68569 = v_68472 & v_68568;
assign v_68570 = v_68407 & v_68566;
assign v_68572 = v_68405 & v_68571;
assign v_68574 = v_68478 & v_68573;
assign v_68575 = v_68404 & v_68571;
assign v_68577 = v_68402 & v_68576;
assign v_68579 = v_68484 & v_68578;
assign v_68580 = v_68401 & v_68576;
assign v_68582 = v_68399 & v_68581;
assign v_68584 = v_68490 & v_68583;
assign v_68585 = v_68398 & v_68581;
assign v_68587 = v_68396 & v_68586;
assign v_68589 = v_68496 & v_68588;
assign v_68590 = v_68395 & v_68586;
assign v_68592 = v_68393 & v_68591;
assign v_68594 = v_68502 & v_68593;
assign v_68595 = v_68392 & v_68591;
assign v_68597 = v_68390 & v_68596;
assign v_68599 = v_68508 & v_68598;
assign v_68600 = v_68389 & v_68596;
assign v_68602 = v_68387 & v_68601;
assign v_68604 = v_68514 & v_68603;
assign v_68605 = v_68386 & v_68601;
assign v_68607 = v_68384 & v_68606;
assign v_68609 = v_68520 & v_68608;
assign v_68610 = v_68383 & v_68606;
assign v_68612 = v_68381 & v_68611;
assign v_68614 = v_68526 & v_68613;
assign v_68615 = v_68380 & v_68611;
assign v_68617 = v_68529;
assign v_68619 = v_68531 & v_68618;
assign v_68620 = v_68619;
assign v_68622 = v_68621;
assign v_68623 = ~v_2103;
assign v_68624 = ~v_66663;
assign v_68625 = v_66663;
assign v_68626 = ~v_2107;
assign v_68627 = ~v_66667;
assign v_68628 = v_66667;
assign v_68629 = ~v_2111;
assign v_68630 = ~v_66671;
assign v_68631 = v_66671;
assign v_68632 = ~v_2115;
assign v_68633 = ~v_66675;
assign v_68634 = v_66675;
assign v_68635 = ~v_66678;
assign v_68636 = ~v_2120;
assign v_68637 = v_2120;
assign v_68638 = ~v_66682;
assign v_68639 = ~v_2124;
assign v_68640 = v_2124;
assign v_68641 = ~v_66686;
assign v_68642 = ~v_2128;
assign v_68643 = v_2128;
assign v_68644 = ~v_66690;
assign v_68645 = ~v_2132;
assign v_68646 = v_2132;
assign v_68647 = ~v_66694;
assign v_68648 = ~v_2136;
assign v_68649 = v_2136;
assign v_68650 = ~v_66698;
assign v_68651 = ~v_2140;
assign v_68652 = v_2140;
assign v_68653 = ~v_66702;
assign v_68654 = ~v_2144;
assign v_68655 = v_2144;
assign v_68656 = ~v_66706;
assign v_68657 = ~v_2148;
assign v_68658 = v_2148;
assign v_68659 = ~v_66710;
assign v_68660 = ~v_2152;
assign v_68661 = v_2152;
assign v_68662 = ~v_66714;
assign v_68663 = ~v_2156;
assign v_68664 = v_2156;
assign v_68665 = ~v_66718;
assign v_68666 = ~v_2160;
assign v_68667 = v_2160;
assign v_68668 = ~v_66722;
assign v_68669 = ~v_2164;
assign v_68670 = v_2164;
assign v_68671 = ~v_66726;
assign v_68672 = ~v_2168;
assign v_68673 = v_68672;
assign v_68675 = v_68674;
assign v_68677 = v_68669 & v_68676;
assign v_68679 = v_66722;
assign v_68681 = v_68678 & v_68680;
assign v_68683 = v_68666 & v_68682;
assign v_68685 = v_66718;
assign v_68687 = v_68684 & v_68686;
assign v_68689 = v_68663 & v_68688;
assign v_68691 = v_66714;
assign v_68693 = v_68690 & v_68692;
assign v_68695 = v_68660 & v_68694;
assign v_68697 = v_66710;
assign v_68699 = v_68696 & v_68698;
assign v_68701 = v_68657 & v_68700;
assign v_68703 = v_66706;
assign v_68705 = v_68702 & v_68704;
assign v_68707 = v_68654 & v_68706;
assign v_68709 = v_66702;
assign v_68711 = v_68708 & v_68710;
assign v_68713 = v_68651 & v_68712;
assign v_68715 = v_66698;
assign v_68717 = v_68714 & v_68716;
assign v_68719 = v_68648 & v_68718;
assign v_68721 = v_66694;
assign v_68723 = v_68720 & v_68722;
assign v_68725 = v_68645 & v_68724;
assign v_68727 = v_66690;
assign v_68729 = v_68726 & v_68728;
assign v_68731 = v_68642 & v_68730;
assign v_68733 = v_66686;
assign v_68735 = v_68732 & v_68734;
assign v_68737 = v_68639 & v_68736;
assign v_68739 = v_66682;
assign v_68741 = v_68738 & v_68740;
assign v_68743 = v_68636 & v_68742;
assign v_68745 = v_66678;
assign v_68747 = v_68744 & v_68746;
assign v_68749 = v_68633 & v_68748;
assign v_68751 = v_2115;
assign v_68753 = v_68750 & v_68752;
assign v_68755 = v_68630 & v_68754;
assign v_68757 = v_2111;
assign v_68759 = v_68756 & v_68758;
assign v_68761 = v_68627 & v_68760;
assign v_68763 = v_2107;
assign v_68765 = v_68762 & v_68764;
assign v_68767 = v_68624 & v_68766;
assign v_68769 = v_2103;
assign v_68771 = v_68768 & v_68770;
assign v_68773 = ~v_68772;
assign v_68775 = v_66726;
assign v_68776 = v_2168;
assign v_68777 = v_68776;
assign v_68778 = v_68775 & v_68777;
assign v_68779 = v_68778;
assign v_68780 = v_68669 & v_68779;
assign v_68782 = v_68679 & v_68781;
assign v_68783 = v_68668 & v_68779;
assign v_68785 = v_68666 & v_68784;
assign v_68787 = v_68685 & v_68786;
assign v_68788 = v_68665 & v_68784;
assign v_68790 = v_68663 & v_68789;
assign v_68792 = v_68691 & v_68791;
assign v_68793 = v_68662 & v_68789;
assign v_68795 = v_68660 & v_68794;
assign v_68797 = v_68697 & v_68796;
assign v_68798 = v_68659 & v_68794;
assign v_68800 = v_68657 & v_68799;
assign v_68802 = v_68703 & v_68801;
assign v_68803 = v_68656 & v_68799;
assign v_68805 = v_68654 & v_68804;
assign v_68807 = v_68709 & v_68806;
assign v_68808 = v_68653 & v_68804;
assign v_68810 = v_68651 & v_68809;
assign v_68812 = v_68715 & v_68811;
assign v_68813 = v_68650 & v_68809;
assign v_68815 = v_68648 & v_68814;
assign v_68817 = v_68721 & v_68816;
assign v_68818 = v_68647 & v_68814;
assign v_68820 = v_68645 & v_68819;
assign v_68822 = v_68727 & v_68821;
assign v_68823 = v_68644 & v_68819;
assign v_68825 = v_68642 & v_68824;
assign v_68827 = v_68733 & v_68826;
assign v_68828 = v_68641 & v_68824;
assign v_68830 = v_68639 & v_68829;
assign v_68832 = v_68739 & v_68831;
assign v_68833 = v_68638 & v_68829;
assign v_68835 = v_68636 & v_68834;
assign v_68837 = v_68745 & v_68836;
assign v_68838 = v_68635 & v_68834;
assign v_68840 = v_68633 & v_68839;
assign v_68842 = v_68751 & v_68841;
assign v_68843 = v_68632 & v_68839;
assign v_68845 = v_68630 & v_68844;
assign v_68847 = v_68757 & v_68846;
assign v_68848 = v_68629 & v_68844;
assign v_68850 = v_68627 & v_68849;
assign v_68852 = v_68763 & v_68851;
assign v_68853 = v_68626 & v_68849;
assign v_68855 = v_68624 & v_68854;
assign v_68857 = v_68769 & v_68856;
assign v_68858 = v_68623 & v_68854;
assign v_68860 = v_68772;
assign v_68862 = v_68774 & v_68861;
assign v_68863 = v_68862;
assign v_68865 = v_68864;
assign v_68866 = ~v_2363;
assign v_68867 = ~v_66663;
assign v_68868 = v_66663;
assign v_68869 = ~v_2367;
assign v_68870 = ~v_66667;
assign v_68871 = v_66667;
assign v_68872 = ~v_2371;
assign v_68873 = ~v_66671;
assign v_68874 = v_66671;
assign v_68875 = ~v_2375;
assign v_68876 = ~v_66675;
assign v_68877 = v_66675;
assign v_68878 = ~v_66678;
assign v_68879 = ~v_2380;
assign v_68880 = v_2380;
assign v_68881 = ~v_66682;
assign v_68882 = ~v_2384;
assign v_68883 = v_2384;
assign v_68884 = ~v_66686;
assign v_68885 = ~v_2388;
assign v_68886 = v_2388;
assign v_68887 = ~v_66690;
assign v_68888 = ~v_2392;
assign v_68889 = v_2392;
assign v_68890 = ~v_66694;
assign v_68891 = ~v_2396;
assign v_68892 = v_2396;
assign v_68893 = ~v_66698;
assign v_68894 = ~v_2400;
assign v_68895 = v_2400;
assign v_68896 = ~v_66702;
assign v_68897 = ~v_2404;
assign v_68898 = v_2404;
assign v_68899 = ~v_66706;
assign v_68900 = ~v_2408;
assign v_68901 = v_2408;
assign v_68902 = ~v_66710;
assign v_68903 = ~v_2412;
assign v_68904 = v_2412;
assign v_68905 = ~v_66714;
assign v_68906 = ~v_2416;
assign v_68907 = v_2416;
assign v_68908 = ~v_66718;
assign v_68909 = ~v_2420;
assign v_68910 = v_2420;
assign v_68911 = ~v_66722;
assign v_68912 = ~v_2424;
assign v_68913 = v_2424;
assign v_68914 = ~v_66726;
assign v_68915 = ~v_2428;
assign v_68916 = v_68915;
assign v_68918 = v_68917;
assign v_68920 = v_68912 & v_68919;
assign v_68922 = v_66722;
assign v_68924 = v_68921 & v_68923;
assign v_68926 = v_68909 & v_68925;
assign v_68928 = v_66718;
assign v_68930 = v_68927 & v_68929;
assign v_68932 = v_68906 & v_68931;
assign v_68934 = v_66714;
assign v_68936 = v_68933 & v_68935;
assign v_68938 = v_68903 & v_68937;
assign v_68940 = v_66710;
assign v_68942 = v_68939 & v_68941;
assign v_68944 = v_68900 & v_68943;
assign v_68946 = v_66706;
assign v_68948 = v_68945 & v_68947;
assign v_68950 = v_68897 & v_68949;
assign v_68952 = v_66702;
assign v_68954 = v_68951 & v_68953;
assign v_68956 = v_68894 & v_68955;
assign v_68958 = v_66698;
assign v_68960 = v_68957 & v_68959;
assign v_68962 = v_68891 & v_68961;
assign v_68964 = v_66694;
assign v_68966 = v_68963 & v_68965;
assign v_68968 = v_68888 & v_68967;
assign v_68970 = v_66690;
assign v_68972 = v_68969 & v_68971;
assign v_68974 = v_68885 & v_68973;
assign v_68976 = v_66686;
assign v_68978 = v_68975 & v_68977;
assign v_68980 = v_68882 & v_68979;
assign v_68982 = v_66682;
assign v_68984 = v_68981 & v_68983;
assign v_68986 = v_68879 & v_68985;
assign v_68988 = v_66678;
assign v_68990 = v_68987 & v_68989;
assign v_68992 = v_68876 & v_68991;
assign v_68994 = v_2375;
assign v_68996 = v_68993 & v_68995;
assign v_68998 = v_68873 & v_68997;
assign v_69000 = v_2371;
assign v_69002 = v_68999 & v_69001;
assign v_69004 = v_68870 & v_69003;
assign v_69006 = v_2367;
assign v_69008 = v_69005 & v_69007;
assign v_69010 = v_68867 & v_69009;
assign v_69012 = v_2363;
assign v_69014 = v_69011 & v_69013;
assign v_69016 = ~v_69015;
assign v_69018 = v_66726;
assign v_69019 = v_2428;
assign v_69020 = v_69019;
assign v_69021 = v_69018 & v_69020;
assign v_69022 = v_69021;
assign v_69023 = v_68912 & v_69022;
assign v_69025 = v_68922 & v_69024;
assign v_69026 = v_68911 & v_69022;
assign v_69028 = v_68909 & v_69027;
assign v_69030 = v_68928 & v_69029;
assign v_69031 = v_68908 & v_69027;
assign v_69033 = v_68906 & v_69032;
assign v_69035 = v_68934 & v_69034;
assign v_69036 = v_68905 & v_69032;
assign v_69038 = v_68903 & v_69037;
assign v_69040 = v_68940 & v_69039;
assign v_69041 = v_68902 & v_69037;
assign v_69043 = v_68900 & v_69042;
assign v_69045 = v_68946 & v_69044;
assign v_69046 = v_68899 & v_69042;
assign v_69048 = v_68897 & v_69047;
assign v_69050 = v_68952 & v_69049;
assign v_69051 = v_68896 & v_69047;
assign v_69053 = v_68894 & v_69052;
assign v_69055 = v_68958 & v_69054;
assign v_69056 = v_68893 & v_69052;
assign v_69058 = v_68891 & v_69057;
assign v_69060 = v_68964 & v_69059;
assign v_69061 = v_68890 & v_69057;
assign v_69063 = v_68888 & v_69062;
assign v_69065 = v_68970 & v_69064;
assign v_69066 = v_68887 & v_69062;
assign v_69068 = v_68885 & v_69067;
assign v_69070 = v_68976 & v_69069;
assign v_69071 = v_68884 & v_69067;
assign v_69073 = v_68882 & v_69072;
assign v_69075 = v_68982 & v_69074;
assign v_69076 = v_68881 & v_69072;
assign v_69078 = v_68879 & v_69077;
assign v_69080 = v_68988 & v_69079;
assign v_69081 = v_68878 & v_69077;
assign v_69083 = v_68876 & v_69082;
assign v_69085 = v_68994 & v_69084;
assign v_69086 = v_68875 & v_69082;
assign v_69088 = v_68873 & v_69087;
assign v_69090 = v_69000 & v_69089;
assign v_69091 = v_68872 & v_69087;
assign v_69093 = v_68870 & v_69092;
assign v_69095 = v_69006 & v_69094;
assign v_69096 = v_68869 & v_69092;
assign v_69098 = v_68867 & v_69097;
assign v_69100 = v_69012 & v_69099;
assign v_69101 = v_68866 & v_69097;
assign v_69103 = v_69015;
assign v_69105 = v_69017 & v_69104;
assign v_69106 = v_69105;
assign v_69108 = v_69107;
assign v_69109 = ~v_2623;
assign v_69110 = ~v_66663;
assign v_69111 = v_66663;
assign v_69112 = ~v_2627;
assign v_69113 = ~v_66667;
assign v_69114 = v_66667;
assign v_69115 = ~v_2631;
assign v_69116 = ~v_66671;
assign v_69117 = v_66671;
assign v_69118 = ~v_2635;
assign v_69119 = ~v_66675;
assign v_69120 = v_66675;
assign v_69121 = ~v_66678;
assign v_69122 = ~v_2640;
assign v_69123 = v_2640;
assign v_69124 = ~v_66682;
assign v_69125 = ~v_2644;
assign v_69126 = v_2644;
assign v_69127 = ~v_66686;
assign v_69128 = ~v_2648;
assign v_69129 = v_2648;
assign v_69130 = ~v_66690;
assign v_69131 = ~v_2652;
assign v_69132 = v_2652;
assign v_69133 = ~v_66694;
assign v_69134 = ~v_2656;
assign v_69135 = v_2656;
assign v_69136 = ~v_66698;
assign v_69137 = ~v_2660;
assign v_69138 = v_2660;
assign v_69139 = ~v_66702;
assign v_69140 = ~v_2664;
assign v_69141 = v_2664;
assign v_69142 = ~v_66706;
assign v_69143 = ~v_2668;
assign v_69144 = v_2668;
assign v_69145 = ~v_66710;
assign v_69146 = ~v_2672;
assign v_69147 = v_2672;
assign v_69148 = ~v_66714;
assign v_69149 = ~v_2676;
assign v_69150 = v_2676;
assign v_69151 = ~v_66718;
assign v_69152 = ~v_2680;
assign v_69153 = v_2680;
assign v_69154 = ~v_66722;
assign v_69155 = ~v_2684;
assign v_69156 = v_2684;
assign v_69157 = ~v_66726;
assign v_69158 = ~v_2688;
assign v_69159 = v_69158;
assign v_69161 = v_69160;
assign v_69163 = v_69155 & v_69162;
assign v_69165 = v_66722;
assign v_69167 = v_69164 & v_69166;
assign v_69169 = v_69152 & v_69168;
assign v_69171 = v_66718;
assign v_69173 = v_69170 & v_69172;
assign v_69175 = v_69149 & v_69174;
assign v_69177 = v_66714;
assign v_69179 = v_69176 & v_69178;
assign v_69181 = v_69146 & v_69180;
assign v_69183 = v_66710;
assign v_69185 = v_69182 & v_69184;
assign v_69187 = v_69143 & v_69186;
assign v_69189 = v_66706;
assign v_69191 = v_69188 & v_69190;
assign v_69193 = v_69140 & v_69192;
assign v_69195 = v_66702;
assign v_69197 = v_69194 & v_69196;
assign v_69199 = v_69137 & v_69198;
assign v_69201 = v_66698;
assign v_69203 = v_69200 & v_69202;
assign v_69205 = v_69134 & v_69204;
assign v_69207 = v_66694;
assign v_69209 = v_69206 & v_69208;
assign v_69211 = v_69131 & v_69210;
assign v_69213 = v_66690;
assign v_69215 = v_69212 & v_69214;
assign v_69217 = v_69128 & v_69216;
assign v_69219 = v_66686;
assign v_69221 = v_69218 & v_69220;
assign v_69223 = v_69125 & v_69222;
assign v_69225 = v_66682;
assign v_69227 = v_69224 & v_69226;
assign v_69229 = v_69122 & v_69228;
assign v_69231 = v_66678;
assign v_69233 = v_69230 & v_69232;
assign v_69235 = v_69119 & v_69234;
assign v_69237 = v_2635;
assign v_69239 = v_69236 & v_69238;
assign v_69241 = v_69116 & v_69240;
assign v_69243 = v_2631;
assign v_69245 = v_69242 & v_69244;
assign v_69247 = v_69113 & v_69246;
assign v_69249 = v_2627;
assign v_69251 = v_69248 & v_69250;
assign v_69253 = v_69110 & v_69252;
assign v_69255 = v_2623;
assign v_69257 = v_69254 & v_69256;
assign v_69259 = ~v_69258;
assign v_69261 = v_66726;
assign v_69262 = v_2688;
assign v_69263 = v_69262;
assign v_69264 = v_69261 & v_69263;
assign v_69265 = v_69264;
assign v_69266 = v_69155 & v_69265;
assign v_69268 = v_69165 & v_69267;
assign v_69269 = v_69154 & v_69265;
assign v_69271 = v_69152 & v_69270;
assign v_69273 = v_69171 & v_69272;
assign v_69274 = v_69151 & v_69270;
assign v_69276 = v_69149 & v_69275;
assign v_69278 = v_69177 & v_69277;
assign v_69279 = v_69148 & v_69275;
assign v_69281 = v_69146 & v_69280;
assign v_69283 = v_69183 & v_69282;
assign v_69284 = v_69145 & v_69280;
assign v_69286 = v_69143 & v_69285;
assign v_69288 = v_69189 & v_69287;
assign v_69289 = v_69142 & v_69285;
assign v_69291 = v_69140 & v_69290;
assign v_69293 = v_69195 & v_69292;
assign v_69294 = v_69139 & v_69290;
assign v_69296 = v_69137 & v_69295;
assign v_69298 = v_69201 & v_69297;
assign v_69299 = v_69136 & v_69295;
assign v_69301 = v_69134 & v_69300;
assign v_69303 = v_69207 & v_69302;
assign v_69304 = v_69133 & v_69300;
assign v_69306 = v_69131 & v_69305;
assign v_69308 = v_69213 & v_69307;
assign v_69309 = v_69130 & v_69305;
assign v_69311 = v_69128 & v_69310;
assign v_69313 = v_69219 & v_69312;
assign v_69314 = v_69127 & v_69310;
assign v_69316 = v_69125 & v_69315;
assign v_69318 = v_69225 & v_69317;
assign v_69319 = v_69124 & v_69315;
assign v_69321 = v_69122 & v_69320;
assign v_69323 = v_69231 & v_69322;
assign v_69324 = v_69121 & v_69320;
assign v_69326 = v_69119 & v_69325;
assign v_69328 = v_69237 & v_69327;
assign v_69329 = v_69118 & v_69325;
assign v_69331 = v_69116 & v_69330;
assign v_69333 = v_69243 & v_69332;
assign v_69334 = v_69115 & v_69330;
assign v_69336 = v_69113 & v_69335;
assign v_69338 = v_69249 & v_69337;
assign v_69339 = v_69112 & v_69335;
assign v_69341 = v_69110 & v_69340;
assign v_69343 = v_69255 & v_69342;
assign v_69344 = v_69109 & v_69340;
assign v_69346 = v_69258;
assign v_69348 = v_69260 & v_69347;
assign v_69349 = v_69348;
assign v_69351 = v_69350;
assign v_69352 = ~v_2883;
assign v_69353 = ~v_66663;
assign v_69354 = v_66663;
assign v_69355 = ~v_2887;
assign v_69356 = ~v_66667;
assign v_69357 = v_66667;
assign v_69358 = ~v_2891;
assign v_69359 = ~v_66671;
assign v_69360 = v_66671;
assign v_69361 = ~v_2895;
assign v_69362 = ~v_66675;
assign v_69363 = v_66675;
assign v_69364 = ~v_66678;
assign v_69365 = ~v_2900;
assign v_69366 = v_2900;
assign v_69367 = ~v_66682;
assign v_69368 = ~v_2904;
assign v_69369 = v_2904;
assign v_69370 = ~v_66686;
assign v_69371 = ~v_2908;
assign v_69372 = v_2908;
assign v_69373 = ~v_66690;
assign v_69374 = ~v_2912;
assign v_69375 = v_2912;
assign v_69376 = ~v_66694;
assign v_69377 = ~v_2916;
assign v_69378 = v_2916;
assign v_69379 = ~v_66698;
assign v_69380 = ~v_2920;
assign v_69381 = v_2920;
assign v_69382 = ~v_66702;
assign v_69383 = ~v_2924;
assign v_69384 = v_2924;
assign v_69385 = ~v_66706;
assign v_69386 = ~v_2928;
assign v_69387 = v_2928;
assign v_69388 = ~v_66710;
assign v_69389 = ~v_2932;
assign v_69390 = v_2932;
assign v_69391 = ~v_66714;
assign v_69392 = ~v_2936;
assign v_69393 = v_2936;
assign v_69394 = ~v_66718;
assign v_69395 = ~v_2940;
assign v_69396 = v_2940;
assign v_69397 = ~v_66722;
assign v_69398 = ~v_2944;
assign v_69399 = v_2944;
assign v_69400 = ~v_66726;
assign v_69401 = ~v_2948;
assign v_69402 = v_69401;
assign v_69404 = v_69403;
assign v_69406 = v_69398 & v_69405;
assign v_69408 = v_66722;
assign v_69410 = v_69407 & v_69409;
assign v_69412 = v_69395 & v_69411;
assign v_69414 = v_66718;
assign v_69416 = v_69413 & v_69415;
assign v_69418 = v_69392 & v_69417;
assign v_69420 = v_66714;
assign v_69422 = v_69419 & v_69421;
assign v_69424 = v_69389 & v_69423;
assign v_69426 = v_66710;
assign v_69428 = v_69425 & v_69427;
assign v_69430 = v_69386 & v_69429;
assign v_69432 = v_66706;
assign v_69434 = v_69431 & v_69433;
assign v_69436 = v_69383 & v_69435;
assign v_69438 = v_66702;
assign v_69440 = v_69437 & v_69439;
assign v_69442 = v_69380 & v_69441;
assign v_69444 = v_66698;
assign v_69446 = v_69443 & v_69445;
assign v_69448 = v_69377 & v_69447;
assign v_69450 = v_66694;
assign v_69452 = v_69449 & v_69451;
assign v_69454 = v_69374 & v_69453;
assign v_69456 = v_66690;
assign v_69458 = v_69455 & v_69457;
assign v_69460 = v_69371 & v_69459;
assign v_69462 = v_66686;
assign v_69464 = v_69461 & v_69463;
assign v_69466 = v_69368 & v_69465;
assign v_69468 = v_66682;
assign v_69470 = v_69467 & v_69469;
assign v_69472 = v_69365 & v_69471;
assign v_69474 = v_66678;
assign v_69476 = v_69473 & v_69475;
assign v_69478 = v_69362 & v_69477;
assign v_69480 = v_2895;
assign v_69482 = v_69479 & v_69481;
assign v_69484 = v_69359 & v_69483;
assign v_69486 = v_2891;
assign v_69488 = v_69485 & v_69487;
assign v_69490 = v_69356 & v_69489;
assign v_69492 = v_2887;
assign v_69494 = v_69491 & v_69493;
assign v_69496 = v_69353 & v_69495;
assign v_69498 = v_2883;
assign v_69500 = v_69497 & v_69499;
assign v_69502 = ~v_69501;
assign v_69504 = v_66726;
assign v_69505 = v_2948;
assign v_69506 = v_69505;
assign v_69507 = v_69504 & v_69506;
assign v_69508 = v_69507;
assign v_69509 = v_69398 & v_69508;
assign v_69511 = v_69408 & v_69510;
assign v_69512 = v_69397 & v_69508;
assign v_69514 = v_69395 & v_69513;
assign v_69516 = v_69414 & v_69515;
assign v_69517 = v_69394 & v_69513;
assign v_69519 = v_69392 & v_69518;
assign v_69521 = v_69420 & v_69520;
assign v_69522 = v_69391 & v_69518;
assign v_69524 = v_69389 & v_69523;
assign v_69526 = v_69426 & v_69525;
assign v_69527 = v_69388 & v_69523;
assign v_69529 = v_69386 & v_69528;
assign v_69531 = v_69432 & v_69530;
assign v_69532 = v_69385 & v_69528;
assign v_69534 = v_69383 & v_69533;
assign v_69536 = v_69438 & v_69535;
assign v_69537 = v_69382 & v_69533;
assign v_69539 = v_69380 & v_69538;
assign v_69541 = v_69444 & v_69540;
assign v_69542 = v_69379 & v_69538;
assign v_69544 = v_69377 & v_69543;
assign v_69546 = v_69450 & v_69545;
assign v_69547 = v_69376 & v_69543;
assign v_69549 = v_69374 & v_69548;
assign v_69551 = v_69456 & v_69550;
assign v_69552 = v_69373 & v_69548;
assign v_69554 = v_69371 & v_69553;
assign v_69556 = v_69462 & v_69555;
assign v_69557 = v_69370 & v_69553;
assign v_69559 = v_69368 & v_69558;
assign v_69561 = v_69468 & v_69560;
assign v_69562 = v_69367 & v_69558;
assign v_69564 = v_69365 & v_69563;
assign v_69566 = v_69474 & v_69565;
assign v_69567 = v_69364 & v_69563;
assign v_69569 = v_69362 & v_69568;
assign v_69571 = v_69480 & v_69570;
assign v_69572 = v_69361 & v_69568;
assign v_69574 = v_69359 & v_69573;
assign v_69576 = v_69486 & v_69575;
assign v_69577 = v_69358 & v_69573;
assign v_69579 = v_69356 & v_69578;
assign v_69581 = v_69492 & v_69580;
assign v_69582 = v_69355 & v_69578;
assign v_69584 = v_69353 & v_69583;
assign v_69586 = v_69498 & v_69585;
assign v_69587 = v_69352 & v_69583;
assign v_69589 = v_69501;
assign v_69591 = v_69503 & v_69590;
assign v_69592 = v_69591;
assign v_69594 = v_69593;
assign v_69595 = ~v_3143;
assign v_69596 = ~v_66663;
assign v_69597 = v_66663;
assign v_69598 = ~v_3147;
assign v_69599 = ~v_66667;
assign v_69600 = v_66667;
assign v_69601 = ~v_3151;
assign v_69602 = ~v_66671;
assign v_69603 = v_66671;
assign v_69604 = ~v_3155;
assign v_69605 = ~v_66675;
assign v_69606 = v_66675;
assign v_69607 = ~v_66678;
assign v_69608 = ~v_3160;
assign v_69609 = v_3160;
assign v_69610 = ~v_66682;
assign v_69611 = ~v_3164;
assign v_69612 = v_3164;
assign v_69613 = ~v_66686;
assign v_69614 = ~v_3168;
assign v_69615 = v_3168;
assign v_69616 = ~v_66690;
assign v_69617 = ~v_3172;
assign v_69618 = v_3172;
assign v_69619 = ~v_66694;
assign v_69620 = ~v_3176;
assign v_69621 = v_3176;
assign v_69622 = ~v_66698;
assign v_69623 = ~v_3180;
assign v_69624 = v_3180;
assign v_69625 = ~v_66702;
assign v_69626 = ~v_3184;
assign v_69627 = v_3184;
assign v_69628 = ~v_66706;
assign v_69629 = ~v_3188;
assign v_69630 = v_3188;
assign v_69631 = ~v_66710;
assign v_69632 = ~v_3192;
assign v_69633 = v_3192;
assign v_69634 = ~v_66714;
assign v_69635 = ~v_3196;
assign v_69636 = v_3196;
assign v_69637 = ~v_66718;
assign v_69638 = ~v_3200;
assign v_69639 = v_3200;
assign v_69640 = ~v_66722;
assign v_69641 = ~v_3204;
assign v_69642 = v_3204;
assign v_69643 = ~v_66726;
assign v_69644 = ~v_3208;
assign v_69645 = v_69644;
assign v_69647 = v_69646;
assign v_69649 = v_69641 & v_69648;
assign v_69651 = v_66722;
assign v_69653 = v_69650 & v_69652;
assign v_69655 = v_69638 & v_69654;
assign v_69657 = v_66718;
assign v_69659 = v_69656 & v_69658;
assign v_69661 = v_69635 & v_69660;
assign v_69663 = v_66714;
assign v_69665 = v_69662 & v_69664;
assign v_69667 = v_69632 & v_69666;
assign v_69669 = v_66710;
assign v_69671 = v_69668 & v_69670;
assign v_69673 = v_69629 & v_69672;
assign v_69675 = v_66706;
assign v_69677 = v_69674 & v_69676;
assign v_69679 = v_69626 & v_69678;
assign v_69681 = v_66702;
assign v_69683 = v_69680 & v_69682;
assign v_69685 = v_69623 & v_69684;
assign v_69687 = v_66698;
assign v_69689 = v_69686 & v_69688;
assign v_69691 = v_69620 & v_69690;
assign v_69693 = v_66694;
assign v_69695 = v_69692 & v_69694;
assign v_69697 = v_69617 & v_69696;
assign v_69699 = v_66690;
assign v_69701 = v_69698 & v_69700;
assign v_69703 = v_69614 & v_69702;
assign v_69705 = v_66686;
assign v_69707 = v_69704 & v_69706;
assign v_69709 = v_69611 & v_69708;
assign v_69711 = v_66682;
assign v_69713 = v_69710 & v_69712;
assign v_69715 = v_69608 & v_69714;
assign v_69717 = v_66678;
assign v_69719 = v_69716 & v_69718;
assign v_69721 = v_69605 & v_69720;
assign v_69723 = v_3155;
assign v_69725 = v_69722 & v_69724;
assign v_69727 = v_69602 & v_69726;
assign v_69729 = v_3151;
assign v_69731 = v_69728 & v_69730;
assign v_69733 = v_69599 & v_69732;
assign v_69735 = v_3147;
assign v_69737 = v_69734 & v_69736;
assign v_69739 = v_69596 & v_69738;
assign v_69741 = v_3143;
assign v_69743 = v_69740 & v_69742;
assign v_69745 = ~v_69744;
assign v_69747 = v_66726;
assign v_69748 = v_3208;
assign v_69749 = v_69748;
assign v_69750 = v_69747 & v_69749;
assign v_69751 = v_69750;
assign v_69752 = v_69641 & v_69751;
assign v_69754 = v_69651 & v_69753;
assign v_69755 = v_69640 & v_69751;
assign v_69757 = v_69638 & v_69756;
assign v_69759 = v_69657 & v_69758;
assign v_69760 = v_69637 & v_69756;
assign v_69762 = v_69635 & v_69761;
assign v_69764 = v_69663 & v_69763;
assign v_69765 = v_69634 & v_69761;
assign v_69767 = v_69632 & v_69766;
assign v_69769 = v_69669 & v_69768;
assign v_69770 = v_69631 & v_69766;
assign v_69772 = v_69629 & v_69771;
assign v_69774 = v_69675 & v_69773;
assign v_69775 = v_69628 & v_69771;
assign v_69777 = v_69626 & v_69776;
assign v_69779 = v_69681 & v_69778;
assign v_69780 = v_69625 & v_69776;
assign v_69782 = v_69623 & v_69781;
assign v_69784 = v_69687 & v_69783;
assign v_69785 = v_69622 & v_69781;
assign v_69787 = v_69620 & v_69786;
assign v_69789 = v_69693 & v_69788;
assign v_69790 = v_69619 & v_69786;
assign v_69792 = v_69617 & v_69791;
assign v_69794 = v_69699 & v_69793;
assign v_69795 = v_69616 & v_69791;
assign v_69797 = v_69614 & v_69796;
assign v_69799 = v_69705 & v_69798;
assign v_69800 = v_69613 & v_69796;
assign v_69802 = v_69611 & v_69801;
assign v_69804 = v_69711 & v_69803;
assign v_69805 = v_69610 & v_69801;
assign v_69807 = v_69608 & v_69806;
assign v_69809 = v_69717 & v_69808;
assign v_69810 = v_69607 & v_69806;
assign v_69812 = v_69605 & v_69811;
assign v_69814 = v_69723 & v_69813;
assign v_69815 = v_69604 & v_69811;
assign v_69817 = v_69602 & v_69816;
assign v_69819 = v_69729 & v_69818;
assign v_69820 = v_69601 & v_69816;
assign v_69822 = v_69599 & v_69821;
assign v_69824 = v_69735 & v_69823;
assign v_69825 = v_69598 & v_69821;
assign v_69827 = v_69596 & v_69826;
assign v_69829 = v_69741 & v_69828;
assign v_69830 = v_69595 & v_69826;
assign v_69832 = v_69744;
assign v_69834 = v_69746 & v_69833;
assign v_69835 = v_69834;
assign v_69837 = v_69836;
assign v_69838 = ~v_3403;
assign v_69839 = ~v_66663;
assign v_69840 = v_66663;
assign v_69841 = ~v_3407;
assign v_69842 = ~v_66667;
assign v_69843 = v_66667;
assign v_69844 = ~v_3411;
assign v_69845 = ~v_66671;
assign v_69846 = v_66671;
assign v_69847 = ~v_3415;
assign v_69848 = ~v_66675;
assign v_69849 = v_66675;
assign v_69850 = ~v_66678;
assign v_69851 = ~v_3420;
assign v_69852 = v_3420;
assign v_69853 = ~v_66682;
assign v_69854 = ~v_3424;
assign v_69855 = v_3424;
assign v_69856 = ~v_66686;
assign v_69857 = ~v_3428;
assign v_69858 = v_3428;
assign v_69859 = ~v_66690;
assign v_69860 = ~v_3432;
assign v_69861 = v_3432;
assign v_69862 = ~v_66694;
assign v_69863 = ~v_3436;
assign v_69864 = v_3436;
assign v_69865 = ~v_66698;
assign v_69866 = ~v_3440;
assign v_69867 = v_3440;
assign v_69868 = ~v_66702;
assign v_69869 = ~v_3444;
assign v_69870 = v_3444;
assign v_69871 = ~v_66706;
assign v_69872 = ~v_3448;
assign v_69873 = v_3448;
assign v_69874 = ~v_66710;
assign v_69875 = ~v_3452;
assign v_69876 = v_3452;
assign v_69877 = ~v_66714;
assign v_69878 = ~v_3456;
assign v_69879 = v_3456;
assign v_69880 = ~v_66718;
assign v_69881 = ~v_3460;
assign v_69882 = v_3460;
assign v_69883 = ~v_66722;
assign v_69884 = ~v_3464;
assign v_69885 = v_3464;
assign v_69886 = ~v_66726;
assign v_69887 = ~v_3468;
assign v_69888 = v_69887;
assign v_69890 = v_69889;
assign v_69892 = v_69884 & v_69891;
assign v_69894 = v_66722;
assign v_69896 = v_69893 & v_69895;
assign v_69898 = v_69881 & v_69897;
assign v_69900 = v_66718;
assign v_69902 = v_69899 & v_69901;
assign v_69904 = v_69878 & v_69903;
assign v_69906 = v_66714;
assign v_69908 = v_69905 & v_69907;
assign v_69910 = v_69875 & v_69909;
assign v_69912 = v_66710;
assign v_69914 = v_69911 & v_69913;
assign v_69916 = v_69872 & v_69915;
assign v_69918 = v_66706;
assign v_69920 = v_69917 & v_69919;
assign v_69922 = v_69869 & v_69921;
assign v_69924 = v_66702;
assign v_69926 = v_69923 & v_69925;
assign v_69928 = v_69866 & v_69927;
assign v_69930 = v_66698;
assign v_69932 = v_69929 & v_69931;
assign v_69934 = v_69863 & v_69933;
assign v_69936 = v_66694;
assign v_69938 = v_69935 & v_69937;
assign v_69940 = v_69860 & v_69939;
assign v_69942 = v_66690;
assign v_69944 = v_69941 & v_69943;
assign v_69946 = v_69857 & v_69945;
assign v_69948 = v_66686;
assign v_69950 = v_69947 & v_69949;
assign v_69952 = v_69854 & v_69951;
assign v_69954 = v_66682;
assign v_69956 = v_69953 & v_69955;
assign v_69958 = v_69851 & v_69957;
assign v_69960 = v_66678;
assign v_69962 = v_69959 & v_69961;
assign v_69964 = v_69848 & v_69963;
assign v_69966 = v_3415;
assign v_69968 = v_69965 & v_69967;
assign v_69970 = v_69845 & v_69969;
assign v_69972 = v_3411;
assign v_69974 = v_69971 & v_69973;
assign v_69976 = v_69842 & v_69975;
assign v_69978 = v_3407;
assign v_69980 = v_69977 & v_69979;
assign v_69982 = v_69839 & v_69981;
assign v_69984 = v_3403;
assign v_69986 = v_69983 & v_69985;
assign v_69988 = ~v_69987;
assign v_69990 = v_66726;
assign v_69991 = v_3468;
assign v_69992 = v_69991;
assign v_69993 = v_69990 & v_69992;
assign v_69994 = v_69993;
assign v_69995 = v_69884 & v_69994;
assign v_69997 = v_69894 & v_69996;
assign v_69998 = v_69883 & v_69994;
assign v_70000 = v_69881 & v_69999;
assign v_70002 = v_69900 & v_70001;
assign v_70003 = v_69880 & v_69999;
assign v_70005 = v_69878 & v_70004;
assign v_70007 = v_69906 & v_70006;
assign v_70008 = v_69877 & v_70004;
assign v_70010 = v_69875 & v_70009;
assign v_70012 = v_69912 & v_70011;
assign v_70013 = v_69874 & v_70009;
assign v_70015 = v_69872 & v_70014;
assign v_70017 = v_69918 & v_70016;
assign v_70018 = v_69871 & v_70014;
assign v_70020 = v_69869 & v_70019;
assign v_70022 = v_69924 & v_70021;
assign v_70023 = v_69868 & v_70019;
assign v_70025 = v_69866 & v_70024;
assign v_70027 = v_69930 & v_70026;
assign v_70028 = v_69865 & v_70024;
assign v_70030 = v_69863 & v_70029;
assign v_70032 = v_69936 & v_70031;
assign v_70033 = v_69862 & v_70029;
assign v_70035 = v_69860 & v_70034;
assign v_70037 = v_69942 & v_70036;
assign v_70038 = v_69859 & v_70034;
assign v_70040 = v_69857 & v_70039;
assign v_70042 = v_69948 & v_70041;
assign v_70043 = v_69856 & v_70039;
assign v_70045 = v_69854 & v_70044;
assign v_70047 = v_69954 & v_70046;
assign v_70048 = v_69853 & v_70044;
assign v_70050 = v_69851 & v_70049;
assign v_70052 = v_69960 & v_70051;
assign v_70053 = v_69850 & v_70049;
assign v_70055 = v_69848 & v_70054;
assign v_70057 = v_69966 & v_70056;
assign v_70058 = v_69847 & v_70054;
assign v_70060 = v_69845 & v_70059;
assign v_70062 = v_69972 & v_70061;
assign v_70063 = v_69844 & v_70059;
assign v_70065 = v_69842 & v_70064;
assign v_70067 = v_69978 & v_70066;
assign v_70068 = v_69841 & v_70064;
assign v_70070 = v_69839 & v_70069;
assign v_70072 = v_69984 & v_70071;
assign v_70073 = v_69838 & v_70069;
assign v_70075 = v_69987;
assign v_70077 = v_69989 & v_70076;
assign v_70078 = v_70077;
assign v_70080 = v_70079;
assign v_70081 = ~v_3663;
assign v_70082 = ~v_66663;
assign v_70083 = v_66663;
assign v_70084 = ~v_3667;
assign v_70085 = ~v_66667;
assign v_70086 = v_66667;
assign v_70087 = ~v_3671;
assign v_70088 = ~v_66671;
assign v_70089 = v_66671;
assign v_70090 = ~v_3675;
assign v_70091 = ~v_66675;
assign v_70092 = v_66675;
assign v_70093 = ~v_66678;
assign v_70094 = ~v_3680;
assign v_70095 = v_3680;
assign v_70096 = ~v_66682;
assign v_70097 = ~v_3684;
assign v_70098 = v_3684;
assign v_70099 = ~v_66686;
assign v_70100 = ~v_3688;
assign v_70101 = v_3688;
assign v_70102 = ~v_66690;
assign v_70103 = ~v_3692;
assign v_70104 = v_3692;
assign v_70105 = ~v_66694;
assign v_70106 = ~v_3696;
assign v_70107 = v_3696;
assign v_70108 = ~v_66698;
assign v_70109 = ~v_3700;
assign v_70110 = v_3700;
assign v_70111 = ~v_66702;
assign v_70112 = ~v_3704;
assign v_70113 = v_3704;
assign v_70114 = ~v_66706;
assign v_70115 = ~v_3708;
assign v_70116 = v_3708;
assign v_70117 = ~v_66710;
assign v_70118 = ~v_3712;
assign v_70119 = v_3712;
assign v_70120 = ~v_66714;
assign v_70121 = ~v_3716;
assign v_70122 = v_3716;
assign v_70123 = ~v_66718;
assign v_70124 = ~v_3720;
assign v_70125 = v_3720;
assign v_70126 = ~v_66722;
assign v_70127 = ~v_3724;
assign v_70128 = v_3724;
assign v_70129 = ~v_66726;
assign v_70130 = ~v_3728;
assign v_70131 = v_70130;
assign v_70133 = v_70132;
assign v_70135 = v_70127 & v_70134;
assign v_70137 = v_66722;
assign v_70139 = v_70136 & v_70138;
assign v_70141 = v_70124 & v_70140;
assign v_70143 = v_66718;
assign v_70145 = v_70142 & v_70144;
assign v_70147 = v_70121 & v_70146;
assign v_70149 = v_66714;
assign v_70151 = v_70148 & v_70150;
assign v_70153 = v_70118 & v_70152;
assign v_70155 = v_66710;
assign v_70157 = v_70154 & v_70156;
assign v_70159 = v_70115 & v_70158;
assign v_70161 = v_66706;
assign v_70163 = v_70160 & v_70162;
assign v_70165 = v_70112 & v_70164;
assign v_70167 = v_66702;
assign v_70169 = v_70166 & v_70168;
assign v_70171 = v_70109 & v_70170;
assign v_70173 = v_66698;
assign v_70175 = v_70172 & v_70174;
assign v_70177 = v_70106 & v_70176;
assign v_70179 = v_66694;
assign v_70181 = v_70178 & v_70180;
assign v_70183 = v_70103 & v_70182;
assign v_70185 = v_66690;
assign v_70187 = v_70184 & v_70186;
assign v_70189 = v_70100 & v_70188;
assign v_70191 = v_66686;
assign v_70193 = v_70190 & v_70192;
assign v_70195 = v_70097 & v_70194;
assign v_70197 = v_66682;
assign v_70199 = v_70196 & v_70198;
assign v_70201 = v_70094 & v_70200;
assign v_70203 = v_66678;
assign v_70205 = v_70202 & v_70204;
assign v_70207 = v_70091 & v_70206;
assign v_70209 = v_3675;
assign v_70211 = v_70208 & v_70210;
assign v_70213 = v_70088 & v_70212;
assign v_70215 = v_3671;
assign v_70217 = v_70214 & v_70216;
assign v_70219 = v_70085 & v_70218;
assign v_70221 = v_3667;
assign v_70223 = v_70220 & v_70222;
assign v_70225 = v_70082 & v_70224;
assign v_70227 = v_3663;
assign v_70229 = v_70226 & v_70228;
assign v_70231 = ~v_70230;
assign v_70233 = v_66726;
assign v_70234 = v_3728;
assign v_70235 = v_70234;
assign v_70236 = v_70233 & v_70235;
assign v_70237 = v_70236;
assign v_70238 = v_70127 & v_70237;
assign v_70240 = v_70137 & v_70239;
assign v_70241 = v_70126 & v_70237;
assign v_70243 = v_70124 & v_70242;
assign v_70245 = v_70143 & v_70244;
assign v_70246 = v_70123 & v_70242;
assign v_70248 = v_70121 & v_70247;
assign v_70250 = v_70149 & v_70249;
assign v_70251 = v_70120 & v_70247;
assign v_70253 = v_70118 & v_70252;
assign v_70255 = v_70155 & v_70254;
assign v_70256 = v_70117 & v_70252;
assign v_70258 = v_70115 & v_70257;
assign v_70260 = v_70161 & v_70259;
assign v_70261 = v_70114 & v_70257;
assign v_70263 = v_70112 & v_70262;
assign v_70265 = v_70167 & v_70264;
assign v_70266 = v_70111 & v_70262;
assign v_70268 = v_70109 & v_70267;
assign v_70270 = v_70173 & v_70269;
assign v_70271 = v_70108 & v_70267;
assign v_70273 = v_70106 & v_70272;
assign v_70275 = v_70179 & v_70274;
assign v_70276 = v_70105 & v_70272;
assign v_70278 = v_70103 & v_70277;
assign v_70280 = v_70185 & v_70279;
assign v_70281 = v_70102 & v_70277;
assign v_70283 = v_70100 & v_70282;
assign v_70285 = v_70191 & v_70284;
assign v_70286 = v_70099 & v_70282;
assign v_70288 = v_70097 & v_70287;
assign v_70290 = v_70197 & v_70289;
assign v_70291 = v_70096 & v_70287;
assign v_70293 = v_70094 & v_70292;
assign v_70295 = v_70203 & v_70294;
assign v_70296 = v_70093 & v_70292;
assign v_70298 = v_70091 & v_70297;
assign v_70300 = v_70209 & v_70299;
assign v_70301 = v_70090 & v_70297;
assign v_70303 = v_70088 & v_70302;
assign v_70305 = v_70215 & v_70304;
assign v_70306 = v_70087 & v_70302;
assign v_70308 = v_70085 & v_70307;
assign v_70310 = v_70221 & v_70309;
assign v_70311 = v_70084 & v_70307;
assign v_70313 = v_70082 & v_70312;
assign v_70315 = v_70227 & v_70314;
assign v_70316 = v_70081 & v_70312;
assign v_70318 = v_70230;
assign v_70320 = v_70232 & v_70319;
assign v_70321 = v_70320;
assign v_70323 = v_70322;
assign v_70324 = ~v_3923;
assign v_70325 = ~v_66663;
assign v_70326 = v_66663;
assign v_70327 = ~v_3927;
assign v_70328 = ~v_66667;
assign v_70329 = v_66667;
assign v_70330 = ~v_3931;
assign v_70331 = ~v_66671;
assign v_70332 = v_66671;
assign v_70333 = ~v_3935;
assign v_70334 = ~v_66675;
assign v_70335 = v_66675;
assign v_70336 = ~v_66678;
assign v_70337 = ~v_3940;
assign v_70338 = v_3940;
assign v_70339 = ~v_66682;
assign v_70340 = ~v_3944;
assign v_70341 = v_3944;
assign v_70342 = ~v_66686;
assign v_70343 = ~v_3948;
assign v_70344 = v_3948;
assign v_70345 = ~v_66690;
assign v_70346 = ~v_3952;
assign v_70347 = v_3952;
assign v_70348 = ~v_66694;
assign v_70349 = ~v_3956;
assign v_70350 = v_3956;
assign v_70351 = ~v_66698;
assign v_70352 = ~v_3960;
assign v_70353 = v_3960;
assign v_70354 = ~v_66702;
assign v_70355 = ~v_3964;
assign v_70356 = v_3964;
assign v_70357 = ~v_66706;
assign v_70358 = ~v_3968;
assign v_70359 = v_3968;
assign v_70360 = ~v_66710;
assign v_70361 = ~v_3972;
assign v_70362 = v_3972;
assign v_70363 = ~v_66714;
assign v_70364 = ~v_3976;
assign v_70365 = v_3976;
assign v_70366 = ~v_66718;
assign v_70367 = ~v_3980;
assign v_70368 = v_3980;
assign v_70369 = ~v_66722;
assign v_70370 = ~v_3984;
assign v_70371 = v_3984;
assign v_70372 = ~v_66726;
assign v_70373 = ~v_3988;
assign v_70374 = v_70373;
assign v_70376 = v_70375;
assign v_70378 = v_70370 & v_70377;
assign v_70380 = v_66722;
assign v_70382 = v_70379 & v_70381;
assign v_70384 = v_70367 & v_70383;
assign v_70386 = v_66718;
assign v_70388 = v_70385 & v_70387;
assign v_70390 = v_70364 & v_70389;
assign v_70392 = v_66714;
assign v_70394 = v_70391 & v_70393;
assign v_70396 = v_70361 & v_70395;
assign v_70398 = v_66710;
assign v_70400 = v_70397 & v_70399;
assign v_70402 = v_70358 & v_70401;
assign v_70404 = v_66706;
assign v_70406 = v_70403 & v_70405;
assign v_70408 = v_70355 & v_70407;
assign v_70410 = v_66702;
assign v_70412 = v_70409 & v_70411;
assign v_70414 = v_70352 & v_70413;
assign v_70416 = v_66698;
assign v_70418 = v_70415 & v_70417;
assign v_70420 = v_70349 & v_70419;
assign v_70422 = v_66694;
assign v_70424 = v_70421 & v_70423;
assign v_70426 = v_70346 & v_70425;
assign v_70428 = v_66690;
assign v_70430 = v_70427 & v_70429;
assign v_70432 = v_70343 & v_70431;
assign v_70434 = v_66686;
assign v_70436 = v_70433 & v_70435;
assign v_70438 = v_70340 & v_70437;
assign v_70440 = v_66682;
assign v_70442 = v_70439 & v_70441;
assign v_70444 = v_70337 & v_70443;
assign v_70446 = v_66678;
assign v_70448 = v_70445 & v_70447;
assign v_70450 = v_70334 & v_70449;
assign v_70452 = v_3935;
assign v_70454 = v_70451 & v_70453;
assign v_70456 = v_70331 & v_70455;
assign v_70458 = v_3931;
assign v_70460 = v_70457 & v_70459;
assign v_70462 = v_70328 & v_70461;
assign v_70464 = v_3927;
assign v_70466 = v_70463 & v_70465;
assign v_70468 = v_70325 & v_70467;
assign v_70470 = v_3923;
assign v_70472 = v_70469 & v_70471;
assign v_70474 = ~v_70473;
assign v_70476 = v_66726;
assign v_70477 = v_3988;
assign v_70478 = v_70477;
assign v_70479 = v_70476 & v_70478;
assign v_70480 = v_70479;
assign v_70481 = v_70370 & v_70480;
assign v_70483 = v_70380 & v_70482;
assign v_70484 = v_70369 & v_70480;
assign v_70486 = v_70367 & v_70485;
assign v_70488 = v_70386 & v_70487;
assign v_70489 = v_70366 & v_70485;
assign v_70491 = v_70364 & v_70490;
assign v_70493 = v_70392 & v_70492;
assign v_70494 = v_70363 & v_70490;
assign v_70496 = v_70361 & v_70495;
assign v_70498 = v_70398 & v_70497;
assign v_70499 = v_70360 & v_70495;
assign v_70501 = v_70358 & v_70500;
assign v_70503 = v_70404 & v_70502;
assign v_70504 = v_70357 & v_70500;
assign v_70506 = v_70355 & v_70505;
assign v_70508 = v_70410 & v_70507;
assign v_70509 = v_70354 & v_70505;
assign v_70511 = v_70352 & v_70510;
assign v_70513 = v_70416 & v_70512;
assign v_70514 = v_70351 & v_70510;
assign v_70516 = v_70349 & v_70515;
assign v_70518 = v_70422 & v_70517;
assign v_70519 = v_70348 & v_70515;
assign v_70521 = v_70346 & v_70520;
assign v_70523 = v_70428 & v_70522;
assign v_70524 = v_70345 & v_70520;
assign v_70526 = v_70343 & v_70525;
assign v_70528 = v_70434 & v_70527;
assign v_70529 = v_70342 & v_70525;
assign v_70531 = v_70340 & v_70530;
assign v_70533 = v_70440 & v_70532;
assign v_70534 = v_70339 & v_70530;
assign v_70536 = v_70337 & v_70535;
assign v_70538 = v_70446 & v_70537;
assign v_70539 = v_70336 & v_70535;
assign v_70541 = v_70334 & v_70540;
assign v_70543 = v_70452 & v_70542;
assign v_70544 = v_70333 & v_70540;
assign v_70546 = v_70331 & v_70545;
assign v_70548 = v_70458 & v_70547;
assign v_70549 = v_70330 & v_70545;
assign v_70551 = v_70328 & v_70550;
assign v_70553 = v_70464 & v_70552;
assign v_70554 = v_70327 & v_70550;
assign v_70556 = v_70325 & v_70555;
assign v_70558 = v_70470 & v_70557;
assign v_70559 = v_70324 & v_70555;
assign v_70561 = v_70473;
assign v_70563 = v_70475 & v_70562;
assign v_70564 = v_70563;
assign v_70566 = v_70565;
assign v_70567 = ~v_4182;
assign v_70568 = ~v_66663;
assign v_70569 = v_66663;
assign v_70570 = ~v_4186;
assign v_70571 = ~v_66667;
assign v_70572 = v_66667;
assign v_70573 = ~v_4190;
assign v_70574 = ~v_66671;
assign v_70575 = v_66671;
assign v_70576 = ~v_4194;
assign v_70577 = ~v_66675;
assign v_70578 = v_66675;
assign v_70579 = ~v_66678;
assign v_70580 = ~v_4199;
assign v_70581 = v_4199;
assign v_70582 = ~v_66682;
assign v_70583 = ~v_4203;
assign v_70584 = v_4203;
assign v_70585 = ~v_66686;
assign v_70586 = ~v_4207;
assign v_70587 = v_4207;
assign v_70588 = ~v_66690;
assign v_70589 = ~v_4211;
assign v_70590 = v_4211;
assign v_70591 = ~v_66694;
assign v_70592 = ~v_4215;
assign v_70593 = v_4215;
assign v_70594 = ~v_66698;
assign v_70595 = ~v_4219;
assign v_70596 = v_4219;
assign v_70597 = ~v_66702;
assign v_70598 = ~v_4223;
assign v_70599 = v_4223;
assign v_70600 = ~v_66706;
assign v_70601 = ~v_4227;
assign v_70602 = v_4227;
assign v_70603 = ~v_66710;
assign v_70604 = ~v_4231;
assign v_70605 = v_4231;
assign v_70606 = ~v_66714;
assign v_70607 = ~v_4235;
assign v_70608 = v_4235;
assign v_70609 = ~v_66718;
assign v_70610 = ~v_4239;
assign v_70611 = v_4239;
assign v_70612 = ~v_66722;
assign v_70613 = ~v_4243;
assign v_70614 = v_4243;
assign v_70615 = ~v_66726;
assign v_70616 = ~v_4247;
assign v_70617 = v_70616;
assign v_70619 = v_70618;
assign v_70621 = v_70613 & v_70620;
assign v_70623 = v_66722;
assign v_70625 = v_70622 & v_70624;
assign v_70627 = v_70610 & v_70626;
assign v_70629 = v_66718;
assign v_70631 = v_70628 & v_70630;
assign v_70633 = v_70607 & v_70632;
assign v_70635 = v_66714;
assign v_70637 = v_70634 & v_70636;
assign v_70639 = v_70604 & v_70638;
assign v_70641 = v_66710;
assign v_70643 = v_70640 & v_70642;
assign v_70645 = v_70601 & v_70644;
assign v_70647 = v_66706;
assign v_70649 = v_70646 & v_70648;
assign v_70651 = v_70598 & v_70650;
assign v_70653 = v_66702;
assign v_70655 = v_70652 & v_70654;
assign v_70657 = v_70595 & v_70656;
assign v_70659 = v_66698;
assign v_70661 = v_70658 & v_70660;
assign v_70663 = v_70592 & v_70662;
assign v_70665 = v_66694;
assign v_70667 = v_70664 & v_70666;
assign v_70669 = v_70589 & v_70668;
assign v_70671 = v_66690;
assign v_70673 = v_70670 & v_70672;
assign v_70675 = v_70586 & v_70674;
assign v_70677 = v_66686;
assign v_70679 = v_70676 & v_70678;
assign v_70681 = v_70583 & v_70680;
assign v_70683 = v_66682;
assign v_70685 = v_70682 & v_70684;
assign v_70687 = v_70580 & v_70686;
assign v_70689 = v_66678;
assign v_70691 = v_70688 & v_70690;
assign v_70693 = v_70577 & v_70692;
assign v_70695 = v_4194;
assign v_70697 = v_70694 & v_70696;
assign v_70699 = v_70574 & v_70698;
assign v_70701 = v_4190;
assign v_70703 = v_70700 & v_70702;
assign v_70705 = v_70571 & v_70704;
assign v_70707 = v_4186;
assign v_70709 = v_70706 & v_70708;
assign v_70711 = v_70568 & v_70710;
assign v_70713 = v_4182;
assign v_70715 = v_70712 & v_70714;
assign v_70717 = ~v_70716;
assign v_70719 = v_66726;
assign v_70720 = v_4247;
assign v_70721 = v_70720;
assign v_70722 = v_70719 & v_70721;
assign v_70723 = v_70722;
assign v_70724 = v_70613 & v_70723;
assign v_70726 = v_70623 & v_70725;
assign v_70727 = v_70612 & v_70723;
assign v_70729 = v_70610 & v_70728;
assign v_70731 = v_70629 & v_70730;
assign v_70732 = v_70609 & v_70728;
assign v_70734 = v_70607 & v_70733;
assign v_70736 = v_70635 & v_70735;
assign v_70737 = v_70606 & v_70733;
assign v_70739 = v_70604 & v_70738;
assign v_70741 = v_70641 & v_70740;
assign v_70742 = v_70603 & v_70738;
assign v_70744 = v_70601 & v_70743;
assign v_70746 = v_70647 & v_70745;
assign v_70747 = v_70600 & v_70743;
assign v_70749 = v_70598 & v_70748;
assign v_70751 = v_70653 & v_70750;
assign v_70752 = v_70597 & v_70748;
assign v_70754 = v_70595 & v_70753;
assign v_70756 = v_70659 & v_70755;
assign v_70757 = v_70594 & v_70753;
assign v_70759 = v_70592 & v_70758;
assign v_70761 = v_70665 & v_70760;
assign v_70762 = v_70591 & v_70758;
assign v_70764 = v_70589 & v_70763;
assign v_70766 = v_70671 & v_70765;
assign v_70767 = v_70588 & v_70763;
assign v_70769 = v_70586 & v_70768;
assign v_70771 = v_70677 & v_70770;
assign v_70772 = v_70585 & v_70768;
assign v_70774 = v_70583 & v_70773;
assign v_70776 = v_70683 & v_70775;
assign v_70777 = v_70582 & v_70773;
assign v_70779 = v_70580 & v_70778;
assign v_70781 = v_70689 & v_70780;
assign v_70782 = v_70579 & v_70778;
assign v_70784 = v_70577 & v_70783;
assign v_70786 = v_70695 & v_70785;
assign v_70787 = v_70576 & v_70783;
assign v_70789 = v_70574 & v_70788;
assign v_70791 = v_70701 & v_70790;
assign v_70792 = v_70573 & v_70788;
assign v_70794 = v_70571 & v_70793;
assign v_70796 = v_70707 & v_70795;
assign v_70797 = v_70570 & v_70793;
assign v_70799 = v_70568 & v_70798;
assign v_70801 = v_70713 & v_70800;
assign v_70802 = v_70567 & v_70798;
assign v_70804 = v_70716;
assign v_70806 = v_70718 & v_70805;
assign v_70807 = v_70806;
assign v_70810 = v_277;
assign v_70811 = v_5 & v_70810;
assign v_70812 = v_190;
assign v_70813 = ~v_5 & v_70812;
assign v_70815 = v_70814;
assign v_70816 = v_535;
assign v_70817 = v_282 & v_70816;
assign v_70818 = v_448;
assign v_70819 = ~v_282 & v_70818;
assign v_70821 = v_70820;
assign v_70822 = v_70815 & v_70821;
assign v_70823 = v_70822;
assign v_70824 = v_795;
assign v_70825 = v_542 & v_70824;
assign v_70826 = v_708;
assign v_70827 = ~v_542 & v_70826;
assign v_70829 = v_70828;
assign v_70830 = v_70823 & v_70829;
assign v_70831 = v_70830;
assign v_70832 = v_1055;
assign v_70833 = v_802 & v_70832;
assign v_70834 = v_968;
assign v_70835 = ~v_802 & v_70834;
assign v_70837 = v_70836;
assign v_70838 = v_70831 & v_70837;
assign v_70839 = v_70838;
assign v_70840 = v_1315;
assign v_70841 = v_1062 & v_70840;
assign v_70842 = v_1228;
assign v_70843 = ~v_1062 & v_70842;
assign v_70845 = v_70844;
assign v_70846 = v_70839 & v_70845;
assign v_70847 = v_70846;
assign v_70848 = v_1575;
assign v_70849 = v_1322 & v_70848;
assign v_70850 = v_1488;
assign v_70851 = ~v_1322 & v_70850;
assign v_70853 = v_70852;
assign v_70854 = v_70847 & v_70853;
assign v_70855 = v_70854;
assign v_70856 = v_1835;
assign v_70857 = v_1582 & v_70856;
assign v_70858 = v_1748;
assign v_70859 = ~v_1582 & v_70858;
assign v_70861 = v_70860;
assign v_70862 = v_70855 & v_70861;
assign v_70863 = v_70862;
assign v_70864 = v_2095;
assign v_70865 = v_1842 & v_70864;
assign v_70866 = v_2008;
assign v_70867 = ~v_1842 & v_70866;
assign v_70869 = v_70868;
assign v_70870 = v_70863 & v_70869;
assign v_70871 = v_70870;
assign v_70872 = v_2355;
assign v_70873 = v_2102 & v_70872;
assign v_70874 = v_2268;
assign v_70875 = ~v_2102 & v_70874;
assign v_70877 = v_70876;
assign v_70878 = v_70871 & v_70877;
assign v_70879 = v_70878;
assign v_70880 = v_2615;
assign v_70881 = v_2362 & v_70880;
assign v_70882 = v_2528;
assign v_70883 = ~v_2362 & v_70882;
assign v_70885 = v_70884;
assign v_70886 = v_70879 & v_70885;
assign v_70887 = v_70886;
assign v_70888 = v_2875;
assign v_70889 = v_2622 & v_70888;
assign v_70890 = v_2788;
assign v_70891 = ~v_2622 & v_70890;
assign v_70893 = v_70892;
assign v_70894 = v_70887 & v_70893;
assign v_70895 = v_70894;
assign v_70896 = v_3135;
assign v_70897 = v_2882 & v_70896;
assign v_70898 = v_3048;
assign v_70899 = ~v_2882 & v_70898;
assign v_70901 = v_70900;
assign v_70902 = v_70895 & v_70901;
assign v_70903 = v_70902;
assign v_70904 = v_3395;
assign v_70905 = v_3142 & v_70904;
assign v_70906 = v_3308;
assign v_70907 = ~v_3142 & v_70906;
assign v_70909 = v_70908;
assign v_70910 = v_70903 & v_70909;
assign v_70911 = v_70910;
assign v_70912 = v_3655;
assign v_70913 = v_3402 & v_70912;
assign v_70914 = v_3568;
assign v_70915 = ~v_3402 & v_70914;
assign v_70917 = v_70916;
assign v_70918 = v_70911 & v_70917;
assign v_70919 = v_70918;
assign v_70920 = v_3915;
assign v_70921 = v_3662 & v_70920;
assign v_70922 = v_3828;
assign v_70923 = ~v_3662 & v_70922;
assign v_70925 = v_70924;
assign v_70926 = v_70919 & v_70925;
assign v_70927 = v_70926;
assign v_70928 = v_4175;
assign v_70929 = v_3922 & v_70928;
assign v_70930 = v_4088;
assign v_70931 = ~v_3922 & v_70930;
assign v_70933 = v_70932;
assign v_70934 = v_70927 & v_70933;
assign v_70935 = v_70934;
assign v_70936 = v_4348;
assign v_70937 = v_4435 & v_70936;
assign v_70938 = ~v_4348;
assign v_70939 = v_4347 & v_70938;
assign v_70941 = v_70940;
assign v_70942 = v_70935 & v_70941;
assign v_70943 = v_70942;
assign v_70944 = v_4695;
assign v_70945 = v_4442 & v_70944;
assign v_70946 = v_4608;
assign v_70947 = ~v_4442 & v_70946;
assign v_70949 = v_70948;
assign v_70950 = v_70943 & v_70949;
assign v_70951 = v_70950;
assign v_70952 = v_4938;
assign v_70953 = v_4702 & v_70952;
assign v_70954 = v_4851;
assign v_70955 = ~v_4702 & v_70954;
assign v_70957 = v_70956;
assign v_70958 = v_70951 & v_70957;
assign v_70959 = v_70958;
assign v_70960 = v_5181;
assign v_70961 = v_4945 & v_70960;
assign v_70962 = v_5094;
assign v_70963 = ~v_4945 & v_70962;
assign v_70965 = v_70964;
assign v_70966 = v_70959 & v_70965;
assign v_70967 = v_70966;
assign v_70968 = v_5424;
assign v_70969 = v_5188 & v_70968;
assign v_70970 = v_5337;
assign v_70971 = ~v_5188 & v_70970;
assign v_70973 = v_70972;
assign v_70974 = v_70967 & v_70973;
assign v_70975 = v_70974;
assign v_70976 = v_5667;
assign v_70977 = v_5431 & v_70976;
assign v_70978 = v_5580;
assign v_70979 = ~v_5431 & v_70978;
assign v_70981 = v_70980;
assign v_70982 = v_70975 & v_70981;
assign v_70983 = v_70982;
assign v_70984 = v_5910;
assign v_70985 = v_5674 & v_70984;
assign v_70986 = v_5823;
assign v_70987 = ~v_5674 & v_70986;
assign v_70989 = v_70988;
assign v_70990 = v_70983 & v_70989;
assign v_70991 = v_70990;
assign v_70992 = v_6153;
assign v_70993 = v_5917 & v_70992;
assign v_70994 = v_6066;
assign v_70995 = ~v_5917 & v_70994;
assign v_70997 = v_70996;
assign v_70998 = v_70991 & v_70997;
assign v_70999 = v_70998;
assign v_71000 = v_6396;
assign v_71001 = v_6160 & v_71000;
assign v_71002 = v_6309;
assign v_71003 = ~v_6160 & v_71002;
assign v_71005 = v_71004;
assign v_71006 = v_70999 & v_71005;
assign v_71007 = v_71006;
assign v_71008 = v_6639;
assign v_71009 = v_6403 & v_71008;
assign v_71010 = v_6552;
assign v_71011 = ~v_6403 & v_71010;
assign v_71013 = v_71012;
assign v_71014 = v_71007 & v_71013;
assign v_71015 = v_71014;
assign v_71016 = v_6882;
assign v_71017 = v_6646 & v_71016;
assign v_71018 = v_6795;
assign v_71019 = ~v_6646 & v_71018;
assign v_71021 = v_71020;
assign v_71022 = v_71015 & v_71021;
assign v_71023 = v_71022;
assign v_71024 = v_7125;
assign v_71025 = v_6889 & v_71024;
assign v_71026 = v_7038;
assign v_71027 = ~v_6889 & v_71026;
assign v_71029 = v_71028;
assign v_71030 = v_71023 & v_71029;
assign v_71031 = v_71030;
assign v_71032 = v_7368;
assign v_71033 = v_7132 & v_71032;
assign v_71034 = v_7281;
assign v_71035 = ~v_7132 & v_71034;
assign v_71037 = v_71036;
assign v_71038 = v_71031 & v_71037;
assign v_71039 = v_71038;
assign v_71040 = v_7611;
assign v_71041 = v_7375 & v_71040;
assign v_71042 = v_7524;
assign v_71043 = ~v_7375 & v_71042;
assign v_71045 = v_71044;
assign v_71046 = v_71039 & v_71045;
assign v_71047 = v_71046;
assign v_71048 = v_7854;
assign v_71049 = v_7618 & v_71048;
assign v_71050 = v_7767;
assign v_71051 = ~v_7618 & v_71050;
assign v_71053 = v_71052;
assign v_71054 = v_71047 & v_71053;
assign v_71055 = v_71054;
assign v_71056 = v_8097;
assign v_71057 = v_7861 & v_71056;
assign v_71058 = v_8010;
assign v_71059 = ~v_7861 & v_71058;
assign v_71061 = v_71060;
assign v_71062 = v_71055 & v_71061;
assign v_71063 = v_71062;
assign v_71064 = v_8340;
assign v_71065 = v_8104 & v_71064;
assign v_71066 = v_8253;
assign v_71067 = ~v_8104 & v_71066;
assign v_71069 = v_71068;
assign v_71070 = v_71063 & v_71069;
assign v_71071 = v_71070;
assign v_71072 = v_8496;
assign v_71073 = v_8583 & v_71072;
assign v_71074 = ~v_8496;
assign v_71075 = v_8495 & v_71074;
assign v_71077 = v_71076;
assign v_71078 = v_71071 & v_71077;
assign v_71079 = v_71078;
assign v_71080 = v_8843;
assign v_71081 = v_8590 & v_71080;
assign v_71082 = v_8756;
assign v_71083 = ~v_8590 & v_71082;
assign v_71085 = v_71084;
assign v_71086 = v_71079 & v_71085;
assign v_71087 = v_71086;
assign v_71088 = v_9086;
assign v_71089 = v_8850 & v_71088;
assign v_71090 = v_8999;
assign v_71091 = ~v_8850 & v_71090;
assign v_71093 = v_71092;
assign v_71094 = v_71087 & v_71093;
assign v_71095 = v_71094;
assign v_71096 = v_9329;
assign v_71097 = v_9093 & v_71096;
assign v_71098 = v_9242;
assign v_71099 = ~v_9093 & v_71098;
assign v_71101 = v_71100;
assign v_71102 = v_71095 & v_71101;
assign v_71103 = v_71102;
assign v_71104 = v_9572;
assign v_71105 = v_9336 & v_71104;
assign v_71106 = v_9485;
assign v_71107 = ~v_9336 & v_71106;
assign v_71109 = v_71108;
assign v_71110 = v_71103 & v_71109;
assign v_71111 = v_71110;
assign v_71112 = v_9815;
assign v_71113 = v_9579 & v_71112;
assign v_71114 = v_9728;
assign v_71115 = ~v_9579 & v_71114;
assign v_71117 = v_71116;
assign v_71118 = v_71111 & v_71117;
assign v_71119 = v_71118;
assign v_71120 = v_10058;
assign v_71121 = v_9822 & v_71120;
assign v_71122 = v_9971;
assign v_71123 = ~v_9822 & v_71122;
assign v_71125 = v_71124;
assign v_71126 = v_71119 & v_71125;
assign v_71127 = v_71126;
assign v_71128 = v_10301;
assign v_71129 = v_10065 & v_71128;
assign v_71130 = v_10214;
assign v_71131 = ~v_10065 & v_71130;
assign v_71133 = v_71132;
assign v_71134 = v_71127 & v_71133;
assign v_71135 = v_71134;
assign v_71136 = v_10544;
assign v_71137 = v_10308 & v_71136;
assign v_71138 = v_10457;
assign v_71139 = ~v_10308 & v_71138;
assign v_71141 = v_71140;
assign v_71142 = v_71135 & v_71141;
assign v_71143 = v_71142;
assign v_71144 = v_10787;
assign v_71145 = v_10551 & v_71144;
assign v_71146 = v_10700;
assign v_71147 = ~v_10551 & v_71146;
assign v_71149 = v_71148;
assign v_71150 = v_71143 & v_71149;
assign v_71151 = v_71150;
assign v_71152 = v_11030;
assign v_71153 = v_10794 & v_71152;
assign v_71154 = v_10943;
assign v_71155 = ~v_10794 & v_71154;
assign v_71157 = v_71156;
assign v_71158 = v_71151 & v_71157;
assign v_71159 = v_71158;
assign v_71160 = v_11273;
assign v_71161 = v_11037 & v_71160;
assign v_71162 = v_11186;
assign v_71163 = ~v_11037 & v_71162;
assign v_71165 = v_71164;
assign v_71166 = v_71159 & v_71165;
assign v_71167 = v_71166;
assign v_71168 = v_11516;
assign v_71169 = v_11280 & v_71168;
assign v_71170 = v_11429;
assign v_71171 = ~v_11280 & v_71170;
assign v_71173 = v_71172;
assign v_71174 = v_71167 & v_71173;
assign v_71175 = v_71174;
assign v_71176 = v_11759;
assign v_71177 = v_11523 & v_71176;
assign v_71178 = v_11672;
assign v_71179 = ~v_11523 & v_71178;
assign v_71181 = v_71180;
assign v_71182 = v_71175 & v_71181;
assign v_71183 = v_71182;
assign v_71184 = v_12002;
assign v_71185 = v_11766 & v_71184;
assign v_71186 = v_11915;
assign v_71187 = ~v_11766 & v_71186;
assign v_71189 = v_71188;
assign v_71190 = v_71183 & v_71189;
assign v_71191 = v_71190;
assign v_71192 = v_12245;
assign v_71193 = v_12009 & v_71192;
assign v_71194 = v_12158;
assign v_71195 = ~v_12009 & v_71194;
assign v_71197 = v_71196;
assign v_71198 = v_71191 & v_71197;
assign v_71199 = v_71198;
assign v_71200 = v_12488;
assign v_71201 = v_12252 & v_71200;
assign v_71202 = v_12401;
assign v_71203 = ~v_12252 & v_71202;
assign v_71205 = v_71204;
assign v_71206 = v_71199 & v_71205;
assign v_71207 = v_71206;
assign v_71208 = v_12644;
assign v_71209 = v_12731 & v_71208;
assign v_71210 = ~v_12644;
assign v_71211 = v_12643 & v_71210;
assign v_71213 = v_71212;
assign v_71214 = v_71207 & v_71213;
assign v_71215 = v_71214;
assign v_71216 = v_12991;
assign v_71217 = v_12738 & v_71216;
assign v_71218 = v_12904;
assign v_71219 = ~v_12738 & v_71218;
assign v_71221 = v_71220;
assign v_71222 = v_71215 & v_71221;
assign v_71223 = v_71222;
assign v_71224 = v_13234;
assign v_71225 = v_12998 & v_71224;
assign v_71226 = v_13147;
assign v_71227 = ~v_12998 & v_71226;
assign v_71229 = v_71228;
assign v_71230 = v_71223 & v_71229;
assign v_71231 = v_71230;
assign v_71232 = v_13477;
assign v_71233 = v_13241 & v_71232;
assign v_71234 = v_13390;
assign v_71235 = ~v_13241 & v_71234;
assign v_71237 = v_71236;
assign v_71238 = v_71231 & v_71237;
assign v_71239 = v_71238;
assign v_71240 = v_13720;
assign v_71241 = v_13484 & v_71240;
assign v_71242 = v_13633;
assign v_71243 = ~v_13484 & v_71242;
assign v_71245 = v_71244;
assign v_71246 = v_71239 & v_71245;
assign v_71247 = v_71246;
assign v_71248 = v_13963;
assign v_71249 = v_13727 & v_71248;
assign v_71250 = v_13876;
assign v_71251 = ~v_13727 & v_71250;
assign v_71253 = v_71252;
assign v_71254 = v_71247 & v_71253;
assign v_71255 = v_71254;
assign v_71256 = v_14206;
assign v_71257 = v_13970 & v_71256;
assign v_71258 = v_14119;
assign v_71259 = ~v_13970 & v_71258;
assign v_71261 = v_71260;
assign v_71262 = v_71255 & v_71261;
assign v_71263 = v_71262;
assign v_71264 = v_14449;
assign v_71265 = v_14213 & v_71264;
assign v_71266 = v_14362;
assign v_71267 = ~v_14213 & v_71266;
assign v_71269 = v_71268;
assign v_71270 = v_71263 & v_71269;
assign v_71271 = v_71270;
assign v_71272 = v_14692;
assign v_71273 = v_14456 & v_71272;
assign v_71274 = v_14605;
assign v_71275 = ~v_14456 & v_71274;
assign v_71277 = v_71276;
assign v_71278 = v_71271 & v_71277;
assign v_71279 = v_71278;
assign v_71280 = v_14935;
assign v_71281 = v_14699 & v_71280;
assign v_71282 = v_14848;
assign v_71283 = ~v_14699 & v_71282;
assign v_71285 = v_71284;
assign v_71286 = v_71279 & v_71285;
assign v_71287 = v_71286;
assign v_71288 = v_15178;
assign v_71289 = v_14942 & v_71288;
assign v_71290 = v_15091;
assign v_71291 = ~v_14942 & v_71290;
assign v_71293 = v_71292;
assign v_71294 = v_71287 & v_71293;
assign v_71295 = v_71294;
assign v_71296 = v_15421;
assign v_71297 = v_15185 & v_71296;
assign v_71298 = v_15334;
assign v_71299 = ~v_15185 & v_71298;
assign v_71301 = v_71300;
assign v_71302 = v_71295 & v_71301;
assign v_71303 = v_71302;
assign v_71304 = v_15664;
assign v_71305 = v_15428 & v_71304;
assign v_71306 = v_15577;
assign v_71307 = ~v_15428 & v_71306;
assign v_71309 = v_71308;
assign v_71310 = v_71303 & v_71309;
assign v_71311 = v_71310;
assign v_71312 = v_15907;
assign v_71313 = v_15671 & v_71312;
assign v_71314 = v_15820;
assign v_71315 = ~v_15671 & v_71314;
assign v_71317 = v_71316;
assign v_71318 = v_71311 & v_71317;
assign v_71319 = v_71318;
assign v_71320 = v_16150;
assign v_71321 = v_15914 & v_71320;
assign v_71322 = v_16063;
assign v_71323 = ~v_15914 & v_71322;
assign v_71325 = v_71324;
assign v_71326 = v_71319 & v_71325;
assign v_71327 = v_71326;
assign v_71328 = v_16393;
assign v_71329 = v_16157 & v_71328;
assign v_71330 = v_16306;
assign v_71331 = ~v_16157 & v_71330;
assign v_71333 = v_71332;
assign v_71334 = v_71327 & v_71333;
assign v_71335 = v_71334;
assign v_71336 = v_16636;
assign v_71337 = v_16400 & v_71336;
assign v_71338 = v_16549;
assign v_71339 = ~v_16400 & v_71338;
assign v_71341 = v_71340;
assign v_71342 = v_71335 & v_71341;
assign v_71343 = v_71342;
assign v_71344 = v_16792;
assign v_71345 = v_16879 & v_71344;
assign v_71346 = ~v_16792;
assign v_71347 = v_16791 & v_71346;
assign v_71349 = v_71348;
assign v_71350 = v_71343 & v_71349;
assign v_71351 = v_71350;
assign v_71352 = v_17139;
assign v_71353 = v_16886 & v_71352;
assign v_71354 = v_17052;
assign v_71355 = ~v_16886 & v_71354;
assign v_71357 = v_71356;
assign v_71358 = v_71351 & v_71357;
assign v_71359 = v_71358;
assign v_71360 = v_17382;
assign v_71361 = v_17146 & v_71360;
assign v_71362 = v_17295;
assign v_71363 = ~v_17146 & v_71362;
assign v_71365 = v_71364;
assign v_71366 = v_71359 & v_71365;
assign v_71367 = v_71366;
assign v_71368 = v_17625;
assign v_71369 = v_17389 & v_71368;
assign v_71370 = v_17538;
assign v_71371 = ~v_17389 & v_71370;
assign v_71373 = v_71372;
assign v_71374 = v_71367 & v_71373;
assign v_71375 = v_71374;
assign v_71376 = v_17868;
assign v_71377 = v_17632 & v_71376;
assign v_71378 = v_17781;
assign v_71379 = ~v_17632 & v_71378;
assign v_71381 = v_71380;
assign v_71382 = v_71375 & v_71381;
assign v_71383 = v_71382;
assign v_71384 = v_18111;
assign v_71385 = v_17875 & v_71384;
assign v_71386 = v_18024;
assign v_71387 = ~v_17875 & v_71386;
assign v_71389 = v_71388;
assign v_71390 = v_71383 & v_71389;
assign v_71391 = v_71390;
assign v_71392 = v_18354;
assign v_71393 = v_18118 & v_71392;
assign v_71394 = v_18267;
assign v_71395 = ~v_18118 & v_71394;
assign v_71397 = v_71396;
assign v_71398 = v_71391 & v_71397;
assign v_71399 = v_71398;
assign v_71400 = v_18597;
assign v_71401 = v_18361 & v_71400;
assign v_71402 = v_18510;
assign v_71403 = ~v_18361 & v_71402;
assign v_71405 = v_71404;
assign v_71406 = v_71399 & v_71405;
assign v_71407 = v_71406;
assign v_71408 = v_18840;
assign v_71409 = v_18604 & v_71408;
assign v_71410 = v_18753;
assign v_71411 = ~v_18604 & v_71410;
assign v_71413 = v_71412;
assign v_71414 = v_71407 & v_71413;
assign v_71415 = v_71414;
assign v_71416 = v_19083;
assign v_71417 = v_18847 & v_71416;
assign v_71418 = v_18996;
assign v_71419 = ~v_18847 & v_71418;
assign v_71421 = v_71420;
assign v_71422 = v_71415 & v_71421;
assign v_71423 = v_71422;
assign v_71424 = v_19326;
assign v_71425 = v_19090 & v_71424;
assign v_71426 = v_19239;
assign v_71427 = ~v_19090 & v_71426;
assign v_71429 = v_71428;
assign v_71430 = v_71423 & v_71429;
assign v_71431 = v_71430;
assign v_71432 = v_19569;
assign v_71433 = v_19333 & v_71432;
assign v_71434 = v_19482;
assign v_71435 = ~v_19333 & v_71434;
assign v_71437 = v_71436;
assign v_71438 = v_71431 & v_71437;
assign v_71439 = v_71438;
assign v_71440 = v_19812;
assign v_71441 = v_19576 & v_71440;
assign v_71442 = v_19725;
assign v_71443 = ~v_19576 & v_71442;
assign v_71445 = v_71444;
assign v_71446 = v_71439 & v_71445;
assign v_71447 = v_71446;
assign v_71448 = v_20055;
assign v_71449 = v_19819 & v_71448;
assign v_71450 = v_19968;
assign v_71451 = ~v_19819 & v_71450;
assign v_71453 = v_71452;
assign v_71454 = v_71447 & v_71453;
assign v_71455 = v_71454;
assign v_71456 = v_20298;
assign v_71457 = v_20062 & v_71456;
assign v_71458 = v_20211;
assign v_71459 = ~v_20062 & v_71458;
assign v_71461 = v_71460;
assign v_71462 = v_71455 & v_71461;
assign v_71463 = v_71462;
assign v_71464 = v_20541;
assign v_71465 = v_20305 & v_71464;
assign v_71466 = v_20454;
assign v_71467 = ~v_20305 & v_71466;
assign v_71469 = v_71468;
assign v_71470 = v_71463 & v_71469;
assign v_71471 = v_71470;
assign v_71472 = v_20784;
assign v_71473 = v_20548 & v_71472;
assign v_71474 = v_20697;
assign v_71475 = ~v_20548 & v_71474;
assign v_71477 = v_71476;
assign v_71478 = v_71471 & v_71477;
assign v_71479 = v_71478;
assign v_71480 = v_20940;
assign v_71481 = v_21027 & v_71480;
assign v_71482 = ~v_20940;
assign v_71483 = v_20939 & v_71482;
assign v_71485 = v_71484;
assign v_71486 = v_71479 & v_71485;
assign v_71487 = v_71486;
assign v_71488 = v_21287;
assign v_71489 = v_21034 & v_71488;
assign v_71490 = v_21200;
assign v_71491 = ~v_21034 & v_71490;
assign v_71493 = v_71492;
assign v_71494 = v_71487 & v_71493;
assign v_71495 = v_71494;
assign v_71496 = v_21530;
assign v_71497 = v_21294 & v_71496;
assign v_71498 = v_21443;
assign v_71499 = ~v_21294 & v_71498;
assign v_71501 = v_71500;
assign v_71502 = v_71495 & v_71501;
assign v_71503 = v_71502;
assign v_71504 = v_21773;
assign v_71505 = v_21537 & v_71504;
assign v_71506 = v_21686;
assign v_71507 = ~v_21537 & v_71506;
assign v_71509 = v_71508;
assign v_71510 = v_71503 & v_71509;
assign v_71511 = v_71510;
assign v_71512 = v_22016;
assign v_71513 = v_21780 & v_71512;
assign v_71514 = v_21929;
assign v_71515 = ~v_21780 & v_71514;
assign v_71517 = v_71516;
assign v_71518 = v_71511 & v_71517;
assign v_71519 = v_71518;
assign v_71520 = v_22259;
assign v_71521 = v_22023 & v_71520;
assign v_71522 = v_22172;
assign v_71523 = ~v_22023 & v_71522;
assign v_71525 = v_71524;
assign v_71526 = v_71519 & v_71525;
assign v_71527 = v_71526;
assign v_71528 = v_22502;
assign v_71529 = v_22266 & v_71528;
assign v_71530 = v_22415;
assign v_71531 = ~v_22266 & v_71530;
assign v_71533 = v_71532;
assign v_71534 = v_71527 & v_71533;
assign v_71535 = v_71534;
assign v_71536 = v_22745;
assign v_71537 = v_22509 & v_71536;
assign v_71538 = v_22658;
assign v_71539 = ~v_22509 & v_71538;
assign v_71541 = v_71540;
assign v_71542 = v_71535 & v_71541;
assign v_71543 = v_71542;
assign v_71544 = v_22988;
assign v_71545 = v_22752 & v_71544;
assign v_71546 = v_22901;
assign v_71547 = ~v_22752 & v_71546;
assign v_71549 = v_71548;
assign v_71550 = v_71543 & v_71549;
assign v_71551 = v_71550;
assign v_71552 = v_23231;
assign v_71553 = v_22995 & v_71552;
assign v_71554 = v_23144;
assign v_71555 = ~v_22995 & v_71554;
assign v_71557 = v_71556;
assign v_71558 = v_71551 & v_71557;
assign v_71559 = v_71558;
assign v_71560 = v_23474;
assign v_71561 = v_23238 & v_71560;
assign v_71562 = v_23387;
assign v_71563 = ~v_23238 & v_71562;
assign v_71565 = v_71564;
assign v_71566 = v_71559 & v_71565;
assign v_71567 = v_71566;
assign v_71568 = v_23717;
assign v_71569 = v_23481 & v_71568;
assign v_71570 = v_23630;
assign v_71571 = ~v_23481 & v_71570;
assign v_71573 = v_71572;
assign v_71574 = v_71567 & v_71573;
assign v_71575 = v_71574;
assign v_71576 = v_23960;
assign v_71577 = v_23724 & v_71576;
assign v_71578 = v_23873;
assign v_71579 = ~v_23724 & v_71578;
assign v_71581 = v_71580;
assign v_71582 = v_71575 & v_71581;
assign v_71583 = v_71582;
assign v_71584 = v_24203;
assign v_71585 = v_23967 & v_71584;
assign v_71586 = v_24116;
assign v_71587 = ~v_23967 & v_71586;
assign v_71589 = v_71588;
assign v_71590 = v_71583 & v_71589;
assign v_71591 = v_71590;
assign v_71592 = v_24446;
assign v_71593 = v_24210 & v_71592;
assign v_71594 = v_24359;
assign v_71595 = ~v_24210 & v_71594;
assign v_71597 = v_71596;
assign v_71598 = v_71591 & v_71597;
assign v_71599 = v_71598;
assign v_71600 = v_24689;
assign v_71601 = v_24453 & v_71600;
assign v_71602 = v_24602;
assign v_71603 = ~v_24453 & v_71602;
assign v_71605 = v_71604;
assign v_71606 = v_71599 & v_71605;
assign v_71607 = v_71606;
assign v_71608 = v_24932;
assign v_71609 = v_24696 & v_71608;
assign v_71610 = v_24845;
assign v_71611 = ~v_24696 & v_71610;
assign v_71613 = v_71612;
assign v_71614 = v_71607 & v_71613;
assign v_71615 = v_71614;
assign v_71616 = v_25088;
assign v_71617 = v_25175 & v_71616;
assign v_71618 = ~v_25088;
assign v_71619 = v_25087 & v_71618;
assign v_71621 = v_71620;
assign v_71622 = v_71615 & v_71621;
assign v_71623 = v_71622;
assign v_71624 = v_25435;
assign v_71625 = v_25182 & v_71624;
assign v_71626 = v_25348;
assign v_71627 = ~v_25182 & v_71626;
assign v_71629 = v_71628;
assign v_71630 = v_71623 & v_71629;
assign v_71631 = v_71630;
assign v_71632 = v_25678;
assign v_71633 = v_25442 & v_71632;
assign v_71634 = v_25591;
assign v_71635 = ~v_25442 & v_71634;
assign v_71637 = v_71636;
assign v_71638 = v_71631 & v_71637;
assign v_71639 = v_71638;
assign v_71640 = v_25921;
assign v_71641 = v_25685 & v_71640;
assign v_71642 = v_25834;
assign v_71643 = ~v_25685 & v_71642;
assign v_71645 = v_71644;
assign v_71646 = v_71639 & v_71645;
assign v_71647 = v_71646;
assign v_71648 = v_26164;
assign v_71649 = v_25928 & v_71648;
assign v_71650 = v_26077;
assign v_71651 = ~v_25928 & v_71650;
assign v_71653 = v_71652;
assign v_71654 = v_71647 & v_71653;
assign v_71655 = v_71654;
assign v_71656 = v_26407;
assign v_71657 = v_26171 & v_71656;
assign v_71658 = v_26320;
assign v_71659 = ~v_26171 & v_71658;
assign v_71661 = v_71660;
assign v_71662 = v_71655 & v_71661;
assign v_71663 = v_71662;
assign v_71664 = v_26650;
assign v_71665 = v_26414 & v_71664;
assign v_71666 = v_26563;
assign v_71667 = ~v_26414 & v_71666;
assign v_71669 = v_71668;
assign v_71670 = v_71663 & v_71669;
assign v_71671 = v_71670;
assign v_71672 = v_26893;
assign v_71673 = v_26657 & v_71672;
assign v_71674 = v_26806;
assign v_71675 = ~v_26657 & v_71674;
assign v_71677 = v_71676;
assign v_71678 = v_71671 & v_71677;
assign v_71679 = v_71678;
assign v_71680 = v_27136;
assign v_71681 = v_26900 & v_71680;
assign v_71682 = v_27049;
assign v_71683 = ~v_26900 & v_71682;
assign v_71685 = v_71684;
assign v_71686 = v_71679 & v_71685;
assign v_71687 = v_71686;
assign v_71688 = v_27379;
assign v_71689 = v_27143 & v_71688;
assign v_71690 = v_27292;
assign v_71691 = ~v_27143 & v_71690;
assign v_71693 = v_71692;
assign v_71694 = v_71687 & v_71693;
assign v_71695 = v_71694;
assign v_71696 = v_27622;
assign v_71697 = v_27386 & v_71696;
assign v_71698 = v_27535;
assign v_71699 = ~v_27386 & v_71698;
assign v_71701 = v_71700;
assign v_71702 = v_71695 & v_71701;
assign v_71703 = v_71702;
assign v_71704 = v_27865;
assign v_71705 = v_27629 & v_71704;
assign v_71706 = v_27778;
assign v_71707 = ~v_27629 & v_71706;
assign v_71709 = v_71708;
assign v_71710 = v_71703 & v_71709;
assign v_71711 = v_71710;
assign v_71712 = v_28108;
assign v_71713 = v_27872 & v_71712;
assign v_71714 = v_28021;
assign v_71715 = ~v_27872 & v_71714;
assign v_71717 = v_71716;
assign v_71718 = v_71711 & v_71717;
assign v_71719 = v_71718;
assign v_71720 = v_28351;
assign v_71721 = v_28115 & v_71720;
assign v_71722 = v_28264;
assign v_71723 = ~v_28115 & v_71722;
assign v_71725 = v_71724;
assign v_71726 = v_71719 & v_71725;
assign v_71727 = v_71726;
assign v_71728 = v_28594;
assign v_71729 = v_28358 & v_71728;
assign v_71730 = v_28507;
assign v_71731 = ~v_28358 & v_71730;
assign v_71733 = v_71732;
assign v_71734 = v_71727 & v_71733;
assign v_71735 = v_71734;
assign v_71736 = v_28837;
assign v_71737 = v_28601 & v_71736;
assign v_71738 = v_28750;
assign v_71739 = ~v_28601 & v_71738;
assign v_71741 = v_71740;
assign v_71742 = v_71735 & v_71741;
assign v_71743 = v_71742;
assign v_71744 = v_29080;
assign v_71745 = v_28844 & v_71744;
assign v_71746 = v_28993;
assign v_71747 = ~v_28844 & v_71746;
assign v_71749 = v_71748;
assign v_71750 = v_71743 & v_71749;
assign v_71751 = v_71750;
assign v_71752 = v_29236;
assign v_71753 = v_29323 & v_71752;
assign v_71754 = ~v_29236;
assign v_71755 = v_29235 & v_71754;
assign v_71757 = v_71756;
assign v_71758 = v_71751 & v_71757;
assign v_71759 = v_71758;
assign v_71760 = v_29583;
assign v_71761 = v_29330 & v_71760;
assign v_71762 = v_29496;
assign v_71763 = ~v_29330 & v_71762;
assign v_71765 = v_71764;
assign v_71766 = v_71759 & v_71765;
assign v_71767 = v_71766;
assign v_71768 = v_29826;
assign v_71769 = v_29590 & v_71768;
assign v_71770 = v_29739;
assign v_71771 = ~v_29590 & v_71770;
assign v_71773 = v_71772;
assign v_71774 = v_71767 & v_71773;
assign v_71775 = v_71774;
assign v_71776 = v_30069;
assign v_71777 = v_29833 & v_71776;
assign v_71778 = v_29982;
assign v_71779 = ~v_29833 & v_71778;
assign v_71781 = v_71780;
assign v_71782 = v_71775 & v_71781;
assign v_71783 = v_71782;
assign v_71784 = v_30312;
assign v_71785 = v_30076 & v_71784;
assign v_71786 = v_30225;
assign v_71787 = ~v_30076 & v_71786;
assign v_71789 = v_71788;
assign v_71790 = v_71783 & v_71789;
assign v_71791 = v_71790;
assign v_71792 = v_30555;
assign v_71793 = v_30319 & v_71792;
assign v_71794 = v_30468;
assign v_71795 = ~v_30319 & v_71794;
assign v_71797 = v_71796;
assign v_71798 = v_71791 & v_71797;
assign v_71799 = v_71798;
assign v_71800 = v_30798;
assign v_71801 = v_30562 & v_71800;
assign v_71802 = v_30711;
assign v_71803 = ~v_30562 & v_71802;
assign v_71805 = v_71804;
assign v_71806 = v_71799 & v_71805;
assign v_71807 = v_71806;
assign v_71808 = v_31041;
assign v_71809 = v_30805 & v_71808;
assign v_71810 = v_30954;
assign v_71811 = ~v_30805 & v_71810;
assign v_71813 = v_71812;
assign v_71814 = v_71807 & v_71813;
assign v_71815 = v_71814;
assign v_71816 = v_31284;
assign v_71817 = v_31048 & v_71816;
assign v_71818 = v_31197;
assign v_71819 = ~v_31048 & v_71818;
assign v_71821 = v_71820;
assign v_71822 = v_71815 & v_71821;
assign v_71823 = v_71822;
assign v_71824 = v_31527;
assign v_71825 = v_31291 & v_71824;
assign v_71826 = v_31440;
assign v_71827 = ~v_31291 & v_71826;
assign v_71829 = v_71828;
assign v_71830 = v_71823 & v_71829;
assign v_71831 = v_71830;
assign v_71832 = v_31770;
assign v_71833 = v_31534 & v_71832;
assign v_71834 = v_31683;
assign v_71835 = ~v_31534 & v_71834;
assign v_71837 = v_71836;
assign v_71838 = v_71831 & v_71837;
assign v_71839 = v_71838;
assign v_71840 = v_32013;
assign v_71841 = v_31777 & v_71840;
assign v_71842 = v_31926;
assign v_71843 = ~v_31777 & v_71842;
assign v_71845 = v_71844;
assign v_71846 = v_71839 & v_71845;
assign v_71847 = v_71846;
assign v_71848 = v_32256;
assign v_71849 = v_32020 & v_71848;
assign v_71850 = v_32169;
assign v_71851 = ~v_32020 & v_71850;
assign v_71853 = v_71852;
assign v_71854 = v_71847 & v_71853;
assign v_71855 = v_71854;
assign v_71856 = v_32499;
assign v_71857 = v_32263 & v_71856;
assign v_71858 = v_32412;
assign v_71859 = ~v_32263 & v_71858;
assign v_71861 = v_71860;
assign v_71862 = v_71855 & v_71861;
assign v_71863 = v_71862;
assign v_71864 = v_32742;
assign v_71865 = v_32506 & v_71864;
assign v_71866 = v_32655;
assign v_71867 = ~v_32506 & v_71866;
assign v_71869 = v_71868;
assign v_71870 = v_71863 & v_71869;
assign v_71871 = v_71870;
assign v_71872 = v_32985;
assign v_71873 = v_32749 & v_71872;
assign v_71874 = v_32898;
assign v_71875 = ~v_32749 & v_71874;
assign v_71877 = v_71876;
assign v_71878 = v_71871 & v_71877;
assign v_71879 = v_71878;
assign v_71880 = v_33228;
assign v_71881 = v_32992 & v_71880;
assign v_71882 = v_33141;
assign v_71883 = ~v_32992 & v_71882;
assign v_71885 = v_71884;
assign v_71886 = v_71879 & v_71885;
assign v_71887 = v_71886;
assign v_71888 = v_33384;
assign v_71889 = v_33471 & v_71888;
assign v_71890 = ~v_33384;
assign v_71891 = v_33383 & v_71890;
assign v_71893 = v_71892;
assign v_71894 = v_71887 & v_71893;
assign v_71895 = v_71894;
assign v_71896 = v_33731;
assign v_71897 = v_33478 & v_71896;
assign v_71898 = v_33644;
assign v_71899 = ~v_33478 & v_71898;
assign v_71901 = v_71900;
assign v_71902 = v_71895 & v_71901;
assign v_71903 = v_71902;
assign v_71904 = v_33974;
assign v_71905 = v_33738 & v_71904;
assign v_71906 = v_33887;
assign v_71907 = ~v_33738 & v_71906;
assign v_71909 = v_71908;
assign v_71910 = v_71903 & v_71909;
assign v_71911 = v_71910;
assign v_71912 = v_34217;
assign v_71913 = v_33981 & v_71912;
assign v_71914 = v_34130;
assign v_71915 = ~v_33981 & v_71914;
assign v_71917 = v_71916;
assign v_71918 = v_71911 & v_71917;
assign v_71919 = v_71918;
assign v_71920 = v_34460;
assign v_71921 = v_34224 & v_71920;
assign v_71922 = v_34373;
assign v_71923 = ~v_34224 & v_71922;
assign v_71925 = v_71924;
assign v_71926 = v_71919 & v_71925;
assign v_71927 = v_71926;
assign v_71928 = v_34703;
assign v_71929 = v_34467 & v_71928;
assign v_71930 = v_34616;
assign v_71931 = ~v_34467 & v_71930;
assign v_71933 = v_71932;
assign v_71934 = v_71927 & v_71933;
assign v_71935 = v_71934;
assign v_71936 = v_34946;
assign v_71937 = v_34710 & v_71936;
assign v_71938 = v_34859;
assign v_71939 = ~v_34710 & v_71938;
assign v_71941 = v_71940;
assign v_71942 = v_71935 & v_71941;
assign v_71943 = v_71942;
assign v_71944 = v_35189;
assign v_71945 = v_34953 & v_71944;
assign v_71946 = v_35102;
assign v_71947 = ~v_34953 & v_71946;
assign v_71949 = v_71948;
assign v_71950 = v_71943 & v_71949;
assign v_71951 = v_71950;
assign v_71952 = v_35432;
assign v_71953 = v_35196 & v_71952;
assign v_71954 = v_35345;
assign v_71955 = ~v_35196 & v_71954;
assign v_71957 = v_71956;
assign v_71958 = v_71951 & v_71957;
assign v_71959 = v_71958;
assign v_71960 = v_35675;
assign v_71961 = v_35439 & v_71960;
assign v_71962 = v_35588;
assign v_71963 = ~v_35439 & v_71962;
assign v_71965 = v_71964;
assign v_71966 = v_71959 & v_71965;
assign v_71967 = v_71966;
assign v_71968 = v_35918;
assign v_71969 = v_35682 & v_71968;
assign v_71970 = v_35831;
assign v_71971 = ~v_35682 & v_71970;
assign v_71973 = v_71972;
assign v_71974 = v_71967 & v_71973;
assign v_71975 = v_71974;
assign v_71976 = v_36161;
assign v_71977 = v_35925 & v_71976;
assign v_71978 = v_36074;
assign v_71979 = ~v_35925 & v_71978;
assign v_71981 = v_71980;
assign v_71982 = v_71975 & v_71981;
assign v_71983 = v_71982;
assign v_71984 = v_36404;
assign v_71985 = v_36168 & v_71984;
assign v_71986 = v_36317;
assign v_71987 = ~v_36168 & v_71986;
assign v_71989 = v_71988;
assign v_71990 = v_71983 & v_71989;
assign v_71991 = v_71990;
assign v_71992 = v_36647;
assign v_71993 = v_36411 & v_71992;
assign v_71994 = v_36560;
assign v_71995 = ~v_36411 & v_71994;
assign v_71997 = v_71996;
assign v_71998 = v_71991 & v_71997;
assign v_71999 = v_71998;
assign v_72000 = v_36890;
assign v_72001 = v_36654 & v_72000;
assign v_72002 = v_36803;
assign v_72003 = ~v_36654 & v_72002;
assign v_72005 = v_72004;
assign v_72006 = v_71999 & v_72005;
assign v_72007 = v_72006;
assign v_72008 = v_37133;
assign v_72009 = v_36897 & v_72008;
assign v_72010 = v_37046;
assign v_72011 = ~v_36897 & v_72010;
assign v_72013 = v_72012;
assign v_72014 = v_72007 & v_72013;
assign v_72015 = v_72014;
assign v_72016 = v_37376;
assign v_72017 = v_37140 & v_72016;
assign v_72018 = v_37289;
assign v_72019 = ~v_37140 & v_72018;
assign v_72021 = v_72020;
assign v_72022 = v_72015 & v_72021;
assign v_72023 = v_72022;
assign v_72024 = v_37532;
assign v_72025 = v_37619 & v_72024;
assign v_72026 = ~v_37532;
assign v_72027 = v_37531 & v_72026;
assign v_72029 = v_72028;
assign v_72030 = v_72023 & v_72029;
assign v_72031 = v_72030;
assign v_72032 = v_37879;
assign v_72033 = v_37626 & v_72032;
assign v_72034 = v_37792;
assign v_72035 = ~v_37626 & v_72034;
assign v_72037 = v_72036;
assign v_72038 = v_72031 & v_72037;
assign v_72039 = v_72038;
assign v_72040 = v_38122;
assign v_72041 = v_37886 & v_72040;
assign v_72042 = v_38035;
assign v_72043 = ~v_37886 & v_72042;
assign v_72045 = v_72044;
assign v_72046 = v_72039 & v_72045;
assign v_72047 = v_72046;
assign v_72048 = v_38365;
assign v_72049 = v_38129 & v_72048;
assign v_72050 = v_38278;
assign v_72051 = ~v_38129 & v_72050;
assign v_72053 = v_72052;
assign v_72054 = v_72047 & v_72053;
assign v_72055 = v_72054;
assign v_72056 = v_38608;
assign v_72057 = v_38372 & v_72056;
assign v_72058 = v_38521;
assign v_72059 = ~v_38372 & v_72058;
assign v_72061 = v_72060;
assign v_72062 = v_72055 & v_72061;
assign v_72063 = v_72062;
assign v_72064 = v_38851;
assign v_72065 = v_38615 & v_72064;
assign v_72066 = v_38764;
assign v_72067 = ~v_38615 & v_72066;
assign v_72069 = v_72068;
assign v_72070 = v_72063 & v_72069;
assign v_72071 = v_72070;
assign v_72072 = v_39094;
assign v_72073 = v_38858 & v_72072;
assign v_72074 = v_39007;
assign v_72075 = ~v_38858 & v_72074;
assign v_72077 = v_72076;
assign v_72078 = v_72071 & v_72077;
assign v_72079 = v_72078;
assign v_72080 = v_39337;
assign v_72081 = v_39101 & v_72080;
assign v_72082 = v_39250;
assign v_72083 = ~v_39101 & v_72082;
assign v_72085 = v_72084;
assign v_72086 = v_72079 & v_72085;
assign v_72087 = v_72086;
assign v_72088 = v_39580;
assign v_72089 = v_39344 & v_72088;
assign v_72090 = v_39493;
assign v_72091 = ~v_39344 & v_72090;
assign v_72093 = v_72092;
assign v_72094 = v_72087 & v_72093;
assign v_72095 = v_72094;
assign v_72096 = v_39823;
assign v_72097 = v_39587 & v_72096;
assign v_72098 = v_39736;
assign v_72099 = ~v_39587 & v_72098;
assign v_72101 = v_72100;
assign v_72102 = v_72095 & v_72101;
assign v_72103 = v_72102;
assign v_72104 = v_40066;
assign v_72105 = v_39830 & v_72104;
assign v_72106 = v_39979;
assign v_72107 = ~v_39830 & v_72106;
assign v_72109 = v_72108;
assign v_72110 = v_72103 & v_72109;
assign v_72111 = v_72110;
assign v_72112 = v_40309;
assign v_72113 = v_40073 & v_72112;
assign v_72114 = v_40222;
assign v_72115 = ~v_40073 & v_72114;
assign v_72117 = v_72116;
assign v_72118 = v_72111 & v_72117;
assign v_72119 = v_72118;
assign v_72120 = v_40552;
assign v_72121 = v_40316 & v_72120;
assign v_72122 = v_40465;
assign v_72123 = ~v_40316 & v_72122;
assign v_72125 = v_72124;
assign v_72126 = v_72119 & v_72125;
assign v_72127 = v_72126;
assign v_72128 = v_40795;
assign v_72129 = v_40559 & v_72128;
assign v_72130 = v_40708;
assign v_72131 = ~v_40559 & v_72130;
assign v_72133 = v_72132;
assign v_72134 = v_72127 & v_72133;
assign v_72135 = v_72134;
assign v_72136 = v_41038;
assign v_72137 = v_40802 & v_72136;
assign v_72138 = v_40951;
assign v_72139 = ~v_40802 & v_72138;
assign v_72141 = v_72140;
assign v_72142 = v_72135 & v_72141;
assign v_72143 = v_72142;
assign v_72144 = v_41281;
assign v_72145 = v_41045 & v_72144;
assign v_72146 = v_41194;
assign v_72147 = ~v_41045 & v_72146;
assign v_72149 = v_72148;
assign v_72150 = v_72143 & v_72149;
assign v_72151 = v_72150;
assign v_72152 = v_41524;
assign v_72153 = v_41288 & v_72152;
assign v_72154 = v_41437;
assign v_72155 = ~v_41288 & v_72154;
assign v_72157 = v_72156;
assign v_72158 = v_72151 & v_72157;
assign v_72159 = v_72158;
assign v_72160 = v_41680;
assign v_72161 = v_41767 & v_72160;
assign v_72162 = ~v_41680;
assign v_72163 = v_41679 & v_72162;
assign v_72165 = v_72164;
assign v_72166 = v_72159 & v_72165;
assign v_72167 = v_72166;
assign v_72168 = v_42027;
assign v_72169 = v_41774 & v_72168;
assign v_72170 = v_41940;
assign v_72171 = ~v_41774 & v_72170;
assign v_72173 = v_72172;
assign v_72174 = v_72167 & v_72173;
assign v_72175 = v_72174;
assign v_72176 = v_42270;
assign v_72177 = v_42034 & v_72176;
assign v_72178 = v_42183;
assign v_72179 = ~v_42034 & v_72178;
assign v_72181 = v_72180;
assign v_72182 = v_72175 & v_72181;
assign v_72183 = v_72182;
assign v_72184 = v_42513;
assign v_72185 = v_42277 & v_72184;
assign v_72186 = v_42426;
assign v_72187 = ~v_42277 & v_72186;
assign v_72189 = v_72188;
assign v_72190 = v_72183 & v_72189;
assign v_72191 = v_72190;
assign v_72192 = v_42756;
assign v_72193 = v_42520 & v_72192;
assign v_72194 = v_42669;
assign v_72195 = ~v_42520 & v_72194;
assign v_72197 = v_72196;
assign v_72198 = v_72191 & v_72197;
assign v_72199 = v_72198;
assign v_72200 = v_42999;
assign v_72201 = v_42763 & v_72200;
assign v_72202 = v_42912;
assign v_72203 = ~v_42763 & v_72202;
assign v_72205 = v_72204;
assign v_72206 = v_72199 & v_72205;
assign v_72207 = v_72206;
assign v_72208 = v_43242;
assign v_72209 = v_43006 & v_72208;
assign v_72210 = v_43155;
assign v_72211 = ~v_43006 & v_72210;
assign v_72213 = v_72212;
assign v_72214 = v_72207 & v_72213;
assign v_72215 = v_72214;
assign v_72216 = v_43485;
assign v_72217 = v_43249 & v_72216;
assign v_72218 = v_43398;
assign v_72219 = ~v_43249 & v_72218;
assign v_72221 = v_72220;
assign v_72222 = v_72215 & v_72221;
assign v_72223 = v_72222;
assign v_72224 = v_43728;
assign v_72225 = v_43492 & v_72224;
assign v_72226 = v_43641;
assign v_72227 = ~v_43492 & v_72226;
assign v_72229 = v_72228;
assign v_72230 = v_72223 & v_72229;
assign v_72231 = v_72230;
assign v_72232 = v_43971;
assign v_72233 = v_43735 & v_72232;
assign v_72234 = v_43884;
assign v_72235 = ~v_43735 & v_72234;
assign v_72237 = v_72236;
assign v_72238 = v_72231 & v_72237;
assign v_72239 = v_72238;
assign v_72240 = v_44214;
assign v_72241 = v_43978 & v_72240;
assign v_72242 = v_44127;
assign v_72243 = ~v_43978 & v_72242;
assign v_72245 = v_72244;
assign v_72246 = v_72239 & v_72245;
assign v_72247 = v_72246;
assign v_72248 = v_44457;
assign v_72249 = v_44221 & v_72248;
assign v_72250 = v_44370;
assign v_72251 = ~v_44221 & v_72250;
assign v_72253 = v_72252;
assign v_72254 = v_72247 & v_72253;
assign v_72255 = v_72254;
assign v_72256 = v_44700;
assign v_72257 = v_44464 & v_72256;
assign v_72258 = v_44613;
assign v_72259 = ~v_44464 & v_72258;
assign v_72261 = v_72260;
assign v_72262 = v_72255 & v_72261;
assign v_72263 = v_72262;
assign v_72264 = v_44943;
assign v_72265 = v_44707 & v_72264;
assign v_72266 = v_44856;
assign v_72267 = ~v_44707 & v_72266;
assign v_72269 = v_72268;
assign v_72270 = v_72263 & v_72269;
assign v_72271 = v_72270;
assign v_72272 = v_45186;
assign v_72273 = v_44950 & v_72272;
assign v_72274 = v_45099;
assign v_72275 = ~v_44950 & v_72274;
assign v_72277 = v_72276;
assign v_72278 = v_72271 & v_72277;
assign v_72279 = v_72278;
assign v_72280 = v_45429;
assign v_72281 = v_45193 & v_72280;
assign v_72282 = v_45342;
assign v_72283 = ~v_45193 & v_72282;
assign v_72285 = v_72284;
assign v_72286 = v_72279 & v_72285;
assign v_72287 = v_72286;
assign v_72288 = v_45672;
assign v_72289 = v_45436 & v_72288;
assign v_72290 = v_45585;
assign v_72291 = ~v_45436 & v_72290;
assign v_72293 = v_72292;
assign v_72294 = v_72287 & v_72293;
assign v_72295 = v_72294;
assign v_72296 = v_45828;
assign v_72297 = v_45915 & v_72296;
assign v_72298 = ~v_45828;
assign v_72299 = v_45827 & v_72298;
assign v_72301 = v_72300;
assign v_72302 = v_72295 & v_72301;
assign v_72303 = v_72302;
assign v_72304 = v_46175;
assign v_72305 = v_45922 & v_72304;
assign v_72306 = v_46088;
assign v_72307 = ~v_45922 & v_72306;
assign v_72309 = v_72308;
assign v_72310 = v_72303 & v_72309;
assign v_72311 = v_72310;
assign v_72312 = v_46418;
assign v_72313 = v_46182 & v_72312;
assign v_72314 = v_46331;
assign v_72315 = ~v_46182 & v_72314;
assign v_72317 = v_72316;
assign v_72318 = v_72311 & v_72317;
assign v_72319 = v_72318;
assign v_72320 = v_46661;
assign v_72321 = v_46425 & v_72320;
assign v_72322 = v_46574;
assign v_72323 = ~v_46425 & v_72322;
assign v_72325 = v_72324;
assign v_72326 = v_72319 & v_72325;
assign v_72327 = v_72326;
assign v_72328 = v_46904;
assign v_72329 = v_46668 & v_72328;
assign v_72330 = v_46817;
assign v_72331 = ~v_46668 & v_72330;
assign v_72333 = v_72332;
assign v_72334 = v_72327 & v_72333;
assign v_72335 = v_72334;
assign v_72336 = v_47147;
assign v_72337 = v_46911 & v_72336;
assign v_72338 = v_47060;
assign v_72339 = ~v_46911 & v_72338;
assign v_72341 = v_72340;
assign v_72342 = v_72335 & v_72341;
assign v_72343 = v_72342;
assign v_72344 = v_47390;
assign v_72345 = v_47154 & v_72344;
assign v_72346 = v_47303;
assign v_72347 = ~v_47154 & v_72346;
assign v_72349 = v_72348;
assign v_72350 = v_72343 & v_72349;
assign v_72351 = v_72350;
assign v_72352 = v_47633;
assign v_72353 = v_47397 & v_72352;
assign v_72354 = v_47546;
assign v_72355 = ~v_47397 & v_72354;
assign v_72357 = v_72356;
assign v_72358 = v_72351 & v_72357;
assign v_72359 = v_72358;
assign v_72360 = v_47876;
assign v_72361 = v_47640 & v_72360;
assign v_72362 = v_47789;
assign v_72363 = ~v_47640 & v_72362;
assign v_72365 = v_72364;
assign v_72366 = v_72359 & v_72365;
assign v_72367 = v_72366;
assign v_72368 = v_48119;
assign v_72369 = v_47883 & v_72368;
assign v_72370 = v_48032;
assign v_72371 = ~v_47883 & v_72370;
assign v_72373 = v_72372;
assign v_72374 = v_72367 & v_72373;
assign v_72375 = v_72374;
assign v_72376 = v_48362;
assign v_72377 = v_48126 & v_72376;
assign v_72378 = v_48275;
assign v_72379 = ~v_48126 & v_72378;
assign v_72381 = v_72380;
assign v_72382 = v_72375 & v_72381;
assign v_72383 = v_72382;
assign v_72384 = v_48605;
assign v_72385 = v_48369 & v_72384;
assign v_72386 = v_48518;
assign v_72387 = ~v_48369 & v_72386;
assign v_72389 = v_72388;
assign v_72390 = v_72383 & v_72389;
assign v_72391 = v_72390;
assign v_72392 = v_48848;
assign v_72393 = v_48612 & v_72392;
assign v_72394 = v_48761;
assign v_72395 = ~v_48612 & v_72394;
assign v_72397 = v_72396;
assign v_72398 = v_72391 & v_72397;
assign v_72399 = v_72398;
assign v_72400 = v_49091;
assign v_72401 = v_48855 & v_72400;
assign v_72402 = v_49004;
assign v_72403 = ~v_48855 & v_72402;
assign v_72405 = v_72404;
assign v_72406 = v_72399 & v_72405;
assign v_72407 = v_72406;
assign v_72408 = v_49334;
assign v_72409 = v_49098 & v_72408;
assign v_72410 = v_49247;
assign v_72411 = ~v_49098 & v_72410;
assign v_72413 = v_72412;
assign v_72414 = v_72407 & v_72413;
assign v_72415 = v_72414;
assign v_72416 = v_49577;
assign v_72417 = v_49341 & v_72416;
assign v_72418 = v_49490;
assign v_72419 = ~v_49341 & v_72418;
assign v_72421 = v_72420;
assign v_72422 = v_72415 & v_72421;
assign v_72423 = v_72422;
assign v_72424 = v_49820;
assign v_72425 = v_49584 & v_72424;
assign v_72426 = v_49733;
assign v_72427 = ~v_49584 & v_72426;
assign v_72429 = v_72428;
assign v_72430 = v_72423 & v_72429;
assign v_72431 = v_72430;
assign v_72432 = v_49976;
assign v_72433 = v_50063 & v_72432;
assign v_72434 = ~v_49976;
assign v_72435 = v_49975 & v_72434;
assign v_72437 = v_72436;
assign v_72438 = v_72431 & v_72437;
assign v_72439 = v_72438;
assign v_72440 = v_50323;
assign v_72441 = v_50070 & v_72440;
assign v_72442 = v_50236;
assign v_72443 = ~v_50070 & v_72442;
assign v_72445 = v_72444;
assign v_72446 = v_72439 & v_72445;
assign v_72447 = v_72446;
assign v_72448 = v_50566;
assign v_72449 = v_50330 & v_72448;
assign v_72450 = v_50479;
assign v_72451 = ~v_50330 & v_72450;
assign v_72453 = v_72452;
assign v_72454 = v_72447 & v_72453;
assign v_72455 = v_72454;
assign v_72456 = v_50809;
assign v_72457 = v_50573 & v_72456;
assign v_72458 = v_50722;
assign v_72459 = ~v_50573 & v_72458;
assign v_72461 = v_72460;
assign v_72462 = v_72455 & v_72461;
assign v_72463 = v_72462;
assign v_72464 = v_51052;
assign v_72465 = v_50816 & v_72464;
assign v_72466 = v_50965;
assign v_72467 = ~v_50816 & v_72466;
assign v_72469 = v_72468;
assign v_72470 = v_72463 & v_72469;
assign v_72471 = v_72470;
assign v_72472 = v_51295;
assign v_72473 = v_51059 & v_72472;
assign v_72474 = v_51208;
assign v_72475 = ~v_51059 & v_72474;
assign v_72477 = v_72476;
assign v_72478 = v_72471 & v_72477;
assign v_72479 = v_72478;
assign v_72480 = v_51538;
assign v_72481 = v_51302 & v_72480;
assign v_72482 = v_51451;
assign v_72483 = ~v_51302 & v_72482;
assign v_72485 = v_72484;
assign v_72486 = v_72479 & v_72485;
assign v_72487 = v_72486;
assign v_72488 = v_51781;
assign v_72489 = v_51545 & v_72488;
assign v_72490 = v_51694;
assign v_72491 = ~v_51545 & v_72490;
assign v_72493 = v_72492;
assign v_72494 = v_72487 & v_72493;
assign v_72495 = v_72494;
assign v_72496 = v_52024;
assign v_72497 = v_51788 & v_72496;
assign v_72498 = v_51937;
assign v_72499 = ~v_51788 & v_72498;
assign v_72501 = v_72500;
assign v_72502 = v_72495 & v_72501;
assign v_72503 = v_72502;
assign v_72504 = v_52267;
assign v_72505 = v_52031 & v_72504;
assign v_72506 = v_52180;
assign v_72507 = ~v_52031 & v_72506;
assign v_72509 = v_72508;
assign v_72510 = v_72503 & v_72509;
assign v_72511 = v_72510;
assign v_72512 = v_52510;
assign v_72513 = v_52274 & v_72512;
assign v_72514 = v_52423;
assign v_72515 = ~v_52274 & v_72514;
assign v_72517 = v_72516;
assign v_72518 = v_72511 & v_72517;
assign v_72519 = v_72518;
assign v_72520 = v_52753;
assign v_72521 = v_52517 & v_72520;
assign v_72522 = v_52666;
assign v_72523 = ~v_52517 & v_72522;
assign v_72525 = v_72524;
assign v_72526 = v_72519 & v_72525;
assign v_72527 = v_72526;
assign v_72528 = v_52996;
assign v_72529 = v_52760 & v_72528;
assign v_72530 = v_52909;
assign v_72531 = ~v_52760 & v_72530;
assign v_72533 = v_72532;
assign v_72534 = v_72527 & v_72533;
assign v_72535 = v_72534;
assign v_72536 = v_53239;
assign v_72537 = v_53003 & v_72536;
assign v_72538 = v_53152;
assign v_72539 = ~v_53003 & v_72538;
assign v_72541 = v_72540;
assign v_72542 = v_72535 & v_72541;
assign v_72543 = v_72542;
assign v_72544 = v_53482;
assign v_72545 = v_53246 & v_72544;
assign v_72546 = v_53395;
assign v_72547 = ~v_53246 & v_72546;
assign v_72549 = v_72548;
assign v_72550 = v_72543 & v_72549;
assign v_72551 = v_72550;
assign v_72552 = v_53725;
assign v_72553 = v_53489 & v_72552;
assign v_72554 = v_53638;
assign v_72555 = ~v_53489 & v_72554;
assign v_72557 = v_72556;
assign v_72558 = v_72551 & v_72557;
assign v_72559 = v_72558;
assign v_72560 = v_53968;
assign v_72561 = v_53732 & v_72560;
assign v_72562 = v_53881;
assign v_72563 = ~v_53732 & v_72562;
assign v_72565 = v_72564;
assign v_72566 = v_72559 & v_72565;
assign v_72567 = v_72566;
assign v_72568 = v_54124;
assign v_72569 = v_54211 & v_72568;
assign v_72570 = ~v_54124;
assign v_72571 = v_54123 & v_72570;
assign v_72573 = v_72572;
assign v_72574 = v_72567 & v_72573;
assign v_72575 = v_72574;
assign v_72576 = v_54471;
assign v_72577 = v_54218 & v_72576;
assign v_72578 = v_54384;
assign v_72579 = ~v_54218 & v_72578;
assign v_72581 = v_72580;
assign v_72582 = v_72575 & v_72581;
assign v_72583 = v_72582;
assign v_72584 = v_54714;
assign v_72585 = v_54478 & v_72584;
assign v_72586 = v_54627;
assign v_72587 = ~v_54478 & v_72586;
assign v_72589 = v_72588;
assign v_72590 = v_72583 & v_72589;
assign v_72591 = v_72590;
assign v_72592 = v_54957;
assign v_72593 = v_54721 & v_72592;
assign v_72594 = v_54870;
assign v_72595 = ~v_54721 & v_72594;
assign v_72597 = v_72596;
assign v_72598 = v_72591 & v_72597;
assign v_72599 = v_72598;
assign v_72600 = v_55200;
assign v_72601 = v_54964 & v_72600;
assign v_72602 = v_55113;
assign v_72603 = ~v_54964 & v_72602;
assign v_72605 = v_72604;
assign v_72606 = v_72599 & v_72605;
assign v_72607 = v_72606;
assign v_72608 = v_55443;
assign v_72609 = v_55207 & v_72608;
assign v_72610 = v_55356;
assign v_72611 = ~v_55207 & v_72610;
assign v_72613 = v_72612;
assign v_72614 = v_72607 & v_72613;
assign v_72615 = v_72614;
assign v_72616 = v_55686;
assign v_72617 = v_55450 & v_72616;
assign v_72618 = v_55599;
assign v_72619 = ~v_55450 & v_72618;
assign v_72621 = v_72620;
assign v_72622 = v_72615 & v_72621;
assign v_72623 = v_72622;
assign v_72624 = v_55929;
assign v_72625 = v_55693 & v_72624;
assign v_72626 = v_55842;
assign v_72627 = ~v_55693 & v_72626;
assign v_72629 = v_72628;
assign v_72630 = v_72623 & v_72629;
assign v_72631 = v_72630;
assign v_72632 = v_56172;
assign v_72633 = v_55936 & v_72632;
assign v_72634 = v_56085;
assign v_72635 = ~v_55936 & v_72634;
assign v_72637 = v_72636;
assign v_72638 = v_72631 & v_72637;
assign v_72639 = v_72638;
assign v_72640 = v_56415;
assign v_72641 = v_56179 & v_72640;
assign v_72642 = v_56328;
assign v_72643 = ~v_56179 & v_72642;
assign v_72645 = v_72644;
assign v_72646 = v_72639 & v_72645;
assign v_72647 = v_72646;
assign v_72648 = v_56658;
assign v_72649 = v_56422 & v_72648;
assign v_72650 = v_56571;
assign v_72651 = ~v_56422 & v_72650;
assign v_72653 = v_72652;
assign v_72654 = v_72647 & v_72653;
assign v_72655 = v_72654;
assign v_72656 = v_56901;
assign v_72657 = v_56665 & v_72656;
assign v_72658 = v_56814;
assign v_72659 = ~v_56665 & v_72658;
assign v_72661 = v_72660;
assign v_72662 = v_72655 & v_72661;
assign v_72663 = v_72662;
assign v_72664 = v_57144;
assign v_72665 = v_56908 & v_72664;
assign v_72666 = v_57057;
assign v_72667 = ~v_56908 & v_72666;
assign v_72669 = v_72668;
assign v_72670 = v_72663 & v_72669;
assign v_72671 = v_72670;
assign v_72672 = v_57387;
assign v_72673 = v_57151 & v_72672;
assign v_72674 = v_57300;
assign v_72675 = ~v_57151 & v_72674;
assign v_72677 = v_72676;
assign v_72678 = v_72671 & v_72677;
assign v_72679 = v_72678;
assign v_72680 = v_57630;
assign v_72681 = v_57394 & v_72680;
assign v_72682 = v_57543;
assign v_72683 = ~v_57394 & v_72682;
assign v_72685 = v_72684;
assign v_72686 = v_72679 & v_72685;
assign v_72687 = v_72686;
assign v_72688 = v_57873;
assign v_72689 = v_57637 & v_72688;
assign v_72690 = v_57786;
assign v_72691 = ~v_57637 & v_72690;
assign v_72693 = v_72692;
assign v_72694 = v_72687 & v_72693;
assign v_72695 = v_72694;
assign v_72696 = v_58116;
assign v_72697 = v_57880 & v_72696;
assign v_72698 = v_58029;
assign v_72699 = ~v_57880 & v_72698;
assign v_72701 = v_72700;
assign v_72702 = v_72695 & v_72701;
assign v_72703 = v_72702;
assign v_72704 = v_58272;
assign v_72705 = v_58359 & v_72704;
assign v_72706 = ~v_58272;
assign v_72707 = v_58271 & v_72706;
assign v_72709 = v_72708;
assign v_72710 = v_72703 & v_72709;
assign v_72711 = v_72710;
assign v_72712 = v_58619;
assign v_72713 = v_58366 & v_72712;
assign v_72714 = v_58532;
assign v_72715 = ~v_58366 & v_72714;
assign v_72717 = v_72716;
assign v_72718 = v_72711 & v_72717;
assign v_72719 = v_72718;
assign v_72720 = v_58862;
assign v_72721 = v_58626 & v_72720;
assign v_72722 = v_58775;
assign v_72723 = ~v_58626 & v_72722;
assign v_72725 = v_72724;
assign v_72726 = v_72719 & v_72725;
assign v_72727 = v_72726;
assign v_72728 = v_59105;
assign v_72729 = v_58869 & v_72728;
assign v_72730 = v_59018;
assign v_72731 = ~v_58869 & v_72730;
assign v_72733 = v_72732;
assign v_72734 = v_72727 & v_72733;
assign v_72735 = v_72734;
assign v_72736 = v_59348;
assign v_72737 = v_59112 & v_72736;
assign v_72738 = v_59261;
assign v_72739 = ~v_59112 & v_72738;
assign v_72741 = v_72740;
assign v_72742 = v_72735 & v_72741;
assign v_72743 = v_72742;
assign v_72744 = v_59591;
assign v_72745 = v_59355 & v_72744;
assign v_72746 = v_59504;
assign v_72747 = ~v_59355 & v_72746;
assign v_72749 = v_72748;
assign v_72750 = v_72743 & v_72749;
assign v_72751 = v_72750;
assign v_72752 = v_59834;
assign v_72753 = v_59598 & v_72752;
assign v_72754 = v_59747;
assign v_72755 = ~v_59598 & v_72754;
assign v_72757 = v_72756;
assign v_72758 = v_72751 & v_72757;
assign v_72759 = v_72758;
assign v_72760 = v_60077;
assign v_72761 = v_59841 & v_72760;
assign v_72762 = v_59990;
assign v_72763 = ~v_59841 & v_72762;
assign v_72765 = v_72764;
assign v_72766 = v_72759 & v_72765;
assign v_72767 = v_72766;
assign v_72768 = v_60320;
assign v_72769 = v_60084 & v_72768;
assign v_72770 = v_60233;
assign v_72771 = ~v_60084 & v_72770;
assign v_72773 = v_72772;
assign v_72774 = v_72767 & v_72773;
assign v_72775 = v_72774;
assign v_72776 = v_60563;
assign v_72777 = v_60327 & v_72776;
assign v_72778 = v_60476;
assign v_72779 = ~v_60327 & v_72778;
assign v_72781 = v_72780;
assign v_72782 = v_72775 & v_72781;
assign v_72783 = v_72782;
assign v_72784 = v_60806;
assign v_72785 = v_60570 & v_72784;
assign v_72786 = v_60719;
assign v_72787 = ~v_60570 & v_72786;
assign v_72789 = v_72788;
assign v_72790 = v_72783 & v_72789;
assign v_72791 = v_72790;
assign v_72792 = v_61049;
assign v_72793 = v_60813 & v_72792;
assign v_72794 = v_60962;
assign v_72795 = ~v_60813 & v_72794;
assign v_72797 = v_72796;
assign v_72798 = v_72791 & v_72797;
assign v_72799 = v_72798;
assign v_72800 = v_61292;
assign v_72801 = v_61056 & v_72800;
assign v_72802 = v_61205;
assign v_72803 = ~v_61056 & v_72802;
assign v_72805 = v_72804;
assign v_72806 = v_72799 & v_72805;
assign v_72807 = v_72806;
assign v_72808 = v_61535;
assign v_72809 = v_61299 & v_72808;
assign v_72810 = v_61448;
assign v_72811 = ~v_61299 & v_72810;
assign v_72813 = v_72812;
assign v_72814 = v_72807 & v_72813;
assign v_72815 = v_72814;
assign v_72816 = v_61778;
assign v_72817 = v_61542 & v_72816;
assign v_72818 = v_61691;
assign v_72819 = ~v_61542 & v_72818;
assign v_72821 = v_72820;
assign v_72822 = v_72815 & v_72821;
assign v_72823 = v_72822;
assign v_72824 = v_62021;
assign v_72825 = v_61785 & v_72824;
assign v_72826 = v_61934;
assign v_72827 = ~v_61785 & v_72826;
assign v_72829 = v_72828;
assign v_72830 = v_72823 & v_72829;
assign v_72831 = v_72830;
assign v_72832 = v_62264;
assign v_72833 = v_62028 & v_72832;
assign v_72834 = v_62177;
assign v_72835 = ~v_62028 & v_72834;
assign v_72837 = v_72836;
assign v_72838 = v_72831 & v_72837;
assign v_72839 = v_72838;
assign v_72840 = v_62420;
assign v_72841 = v_62507 & v_72840;
assign v_72842 = ~v_62420;
assign v_72843 = v_62419 & v_72842;
assign v_72845 = v_72844;
assign v_72846 = v_72839 & v_72845;
assign v_72847 = v_72846;
assign v_72848 = v_62767;
assign v_72849 = v_62514 & v_72848;
assign v_72850 = v_62680;
assign v_72851 = ~v_62514 & v_72850;
assign v_72853 = v_72852;
assign v_72854 = v_72847 & v_72853;
assign v_72855 = v_72854;
assign v_72856 = v_63010;
assign v_72857 = v_62774 & v_72856;
assign v_72858 = v_62923;
assign v_72859 = ~v_62774 & v_72858;
assign v_72861 = v_72860;
assign v_72862 = v_72855 & v_72861;
assign v_72863 = v_72862;
assign v_72864 = v_63253;
assign v_72865 = v_63017 & v_72864;
assign v_72866 = v_63166;
assign v_72867 = ~v_63017 & v_72866;
assign v_72869 = v_72868;
assign v_72870 = v_72863 & v_72869;
assign v_72871 = v_72870;
assign v_72872 = v_63496;
assign v_72873 = v_63260 & v_72872;
assign v_72874 = v_63409;
assign v_72875 = ~v_63260 & v_72874;
assign v_72877 = v_72876;
assign v_72878 = v_72871 & v_72877;
assign v_72879 = v_72878;
assign v_72880 = v_63739;
assign v_72881 = v_63503 & v_72880;
assign v_72882 = v_63652;
assign v_72883 = ~v_63503 & v_72882;
assign v_72885 = v_72884;
assign v_72886 = v_72879 & v_72885;
assign v_72887 = v_72886;
assign v_72888 = v_63982;
assign v_72889 = v_63746 & v_72888;
assign v_72890 = v_63895;
assign v_72891 = ~v_63746 & v_72890;
assign v_72893 = v_72892;
assign v_72894 = v_72887 & v_72893;
assign v_72895 = v_72894;
assign v_72896 = v_64225;
assign v_72897 = v_63989 & v_72896;
assign v_72898 = v_64138;
assign v_72899 = ~v_63989 & v_72898;
assign v_72901 = v_72900;
assign v_72902 = v_72895 & v_72901;
assign v_72903 = v_72902;
assign v_72904 = v_64468;
assign v_72905 = v_64232 & v_72904;
assign v_72906 = v_64381;
assign v_72907 = ~v_64232 & v_72906;
assign v_72909 = v_72908;
assign v_72910 = v_72903 & v_72909;
assign v_72911 = v_72910;
assign v_72912 = v_64711;
assign v_72913 = v_64475 & v_72912;
assign v_72914 = v_64624;
assign v_72915 = ~v_64475 & v_72914;
assign v_72917 = v_72916;
assign v_72918 = v_72911 & v_72917;
assign v_72919 = v_72918;
assign v_72920 = v_64954;
assign v_72921 = v_64718 & v_72920;
assign v_72922 = v_64867;
assign v_72923 = ~v_64718 & v_72922;
assign v_72925 = v_72924;
assign v_72926 = v_72919 & v_72925;
assign v_72927 = v_72926;
assign v_72928 = v_65197;
assign v_72929 = v_64961 & v_72928;
assign v_72930 = v_65110;
assign v_72931 = ~v_64961 & v_72930;
assign v_72933 = v_72932;
assign v_72934 = v_72927 & v_72933;
assign v_72935 = v_72934;
assign v_72936 = v_65440;
assign v_72937 = v_65204 & v_72936;
assign v_72938 = v_65353;
assign v_72939 = ~v_65204 & v_72938;
assign v_72941 = v_72940;
assign v_72942 = v_72935 & v_72941;
assign v_72943 = v_72942;
assign v_72944 = v_65683;
assign v_72945 = v_65447 & v_72944;
assign v_72946 = v_65596;
assign v_72947 = ~v_65447 & v_72946;
assign v_72949 = v_72948;
assign v_72950 = v_72943 & v_72949;
assign v_72951 = v_72950;
assign v_72952 = v_65926;
assign v_72953 = v_65690 & v_72952;
assign v_72954 = v_65839;
assign v_72955 = ~v_65690 & v_72954;
assign v_72957 = v_72956;
assign v_72958 = v_72951 & v_72957;
assign v_72959 = v_72958;
assign v_72960 = v_66169;
assign v_72961 = v_65933 & v_72960;
assign v_72962 = v_66082;
assign v_72963 = ~v_65933 & v_72962;
assign v_72965 = v_72964;
assign v_72966 = v_72959 & v_72965;
assign v_72967 = v_72966;
assign v_72968 = v_66412;
assign v_72969 = v_66176 & v_72968;
assign v_72970 = v_66325;
assign v_72971 = ~v_66176 & v_72970;
assign v_72973 = v_72972;
assign v_72974 = v_72967 & v_72973;
assign v_72975 = v_72974;
assign v_72976 = v_66568;
assign v_72977 = v_66655 & v_72976;
assign v_72978 = ~v_66568;
assign v_72979 = v_66567 & v_72978;
assign v_72981 = v_72980;
assign v_72982 = v_72975 & v_72981;
assign v_72983 = v_72982;
assign v_72984 = v_66828;
assign v_72985 = v_66915 & v_72984;
assign v_72986 = ~v_66828;
assign v_72987 = v_66827 & v_72986;
assign v_72989 = v_72988;
assign v_72990 = v_72983 & v_72989;
assign v_72991 = v_72990;
assign v_72992 = v_67071;
assign v_72993 = v_67158 & v_72992;
assign v_72994 = ~v_67071;
assign v_72995 = v_67070 & v_72994;
assign v_72997 = v_72996;
assign v_72998 = v_72991 & v_72997;
assign v_72999 = v_72998;
assign v_73000 = v_67314;
assign v_73001 = v_67401 & v_73000;
assign v_73002 = ~v_67314;
assign v_73003 = v_67313 & v_73002;
assign v_73005 = v_73004;
assign v_73006 = v_72999 & v_73005;
assign v_73007 = v_73006;
assign v_73008 = v_67557;
assign v_73009 = v_67644 & v_73008;
assign v_73010 = ~v_67557;
assign v_73011 = v_67556 & v_73010;
assign v_73013 = v_73012;
assign v_73014 = v_73007 & v_73013;
assign v_73015 = v_73014;
assign v_73016 = v_67800;
assign v_73017 = v_67887 & v_73016;
assign v_73018 = ~v_67800;
assign v_73019 = v_67799 & v_73018;
assign v_73021 = v_73020;
assign v_73022 = v_73015 & v_73021;
assign v_73023 = v_73022;
assign v_73024 = v_68043;
assign v_73025 = v_68130 & v_73024;
assign v_73026 = ~v_68043;
assign v_73027 = v_68042 & v_73026;
assign v_73029 = v_73028;
assign v_73030 = v_73023 & v_73029;
assign v_73031 = v_73030;
assign v_73032 = v_68286;
assign v_73033 = v_68373 & v_73032;
assign v_73034 = ~v_68286;
assign v_73035 = v_68285 & v_73034;
assign v_73037 = v_73036;
assign v_73038 = v_73031 & v_73037;
assign v_73039 = v_73038;
assign v_73040 = v_68529;
assign v_73041 = v_68616 & v_73040;
assign v_73042 = ~v_68529;
assign v_73043 = v_68528 & v_73042;
assign v_73045 = v_73044;
assign v_73046 = v_73039 & v_73045;
assign v_73047 = v_73046;
assign v_73048 = v_68772;
assign v_73049 = v_68859 & v_73048;
assign v_73050 = ~v_68772;
assign v_73051 = v_68771 & v_73050;
assign v_73053 = v_73052;
assign v_73054 = v_73047 & v_73053;
assign v_73055 = v_73054;
assign v_73056 = v_69015;
assign v_73057 = v_69102 & v_73056;
assign v_73058 = ~v_69015;
assign v_73059 = v_69014 & v_73058;
assign v_73061 = v_73060;
assign v_73062 = v_73055 & v_73061;
assign v_73063 = v_73062;
assign v_73064 = v_69258;
assign v_73065 = v_69345 & v_73064;
assign v_73066 = ~v_69258;
assign v_73067 = v_69257 & v_73066;
assign v_73069 = v_73068;
assign v_73070 = v_73063 & v_73069;
assign v_73071 = v_73070;
assign v_73072 = v_69501;
assign v_73073 = v_69588 & v_73072;
assign v_73074 = ~v_69501;
assign v_73075 = v_69500 & v_73074;
assign v_73077 = v_73076;
assign v_73078 = v_73071 & v_73077;
assign v_73079 = v_73078;
assign v_73080 = v_69744;
assign v_73081 = v_69831 & v_73080;
assign v_73082 = ~v_69744;
assign v_73083 = v_69743 & v_73082;
assign v_73085 = v_73084;
assign v_73086 = v_73079 & v_73085;
assign v_73087 = v_73086;
assign v_73088 = v_69987;
assign v_73089 = v_70074 & v_73088;
assign v_73090 = ~v_69987;
assign v_73091 = v_69986 & v_73090;
assign v_73093 = v_73092;
assign v_73094 = v_73087 & v_73093;
assign v_73095 = v_73094;
assign v_73096 = v_70230;
assign v_73097 = v_70317 & v_73096;
assign v_73098 = ~v_70230;
assign v_73099 = v_70229 & v_73098;
assign v_73101 = v_73100;
assign v_73102 = v_73095 & v_73101;
assign v_73103 = v_73102;
assign v_73104 = v_70473;
assign v_73105 = v_70560 & v_73104;
assign v_73106 = ~v_70473;
assign v_73107 = v_70472 & v_73106;
assign v_73109 = v_73108;
assign v_73110 = v_73103 & v_73109;
assign v_73111 = v_73110;
assign v_73112 = v_70716;
assign v_73113 = v_70803 & v_73112;
assign v_73114 = ~v_70716;
assign v_73115 = v_70715 & v_73114;
assign v_73117 = v_73116;
assign v_73118 = v_73111 & v_73117;
assign v_73120 = ~v_4;
assign v_73121 = v_73120;
assign v_73122 = v_70809 & v_73119 & v_73121;
assign v_93 = v_89 | v_92;
assign v_95 = v_87 | v_94;
assign v_97 = v_84 | v_96;
assign v_99 = v_94 | v_98;
assign v_101 = v_82 | v_100;
assign v_103 = v_79 | v_102;
assign v_105 = v_100 | v_104;
assign v_107 = v_77 | v_106;
assign v_109 = v_74 | v_108;
assign v_111 = v_106 | v_110;
assign v_113 = v_72 | v_112;
assign v_115 = v_69 | v_114;
assign v_117 = v_112 | v_116;
assign v_119 = v_67 | v_118;
assign v_121 = v_64 | v_120;
assign v_123 = v_118 | v_122;
assign v_125 = v_62 | v_124;
assign v_127 = v_59 | v_126;
assign v_129 = v_124 | v_128;
assign v_131 = v_57 | v_130;
assign v_133 = v_54 | v_132;
assign v_135 = v_130 | v_134;
assign v_137 = v_52 | v_136;
assign v_139 = v_49 | v_138;
assign v_141 = v_136 | v_140;
assign v_143 = v_47 | v_142;
assign v_145 = v_44 | v_144;
assign v_147 = v_142 | v_146;
assign v_149 = v_42 | v_148;
assign v_151 = v_39 | v_150;
assign v_153 = v_148 | v_152;
assign v_155 = v_37 | v_154;
assign v_157 = v_34 | v_156;
assign v_159 = v_154 | v_158;
assign v_161 = v_32 | v_160;
assign v_163 = v_29 | v_162;
assign v_165 = v_160 | v_164;
assign v_167 = v_27 | v_166;
assign v_169 = v_24 | v_168;
assign v_171 = v_166 | v_170;
assign v_173 = v_22 | v_172;
assign v_175 = v_19 | v_174;
assign v_177 = v_172 | v_176;
assign v_179 = v_17 | v_178;
assign v_181 = v_14 | v_180;
assign v_183 = v_178 | v_182;
assign v_185 = v_12 | v_184;
assign v_187 = v_8 | v_186;
assign v_189 = v_184 | v_188;
assign v_192 = ~v_5 | v_191;
assign v_199 = v_87 | v_198;
assign v_202 = v_200 | v_201;
assign v_204 = v_82 | v_203;
assign v_207 = v_205 | v_206;
assign v_209 = v_77 | v_208;
assign v_212 = v_210 | v_211;
assign v_214 = v_72 | v_213;
assign v_217 = v_215 | v_216;
assign v_219 = v_67 | v_218;
assign v_222 = v_220 | v_221;
assign v_224 = v_62 | v_223;
assign v_227 = v_225 | v_226;
assign v_229 = v_57 | v_228;
assign v_232 = v_230 | v_231;
assign v_234 = v_52 | v_233;
assign v_237 = v_235 | v_236;
assign v_239 = v_47 | v_238;
assign v_242 = v_240 | v_241;
assign v_244 = v_42 | v_243;
assign v_247 = v_245 | v_246;
assign v_249 = v_37 | v_248;
assign v_252 = v_250 | v_251;
assign v_254 = v_32 | v_253;
assign v_257 = v_255 | v_256;
assign v_259 = v_27 | v_258;
assign v_262 = v_260 | v_261;
assign v_264 = v_22 | v_263;
assign v_267 = v_265 | v_266;
assign v_269 = v_17 | v_268;
assign v_272 = v_270 | v_271;
assign v_274 = v_12 | v_273;
assign v_277 = v_275 | v_276;
assign v_279 = v_5 | v_278;
assign v_351 = v_347 | v_350;
assign v_353 = v_346 | v_352;
assign v_355 = v_343 | v_354;
assign v_357 = v_352 | v_356;
assign v_359 = v_342 | v_358;
assign v_361 = v_339 | v_360;
assign v_363 = v_358 | v_362;
assign v_365 = v_338 | v_364;
assign v_367 = v_335 | v_366;
assign v_369 = v_364 | v_368;
assign v_371 = v_334 | v_370;
assign v_373 = v_331 | v_372;
assign v_375 = v_370 | v_374;
assign v_377 = v_330 | v_376;
assign v_379 = v_327 | v_378;
assign v_381 = v_376 | v_380;
assign v_383 = v_326 | v_382;
assign v_385 = v_323 | v_384;
assign v_387 = v_382 | v_386;
assign v_389 = v_322 | v_388;
assign v_391 = v_319 | v_390;
assign v_393 = v_388 | v_392;
assign v_395 = v_318 | v_394;
assign v_397 = v_315 | v_396;
assign v_399 = v_394 | v_398;
assign v_401 = v_314 | v_400;
assign v_403 = v_311 | v_402;
assign v_405 = v_400 | v_404;
assign v_407 = v_310 | v_406;
assign v_409 = v_307 | v_408;
assign v_411 = v_406 | v_410;
assign v_413 = v_306 | v_412;
assign v_415 = v_303 | v_414;
assign v_417 = v_412 | v_416;
assign v_419 = v_302 | v_418;
assign v_421 = v_299 | v_420;
assign v_423 = v_418 | v_422;
assign v_425 = v_298 | v_424;
assign v_427 = v_296 | v_426;
assign v_429 = v_424 | v_428;
assign v_431 = v_294 | v_430;
assign v_433 = v_292 | v_432;
assign v_435 = v_430 | v_434;
assign v_437 = v_290 | v_436;
assign v_439 = v_288 | v_438;
assign v_441 = v_436 | v_440;
assign v_443 = v_286 | v_442;
assign v_445 = v_284 | v_444;
assign v_447 = v_442 | v_446;
assign v_450 = ~v_282 | v_449;
assign v_457 = v_346 | v_456;
assign v_460 = v_458 | v_459;
assign v_462 = v_342 | v_461;
assign v_465 = v_463 | v_464;
assign v_467 = v_338 | v_466;
assign v_470 = v_468 | v_469;
assign v_472 = v_334 | v_471;
assign v_475 = v_473 | v_474;
assign v_477 = v_330 | v_476;
assign v_480 = v_478 | v_479;
assign v_482 = v_326 | v_481;
assign v_485 = v_483 | v_484;
assign v_487 = v_322 | v_486;
assign v_490 = v_488 | v_489;
assign v_492 = v_318 | v_491;
assign v_495 = v_493 | v_494;
assign v_497 = v_314 | v_496;
assign v_500 = v_498 | v_499;
assign v_502 = v_310 | v_501;
assign v_505 = v_503 | v_504;
assign v_507 = v_306 | v_506;
assign v_510 = v_508 | v_509;
assign v_512 = v_302 | v_511;
assign v_515 = v_513 | v_514;
assign v_517 = v_298 | v_516;
assign v_520 = v_518 | v_519;
assign v_522 = v_294 | v_521;
assign v_525 = v_523 | v_524;
assign v_527 = v_290 | v_526;
assign v_530 = v_528 | v_529;
assign v_532 = v_286 | v_531;
assign v_535 = v_533 | v_534;
assign v_537 = v_282 | v_536;
assign v_540 = v_281 | v_539;
assign v_611 = v_607 | v_610;
assign v_613 = v_606 | v_612;
assign v_615 = v_603 | v_614;
assign v_617 = v_612 | v_616;
assign v_619 = v_602 | v_618;
assign v_621 = v_599 | v_620;
assign v_623 = v_618 | v_622;
assign v_625 = v_598 | v_624;
assign v_627 = v_595 | v_626;
assign v_629 = v_624 | v_628;
assign v_631 = v_594 | v_630;
assign v_633 = v_591 | v_632;
assign v_635 = v_630 | v_634;
assign v_637 = v_590 | v_636;
assign v_639 = v_587 | v_638;
assign v_641 = v_636 | v_640;
assign v_643 = v_586 | v_642;
assign v_645 = v_583 | v_644;
assign v_647 = v_642 | v_646;
assign v_649 = v_582 | v_648;
assign v_651 = v_579 | v_650;
assign v_653 = v_648 | v_652;
assign v_655 = v_578 | v_654;
assign v_657 = v_575 | v_656;
assign v_659 = v_654 | v_658;
assign v_661 = v_574 | v_660;
assign v_663 = v_571 | v_662;
assign v_665 = v_660 | v_664;
assign v_667 = v_570 | v_666;
assign v_669 = v_567 | v_668;
assign v_671 = v_666 | v_670;
assign v_673 = v_566 | v_672;
assign v_675 = v_563 | v_674;
assign v_677 = v_672 | v_676;
assign v_679 = v_562 | v_678;
assign v_681 = v_559 | v_680;
assign v_683 = v_678 | v_682;
assign v_685 = v_558 | v_684;
assign v_687 = v_556 | v_686;
assign v_689 = v_684 | v_688;
assign v_691 = v_554 | v_690;
assign v_693 = v_552 | v_692;
assign v_695 = v_690 | v_694;
assign v_697 = v_550 | v_696;
assign v_699 = v_548 | v_698;
assign v_701 = v_696 | v_700;
assign v_703 = v_546 | v_702;
assign v_705 = v_544 | v_704;
assign v_707 = v_702 | v_706;
assign v_710 = ~v_542 | v_709;
assign v_717 = v_606 | v_716;
assign v_720 = v_718 | v_719;
assign v_722 = v_602 | v_721;
assign v_725 = v_723 | v_724;
assign v_727 = v_598 | v_726;
assign v_730 = v_728 | v_729;
assign v_732 = v_594 | v_731;
assign v_735 = v_733 | v_734;
assign v_737 = v_590 | v_736;
assign v_740 = v_738 | v_739;
assign v_742 = v_586 | v_741;
assign v_745 = v_743 | v_744;
assign v_747 = v_582 | v_746;
assign v_750 = v_748 | v_749;
assign v_752 = v_578 | v_751;
assign v_755 = v_753 | v_754;
assign v_757 = v_574 | v_756;
assign v_760 = v_758 | v_759;
assign v_762 = v_570 | v_761;
assign v_765 = v_763 | v_764;
assign v_767 = v_566 | v_766;
assign v_770 = v_768 | v_769;
assign v_772 = v_562 | v_771;
assign v_775 = v_773 | v_774;
assign v_777 = v_558 | v_776;
assign v_780 = v_778 | v_779;
assign v_782 = v_554 | v_781;
assign v_785 = v_783 | v_784;
assign v_787 = v_550 | v_786;
assign v_790 = v_788 | v_789;
assign v_792 = v_546 | v_791;
assign v_795 = v_793 | v_794;
assign v_797 = v_542 | v_796;
assign v_800 = v_541 | v_799;
assign v_871 = v_867 | v_870;
assign v_873 = v_866 | v_872;
assign v_875 = v_863 | v_874;
assign v_877 = v_872 | v_876;
assign v_879 = v_862 | v_878;
assign v_881 = v_859 | v_880;
assign v_883 = v_878 | v_882;
assign v_885 = v_858 | v_884;
assign v_887 = v_855 | v_886;
assign v_889 = v_884 | v_888;
assign v_891 = v_854 | v_890;
assign v_893 = v_851 | v_892;
assign v_895 = v_890 | v_894;
assign v_897 = v_850 | v_896;
assign v_899 = v_847 | v_898;
assign v_901 = v_896 | v_900;
assign v_903 = v_846 | v_902;
assign v_905 = v_843 | v_904;
assign v_907 = v_902 | v_906;
assign v_909 = v_842 | v_908;
assign v_911 = v_839 | v_910;
assign v_913 = v_908 | v_912;
assign v_915 = v_838 | v_914;
assign v_917 = v_835 | v_916;
assign v_919 = v_914 | v_918;
assign v_921 = v_834 | v_920;
assign v_923 = v_831 | v_922;
assign v_925 = v_920 | v_924;
assign v_927 = v_830 | v_926;
assign v_929 = v_827 | v_928;
assign v_931 = v_926 | v_930;
assign v_933 = v_826 | v_932;
assign v_935 = v_823 | v_934;
assign v_937 = v_932 | v_936;
assign v_939 = v_822 | v_938;
assign v_941 = v_819 | v_940;
assign v_943 = v_938 | v_942;
assign v_945 = v_818 | v_944;
assign v_947 = v_816 | v_946;
assign v_949 = v_944 | v_948;
assign v_951 = v_814 | v_950;
assign v_953 = v_812 | v_952;
assign v_955 = v_950 | v_954;
assign v_957 = v_810 | v_956;
assign v_959 = v_808 | v_958;
assign v_961 = v_956 | v_960;
assign v_963 = v_806 | v_962;
assign v_965 = v_804 | v_964;
assign v_967 = v_962 | v_966;
assign v_970 = ~v_802 | v_969;
assign v_977 = v_866 | v_976;
assign v_980 = v_978 | v_979;
assign v_982 = v_862 | v_981;
assign v_985 = v_983 | v_984;
assign v_987 = v_858 | v_986;
assign v_990 = v_988 | v_989;
assign v_992 = v_854 | v_991;
assign v_995 = v_993 | v_994;
assign v_997 = v_850 | v_996;
assign v_1000 = v_998 | v_999;
assign v_1002 = v_846 | v_1001;
assign v_1005 = v_1003 | v_1004;
assign v_1007 = v_842 | v_1006;
assign v_1010 = v_1008 | v_1009;
assign v_1012 = v_838 | v_1011;
assign v_1015 = v_1013 | v_1014;
assign v_1017 = v_834 | v_1016;
assign v_1020 = v_1018 | v_1019;
assign v_1022 = v_830 | v_1021;
assign v_1025 = v_1023 | v_1024;
assign v_1027 = v_826 | v_1026;
assign v_1030 = v_1028 | v_1029;
assign v_1032 = v_822 | v_1031;
assign v_1035 = v_1033 | v_1034;
assign v_1037 = v_818 | v_1036;
assign v_1040 = v_1038 | v_1039;
assign v_1042 = v_814 | v_1041;
assign v_1045 = v_1043 | v_1044;
assign v_1047 = v_810 | v_1046;
assign v_1050 = v_1048 | v_1049;
assign v_1052 = v_806 | v_1051;
assign v_1055 = v_1053 | v_1054;
assign v_1057 = v_802 | v_1056;
assign v_1060 = v_801 | v_1059;
assign v_1131 = v_1127 | v_1130;
assign v_1133 = v_1126 | v_1132;
assign v_1135 = v_1123 | v_1134;
assign v_1137 = v_1132 | v_1136;
assign v_1139 = v_1122 | v_1138;
assign v_1141 = v_1119 | v_1140;
assign v_1143 = v_1138 | v_1142;
assign v_1145 = v_1118 | v_1144;
assign v_1147 = v_1115 | v_1146;
assign v_1149 = v_1144 | v_1148;
assign v_1151 = v_1114 | v_1150;
assign v_1153 = v_1111 | v_1152;
assign v_1155 = v_1150 | v_1154;
assign v_1157 = v_1110 | v_1156;
assign v_1159 = v_1107 | v_1158;
assign v_1161 = v_1156 | v_1160;
assign v_1163 = v_1106 | v_1162;
assign v_1165 = v_1103 | v_1164;
assign v_1167 = v_1162 | v_1166;
assign v_1169 = v_1102 | v_1168;
assign v_1171 = v_1099 | v_1170;
assign v_1173 = v_1168 | v_1172;
assign v_1175 = v_1098 | v_1174;
assign v_1177 = v_1095 | v_1176;
assign v_1179 = v_1174 | v_1178;
assign v_1181 = v_1094 | v_1180;
assign v_1183 = v_1091 | v_1182;
assign v_1185 = v_1180 | v_1184;
assign v_1187 = v_1090 | v_1186;
assign v_1189 = v_1087 | v_1188;
assign v_1191 = v_1186 | v_1190;
assign v_1193 = v_1086 | v_1192;
assign v_1195 = v_1083 | v_1194;
assign v_1197 = v_1192 | v_1196;
assign v_1199 = v_1082 | v_1198;
assign v_1201 = v_1079 | v_1200;
assign v_1203 = v_1198 | v_1202;
assign v_1205 = v_1078 | v_1204;
assign v_1207 = v_1076 | v_1206;
assign v_1209 = v_1204 | v_1208;
assign v_1211 = v_1074 | v_1210;
assign v_1213 = v_1072 | v_1212;
assign v_1215 = v_1210 | v_1214;
assign v_1217 = v_1070 | v_1216;
assign v_1219 = v_1068 | v_1218;
assign v_1221 = v_1216 | v_1220;
assign v_1223 = v_1066 | v_1222;
assign v_1225 = v_1064 | v_1224;
assign v_1227 = v_1222 | v_1226;
assign v_1230 = ~v_1062 | v_1229;
assign v_1237 = v_1126 | v_1236;
assign v_1240 = v_1238 | v_1239;
assign v_1242 = v_1122 | v_1241;
assign v_1245 = v_1243 | v_1244;
assign v_1247 = v_1118 | v_1246;
assign v_1250 = v_1248 | v_1249;
assign v_1252 = v_1114 | v_1251;
assign v_1255 = v_1253 | v_1254;
assign v_1257 = v_1110 | v_1256;
assign v_1260 = v_1258 | v_1259;
assign v_1262 = v_1106 | v_1261;
assign v_1265 = v_1263 | v_1264;
assign v_1267 = v_1102 | v_1266;
assign v_1270 = v_1268 | v_1269;
assign v_1272 = v_1098 | v_1271;
assign v_1275 = v_1273 | v_1274;
assign v_1277 = v_1094 | v_1276;
assign v_1280 = v_1278 | v_1279;
assign v_1282 = v_1090 | v_1281;
assign v_1285 = v_1283 | v_1284;
assign v_1287 = v_1086 | v_1286;
assign v_1290 = v_1288 | v_1289;
assign v_1292 = v_1082 | v_1291;
assign v_1295 = v_1293 | v_1294;
assign v_1297 = v_1078 | v_1296;
assign v_1300 = v_1298 | v_1299;
assign v_1302 = v_1074 | v_1301;
assign v_1305 = v_1303 | v_1304;
assign v_1307 = v_1070 | v_1306;
assign v_1310 = v_1308 | v_1309;
assign v_1312 = v_1066 | v_1311;
assign v_1315 = v_1313 | v_1314;
assign v_1317 = v_1062 | v_1316;
assign v_1320 = v_1061 | v_1319;
assign v_1391 = v_1387 | v_1390;
assign v_1393 = v_1386 | v_1392;
assign v_1395 = v_1383 | v_1394;
assign v_1397 = v_1392 | v_1396;
assign v_1399 = v_1382 | v_1398;
assign v_1401 = v_1379 | v_1400;
assign v_1403 = v_1398 | v_1402;
assign v_1405 = v_1378 | v_1404;
assign v_1407 = v_1375 | v_1406;
assign v_1409 = v_1404 | v_1408;
assign v_1411 = v_1374 | v_1410;
assign v_1413 = v_1371 | v_1412;
assign v_1415 = v_1410 | v_1414;
assign v_1417 = v_1370 | v_1416;
assign v_1419 = v_1367 | v_1418;
assign v_1421 = v_1416 | v_1420;
assign v_1423 = v_1366 | v_1422;
assign v_1425 = v_1363 | v_1424;
assign v_1427 = v_1422 | v_1426;
assign v_1429 = v_1362 | v_1428;
assign v_1431 = v_1359 | v_1430;
assign v_1433 = v_1428 | v_1432;
assign v_1435 = v_1358 | v_1434;
assign v_1437 = v_1355 | v_1436;
assign v_1439 = v_1434 | v_1438;
assign v_1441 = v_1354 | v_1440;
assign v_1443 = v_1351 | v_1442;
assign v_1445 = v_1440 | v_1444;
assign v_1447 = v_1350 | v_1446;
assign v_1449 = v_1347 | v_1448;
assign v_1451 = v_1446 | v_1450;
assign v_1453 = v_1346 | v_1452;
assign v_1455 = v_1343 | v_1454;
assign v_1457 = v_1452 | v_1456;
assign v_1459 = v_1342 | v_1458;
assign v_1461 = v_1339 | v_1460;
assign v_1463 = v_1458 | v_1462;
assign v_1465 = v_1338 | v_1464;
assign v_1467 = v_1336 | v_1466;
assign v_1469 = v_1464 | v_1468;
assign v_1471 = v_1334 | v_1470;
assign v_1473 = v_1332 | v_1472;
assign v_1475 = v_1470 | v_1474;
assign v_1477 = v_1330 | v_1476;
assign v_1479 = v_1328 | v_1478;
assign v_1481 = v_1476 | v_1480;
assign v_1483 = v_1326 | v_1482;
assign v_1485 = v_1324 | v_1484;
assign v_1487 = v_1482 | v_1486;
assign v_1490 = ~v_1322 | v_1489;
assign v_1497 = v_1386 | v_1496;
assign v_1500 = v_1498 | v_1499;
assign v_1502 = v_1382 | v_1501;
assign v_1505 = v_1503 | v_1504;
assign v_1507 = v_1378 | v_1506;
assign v_1510 = v_1508 | v_1509;
assign v_1512 = v_1374 | v_1511;
assign v_1515 = v_1513 | v_1514;
assign v_1517 = v_1370 | v_1516;
assign v_1520 = v_1518 | v_1519;
assign v_1522 = v_1366 | v_1521;
assign v_1525 = v_1523 | v_1524;
assign v_1527 = v_1362 | v_1526;
assign v_1530 = v_1528 | v_1529;
assign v_1532 = v_1358 | v_1531;
assign v_1535 = v_1533 | v_1534;
assign v_1537 = v_1354 | v_1536;
assign v_1540 = v_1538 | v_1539;
assign v_1542 = v_1350 | v_1541;
assign v_1545 = v_1543 | v_1544;
assign v_1547 = v_1346 | v_1546;
assign v_1550 = v_1548 | v_1549;
assign v_1552 = v_1342 | v_1551;
assign v_1555 = v_1553 | v_1554;
assign v_1557 = v_1338 | v_1556;
assign v_1560 = v_1558 | v_1559;
assign v_1562 = v_1334 | v_1561;
assign v_1565 = v_1563 | v_1564;
assign v_1567 = v_1330 | v_1566;
assign v_1570 = v_1568 | v_1569;
assign v_1572 = v_1326 | v_1571;
assign v_1575 = v_1573 | v_1574;
assign v_1577 = v_1322 | v_1576;
assign v_1580 = v_1321 | v_1579;
assign v_1651 = v_1647 | v_1650;
assign v_1653 = v_1646 | v_1652;
assign v_1655 = v_1643 | v_1654;
assign v_1657 = v_1652 | v_1656;
assign v_1659 = v_1642 | v_1658;
assign v_1661 = v_1639 | v_1660;
assign v_1663 = v_1658 | v_1662;
assign v_1665 = v_1638 | v_1664;
assign v_1667 = v_1635 | v_1666;
assign v_1669 = v_1664 | v_1668;
assign v_1671 = v_1634 | v_1670;
assign v_1673 = v_1631 | v_1672;
assign v_1675 = v_1670 | v_1674;
assign v_1677 = v_1630 | v_1676;
assign v_1679 = v_1627 | v_1678;
assign v_1681 = v_1676 | v_1680;
assign v_1683 = v_1626 | v_1682;
assign v_1685 = v_1623 | v_1684;
assign v_1687 = v_1682 | v_1686;
assign v_1689 = v_1622 | v_1688;
assign v_1691 = v_1619 | v_1690;
assign v_1693 = v_1688 | v_1692;
assign v_1695 = v_1618 | v_1694;
assign v_1697 = v_1615 | v_1696;
assign v_1699 = v_1694 | v_1698;
assign v_1701 = v_1614 | v_1700;
assign v_1703 = v_1611 | v_1702;
assign v_1705 = v_1700 | v_1704;
assign v_1707 = v_1610 | v_1706;
assign v_1709 = v_1607 | v_1708;
assign v_1711 = v_1706 | v_1710;
assign v_1713 = v_1606 | v_1712;
assign v_1715 = v_1603 | v_1714;
assign v_1717 = v_1712 | v_1716;
assign v_1719 = v_1602 | v_1718;
assign v_1721 = v_1599 | v_1720;
assign v_1723 = v_1718 | v_1722;
assign v_1725 = v_1598 | v_1724;
assign v_1727 = v_1596 | v_1726;
assign v_1729 = v_1724 | v_1728;
assign v_1731 = v_1594 | v_1730;
assign v_1733 = v_1592 | v_1732;
assign v_1735 = v_1730 | v_1734;
assign v_1737 = v_1590 | v_1736;
assign v_1739 = v_1588 | v_1738;
assign v_1741 = v_1736 | v_1740;
assign v_1743 = v_1586 | v_1742;
assign v_1745 = v_1584 | v_1744;
assign v_1747 = v_1742 | v_1746;
assign v_1750 = ~v_1582 | v_1749;
assign v_1757 = v_1646 | v_1756;
assign v_1760 = v_1758 | v_1759;
assign v_1762 = v_1642 | v_1761;
assign v_1765 = v_1763 | v_1764;
assign v_1767 = v_1638 | v_1766;
assign v_1770 = v_1768 | v_1769;
assign v_1772 = v_1634 | v_1771;
assign v_1775 = v_1773 | v_1774;
assign v_1777 = v_1630 | v_1776;
assign v_1780 = v_1778 | v_1779;
assign v_1782 = v_1626 | v_1781;
assign v_1785 = v_1783 | v_1784;
assign v_1787 = v_1622 | v_1786;
assign v_1790 = v_1788 | v_1789;
assign v_1792 = v_1618 | v_1791;
assign v_1795 = v_1793 | v_1794;
assign v_1797 = v_1614 | v_1796;
assign v_1800 = v_1798 | v_1799;
assign v_1802 = v_1610 | v_1801;
assign v_1805 = v_1803 | v_1804;
assign v_1807 = v_1606 | v_1806;
assign v_1810 = v_1808 | v_1809;
assign v_1812 = v_1602 | v_1811;
assign v_1815 = v_1813 | v_1814;
assign v_1817 = v_1598 | v_1816;
assign v_1820 = v_1818 | v_1819;
assign v_1822 = v_1594 | v_1821;
assign v_1825 = v_1823 | v_1824;
assign v_1827 = v_1590 | v_1826;
assign v_1830 = v_1828 | v_1829;
assign v_1832 = v_1586 | v_1831;
assign v_1835 = v_1833 | v_1834;
assign v_1837 = v_1582 | v_1836;
assign v_1840 = v_1581 | v_1839;
assign v_1911 = v_1907 | v_1910;
assign v_1913 = v_1906 | v_1912;
assign v_1915 = v_1903 | v_1914;
assign v_1917 = v_1912 | v_1916;
assign v_1919 = v_1902 | v_1918;
assign v_1921 = v_1899 | v_1920;
assign v_1923 = v_1918 | v_1922;
assign v_1925 = v_1898 | v_1924;
assign v_1927 = v_1895 | v_1926;
assign v_1929 = v_1924 | v_1928;
assign v_1931 = v_1894 | v_1930;
assign v_1933 = v_1891 | v_1932;
assign v_1935 = v_1930 | v_1934;
assign v_1937 = v_1890 | v_1936;
assign v_1939 = v_1887 | v_1938;
assign v_1941 = v_1936 | v_1940;
assign v_1943 = v_1886 | v_1942;
assign v_1945 = v_1883 | v_1944;
assign v_1947 = v_1942 | v_1946;
assign v_1949 = v_1882 | v_1948;
assign v_1951 = v_1879 | v_1950;
assign v_1953 = v_1948 | v_1952;
assign v_1955 = v_1878 | v_1954;
assign v_1957 = v_1875 | v_1956;
assign v_1959 = v_1954 | v_1958;
assign v_1961 = v_1874 | v_1960;
assign v_1963 = v_1871 | v_1962;
assign v_1965 = v_1960 | v_1964;
assign v_1967 = v_1870 | v_1966;
assign v_1969 = v_1867 | v_1968;
assign v_1971 = v_1966 | v_1970;
assign v_1973 = v_1866 | v_1972;
assign v_1975 = v_1863 | v_1974;
assign v_1977 = v_1972 | v_1976;
assign v_1979 = v_1862 | v_1978;
assign v_1981 = v_1859 | v_1980;
assign v_1983 = v_1978 | v_1982;
assign v_1985 = v_1858 | v_1984;
assign v_1987 = v_1856 | v_1986;
assign v_1989 = v_1984 | v_1988;
assign v_1991 = v_1854 | v_1990;
assign v_1993 = v_1852 | v_1992;
assign v_1995 = v_1990 | v_1994;
assign v_1997 = v_1850 | v_1996;
assign v_1999 = v_1848 | v_1998;
assign v_2001 = v_1996 | v_2000;
assign v_2003 = v_1846 | v_2002;
assign v_2005 = v_1844 | v_2004;
assign v_2007 = v_2002 | v_2006;
assign v_2010 = ~v_1842 | v_2009;
assign v_2017 = v_1906 | v_2016;
assign v_2020 = v_2018 | v_2019;
assign v_2022 = v_1902 | v_2021;
assign v_2025 = v_2023 | v_2024;
assign v_2027 = v_1898 | v_2026;
assign v_2030 = v_2028 | v_2029;
assign v_2032 = v_1894 | v_2031;
assign v_2035 = v_2033 | v_2034;
assign v_2037 = v_1890 | v_2036;
assign v_2040 = v_2038 | v_2039;
assign v_2042 = v_1886 | v_2041;
assign v_2045 = v_2043 | v_2044;
assign v_2047 = v_1882 | v_2046;
assign v_2050 = v_2048 | v_2049;
assign v_2052 = v_1878 | v_2051;
assign v_2055 = v_2053 | v_2054;
assign v_2057 = v_1874 | v_2056;
assign v_2060 = v_2058 | v_2059;
assign v_2062 = v_1870 | v_2061;
assign v_2065 = v_2063 | v_2064;
assign v_2067 = v_1866 | v_2066;
assign v_2070 = v_2068 | v_2069;
assign v_2072 = v_1862 | v_2071;
assign v_2075 = v_2073 | v_2074;
assign v_2077 = v_1858 | v_2076;
assign v_2080 = v_2078 | v_2079;
assign v_2082 = v_1854 | v_2081;
assign v_2085 = v_2083 | v_2084;
assign v_2087 = v_1850 | v_2086;
assign v_2090 = v_2088 | v_2089;
assign v_2092 = v_1846 | v_2091;
assign v_2095 = v_2093 | v_2094;
assign v_2097 = v_1842 | v_2096;
assign v_2100 = v_1841 | v_2099;
assign v_2171 = v_2167 | v_2170;
assign v_2173 = v_2166 | v_2172;
assign v_2175 = v_2163 | v_2174;
assign v_2177 = v_2172 | v_2176;
assign v_2179 = v_2162 | v_2178;
assign v_2181 = v_2159 | v_2180;
assign v_2183 = v_2178 | v_2182;
assign v_2185 = v_2158 | v_2184;
assign v_2187 = v_2155 | v_2186;
assign v_2189 = v_2184 | v_2188;
assign v_2191 = v_2154 | v_2190;
assign v_2193 = v_2151 | v_2192;
assign v_2195 = v_2190 | v_2194;
assign v_2197 = v_2150 | v_2196;
assign v_2199 = v_2147 | v_2198;
assign v_2201 = v_2196 | v_2200;
assign v_2203 = v_2146 | v_2202;
assign v_2205 = v_2143 | v_2204;
assign v_2207 = v_2202 | v_2206;
assign v_2209 = v_2142 | v_2208;
assign v_2211 = v_2139 | v_2210;
assign v_2213 = v_2208 | v_2212;
assign v_2215 = v_2138 | v_2214;
assign v_2217 = v_2135 | v_2216;
assign v_2219 = v_2214 | v_2218;
assign v_2221 = v_2134 | v_2220;
assign v_2223 = v_2131 | v_2222;
assign v_2225 = v_2220 | v_2224;
assign v_2227 = v_2130 | v_2226;
assign v_2229 = v_2127 | v_2228;
assign v_2231 = v_2226 | v_2230;
assign v_2233 = v_2126 | v_2232;
assign v_2235 = v_2123 | v_2234;
assign v_2237 = v_2232 | v_2236;
assign v_2239 = v_2122 | v_2238;
assign v_2241 = v_2119 | v_2240;
assign v_2243 = v_2238 | v_2242;
assign v_2245 = v_2118 | v_2244;
assign v_2247 = v_2116 | v_2246;
assign v_2249 = v_2244 | v_2248;
assign v_2251 = v_2114 | v_2250;
assign v_2253 = v_2112 | v_2252;
assign v_2255 = v_2250 | v_2254;
assign v_2257 = v_2110 | v_2256;
assign v_2259 = v_2108 | v_2258;
assign v_2261 = v_2256 | v_2260;
assign v_2263 = v_2106 | v_2262;
assign v_2265 = v_2104 | v_2264;
assign v_2267 = v_2262 | v_2266;
assign v_2270 = ~v_2102 | v_2269;
assign v_2277 = v_2166 | v_2276;
assign v_2280 = v_2278 | v_2279;
assign v_2282 = v_2162 | v_2281;
assign v_2285 = v_2283 | v_2284;
assign v_2287 = v_2158 | v_2286;
assign v_2290 = v_2288 | v_2289;
assign v_2292 = v_2154 | v_2291;
assign v_2295 = v_2293 | v_2294;
assign v_2297 = v_2150 | v_2296;
assign v_2300 = v_2298 | v_2299;
assign v_2302 = v_2146 | v_2301;
assign v_2305 = v_2303 | v_2304;
assign v_2307 = v_2142 | v_2306;
assign v_2310 = v_2308 | v_2309;
assign v_2312 = v_2138 | v_2311;
assign v_2315 = v_2313 | v_2314;
assign v_2317 = v_2134 | v_2316;
assign v_2320 = v_2318 | v_2319;
assign v_2322 = v_2130 | v_2321;
assign v_2325 = v_2323 | v_2324;
assign v_2327 = v_2126 | v_2326;
assign v_2330 = v_2328 | v_2329;
assign v_2332 = v_2122 | v_2331;
assign v_2335 = v_2333 | v_2334;
assign v_2337 = v_2118 | v_2336;
assign v_2340 = v_2338 | v_2339;
assign v_2342 = v_2114 | v_2341;
assign v_2345 = v_2343 | v_2344;
assign v_2347 = v_2110 | v_2346;
assign v_2350 = v_2348 | v_2349;
assign v_2352 = v_2106 | v_2351;
assign v_2355 = v_2353 | v_2354;
assign v_2357 = v_2102 | v_2356;
assign v_2360 = v_2101 | v_2359;
assign v_2431 = v_2427 | v_2430;
assign v_2433 = v_2426 | v_2432;
assign v_2435 = v_2423 | v_2434;
assign v_2437 = v_2432 | v_2436;
assign v_2439 = v_2422 | v_2438;
assign v_2441 = v_2419 | v_2440;
assign v_2443 = v_2438 | v_2442;
assign v_2445 = v_2418 | v_2444;
assign v_2447 = v_2415 | v_2446;
assign v_2449 = v_2444 | v_2448;
assign v_2451 = v_2414 | v_2450;
assign v_2453 = v_2411 | v_2452;
assign v_2455 = v_2450 | v_2454;
assign v_2457 = v_2410 | v_2456;
assign v_2459 = v_2407 | v_2458;
assign v_2461 = v_2456 | v_2460;
assign v_2463 = v_2406 | v_2462;
assign v_2465 = v_2403 | v_2464;
assign v_2467 = v_2462 | v_2466;
assign v_2469 = v_2402 | v_2468;
assign v_2471 = v_2399 | v_2470;
assign v_2473 = v_2468 | v_2472;
assign v_2475 = v_2398 | v_2474;
assign v_2477 = v_2395 | v_2476;
assign v_2479 = v_2474 | v_2478;
assign v_2481 = v_2394 | v_2480;
assign v_2483 = v_2391 | v_2482;
assign v_2485 = v_2480 | v_2484;
assign v_2487 = v_2390 | v_2486;
assign v_2489 = v_2387 | v_2488;
assign v_2491 = v_2486 | v_2490;
assign v_2493 = v_2386 | v_2492;
assign v_2495 = v_2383 | v_2494;
assign v_2497 = v_2492 | v_2496;
assign v_2499 = v_2382 | v_2498;
assign v_2501 = v_2379 | v_2500;
assign v_2503 = v_2498 | v_2502;
assign v_2505 = v_2378 | v_2504;
assign v_2507 = v_2376 | v_2506;
assign v_2509 = v_2504 | v_2508;
assign v_2511 = v_2374 | v_2510;
assign v_2513 = v_2372 | v_2512;
assign v_2515 = v_2510 | v_2514;
assign v_2517 = v_2370 | v_2516;
assign v_2519 = v_2368 | v_2518;
assign v_2521 = v_2516 | v_2520;
assign v_2523 = v_2366 | v_2522;
assign v_2525 = v_2364 | v_2524;
assign v_2527 = v_2522 | v_2526;
assign v_2530 = ~v_2362 | v_2529;
assign v_2537 = v_2426 | v_2536;
assign v_2540 = v_2538 | v_2539;
assign v_2542 = v_2422 | v_2541;
assign v_2545 = v_2543 | v_2544;
assign v_2547 = v_2418 | v_2546;
assign v_2550 = v_2548 | v_2549;
assign v_2552 = v_2414 | v_2551;
assign v_2555 = v_2553 | v_2554;
assign v_2557 = v_2410 | v_2556;
assign v_2560 = v_2558 | v_2559;
assign v_2562 = v_2406 | v_2561;
assign v_2565 = v_2563 | v_2564;
assign v_2567 = v_2402 | v_2566;
assign v_2570 = v_2568 | v_2569;
assign v_2572 = v_2398 | v_2571;
assign v_2575 = v_2573 | v_2574;
assign v_2577 = v_2394 | v_2576;
assign v_2580 = v_2578 | v_2579;
assign v_2582 = v_2390 | v_2581;
assign v_2585 = v_2583 | v_2584;
assign v_2587 = v_2386 | v_2586;
assign v_2590 = v_2588 | v_2589;
assign v_2592 = v_2382 | v_2591;
assign v_2595 = v_2593 | v_2594;
assign v_2597 = v_2378 | v_2596;
assign v_2600 = v_2598 | v_2599;
assign v_2602 = v_2374 | v_2601;
assign v_2605 = v_2603 | v_2604;
assign v_2607 = v_2370 | v_2606;
assign v_2610 = v_2608 | v_2609;
assign v_2612 = v_2366 | v_2611;
assign v_2615 = v_2613 | v_2614;
assign v_2617 = v_2362 | v_2616;
assign v_2620 = v_2361 | v_2619;
assign v_2691 = v_2687 | v_2690;
assign v_2693 = v_2686 | v_2692;
assign v_2695 = v_2683 | v_2694;
assign v_2697 = v_2692 | v_2696;
assign v_2699 = v_2682 | v_2698;
assign v_2701 = v_2679 | v_2700;
assign v_2703 = v_2698 | v_2702;
assign v_2705 = v_2678 | v_2704;
assign v_2707 = v_2675 | v_2706;
assign v_2709 = v_2704 | v_2708;
assign v_2711 = v_2674 | v_2710;
assign v_2713 = v_2671 | v_2712;
assign v_2715 = v_2710 | v_2714;
assign v_2717 = v_2670 | v_2716;
assign v_2719 = v_2667 | v_2718;
assign v_2721 = v_2716 | v_2720;
assign v_2723 = v_2666 | v_2722;
assign v_2725 = v_2663 | v_2724;
assign v_2727 = v_2722 | v_2726;
assign v_2729 = v_2662 | v_2728;
assign v_2731 = v_2659 | v_2730;
assign v_2733 = v_2728 | v_2732;
assign v_2735 = v_2658 | v_2734;
assign v_2737 = v_2655 | v_2736;
assign v_2739 = v_2734 | v_2738;
assign v_2741 = v_2654 | v_2740;
assign v_2743 = v_2651 | v_2742;
assign v_2745 = v_2740 | v_2744;
assign v_2747 = v_2650 | v_2746;
assign v_2749 = v_2647 | v_2748;
assign v_2751 = v_2746 | v_2750;
assign v_2753 = v_2646 | v_2752;
assign v_2755 = v_2643 | v_2754;
assign v_2757 = v_2752 | v_2756;
assign v_2759 = v_2642 | v_2758;
assign v_2761 = v_2639 | v_2760;
assign v_2763 = v_2758 | v_2762;
assign v_2765 = v_2638 | v_2764;
assign v_2767 = v_2636 | v_2766;
assign v_2769 = v_2764 | v_2768;
assign v_2771 = v_2634 | v_2770;
assign v_2773 = v_2632 | v_2772;
assign v_2775 = v_2770 | v_2774;
assign v_2777 = v_2630 | v_2776;
assign v_2779 = v_2628 | v_2778;
assign v_2781 = v_2776 | v_2780;
assign v_2783 = v_2626 | v_2782;
assign v_2785 = v_2624 | v_2784;
assign v_2787 = v_2782 | v_2786;
assign v_2790 = ~v_2622 | v_2789;
assign v_2797 = v_2686 | v_2796;
assign v_2800 = v_2798 | v_2799;
assign v_2802 = v_2682 | v_2801;
assign v_2805 = v_2803 | v_2804;
assign v_2807 = v_2678 | v_2806;
assign v_2810 = v_2808 | v_2809;
assign v_2812 = v_2674 | v_2811;
assign v_2815 = v_2813 | v_2814;
assign v_2817 = v_2670 | v_2816;
assign v_2820 = v_2818 | v_2819;
assign v_2822 = v_2666 | v_2821;
assign v_2825 = v_2823 | v_2824;
assign v_2827 = v_2662 | v_2826;
assign v_2830 = v_2828 | v_2829;
assign v_2832 = v_2658 | v_2831;
assign v_2835 = v_2833 | v_2834;
assign v_2837 = v_2654 | v_2836;
assign v_2840 = v_2838 | v_2839;
assign v_2842 = v_2650 | v_2841;
assign v_2845 = v_2843 | v_2844;
assign v_2847 = v_2646 | v_2846;
assign v_2850 = v_2848 | v_2849;
assign v_2852 = v_2642 | v_2851;
assign v_2855 = v_2853 | v_2854;
assign v_2857 = v_2638 | v_2856;
assign v_2860 = v_2858 | v_2859;
assign v_2862 = v_2634 | v_2861;
assign v_2865 = v_2863 | v_2864;
assign v_2867 = v_2630 | v_2866;
assign v_2870 = v_2868 | v_2869;
assign v_2872 = v_2626 | v_2871;
assign v_2875 = v_2873 | v_2874;
assign v_2877 = v_2622 | v_2876;
assign v_2880 = v_2621 | v_2879;
assign v_2951 = v_2947 | v_2950;
assign v_2953 = v_2946 | v_2952;
assign v_2955 = v_2943 | v_2954;
assign v_2957 = v_2952 | v_2956;
assign v_2959 = v_2942 | v_2958;
assign v_2961 = v_2939 | v_2960;
assign v_2963 = v_2958 | v_2962;
assign v_2965 = v_2938 | v_2964;
assign v_2967 = v_2935 | v_2966;
assign v_2969 = v_2964 | v_2968;
assign v_2971 = v_2934 | v_2970;
assign v_2973 = v_2931 | v_2972;
assign v_2975 = v_2970 | v_2974;
assign v_2977 = v_2930 | v_2976;
assign v_2979 = v_2927 | v_2978;
assign v_2981 = v_2976 | v_2980;
assign v_2983 = v_2926 | v_2982;
assign v_2985 = v_2923 | v_2984;
assign v_2987 = v_2982 | v_2986;
assign v_2989 = v_2922 | v_2988;
assign v_2991 = v_2919 | v_2990;
assign v_2993 = v_2988 | v_2992;
assign v_2995 = v_2918 | v_2994;
assign v_2997 = v_2915 | v_2996;
assign v_2999 = v_2994 | v_2998;
assign v_3001 = v_2914 | v_3000;
assign v_3003 = v_2911 | v_3002;
assign v_3005 = v_3000 | v_3004;
assign v_3007 = v_2910 | v_3006;
assign v_3009 = v_2907 | v_3008;
assign v_3011 = v_3006 | v_3010;
assign v_3013 = v_2906 | v_3012;
assign v_3015 = v_2903 | v_3014;
assign v_3017 = v_3012 | v_3016;
assign v_3019 = v_2902 | v_3018;
assign v_3021 = v_2899 | v_3020;
assign v_3023 = v_3018 | v_3022;
assign v_3025 = v_2898 | v_3024;
assign v_3027 = v_2896 | v_3026;
assign v_3029 = v_3024 | v_3028;
assign v_3031 = v_2894 | v_3030;
assign v_3033 = v_2892 | v_3032;
assign v_3035 = v_3030 | v_3034;
assign v_3037 = v_2890 | v_3036;
assign v_3039 = v_2888 | v_3038;
assign v_3041 = v_3036 | v_3040;
assign v_3043 = v_2886 | v_3042;
assign v_3045 = v_2884 | v_3044;
assign v_3047 = v_3042 | v_3046;
assign v_3050 = ~v_2882 | v_3049;
assign v_3057 = v_2946 | v_3056;
assign v_3060 = v_3058 | v_3059;
assign v_3062 = v_2942 | v_3061;
assign v_3065 = v_3063 | v_3064;
assign v_3067 = v_2938 | v_3066;
assign v_3070 = v_3068 | v_3069;
assign v_3072 = v_2934 | v_3071;
assign v_3075 = v_3073 | v_3074;
assign v_3077 = v_2930 | v_3076;
assign v_3080 = v_3078 | v_3079;
assign v_3082 = v_2926 | v_3081;
assign v_3085 = v_3083 | v_3084;
assign v_3087 = v_2922 | v_3086;
assign v_3090 = v_3088 | v_3089;
assign v_3092 = v_2918 | v_3091;
assign v_3095 = v_3093 | v_3094;
assign v_3097 = v_2914 | v_3096;
assign v_3100 = v_3098 | v_3099;
assign v_3102 = v_2910 | v_3101;
assign v_3105 = v_3103 | v_3104;
assign v_3107 = v_2906 | v_3106;
assign v_3110 = v_3108 | v_3109;
assign v_3112 = v_2902 | v_3111;
assign v_3115 = v_3113 | v_3114;
assign v_3117 = v_2898 | v_3116;
assign v_3120 = v_3118 | v_3119;
assign v_3122 = v_2894 | v_3121;
assign v_3125 = v_3123 | v_3124;
assign v_3127 = v_2890 | v_3126;
assign v_3130 = v_3128 | v_3129;
assign v_3132 = v_2886 | v_3131;
assign v_3135 = v_3133 | v_3134;
assign v_3137 = v_2882 | v_3136;
assign v_3140 = v_2881 | v_3139;
assign v_3211 = v_3207 | v_3210;
assign v_3213 = v_3206 | v_3212;
assign v_3215 = v_3203 | v_3214;
assign v_3217 = v_3212 | v_3216;
assign v_3219 = v_3202 | v_3218;
assign v_3221 = v_3199 | v_3220;
assign v_3223 = v_3218 | v_3222;
assign v_3225 = v_3198 | v_3224;
assign v_3227 = v_3195 | v_3226;
assign v_3229 = v_3224 | v_3228;
assign v_3231 = v_3194 | v_3230;
assign v_3233 = v_3191 | v_3232;
assign v_3235 = v_3230 | v_3234;
assign v_3237 = v_3190 | v_3236;
assign v_3239 = v_3187 | v_3238;
assign v_3241 = v_3236 | v_3240;
assign v_3243 = v_3186 | v_3242;
assign v_3245 = v_3183 | v_3244;
assign v_3247 = v_3242 | v_3246;
assign v_3249 = v_3182 | v_3248;
assign v_3251 = v_3179 | v_3250;
assign v_3253 = v_3248 | v_3252;
assign v_3255 = v_3178 | v_3254;
assign v_3257 = v_3175 | v_3256;
assign v_3259 = v_3254 | v_3258;
assign v_3261 = v_3174 | v_3260;
assign v_3263 = v_3171 | v_3262;
assign v_3265 = v_3260 | v_3264;
assign v_3267 = v_3170 | v_3266;
assign v_3269 = v_3167 | v_3268;
assign v_3271 = v_3266 | v_3270;
assign v_3273 = v_3166 | v_3272;
assign v_3275 = v_3163 | v_3274;
assign v_3277 = v_3272 | v_3276;
assign v_3279 = v_3162 | v_3278;
assign v_3281 = v_3159 | v_3280;
assign v_3283 = v_3278 | v_3282;
assign v_3285 = v_3158 | v_3284;
assign v_3287 = v_3156 | v_3286;
assign v_3289 = v_3284 | v_3288;
assign v_3291 = v_3154 | v_3290;
assign v_3293 = v_3152 | v_3292;
assign v_3295 = v_3290 | v_3294;
assign v_3297 = v_3150 | v_3296;
assign v_3299 = v_3148 | v_3298;
assign v_3301 = v_3296 | v_3300;
assign v_3303 = v_3146 | v_3302;
assign v_3305 = v_3144 | v_3304;
assign v_3307 = v_3302 | v_3306;
assign v_3310 = ~v_3142 | v_3309;
assign v_3317 = v_3206 | v_3316;
assign v_3320 = v_3318 | v_3319;
assign v_3322 = v_3202 | v_3321;
assign v_3325 = v_3323 | v_3324;
assign v_3327 = v_3198 | v_3326;
assign v_3330 = v_3328 | v_3329;
assign v_3332 = v_3194 | v_3331;
assign v_3335 = v_3333 | v_3334;
assign v_3337 = v_3190 | v_3336;
assign v_3340 = v_3338 | v_3339;
assign v_3342 = v_3186 | v_3341;
assign v_3345 = v_3343 | v_3344;
assign v_3347 = v_3182 | v_3346;
assign v_3350 = v_3348 | v_3349;
assign v_3352 = v_3178 | v_3351;
assign v_3355 = v_3353 | v_3354;
assign v_3357 = v_3174 | v_3356;
assign v_3360 = v_3358 | v_3359;
assign v_3362 = v_3170 | v_3361;
assign v_3365 = v_3363 | v_3364;
assign v_3367 = v_3166 | v_3366;
assign v_3370 = v_3368 | v_3369;
assign v_3372 = v_3162 | v_3371;
assign v_3375 = v_3373 | v_3374;
assign v_3377 = v_3158 | v_3376;
assign v_3380 = v_3378 | v_3379;
assign v_3382 = v_3154 | v_3381;
assign v_3385 = v_3383 | v_3384;
assign v_3387 = v_3150 | v_3386;
assign v_3390 = v_3388 | v_3389;
assign v_3392 = v_3146 | v_3391;
assign v_3395 = v_3393 | v_3394;
assign v_3397 = v_3142 | v_3396;
assign v_3400 = v_3141 | v_3399;
assign v_3471 = v_3467 | v_3470;
assign v_3473 = v_3466 | v_3472;
assign v_3475 = v_3463 | v_3474;
assign v_3477 = v_3472 | v_3476;
assign v_3479 = v_3462 | v_3478;
assign v_3481 = v_3459 | v_3480;
assign v_3483 = v_3478 | v_3482;
assign v_3485 = v_3458 | v_3484;
assign v_3487 = v_3455 | v_3486;
assign v_3489 = v_3484 | v_3488;
assign v_3491 = v_3454 | v_3490;
assign v_3493 = v_3451 | v_3492;
assign v_3495 = v_3490 | v_3494;
assign v_3497 = v_3450 | v_3496;
assign v_3499 = v_3447 | v_3498;
assign v_3501 = v_3496 | v_3500;
assign v_3503 = v_3446 | v_3502;
assign v_3505 = v_3443 | v_3504;
assign v_3507 = v_3502 | v_3506;
assign v_3509 = v_3442 | v_3508;
assign v_3511 = v_3439 | v_3510;
assign v_3513 = v_3508 | v_3512;
assign v_3515 = v_3438 | v_3514;
assign v_3517 = v_3435 | v_3516;
assign v_3519 = v_3514 | v_3518;
assign v_3521 = v_3434 | v_3520;
assign v_3523 = v_3431 | v_3522;
assign v_3525 = v_3520 | v_3524;
assign v_3527 = v_3430 | v_3526;
assign v_3529 = v_3427 | v_3528;
assign v_3531 = v_3526 | v_3530;
assign v_3533 = v_3426 | v_3532;
assign v_3535 = v_3423 | v_3534;
assign v_3537 = v_3532 | v_3536;
assign v_3539 = v_3422 | v_3538;
assign v_3541 = v_3419 | v_3540;
assign v_3543 = v_3538 | v_3542;
assign v_3545 = v_3418 | v_3544;
assign v_3547 = v_3416 | v_3546;
assign v_3549 = v_3544 | v_3548;
assign v_3551 = v_3414 | v_3550;
assign v_3553 = v_3412 | v_3552;
assign v_3555 = v_3550 | v_3554;
assign v_3557 = v_3410 | v_3556;
assign v_3559 = v_3408 | v_3558;
assign v_3561 = v_3556 | v_3560;
assign v_3563 = v_3406 | v_3562;
assign v_3565 = v_3404 | v_3564;
assign v_3567 = v_3562 | v_3566;
assign v_3570 = ~v_3402 | v_3569;
assign v_3577 = v_3466 | v_3576;
assign v_3580 = v_3578 | v_3579;
assign v_3582 = v_3462 | v_3581;
assign v_3585 = v_3583 | v_3584;
assign v_3587 = v_3458 | v_3586;
assign v_3590 = v_3588 | v_3589;
assign v_3592 = v_3454 | v_3591;
assign v_3595 = v_3593 | v_3594;
assign v_3597 = v_3450 | v_3596;
assign v_3600 = v_3598 | v_3599;
assign v_3602 = v_3446 | v_3601;
assign v_3605 = v_3603 | v_3604;
assign v_3607 = v_3442 | v_3606;
assign v_3610 = v_3608 | v_3609;
assign v_3612 = v_3438 | v_3611;
assign v_3615 = v_3613 | v_3614;
assign v_3617 = v_3434 | v_3616;
assign v_3620 = v_3618 | v_3619;
assign v_3622 = v_3430 | v_3621;
assign v_3625 = v_3623 | v_3624;
assign v_3627 = v_3426 | v_3626;
assign v_3630 = v_3628 | v_3629;
assign v_3632 = v_3422 | v_3631;
assign v_3635 = v_3633 | v_3634;
assign v_3637 = v_3418 | v_3636;
assign v_3640 = v_3638 | v_3639;
assign v_3642 = v_3414 | v_3641;
assign v_3645 = v_3643 | v_3644;
assign v_3647 = v_3410 | v_3646;
assign v_3650 = v_3648 | v_3649;
assign v_3652 = v_3406 | v_3651;
assign v_3655 = v_3653 | v_3654;
assign v_3657 = v_3402 | v_3656;
assign v_3660 = v_3401 | v_3659;
assign v_3731 = v_3727 | v_3730;
assign v_3733 = v_3726 | v_3732;
assign v_3735 = v_3723 | v_3734;
assign v_3737 = v_3732 | v_3736;
assign v_3739 = v_3722 | v_3738;
assign v_3741 = v_3719 | v_3740;
assign v_3743 = v_3738 | v_3742;
assign v_3745 = v_3718 | v_3744;
assign v_3747 = v_3715 | v_3746;
assign v_3749 = v_3744 | v_3748;
assign v_3751 = v_3714 | v_3750;
assign v_3753 = v_3711 | v_3752;
assign v_3755 = v_3750 | v_3754;
assign v_3757 = v_3710 | v_3756;
assign v_3759 = v_3707 | v_3758;
assign v_3761 = v_3756 | v_3760;
assign v_3763 = v_3706 | v_3762;
assign v_3765 = v_3703 | v_3764;
assign v_3767 = v_3762 | v_3766;
assign v_3769 = v_3702 | v_3768;
assign v_3771 = v_3699 | v_3770;
assign v_3773 = v_3768 | v_3772;
assign v_3775 = v_3698 | v_3774;
assign v_3777 = v_3695 | v_3776;
assign v_3779 = v_3774 | v_3778;
assign v_3781 = v_3694 | v_3780;
assign v_3783 = v_3691 | v_3782;
assign v_3785 = v_3780 | v_3784;
assign v_3787 = v_3690 | v_3786;
assign v_3789 = v_3687 | v_3788;
assign v_3791 = v_3786 | v_3790;
assign v_3793 = v_3686 | v_3792;
assign v_3795 = v_3683 | v_3794;
assign v_3797 = v_3792 | v_3796;
assign v_3799 = v_3682 | v_3798;
assign v_3801 = v_3679 | v_3800;
assign v_3803 = v_3798 | v_3802;
assign v_3805 = v_3678 | v_3804;
assign v_3807 = v_3676 | v_3806;
assign v_3809 = v_3804 | v_3808;
assign v_3811 = v_3674 | v_3810;
assign v_3813 = v_3672 | v_3812;
assign v_3815 = v_3810 | v_3814;
assign v_3817 = v_3670 | v_3816;
assign v_3819 = v_3668 | v_3818;
assign v_3821 = v_3816 | v_3820;
assign v_3823 = v_3666 | v_3822;
assign v_3825 = v_3664 | v_3824;
assign v_3827 = v_3822 | v_3826;
assign v_3830 = ~v_3662 | v_3829;
assign v_3837 = v_3726 | v_3836;
assign v_3840 = v_3838 | v_3839;
assign v_3842 = v_3722 | v_3841;
assign v_3845 = v_3843 | v_3844;
assign v_3847 = v_3718 | v_3846;
assign v_3850 = v_3848 | v_3849;
assign v_3852 = v_3714 | v_3851;
assign v_3855 = v_3853 | v_3854;
assign v_3857 = v_3710 | v_3856;
assign v_3860 = v_3858 | v_3859;
assign v_3862 = v_3706 | v_3861;
assign v_3865 = v_3863 | v_3864;
assign v_3867 = v_3702 | v_3866;
assign v_3870 = v_3868 | v_3869;
assign v_3872 = v_3698 | v_3871;
assign v_3875 = v_3873 | v_3874;
assign v_3877 = v_3694 | v_3876;
assign v_3880 = v_3878 | v_3879;
assign v_3882 = v_3690 | v_3881;
assign v_3885 = v_3883 | v_3884;
assign v_3887 = v_3686 | v_3886;
assign v_3890 = v_3888 | v_3889;
assign v_3892 = v_3682 | v_3891;
assign v_3895 = v_3893 | v_3894;
assign v_3897 = v_3678 | v_3896;
assign v_3900 = v_3898 | v_3899;
assign v_3902 = v_3674 | v_3901;
assign v_3905 = v_3903 | v_3904;
assign v_3907 = v_3670 | v_3906;
assign v_3910 = v_3908 | v_3909;
assign v_3912 = v_3666 | v_3911;
assign v_3915 = v_3913 | v_3914;
assign v_3917 = v_3662 | v_3916;
assign v_3920 = v_3661 | v_3919;
assign v_3991 = v_3987 | v_3990;
assign v_3993 = v_3986 | v_3992;
assign v_3995 = v_3983 | v_3994;
assign v_3997 = v_3992 | v_3996;
assign v_3999 = v_3982 | v_3998;
assign v_4001 = v_3979 | v_4000;
assign v_4003 = v_3998 | v_4002;
assign v_4005 = v_3978 | v_4004;
assign v_4007 = v_3975 | v_4006;
assign v_4009 = v_4004 | v_4008;
assign v_4011 = v_3974 | v_4010;
assign v_4013 = v_3971 | v_4012;
assign v_4015 = v_4010 | v_4014;
assign v_4017 = v_3970 | v_4016;
assign v_4019 = v_3967 | v_4018;
assign v_4021 = v_4016 | v_4020;
assign v_4023 = v_3966 | v_4022;
assign v_4025 = v_3963 | v_4024;
assign v_4027 = v_4022 | v_4026;
assign v_4029 = v_3962 | v_4028;
assign v_4031 = v_3959 | v_4030;
assign v_4033 = v_4028 | v_4032;
assign v_4035 = v_3958 | v_4034;
assign v_4037 = v_3955 | v_4036;
assign v_4039 = v_4034 | v_4038;
assign v_4041 = v_3954 | v_4040;
assign v_4043 = v_3951 | v_4042;
assign v_4045 = v_4040 | v_4044;
assign v_4047 = v_3950 | v_4046;
assign v_4049 = v_3947 | v_4048;
assign v_4051 = v_4046 | v_4050;
assign v_4053 = v_3946 | v_4052;
assign v_4055 = v_3943 | v_4054;
assign v_4057 = v_4052 | v_4056;
assign v_4059 = v_3942 | v_4058;
assign v_4061 = v_3939 | v_4060;
assign v_4063 = v_4058 | v_4062;
assign v_4065 = v_3938 | v_4064;
assign v_4067 = v_3936 | v_4066;
assign v_4069 = v_4064 | v_4068;
assign v_4071 = v_3934 | v_4070;
assign v_4073 = v_3932 | v_4072;
assign v_4075 = v_4070 | v_4074;
assign v_4077 = v_3930 | v_4076;
assign v_4079 = v_3928 | v_4078;
assign v_4081 = v_4076 | v_4080;
assign v_4083 = v_3926 | v_4082;
assign v_4085 = v_3924 | v_4084;
assign v_4087 = v_4082 | v_4086;
assign v_4090 = ~v_3922 | v_4089;
assign v_4097 = v_3986 | v_4096;
assign v_4100 = v_4098 | v_4099;
assign v_4102 = v_3982 | v_4101;
assign v_4105 = v_4103 | v_4104;
assign v_4107 = v_3978 | v_4106;
assign v_4110 = v_4108 | v_4109;
assign v_4112 = v_3974 | v_4111;
assign v_4115 = v_4113 | v_4114;
assign v_4117 = v_3970 | v_4116;
assign v_4120 = v_4118 | v_4119;
assign v_4122 = v_3966 | v_4121;
assign v_4125 = v_4123 | v_4124;
assign v_4127 = v_3962 | v_4126;
assign v_4130 = v_4128 | v_4129;
assign v_4132 = v_3958 | v_4131;
assign v_4135 = v_4133 | v_4134;
assign v_4137 = v_3954 | v_4136;
assign v_4140 = v_4138 | v_4139;
assign v_4142 = v_3950 | v_4141;
assign v_4145 = v_4143 | v_4144;
assign v_4147 = v_3946 | v_4146;
assign v_4150 = v_4148 | v_4149;
assign v_4152 = v_3942 | v_4151;
assign v_4155 = v_4153 | v_4154;
assign v_4157 = v_3938 | v_4156;
assign v_4160 = v_4158 | v_4159;
assign v_4162 = v_3934 | v_4161;
assign v_4165 = v_4163 | v_4164;
assign v_4167 = v_3930 | v_4166;
assign v_4170 = v_4168 | v_4169;
assign v_4172 = v_3926 | v_4171;
assign v_4175 = v_4173 | v_4174;
assign v_4177 = v_3922 | v_4176;
assign v_4180 = v_3921 | v_4179;
assign v_4250 = v_4246 | v_4249;
assign v_4252 = v_4245 | v_4251;
assign v_4254 = v_4242 | v_4253;
assign v_4256 = v_4251 | v_4255;
assign v_4258 = v_4241 | v_4257;
assign v_4260 = v_4238 | v_4259;
assign v_4262 = v_4257 | v_4261;
assign v_4264 = v_4237 | v_4263;
assign v_4266 = v_4234 | v_4265;
assign v_4268 = v_4263 | v_4267;
assign v_4270 = v_4233 | v_4269;
assign v_4272 = v_4230 | v_4271;
assign v_4274 = v_4269 | v_4273;
assign v_4276 = v_4229 | v_4275;
assign v_4278 = v_4226 | v_4277;
assign v_4280 = v_4275 | v_4279;
assign v_4282 = v_4225 | v_4281;
assign v_4284 = v_4222 | v_4283;
assign v_4286 = v_4281 | v_4285;
assign v_4288 = v_4221 | v_4287;
assign v_4290 = v_4218 | v_4289;
assign v_4292 = v_4287 | v_4291;
assign v_4294 = v_4217 | v_4293;
assign v_4296 = v_4214 | v_4295;
assign v_4298 = v_4293 | v_4297;
assign v_4300 = v_4213 | v_4299;
assign v_4302 = v_4210 | v_4301;
assign v_4304 = v_4299 | v_4303;
assign v_4306 = v_4209 | v_4305;
assign v_4308 = v_4206 | v_4307;
assign v_4310 = v_4305 | v_4309;
assign v_4312 = v_4205 | v_4311;
assign v_4314 = v_4202 | v_4313;
assign v_4316 = v_4311 | v_4315;
assign v_4318 = v_4201 | v_4317;
assign v_4320 = v_4198 | v_4319;
assign v_4322 = v_4317 | v_4321;
assign v_4324 = v_4197 | v_4323;
assign v_4326 = v_4195 | v_4325;
assign v_4328 = v_4323 | v_4327;
assign v_4330 = v_4193 | v_4329;
assign v_4332 = v_4191 | v_4331;
assign v_4334 = v_4329 | v_4333;
assign v_4336 = v_4189 | v_4335;
assign v_4338 = v_4187 | v_4337;
assign v_4340 = v_4335 | v_4339;
assign v_4342 = v_4185 | v_4341;
assign v_4344 = v_4183 | v_4343;
assign v_4346 = v_4341 | v_4345;
assign v_4350 = v_4347 | v_4349;
assign v_4357 = v_4245 | v_4356;
assign v_4360 = v_4358 | v_4359;
assign v_4362 = v_4241 | v_4361;
assign v_4365 = v_4363 | v_4364;
assign v_4367 = v_4237 | v_4366;
assign v_4370 = v_4368 | v_4369;
assign v_4372 = v_4233 | v_4371;
assign v_4375 = v_4373 | v_4374;
assign v_4377 = v_4229 | v_4376;
assign v_4380 = v_4378 | v_4379;
assign v_4382 = v_4225 | v_4381;
assign v_4385 = v_4383 | v_4384;
assign v_4387 = v_4221 | v_4386;
assign v_4390 = v_4388 | v_4389;
assign v_4392 = v_4217 | v_4391;
assign v_4395 = v_4393 | v_4394;
assign v_4397 = v_4213 | v_4396;
assign v_4400 = v_4398 | v_4399;
assign v_4402 = v_4209 | v_4401;
assign v_4405 = v_4403 | v_4404;
assign v_4407 = v_4205 | v_4406;
assign v_4410 = v_4408 | v_4409;
assign v_4412 = v_4201 | v_4411;
assign v_4415 = v_4413 | v_4414;
assign v_4417 = v_4197 | v_4416;
assign v_4420 = v_4418 | v_4419;
assign v_4422 = v_4193 | v_4421;
assign v_4425 = v_4423 | v_4424;
assign v_4427 = v_4189 | v_4426;
assign v_4430 = v_4428 | v_4429;
assign v_4432 = v_4185 | v_4431;
assign v_4435 = v_4433 | v_4434;
assign v_4437 = v_4435 | v_4436;
assign v_4440 = v_4181 | v_4439;
assign v_4511 = v_4508 | v_4510;
assign v_4513 = v_4506 | v_4512;
assign v_4515 = v_4504 | v_4514;
assign v_4517 = v_4512 | v_4516;
assign v_4519 = v_4502 | v_4518;
assign v_4521 = v_4500 | v_4520;
assign v_4523 = v_4518 | v_4522;
assign v_4525 = v_4498 | v_4524;
assign v_4527 = v_4496 | v_4526;
assign v_4529 = v_4524 | v_4528;
assign v_4531 = v_4494 | v_4530;
assign v_4533 = v_4492 | v_4532;
assign v_4535 = v_4530 | v_4534;
assign v_4537 = v_4490 | v_4536;
assign v_4539 = v_4488 | v_4538;
assign v_4541 = v_4536 | v_4540;
assign v_4543 = v_4486 | v_4542;
assign v_4545 = v_4484 | v_4544;
assign v_4547 = v_4542 | v_4546;
assign v_4549 = v_4482 | v_4548;
assign v_4551 = v_4480 | v_4550;
assign v_4553 = v_4548 | v_4552;
assign v_4555 = v_4478 | v_4554;
assign v_4557 = v_4476 | v_4556;
assign v_4559 = v_4554 | v_4558;
assign v_4561 = v_4474 | v_4560;
assign v_4563 = v_4472 | v_4562;
assign v_4565 = v_4560 | v_4564;
assign v_4567 = v_4470 | v_4566;
assign v_4569 = v_4468 | v_4568;
assign v_4571 = v_4566 | v_4570;
assign v_4573 = v_4466 | v_4572;
assign v_4575 = v_4464 | v_4574;
assign v_4577 = v_4572 | v_4576;
assign v_4579 = v_4462 | v_4578;
assign v_4581 = v_4460 | v_4580;
assign v_4583 = v_4578 | v_4582;
assign v_4585 = v_4458 | v_4584;
assign v_4587 = v_4455 | v_4586;
assign v_4589 = v_4584 | v_4588;
assign v_4591 = v_4454 | v_4590;
assign v_4593 = v_4451 | v_4592;
assign v_4595 = v_4590 | v_4594;
assign v_4597 = v_4450 | v_4596;
assign v_4599 = v_4447 | v_4598;
assign v_4601 = v_4596 | v_4600;
assign v_4603 = v_4446 | v_4602;
assign v_4605 = v_4443 | v_4604;
assign v_4607 = v_4602 | v_4606;
assign v_4610 = ~v_4442 | v_4609;
assign v_4617 = v_4506 | v_4616;
assign v_4620 = v_4618 | v_4619;
assign v_4622 = v_4502 | v_4621;
assign v_4625 = v_4623 | v_4624;
assign v_4627 = v_4498 | v_4626;
assign v_4630 = v_4628 | v_4629;
assign v_4632 = v_4494 | v_4631;
assign v_4635 = v_4633 | v_4634;
assign v_4637 = v_4490 | v_4636;
assign v_4640 = v_4638 | v_4639;
assign v_4642 = v_4486 | v_4641;
assign v_4645 = v_4643 | v_4644;
assign v_4647 = v_4482 | v_4646;
assign v_4650 = v_4648 | v_4649;
assign v_4652 = v_4478 | v_4651;
assign v_4655 = v_4653 | v_4654;
assign v_4657 = v_4474 | v_4656;
assign v_4660 = v_4658 | v_4659;
assign v_4662 = v_4470 | v_4661;
assign v_4665 = v_4663 | v_4664;
assign v_4667 = v_4466 | v_4666;
assign v_4670 = v_4668 | v_4669;
assign v_4672 = v_4462 | v_4671;
assign v_4675 = v_4673 | v_4674;
assign v_4677 = v_4458 | v_4676;
assign v_4680 = v_4678 | v_4679;
assign v_4682 = v_4454 | v_4681;
assign v_4685 = v_4683 | v_4684;
assign v_4687 = v_4450 | v_4686;
assign v_4690 = v_4688 | v_4689;
assign v_4692 = v_4446 | v_4691;
assign v_4695 = v_4693 | v_4694;
assign v_4697 = v_4442 | v_4696;
assign v_4700 = v_4441 | v_4699;
assign v_4754 = v_4751 | v_4753;
assign v_4756 = v_4750 | v_4755;
assign v_4758 = v_4748 | v_4757;
assign v_4760 = v_4755 | v_4759;
assign v_4762 = v_4747 | v_4761;
assign v_4764 = v_4745 | v_4763;
assign v_4766 = v_4761 | v_4765;
assign v_4768 = v_4744 | v_4767;
assign v_4770 = v_4742 | v_4769;
assign v_4772 = v_4767 | v_4771;
assign v_4774 = v_4741 | v_4773;
assign v_4776 = v_4739 | v_4775;
assign v_4778 = v_4773 | v_4777;
assign v_4780 = v_4738 | v_4779;
assign v_4782 = v_4736 | v_4781;
assign v_4784 = v_4779 | v_4783;
assign v_4786 = v_4735 | v_4785;
assign v_4788 = v_4733 | v_4787;
assign v_4790 = v_4785 | v_4789;
assign v_4792 = v_4732 | v_4791;
assign v_4794 = v_4730 | v_4793;
assign v_4796 = v_4791 | v_4795;
assign v_4798 = v_4729 | v_4797;
assign v_4800 = v_4727 | v_4799;
assign v_4802 = v_4797 | v_4801;
assign v_4804 = v_4726 | v_4803;
assign v_4806 = v_4724 | v_4805;
assign v_4808 = v_4803 | v_4807;
assign v_4810 = v_4723 | v_4809;
assign v_4812 = v_4721 | v_4811;
assign v_4814 = v_4809 | v_4813;
assign v_4816 = v_4720 | v_4815;
assign v_4818 = v_4718 | v_4817;
assign v_4820 = v_4815 | v_4819;
assign v_4822 = v_4717 | v_4821;
assign v_4824 = v_4715 | v_4823;
assign v_4826 = v_4821 | v_4825;
assign v_4828 = v_4714 | v_4827;
assign v_4830 = v_4712 | v_4829;
assign v_4832 = v_4827 | v_4831;
assign v_4834 = v_4711 | v_4833;
assign v_4836 = v_4709 | v_4835;
assign v_4838 = v_4833 | v_4837;
assign v_4840 = v_4708 | v_4839;
assign v_4842 = v_4706 | v_4841;
assign v_4844 = v_4839 | v_4843;
assign v_4846 = v_4705 | v_4845;
assign v_4848 = v_4703 | v_4847;
assign v_4850 = v_4845 | v_4849;
assign v_4853 = ~v_4702 | v_4852;
assign v_4860 = v_4750 | v_4859;
assign v_4863 = v_4861 | v_4862;
assign v_4865 = v_4747 | v_4864;
assign v_4868 = v_4866 | v_4867;
assign v_4870 = v_4744 | v_4869;
assign v_4873 = v_4871 | v_4872;
assign v_4875 = v_4741 | v_4874;
assign v_4878 = v_4876 | v_4877;
assign v_4880 = v_4738 | v_4879;
assign v_4883 = v_4881 | v_4882;
assign v_4885 = v_4735 | v_4884;
assign v_4888 = v_4886 | v_4887;
assign v_4890 = v_4732 | v_4889;
assign v_4893 = v_4891 | v_4892;
assign v_4895 = v_4729 | v_4894;
assign v_4898 = v_4896 | v_4897;
assign v_4900 = v_4726 | v_4899;
assign v_4903 = v_4901 | v_4902;
assign v_4905 = v_4723 | v_4904;
assign v_4908 = v_4906 | v_4907;
assign v_4910 = v_4720 | v_4909;
assign v_4913 = v_4911 | v_4912;
assign v_4915 = v_4717 | v_4914;
assign v_4918 = v_4916 | v_4917;
assign v_4920 = v_4714 | v_4919;
assign v_4923 = v_4921 | v_4922;
assign v_4925 = v_4711 | v_4924;
assign v_4928 = v_4926 | v_4927;
assign v_4930 = v_4708 | v_4929;
assign v_4933 = v_4931 | v_4932;
assign v_4935 = v_4705 | v_4934;
assign v_4938 = v_4936 | v_4937;
assign v_4940 = v_4702 | v_4939;
assign v_4943 = v_4701 | v_4942;
assign v_4997 = v_4994 | v_4996;
assign v_4999 = v_4993 | v_4998;
assign v_5001 = v_4991 | v_5000;
assign v_5003 = v_4998 | v_5002;
assign v_5005 = v_4990 | v_5004;
assign v_5007 = v_4988 | v_5006;
assign v_5009 = v_5004 | v_5008;
assign v_5011 = v_4987 | v_5010;
assign v_5013 = v_4985 | v_5012;
assign v_5015 = v_5010 | v_5014;
assign v_5017 = v_4984 | v_5016;
assign v_5019 = v_4982 | v_5018;
assign v_5021 = v_5016 | v_5020;
assign v_5023 = v_4981 | v_5022;
assign v_5025 = v_4979 | v_5024;
assign v_5027 = v_5022 | v_5026;
assign v_5029 = v_4978 | v_5028;
assign v_5031 = v_4976 | v_5030;
assign v_5033 = v_5028 | v_5032;
assign v_5035 = v_4975 | v_5034;
assign v_5037 = v_4973 | v_5036;
assign v_5039 = v_5034 | v_5038;
assign v_5041 = v_4972 | v_5040;
assign v_5043 = v_4970 | v_5042;
assign v_5045 = v_5040 | v_5044;
assign v_5047 = v_4969 | v_5046;
assign v_5049 = v_4967 | v_5048;
assign v_5051 = v_5046 | v_5050;
assign v_5053 = v_4966 | v_5052;
assign v_5055 = v_4964 | v_5054;
assign v_5057 = v_5052 | v_5056;
assign v_5059 = v_4963 | v_5058;
assign v_5061 = v_4961 | v_5060;
assign v_5063 = v_5058 | v_5062;
assign v_5065 = v_4960 | v_5064;
assign v_5067 = v_4958 | v_5066;
assign v_5069 = v_5064 | v_5068;
assign v_5071 = v_4957 | v_5070;
assign v_5073 = v_4955 | v_5072;
assign v_5075 = v_5070 | v_5074;
assign v_5077 = v_4954 | v_5076;
assign v_5079 = v_4952 | v_5078;
assign v_5081 = v_5076 | v_5080;
assign v_5083 = v_4951 | v_5082;
assign v_5085 = v_4949 | v_5084;
assign v_5087 = v_5082 | v_5086;
assign v_5089 = v_4948 | v_5088;
assign v_5091 = v_4946 | v_5090;
assign v_5093 = v_5088 | v_5092;
assign v_5096 = ~v_4945 | v_5095;
assign v_5103 = v_4993 | v_5102;
assign v_5106 = v_5104 | v_5105;
assign v_5108 = v_4990 | v_5107;
assign v_5111 = v_5109 | v_5110;
assign v_5113 = v_4987 | v_5112;
assign v_5116 = v_5114 | v_5115;
assign v_5118 = v_4984 | v_5117;
assign v_5121 = v_5119 | v_5120;
assign v_5123 = v_4981 | v_5122;
assign v_5126 = v_5124 | v_5125;
assign v_5128 = v_4978 | v_5127;
assign v_5131 = v_5129 | v_5130;
assign v_5133 = v_4975 | v_5132;
assign v_5136 = v_5134 | v_5135;
assign v_5138 = v_4972 | v_5137;
assign v_5141 = v_5139 | v_5140;
assign v_5143 = v_4969 | v_5142;
assign v_5146 = v_5144 | v_5145;
assign v_5148 = v_4966 | v_5147;
assign v_5151 = v_5149 | v_5150;
assign v_5153 = v_4963 | v_5152;
assign v_5156 = v_5154 | v_5155;
assign v_5158 = v_4960 | v_5157;
assign v_5161 = v_5159 | v_5160;
assign v_5163 = v_4957 | v_5162;
assign v_5166 = v_5164 | v_5165;
assign v_5168 = v_4954 | v_5167;
assign v_5171 = v_5169 | v_5170;
assign v_5173 = v_4951 | v_5172;
assign v_5176 = v_5174 | v_5175;
assign v_5178 = v_4948 | v_5177;
assign v_5181 = v_5179 | v_5180;
assign v_5183 = v_4945 | v_5182;
assign v_5186 = v_4944 | v_5185;
assign v_5240 = v_5237 | v_5239;
assign v_5242 = v_5236 | v_5241;
assign v_5244 = v_5234 | v_5243;
assign v_5246 = v_5241 | v_5245;
assign v_5248 = v_5233 | v_5247;
assign v_5250 = v_5231 | v_5249;
assign v_5252 = v_5247 | v_5251;
assign v_5254 = v_5230 | v_5253;
assign v_5256 = v_5228 | v_5255;
assign v_5258 = v_5253 | v_5257;
assign v_5260 = v_5227 | v_5259;
assign v_5262 = v_5225 | v_5261;
assign v_5264 = v_5259 | v_5263;
assign v_5266 = v_5224 | v_5265;
assign v_5268 = v_5222 | v_5267;
assign v_5270 = v_5265 | v_5269;
assign v_5272 = v_5221 | v_5271;
assign v_5274 = v_5219 | v_5273;
assign v_5276 = v_5271 | v_5275;
assign v_5278 = v_5218 | v_5277;
assign v_5280 = v_5216 | v_5279;
assign v_5282 = v_5277 | v_5281;
assign v_5284 = v_5215 | v_5283;
assign v_5286 = v_5213 | v_5285;
assign v_5288 = v_5283 | v_5287;
assign v_5290 = v_5212 | v_5289;
assign v_5292 = v_5210 | v_5291;
assign v_5294 = v_5289 | v_5293;
assign v_5296 = v_5209 | v_5295;
assign v_5298 = v_5207 | v_5297;
assign v_5300 = v_5295 | v_5299;
assign v_5302 = v_5206 | v_5301;
assign v_5304 = v_5204 | v_5303;
assign v_5306 = v_5301 | v_5305;
assign v_5308 = v_5203 | v_5307;
assign v_5310 = v_5201 | v_5309;
assign v_5312 = v_5307 | v_5311;
assign v_5314 = v_5200 | v_5313;
assign v_5316 = v_5198 | v_5315;
assign v_5318 = v_5313 | v_5317;
assign v_5320 = v_5197 | v_5319;
assign v_5322 = v_5195 | v_5321;
assign v_5324 = v_5319 | v_5323;
assign v_5326 = v_5194 | v_5325;
assign v_5328 = v_5192 | v_5327;
assign v_5330 = v_5325 | v_5329;
assign v_5332 = v_5191 | v_5331;
assign v_5334 = v_5189 | v_5333;
assign v_5336 = v_5331 | v_5335;
assign v_5339 = ~v_5188 | v_5338;
assign v_5346 = v_5236 | v_5345;
assign v_5349 = v_5347 | v_5348;
assign v_5351 = v_5233 | v_5350;
assign v_5354 = v_5352 | v_5353;
assign v_5356 = v_5230 | v_5355;
assign v_5359 = v_5357 | v_5358;
assign v_5361 = v_5227 | v_5360;
assign v_5364 = v_5362 | v_5363;
assign v_5366 = v_5224 | v_5365;
assign v_5369 = v_5367 | v_5368;
assign v_5371 = v_5221 | v_5370;
assign v_5374 = v_5372 | v_5373;
assign v_5376 = v_5218 | v_5375;
assign v_5379 = v_5377 | v_5378;
assign v_5381 = v_5215 | v_5380;
assign v_5384 = v_5382 | v_5383;
assign v_5386 = v_5212 | v_5385;
assign v_5389 = v_5387 | v_5388;
assign v_5391 = v_5209 | v_5390;
assign v_5394 = v_5392 | v_5393;
assign v_5396 = v_5206 | v_5395;
assign v_5399 = v_5397 | v_5398;
assign v_5401 = v_5203 | v_5400;
assign v_5404 = v_5402 | v_5403;
assign v_5406 = v_5200 | v_5405;
assign v_5409 = v_5407 | v_5408;
assign v_5411 = v_5197 | v_5410;
assign v_5414 = v_5412 | v_5413;
assign v_5416 = v_5194 | v_5415;
assign v_5419 = v_5417 | v_5418;
assign v_5421 = v_5191 | v_5420;
assign v_5424 = v_5422 | v_5423;
assign v_5426 = v_5188 | v_5425;
assign v_5429 = v_5187 | v_5428;
assign v_5483 = v_5480 | v_5482;
assign v_5485 = v_5479 | v_5484;
assign v_5487 = v_5477 | v_5486;
assign v_5489 = v_5484 | v_5488;
assign v_5491 = v_5476 | v_5490;
assign v_5493 = v_5474 | v_5492;
assign v_5495 = v_5490 | v_5494;
assign v_5497 = v_5473 | v_5496;
assign v_5499 = v_5471 | v_5498;
assign v_5501 = v_5496 | v_5500;
assign v_5503 = v_5470 | v_5502;
assign v_5505 = v_5468 | v_5504;
assign v_5507 = v_5502 | v_5506;
assign v_5509 = v_5467 | v_5508;
assign v_5511 = v_5465 | v_5510;
assign v_5513 = v_5508 | v_5512;
assign v_5515 = v_5464 | v_5514;
assign v_5517 = v_5462 | v_5516;
assign v_5519 = v_5514 | v_5518;
assign v_5521 = v_5461 | v_5520;
assign v_5523 = v_5459 | v_5522;
assign v_5525 = v_5520 | v_5524;
assign v_5527 = v_5458 | v_5526;
assign v_5529 = v_5456 | v_5528;
assign v_5531 = v_5526 | v_5530;
assign v_5533 = v_5455 | v_5532;
assign v_5535 = v_5453 | v_5534;
assign v_5537 = v_5532 | v_5536;
assign v_5539 = v_5452 | v_5538;
assign v_5541 = v_5450 | v_5540;
assign v_5543 = v_5538 | v_5542;
assign v_5545 = v_5449 | v_5544;
assign v_5547 = v_5447 | v_5546;
assign v_5549 = v_5544 | v_5548;
assign v_5551 = v_5446 | v_5550;
assign v_5553 = v_5444 | v_5552;
assign v_5555 = v_5550 | v_5554;
assign v_5557 = v_5443 | v_5556;
assign v_5559 = v_5441 | v_5558;
assign v_5561 = v_5556 | v_5560;
assign v_5563 = v_5440 | v_5562;
assign v_5565 = v_5438 | v_5564;
assign v_5567 = v_5562 | v_5566;
assign v_5569 = v_5437 | v_5568;
assign v_5571 = v_5435 | v_5570;
assign v_5573 = v_5568 | v_5572;
assign v_5575 = v_5434 | v_5574;
assign v_5577 = v_5432 | v_5576;
assign v_5579 = v_5574 | v_5578;
assign v_5582 = ~v_5431 | v_5581;
assign v_5589 = v_5479 | v_5588;
assign v_5592 = v_5590 | v_5591;
assign v_5594 = v_5476 | v_5593;
assign v_5597 = v_5595 | v_5596;
assign v_5599 = v_5473 | v_5598;
assign v_5602 = v_5600 | v_5601;
assign v_5604 = v_5470 | v_5603;
assign v_5607 = v_5605 | v_5606;
assign v_5609 = v_5467 | v_5608;
assign v_5612 = v_5610 | v_5611;
assign v_5614 = v_5464 | v_5613;
assign v_5617 = v_5615 | v_5616;
assign v_5619 = v_5461 | v_5618;
assign v_5622 = v_5620 | v_5621;
assign v_5624 = v_5458 | v_5623;
assign v_5627 = v_5625 | v_5626;
assign v_5629 = v_5455 | v_5628;
assign v_5632 = v_5630 | v_5631;
assign v_5634 = v_5452 | v_5633;
assign v_5637 = v_5635 | v_5636;
assign v_5639 = v_5449 | v_5638;
assign v_5642 = v_5640 | v_5641;
assign v_5644 = v_5446 | v_5643;
assign v_5647 = v_5645 | v_5646;
assign v_5649 = v_5443 | v_5648;
assign v_5652 = v_5650 | v_5651;
assign v_5654 = v_5440 | v_5653;
assign v_5657 = v_5655 | v_5656;
assign v_5659 = v_5437 | v_5658;
assign v_5662 = v_5660 | v_5661;
assign v_5664 = v_5434 | v_5663;
assign v_5667 = v_5665 | v_5666;
assign v_5669 = v_5431 | v_5668;
assign v_5672 = v_5430 | v_5671;
assign v_5726 = v_5723 | v_5725;
assign v_5728 = v_5722 | v_5727;
assign v_5730 = v_5720 | v_5729;
assign v_5732 = v_5727 | v_5731;
assign v_5734 = v_5719 | v_5733;
assign v_5736 = v_5717 | v_5735;
assign v_5738 = v_5733 | v_5737;
assign v_5740 = v_5716 | v_5739;
assign v_5742 = v_5714 | v_5741;
assign v_5744 = v_5739 | v_5743;
assign v_5746 = v_5713 | v_5745;
assign v_5748 = v_5711 | v_5747;
assign v_5750 = v_5745 | v_5749;
assign v_5752 = v_5710 | v_5751;
assign v_5754 = v_5708 | v_5753;
assign v_5756 = v_5751 | v_5755;
assign v_5758 = v_5707 | v_5757;
assign v_5760 = v_5705 | v_5759;
assign v_5762 = v_5757 | v_5761;
assign v_5764 = v_5704 | v_5763;
assign v_5766 = v_5702 | v_5765;
assign v_5768 = v_5763 | v_5767;
assign v_5770 = v_5701 | v_5769;
assign v_5772 = v_5699 | v_5771;
assign v_5774 = v_5769 | v_5773;
assign v_5776 = v_5698 | v_5775;
assign v_5778 = v_5696 | v_5777;
assign v_5780 = v_5775 | v_5779;
assign v_5782 = v_5695 | v_5781;
assign v_5784 = v_5693 | v_5783;
assign v_5786 = v_5781 | v_5785;
assign v_5788 = v_5692 | v_5787;
assign v_5790 = v_5690 | v_5789;
assign v_5792 = v_5787 | v_5791;
assign v_5794 = v_5689 | v_5793;
assign v_5796 = v_5687 | v_5795;
assign v_5798 = v_5793 | v_5797;
assign v_5800 = v_5686 | v_5799;
assign v_5802 = v_5684 | v_5801;
assign v_5804 = v_5799 | v_5803;
assign v_5806 = v_5683 | v_5805;
assign v_5808 = v_5681 | v_5807;
assign v_5810 = v_5805 | v_5809;
assign v_5812 = v_5680 | v_5811;
assign v_5814 = v_5678 | v_5813;
assign v_5816 = v_5811 | v_5815;
assign v_5818 = v_5677 | v_5817;
assign v_5820 = v_5675 | v_5819;
assign v_5822 = v_5817 | v_5821;
assign v_5825 = ~v_5674 | v_5824;
assign v_5832 = v_5722 | v_5831;
assign v_5835 = v_5833 | v_5834;
assign v_5837 = v_5719 | v_5836;
assign v_5840 = v_5838 | v_5839;
assign v_5842 = v_5716 | v_5841;
assign v_5845 = v_5843 | v_5844;
assign v_5847 = v_5713 | v_5846;
assign v_5850 = v_5848 | v_5849;
assign v_5852 = v_5710 | v_5851;
assign v_5855 = v_5853 | v_5854;
assign v_5857 = v_5707 | v_5856;
assign v_5860 = v_5858 | v_5859;
assign v_5862 = v_5704 | v_5861;
assign v_5865 = v_5863 | v_5864;
assign v_5867 = v_5701 | v_5866;
assign v_5870 = v_5868 | v_5869;
assign v_5872 = v_5698 | v_5871;
assign v_5875 = v_5873 | v_5874;
assign v_5877 = v_5695 | v_5876;
assign v_5880 = v_5878 | v_5879;
assign v_5882 = v_5692 | v_5881;
assign v_5885 = v_5883 | v_5884;
assign v_5887 = v_5689 | v_5886;
assign v_5890 = v_5888 | v_5889;
assign v_5892 = v_5686 | v_5891;
assign v_5895 = v_5893 | v_5894;
assign v_5897 = v_5683 | v_5896;
assign v_5900 = v_5898 | v_5899;
assign v_5902 = v_5680 | v_5901;
assign v_5905 = v_5903 | v_5904;
assign v_5907 = v_5677 | v_5906;
assign v_5910 = v_5908 | v_5909;
assign v_5912 = v_5674 | v_5911;
assign v_5915 = v_5673 | v_5914;
assign v_5969 = v_5966 | v_5968;
assign v_5971 = v_5965 | v_5970;
assign v_5973 = v_5963 | v_5972;
assign v_5975 = v_5970 | v_5974;
assign v_5977 = v_5962 | v_5976;
assign v_5979 = v_5960 | v_5978;
assign v_5981 = v_5976 | v_5980;
assign v_5983 = v_5959 | v_5982;
assign v_5985 = v_5957 | v_5984;
assign v_5987 = v_5982 | v_5986;
assign v_5989 = v_5956 | v_5988;
assign v_5991 = v_5954 | v_5990;
assign v_5993 = v_5988 | v_5992;
assign v_5995 = v_5953 | v_5994;
assign v_5997 = v_5951 | v_5996;
assign v_5999 = v_5994 | v_5998;
assign v_6001 = v_5950 | v_6000;
assign v_6003 = v_5948 | v_6002;
assign v_6005 = v_6000 | v_6004;
assign v_6007 = v_5947 | v_6006;
assign v_6009 = v_5945 | v_6008;
assign v_6011 = v_6006 | v_6010;
assign v_6013 = v_5944 | v_6012;
assign v_6015 = v_5942 | v_6014;
assign v_6017 = v_6012 | v_6016;
assign v_6019 = v_5941 | v_6018;
assign v_6021 = v_5939 | v_6020;
assign v_6023 = v_6018 | v_6022;
assign v_6025 = v_5938 | v_6024;
assign v_6027 = v_5936 | v_6026;
assign v_6029 = v_6024 | v_6028;
assign v_6031 = v_5935 | v_6030;
assign v_6033 = v_5933 | v_6032;
assign v_6035 = v_6030 | v_6034;
assign v_6037 = v_5932 | v_6036;
assign v_6039 = v_5930 | v_6038;
assign v_6041 = v_6036 | v_6040;
assign v_6043 = v_5929 | v_6042;
assign v_6045 = v_5927 | v_6044;
assign v_6047 = v_6042 | v_6046;
assign v_6049 = v_5926 | v_6048;
assign v_6051 = v_5924 | v_6050;
assign v_6053 = v_6048 | v_6052;
assign v_6055 = v_5923 | v_6054;
assign v_6057 = v_5921 | v_6056;
assign v_6059 = v_6054 | v_6058;
assign v_6061 = v_5920 | v_6060;
assign v_6063 = v_5918 | v_6062;
assign v_6065 = v_6060 | v_6064;
assign v_6068 = ~v_5917 | v_6067;
assign v_6075 = v_5965 | v_6074;
assign v_6078 = v_6076 | v_6077;
assign v_6080 = v_5962 | v_6079;
assign v_6083 = v_6081 | v_6082;
assign v_6085 = v_5959 | v_6084;
assign v_6088 = v_6086 | v_6087;
assign v_6090 = v_5956 | v_6089;
assign v_6093 = v_6091 | v_6092;
assign v_6095 = v_5953 | v_6094;
assign v_6098 = v_6096 | v_6097;
assign v_6100 = v_5950 | v_6099;
assign v_6103 = v_6101 | v_6102;
assign v_6105 = v_5947 | v_6104;
assign v_6108 = v_6106 | v_6107;
assign v_6110 = v_5944 | v_6109;
assign v_6113 = v_6111 | v_6112;
assign v_6115 = v_5941 | v_6114;
assign v_6118 = v_6116 | v_6117;
assign v_6120 = v_5938 | v_6119;
assign v_6123 = v_6121 | v_6122;
assign v_6125 = v_5935 | v_6124;
assign v_6128 = v_6126 | v_6127;
assign v_6130 = v_5932 | v_6129;
assign v_6133 = v_6131 | v_6132;
assign v_6135 = v_5929 | v_6134;
assign v_6138 = v_6136 | v_6137;
assign v_6140 = v_5926 | v_6139;
assign v_6143 = v_6141 | v_6142;
assign v_6145 = v_5923 | v_6144;
assign v_6148 = v_6146 | v_6147;
assign v_6150 = v_5920 | v_6149;
assign v_6153 = v_6151 | v_6152;
assign v_6155 = v_5917 | v_6154;
assign v_6158 = v_5916 | v_6157;
assign v_6212 = v_6209 | v_6211;
assign v_6214 = v_6208 | v_6213;
assign v_6216 = v_6206 | v_6215;
assign v_6218 = v_6213 | v_6217;
assign v_6220 = v_6205 | v_6219;
assign v_6222 = v_6203 | v_6221;
assign v_6224 = v_6219 | v_6223;
assign v_6226 = v_6202 | v_6225;
assign v_6228 = v_6200 | v_6227;
assign v_6230 = v_6225 | v_6229;
assign v_6232 = v_6199 | v_6231;
assign v_6234 = v_6197 | v_6233;
assign v_6236 = v_6231 | v_6235;
assign v_6238 = v_6196 | v_6237;
assign v_6240 = v_6194 | v_6239;
assign v_6242 = v_6237 | v_6241;
assign v_6244 = v_6193 | v_6243;
assign v_6246 = v_6191 | v_6245;
assign v_6248 = v_6243 | v_6247;
assign v_6250 = v_6190 | v_6249;
assign v_6252 = v_6188 | v_6251;
assign v_6254 = v_6249 | v_6253;
assign v_6256 = v_6187 | v_6255;
assign v_6258 = v_6185 | v_6257;
assign v_6260 = v_6255 | v_6259;
assign v_6262 = v_6184 | v_6261;
assign v_6264 = v_6182 | v_6263;
assign v_6266 = v_6261 | v_6265;
assign v_6268 = v_6181 | v_6267;
assign v_6270 = v_6179 | v_6269;
assign v_6272 = v_6267 | v_6271;
assign v_6274 = v_6178 | v_6273;
assign v_6276 = v_6176 | v_6275;
assign v_6278 = v_6273 | v_6277;
assign v_6280 = v_6175 | v_6279;
assign v_6282 = v_6173 | v_6281;
assign v_6284 = v_6279 | v_6283;
assign v_6286 = v_6172 | v_6285;
assign v_6288 = v_6170 | v_6287;
assign v_6290 = v_6285 | v_6289;
assign v_6292 = v_6169 | v_6291;
assign v_6294 = v_6167 | v_6293;
assign v_6296 = v_6291 | v_6295;
assign v_6298 = v_6166 | v_6297;
assign v_6300 = v_6164 | v_6299;
assign v_6302 = v_6297 | v_6301;
assign v_6304 = v_6163 | v_6303;
assign v_6306 = v_6161 | v_6305;
assign v_6308 = v_6303 | v_6307;
assign v_6311 = ~v_6160 | v_6310;
assign v_6318 = v_6208 | v_6317;
assign v_6321 = v_6319 | v_6320;
assign v_6323 = v_6205 | v_6322;
assign v_6326 = v_6324 | v_6325;
assign v_6328 = v_6202 | v_6327;
assign v_6331 = v_6329 | v_6330;
assign v_6333 = v_6199 | v_6332;
assign v_6336 = v_6334 | v_6335;
assign v_6338 = v_6196 | v_6337;
assign v_6341 = v_6339 | v_6340;
assign v_6343 = v_6193 | v_6342;
assign v_6346 = v_6344 | v_6345;
assign v_6348 = v_6190 | v_6347;
assign v_6351 = v_6349 | v_6350;
assign v_6353 = v_6187 | v_6352;
assign v_6356 = v_6354 | v_6355;
assign v_6358 = v_6184 | v_6357;
assign v_6361 = v_6359 | v_6360;
assign v_6363 = v_6181 | v_6362;
assign v_6366 = v_6364 | v_6365;
assign v_6368 = v_6178 | v_6367;
assign v_6371 = v_6369 | v_6370;
assign v_6373 = v_6175 | v_6372;
assign v_6376 = v_6374 | v_6375;
assign v_6378 = v_6172 | v_6377;
assign v_6381 = v_6379 | v_6380;
assign v_6383 = v_6169 | v_6382;
assign v_6386 = v_6384 | v_6385;
assign v_6388 = v_6166 | v_6387;
assign v_6391 = v_6389 | v_6390;
assign v_6393 = v_6163 | v_6392;
assign v_6396 = v_6394 | v_6395;
assign v_6398 = v_6160 | v_6397;
assign v_6401 = v_6159 | v_6400;
assign v_6455 = v_6452 | v_6454;
assign v_6457 = v_6451 | v_6456;
assign v_6459 = v_6449 | v_6458;
assign v_6461 = v_6456 | v_6460;
assign v_6463 = v_6448 | v_6462;
assign v_6465 = v_6446 | v_6464;
assign v_6467 = v_6462 | v_6466;
assign v_6469 = v_6445 | v_6468;
assign v_6471 = v_6443 | v_6470;
assign v_6473 = v_6468 | v_6472;
assign v_6475 = v_6442 | v_6474;
assign v_6477 = v_6440 | v_6476;
assign v_6479 = v_6474 | v_6478;
assign v_6481 = v_6439 | v_6480;
assign v_6483 = v_6437 | v_6482;
assign v_6485 = v_6480 | v_6484;
assign v_6487 = v_6436 | v_6486;
assign v_6489 = v_6434 | v_6488;
assign v_6491 = v_6486 | v_6490;
assign v_6493 = v_6433 | v_6492;
assign v_6495 = v_6431 | v_6494;
assign v_6497 = v_6492 | v_6496;
assign v_6499 = v_6430 | v_6498;
assign v_6501 = v_6428 | v_6500;
assign v_6503 = v_6498 | v_6502;
assign v_6505 = v_6427 | v_6504;
assign v_6507 = v_6425 | v_6506;
assign v_6509 = v_6504 | v_6508;
assign v_6511 = v_6424 | v_6510;
assign v_6513 = v_6422 | v_6512;
assign v_6515 = v_6510 | v_6514;
assign v_6517 = v_6421 | v_6516;
assign v_6519 = v_6419 | v_6518;
assign v_6521 = v_6516 | v_6520;
assign v_6523 = v_6418 | v_6522;
assign v_6525 = v_6416 | v_6524;
assign v_6527 = v_6522 | v_6526;
assign v_6529 = v_6415 | v_6528;
assign v_6531 = v_6413 | v_6530;
assign v_6533 = v_6528 | v_6532;
assign v_6535 = v_6412 | v_6534;
assign v_6537 = v_6410 | v_6536;
assign v_6539 = v_6534 | v_6538;
assign v_6541 = v_6409 | v_6540;
assign v_6543 = v_6407 | v_6542;
assign v_6545 = v_6540 | v_6544;
assign v_6547 = v_6406 | v_6546;
assign v_6549 = v_6404 | v_6548;
assign v_6551 = v_6546 | v_6550;
assign v_6554 = ~v_6403 | v_6553;
assign v_6561 = v_6451 | v_6560;
assign v_6564 = v_6562 | v_6563;
assign v_6566 = v_6448 | v_6565;
assign v_6569 = v_6567 | v_6568;
assign v_6571 = v_6445 | v_6570;
assign v_6574 = v_6572 | v_6573;
assign v_6576 = v_6442 | v_6575;
assign v_6579 = v_6577 | v_6578;
assign v_6581 = v_6439 | v_6580;
assign v_6584 = v_6582 | v_6583;
assign v_6586 = v_6436 | v_6585;
assign v_6589 = v_6587 | v_6588;
assign v_6591 = v_6433 | v_6590;
assign v_6594 = v_6592 | v_6593;
assign v_6596 = v_6430 | v_6595;
assign v_6599 = v_6597 | v_6598;
assign v_6601 = v_6427 | v_6600;
assign v_6604 = v_6602 | v_6603;
assign v_6606 = v_6424 | v_6605;
assign v_6609 = v_6607 | v_6608;
assign v_6611 = v_6421 | v_6610;
assign v_6614 = v_6612 | v_6613;
assign v_6616 = v_6418 | v_6615;
assign v_6619 = v_6617 | v_6618;
assign v_6621 = v_6415 | v_6620;
assign v_6624 = v_6622 | v_6623;
assign v_6626 = v_6412 | v_6625;
assign v_6629 = v_6627 | v_6628;
assign v_6631 = v_6409 | v_6630;
assign v_6634 = v_6632 | v_6633;
assign v_6636 = v_6406 | v_6635;
assign v_6639 = v_6637 | v_6638;
assign v_6641 = v_6403 | v_6640;
assign v_6644 = v_6402 | v_6643;
assign v_6698 = v_6695 | v_6697;
assign v_6700 = v_6694 | v_6699;
assign v_6702 = v_6692 | v_6701;
assign v_6704 = v_6699 | v_6703;
assign v_6706 = v_6691 | v_6705;
assign v_6708 = v_6689 | v_6707;
assign v_6710 = v_6705 | v_6709;
assign v_6712 = v_6688 | v_6711;
assign v_6714 = v_6686 | v_6713;
assign v_6716 = v_6711 | v_6715;
assign v_6718 = v_6685 | v_6717;
assign v_6720 = v_6683 | v_6719;
assign v_6722 = v_6717 | v_6721;
assign v_6724 = v_6682 | v_6723;
assign v_6726 = v_6680 | v_6725;
assign v_6728 = v_6723 | v_6727;
assign v_6730 = v_6679 | v_6729;
assign v_6732 = v_6677 | v_6731;
assign v_6734 = v_6729 | v_6733;
assign v_6736 = v_6676 | v_6735;
assign v_6738 = v_6674 | v_6737;
assign v_6740 = v_6735 | v_6739;
assign v_6742 = v_6673 | v_6741;
assign v_6744 = v_6671 | v_6743;
assign v_6746 = v_6741 | v_6745;
assign v_6748 = v_6670 | v_6747;
assign v_6750 = v_6668 | v_6749;
assign v_6752 = v_6747 | v_6751;
assign v_6754 = v_6667 | v_6753;
assign v_6756 = v_6665 | v_6755;
assign v_6758 = v_6753 | v_6757;
assign v_6760 = v_6664 | v_6759;
assign v_6762 = v_6662 | v_6761;
assign v_6764 = v_6759 | v_6763;
assign v_6766 = v_6661 | v_6765;
assign v_6768 = v_6659 | v_6767;
assign v_6770 = v_6765 | v_6769;
assign v_6772 = v_6658 | v_6771;
assign v_6774 = v_6656 | v_6773;
assign v_6776 = v_6771 | v_6775;
assign v_6778 = v_6655 | v_6777;
assign v_6780 = v_6653 | v_6779;
assign v_6782 = v_6777 | v_6781;
assign v_6784 = v_6652 | v_6783;
assign v_6786 = v_6650 | v_6785;
assign v_6788 = v_6783 | v_6787;
assign v_6790 = v_6649 | v_6789;
assign v_6792 = v_6647 | v_6791;
assign v_6794 = v_6789 | v_6793;
assign v_6797 = ~v_6646 | v_6796;
assign v_6804 = v_6694 | v_6803;
assign v_6807 = v_6805 | v_6806;
assign v_6809 = v_6691 | v_6808;
assign v_6812 = v_6810 | v_6811;
assign v_6814 = v_6688 | v_6813;
assign v_6817 = v_6815 | v_6816;
assign v_6819 = v_6685 | v_6818;
assign v_6822 = v_6820 | v_6821;
assign v_6824 = v_6682 | v_6823;
assign v_6827 = v_6825 | v_6826;
assign v_6829 = v_6679 | v_6828;
assign v_6832 = v_6830 | v_6831;
assign v_6834 = v_6676 | v_6833;
assign v_6837 = v_6835 | v_6836;
assign v_6839 = v_6673 | v_6838;
assign v_6842 = v_6840 | v_6841;
assign v_6844 = v_6670 | v_6843;
assign v_6847 = v_6845 | v_6846;
assign v_6849 = v_6667 | v_6848;
assign v_6852 = v_6850 | v_6851;
assign v_6854 = v_6664 | v_6853;
assign v_6857 = v_6855 | v_6856;
assign v_6859 = v_6661 | v_6858;
assign v_6862 = v_6860 | v_6861;
assign v_6864 = v_6658 | v_6863;
assign v_6867 = v_6865 | v_6866;
assign v_6869 = v_6655 | v_6868;
assign v_6872 = v_6870 | v_6871;
assign v_6874 = v_6652 | v_6873;
assign v_6877 = v_6875 | v_6876;
assign v_6879 = v_6649 | v_6878;
assign v_6882 = v_6880 | v_6881;
assign v_6884 = v_6646 | v_6883;
assign v_6887 = v_6645 | v_6886;
assign v_6941 = v_6938 | v_6940;
assign v_6943 = v_6937 | v_6942;
assign v_6945 = v_6935 | v_6944;
assign v_6947 = v_6942 | v_6946;
assign v_6949 = v_6934 | v_6948;
assign v_6951 = v_6932 | v_6950;
assign v_6953 = v_6948 | v_6952;
assign v_6955 = v_6931 | v_6954;
assign v_6957 = v_6929 | v_6956;
assign v_6959 = v_6954 | v_6958;
assign v_6961 = v_6928 | v_6960;
assign v_6963 = v_6926 | v_6962;
assign v_6965 = v_6960 | v_6964;
assign v_6967 = v_6925 | v_6966;
assign v_6969 = v_6923 | v_6968;
assign v_6971 = v_6966 | v_6970;
assign v_6973 = v_6922 | v_6972;
assign v_6975 = v_6920 | v_6974;
assign v_6977 = v_6972 | v_6976;
assign v_6979 = v_6919 | v_6978;
assign v_6981 = v_6917 | v_6980;
assign v_6983 = v_6978 | v_6982;
assign v_6985 = v_6916 | v_6984;
assign v_6987 = v_6914 | v_6986;
assign v_6989 = v_6984 | v_6988;
assign v_6991 = v_6913 | v_6990;
assign v_6993 = v_6911 | v_6992;
assign v_6995 = v_6990 | v_6994;
assign v_6997 = v_6910 | v_6996;
assign v_6999 = v_6908 | v_6998;
assign v_7001 = v_6996 | v_7000;
assign v_7003 = v_6907 | v_7002;
assign v_7005 = v_6905 | v_7004;
assign v_7007 = v_7002 | v_7006;
assign v_7009 = v_6904 | v_7008;
assign v_7011 = v_6902 | v_7010;
assign v_7013 = v_7008 | v_7012;
assign v_7015 = v_6901 | v_7014;
assign v_7017 = v_6899 | v_7016;
assign v_7019 = v_7014 | v_7018;
assign v_7021 = v_6898 | v_7020;
assign v_7023 = v_6896 | v_7022;
assign v_7025 = v_7020 | v_7024;
assign v_7027 = v_6895 | v_7026;
assign v_7029 = v_6893 | v_7028;
assign v_7031 = v_7026 | v_7030;
assign v_7033 = v_6892 | v_7032;
assign v_7035 = v_6890 | v_7034;
assign v_7037 = v_7032 | v_7036;
assign v_7040 = ~v_6889 | v_7039;
assign v_7047 = v_6937 | v_7046;
assign v_7050 = v_7048 | v_7049;
assign v_7052 = v_6934 | v_7051;
assign v_7055 = v_7053 | v_7054;
assign v_7057 = v_6931 | v_7056;
assign v_7060 = v_7058 | v_7059;
assign v_7062 = v_6928 | v_7061;
assign v_7065 = v_7063 | v_7064;
assign v_7067 = v_6925 | v_7066;
assign v_7070 = v_7068 | v_7069;
assign v_7072 = v_6922 | v_7071;
assign v_7075 = v_7073 | v_7074;
assign v_7077 = v_6919 | v_7076;
assign v_7080 = v_7078 | v_7079;
assign v_7082 = v_6916 | v_7081;
assign v_7085 = v_7083 | v_7084;
assign v_7087 = v_6913 | v_7086;
assign v_7090 = v_7088 | v_7089;
assign v_7092 = v_6910 | v_7091;
assign v_7095 = v_7093 | v_7094;
assign v_7097 = v_6907 | v_7096;
assign v_7100 = v_7098 | v_7099;
assign v_7102 = v_6904 | v_7101;
assign v_7105 = v_7103 | v_7104;
assign v_7107 = v_6901 | v_7106;
assign v_7110 = v_7108 | v_7109;
assign v_7112 = v_6898 | v_7111;
assign v_7115 = v_7113 | v_7114;
assign v_7117 = v_6895 | v_7116;
assign v_7120 = v_7118 | v_7119;
assign v_7122 = v_6892 | v_7121;
assign v_7125 = v_7123 | v_7124;
assign v_7127 = v_6889 | v_7126;
assign v_7130 = v_6888 | v_7129;
assign v_7184 = v_7181 | v_7183;
assign v_7186 = v_7180 | v_7185;
assign v_7188 = v_7178 | v_7187;
assign v_7190 = v_7185 | v_7189;
assign v_7192 = v_7177 | v_7191;
assign v_7194 = v_7175 | v_7193;
assign v_7196 = v_7191 | v_7195;
assign v_7198 = v_7174 | v_7197;
assign v_7200 = v_7172 | v_7199;
assign v_7202 = v_7197 | v_7201;
assign v_7204 = v_7171 | v_7203;
assign v_7206 = v_7169 | v_7205;
assign v_7208 = v_7203 | v_7207;
assign v_7210 = v_7168 | v_7209;
assign v_7212 = v_7166 | v_7211;
assign v_7214 = v_7209 | v_7213;
assign v_7216 = v_7165 | v_7215;
assign v_7218 = v_7163 | v_7217;
assign v_7220 = v_7215 | v_7219;
assign v_7222 = v_7162 | v_7221;
assign v_7224 = v_7160 | v_7223;
assign v_7226 = v_7221 | v_7225;
assign v_7228 = v_7159 | v_7227;
assign v_7230 = v_7157 | v_7229;
assign v_7232 = v_7227 | v_7231;
assign v_7234 = v_7156 | v_7233;
assign v_7236 = v_7154 | v_7235;
assign v_7238 = v_7233 | v_7237;
assign v_7240 = v_7153 | v_7239;
assign v_7242 = v_7151 | v_7241;
assign v_7244 = v_7239 | v_7243;
assign v_7246 = v_7150 | v_7245;
assign v_7248 = v_7148 | v_7247;
assign v_7250 = v_7245 | v_7249;
assign v_7252 = v_7147 | v_7251;
assign v_7254 = v_7145 | v_7253;
assign v_7256 = v_7251 | v_7255;
assign v_7258 = v_7144 | v_7257;
assign v_7260 = v_7142 | v_7259;
assign v_7262 = v_7257 | v_7261;
assign v_7264 = v_7141 | v_7263;
assign v_7266 = v_7139 | v_7265;
assign v_7268 = v_7263 | v_7267;
assign v_7270 = v_7138 | v_7269;
assign v_7272 = v_7136 | v_7271;
assign v_7274 = v_7269 | v_7273;
assign v_7276 = v_7135 | v_7275;
assign v_7278 = v_7133 | v_7277;
assign v_7280 = v_7275 | v_7279;
assign v_7283 = ~v_7132 | v_7282;
assign v_7290 = v_7180 | v_7289;
assign v_7293 = v_7291 | v_7292;
assign v_7295 = v_7177 | v_7294;
assign v_7298 = v_7296 | v_7297;
assign v_7300 = v_7174 | v_7299;
assign v_7303 = v_7301 | v_7302;
assign v_7305 = v_7171 | v_7304;
assign v_7308 = v_7306 | v_7307;
assign v_7310 = v_7168 | v_7309;
assign v_7313 = v_7311 | v_7312;
assign v_7315 = v_7165 | v_7314;
assign v_7318 = v_7316 | v_7317;
assign v_7320 = v_7162 | v_7319;
assign v_7323 = v_7321 | v_7322;
assign v_7325 = v_7159 | v_7324;
assign v_7328 = v_7326 | v_7327;
assign v_7330 = v_7156 | v_7329;
assign v_7333 = v_7331 | v_7332;
assign v_7335 = v_7153 | v_7334;
assign v_7338 = v_7336 | v_7337;
assign v_7340 = v_7150 | v_7339;
assign v_7343 = v_7341 | v_7342;
assign v_7345 = v_7147 | v_7344;
assign v_7348 = v_7346 | v_7347;
assign v_7350 = v_7144 | v_7349;
assign v_7353 = v_7351 | v_7352;
assign v_7355 = v_7141 | v_7354;
assign v_7358 = v_7356 | v_7357;
assign v_7360 = v_7138 | v_7359;
assign v_7363 = v_7361 | v_7362;
assign v_7365 = v_7135 | v_7364;
assign v_7368 = v_7366 | v_7367;
assign v_7370 = v_7132 | v_7369;
assign v_7373 = v_7131 | v_7372;
assign v_7427 = v_7424 | v_7426;
assign v_7429 = v_7423 | v_7428;
assign v_7431 = v_7421 | v_7430;
assign v_7433 = v_7428 | v_7432;
assign v_7435 = v_7420 | v_7434;
assign v_7437 = v_7418 | v_7436;
assign v_7439 = v_7434 | v_7438;
assign v_7441 = v_7417 | v_7440;
assign v_7443 = v_7415 | v_7442;
assign v_7445 = v_7440 | v_7444;
assign v_7447 = v_7414 | v_7446;
assign v_7449 = v_7412 | v_7448;
assign v_7451 = v_7446 | v_7450;
assign v_7453 = v_7411 | v_7452;
assign v_7455 = v_7409 | v_7454;
assign v_7457 = v_7452 | v_7456;
assign v_7459 = v_7408 | v_7458;
assign v_7461 = v_7406 | v_7460;
assign v_7463 = v_7458 | v_7462;
assign v_7465 = v_7405 | v_7464;
assign v_7467 = v_7403 | v_7466;
assign v_7469 = v_7464 | v_7468;
assign v_7471 = v_7402 | v_7470;
assign v_7473 = v_7400 | v_7472;
assign v_7475 = v_7470 | v_7474;
assign v_7477 = v_7399 | v_7476;
assign v_7479 = v_7397 | v_7478;
assign v_7481 = v_7476 | v_7480;
assign v_7483 = v_7396 | v_7482;
assign v_7485 = v_7394 | v_7484;
assign v_7487 = v_7482 | v_7486;
assign v_7489 = v_7393 | v_7488;
assign v_7491 = v_7391 | v_7490;
assign v_7493 = v_7488 | v_7492;
assign v_7495 = v_7390 | v_7494;
assign v_7497 = v_7388 | v_7496;
assign v_7499 = v_7494 | v_7498;
assign v_7501 = v_7387 | v_7500;
assign v_7503 = v_7385 | v_7502;
assign v_7505 = v_7500 | v_7504;
assign v_7507 = v_7384 | v_7506;
assign v_7509 = v_7382 | v_7508;
assign v_7511 = v_7506 | v_7510;
assign v_7513 = v_7381 | v_7512;
assign v_7515 = v_7379 | v_7514;
assign v_7517 = v_7512 | v_7516;
assign v_7519 = v_7378 | v_7518;
assign v_7521 = v_7376 | v_7520;
assign v_7523 = v_7518 | v_7522;
assign v_7526 = ~v_7375 | v_7525;
assign v_7533 = v_7423 | v_7532;
assign v_7536 = v_7534 | v_7535;
assign v_7538 = v_7420 | v_7537;
assign v_7541 = v_7539 | v_7540;
assign v_7543 = v_7417 | v_7542;
assign v_7546 = v_7544 | v_7545;
assign v_7548 = v_7414 | v_7547;
assign v_7551 = v_7549 | v_7550;
assign v_7553 = v_7411 | v_7552;
assign v_7556 = v_7554 | v_7555;
assign v_7558 = v_7408 | v_7557;
assign v_7561 = v_7559 | v_7560;
assign v_7563 = v_7405 | v_7562;
assign v_7566 = v_7564 | v_7565;
assign v_7568 = v_7402 | v_7567;
assign v_7571 = v_7569 | v_7570;
assign v_7573 = v_7399 | v_7572;
assign v_7576 = v_7574 | v_7575;
assign v_7578 = v_7396 | v_7577;
assign v_7581 = v_7579 | v_7580;
assign v_7583 = v_7393 | v_7582;
assign v_7586 = v_7584 | v_7585;
assign v_7588 = v_7390 | v_7587;
assign v_7591 = v_7589 | v_7590;
assign v_7593 = v_7387 | v_7592;
assign v_7596 = v_7594 | v_7595;
assign v_7598 = v_7384 | v_7597;
assign v_7601 = v_7599 | v_7600;
assign v_7603 = v_7381 | v_7602;
assign v_7606 = v_7604 | v_7605;
assign v_7608 = v_7378 | v_7607;
assign v_7611 = v_7609 | v_7610;
assign v_7613 = v_7375 | v_7612;
assign v_7616 = v_7374 | v_7615;
assign v_7670 = v_7667 | v_7669;
assign v_7672 = v_7666 | v_7671;
assign v_7674 = v_7664 | v_7673;
assign v_7676 = v_7671 | v_7675;
assign v_7678 = v_7663 | v_7677;
assign v_7680 = v_7661 | v_7679;
assign v_7682 = v_7677 | v_7681;
assign v_7684 = v_7660 | v_7683;
assign v_7686 = v_7658 | v_7685;
assign v_7688 = v_7683 | v_7687;
assign v_7690 = v_7657 | v_7689;
assign v_7692 = v_7655 | v_7691;
assign v_7694 = v_7689 | v_7693;
assign v_7696 = v_7654 | v_7695;
assign v_7698 = v_7652 | v_7697;
assign v_7700 = v_7695 | v_7699;
assign v_7702 = v_7651 | v_7701;
assign v_7704 = v_7649 | v_7703;
assign v_7706 = v_7701 | v_7705;
assign v_7708 = v_7648 | v_7707;
assign v_7710 = v_7646 | v_7709;
assign v_7712 = v_7707 | v_7711;
assign v_7714 = v_7645 | v_7713;
assign v_7716 = v_7643 | v_7715;
assign v_7718 = v_7713 | v_7717;
assign v_7720 = v_7642 | v_7719;
assign v_7722 = v_7640 | v_7721;
assign v_7724 = v_7719 | v_7723;
assign v_7726 = v_7639 | v_7725;
assign v_7728 = v_7637 | v_7727;
assign v_7730 = v_7725 | v_7729;
assign v_7732 = v_7636 | v_7731;
assign v_7734 = v_7634 | v_7733;
assign v_7736 = v_7731 | v_7735;
assign v_7738 = v_7633 | v_7737;
assign v_7740 = v_7631 | v_7739;
assign v_7742 = v_7737 | v_7741;
assign v_7744 = v_7630 | v_7743;
assign v_7746 = v_7628 | v_7745;
assign v_7748 = v_7743 | v_7747;
assign v_7750 = v_7627 | v_7749;
assign v_7752 = v_7625 | v_7751;
assign v_7754 = v_7749 | v_7753;
assign v_7756 = v_7624 | v_7755;
assign v_7758 = v_7622 | v_7757;
assign v_7760 = v_7755 | v_7759;
assign v_7762 = v_7621 | v_7761;
assign v_7764 = v_7619 | v_7763;
assign v_7766 = v_7761 | v_7765;
assign v_7769 = ~v_7618 | v_7768;
assign v_7776 = v_7666 | v_7775;
assign v_7779 = v_7777 | v_7778;
assign v_7781 = v_7663 | v_7780;
assign v_7784 = v_7782 | v_7783;
assign v_7786 = v_7660 | v_7785;
assign v_7789 = v_7787 | v_7788;
assign v_7791 = v_7657 | v_7790;
assign v_7794 = v_7792 | v_7793;
assign v_7796 = v_7654 | v_7795;
assign v_7799 = v_7797 | v_7798;
assign v_7801 = v_7651 | v_7800;
assign v_7804 = v_7802 | v_7803;
assign v_7806 = v_7648 | v_7805;
assign v_7809 = v_7807 | v_7808;
assign v_7811 = v_7645 | v_7810;
assign v_7814 = v_7812 | v_7813;
assign v_7816 = v_7642 | v_7815;
assign v_7819 = v_7817 | v_7818;
assign v_7821 = v_7639 | v_7820;
assign v_7824 = v_7822 | v_7823;
assign v_7826 = v_7636 | v_7825;
assign v_7829 = v_7827 | v_7828;
assign v_7831 = v_7633 | v_7830;
assign v_7834 = v_7832 | v_7833;
assign v_7836 = v_7630 | v_7835;
assign v_7839 = v_7837 | v_7838;
assign v_7841 = v_7627 | v_7840;
assign v_7844 = v_7842 | v_7843;
assign v_7846 = v_7624 | v_7845;
assign v_7849 = v_7847 | v_7848;
assign v_7851 = v_7621 | v_7850;
assign v_7854 = v_7852 | v_7853;
assign v_7856 = v_7618 | v_7855;
assign v_7859 = v_7617 | v_7858;
assign v_7913 = v_7910 | v_7912;
assign v_7915 = v_7909 | v_7914;
assign v_7917 = v_7907 | v_7916;
assign v_7919 = v_7914 | v_7918;
assign v_7921 = v_7906 | v_7920;
assign v_7923 = v_7904 | v_7922;
assign v_7925 = v_7920 | v_7924;
assign v_7927 = v_7903 | v_7926;
assign v_7929 = v_7901 | v_7928;
assign v_7931 = v_7926 | v_7930;
assign v_7933 = v_7900 | v_7932;
assign v_7935 = v_7898 | v_7934;
assign v_7937 = v_7932 | v_7936;
assign v_7939 = v_7897 | v_7938;
assign v_7941 = v_7895 | v_7940;
assign v_7943 = v_7938 | v_7942;
assign v_7945 = v_7894 | v_7944;
assign v_7947 = v_7892 | v_7946;
assign v_7949 = v_7944 | v_7948;
assign v_7951 = v_7891 | v_7950;
assign v_7953 = v_7889 | v_7952;
assign v_7955 = v_7950 | v_7954;
assign v_7957 = v_7888 | v_7956;
assign v_7959 = v_7886 | v_7958;
assign v_7961 = v_7956 | v_7960;
assign v_7963 = v_7885 | v_7962;
assign v_7965 = v_7883 | v_7964;
assign v_7967 = v_7962 | v_7966;
assign v_7969 = v_7882 | v_7968;
assign v_7971 = v_7880 | v_7970;
assign v_7973 = v_7968 | v_7972;
assign v_7975 = v_7879 | v_7974;
assign v_7977 = v_7877 | v_7976;
assign v_7979 = v_7974 | v_7978;
assign v_7981 = v_7876 | v_7980;
assign v_7983 = v_7874 | v_7982;
assign v_7985 = v_7980 | v_7984;
assign v_7987 = v_7873 | v_7986;
assign v_7989 = v_7871 | v_7988;
assign v_7991 = v_7986 | v_7990;
assign v_7993 = v_7870 | v_7992;
assign v_7995 = v_7868 | v_7994;
assign v_7997 = v_7992 | v_7996;
assign v_7999 = v_7867 | v_7998;
assign v_8001 = v_7865 | v_8000;
assign v_8003 = v_7998 | v_8002;
assign v_8005 = v_7864 | v_8004;
assign v_8007 = v_7862 | v_8006;
assign v_8009 = v_8004 | v_8008;
assign v_8012 = ~v_7861 | v_8011;
assign v_8019 = v_7909 | v_8018;
assign v_8022 = v_8020 | v_8021;
assign v_8024 = v_7906 | v_8023;
assign v_8027 = v_8025 | v_8026;
assign v_8029 = v_7903 | v_8028;
assign v_8032 = v_8030 | v_8031;
assign v_8034 = v_7900 | v_8033;
assign v_8037 = v_8035 | v_8036;
assign v_8039 = v_7897 | v_8038;
assign v_8042 = v_8040 | v_8041;
assign v_8044 = v_7894 | v_8043;
assign v_8047 = v_8045 | v_8046;
assign v_8049 = v_7891 | v_8048;
assign v_8052 = v_8050 | v_8051;
assign v_8054 = v_7888 | v_8053;
assign v_8057 = v_8055 | v_8056;
assign v_8059 = v_7885 | v_8058;
assign v_8062 = v_8060 | v_8061;
assign v_8064 = v_7882 | v_8063;
assign v_8067 = v_8065 | v_8066;
assign v_8069 = v_7879 | v_8068;
assign v_8072 = v_8070 | v_8071;
assign v_8074 = v_7876 | v_8073;
assign v_8077 = v_8075 | v_8076;
assign v_8079 = v_7873 | v_8078;
assign v_8082 = v_8080 | v_8081;
assign v_8084 = v_7870 | v_8083;
assign v_8087 = v_8085 | v_8086;
assign v_8089 = v_7867 | v_8088;
assign v_8092 = v_8090 | v_8091;
assign v_8094 = v_7864 | v_8093;
assign v_8097 = v_8095 | v_8096;
assign v_8099 = v_7861 | v_8098;
assign v_8102 = v_7860 | v_8101;
assign v_8156 = v_8153 | v_8155;
assign v_8158 = v_8152 | v_8157;
assign v_8160 = v_8150 | v_8159;
assign v_8162 = v_8157 | v_8161;
assign v_8164 = v_8149 | v_8163;
assign v_8166 = v_8147 | v_8165;
assign v_8168 = v_8163 | v_8167;
assign v_8170 = v_8146 | v_8169;
assign v_8172 = v_8144 | v_8171;
assign v_8174 = v_8169 | v_8173;
assign v_8176 = v_8143 | v_8175;
assign v_8178 = v_8141 | v_8177;
assign v_8180 = v_8175 | v_8179;
assign v_8182 = v_8140 | v_8181;
assign v_8184 = v_8138 | v_8183;
assign v_8186 = v_8181 | v_8185;
assign v_8188 = v_8137 | v_8187;
assign v_8190 = v_8135 | v_8189;
assign v_8192 = v_8187 | v_8191;
assign v_8194 = v_8134 | v_8193;
assign v_8196 = v_8132 | v_8195;
assign v_8198 = v_8193 | v_8197;
assign v_8200 = v_8131 | v_8199;
assign v_8202 = v_8129 | v_8201;
assign v_8204 = v_8199 | v_8203;
assign v_8206 = v_8128 | v_8205;
assign v_8208 = v_8126 | v_8207;
assign v_8210 = v_8205 | v_8209;
assign v_8212 = v_8125 | v_8211;
assign v_8214 = v_8123 | v_8213;
assign v_8216 = v_8211 | v_8215;
assign v_8218 = v_8122 | v_8217;
assign v_8220 = v_8120 | v_8219;
assign v_8222 = v_8217 | v_8221;
assign v_8224 = v_8119 | v_8223;
assign v_8226 = v_8117 | v_8225;
assign v_8228 = v_8223 | v_8227;
assign v_8230 = v_8116 | v_8229;
assign v_8232 = v_8114 | v_8231;
assign v_8234 = v_8229 | v_8233;
assign v_8236 = v_8113 | v_8235;
assign v_8238 = v_8111 | v_8237;
assign v_8240 = v_8235 | v_8239;
assign v_8242 = v_8110 | v_8241;
assign v_8244 = v_8108 | v_8243;
assign v_8246 = v_8241 | v_8245;
assign v_8248 = v_8107 | v_8247;
assign v_8250 = v_8105 | v_8249;
assign v_8252 = v_8247 | v_8251;
assign v_8255 = ~v_8104 | v_8254;
assign v_8262 = v_8152 | v_8261;
assign v_8265 = v_8263 | v_8264;
assign v_8267 = v_8149 | v_8266;
assign v_8270 = v_8268 | v_8269;
assign v_8272 = v_8146 | v_8271;
assign v_8275 = v_8273 | v_8274;
assign v_8277 = v_8143 | v_8276;
assign v_8280 = v_8278 | v_8279;
assign v_8282 = v_8140 | v_8281;
assign v_8285 = v_8283 | v_8284;
assign v_8287 = v_8137 | v_8286;
assign v_8290 = v_8288 | v_8289;
assign v_8292 = v_8134 | v_8291;
assign v_8295 = v_8293 | v_8294;
assign v_8297 = v_8131 | v_8296;
assign v_8300 = v_8298 | v_8299;
assign v_8302 = v_8128 | v_8301;
assign v_8305 = v_8303 | v_8304;
assign v_8307 = v_8125 | v_8306;
assign v_8310 = v_8308 | v_8309;
assign v_8312 = v_8122 | v_8311;
assign v_8315 = v_8313 | v_8314;
assign v_8317 = v_8119 | v_8316;
assign v_8320 = v_8318 | v_8319;
assign v_8322 = v_8116 | v_8321;
assign v_8325 = v_8323 | v_8324;
assign v_8327 = v_8113 | v_8326;
assign v_8330 = v_8328 | v_8329;
assign v_8332 = v_8110 | v_8331;
assign v_8335 = v_8333 | v_8334;
assign v_8337 = v_8107 | v_8336;
assign v_8340 = v_8338 | v_8339;
assign v_8342 = v_8104 | v_8341;
assign v_8345 = v_8103 | v_8344;
assign v_8398 = v_8395 | v_8397;
assign v_8400 = v_8394 | v_8399;
assign v_8402 = v_8392 | v_8401;
assign v_8404 = v_8399 | v_8403;
assign v_8406 = v_8391 | v_8405;
assign v_8408 = v_8389 | v_8407;
assign v_8410 = v_8405 | v_8409;
assign v_8412 = v_8388 | v_8411;
assign v_8414 = v_8386 | v_8413;
assign v_8416 = v_8411 | v_8415;
assign v_8418 = v_8385 | v_8417;
assign v_8420 = v_8383 | v_8419;
assign v_8422 = v_8417 | v_8421;
assign v_8424 = v_8382 | v_8423;
assign v_8426 = v_8380 | v_8425;
assign v_8428 = v_8423 | v_8427;
assign v_8430 = v_8379 | v_8429;
assign v_8432 = v_8377 | v_8431;
assign v_8434 = v_8429 | v_8433;
assign v_8436 = v_8376 | v_8435;
assign v_8438 = v_8374 | v_8437;
assign v_8440 = v_8435 | v_8439;
assign v_8442 = v_8373 | v_8441;
assign v_8444 = v_8371 | v_8443;
assign v_8446 = v_8441 | v_8445;
assign v_8448 = v_8370 | v_8447;
assign v_8450 = v_8368 | v_8449;
assign v_8452 = v_8447 | v_8451;
assign v_8454 = v_8367 | v_8453;
assign v_8456 = v_8365 | v_8455;
assign v_8458 = v_8453 | v_8457;
assign v_8460 = v_8364 | v_8459;
assign v_8462 = v_8362 | v_8461;
assign v_8464 = v_8459 | v_8463;
assign v_8466 = v_8361 | v_8465;
assign v_8468 = v_8359 | v_8467;
assign v_8470 = v_8465 | v_8469;
assign v_8472 = v_8358 | v_8471;
assign v_8474 = v_8356 | v_8473;
assign v_8476 = v_8471 | v_8475;
assign v_8478 = v_8355 | v_8477;
assign v_8480 = v_8353 | v_8479;
assign v_8482 = v_8477 | v_8481;
assign v_8484 = v_8352 | v_8483;
assign v_8486 = v_8350 | v_8485;
assign v_8488 = v_8483 | v_8487;
assign v_8490 = v_8349 | v_8489;
assign v_8492 = v_8347 | v_8491;
assign v_8494 = v_8489 | v_8493;
assign v_8498 = v_8495 | v_8497;
assign v_8505 = v_8394 | v_8504;
assign v_8508 = v_8506 | v_8507;
assign v_8510 = v_8391 | v_8509;
assign v_8513 = v_8511 | v_8512;
assign v_8515 = v_8388 | v_8514;
assign v_8518 = v_8516 | v_8517;
assign v_8520 = v_8385 | v_8519;
assign v_8523 = v_8521 | v_8522;
assign v_8525 = v_8382 | v_8524;
assign v_8528 = v_8526 | v_8527;
assign v_8530 = v_8379 | v_8529;
assign v_8533 = v_8531 | v_8532;
assign v_8535 = v_8376 | v_8534;
assign v_8538 = v_8536 | v_8537;
assign v_8540 = v_8373 | v_8539;
assign v_8543 = v_8541 | v_8542;
assign v_8545 = v_8370 | v_8544;
assign v_8548 = v_8546 | v_8547;
assign v_8550 = v_8367 | v_8549;
assign v_8553 = v_8551 | v_8552;
assign v_8555 = v_8364 | v_8554;
assign v_8558 = v_8556 | v_8557;
assign v_8560 = v_8361 | v_8559;
assign v_8563 = v_8561 | v_8562;
assign v_8565 = v_8358 | v_8564;
assign v_8568 = v_8566 | v_8567;
assign v_8570 = v_8355 | v_8569;
assign v_8573 = v_8571 | v_8572;
assign v_8575 = v_8352 | v_8574;
assign v_8578 = v_8576 | v_8577;
assign v_8580 = v_8349 | v_8579;
assign v_8583 = v_8581 | v_8582;
assign v_8585 = v_8583 | v_8584;
assign v_8588 = v_8346 | v_8587;
assign v_8659 = v_8656 | v_8658;
assign v_8661 = v_8654 | v_8660;
assign v_8663 = v_8652 | v_8662;
assign v_8665 = v_8660 | v_8664;
assign v_8667 = v_8650 | v_8666;
assign v_8669 = v_8648 | v_8668;
assign v_8671 = v_8666 | v_8670;
assign v_8673 = v_8646 | v_8672;
assign v_8675 = v_8644 | v_8674;
assign v_8677 = v_8672 | v_8676;
assign v_8679 = v_8642 | v_8678;
assign v_8681 = v_8640 | v_8680;
assign v_8683 = v_8678 | v_8682;
assign v_8685 = v_8638 | v_8684;
assign v_8687 = v_8636 | v_8686;
assign v_8689 = v_8684 | v_8688;
assign v_8691 = v_8634 | v_8690;
assign v_8693 = v_8632 | v_8692;
assign v_8695 = v_8690 | v_8694;
assign v_8697 = v_8630 | v_8696;
assign v_8699 = v_8628 | v_8698;
assign v_8701 = v_8696 | v_8700;
assign v_8703 = v_8626 | v_8702;
assign v_8705 = v_8624 | v_8704;
assign v_8707 = v_8702 | v_8706;
assign v_8709 = v_8622 | v_8708;
assign v_8711 = v_8620 | v_8710;
assign v_8713 = v_8708 | v_8712;
assign v_8715 = v_8618 | v_8714;
assign v_8717 = v_8616 | v_8716;
assign v_8719 = v_8714 | v_8718;
assign v_8721 = v_8614 | v_8720;
assign v_8723 = v_8612 | v_8722;
assign v_8725 = v_8720 | v_8724;
assign v_8727 = v_8610 | v_8726;
assign v_8729 = v_8608 | v_8728;
assign v_8731 = v_8726 | v_8730;
assign v_8733 = v_8606 | v_8732;
assign v_8735 = v_8603 | v_8734;
assign v_8737 = v_8732 | v_8736;
assign v_8739 = v_8602 | v_8738;
assign v_8741 = v_8599 | v_8740;
assign v_8743 = v_8738 | v_8742;
assign v_8745 = v_8598 | v_8744;
assign v_8747 = v_8595 | v_8746;
assign v_8749 = v_8744 | v_8748;
assign v_8751 = v_8594 | v_8750;
assign v_8753 = v_8591 | v_8752;
assign v_8755 = v_8750 | v_8754;
assign v_8758 = ~v_8590 | v_8757;
assign v_8765 = v_8654 | v_8764;
assign v_8768 = v_8766 | v_8767;
assign v_8770 = v_8650 | v_8769;
assign v_8773 = v_8771 | v_8772;
assign v_8775 = v_8646 | v_8774;
assign v_8778 = v_8776 | v_8777;
assign v_8780 = v_8642 | v_8779;
assign v_8783 = v_8781 | v_8782;
assign v_8785 = v_8638 | v_8784;
assign v_8788 = v_8786 | v_8787;
assign v_8790 = v_8634 | v_8789;
assign v_8793 = v_8791 | v_8792;
assign v_8795 = v_8630 | v_8794;
assign v_8798 = v_8796 | v_8797;
assign v_8800 = v_8626 | v_8799;
assign v_8803 = v_8801 | v_8802;
assign v_8805 = v_8622 | v_8804;
assign v_8808 = v_8806 | v_8807;
assign v_8810 = v_8618 | v_8809;
assign v_8813 = v_8811 | v_8812;
assign v_8815 = v_8614 | v_8814;
assign v_8818 = v_8816 | v_8817;
assign v_8820 = v_8610 | v_8819;
assign v_8823 = v_8821 | v_8822;
assign v_8825 = v_8606 | v_8824;
assign v_8828 = v_8826 | v_8827;
assign v_8830 = v_8602 | v_8829;
assign v_8833 = v_8831 | v_8832;
assign v_8835 = v_8598 | v_8834;
assign v_8838 = v_8836 | v_8837;
assign v_8840 = v_8594 | v_8839;
assign v_8843 = v_8841 | v_8842;
assign v_8845 = v_8590 | v_8844;
assign v_8848 = v_8589 | v_8847;
assign v_8902 = v_8899 | v_8901;
assign v_8904 = v_8898 | v_8903;
assign v_8906 = v_8896 | v_8905;
assign v_8908 = v_8903 | v_8907;
assign v_8910 = v_8895 | v_8909;
assign v_8912 = v_8893 | v_8911;
assign v_8914 = v_8909 | v_8913;
assign v_8916 = v_8892 | v_8915;
assign v_8918 = v_8890 | v_8917;
assign v_8920 = v_8915 | v_8919;
assign v_8922 = v_8889 | v_8921;
assign v_8924 = v_8887 | v_8923;
assign v_8926 = v_8921 | v_8925;
assign v_8928 = v_8886 | v_8927;
assign v_8930 = v_8884 | v_8929;
assign v_8932 = v_8927 | v_8931;
assign v_8934 = v_8883 | v_8933;
assign v_8936 = v_8881 | v_8935;
assign v_8938 = v_8933 | v_8937;
assign v_8940 = v_8880 | v_8939;
assign v_8942 = v_8878 | v_8941;
assign v_8944 = v_8939 | v_8943;
assign v_8946 = v_8877 | v_8945;
assign v_8948 = v_8875 | v_8947;
assign v_8950 = v_8945 | v_8949;
assign v_8952 = v_8874 | v_8951;
assign v_8954 = v_8872 | v_8953;
assign v_8956 = v_8951 | v_8955;
assign v_8958 = v_8871 | v_8957;
assign v_8960 = v_8869 | v_8959;
assign v_8962 = v_8957 | v_8961;
assign v_8964 = v_8868 | v_8963;
assign v_8966 = v_8866 | v_8965;
assign v_8968 = v_8963 | v_8967;
assign v_8970 = v_8865 | v_8969;
assign v_8972 = v_8863 | v_8971;
assign v_8974 = v_8969 | v_8973;
assign v_8976 = v_8862 | v_8975;
assign v_8978 = v_8860 | v_8977;
assign v_8980 = v_8975 | v_8979;
assign v_8982 = v_8859 | v_8981;
assign v_8984 = v_8857 | v_8983;
assign v_8986 = v_8981 | v_8985;
assign v_8988 = v_8856 | v_8987;
assign v_8990 = v_8854 | v_8989;
assign v_8992 = v_8987 | v_8991;
assign v_8994 = v_8853 | v_8993;
assign v_8996 = v_8851 | v_8995;
assign v_8998 = v_8993 | v_8997;
assign v_9001 = ~v_8850 | v_9000;
assign v_9008 = v_8898 | v_9007;
assign v_9011 = v_9009 | v_9010;
assign v_9013 = v_8895 | v_9012;
assign v_9016 = v_9014 | v_9015;
assign v_9018 = v_8892 | v_9017;
assign v_9021 = v_9019 | v_9020;
assign v_9023 = v_8889 | v_9022;
assign v_9026 = v_9024 | v_9025;
assign v_9028 = v_8886 | v_9027;
assign v_9031 = v_9029 | v_9030;
assign v_9033 = v_8883 | v_9032;
assign v_9036 = v_9034 | v_9035;
assign v_9038 = v_8880 | v_9037;
assign v_9041 = v_9039 | v_9040;
assign v_9043 = v_8877 | v_9042;
assign v_9046 = v_9044 | v_9045;
assign v_9048 = v_8874 | v_9047;
assign v_9051 = v_9049 | v_9050;
assign v_9053 = v_8871 | v_9052;
assign v_9056 = v_9054 | v_9055;
assign v_9058 = v_8868 | v_9057;
assign v_9061 = v_9059 | v_9060;
assign v_9063 = v_8865 | v_9062;
assign v_9066 = v_9064 | v_9065;
assign v_9068 = v_8862 | v_9067;
assign v_9071 = v_9069 | v_9070;
assign v_9073 = v_8859 | v_9072;
assign v_9076 = v_9074 | v_9075;
assign v_9078 = v_8856 | v_9077;
assign v_9081 = v_9079 | v_9080;
assign v_9083 = v_8853 | v_9082;
assign v_9086 = v_9084 | v_9085;
assign v_9088 = v_8850 | v_9087;
assign v_9091 = v_8849 | v_9090;
assign v_9145 = v_9142 | v_9144;
assign v_9147 = v_9141 | v_9146;
assign v_9149 = v_9139 | v_9148;
assign v_9151 = v_9146 | v_9150;
assign v_9153 = v_9138 | v_9152;
assign v_9155 = v_9136 | v_9154;
assign v_9157 = v_9152 | v_9156;
assign v_9159 = v_9135 | v_9158;
assign v_9161 = v_9133 | v_9160;
assign v_9163 = v_9158 | v_9162;
assign v_9165 = v_9132 | v_9164;
assign v_9167 = v_9130 | v_9166;
assign v_9169 = v_9164 | v_9168;
assign v_9171 = v_9129 | v_9170;
assign v_9173 = v_9127 | v_9172;
assign v_9175 = v_9170 | v_9174;
assign v_9177 = v_9126 | v_9176;
assign v_9179 = v_9124 | v_9178;
assign v_9181 = v_9176 | v_9180;
assign v_9183 = v_9123 | v_9182;
assign v_9185 = v_9121 | v_9184;
assign v_9187 = v_9182 | v_9186;
assign v_9189 = v_9120 | v_9188;
assign v_9191 = v_9118 | v_9190;
assign v_9193 = v_9188 | v_9192;
assign v_9195 = v_9117 | v_9194;
assign v_9197 = v_9115 | v_9196;
assign v_9199 = v_9194 | v_9198;
assign v_9201 = v_9114 | v_9200;
assign v_9203 = v_9112 | v_9202;
assign v_9205 = v_9200 | v_9204;
assign v_9207 = v_9111 | v_9206;
assign v_9209 = v_9109 | v_9208;
assign v_9211 = v_9206 | v_9210;
assign v_9213 = v_9108 | v_9212;
assign v_9215 = v_9106 | v_9214;
assign v_9217 = v_9212 | v_9216;
assign v_9219 = v_9105 | v_9218;
assign v_9221 = v_9103 | v_9220;
assign v_9223 = v_9218 | v_9222;
assign v_9225 = v_9102 | v_9224;
assign v_9227 = v_9100 | v_9226;
assign v_9229 = v_9224 | v_9228;
assign v_9231 = v_9099 | v_9230;
assign v_9233 = v_9097 | v_9232;
assign v_9235 = v_9230 | v_9234;
assign v_9237 = v_9096 | v_9236;
assign v_9239 = v_9094 | v_9238;
assign v_9241 = v_9236 | v_9240;
assign v_9244 = ~v_9093 | v_9243;
assign v_9251 = v_9141 | v_9250;
assign v_9254 = v_9252 | v_9253;
assign v_9256 = v_9138 | v_9255;
assign v_9259 = v_9257 | v_9258;
assign v_9261 = v_9135 | v_9260;
assign v_9264 = v_9262 | v_9263;
assign v_9266 = v_9132 | v_9265;
assign v_9269 = v_9267 | v_9268;
assign v_9271 = v_9129 | v_9270;
assign v_9274 = v_9272 | v_9273;
assign v_9276 = v_9126 | v_9275;
assign v_9279 = v_9277 | v_9278;
assign v_9281 = v_9123 | v_9280;
assign v_9284 = v_9282 | v_9283;
assign v_9286 = v_9120 | v_9285;
assign v_9289 = v_9287 | v_9288;
assign v_9291 = v_9117 | v_9290;
assign v_9294 = v_9292 | v_9293;
assign v_9296 = v_9114 | v_9295;
assign v_9299 = v_9297 | v_9298;
assign v_9301 = v_9111 | v_9300;
assign v_9304 = v_9302 | v_9303;
assign v_9306 = v_9108 | v_9305;
assign v_9309 = v_9307 | v_9308;
assign v_9311 = v_9105 | v_9310;
assign v_9314 = v_9312 | v_9313;
assign v_9316 = v_9102 | v_9315;
assign v_9319 = v_9317 | v_9318;
assign v_9321 = v_9099 | v_9320;
assign v_9324 = v_9322 | v_9323;
assign v_9326 = v_9096 | v_9325;
assign v_9329 = v_9327 | v_9328;
assign v_9331 = v_9093 | v_9330;
assign v_9334 = v_9092 | v_9333;
assign v_9388 = v_9385 | v_9387;
assign v_9390 = v_9384 | v_9389;
assign v_9392 = v_9382 | v_9391;
assign v_9394 = v_9389 | v_9393;
assign v_9396 = v_9381 | v_9395;
assign v_9398 = v_9379 | v_9397;
assign v_9400 = v_9395 | v_9399;
assign v_9402 = v_9378 | v_9401;
assign v_9404 = v_9376 | v_9403;
assign v_9406 = v_9401 | v_9405;
assign v_9408 = v_9375 | v_9407;
assign v_9410 = v_9373 | v_9409;
assign v_9412 = v_9407 | v_9411;
assign v_9414 = v_9372 | v_9413;
assign v_9416 = v_9370 | v_9415;
assign v_9418 = v_9413 | v_9417;
assign v_9420 = v_9369 | v_9419;
assign v_9422 = v_9367 | v_9421;
assign v_9424 = v_9419 | v_9423;
assign v_9426 = v_9366 | v_9425;
assign v_9428 = v_9364 | v_9427;
assign v_9430 = v_9425 | v_9429;
assign v_9432 = v_9363 | v_9431;
assign v_9434 = v_9361 | v_9433;
assign v_9436 = v_9431 | v_9435;
assign v_9438 = v_9360 | v_9437;
assign v_9440 = v_9358 | v_9439;
assign v_9442 = v_9437 | v_9441;
assign v_9444 = v_9357 | v_9443;
assign v_9446 = v_9355 | v_9445;
assign v_9448 = v_9443 | v_9447;
assign v_9450 = v_9354 | v_9449;
assign v_9452 = v_9352 | v_9451;
assign v_9454 = v_9449 | v_9453;
assign v_9456 = v_9351 | v_9455;
assign v_9458 = v_9349 | v_9457;
assign v_9460 = v_9455 | v_9459;
assign v_9462 = v_9348 | v_9461;
assign v_9464 = v_9346 | v_9463;
assign v_9466 = v_9461 | v_9465;
assign v_9468 = v_9345 | v_9467;
assign v_9470 = v_9343 | v_9469;
assign v_9472 = v_9467 | v_9471;
assign v_9474 = v_9342 | v_9473;
assign v_9476 = v_9340 | v_9475;
assign v_9478 = v_9473 | v_9477;
assign v_9480 = v_9339 | v_9479;
assign v_9482 = v_9337 | v_9481;
assign v_9484 = v_9479 | v_9483;
assign v_9487 = ~v_9336 | v_9486;
assign v_9494 = v_9384 | v_9493;
assign v_9497 = v_9495 | v_9496;
assign v_9499 = v_9381 | v_9498;
assign v_9502 = v_9500 | v_9501;
assign v_9504 = v_9378 | v_9503;
assign v_9507 = v_9505 | v_9506;
assign v_9509 = v_9375 | v_9508;
assign v_9512 = v_9510 | v_9511;
assign v_9514 = v_9372 | v_9513;
assign v_9517 = v_9515 | v_9516;
assign v_9519 = v_9369 | v_9518;
assign v_9522 = v_9520 | v_9521;
assign v_9524 = v_9366 | v_9523;
assign v_9527 = v_9525 | v_9526;
assign v_9529 = v_9363 | v_9528;
assign v_9532 = v_9530 | v_9531;
assign v_9534 = v_9360 | v_9533;
assign v_9537 = v_9535 | v_9536;
assign v_9539 = v_9357 | v_9538;
assign v_9542 = v_9540 | v_9541;
assign v_9544 = v_9354 | v_9543;
assign v_9547 = v_9545 | v_9546;
assign v_9549 = v_9351 | v_9548;
assign v_9552 = v_9550 | v_9551;
assign v_9554 = v_9348 | v_9553;
assign v_9557 = v_9555 | v_9556;
assign v_9559 = v_9345 | v_9558;
assign v_9562 = v_9560 | v_9561;
assign v_9564 = v_9342 | v_9563;
assign v_9567 = v_9565 | v_9566;
assign v_9569 = v_9339 | v_9568;
assign v_9572 = v_9570 | v_9571;
assign v_9574 = v_9336 | v_9573;
assign v_9577 = v_9335 | v_9576;
assign v_9631 = v_9628 | v_9630;
assign v_9633 = v_9627 | v_9632;
assign v_9635 = v_9625 | v_9634;
assign v_9637 = v_9632 | v_9636;
assign v_9639 = v_9624 | v_9638;
assign v_9641 = v_9622 | v_9640;
assign v_9643 = v_9638 | v_9642;
assign v_9645 = v_9621 | v_9644;
assign v_9647 = v_9619 | v_9646;
assign v_9649 = v_9644 | v_9648;
assign v_9651 = v_9618 | v_9650;
assign v_9653 = v_9616 | v_9652;
assign v_9655 = v_9650 | v_9654;
assign v_9657 = v_9615 | v_9656;
assign v_9659 = v_9613 | v_9658;
assign v_9661 = v_9656 | v_9660;
assign v_9663 = v_9612 | v_9662;
assign v_9665 = v_9610 | v_9664;
assign v_9667 = v_9662 | v_9666;
assign v_9669 = v_9609 | v_9668;
assign v_9671 = v_9607 | v_9670;
assign v_9673 = v_9668 | v_9672;
assign v_9675 = v_9606 | v_9674;
assign v_9677 = v_9604 | v_9676;
assign v_9679 = v_9674 | v_9678;
assign v_9681 = v_9603 | v_9680;
assign v_9683 = v_9601 | v_9682;
assign v_9685 = v_9680 | v_9684;
assign v_9687 = v_9600 | v_9686;
assign v_9689 = v_9598 | v_9688;
assign v_9691 = v_9686 | v_9690;
assign v_9693 = v_9597 | v_9692;
assign v_9695 = v_9595 | v_9694;
assign v_9697 = v_9692 | v_9696;
assign v_9699 = v_9594 | v_9698;
assign v_9701 = v_9592 | v_9700;
assign v_9703 = v_9698 | v_9702;
assign v_9705 = v_9591 | v_9704;
assign v_9707 = v_9589 | v_9706;
assign v_9709 = v_9704 | v_9708;
assign v_9711 = v_9588 | v_9710;
assign v_9713 = v_9586 | v_9712;
assign v_9715 = v_9710 | v_9714;
assign v_9717 = v_9585 | v_9716;
assign v_9719 = v_9583 | v_9718;
assign v_9721 = v_9716 | v_9720;
assign v_9723 = v_9582 | v_9722;
assign v_9725 = v_9580 | v_9724;
assign v_9727 = v_9722 | v_9726;
assign v_9730 = ~v_9579 | v_9729;
assign v_9737 = v_9627 | v_9736;
assign v_9740 = v_9738 | v_9739;
assign v_9742 = v_9624 | v_9741;
assign v_9745 = v_9743 | v_9744;
assign v_9747 = v_9621 | v_9746;
assign v_9750 = v_9748 | v_9749;
assign v_9752 = v_9618 | v_9751;
assign v_9755 = v_9753 | v_9754;
assign v_9757 = v_9615 | v_9756;
assign v_9760 = v_9758 | v_9759;
assign v_9762 = v_9612 | v_9761;
assign v_9765 = v_9763 | v_9764;
assign v_9767 = v_9609 | v_9766;
assign v_9770 = v_9768 | v_9769;
assign v_9772 = v_9606 | v_9771;
assign v_9775 = v_9773 | v_9774;
assign v_9777 = v_9603 | v_9776;
assign v_9780 = v_9778 | v_9779;
assign v_9782 = v_9600 | v_9781;
assign v_9785 = v_9783 | v_9784;
assign v_9787 = v_9597 | v_9786;
assign v_9790 = v_9788 | v_9789;
assign v_9792 = v_9594 | v_9791;
assign v_9795 = v_9793 | v_9794;
assign v_9797 = v_9591 | v_9796;
assign v_9800 = v_9798 | v_9799;
assign v_9802 = v_9588 | v_9801;
assign v_9805 = v_9803 | v_9804;
assign v_9807 = v_9585 | v_9806;
assign v_9810 = v_9808 | v_9809;
assign v_9812 = v_9582 | v_9811;
assign v_9815 = v_9813 | v_9814;
assign v_9817 = v_9579 | v_9816;
assign v_9820 = v_9578 | v_9819;
assign v_9874 = v_9871 | v_9873;
assign v_9876 = v_9870 | v_9875;
assign v_9878 = v_9868 | v_9877;
assign v_9880 = v_9875 | v_9879;
assign v_9882 = v_9867 | v_9881;
assign v_9884 = v_9865 | v_9883;
assign v_9886 = v_9881 | v_9885;
assign v_9888 = v_9864 | v_9887;
assign v_9890 = v_9862 | v_9889;
assign v_9892 = v_9887 | v_9891;
assign v_9894 = v_9861 | v_9893;
assign v_9896 = v_9859 | v_9895;
assign v_9898 = v_9893 | v_9897;
assign v_9900 = v_9858 | v_9899;
assign v_9902 = v_9856 | v_9901;
assign v_9904 = v_9899 | v_9903;
assign v_9906 = v_9855 | v_9905;
assign v_9908 = v_9853 | v_9907;
assign v_9910 = v_9905 | v_9909;
assign v_9912 = v_9852 | v_9911;
assign v_9914 = v_9850 | v_9913;
assign v_9916 = v_9911 | v_9915;
assign v_9918 = v_9849 | v_9917;
assign v_9920 = v_9847 | v_9919;
assign v_9922 = v_9917 | v_9921;
assign v_9924 = v_9846 | v_9923;
assign v_9926 = v_9844 | v_9925;
assign v_9928 = v_9923 | v_9927;
assign v_9930 = v_9843 | v_9929;
assign v_9932 = v_9841 | v_9931;
assign v_9934 = v_9929 | v_9933;
assign v_9936 = v_9840 | v_9935;
assign v_9938 = v_9838 | v_9937;
assign v_9940 = v_9935 | v_9939;
assign v_9942 = v_9837 | v_9941;
assign v_9944 = v_9835 | v_9943;
assign v_9946 = v_9941 | v_9945;
assign v_9948 = v_9834 | v_9947;
assign v_9950 = v_9832 | v_9949;
assign v_9952 = v_9947 | v_9951;
assign v_9954 = v_9831 | v_9953;
assign v_9956 = v_9829 | v_9955;
assign v_9958 = v_9953 | v_9957;
assign v_9960 = v_9828 | v_9959;
assign v_9962 = v_9826 | v_9961;
assign v_9964 = v_9959 | v_9963;
assign v_9966 = v_9825 | v_9965;
assign v_9968 = v_9823 | v_9967;
assign v_9970 = v_9965 | v_9969;
assign v_9973 = ~v_9822 | v_9972;
assign v_9980 = v_9870 | v_9979;
assign v_9983 = v_9981 | v_9982;
assign v_9985 = v_9867 | v_9984;
assign v_9988 = v_9986 | v_9987;
assign v_9990 = v_9864 | v_9989;
assign v_9993 = v_9991 | v_9992;
assign v_9995 = v_9861 | v_9994;
assign v_9998 = v_9996 | v_9997;
assign v_10000 = v_9858 | v_9999;
assign v_10003 = v_10001 | v_10002;
assign v_10005 = v_9855 | v_10004;
assign v_10008 = v_10006 | v_10007;
assign v_10010 = v_9852 | v_10009;
assign v_10013 = v_10011 | v_10012;
assign v_10015 = v_9849 | v_10014;
assign v_10018 = v_10016 | v_10017;
assign v_10020 = v_9846 | v_10019;
assign v_10023 = v_10021 | v_10022;
assign v_10025 = v_9843 | v_10024;
assign v_10028 = v_10026 | v_10027;
assign v_10030 = v_9840 | v_10029;
assign v_10033 = v_10031 | v_10032;
assign v_10035 = v_9837 | v_10034;
assign v_10038 = v_10036 | v_10037;
assign v_10040 = v_9834 | v_10039;
assign v_10043 = v_10041 | v_10042;
assign v_10045 = v_9831 | v_10044;
assign v_10048 = v_10046 | v_10047;
assign v_10050 = v_9828 | v_10049;
assign v_10053 = v_10051 | v_10052;
assign v_10055 = v_9825 | v_10054;
assign v_10058 = v_10056 | v_10057;
assign v_10060 = v_9822 | v_10059;
assign v_10063 = v_9821 | v_10062;
assign v_10117 = v_10114 | v_10116;
assign v_10119 = v_10113 | v_10118;
assign v_10121 = v_10111 | v_10120;
assign v_10123 = v_10118 | v_10122;
assign v_10125 = v_10110 | v_10124;
assign v_10127 = v_10108 | v_10126;
assign v_10129 = v_10124 | v_10128;
assign v_10131 = v_10107 | v_10130;
assign v_10133 = v_10105 | v_10132;
assign v_10135 = v_10130 | v_10134;
assign v_10137 = v_10104 | v_10136;
assign v_10139 = v_10102 | v_10138;
assign v_10141 = v_10136 | v_10140;
assign v_10143 = v_10101 | v_10142;
assign v_10145 = v_10099 | v_10144;
assign v_10147 = v_10142 | v_10146;
assign v_10149 = v_10098 | v_10148;
assign v_10151 = v_10096 | v_10150;
assign v_10153 = v_10148 | v_10152;
assign v_10155 = v_10095 | v_10154;
assign v_10157 = v_10093 | v_10156;
assign v_10159 = v_10154 | v_10158;
assign v_10161 = v_10092 | v_10160;
assign v_10163 = v_10090 | v_10162;
assign v_10165 = v_10160 | v_10164;
assign v_10167 = v_10089 | v_10166;
assign v_10169 = v_10087 | v_10168;
assign v_10171 = v_10166 | v_10170;
assign v_10173 = v_10086 | v_10172;
assign v_10175 = v_10084 | v_10174;
assign v_10177 = v_10172 | v_10176;
assign v_10179 = v_10083 | v_10178;
assign v_10181 = v_10081 | v_10180;
assign v_10183 = v_10178 | v_10182;
assign v_10185 = v_10080 | v_10184;
assign v_10187 = v_10078 | v_10186;
assign v_10189 = v_10184 | v_10188;
assign v_10191 = v_10077 | v_10190;
assign v_10193 = v_10075 | v_10192;
assign v_10195 = v_10190 | v_10194;
assign v_10197 = v_10074 | v_10196;
assign v_10199 = v_10072 | v_10198;
assign v_10201 = v_10196 | v_10200;
assign v_10203 = v_10071 | v_10202;
assign v_10205 = v_10069 | v_10204;
assign v_10207 = v_10202 | v_10206;
assign v_10209 = v_10068 | v_10208;
assign v_10211 = v_10066 | v_10210;
assign v_10213 = v_10208 | v_10212;
assign v_10216 = ~v_10065 | v_10215;
assign v_10223 = v_10113 | v_10222;
assign v_10226 = v_10224 | v_10225;
assign v_10228 = v_10110 | v_10227;
assign v_10231 = v_10229 | v_10230;
assign v_10233 = v_10107 | v_10232;
assign v_10236 = v_10234 | v_10235;
assign v_10238 = v_10104 | v_10237;
assign v_10241 = v_10239 | v_10240;
assign v_10243 = v_10101 | v_10242;
assign v_10246 = v_10244 | v_10245;
assign v_10248 = v_10098 | v_10247;
assign v_10251 = v_10249 | v_10250;
assign v_10253 = v_10095 | v_10252;
assign v_10256 = v_10254 | v_10255;
assign v_10258 = v_10092 | v_10257;
assign v_10261 = v_10259 | v_10260;
assign v_10263 = v_10089 | v_10262;
assign v_10266 = v_10264 | v_10265;
assign v_10268 = v_10086 | v_10267;
assign v_10271 = v_10269 | v_10270;
assign v_10273 = v_10083 | v_10272;
assign v_10276 = v_10274 | v_10275;
assign v_10278 = v_10080 | v_10277;
assign v_10281 = v_10279 | v_10280;
assign v_10283 = v_10077 | v_10282;
assign v_10286 = v_10284 | v_10285;
assign v_10288 = v_10074 | v_10287;
assign v_10291 = v_10289 | v_10290;
assign v_10293 = v_10071 | v_10292;
assign v_10296 = v_10294 | v_10295;
assign v_10298 = v_10068 | v_10297;
assign v_10301 = v_10299 | v_10300;
assign v_10303 = v_10065 | v_10302;
assign v_10306 = v_10064 | v_10305;
assign v_10360 = v_10357 | v_10359;
assign v_10362 = v_10356 | v_10361;
assign v_10364 = v_10354 | v_10363;
assign v_10366 = v_10361 | v_10365;
assign v_10368 = v_10353 | v_10367;
assign v_10370 = v_10351 | v_10369;
assign v_10372 = v_10367 | v_10371;
assign v_10374 = v_10350 | v_10373;
assign v_10376 = v_10348 | v_10375;
assign v_10378 = v_10373 | v_10377;
assign v_10380 = v_10347 | v_10379;
assign v_10382 = v_10345 | v_10381;
assign v_10384 = v_10379 | v_10383;
assign v_10386 = v_10344 | v_10385;
assign v_10388 = v_10342 | v_10387;
assign v_10390 = v_10385 | v_10389;
assign v_10392 = v_10341 | v_10391;
assign v_10394 = v_10339 | v_10393;
assign v_10396 = v_10391 | v_10395;
assign v_10398 = v_10338 | v_10397;
assign v_10400 = v_10336 | v_10399;
assign v_10402 = v_10397 | v_10401;
assign v_10404 = v_10335 | v_10403;
assign v_10406 = v_10333 | v_10405;
assign v_10408 = v_10403 | v_10407;
assign v_10410 = v_10332 | v_10409;
assign v_10412 = v_10330 | v_10411;
assign v_10414 = v_10409 | v_10413;
assign v_10416 = v_10329 | v_10415;
assign v_10418 = v_10327 | v_10417;
assign v_10420 = v_10415 | v_10419;
assign v_10422 = v_10326 | v_10421;
assign v_10424 = v_10324 | v_10423;
assign v_10426 = v_10421 | v_10425;
assign v_10428 = v_10323 | v_10427;
assign v_10430 = v_10321 | v_10429;
assign v_10432 = v_10427 | v_10431;
assign v_10434 = v_10320 | v_10433;
assign v_10436 = v_10318 | v_10435;
assign v_10438 = v_10433 | v_10437;
assign v_10440 = v_10317 | v_10439;
assign v_10442 = v_10315 | v_10441;
assign v_10444 = v_10439 | v_10443;
assign v_10446 = v_10314 | v_10445;
assign v_10448 = v_10312 | v_10447;
assign v_10450 = v_10445 | v_10449;
assign v_10452 = v_10311 | v_10451;
assign v_10454 = v_10309 | v_10453;
assign v_10456 = v_10451 | v_10455;
assign v_10459 = ~v_10308 | v_10458;
assign v_10466 = v_10356 | v_10465;
assign v_10469 = v_10467 | v_10468;
assign v_10471 = v_10353 | v_10470;
assign v_10474 = v_10472 | v_10473;
assign v_10476 = v_10350 | v_10475;
assign v_10479 = v_10477 | v_10478;
assign v_10481 = v_10347 | v_10480;
assign v_10484 = v_10482 | v_10483;
assign v_10486 = v_10344 | v_10485;
assign v_10489 = v_10487 | v_10488;
assign v_10491 = v_10341 | v_10490;
assign v_10494 = v_10492 | v_10493;
assign v_10496 = v_10338 | v_10495;
assign v_10499 = v_10497 | v_10498;
assign v_10501 = v_10335 | v_10500;
assign v_10504 = v_10502 | v_10503;
assign v_10506 = v_10332 | v_10505;
assign v_10509 = v_10507 | v_10508;
assign v_10511 = v_10329 | v_10510;
assign v_10514 = v_10512 | v_10513;
assign v_10516 = v_10326 | v_10515;
assign v_10519 = v_10517 | v_10518;
assign v_10521 = v_10323 | v_10520;
assign v_10524 = v_10522 | v_10523;
assign v_10526 = v_10320 | v_10525;
assign v_10529 = v_10527 | v_10528;
assign v_10531 = v_10317 | v_10530;
assign v_10534 = v_10532 | v_10533;
assign v_10536 = v_10314 | v_10535;
assign v_10539 = v_10537 | v_10538;
assign v_10541 = v_10311 | v_10540;
assign v_10544 = v_10542 | v_10543;
assign v_10546 = v_10308 | v_10545;
assign v_10549 = v_10307 | v_10548;
assign v_10603 = v_10600 | v_10602;
assign v_10605 = v_10599 | v_10604;
assign v_10607 = v_10597 | v_10606;
assign v_10609 = v_10604 | v_10608;
assign v_10611 = v_10596 | v_10610;
assign v_10613 = v_10594 | v_10612;
assign v_10615 = v_10610 | v_10614;
assign v_10617 = v_10593 | v_10616;
assign v_10619 = v_10591 | v_10618;
assign v_10621 = v_10616 | v_10620;
assign v_10623 = v_10590 | v_10622;
assign v_10625 = v_10588 | v_10624;
assign v_10627 = v_10622 | v_10626;
assign v_10629 = v_10587 | v_10628;
assign v_10631 = v_10585 | v_10630;
assign v_10633 = v_10628 | v_10632;
assign v_10635 = v_10584 | v_10634;
assign v_10637 = v_10582 | v_10636;
assign v_10639 = v_10634 | v_10638;
assign v_10641 = v_10581 | v_10640;
assign v_10643 = v_10579 | v_10642;
assign v_10645 = v_10640 | v_10644;
assign v_10647 = v_10578 | v_10646;
assign v_10649 = v_10576 | v_10648;
assign v_10651 = v_10646 | v_10650;
assign v_10653 = v_10575 | v_10652;
assign v_10655 = v_10573 | v_10654;
assign v_10657 = v_10652 | v_10656;
assign v_10659 = v_10572 | v_10658;
assign v_10661 = v_10570 | v_10660;
assign v_10663 = v_10658 | v_10662;
assign v_10665 = v_10569 | v_10664;
assign v_10667 = v_10567 | v_10666;
assign v_10669 = v_10664 | v_10668;
assign v_10671 = v_10566 | v_10670;
assign v_10673 = v_10564 | v_10672;
assign v_10675 = v_10670 | v_10674;
assign v_10677 = v_10563 | v_10676;
assign v_10679 = v_10561 | v_10678;
assign v_10681 = v_10676 | v_10680;
assign v_10683 = v_10560 | v_10682;
assign v_10685 = v_10558 | v_10684;
assign v_10687 = v_10682 | v_10686;
assign v_10689 = v_10557 | v_10688;
assign v_10691 = v_10555 | v_10690;
assign v_10693 = v_10688 | v_10692;
assign v_10695 = v_10554 | v_10694;
assign v_10697 = v_10552 | v_10696;
assign v_10699 = v_10694 | v_10698;
assign v_10702 = ~v_10551 | v_10701;
assign v_10709 = v_10599 | v_10708;
assign v_10712 = v_10710 | v_10711;
assign v_10714 = v_10596 | v_10713;
assign v_10717 = v_10715 | v_10716;
assign v_10719 = v_10593 | v_10718;
assign v_10722 = v_10720 | v_10721;
assign v_10724 = v_10590 | v_10723;
assign v_10727 = v_10725 | v_10726;
assign v_10729 = v_10587 | v_10728;
assign v_10732 = v_10730 | v_10731;
assign v_10734 = v_10584 | v_10733;
assign v_10737 = v_10735 | v_10736;
assign v_10739 = v_10581 | v_10738;
assign v_10742 = v_10740 | v_10741;
assign v_10744 = v_10578 | v_10743;
assign v_10747 = v_10745 | v_10746;
assign v_10749 = v_10575 | v_10748;
assign v_10752 = v_10750 | v_10751;
assign v_10754 = v_10572 | v_10753;
assign v_10757 = v_10755 | v_10756;
assign v_10759 = v_10569 | v_10758;
assign v_10762 = v_10760 | v_10761;
assign v_10764 = v_10566 | v_10763;
assign v_10767 = v_10765 | v_10766;
assign v_10769 = v_10563 | v_10768;
assign v_10772 = v_10770 | v_10771;
assign v_10774 = v_10560 | v_10773;
assign v_10777 = v_10775 | v_10776;
assign v_10779 = v_10557 | v_10778;
assign v_10782 = v_10780 | v_10781;
assign v_10784 = v_10554 | v_10783;
assign v_10787 = v_10785 | v_10786;
assign v_10789 = v_10551 | v_10788;
assign v_10792 = v_10550 | v_10791;
assign v_10846 = v_10843 | v_10845;
assign v_10848 = v_10842 | v_10847;
assign v_10850 = v_10840 | v_10849;
assign v_10852 = v_10847 | v_10851;
assign v_10854 = v_10839 | v_10853;
assign v_10856 = v_10837 | v_10855;
assign v_10858 = v_10853 | v_10857;
assign v_10860 = v_10836 | v_10859;
assign v_10862 = v_10834 | v_10861;
assign v_10864 = v_10859 | v_10863;
assign v_10866 = v_10833 | v_10865;
assign v_10868 = v_10831 | v_10867;
assign v_10870 = v_10865 | v_10869;
assign v_10872 = v_10830 | v_10871;
assign v_10874 = v_10828 | v_10873;
assign v_10876 = v_10871 | v_10875;
assign v_10878 = v_10827 | v_10877;
assign v_10880 = v_10825 | v_10879;
assign v_10882 = v_10877 | v_10881;
assign v_10884 = v_10824 | v_10883;
assign v_10886 = v_10822 | v_10885;
assign v_10888 = v_10883 | v_10887;
assign v_10890 = v_10821 | v_10889;
assign v_10892 = v_10819 | v_10891;
assign v_10894 = v_10889 | v_10893;
assign v_10896 = v_10818 | v_10895;
assign v_10898 = v_10816 | v_10897;
assign v_10900 = v_10895 | v_10899;
assign v_10902 = v_10815 | v_10901;
assign v_10904 = v_10813 | v_10903;
assign v_10906 = v_10901 | v_10905;
assign v_10908 = v_10812 | v_10907;
assign v_10910 = v_10810 | v_10909;
assign v_10912 = v_10907 | v_10911;
assign v_10914 = v_10809 | v_10913;
assign v_10916 = v_10807 | v_10915;
assign v_10918 = v_10913 | v_10917;
assign v_10920 = v_10806 | v_10919;
assign v_10922 = v_10804 | v_10921;
assign v_10924 = v_10919 | v_10923;
assign v_10926 = v_10803 | v_10925;
assign v_10928 = v_10801 | v_10927;
assign v_10930 = v_10925 | v_10929;
assign v_10932 = v_10800 | v_10931;
assign v_10934 = v_10798 | v_10933;
assign v_10936 = v_10931 | v_10935;
assign v_10938 = v_10797 | v_10937;
assign v_10940 = v_10795 | v_10939;
assign v_10942 = v_10937 | v_10941;
assign v_10945 = ~v_10794 | v_10944;
assign v_10952 = v_10842 | v_10951;
assign v_10955 = v_10953 | v_10954;
assign v_10957 = v_10839 | v_10956;
assign v_10960 = v_10958 | v_10959;
assign v_10962 = v_10836 | v_10961;
assign v_10965 = v_10963 | v_10964;
assign v_10967 = v_10833 | v_10966;
assign v_10970 = v_10968 | v_10969;
assign v_10972 = v_10830 | v_10971;
assign v_10975 = v_10973 | v_10974;
assign v_10977 = v_10827 | v_10976;
assign v_10980 = v_10978 | v_10979;
assign v_10982 = v_10824 | v_10981;
assign v_10985 = v_10983 | v_10984;
assign v_10987 = v_10821 | v_10986;
assign v_10990 = v_10988 | v_10989;
assign v_10992 = v_10818 | v_10991;
assign v_10995 = v_10993 | v_10994;
assign v_10997 = v_10815 | v_10996;
assign v_11000 = v_10998 | v_10999;
assign v_11002 = v_10812 | v_11001;
assign v_11005 = v_11003 | v_11004;
assign v_11007 = v_10809 | v_11006;
assign v_11010 = v_11008 | v_11009;
assign v_11012 = v_10806 | v_11011;
assign v_11015 = v_11013 | v_11014;
assign v_11017 = v_10803 | v_11016;
assign v_11020 = v_11018 | v_11019;
assign v_11022 = v_10800 | v_11021;
assign v_11025 = v_11023 | v_11024;
assign v_11027 = v_10797 | v_11026;
assign v_11030 = v_11028 | v_11029;
assign v_11032 = v_10794 | v_11031;
assign v_11035 = v_10793 | v_11034;
assign v_11089 = v_11086 | v_11088;
assign v_11091 = v_11085 | v_11090;
assign v_11093 = v_11083 | v_11092;
assign v_11095 = v_11090 | v_11094;
assign v_11097 = v_11082 | v_11096;
assign v_11099 = v_11080 | v_11098;
assign v_11101 = v_11096 | v_11100;
assign v_11103 = v_11079 | v_11102;
assign v_11105 = v_11077 | v_11104;
assign v_11107 = v_11102 | v_11106;
assign v_11109 = v_11076 | v_11108;
assign v_11111 = v_11074 | v_11110;
assign v_11113 = v_11108 | v_11112;
assign v_11115 = v_11073 | v_11114;
assign v_11117 = v_11071 | v_11116;
assign v_11119 = v_11114 | v_11118;
assign v_11121 = v_11070 | v_11120;
assign v_11123 = v_11068 | v_11122;
assign v_11125 = v_11120 | v_11124;
assign v_11127 = v_11067 | v_11126;
assign v_11129 = v_11065 | v_11128;
assign v_11131 = v_11126 | v_11130;
assign v_11133 = v_11064 | v_11132;
assign v_11135 = v_11062 | v_11134;
assign v_11137 = v_11132 | v_11136;
assign v_11139 = v_11061 | v_11138;
assign v_11141 = v_11059 | v_11140;
assign v_11143 = v_11138 | v_11142;
assign v_11145 = v_11058 | v_11144;
assign v_11147 = v_11056 | v_11146;
assign v_11149 = v_11144 | v_11148;
assign v_11151 = v_11055 | v_11150;
assign v_11153 = v_11053 | v_11152;
assign v_11155 = v_11150 | v_11154;
assign v_11157 = v_11052 | v_11156;
assign v_11159 = v_11050 | v_11158;
assign v_11161 = v_11156 | v_11160;
assign v_11163 = v_11049 | v_11162;
assign v_11165 = v_11047 | v_11164;
assign v_11167 = v_11162 | v_11166;
assign v_11169 = v_11046 | v_11168;
assign v_11171 = v_11044 | v_11170;
assign v_11173 = v_11168 | v_11172;
assign v_11175 = v_11043 | v_11174;
assign v_11177 = v_11041 | v_11176;
assign v_11179 = v_11174 | v_11178;
assign v_11181 = v_11040 | v_11180;
assign v_11183 = v_11038 | v_11182;
assign v_11185 = v_11180 | v_11184;
assign v_11188 = ~v_11037 | v_11187;
assign v_11195 = v_11085 | v_11194;
assign v_11198 = v_11196 | v_11197;
assign v_11200 = v_11082 | v_11199;
assign v_11203 = v_11201 | v_11202;
assign v_11205 = v_11079 | v_11204;
assign v_11208 = v_11206 | v_11207;
assign v_11210 = v_11076 | v_11209;
assign v_11213 = v_11211 | v_11212;
assign v_11215 = v_11073 | v_11214;
assign v_11218 = v_11216 | v_11217;
assign v_11220 = v_11070 | v_11219;
assign v_11223 = v_11221 | v_11222;
assign v_11225 = v_11067 | v_11224;
assign v_11228 = v_11226 | v_11227;
assign v_11230 = v_11064 | v_11229;
assign v_11233 = v_11231 | v_11232;
assign v_11235 = v_11061 | v_11234;
assign v_11238 = v_11236 | v_11237;
assign v_11240 = v_11058 | v_11239;
assign v_11243 = v_11241 | v_11242;
assign v_11245 = v_11055 | v_11244;
assign v_11248 = v_11246 | v_11247;
assign v_11250 = v_11052 | v_11249;
assign v_11253 = v_11251 | v_11252;
assign v_11255 = v_11049 | v_11254;
assign v_11258 = v_11256 | v_11257;
assign v_11260 = v_11046 | v_11259;
assign v_11263 = v_11261 | v_11262;
assign v_11265 = v_11043 | v_11264;
assign v_11268 = v_11266 | v_11267;
assign v_11270 = v_11040 | v_11269;
assign v_11273 = v_11271 | v_11272;
assign v_11275 = v_11037 | v_11274;
assign v_11278 = v_11036 | v_11277;
assign v_11332 = v_11329 | v_11331;
assign v_11334 = v_11328 | v_11333;
assign v_11336 = v_11326 | v_11335;
assign v_11338 = v_11333 | v_11337;
assign v_11340 = v_11325 | v_11339;
assign v_11342 = v_11323 | v_11341;
assign v_11344 = v_11339 | v_11343;
assign v_11346 = v_11322 | v_11345;
assign v_11348 = v_11320 | v_11347;
assign v_11350 = v_11345 | v_11349;
assign v_11352 = v_11319 | v_11351;
assign v_11354 = v_11317 | v_11353;
assign v_11356 = v_11351 | v_11355;
assign v_11358 = v_11316 | v_11357;
assign v_11360 = v_11314 | v_11359;
assign v_11362 = v_11357 | v_11361;
assign v_11364 = v_11313 | v_11363;
assign v_11366 = v_11311 | v_11365;
assign v_11368 = v_11363 | v_11367;
assign v_11370 = v_11310 | v_11369;
assign v_11372 = v_11308 | v_11371;
assign v_11374 = v_11369 | v_11373;
assign v_11376 = v_11307 | v_11375;
assign v_11378 = v_11305 | v_11377;
assign v_11380 = v_11375 | v_11379;
assign v_11382 = v_11304 | v_11381;
assign v_11384 = v_11302 | v_11383;
assign v_11386 = v_11381 | v_11385;
assign v_11388 = v_11301 | v_11387;
assign v_11390 = v_11299 | v_11389;
assign v_11392 = v_11387 | v_11391;
assign v_11394 = v_11298 | v_11393;
assign v_11396 = v_11296 | v_11395;
assign v_11398 = v_11393 | v_11397;
assign v_11400 = v_11295 | v_11399;
assign v_11402 = v_11293 | v_11401;
assign v_11404 = v_11399 | v_11403;
assign v_11406 = v_11292 | v_11405;
assign v_11408 = v_11290 | v_11407;
assign v_11410 = v_11405 | v_11409;
assign v_11412 = v_11289 | v_11411;
assign v_11414 = v_11287 | v_11413;
assign v_11416 = v_11411 | v_11415;
assign v_11418 = v_11286 | v_11417;
assign v_11420 = v_11284 | v_11419;
assign v_11422 = v_11417 | v_11421;
assign v_11424 = v_11283 | v_11423;
assign v_11426 = v_11281 | v_11425;
assign v_11428 = v_11423 | v_11427;
assign v_11431 = ~v_11280 | v_11430;
assign v_11438 = v_11328 | v_11437;
assign v_11441 = v_11439 | v_11440;
assign v_11443 = v_11325 | v_11442;
assign v_11446 = v_11444 | v_11445;
assign v_11448 = v_11322 | v_11447;
assign v_11451 = v_11449 | v_11450;
assign v_11453 = v_11319 | v_11452;
assign v_11456 = v_11454 | v_11455;
assign v_11458 = v_11316 | v_11457;
assign v_11461 = v_11459 | v_11460;
assign v_11463 = v_11313 | v_11462;
assign v_11466 = v_11464 | v_11465;
assign v_11468 = v_11310 | v_11467;
assign v_11471 = v_11469 | v_11470;
assign v_11473 = v_11307 | v_11472;
assign v_11476 = v_11474 | v_11475;
assign v_11478 = v_11304 | v_11477;
assign v_11481 = v_11479 | v_11480;
assign v_11483 = v_11301 | v_11482;
assign v_11486 = v_11484 | v_11485;
assign v_11488 = v_11298 | v_11487;
assign v_11491 = v_11489 | v_11490;
assign v_11493 = v_11295 | v_11492;
assign v_11496 = v_11494 | v_11495;
assign v_11498 = v_11292 | v_11497;
assign v_11501 = v_11499 | v_11500;
assign v_11503 = v_11289 | v_11502;
assign v_11506 = v_11504 | v_11505;
assign v_11508 = v_11286 | v_11507;
assign v_11511 = v_11509 | v_11510;
assign v_11513 = v_11283 | v_11512;
assign v_11516 = v_11514 | v_11515;
assign v_11518 = v_11280 | v_11517;
assign v_11521 = v_11279 | v_11520;
assign v_11575 = v_11572 | v_11574;
assign v_11577 = v_11571 | v_11576;
assign v_11579 = v_11569 | v_11578;
assign v_11581 = v_11576 | v_11580;
assign v_11583 = v_11568 | v_11582;
assign v_11585 = v_11566 | v_11584;
assign v_11587 = v_11582 | v_11586;
assign v_11589 = v_11565 | v_11588;
assign v_11591 = v_11563 | v_11590;
assign v_11593 = v_11588 | v_11592;
assign v_11595 = v_11562 | v_11594;
assign v_11597 = v_11560 | v_11596;
assign v_11599 = v_11594 | v_11598;
assign v_11601 = v_11559 | v_11600;
assign v_11603 = v_11557 | v_11602;
assign v_11605 = v_11600 | v_11604;
assign v_11607 = v_11556 | v_11606;
assign v_11609 = v_11554 | v_11608;
assign v_11611 = v_11606 | v_11610;
assign v_11613 = v_11553 | v_11612;
assign v_11615 = v_11551 | v_11614;
assign v_11617 = v_11612 | v_11616;
assign v_11619 = v_11550 | v_11618;
assign v_11621 = v_11548 | v_11620;
assign v_11623 = v_11618 | v_11622;
assign v_11625 = v_11547 | v_11624;
assign v_11627 = v_11545 | v_11626;
assign v_11629 = v_11624 | v_11628;
assign v_11631 = v_11544 | v_11630;
assign v_11633 = v_11542 | v_11632;
assign v_11635 = v_11630 | v_11634;
assign v_11637 = v_11541 | v_11636;
assign v_11639 = v_11539 | v_11638;
assign v_11641 = v_11636 | v_11640;
assign v_11643 = v_11538 | v_11642;
assign v_11645 = v_11536 | v_11644;
assign v_11647 = v_11642 | v_11646;
assign v_11649 = v_11535 | v_11648;
assign v_11651 = v_11533 | v_11650;
assign v_11653 = v_11648 | v_11652;
assign v_11655 = v_11532 | v_11654;
assign v_11657 = v_11530 | v_11656;
assign v_11659 = v_11654 | v_11658;
assign v_11661 = v_11529 | v_11660;
assign v_11663 = v_11527 | v_11662;
assign v_11665 = v_11660 | v_11664;
assign v_11667 = v_11526 | v_11666;
assign v_11669 = v_11524 | v_11668;
assign v_11671 = v_11666 | v_11670;
assign v_11674 = ~v_11523 | v_11673;
assign v_11681 = v_11571 | v_11680;
assign v_11684 = v_11682 | v_11683;
assign v_11686 = v_11568 | v_11685;
assign v_11689 = v_11687 | v_11688;
assign v_11691 = v_11565 | v_11690;
assign v_11694 = v_11692 | v_11693;
assign v_11696 = v_11562 | v_11695;
assign v_11699 = v_11697 | v_11698;
assign v_11701 = v_11559 | v_11700;
assign v_11704 = v_11702 | v_11703;
assign v_11706 = v_11556 | v_11705;
assign v_11709 = v_11707 | v_11708;
assign v_11711 = v_11553 | v_11710;
assign v_11714 = v_11712 | v_11713;
assign v_11716 = v_11550 | v_11715;
assign v_11719 = v_11717 | v_11718;
assign v_11721 = v_11547 | v_11720;
assign v_11724 = v_11722 | v_11723;
assign v_11726 = v_11544 | v_11725;
assign v_11729 = v_11727 | v_11728;
assign v_11731 = v_11541 | v_11730;
assign v_11734 = v_11732 | v_11733;
assign v_11736 = v_11538 | v_11735;
assign v_11739 = v_11737 | v_11738;
assign v_11741 = v_11535 | v_11740;
assign v_11744 = v_11742 | v_11743;
assign v_11746 = v_11532 | v_11745;
assign v_11749 = v_11747 | v_11748;
assign v_11751 = v_11529 | v_11750;
assign v_11754 = v_11752 | v_11753;
assign v_11756 = v_11526 | v_11755;
assign v_11759 = v_11757 | v_11758;
assign v_11761 = v_11523 | v_11760;
assign v_11764 = v_11522 | v_11763;
assign v_11818 = v_11815 | v_11817;
assign v_11820 = v_11814 | v_11819;
assign v_11822 = v_11812 | v_11821;
assign v_11824 = v_11819 | v_11823;
assign v_11826 = v_11811 | v_11825;
assign v_11828 = v_11809 | v_11827;
assign v_11830 = v_11825 | v_11829;
assign v_11832 = v_11808 | v_11831;
assign v_11834 = v_11806 | v_11833;
assign v_11836 = v_11831 | v_11835;
assign v_11838 = v_11805 | v_11837;
assign v_11840 = v_11803 | v_11839;
assign v_11842 = v_11837 | v_11841;
assign v_11844 = v_11802 | v_11843;
assign v_11846 = v_11800 | v_11845;
assign v_11848 = v_11843 | v_11847;
assign v_11850 = v_11799 | v_11849;
assign v_11852 = v_11797 | v_11851;
assign v_11854 = v_11849 | v_11853;
assign v_11856 = v_11796 | v_11855;
assign v_11858 = v_11794 | v_11857;
assign v_11860 = v_11855 | v_11859;
assign v_11862 = v_11793 | v_11861;
assign v_11864 = v_11791 | v_11863;
assign v_11866 = v_11861 | v_11865;
assign v_11868 = v_11790 | v_11867;
assign v_11870 = v_11788 | v_11869;
assign v_11872 = v_11867 | v_11871;
assign v_11874 = v_11787 | v_11873;
assign v_11876 = v_11785 | v_11875;
assign v_11878 = v_11873 | v_11877;
assign v_11880 = v_11784 | v_11879;
assign v_11882 = v_11782 | v_11881;
assign v_11884 = v_11879 | v_11883;
assign v_11886 = v_11781 | v_11885;
assign v_11888 = v_11779 | v_11887;
assign v_11890 = v_11885 | v_11889;
assign v_11892 = v_11778 | v_11891;
assign v_11894 = v_11776 | v_11893;
assign v_11896 = v_11891 | v_11895;
assign v_11898 = v_11775 | v_11897;
assign v_11900 = v_11773 | v_11899;
assign v_11902 = v_11897 | v_11901;
assign v_11904 = v_11772 | v_11903;
assign v_11906 = v_11770 | v_11905;
assign v_11908 = v_11903 | v_11907;
assign v_11910 = v_11769 | v_11909;
assign v_11912 = v_11767 | v_11911;
assign v_11914 = v_11909 | v_11913;
assign v_11917 = ~v_11766 | v_11916;
assign v_11924 = v_11814 | v_11923;
assign v_11927 = v_11925 | v_11926;
assign v_11929 = v_11811 | v_11928;
assign v_11932 = v_11930 | v_11931;
assign v_11934 = v_11808 | v_11933;
assign v_11937 = v_11935 | v_11936;
assign v_11939 = v_11805 | v_11938;
assign v_11942 = v_11940 | v_11941;
assign v_11944 = v_11802 | v_11943;
assign v_11947 = v_11945 | v_11946;
assign v_11949 = v_11799 | v_11948;
assign v_11952 = v_11950 | v_11951;
assign v_11954 = v_11796 | v_11953;
assign v_11957 = v_11955 | v_11956;
assign v_11959 = v_11793 | v_11958;
assign v_11962 = v_11960 | v_11961;
assign v_11964 = v_11790 | v_11963;
assign v_11967 = v_11965 | v_11966;
assign v_11969 = v_11787 | v_11968;
assign v_11972 = v_11970 | v_11971;
assign v_11974 = v_11784 | v_11973;
assign v_11977 = v_11975 | v_11976;
assign v_11979 = v_11781 | v_11978;
assign v_11982 = v_11980 | v_11981;
assign v_11984 = v_11778 | v_11983;
assign v_11987 = v_11985 | v_11986;
assign v_11989 = v_11775 | v_11988;
assign v_11992 = v_11990 | v_11991;
assign v_11994 = v_11772 | v_11993;
assign v_11997 = v_11995 | v_11996;
assign v_11999 = v_11769 | v_11998;
assign v_12002 = v_12000 | v_12001;
assign v_12004 = v_11766 | v_12003;
assign v_12007 = v_11765 | v_12006;
assign v_12061 = v_12058 | v_12060;
assign v_12063 = v_12057 | v_12062;
assign v_12065 = v_12055 | v_12064;
assign v_12067 = v_12062 | v_12066;
assign v_12069 = v_12054 | v_12068;
assign v_12071 = v_12052 | v_12070;
assign v_12073 = v_12068 | v_12072;
assign v_12075 = v_12051 | v_12074;
assign v_12077 = v_12049 | v_12076;
assign v_12079 = v_12074 | v_12078;
assign v_12081 = v_12048 | v_12080;
assign v_12083 = v_12046 | v_12082;
assign v_12085 = v_12080 | v_12084;
assign v_12087 = v_12045 | v_12086;
assign v_12089 = v_12043 | v_12088;
assign v_12091 = v_12086 | v_12090;
assign v_12093 = v_12042 | v_12092;
assign v_12095 = v_12040 | v_12094;
assign v_12097 = v_12092 | v_12096;
assign v_12099 = v_12039 | v_12098;
assign v_12101 = v_12037 | v_12100;
assign v_12103 = v_12098 | v_12102;
assign v_12105 = v_12036 | v_12104;
assign v_12107 = v_12034 | v_12106;
assign v_12109 = v_12104 | v_12108;
assign v_12111 = v_12033 | v_12110;
assign v_12113 = v_12031 | v_12112;
assign v_12115 = v_12110 | v_12114;
assign v_12117 = v_12030 | v_12116;
assign v_12119 = v_12028 | v_12118;
assign v_12121 = v_12116 | v_12120;
assign v_12123 = v_12027 | v_12122;
assign v_12125 = v_12025 | v_12124;
assign v_12127 = v_12122 | v_12126;
assign v_12129 = v_12024 | v_12128;
assign v_12131 = v_12022 | v_12130;
assign v_12133 = v_12128 | v_12132;
assign v_12135 = v_12021 | v_12134;
assign v_12137 = v_12019 | v_12136;
assign v_12139 = v_12134 | v_12138;
assign v_12141 = v_12018 | v_12140;
assign v_12143 = v_12016 | v_12142;
assign v_12145 = v_12140 | v_12144;
assign v_12147 = v_12015 | v_12146;
assign v_12149 = v_12013 | v_12148;
assign v_12151 = v_12146 | v_12150;
assign v_12153 = v_12012 | v_12152;
assign v_12155 = v_12010 | v_12154;
assign v_12157 = v_12152 | v_12156;
assign v_12160 = ~v_12009 | v_12159;
assign v_12167 = v_12057 | v_12166;
assign v_12170 = v_12168 | v_12169;
assign v_12172 = v_12054 | v_12171;
assign v_12175 = v_12173 | v_12174;
assign v_12177 = v_12051 | v_12176;
assign v_12180 = v_12178 | v_12179;
assign v_12182 = v_12048 | v_12181;
assign v_12185 = v_12183 | v_12184;
assign v_12187 = v_12045 | v_12186;
assign v_12190 = v_12188 | v_12189;
assign v_12192 = v_12042 | v_12191;
assign v_12195 = v_12193 | v_12194;
assign v_12197 = v_12039 | v_12196;
assign v_12200 = v_12198 | v_12199;
assign v_12202 = v_12036 | v_12201;
assign v_12205 = v_12203 | v_12204;
assign v_12207 = v_12033 | v_12206;
assign v_12210 = v_12208 | v_12209;
assign v_12212 = v_12030 | v_12211;
assign v_12215 = v_12213 | v_12214;
assign v_12217 = v_12027 | v_12216;
assign v_12220 = v_12218 | v_12219;
assign v_12222 = v_12024 | v_12221;
assign v_12225 = v_12223 | v_12224;
assign v_12227 = v_12021 | v_12226;
assign v_12230 = v_12228 | v_12229;
assign v_12232 = v_12018 | v_12231;
assign v_12235 = v_12233 | v_12234;
assign v_12237 = v_12015 | v_12236;
assign v_12240 = v_12238 | v_12239;
assign v_12242 = v_12012 | v_12241;
assign v_12245 = v_12243 | v_12244;
assign v_12247 = v_12009 | v_12246;
assign v_12250 = v_12008 | v_12249;
assign v_12304 = v_12301 | v_12303;
assign v_12306 = v_12300 | v_12305;
assign v_12308 = v_12298 | v_12307;
assign v_12310 = v_12305 | v_12309;
assign v_12312 = v_12297 | v_12311;
assign v_12314 = v_12295 | v_12313;
assign v_12316 = v_12311 | v_12315;
assign v_12318 = v_12294 | v_12317;
assign v_12320 = v_12292 | v_12319;
assign v_12322 = v_12317 | v_12321;
assign v_12324 = v_12291 | v_12323;
assign v_12326 = v_12289 | v_12325;
assign v_12328 = v_12323 | v_12327;
assign v_12330 = v_12288 | v_12329;
assign v_12332 = v_12286 | v_12331;
assign v_12334 = v_12329 | v_12333;
assign v_12336 = v_12285 | v_12335;
assign v_12338 = v_12283 | v_12337;
assign v_12340 = v_12335 | v_12339;
assign v_12342 = v_12282 | v_12341;
assign v_12344 = v_12280 | v_12343;
assign v_12346 = v_12341 | v_12345;
assign v_12348 = v_12279 | v_12347;
assign v_12350 = v_12277 | v_12349;
assign v_12352 = v_12347 | v_12351;
assign v_12354 = v_12276 | v_12353;
assign v_12356 = v_12274 | v_12355;
assign v_12358 = v_12353 | v_12357;
assign v_12360 = v_12273 | v_12359;
assign v_12362 = v_12271 | v_12361;
assign v_12364 = v_12359 | v_12363;
assign v_12366 = v_12270 | v_12365;
assign v_12368 = v_12268 | v_12367;
assign v_12370 = v_12365 | v_12369;
assign v_12372 = v_12267 | v_12371;
assign v_12374 = v_12265 | v_12373;
assign v_12376 = v_12371 | v_12375;
assign v_12378 = v_12264 | v_12377;
assign v_12380 = v_12262 | v_12379;
assign v_12382 = v_12377 | v_12381;
assign v_12384 = v_12261 | v_12383;
assign v_12386 = v_12259 | v_12385;
assign v_12388 = v_12383 | v_12387;
assign v_12390 = v_12258 | v_12389;
assign v_12392 = v_12256 | v_12391;
assign v_12394 = v_12389 | v_12393;
assign v_12396 = v_12255 | v_12395;
assign v_12398 = v_12253 | v_12397;
assign v_12400 = v_12395 | v_12399;
assign v_12403 = ~v_12252 | v_12402;
assign v_12410 = v_12300 | v_12409;
assign v_12413 = v_12411 | v_12412;
assign v_12415 = v_12297 | v_12414;
assign v_12418 = v_12416 | v_12417;
assign v_12420 = v_12294 | v_12419;
assign v_12423 = v_12421 | v_12422;
assign v_12425 = v_12291 | v_12424;
assign v_12428 = v_12426 | v_12427;
assign v_12430 = v_12288 | v_12429;
assign v_12433 = v_12431 | v_12432;
assign v_12435 = v_12285 | v_12434;
assign v_12438 = v_12436 | v_12437;
assign v_12440 = v_12282 | v_12439;
assign v_12443 = v_12441 | v_12442;
assign v_12445 = v_12279 | v_12444;
assign v_12448 = v_12446 | v_12447;
assign v_12450 = v_12276 | v_12449;
assign v_12453 = v_12451 | v_12452;
assign v_12455 = v_12273 | v_12454;
assign v_12458 = v_12456 | v_12457;
assign v_12460 = v_12270 | v_12459;
assign v_12463 = v_12461 | v_12462;
assign v_12465 = v_12267 | v_12464;
assign v_12468 = v_12466 | v_12467;
assign v_12470 = v_12264 | v_12469;
assign v_12473 = v_12471 | v_12472;
assign v_12475 = v_12261 | v_12474;
assign v_12478 = v_12476 | v_12477;
assign v_12480 = v_12258 | v_12479;
assign v_12483 = v_12481 | v_12482;
assign v_12485 = v_12255 | v_12484;
assign v_12488 = v_12486 | v_12487;
assign v_12490 = v_12252 | v_12489;
assign v_12493 = v_12251 | v_12492;
assign v_12546 = v_12543 | v_12545;
assign v_12548 = v_12542 | v_12547;
assign v_12550 = v_12540 | v_12549;
assign v_12552 = v_12547 | v_12551;
assign v_12554 = v_12539 | v_12553;
assign v_12556 = v_12537 | v_12555;
assign v_12558 = v_12553 | v_12557;
assign v_12560 = v_12536 | v_12559;
assign v_12562 = v_12534 | v_12561;
assign v_12564 = v_12559 | v_12563;
assign v_12566 = v_12533 | v_12565;
assign v_12568 = v_12531 | v_12567;
assign v_12570 = v_12565 | v_12569;
assign v_12572 = v_12530 | v_12571;
assign v_12574 = v_12528 | v_12573;
assign v_12576 = v_12571 | v_12575;
assign v_12578 = v_12527 | v_12577;
assign v_12580 = v_12525 | v_12579;
assign v_12582 = v_12577 | v_12581;
assign v_12584 = v_12524 | v_12583;
assign v_12586 = v_12522 | v_12585;
assign v_12588 = v_12583 | v_12587;
assign v_12590 = v_12521 | v_12589;
assign v_12592 = v_12519 | v_12591;
assign v_12594 = v_12589 | v_12593;
assign v_12596 = v_12518 | v_12595;
assign v_12598 = v_12516 | v_12597;
assign v_12600 = v_12595 | v_12599;
assign v_12602 = v_12515 | v_12601;
assign v_12604 = v_12513 | v_12603;
assign v_12606 = v_12601 | v_12605;
assign v_12608 = v_12512 | v_12607;
assign v_12610 = v_12510 | v_12609;
assign v_12612 = v_12607 | v_12611;
assign v_12614 = v_12509 | v_12613;
assign v_12616 = v_12507 | v_12615;
assign v_12618 = v_12613 | v_12617;
assign v_12620 = v_12506 | v_12619;
assign v_12622 = v_12504 | v_12621;
assign v_12624 = v_12619 | v_12623;
assign v_12626 = v_12503 | v_12625;
assign v_12628 = v_12501 | v_12627;
assign v_12630 = v_12625 | v_12629;
assign v_12632 = v_12500 | v_12631;
assign v_12634 = v_12498 | v_12633;
assign v_12636 = v_12631 | v_12635;
assign v_12638 = v_12497 | v_12637;
assign v_12640 = v_12495 | v_12639;
assign v_12642 = v_12637 | v_12641;
assign v_12646 = v_12643 | v_12645;
assign v_12653 = v_12542 | v_12652;
assign v_12656 = v_12654 | v_12655;
assign v_12658 = v_12539 | v_12657;
assign v_12661 = v_12659 | v_12660;
assign v_12663 = v_12536 | v_12662;
assign v_12666 = v_12664 | v_12665;
assign v_12668 = v_12533 | v_12667;
assign v_12671 = v_12669 | v_12670;
assign v_12673 = v_12530 | v_12672;
assign v_12676 = v_12674 | v_12675;
assign v_12678 = v_12527 | v_12677;
assign v_12681 = v_12679 | v_12680;
assign v_12683 = v_12524 | v_12682;
assign v_12686 = v_12684 | v_12685;
assign v_12688 = v_12521 | v_12687;
assign v_12691 = v_12689 | v_12690;
assign v_12693 = v_12518 | v_12692;
assign v_12696 = v_12694 | v_12695;
assign v_12698 = v_12515 | v_12697;
assign v_12701 = v_12699 | v_12700;
assign v_12703 = v_12512 | v_12702;
assign v_12706 = v_12704 | v_12705;
assign v_12708 = v_12509 | v_12707;
assign v_12711 = v_12709 | v_12710;
assign v_12713 = v_12506 | v_12712;
assign v_12716 = v_12714 | v_12715;
assign v_12718 = v_12503 | v_12717;
assign v_12721 = v_12719 | v_12720;
assign v_12723 = v_12500 | v_12722;
assign v_12726 = v_12724 | v_12725;
assign v_12728 = v_12497 | v_12727;
assign v_12731 = v_12729 | v_12730;
assign v_12733 = v_12731 | v_12732;
assign v_12736 = v_12494 | v_12735;
assign v_12807 = v_12804 | v_12806;
assign v_12809 = v_12802 | v_12808;
assign v_12811 = v_12800 | v_12810;
assign v_12813 = v_12808 | v_12812;
assign v_12815 = v_12798 | v_12814;
assign v_12817 = v_12796 | v_12816;
assign v_12819 = v_12814 | v_12818;
assign v_12821 = v_12794 | v_12820;
assign v_12823 = v_12792 | v_12822;
assign v_12825 = v_12820 | v_12824;
assign v_12827 = v_12790 | v_12826;
assign v_12829 = v_12788 | v_12828;
assign v_12831 = v_12826 | v_12830;
assign v_12833 = v_12786 | v_12832;
assign v_12835 = v_12784 | v_12834;
assign v_12837 = v_12832 | v_12836;
assign v_12839 = v_12782 | v_12838;
assign v_12841 = v_12780 | v_12840;
assign v_12843 = v_12838 | v_12842;
assign v_12845 = v_12778 | v_12844;
assign v_12847 = v_12776 | v_12846;
assign v_12849 = v_12844 | v_12848;
assign v_12851 = v_12774 | v_12850;
assign v_12853 = v_12772 | v_12852;
assign v_12855 = v_12850 | v_12854;
assign v_12857 = v_12770 | v_12856;
assign v_12859 = v_12768 | v_12858;
assign v_12861 = v_12856 | v_12860;
assign v_12863 = v_12766 | v_12862;
assign v_12865 = v_12764 | v_12864;
assign v_12867 = v_12862 | v_12866;
assign v_12869 = v_12762 | v_12868;
assign v_12871 = v_12760 | v_12870;
assign v_12873 = v_12868 | v_12872;
assign v_12875 = v_12758 | v_12874;
assign v_12877 = v_12756 | v_12876;
assign v_12879 = v_12874 | v_12878;
assign v_12881 = v_12754 | v_12880;
assign v_12883 = v_12751 | v_12882;
assign v_12885 = v_12880 | v_12884;
assign v_12887 = v_12750 | v_12886;
assign v_12889 = v_12747 | v_12888;
assign v_12891 = v_12886 | v_12890;
assign v_12893 = v_12746 | v_12892;
assign v_12895 = v_12743 | v_12894;
assign v_12897 = v_12892 | v_12896;
assign v_12899 = v_12742 | v_12898;
assign v_12901 = v_12739 | v_12900;
assign v_12903 = v_12898 | v_12902;
assign v_12906 = ~v_12738 | v_12905;
assign v_12913 = v_12802 | v_12912;
assign v_12916 = v_12914 | v_12915;
assign v_12918 = v_12798 | v_12917;
assign v_12921 = v_12919 | v_12920;
assign v_12923 = v_12794 | v_12922;
assign v_12926 = v_12924 | v_12925;
assign v_12928 = v_12790 | v_12927;
assign v_12931 = v_12929 | v_12930;
assign v_12933 = v_12786 | v_12932;
assign v_12936 = v_12934 | v_12935;
assign v_12938 = v_12782 | v_12937;
assign v_12941 = v_12939 | v_12940;
assign v_12943 = v_12778 | v_12942;
assign v_12946 = v_12944 | v_12945;
assign v_12948 = v_12774 | v_12947;
assign v_12951 = v_12949 | v_12950;
assign v_12953 = v_12770 | v_12952;
assign v_12956 = v_12954 | v_12955;
assign v_12958 = v_12766 | v_12957;
assign v_12961 = v_12959 | v_12960;
assign v_12963 = v_12762 | v_12962;
assign v_12966 = v_12964 | v_12965;
assign v_12968 = v_12758 | v_12967;
assign v_12971 = v_12969 | v_12970;
assign v_12973 = v_12754 | v_12972;
assign v_12976 = v_12974 | v_12975;
assign v_12978 = v_12750 | v_12977;
assign v_12981 = v_12979 | v_12980;
assign v_12983 = v_12746 | v_12982;
assign v_12986 = v_12984 | v_12985;
assign v_12988 = v_12742 | v_12987;
assign v_12991 = v_12989 | v_12990;
assign v_12993 = v_12738 | v_12992;
assign v_12996 = v_12737 | v_12995;
assign v_13050 = v_13047 | v_13049;
assign v_13052 = v_13046 | v_13051;
assign v_13054 = v_13044 | v_13053;
assign v_13056 = v_13051 | v_13055;
assign v_13058 = v_13043 | v_13057;
assign v_13060 = v_13041 | v_13059;
assign v_13062 = v_13057 | v_13061;
assign v_13064 = v_13040 | v_13063;
assign v_13066 = v_13038 | v_13065;
assign v_13068 = v_13063 | v_13067;
assign v_13070 = v_13037 | v_13069;
assign v_13072 = v_13035 | v_13071;
assign v_13074 = v_13069 | v_13073;
assign v_13076 = v_13034 | v_13075;
assign v_13078 = v_13032 | v_13077;
assign v_13080 = v_13075 | v_13079;
assign v_13082 = v_13031 | v_13081;
assign v_13084 = v_13029 | v_13083;
assign v_13086 = v_13081 | v_13085;
assign v_13088 = v_13028 | v_13087;
assign v_13090 = v_13026 | v_13089;
assign v_13092 = v_13087 | v_13091;
assign v_13094 = v_13025 | v_13093;
assign v_13096 = v_13023 | v_13095;
assign v_13098 = v_13093 | v_13097;
assign v_13100 = v_13022 | v_13099;
assign v_13102 = v_13020 | v_13101;
assign v_13104 = v_13099 | v_13103;
assign v_13106 = v_13019 | v_13105;
assign v_13108 = v_13017 | v_13107;
assign v_13110 = v_13105 | v_13109;
assign v_13112 = v_13016 | v_13111;
assign v_13114 = v_13014 | v_13113;
assign v_13116 = v_13111 | v_13115;
assign v_13118 = v_13013 | v_13117;
assign v_13120 = v_13011 | v_13119;
assign v_13122 = v_13117 | v_13121;
assign v_13124 = v_13010 | v_13123;
assign v_13126 = v_13008 | v_13125;
assign v_13128 = v_13123 | v_13127;
assign v_13130 = v_13007 | v_13129;
assign v_13132 = v_13005 | v_13131;
assign v_13134 = v_13129 | v_13133;
assign v_13136 = v_13004 | v_13135;
assign v_13138 = v_13002 | v_13137;
assign v_13140 = v_13135 | v_13139;
assign v_13142 = v_13001 | v_13141;
assign v_13144 = v_12999 | v_13143;
assign v_13146 = v_13141 | v_13145;
assign v_13149 = ~v_12998 | v_13148;
assign v_13156 = v_13046 | v_13155;
assign v_13159 = v_13157 | v_13158;
assign v_13161 = v_13043 | v_13160;
assign v_13164 = v_13162 | v_13163;
assign v_13166 = v_13040 | v_13165;
assign v_13169 = v_13167 | v_13168;
assign v_13171 = v_13037 | v_13170;
assign v_13174 = v_13172 | v_13173;
assign v_13176 = v_13034 | v_13175;
assign v_13179 = v_13177 | v_13178;
assign v_13181 = v_13031 | v_13180;
assign v_13184 = v_13182 | v_13183;
assign v_13186 = v_13028 | v_13185;
assign v_13189 = v_13187 | v_13188;
assign v_13191 = v_13025 | v_13190;
assign v_13194 = v_13192 | v_13193;
assign v_13196 = v_13022 | v_13195;
assign v_13199 = v_13197 | v_13198;
assign v_13201 = v_13019 | v_13200;
assign v_13204 = v_13202 | v_13203;
assign v_13206 = v_13016 | v_13205;
assign v_13209 = v_13207 | v_13208;
assign v_13211 = v_13013 | v_13210;
assign v_13214 = v_13212 | v_13213;
assign v_13216 = v_13010 | v_13215;
assign v_13219 = v_13217 | v_13218;
assign v_13221 = v_13007 | v_13220;
assign v_13224 = v_13222 | v_13223;
assign v_13226 = v_13004 | v_13225;
assign v_13229 = v_13227 | v_13228;
assign v_13231 = v_13001 | v_13230;
assign v_13234 = v_13232 | v_13233;
assign v_13236 = v_12998 | v_13235;
assign v_13239 = v_12997 | v_13238;
assign v_13293 = v_13290 | v_13292;
assign v_13295 = v_13289 | v_13294;
assign v_13297 = v_13287 | v_13296;
assign v_13299 = v_13294 | v_13298;
assign v_13301 = v_13286 | v_13300;
assign v_13303 = v_13284 | v_13302;
assign v_13305 = v_13300 | v_13304;
assign v_13307 = v_13283 | v_13306;
assign v_13309 = v_13281 | v_13308;
assign v_13311 = v_13306 | v_13310;
assign v_13313 = v_13280 | v_13312;
assign v_13315 = v_13278 | v_13314;
assign v_13317 = v_13312 | v_13316;
assign v_13319 = v_13277 | v_13318;
assign v_13321 = v_13275 | v_13320;
assign v_13323 = v_13318 | v_13322;
assign v_13325 = v_13274 | v_13324;
assign v_13327 = v_13272 | v_13326;
assign v_13329 = v_13324 | v_13328;
assign v_13331 = v_13271 | v_13330;
assign v_13333 = v_13269 | v_13332;
assign v_13335 = v_13330 | v_13334;
assign v_13337 = v_13268 | v_13336;
assign v_13339 = v_13266 | v_13338;
assign v_13341 = v_13336 | v_13340;
assign v_13343 = v_13265 | v_13342;
assign v_13345 = v_13263 | v_13344;
assign v_13347 = v_13342 | v_13346;
assign v_13349 = v_13262 | v_13348;
assign v_13351 = v_13260 | v_13350;
assign v_13353 = v_13348 | v_13352;
assign v_13355 = v_13259 | v_13354;
assign v_13357 = v_13257 | v_13356;
assign v_13359 = v_13354 | v_13358;
assign v_13361 = v_13256 | v_13360;
assign v_13363 = v_13254 | v_13362;
assign v_13365 = v_13360 | v_13364;
assign v_13367 = v_13253 | v_13366;
assign v_13369 = v_13251 | v_13368;
assign v_13371 = v_13366 | v_13370;
assign v_13373 = v_13250 | v_13372;
assign v_13375 = v_13248 | v_13374;
assign v_13377 = v_13372 | v_13376;
assign v_13379 = v_13247 | v_13378;
assign v_13381 = v_13245 | v_13380;
assign v_13383 = v_13378 | v_13382;
assign v_13385 = v_13244 | v_13384;
assign v_13387 = v_13242 | v_13386;
assign v_13389 = v_13384 | v_13388;
assign v_13392 = ~v_13241 | v_13391;
assign v_13399 = v_13289 | v_13398;
assign v_13402 = v_13400 | v_13401;
assign v_13404 = v_13286 | v_13403;
assign v_13407 = v_13405 | v_13406;
assign v_13409 = v_13283 | v_13408;
assign v_13412 = v_13410 | v_13411;
assign v_13414 = v_13280 | v_13413;
assign v_13417 = v_13415 | v_13416;
assign v_13419 = v_13277 | v_13418;
assign v_13422 = v_13420 | v_13421;
assign v_13424 = v_13274 | v_13423;
assign v_13427 = v_13425 | v_13426;
assign v_13429 = v_13271 | v_13428;
assign v_13432 = v_13430 | v_13431;
assign v_13434 = v_13268 | v_13433;
assign v_13437 = v_13435 | v_13436;
assign v_13439 = v_13265 | v_13438;
assign v_13442 = v_13440 | v_13441;
assign v_13444 = v_13262 | v_13443;
assign v_13447 = v_13445 | v_13446;
assign v_13449 = v_13259 | v_13448;
assign v_13452 = v_13450 | v_13451;
assign v_13454 = v_13256 | v_13453;
assign v_13457 = v_13455 | v_13456;
assign v_13459 = v_13253 | v_13458;
assign v_13462 = v_13460 | v_13461;
assign v_13464 = v_13250 | v_13463;
assign v_13467 = v_13465 | v_13466;
assign v_13469 = v_13247 | v_13468;
assign v_13472 = v_13470 | v_13471;
assign v_13474 = v_13244 | v_13473;
assign v_13477 = v_13475 | v_13476;
assign v_13479 = v_13241 | v_13478;
assign v_13482 = v_13240 | v_13481;
assign v_13536 = v_13533 | v_13535;
assign v_13538 = v_13532 | v_13537;
assign v_13540 = v_13530 | v_13539;
assign v_13542 = v_13537 | v_13541;
assign v_13544 = v_13529 | v_13543;
assign v_13546 = v_13527 | v_13545;
assign v_13548 = v_13543 | v_13547;
assign v_13550 = v_13526 | v_13549;
assign v_13552 = v_13524 | v_13551;
assign v_13554 = v_13549 | v_13553;
assign v_13556 = v_13523 | v_13555;
assign v_13558 = v_13521 | v_13557;
assign v_13560 = v_13555 | v_13559;
assign v_13562 = v_13520 | v_13561;
assign v_13564 = v_13518 | v_13563;
assign v_13566 = v_13561 | v_13565;
assign v_13568 = v_13517 | v_13567;
assign v_13570 = v_13515 | v_13569;
assign v_13572 = v_13567 | v_13571;
assign v_13574 = v_13514 | v_13573;
assign v_13576 = v_13512 | v_13575;
assign v_13578 = v_13573 | v_13577;
assign v_13580 = v_13511 | v_13579;
assign v_13582 = v_13509 | v_13581;
assign v_13584 = v_13579 | v_13583;
assign v_13586 = v_13508 | v_13585;
assign v_13588 = v_13506 | v_13587;
assign v_13590 = v_13585 | v_13589;
assign v_13592 = v_13505 | v_13591;
assign v_13594 = v_13503 | v_13593;
assign v_13596 = v_13591 | v_13595;
assign v_13598 = v_13502 | v_13597;
assign v_13600 = v_13500 | v_13599;
assign v_13602 = v_13597 | v_13601;
assign v_13604 = v_13499 | v_13603;
assign v_13606 = v_13497 | v_13605;
assign v_13608 = v_13603 | v_13607;
assign v_13610 = v_13496 | v_13609;
assign v_13612 = v_13494 | v_13611;
assign v_13614 = v_13609 | v_13613;
assign v_13616 = v_13493 | v_13615;
assign v_13618 = v_13491 | v_13617;
assign v_13620 = v_13615 | v_13619;
assign v_13622 = v_13490 | v_13621;
assign v_13624 = v_13488 | v_13623;
assign v_13626 = v_13621 | v_13625;
assign v_13628 = v_13487 | v_13627;
assign v_13630 = v_13485 | v_13629;
assign v_13632 = v_13627 | v_13631;
assign v_13635 = ~v_13484 | v_13634;
assign v_13642 = v_13532 | v_13641;
assign v_13645 = v_13643 | v_13644;
assign v_13647 = v_13529 | v_13646;
assign v_13650 = v_13648 | v_13649;
assign v_13652 = v_13526 | v_13651;
assign v_13655 = v_13653 | v_13654;
assign v_13657 = v_13523 | v_13656;
assign v_13660 = v_13658 | v_13659;
assign v_13662 = v_13520 | v_13661;
assign v_13665 = v_13663 | v_13664;
assign v_13667 = v_13517 | v_13666;
assign v_13670 = v_13668 | v_13669;
assign v_13672 = v_13514 | v_13671;
assign v_13675 = v_13673 | v_13674;
assign v_13677 = v_13511 | v_13676;
assign v_13680 = v_13678 | v_13679;
assign v_13682 = v_13508 | v_13681;
assign v_13685 = v_13683 | v_13684;
assign v_13687 = v_13505 | v_13686;
assign v_13690 = v_13688 | v_13689;
assign v_13692 = v_13502 | v_13691;
assign v_13695 = v_13693 | v_13694;
assign v_13697 = v_13499 | v_13696;
assign v_13700 = v_13698 | v_13699;
assign v_13702 = v_13496 | v_13701;
assign v_13705 = v_13703 | v_13704;
assign v_13707 = v_13493 | v_13706;
assign v_13710 = v_13708 | v_13709;
assign v_13712 = v_13490 | v_13711;
assign v_13715 = v_13713 | v_13714;
assign v_13717 = v_13487 | v_13716;
assign v_13720 = v_13718 | v_13719;
assign v_13722 = v_13484 | v_13721;
assign v_13725 = v_13483 | v_13724;
assign v_13779 = v_13776 | v_13778;
assign v_13781 = v_13775 | v_13780;
assign v_13783 = v_13773 | v_13782;
assign v_13785 = v_13780 | v_13784;
assign v_13787 = v_13772 | v_13786;
assign v_13789 = v_13770 | v_13788;
assign v_13791 = v_13786 | v_13790;
assign v_13793 = v_13769 | v_13792;
assign v_13795 = v_13767 | v_13794;
assign v_13797 = v_13792 | v_13796;
assign v_13799 = v_13766 | v_13798;
assign v_13801 = v_13764 | v_13800;
assign v_13803 = v_13798 | v_13802;
assign v_13805 = v_13763 | v_13804;
assign v_13807 = v_13761 | v_13806;
assign v_13809 = v_13804 | v_13808;
assign v_13811 = v_13760 | v_13810;
assign v_13813 = v_13758 | v_13812;
assign v_13815 = v_13810 | v_13814;
assign v_13817 = v_13757 | v_13816;
assign v_13819 = v_13755 | v_13818;
assign v_13821 = v_13816 | v_13820;
assign v_13823 = v_13754 | v_13822;
assign v_13825 = v_13752 | v_13824;
assign v_13827 = v_13822 | v_13826;
assign v_13829 = v_13751 | v_13828;
assign v_13831 = v_13749 | v_13830;
assign v_13833 = v_13828 | v_13832;
assign v_13835 = v_13748 | v_13834;
assign v_13837 = v_13746 | v_13836;
assign v_13839 = v_13834 | v_13838;
assign v_13841 = v_13745 | v_13840;
assign v_13843 = v_13743 | v_13842;
assign v_13845 = v_13840 | v_13844;
assign v_13847 = v_13742 | v_13846;
assign v_13849 = v_13740 | v_13848;
assign v_13851 = v_13846 | v_13850;
assign v_13853 = v_13739 | v_13852;
assign v_13855 = v_13737 | v_13854;
assign v_13857 = v_13852 | v_13856;
assign v_13859 = v_13736 | v_13858;
assign v_13861 = v_13734 | v_13860;
assign v_13863 = v_13858 | v_13862;
assign v_13865 = v_13733 | v_13864;
assign v_13867 = v_13731 | v_13866;
assign v_13869 = v_13864 | v_13868;
assign v_13871 = v_13730 | v_13870;
assign v_13873 = v_13728 | v_13872;
assign v_13875 = v_13870 | v_13874;
assign v_13878 = ~v_13727 | v_13877;
assign v_13885 = v_13775 | v_13884;
assign v_13888 = v_13886 | v_13887;
assign v_13890 = v_13772 | v_13889;
assign v_13893 = v_13891 | v_13892;
assign v_13895 = v_13769 | v_13894;
assign v_13898 = v_13896 | v_13897;
assign v_13900 = v_13766 | v_13899;
assign v_13903 = v_13901 | v_13902;
assign v_13905 = v_13763 | v_13904;
assign v_13908 = v_13906 | v_13907;
assign v_13910 = v_13760 | v_13909;
assign v_13913 = v_13911 | v_13912;
assign v_13915 = v_13757 | v_13914;
assign v_13918 = v_13916 | v_13917;
assign v_13920 = v_13754 | v_13919;
assign v_13923 = v_13921 | v_13922;
assign v_13925 = v_13751 | v_13924;
assign v_13928 = v_13926 | v_13927;
assign v_13930 = v_13748 | v_13929;
assign v_13933 = v_13931 | v_13932;
assign v_13935 = v_13745 | v_13934;
assign v_13938 = v_13936 | v_13937;
assign v_13940 = v_13742 | v_13939;
assign v_13943 = v_13941 | v_13942;
assign v_13945 = v_13739 | v_13944;
assign v_13948 = v_13946 | v_13947;
assign v_13950 = v_13736 | v_13949;
assign v_13953 = v_13951 | v_13952;
assign v_13955 = v_13733 | v_13954;
assign v_13958 = v_13956 | v_13957;
assign v_13960 = v_13730 | v_13959;
assign v_13963 = v_13961 | v_13962;
assign v_13965 = v_13727 | v_13964;
assign v_13968 = v_13726 | v_13967;
assign v_14022 = v_14019 | v_14021;
assign v_14024 = v_14018 | v_14023;
assign v_14026 = v_14016 | v_14025;
assign v_14028 = v_14023 | v_14027;
assign v_14030 = v_14015 | v_14029;
assign v_14032 = v_14013 | v_14031;
assign v_14034 = v_14029 | v_14033;
assign v_14036 = v_14012 | v_14035;
assign v_14038 = v_14010 | v_14037;
assign v_14040 = v_14035 | v_14039;
assign v_14042 = v_14009 | v_14041;
assign v_14044 = v_14007 | v_14043;
assign v_14046 = v_14041 | v_14045;
assign v_14048 = v_14006 | v_14047;
assign v_14050 = v_14004 | v_14049;
assign v_14052 = v_14047 | v_14051;
assign v_14054 = v_14003 | v_14053;
assign v_14056 = v_14001 | v_14055;
assign v_14058 = v_14053 | v_14057;
assign v_14060 = v_14000 | v_14059;
assign v_14062 = v_13998 | v_14061;
assign v_14064 = v_14059 | v_14063;
assign v_14066 = v_13997 | v_14065;
assign v_14068 = v_13995 | v_14067;
assign v_14070 = v_14065 | v_14069;
assign v_14072 = v_13994 | v_14071;
assign v_14074 = v_13992 | v_14073;
assign v_14076 = v_14071 | v_14075;
assign v_14078 = v_13991 | v_14077;
assign v_14080 = v_13989 | v_14079;
assign v_14082 = v_14077 | v_14081;
assign v_14084 = v_13988 | v_14083;
assign v_14086 = v_13986 | v_14085;
assign v_14088 = v_14083 | v_14087;
assign v_14090 = v_13985 | v_14089;
assign v_14092 = v_13983 | v_14091;
assign v_14094 = v_14089 | v_14093;
assign v_14096 = v_13982 | v_14095;
assign v_14098 = v_13980 | v_14097;
assign v_14100 = v_14095 | v_14099;
assign v_14102 = v_13979 | v_14101;
assign v_14104 = v_13977 | v_14103;
assign v_14106 = v_14101 | v_14105;
assign v_14108 = v_13976 | v_14107;
assign v_14110 = v_13974 | v_14109;
assign v_14112 = v_14107 | v_14111;
assign v_14114 = v_13973 | v_14113;
assign v_14116 = v_13971 | v_14115;
assign v_14118 = v_14113 | v_14117;
assign v_14121 = ~v_13970 | v_14120;
assign v_14128 = v_14018 | v_14127;
assign v_14131 = v_14129 | v_14130;
assign v_14133 = v_14015 | v_14132;
assign v_14136 = v_14134 | v_14135;
assign v_14138 = v_14012 | v_14137;
assign v_14141 = v_14139 | v_14140;
assign v_14143 = v_14009 | v_14142;
assign v_14146 = v_14144 | v_14145;
assign v_14148 = v_14006 | v_14147;
assign v_14151 = v_14149 | v_14150;
assign v_14153 = v_14003 | v_14152;
assign v_14156 = v_14154 | v_14155;
assign v_14158 = v_14000 | v_14157;
assign v_14161 = v_14159 | v_14160;
assign v_14163 = v_13997 | v_14162;
assign v_14166 = v_14164 | v_14165;
assign v_14168 = v_13994 | v_14167;
assign v_14171 = v_14169 | v_14170;
assign v_14173 = v_13991 | v_14172;
assign v_14176 = v_14174 | v_14175;
assign v_14178 = v_13988 | v_14177;
assign v_14181 = v_14179 | v_14180;
assign v_14183 = v_13985 | v_14182;
assign v_14186 = v_14184 | v_14185;
assign v_14188 = v_13982 | v_14187;
assign v_14191 = v_14189 | v_14190;
assign v_14193 = v_13979 | v_14192;
assign v_14196 = v_14194 | v_14195;
assign v_14198 = v_13976 | v_14197;
assign v_14201 = v_14199 | v_14200;
assign v_14203 = v_13973 | v_14202;
assign v_14206 = v_14204 | v_14205;
assign v_14208 = v_13970 | v_14207;
assign v_14211 = v_13969 | v_14210;
assign v_14265 = v_14262 | v_14264;
assign v_14267 = v_14261 | v_14266;
assign v_14269 = v_14259 | v_14268;
assign v_14271 = v_14266 | v_14270;
assign v_14273 = v_14258 | v_14272;
assign v_14275 = v_14256 | v_14274;
assign v_14277 = v_14272 | v_14276;
assign v_14279 = v_14255 | v_14278;
assign v_14281 = v_14253 | v_14280;
assign v_14283 = v_14278 | v_14282;
assign v_14285 = v_14252 | v_14284;
assign v_14287 = v_14250 | v_14286;
assign v_14289 = v_14284 | v_14288;
assign v_14291 = v_14249 | v_14290;
assign v_14293 = v_14247 | v_14292;
assign v_14295 = v_14290 | v_14294;
assign v_14297 = v_14246 | v_14296;
assign v_14299 = v_14244 | v_14298;
assign v_14301 = v_14296 | v_14300;
assign v_14303 = v_14243 | v_14302;
assign v_14305 = v_14241 | v_14304;
assign v_14307 = v_14302 | v_14306;
assign v_14309 = v_14240 | v_14308;
assign v_14311 = v_14238 | v_14310;
assign v_14313 = v_14308 | v_14312;
assign v_14315 = v_14237 | v_14314;
assign v_14317 = v_14235 | v_14316;
assign v_14319 = v_14314 | v_14318;
assign v_14321 = v_14234 | v_14320;
assign v_14323 = v_14232 | v_14322;
assign v_14325 = v_14320 | v_14324;
assign v_14327 = v_14231 | v_14326;
assign v_14329 = v_14229 | v_14328;
assign v_14331 = v_14326 | v_14330;
assign v_14333 = v_14228 | v_14332;
assign v_14335 = v_14226 | v_14334;
assign v_14337 = v_14332 | v_14336;
assign v_14339 = v_14225 | v_14338;
assign v_14341 = v_14223 | v_14340;
assign v_14343 = v_14338 | v_14342;
assign v_14345 = v_14222 | v_14344;
assign v_14347 = v_14220 | v_14346;
assign v_14349 = v_14344 | v_14348;
assign v_14351 = v_14219 | v_14350;
assign v_14353 = v_14217 | v_14352;
assign v_14355 = v_14350 | v_14354;
assign v_14357 = v_14216 | v_14356;
assign v_14359 = v_14214 | v_14358;
assign v_14361 = v_14356 | v_14360;
assign v_14364 = ~v_14213 | v_14363;
assign v_14371 = v_14261 | v_14370;
assign v_14374 = v_14372 | v_14373;
assign v_14376 = v_14258 | v_14375;
assign v_14379 = v_14377 | v_14378;
assign v_14381 = v_14255 | v_14380;
assign v_14384 = v_14382 | v_14383;
assign v_14386 = v_14252 | v_14385;
assign v_14389 = v_14387 | v_14388;
assign v_14391 = v_14249 | v_14390;
assign v_14394 = v_14392 | v_14393;
assign v_14396 = v_14246 | v_14395;
assign v_14399 = v_14397 | v_14398;
assign v_14401 = v_14243 | v_14400;
assign v_14404 = v_14402 | v_14403;
assign v_14406 = v_14240 | v_14405;
assign v_14409 = v_14407 | v_14408;
assign v_14411 = v_14237 | v_14410;
assign v_14414 = v_14412 | v_14413;
assign v_14416 = v_14234 | v_14415;
assign v_14419 = v_14417 | v_14418;
assign v_14421 = v_14231 | v_14420;
assign v_14424 = v_14422 | v_14423;
assign v_14426 = v_14228 | v_14425;
assign v_14429 = v_14427 | v_14428;
assign v_14431 = v_14225 | v_14430;
assign v_14434 = v_14432 | v_14433;
assign v_14436 = v_14222 | v_14435;
assign v_14439 = v_14437 | v_14438;
assign v_14441 = v_14219 | v_14440;
assign v_14444 = v_14442 | v_14443;
assign v_14446 = v_14216 | v_14445;
assign v_14449 = v_14447 | v_14448;
assign v_14451 = v_14213 | v_14450;
assign v_14454 = v_14212 | v_14453;
assign v_14508 = v_14505 | v_14507;
assign v_14510 = v_14504 | v_14509;
assign v_14512 = v_14502 | v_14511;
assign v_14514 = v_14509 | v_14513;
assign v_14516 = v_14501 | v_14515;
assign v_14518 = v_14499 | v_14517;
assign v_14520 = v_14515 | v_14519;
assign v_14522 = v_14498 | v_14521;
assign v_14524 = v_14496 | v_14523;
assign v_14526 = v_14521 | v_14525;
assign v_14528 = v_14495 | v_14527;
assign v_14530 = v_14493 | v_14529;
assign v_14532 = v_14527 | v_14531;
assign v_14534 = v_14492 | v_14533;
assign v_14536 = v_14490 | v_14535;
assign v_14538 = v_14533 | v_14537;
assign v_14540 = v_14489 | v_14539;
assign v_14542 = v_14487 | v_14541;
assign v_14544 = v_14539 | v_14543;
assign v_14546 = v_14486 | v_14545;
assign v_14548 = v_14484 | v_14547;
assign v_14550 = v_14545 | v_14549;
assign v_14552 = v_14483 | v_14551;
assign v_14554 = v_14481 | v_14553;
assign v_14556 = v_14551 | v_14555;
assign v_14558 = v_14480 | v_14557;
assign v_14560 = v_14478 | v_14559;
assign v_14562 = v_14557 | v_14561;
assign v_14564 = v_14477 | v_14563;
assign v_14566 = v_14475 | v_14565;
assign v_14568 = v_14563 | v_14567;
assign v_14570 = v_14474 | v_14569;
assign v_14572 = v_14472 | v_14571;
assign v_14574 = v_14569 | v_14573;
assign v_14576 = v_14471 | v_14575;
assign v_14578 = v_14469 | v_14577;
assign v_14580 = v_14575 | v_14579;
assign v_14582 = v_14468 | v_14581;
assign v_14584 = v_14466 | v_14583;
assign v_14586 = v_14581 | v_14585;
assign v_14588 = v_14465 | v_14587;
assign v_14590 = v_14463 | v_14589;
assign v_14592 = v_14587 | v_14591;
assign v_14594 = v_14462 | v_14593;
assign v_14596 = v_14460 | v_14595;
assign v_14598 = v_14593 | v_14597;
assign v_14600 = v_14459 | v_14599;
assign v_14602 = v_14457 | v_14601;
assign v_14604 = v_14599 | v_14603;
assign v_14607 = ~v_14456 | v_14606;
assign v_14614 = v_14504 | v_14613;
assign v_14617 = v_14615 | v_14616;
assign v_14619 = v_14501 | v_14618;
assign v_14622 = v_14620 | v_14621;
assign v_14624 = v_14498 | v_14623;
assign v_14627 = v_14625 | v_14626;
assign v_14629 = v_14495 | v_14628;
assign v_14632 = v_14630 | v_14631;
assign v_14634 = v_14492 | v_14633;
assign v_14637 = v_14635 | v_14636;
assign v_14639 = v_14489 | v_14638;
assign v_14642 = v_14640 | v_14641;
assign v_14644 = v_14486 | v_14643;
assign v_14647 = v_14645 | v_14646;
assign v_14649 = v_14483 | v_14648;
assign v_14652 = v_14650 | v_14651;
assign v_14654 = v_14480 | v_14653;
assign v_14657 = v_14655 | v_14656;
assign v_14659 = v_14477 | v_14658;
assign v_14662 = v_14660 | v_14661;
assign v_14664 = v_14474 | v_14663;
assign v_14667 = v_14665 | v_14666;
assign v_14669 = v_14471 | v_14668;
assign v_14672 = v_14670 | v_14671;
assign v_14674 = v_14468 | v_14673;
assign v_14677 = v_14675 | v_14676;
assign v_14679 = v_14465 | v_14678;
assign v_14682 = v_14680 | v_14681;
assign v_14684 = v_14462 | v_14683;
assign v_14687 = v_14685 | v_14686;
assign v_14689 = v_14459 | v_14688;
assign v_14692 = v_14690 | v_14691;
assign v_14694 = v_14456 | v_14693;
assign v_14697 = v_14455 | v_14696;
assign v_14751 = v_14748 | v_14750;
assign v_14753 = v_14747 | v_14752;
assign v_14755 = v_14745 | v_14754;
assign v_14757 = v_14752 | v_14756;
assign v_14759 = v_14744 | v_14758;
assign v_14761 = v_14742 | v_14760;
assign v_14763 = v_14758 | v_14762;
assign v_14765 = v_14741 | v_14764;
assign v_14767 = v_14739 | v_14766;
assign v_14769 = v_14764 | v_14768;
assign v_14771 = v_14738 | v_14770;
assign v_14773 = v_14736 | v_14772;
assign v_14775 = v_14770 | v_14774;
assign v_14777 = v_14735 | v_14776;
assign v_14779 = v_14733 | v_14778;
assign v_14781 = v_14776 | v_14780;
assign v_14783 = v_14732 | v_14782;
assign v_14785 = v_14730 | v_14784;
assign v_14787 = v_14782 | v_14786;
assign v_14789 = v_14729 | v_14788;
assign v_14791 = v_14727 | v_14790;
assign v_14793 = v_14788 | v_14792;
assign v_14795 = v_14726 | v_14794;
assign v_14797 = v_14724 | v_14796;
assign v_14799 = v_14794 | v_14798;
assign v_14801 = v_14723 | v_14800;
assign v_14803 = v_14721 | v_14802;
assign v_14805 = v_14800 | v_14804;
assign v_14807 = v_14720 | v_14806;
assign v_14809 = v_14718 | v_14808;
assign v_14811 = v_14806 | v_14810;
assign v_14813 = v_14717 | v_14812;
assign v_14815 = v_14715 | v_14814;
assign v_14817 = v_14812 | v_14816;
assign v_14819 = v_14714 | v_14818;
assign v_14821 = v_14712 | v_14820;
assign v_14823 = v_14818 | v_14822;
assign v_14825 = v_14711 | v_14824;
assign v_14827 = v_14709 | v_14826;
assign v_14829 = v_14824 | v_14828;
assign v_14831 = v_14708 | v_14830;
assign v_14833 = v_14706 | v_14832;
assign v_14835 = v_14830 | v_14834;
assign v_14837 = v_14705 | v_14836;
assign v_14839 = v_14703 | v_14838;
assign v_14841 = v_14836 | v_14840;
assign v_14843 = v_14702 | v_14842;
assign v_14845 = v_14700 | v_14844;
assign v_14847 = v_14842 | v_14846;
assign v_14850 = ~v_14699 | v_14849;
assign v_14857 = v_14747 | v_14856;
assign v_14860 = v_14858 | v_14859;
assign v_14862 = v_14744 | v_14861;
assign v_14865 = v_14863 | v_14864;
assign v_14867 = v_14741 | v_14866;
assign v_14870 = v_14868 | v_14869;
assign v_14872 = v_14738 | v_14871;
assign v_14875 = v_14873 | v_14874;
assign v_14877 = v_14735 | v_14876;
assign v_14880 = v_14878 | v_14879;
assign v_14882 = v_14732 | v_14881;
assign v_14885 = v_14883 | v_14884;
assign v_14887 = v_14729 | v_14886;
assign v_14890 = v_14888 | v_14889;
assign v_14892 = v_14726 | v_14891;
assign v_14895 = v_14893 | v_14894;
assign v_14897 = v_14723 | v_14896;
assign v_14900 = v_14898 | v_14899;
assign v_14902 = v_14720 | v_14901;
assign v_14905 = v_14903 | v_14904;
assign v_14907 = v_14717 | v_14906;
assign v_14910 = v_14908 | v_14909;
assign v_14912 = v_14714 | v_14911;
assign v_14915 = v_14913 | v_14914;
assign v_14917 = v_14711 | v_14916;
assign v_14920 = v_14918 | v_14919;
assign v_14922 = v_14708 | v_14921;
assign v_14925 = v_14923 | v_14924;
assign v_14927 = v_14705 | v_14926;
assign v_14930 = v_14928 | v_14929;
assign v_14932 = v_14702 | v_14931;
assign v_14935 = v_14933 | v_14934;
assign v_14937 = v_14699 | v_14936;
assign v_14940 = v_14698 | v_14939;
assign v_14994 = v_14991 | v_14993;
assign v_14996 = v_14990 | v_14995;
assign v_14998 = v_14988 | v_14997;
assign v_15000 = v_14995 | v_14999;
assign v_15002 = v_14987 | v_15001;
assign v_15004 = v_14985 | v_15003;
assign v_15006 = v_15001 | v_15005;
assign v_15008 = v_14984 | v_15007;
assign v_15010 = v_14982 | v_15009;
assign v_15012 = v_15007 | v_15011;
assign v_15014 = v_14981 | v_15013;
assign v_15016 = v_14979 | v_15015;
assign v_15018 = v_15013 | v_15017;
assign v_15020 = v_14978 | v_15019;
assign v_15022 = v_14976 | v_15021;
assign v_15024 = v_15019 | v_15023;
assign v_15026 = v_14975 | v_15025;
assign v_15028 = v_14973 | v_15027;
assign v_15030 = v_15025 | v_15029;
assign v_15032 = v_14972 | v_15031;
assign v_15034 = v_14970 | v_15033;
assign v_15036 = v_15031 | v_15035;
assign v_15038 = v_14969 | v_15037;
assign v_15040 = v_14967 | v_15039;
assign v_15042 = v_15037 | v_15041;
assign v_15044 = v_14966 | v_15043;
assign v_15046 = v_14964 | v_15045;
assign v_15048 = v_15043 | v_15047;
assign v_15050 = v_14963 | v_15049;
assign v_15052 = v_14961 | v_15051;
assign v_15054 = v_15049 | v_15053;
assign v_15056 = v_14960 | v_15055;
assign v_15058 = v_14958 | v_15057;
assign v_15060 = v_15055 | v_15059;
assign v_15062 = v_14957 | v_15061;
assign v_15064 = v_14955 | v_15063;
assign v_15066 = v_15061 | v_15065;
assign v_15068 = v_14954 | v_15067;
assign v_15070 = v_14952 | v_15069;
assign v_15072 = v_15067 | v_15071;
assign v_15074 = v_14951 | v_15073;
assign v_15076 = v_14949 | v_15075;
assign v_15078 = v_15073 | v_15077;
assign v_15080 = v_14948 | v_15079;
assign v_15082 = v_14946 | v_15081;
assign v_15084 = v_15079 | v_15083;
assign v_15086 = v_14945 | v_15085;
assign v_15088 = v_14943 | v_15087;
assign v_15090 = v_15085 | v_15089;
assign v_15093 = ~v_14942 | v_15092;
assign v_15100 = v_14990 | v_15099;
assign v_15103 = v_15101 | v_15102;
assign v_15105 = v_14987 | v_15104;
assign v_15108 = v_15106 | v_15107;
assign v_15110 = v_14984 | v_15109;
assign v_15113 = v_15111 | v_15112;
assign v_15115 = v_14981 | v_15114;
assign v_15118 = v_15116 | v_15117;
assign v_15120 = v_14978 | v_15119;
assign v_15123 = v_15121 | v_15122;
assign v_15125 = v_14975 | v_15124;
assign v_15128 = v_15126 | v_15127;
assign v_15130 = v_14972 | v_15129;
assign v_15133 = v_15131 | v_15132;
assign v_15135 = v_14969 | v_15134;
assign v_15138 = v_15136 | v_15137;
assign v_15140 = v_14966 | v_15139;
assign v_15143 = v_15141 | v_15142;
assign v_15145 = v_14963 | v_15144;
assign v_15148 = v_15146 | v_15147;
assign v_15150 = v_14960 | v_15149;
assign v_15153 = v_15151 | v_15152;
assign v_15155 = v_14957 | v_15154;
assign v_15158 = v_15156 | v_15157;
assign v_15160 = v_14954 | v_15159;
assign v_15163 = v_15161 | v_15162;
assign v_15165 = v_14951 | v_15164;
assign v_15168 = v_15166 | v_15167;
assign v_15170 = v_14948 | v_15169;
assign v_15173 = v_15171 | v_15172;
assign v_15175 = v_14945 | v_15174;
assign v_15178 = v_15176 | v_15177;
assign v_15180 = v_14942 | v_15179;
assign v_15183 = v_14941 | v_15182;
assign v_15237 = v_15234 | v_15236;
assign v_15239 = v_15233 | v_15238;
assign v_15241 = v_15231 | v_15240;
assign v_15243 = v_15238 | v_15242;
assign v_15245 = v_15230 | v_15244;
assign v_15247 = v_15228 | v_15246;
assign v_15249 = v_15244 | v_15248;
assign v_15251 = v_15227 | v_15250;
assign v_15253 = v_15225 | v_15252;
assign v_15255 = v_15250 | v_15254;
assign v_15257 = v_15224 | v_15256;
assign v_15259 = v_15222 | v_15258;
assign v_15261 = v_15256 | v_15260;
assign v_15263 = v_15221 | v_15262;
assign v_15265 = v_15219 | v_15264;
assign v_15267 = v_15262 | v_15266;
assign v_15269 = v_15218 | v_15268;
assign v_15271 = v_15216 | v_15270;
assign v_15273 = v_15268 | v_15272;
assign v_15275 = v_15215 | v_15274;
assign v_15277 = v_15213 | v_15276;
assign v_15279 = v_15274 | v_15278;
assign v_15281 = v_15212 | v_15280;
assign v_15283 = v_15210 | v_15282;
assign v_15285 = v_15280 | v_15284;
assign v_15287 = v_15209 | v_15286;
assign v_15289 = v_15207 | v_15288;
assign v_15291 = v_15286 | v_15290;
assign v_15293 = v_15206 | v_15292;
assign v_15295 = v_15204 | v_15294;
assign v_15297 = v_15292 | v_15296;
assign v_15299 = v_15203 | v_15298;
assign v_15301 = v_15201 | v_15300;
assign v_15303 = v_15298 | v_15302;
assign v_15305 = v_15200 | v_15304;
assign v_15307 = v_15198 | v_15306;
assign v_15309 = v_15304 | v_15308;
assign v_15311 = v_15197 | v_15310;
assign v_15313 = v_15195 | v_15312;
assign v_15315 = v_15310 | v_15314;
assign v_15317 = v_15194 | v_15316;
assign v_15319 = v_15192 | v_15318;
assign v_15321 = v_15316 | v_15320;
assign v_15323 = v_15191 | v_15322;
assign v_15325 = v_15189 | v_15324;
assign v_15327 = v_15322 | v_15326;
assign v_15329 = v_15188 | v_15328;
assign v_15331 = v_15186 | v_15330;
assign v_15333 = v_15328 | v_15332;
assign v_15336 = ~v_15185 | v_15335;
assign v_15343 = v_15233 | v_15342;
assign v_15346 = v_15344 | v_15345;
assign v_15348 = v_15230 | v_15347;
assign v_15351 = v_15349 | v_15350;
assign v_15353 = v_15227 | v_15352;
assign v_15356 = v_15354 | v_15355;
assign v_15358 = v_15224 | v_15357;
assign v_15361 = v_15359 | v_15360;
assign v_15363 = v_15221 | v_15362;
assign v_15366 = v_15364 | v_15365;
assign v_15368 = v_15218 | v_15367;
assign v_15371 = v_15369 | v_15370;
assign v_15373 = v_15215 | v_15372;
assign v_15376 = v_15374 | v_15375;
assign v_15378 = v_15212 | v_15377;
assign v_15381 = v_15379 | v_15380;
assign v_15383 = v_15209 | v_15382;
assign v_15386 = v_15384 | v_15385;
assign v_15388 = v_15206 | v_15387;
assign v_15391 = v_15389 | v_15390;
assign v_15393 = v_15203 | v_15392;
assign v_15396 = v_15394 | v_15395;
assign v_15398 = v_15200 | v_15397;
assign v_15401 = v_15399 | v_15400;
assign v_15403 = v_15197 | v_15402;
assign v_15406 = v_15404 | v_15405;
assign v_15408 = v_15194 | v_15407;
assign v_15411 = v_15409 | v_15410;
assign v_15413 = v_15191 | v_15412;
assign v_15416 = v_15414 | v_15415;
assign v_15418 = v_15188 | v_15417;
assign v_15421 = v_15419 | v_15420;
assign v_15423 = v_15185 | v_15422;
assign v_15426 = v_15184 | v_15425;
assign v_15480 = v_15477 | v_15479;
assign v_15482 = v_15476 | v_15481;
assign v_15484 = v_15474 | v_15483;
assign v_15486 = v_15481 | v_15485;
assign v_15488 = v_15473 | v_15487;
assign v_15490 = v_15471 | v_15489;
assign v_15492 = v_15487 | v_15491;
assign v_15494 = v_15470 | v_15493;
assign v_15496 = v_15468 | v_15495;
assign v_15498 = v_15493 | v_15497;
assign v_15500 = v_15467 | v_15499;
assign v_15502 = v_15465 | v_15501;
assign v_15504 = v_15499 | v_15503;
assign v_15506 = v_15464 | v_15505;
assign v_15508 = v_15462 | v_15507;
assign v_15510 = v_15505 | v_15509;
assign v_15512 = v_15461 | v_15511;
assign v_15514 = v_15459 | v_15513;
assign v_15516 = v_15511 | v_15515;
assign v_15518 = v_15458 | v_15517;
assign v_15520 = v_15456 | v_15519;
assign v_15522 = v_15517 | v_15521;
assign v_15524 = v_15455 | v_15523;
assign v_15526 = v_15453 | v_15525;
assign v_15528 = v_15523 | v_15527;
assign v_15530 = v_15452 | v_15529;
assign v_15532 = v_15450 | v_15531;
assign v_15534 = v_15529 | v_15533;
assign v_15536 = v_15449 | v_15535;
assign v_15538 = v_15447 | v_15537;
assign v_15540 = v_15535 | v_15539;
assign v_15542 = v_15446 | v_15541;
assign v_15544 = v_15444 | v_15543;
assign v_15546 = v_15541 | v_15545;
assign v_15548 = v_15443 | v_15547;
assign v_15550 = v_15441 | v_15549;
assign v_15552 = v_15547 | v_15551;
assign v_15554 = v_15440 | v_15553;
assign v_15556 = v_15438 | v_15555;
assign v_15558 = v_15553 | v_15557;
assign v_15560 = v_15437 | v_15559;
assign v_15562 = v_15435 | v_15561;
assign v_15564 = v_15559 | v_15563;
assign v_15566 = v_15434 | v_15565;
assign v_15568 = v_15432 | v_15567;
assign v_15570 = v_15565 | v_15569;
assign v_15572 = v_15431 | v_15571;
assign v_15574 = v_15429 | v_15573;
assign v_15576 = v_15571 | v_15575;
assign v_15579 = ~v_15428 | v_15578;
assign v_15586 = v_15476 | v_15585;
assign v_15589 = v_15587 | v_15588;
assign v_15591 = v_15473 | v_15590;
assign v_15594 = v_15592 | v_15593;
assign v_15596 = v_15470 | v_15595;
assign v_15599 = v_15597 | v_15598;
assign v_15601 = v_15467 | v_15600;
assign v_15604 = v_15602 | v_15603;
assign v_15606 = v_15464 | v_15605;
assign v_15609 = v_15607 | v_15608;
assign v_15611 = v_15461 | v_15610;
assign v_15614 = v_15612 | v_15613;
assign v_15616 = v_15458 | v_15615;
assign v_15619 = v_15617 | v_15618;
assign v_15621 = v_15455 | v_15620;
assign v_15624 = v_15622 | v_15623;
assign v_15626 = v_15452 | v_15625;
assign v_15629 = v_15627 | v_15628;
assign v_15631 = v_15449 | v_15630;
assign v_15634 = v_15632 | v_15633;
assign v_15636 = v_15446 | v_15635;
assign v_15639 = v_15637 | v_15638;
assign v_15641 = v_15443 | v_15640;
assign v_15644 = v_15642 | v_15643;
assign v_15646 = v_15440 | v_15645;
assign v_15649 = v_15647 | v_15648;
assign v_15651 = v_15437 | v_15650;
assign v_15654 = v_15652 | v_15653;
assign v_15656 = v_15434 | v_15655;
assign v_15659 = v_15657 | v_15658;
assign v_15661 = v_15431 | v_15660;
assign v_15664 = v_15662 | v_15663;
assign v_15666 = v_15428 | v_15665;
assign v_15669 = v_15427 | v_15668;
assign v_15723 = v_15720 | v_15722;
assign v_15725 = v_15719 | v_15724;
assign v_15727 = v_15717 | v_15726;
assign v_15729 = v_15724 | v_15728;
assign v_15731 = v_15716 | v_15730;
assign v_15733 = v_15714 | v_15732;
assign v_15735 = v_15730 | v_15734;
assign v_15737 = v_15713 | v_15736;
assign v_15739 = v_15711 | v_15738;
assign v_15741 = v_15736 | v_15740;
assign v_15743 = v_15710 | v_15742;
assign v_15745 = v_15708 | v_15744;
assign v_15747 = v_15742 | v_15746;
assign v_15749 = v_15707 | v_15748;
assign v_15751 = v_15705 | v_15750;
assign v_15753 = v_15748 | v_15752;
assign v_15755 = v_15704 | v_15754;
assign v_15757 = v_15702 | v_15756;
assign v_15759 = v_15754 | v_15758;
assign v_15761 = v_15701 | v_15760;
assign v_15763 = v_15699 | v_15762;
assign v_15765 = v_15760 | v_15764;
assign v_15767 = v_15698 | v_15766;
assign v_15769 = v_15696 | v_15768;
assign v_15771 = v_15766 | v_15770;
assign v_15773 = v_15695 | v_15772;
assign v_15775 = v_15693 | v_15774;
assign v_15777 = v_15772 | v_15776;
assign v_15779 = v_15692 | v_15778;
assign v_15781 = v_15690 | v_15780;
assign v_15783 = v_15778 | v_15782;
assign v_15785 = v_15689 | v_15784;
assign v_15787 = v_15687 | v_15786;
assign v_15789 = v_15784 | v_15788;
assign v_15791 = v_15686 | v_15790;
assign v_15793 = v_15684 | v_15792;
assign v_15795 = v_15790 | v_15794;
assign v_15797 = v_15683 | v_15796;
assign v_15799 = v_15681 | v_15798;
assign v_15801 = v_15796 | v_15800;
assign v_15803 = v_15680 | v_15802;
assign v_15805 = v_15678 | v_15804;
assign v_15807 = v_15802 | v_15806;
assign v_15809 = v_15677 | v_15808;
assign v_15811 = v_15675 | v_15810;
assign v_15813 = v_15808 | v_15812;
assign v_15815 = v_15674 | v_15814;
assign v_15817 = v_15672 | v_15816;
assign v_15819 = v_15814 | v_15818;
assign v_15822 = ~v_15671 | v_15821;
assign v_15829 = v_15719 | v_15828;
assign v_15832 = v_15830 | v_15831;
assign v_15834 = v_15716 | v_15833;
assign v_15837 = v_15835 | v_15836;
assign v_15839 = v_15713 | v_15838;
assign v_15842 = v_15840 | v_15841;
assign v_15844 = v_15710 | v_15843;
assign v_15847 = v_15845 | v_15846;
assign v_15849 = v_15707 | v_15848;
assign v_15852 = v_15850 | v_15851;
assign v_15854 = v_15704 | v_15853;
assign v_15857 = v_15855 | v_15856;
assign v_15859 = v_15701 | v_15858;
assign v_15862 = v_15860 | v_15861;
assign v_15864 = v_15698 | v_15863;
assign v_15867 = v_15865 | v_15866;
assign v_15869 = v_15695 | v_15868;
assign v_15872 = v_15870 | v_15871;
assign v_15874 = v_15692 | v_15873;
assign v_15877 = v_15875 | v_15876;
assign v_15879 = v_15689 | v_15878;
assign v_15882 = v_15880 | v_15881;
assign v_15884 = v_15686 | v_15883;
assign v_15887 = v_15885 | v_15886;
assign v_15889 = v_15683 | v_15888;
assign v_15892 = v_15890 | v_15891;
assign v_15894 = v_15680 | v_15893;
assign v_15897 = v_15895 | v_15896;
assign v_15899 = v_15677 | v_15898;
assign v_15902 = v_15900 | v_15901;
assign v_15904 = v_15674 | v_15903;
assign v_15907 = v_15905 | v_15906;
assign v_15909 = v_15671 | v_15908;
assign v_15912 = v_15670 | v_15911;
assign v_15966 = v_15963 | v_15965;
assign v_15968 = v_15962 | v_15967;
assign v_15970 = v_15960 | v_15969;
assign v_15972 = v_15967 | v_15971;
assign v_15974 = v_15959 | v_15973;
assign v_15976 = v_15957 | v_15975;
assign v_15978 = v_15973 | v_15977;
assign v_15980 = v_15956 | v_15979;
assign v_15982 = v_15954 | v_15981;
assign v_15984 = v_15979 | v_15983;
assign v_15986 = v_15953 | v_15985;
assign v_15988 = v_15951 | v_15987;
assign v_15990 = v_15985 | v_15989;
assign v_15992 = v_15950 | v_15991;
assign v_15994 = v_15948 | v_15993;
assign v_15996 = v_15991 | v_15995;
assign v_15998 = v_15947 | v_15997;
assign v_16000 = v_15945 | v_15999;
assign v_16002 = v_15997 | v_16001;
assign v_16004 = v_15944 | v_16003;
assign v_16006 = v_15942 | v_16005;
assign v_16008 = v_16003 | v_16007;
assign v_16010 = v_15941 | v_16009;
assign v_16012 = v_15939 | v_16011;
assign v_16014 = v_16009 | v_16013;
assign v_16016 = v_15938 | v_16015;
assign v_16018 = v_15936 | v_16017;
assign v_16020 = v_16015 | v_16019;
assign v_16022 = v_15935 | v_16021;
assign v_16024 = v_15933 | v_16023;
assign v_16026 = v_16021 | v_16025;
assign v_16028 = v_15932 | v_16027;
assign v_16030 = v_15930 | v_16029;
assign v_16032 = v_16027 | v_16031;
assign v_16034 = v_15929 | v_16033;
assign v_16036 = v_15927 | v_16035;
assign v_16038 = v_16033 | v_16037;
assign v_16040 = v_15926 | v_16039;
assign v_16042 = v_15924 | v_16041;
assign v_16044 = v_16039 | v_16043;
assign v_16046 = v_15923 | v_16045;
assign v_16048 = v_15921 | v_16047;
assign v_16050 = v_16045 | v_16049;
assign v_16052 = v_15920 | v_16051;
assign v_16054 = v_15918 | v_16053;
assign v_16056 = v_16051 | v_16055;
assign v_16058 = v_15917 | v_16057;
assign v_16060 = v_15915 | v_16059;
assign v_16062 = v_16057 | v_16061;
assign v_16065 = ~v_15914 | v_16064;
assign v_16072 = v_15962 | v_16071;
assign v_16075 = v_16073 | v_16074;
assign v_16077 = v_15959 | v_16076;
assign v_16080 = v_16078 | v_16079;
assign v_16082 = v_15956 | v_16081;
assign v_16085 = v_16083 | v_16084;
assign v_16087 = v_15953 | v_16086;
assign v_16090 = v_16088 | v_16089;
assign v_16092 = v_15950 | v_16091;
assign v_16095 = v_16093 | v_16094;
assign v_16097 = v_15947 | v_16096;
assign v_16100 = v_16098 | v_16099;
assign v_16102 = v_15944 | v_16101;
assign v_16105 = v_16103 | v_16104;
assign v_16107 = v_15941 | v_16106;
assign v_16110 = v_16108 | v_16109;
assign v_16112 = v_15938 | v_16111;
assign v_16115 = v_16113 | v_16114;
assign v_16117 = v_15935 | v_16116;
assign v_16120 = v_16118 | v_16119;
assign v_16122 = v_15932 | v_16121;
assign v_16125 = v_16123 | v_16124;
assign v_16127 = v_15929 | v_16126;
assign v_16130 = v_16128 | v_16129;
assign v_16132 = v_15926 | v_16131;
assign v_16135 = v_16133 | v_16134;
assign v_16137 = v_15923 | v_16136;
assign v_16140 = v_16138 | v_16139;
assign v_16142 = v_15920 | v_16141;
assign v_16145 = v_16143 | v_16144;
assign v_16147 = v_15917 | v_16146;
assign v_16150 = v_16148 | v_16149;
assign v_16152 = v_15914 | v_16151;
assign v_16155 = v_15913 | v_16154;
assign v_16209 = v_16206 | v_16208;
assign v_16211 = v_16205 | v_16210;
assign v_16213 = v_16203 | v_16212;
assign v_16215 = v_16210 | v_16214;
assign v_16217 = v_16202 | v_16216;
assign v_16219 = v_16200 | v_16218;
assign v_16221 = v_16216 | v_16220;
assign v_16223 = v_16199 | v_16222;
assign v_16225 = v_16197 | v_16224;
assign v_16227 = v_16222 | v_16226;
assign v_16229 = v_16196 | v_16228;
assign v_16231 = v_16194 | v_16230;
assign v_16233 = v_16228 | v_16232;
assign v_16235 = v_16193 | v_16234;
assign v_16237 = v_16191 | v_16236;
assign v_16239 = v_16234 | v_16238;
assign v_16241 = v_16190 | v_16240;
assign v_16243 = v_16188 | v_16242;
assign v_16245 = v_16240 | v_16244;
assign v_16247 = v_16187 | v_16246;
assign v_16249 = v_16185 | v_16248;
assign v_16251 = v_16246 | v_16250;
assign v_16253 = v_16184 | v_16252;
assign v_16255 = v_16182 | v_16254;
assign v_16257 = v_16252 | v_16256;
assign v_16259 = v_16181 | v_16258;
assign v_16261 = v_16179 | v_16260;
assign v_16263 = v_16258 | v_16262;
assign v_16265 = v_16178 | v_16264;
assign v_16267 = v_16176 | v_16266;
assign v_16269 = v_16264 | v_16268;
assign v_16271 = v_16175 | v_16270;
assign v_16273 = v_16173 | v_16272;
assign v_16275 = v_16270 | v_16274;
assign v_16277 = v_16172 | v_16276;
assign v_16279 = v_16170 | v_16278;
assign v_16281 = v_16276 | v_16280;
assign v_16283 = v_16169 | v_16282;
assign v_16285 = v_16167 | v_16284;
assign v_16287 = v_16282 | v_16286;
assign v_16289 = v_16166 | v_16288;
assign v_16291 = v_16164 | v_16290;
assign v_16293 = v_16288 | v_16292;
assign v_16295 = v_16163 | v_16294;
assign v_16297 = v_16161 | v_16296;
assign v_16299 = v_16294 | v_16298;
assign v_16301 = v_16160 | v_16300;
assign v_16303 = v_16158 | v_16302;
assign v_16305 = v_16300 | v_16304;
assign v_16308 = ~v_16157 | v_16307;
assign v_16315 = v_16205 | v_16314;
assign v_16318 = v_16316 | v_16317;
assign v_16320 = v_16202 | v_16319;
assign v_16323 = v_16321 | v_16322;
assign v_16325 = v_16199 | v_16324;
assign v_16328 = v_16326 | v_16327;
assign v_16330 = v_16196 | v_16329;
assign v_16333 = v_16331 | v_16332;
assign v_16335 = v_16193 | v_16334;
assign v_16338 = v_16336 | v_16337;
assign v_16340 = v_16190 | v_16339;
assign v_16343 = v_16341 | v_16342;
assign v_16345 = v_16187 | v_16344;
assign v_16348 = v_16346 | v_16347;
assign v_16350 = v_16184 | v_16349;
assign v_16353 = v_16351 | v_16352;
assign v_16355 = v_16181 | v_16354;
assign v_16358 = v_16356 | v_16357;
assign v_16360 = v_16178 | v_16359;
assign v_16363 = v_16361 | v_16362;
assign v_16365 = v_16175 | v_16364;
assign v_16368 = v_16366 | v_16367;
assign v_16370 = v_16172 | v_16369;
assign v_16373 = v_16371 | v_16372;
assign v_16375 = v_16169 | v_16374;
assign v_16378 = v_16376 | v_16377;
assign v_16380 = v_16166 | v_16379;
assign v_16383 = v_16381 | v_16382;
assign v_16385 = v_16163 | v_16384;
assign v_16388 = v_16386 | v_16387;
assign v_16390 = v_16160 | v_16389;
assign v_16393 = v_16391 | v_16392;
assign v_16395 = v_16157 | v_16394;
assign v_16398 = v_16156 | v_16397;
assign v_16452 = v_16449 | v_16451;
assign v_16454 = v_16448 | v_16453;
assign v_16456 = v_16446 | v_16455;
assign v_16458 = v_16453 | v_16457;
assign v_16460 = v_16445 | v_16459;
assign v_16462 = v_16443 | v_16461;
assign v_16464 = v_16459 | v_16463;
assign v_16466 = v_16442 | v_16465;
assign v_16468 = v_16440 | v_16467;
assign v_16470 = v_16465 | v_16469;
assign v_16472 = v_16439 | v_16471;
assign v_16474 = v_16437 | v_16473;
assign v_16476 = v_16471 | v_16475;
assign v_16478 = v_16436 | v_16477;
assign v_16480 = v_16434 | v_16479;
assign v_16482 = v_16477 | v_16481;
assign v_16484 = v_16433 | v_16483;
assign v_16486 = v_16431 | v_16485;
assign v_16488 = v_16483 | v_16487;
assign v_16490 = v_16430 | v_16489;
assign v_16492 = v_16428 | v_16491;
assign v_16494 = v_16489 | v_16493;
assign v_16496 = v_16427 | v_16495;
assign v_16498 = v_16425 | v_16497;
assign v_16500 = v_16495 | v_16499;
assign v_16502 = v_16424 | v_16501;
assign v_16504 = v_16422 | v_16503;
assign v_16506 = v_16501 | v_16505;
assign v_16508 = v_16421 | v_16507;
assign v_16510 = v_16419 | v_16509;
assign v_16512 = v_16507 | v_16511;
assign v_16514 = v_16418 | v_16513;
assign v_16516 = v_16416 | v_16515;
assign v_16518 = v_16513 | v_16517;
assign v_16520 = v_16415 | v_16519;
assign v_16522 = v_16413 | v_16521;
assign v_16524 = v_16519 | v_16523;
assign v_16526 = v_16412 | v_16525;
assign v_16528 = v_16410 | v_16527;
assign v_16530 = v_16525 | v_16529;
assign v_16532 = v_16409 | v_16531;
assign v_16534 = v_16407 | v_16533;
assign v_16536 = v_16531 | v_16535;
assign v_16538 = v_16406 | v_16537;
assign v_16540 = v_16404 | v_16539;
assign v_16542 = v_16537 | v_16541;
assign v_16544 = v_16403 | v_16543;
assign v_16546 = v_16401 | v_16545;
assign v_16548 = v_16543 | v_16547;
assign v_16551 = ~v_16400 | v_16550;
assign v_16558 = v_16448 | v_16557;
assign v_16561 = v_16559 | v_16560;
assign v_16563 = v_16445 | v_16562;
assign v_16566 = v_16564 | v_16565;
assign v_16568 = v_16442 | v_16567;
assign v_16571 = v_16569 | v_16570;
assign v_16573 = v_16439 | v_16572;
assign v_16576 = v_16574 | v_16575;
assign v_16578 = v_16436 | v_16577;
assign v_16581 = v_16579 | v_16580;
assign v_16583 = v_16433 | v_16582;
assign v_16586 = v_16584 | v_16585;
assign v_16588 = v_16430 | v_16587;
assign v_16591 = v_16589 | v_16590;
assign v_16593 = v_16427 | v_16592;
assign v_16596 = v_16594 | v_16595;
assign v_16598 = v_16424 | v_16597;
assign v_16601 = v_16599 | v_16600;
assign v_16603 = v_16421 | v_16602;
assign v_16606 = v_16604 | v_16605;
assign v_16608 = v_16418 | v_16607;
assign v_16611 = v_16609 | v_16610;
assign v_16613 = v_16415 | v_16612;
assign v_16616 = v_16614 | v_16615;
assign v_16618 = v_16412 | v_16617;
assign v_16621 = v_16619 | v_16620;
assign v_16623 = v_16409 | v_16622;
assign v_16626 = v_16624 | v_16625;
assign v_16628 = v_16406 | v_16627;
assign v_16631 = v_16629 | v_16630;
assign v_16633 = v_16403 | v_16632;
assign v_16636 = v_16634 | v_16635;
assign v_16638 = v_16400 | v_16637;
assign v_16641 = v_16399 | v_16640;
assign v_16694 = v_16691 | v_16693;
assign v_16696 = v_16690 | v_16695;
assign v_16698 = v_16688 | v_16697;
assign v_16700 = v_16695 | v_16699;
assign v_16702 = v_16687 | v_16701;
assign v_16704 = v_16685 | v_16703;
assign v_16706 = v_16701 | v_16705;
assign v_16708 = v_16684 | v_16707;
assign v_16710 = v_16682 | v_16709;
assign v_16712 = v_16707 | v_16711;
assign v_16714 = v_16681 | v_16713;
assign v_16716 = v_16679 | v_16715;
assign v_16718 = v_16713 | v_16717;
assign v_16720 = v_16678 | v_16719;
assign v_16722 = v_16676 | v_16721;
assign v_16724 = v_16719 | v_16723;
assign v_16726 = v_16675 | v_16725;
assign v_16728 = v_16673 | v_16727;
assign v_16730 = v_16725 | v_16729;
assign v_16732 = v_16672 | v_16731;
assign v_16734 = v_16670 | v_16733;
assign v_16736 = v_16731 | v_16735;
assign v_16738 = v_16669 | v_16737;
assign v_16740 = v_16667 | v_16739;
assign v_16742 = v_16737 | v_16741;
assign v_16744 = v_16666 | v_16743;
assign v_16746 = v_16664 | v_16745;
assign v_16748 = v_16743 | v_16747;
assign v_16750 = v_16663 | v_16749;
assign v_16752 = v_16661 | v_16751;
assign v_16754 = v_16749 | v_16753;
assign v_16756 = v_16660 | v_16755;
assign v_16758 = v_16658 | v_16757;
assign v_16760 = v_16755 | v_16759;
assign v_16762 = v_16657 | v_16761;
assign v_16764 = v_16655 | v_16763;
assign v_16766 = v_16761 | v_16765;
assign v_16768 = v_16654 | v_16767;
assign v_16770 = v_16652 | v_16769;
assign v_16772 = v_16767 | v_16771;
assign v_16774 = v_16651 | v_16773;
assign v_16776 = v_16649 | v_16775;
assign v_16778 = v_16773 | v_16777;
assign v_16780 = v_16648 | v_16779;
assign v_16782 = v_16646 | v_16781;
assign v_16784 = v_16779 | v_16783;
assign v_16786 = v_16645 | v_16785;
assign v_16788 = v_16643 | v_16787;
assign v_16790 = v_16785 | v_16789;
assign v_16794 = v_16791 | v_16793;
assign v_16801 = v_16690 | v_16800;
assign v_16804 = v_16802 | v_16803;
assign v_16806 = v_16687 | v_16805;
assign v_16809 = v_16807 | v_16808;
assign v_16811 = v_16684 | v_16810;
assign v_16814 = v_16812 | v_16813;
assign v_16816 = v_16681 | v_16815;
assign v_16819 = v_16817 | v_16818;
assign v_16821 = v_16678 | v_16820;
assign v_16824 = v_16822 | v_16823;
assign v_16826 = v_16675 | v_16825;
assign v_16829 = v_16827 | v_16828;
assign v_16831 = v_16672 | v_16830;
assign v_16834 = v_16832 | v_16833;
assign v_16836 = v_16669 | v_16835;
assign v_16839 = v_16837 | v_16838;
assign v_16841 = v_16666 | v_16840;
assign v_16844 = v_16842 | v_16843;
assign v_16846 = v_16663 | v_16845;
assign v_16849 = v_16847 | v_16848;
assign v_16851 = v_16660 | v_16850;
assign v_16854 = v_16852 | v_16853;
assign v_16856 = v_16657 | v_16855;
assign v_16859 = v_16857 | v_16858;
assign v_16861 = v_16654 | v_16860;
assign v_16864 = v_16862 | v_16863;
assign v_16866 = v_16651 | v_16865;
assign v_16869 = v_16867 | v_16868;
assign v_16871 = v_16648 | v_16870;
assign v_16874 = v_16872 | v_16873;
assign v_16876 = v_16645 | v_16875;
assign v_16879 = v_16877 | v_16878;
assign v_16881 = v_16879 | v_16880;
assign v_16884 = v_16642 | v_16883;
assign v_16955 = v_16952 | v_16954;
assign v_16957 = v_16950 | v_16956;
assign v_16959 = v_16948 | v_16958;
assign v_16961 = v_16956 | v_16960;
assign v_16963 = v_16946 | v_16962;
assign v_16965 = v_16944 | v_16964;
assign v_16967 = v_16962 | v_16966;
assign v_16969 = v_16942 | v_16968;
assign v_16971 = v_16940 | v_16970;
assign v_16973 = v_16968 | v_16972;
assign v_16975 = v_16938 | v_16974;
assign v_16977 = v_16936 | v_16976;
assign v_16979 = v_16974 | v_16978;
assign v_16981 = v_16934 | v_16980;
assign v_16983 = v_16932 | v_16982;
assign v_16985 = v_16980 | v_16984;
assign v_16987 = v_16930 | v_16986;
assign v_16989 = v_16928 | v_16988;
assign v_16991 = v_16986 | v_16990;
assign v_16993 = v_16926 | v_16992;
assign v_16995 = v_16924 | v_16994;
assign v_16997 = v_16992 | v_16996;
assign v_16999 = v_16922 | v_16998;
assign v_17001 = v_16920 | v_17000;
assign v_17003 = v_16998 | v_17002;
assign v_17005 = v_16918 | v_17004;
assign v_17007 = v_16916 | v_17006;
assign v_17009 = v_17004 | v_17008;
assign v_17011 = v_16914 | v_17010;
assign v_17013 = v_16912 | v_17012;
assign v_17015 = v_17010 | v_17014;
assign v_17017 = v_16910 | v_17016;
assign v_17019 = v_16908 | v_17018;
assign v_17021 = v_17016 | v_17020;
assign v_17023 = v_16906 | v_17022;
assign v_17025 = v_16904 | v_17024;
assign v_17027 = v_17022 | v_17026;
assign v_17029 = v_16902 | v_17028;
assign v_17031 = v_16899 | v_17030;
assign v_17033 = v_17028 | v_17032;
assign v_17035 = v_16898 | v_17034;
assign v_17037 = v_16895 | v_17036;
assign v_17039 = v_17034 | v_17038;
assign v_17041 = v_16894 | v_17040;
assign v_17043 = v_16891 | v_17042;
assign v_17045 = v_17040 | v_17044;
assign v_17047 = v_16890 | v_17046;
assign v_17049 = v_16887 | v_17048;
assign v_17051 = v_17046 | v_17050;
assign v_17054 = ~v_16886 | v_17053;
assign v_17061 = v_16950 | v_17060;
assign v_17064 = v_17062 | v_17063;
assign v_17066 = v_16946 | v_17065;
assign v_17069 = v_17067 | v_17068;
assign v_17071 = v_16942 | v_17070;
assign v_17074 = v_17072 | v_17073;
assign v_17076 = v_16938 | v_17075;
assign v_17079 = v_17077 | v_17078;
assign v_17081 = v_16934 | v_17080;
assign v_17084 = v_17082 | v_17083;
assign v_17086 = v_16930 | v_17085;
assign v_17089 = v_17087 | v_17088;
assign v_17091 = v_16926 | v_17090;
assign v_17094 = v_17092 | v_17093;
assign v_17096 = v_16922 | v_17095;
assign v_17099 = v_17097 | v_17098;
assign v_17101 = v_16918 | v_17100;
assign v_17104 = v_17102 | v_17103;
assign v_17106 = v_16914 | v_17105;
assign v_17109 = v_17107 | v_17108;
assign v_17111 = v_16910 | v_17110;
assign v_17114 = v_17112 | v_17113;
assign v_17116 = v_16906 | v_17115;
assign v_17119 = v_17117 | v_17118;
assign v_17121 = v_16902 | v_17120;
assign v_17124 = v_17122 | v_17123;
assign v_17126 = v_16898 | v_17125;
assign v_17129 = v_17127 | v_17128;
assign v_17131 = v_16894 | v_17130;
assign v_17134 = v_17132 | v_17133;
assign v_17136 = v_16890 | v_17135;
assign v_17139 = v_17137 | v_17138;
assign v_17141 = v_16886 | v_17140;
assign v_17144 = v_16885 | v_17143;
assign v_17198 = v_17195 | v_17197;
assign v_17200 = v_17194 | v_17199;
assign v_17202 = v_17192 | v_17201;
assign v_17204 = v_17199 | v_17203;
assign v_17206 = v_17191 | v_17205;
assign v_17208 = v_17189 | v_17207;
assign v_17210 = v_17205 | v_17209;
assign v_17212 = v_17188 | v_17211;
assign v_17214 = v_17186 | v_17213;
assign v_17216 = v_17211 | v_17215;
assign v_17218 = v_17185 | v_17217;
assign v_17220 = v_17183 | v_17219;
assign v_17222 = v_17217 | v_17221;
assign v_17224 = v_17182 | v_17223;
assign v_17226 = v_17180 | v_17225;
assign v_17228 = v_17223 | v_17227;
assign v_17230 = v_17179 | v_17229;
assign v_17232 = v_17177 | v_17231;
assign v_17234 = v_17229 | v_17233;
assign v_17236 = v_17176 | v_17235;
assign v_17238 = v_17174 | v_17237;
assign v_17240 = v_17235 | v_17239;
assign v_17242 = v_17173 | v_17241;
assign v_17244 = v_17171 | v_17243;
assign v_17246 = v_17241 | v_17245;
assign v_17248 = v_17170 | v_17247;
assign v_17250 = v_17168 | v_17249;
assign v_17252 = v_17247 | v_17251;
assign v_17254 = v_17167 | v_17253;
assign v_17256 = v_17165 | v_17255;
assign v_17258 = v_17253 | v_17257;
assign v_17260 = v_17164 | v_17259;
assign v_17262 = v_17162 | v_17261;
assign v_17264 = v_17259 | v_17263;
assign v_17266 = v_17161 | v_17265;
assign v_17268 = v_17159 | v_17267;
assign v_17270 = v_17265 | v_17269;
assign v_17272 = v_17158 | v_17271;
assign v_17274 = v_17156 | v_17273;
assign v_17276 = v_17271 | v_17275;
assign v_17278 = v_17155 | v_17277;
assign v_17280 = v_17153 | v_17279;
assign v_17282 = v_17277 | v_17281;
assign v_17284 = v_17152 | v_17283;
assign v_17286 = v_17150 | v_17285;
assign v_17288 = v_17283 | v_17287;
assign v_17290 = v_17149 | v_17289;
assign v_17292 = v_17147 | v_17291;
assign v_17294 = v_17289 | v_17293;
assign v_17297 = ~v_17146 | v_17296;
assign v_17304 = v_17194 | v_17303;
assign v_17307 = v_17305 | v_17306;
assign v_17309 = v_17191 | v_17308;
assign v_17312 = v_17310 | v_17311;
assign v_17314 = v_17188 | v_17313;
assign v_17317 = v_17315 | v_17316;
assign v_17319 = v_17185 | v_17318;
assign v_17322 = v_17320 | v_17321;
assign v_17324 = v_17182 | v_17323;
assign v_17327 = v_17325 | v_17326;
assign v_17329 = v_17179 | v_17328;
assign v_17332 = v_17330 | v_17331;
assign v_17334 = v_17176 | v_17333;
assign v_17337 = v_17335 | v_17336;
assign v_17339 = v_17173 | v_17338;
assign v_17342 = v_17340 | v_17341;
assign v_17344 = v_17170 | v_17343;
assign v_17347 = v_17345 | v_17346;
assign v_17349 = v_17167 | v_17348;
assign v_17352 = v_17350 | v_17351;
assign v_17354 = v_17164 | v_17353;
assign v_17357 = v_17355 | v_17356;
assign v_17359 = v_17161 | v_17358;
assign v_17362 = v_17360 | v_17361;
assign v_17364 = v_17158 | v_17363;
assign v_17367 = v_17365 | v_17366;
assign v_17369 = v_17155 | v_17368;
assign v_17372 = v_17370 | v_17371;
assign v_17374 = v_17152 | v_17373;
assign v_17377 = v_17375 | v_17376;
assign v_17379 = v_17149 | v_17378;
assign v_17382 = v_17380 | v_17381;
assign v_17384 = v_17146 | v_17383;
assign v_17387 = v_17145 | v_17386;
assign v_17441 = v_17438 | v_17440;
assign v_17443 = v_17437 | v_17442;
assign v_17445 = v_17435 | v_17444;
assign v_17447 = v_17442 | v_17446;
assign v_17449 = v_17434 | v_17448;
assign v_17451 = v_17432 | v_17450;
assign v_17453 = v_17448 | v_17452;
assign v_17455 = v_17431 | v_17454;
assign v_17457 = v_17429 | v_17456;
assign v_17459 = v_17454 | v_17458;
assign v_17461 = v_17428 | v_17460;
assign v_17463 = v_17426 | v_17462;
assign v_17465 = v_17460 | v_17464;
assign v_17467 = v_17425 | v_17466;
assign v_17469 = v_17423 | v_17468;
assign v_17471 = v_17466 | v_17470;
assign v_17473 = v_17422 | v_17472;
assign v_17475 = v_17420 | v_17474;
assign v_17477 = v_17472 | v_17476;
assign v_17479 = v_17419 | v_17478;
assign v_17481 = v_17417 | v_17480;
assign v_17483 = v_17478 | v_17482;
assign v_17485 = v_17416 | v_17484;
assign v_17487 = v_17414 | v_17486;
assign v_17489 = v_17484 | v_17488;
assign v_17491 = v_17413 | v_17490;
assign v_17493 = v_17411 | v_17492;
assign v_17495 = v_17490 | v_17494;
assign v_17497 = v_17410 | v_17496;
assign v_17499 = v_17408 | v_17498;
assign v_17501 = v_17496 | v_17500;
assign v_17503 = v_17407 | v_17502;
assign v_17505 = v_17405 | v_17504;
assign v_17507 = v_17502 | v_17506;
assign v_17509 = v_17404 | v_17508;
assign v_17511 = v_17402 | v_17510;
assign v_17513 = v_17508 | v_17512;
assign v_17515 = v_17401 | v_17514;
assign v_17517 = v_17399 | v_17516;
assign v_17519 = v_17514 | v_17518;
assign v_17521 = v_17398 | v_17520;
assign v_17523 = v_17396 | v_17522;
assign v_17525 = v_17520 | v_17524;
assign v_17527 = v_17395 | v_17526;
assign v_17529 = v_17393 | v_17528;
assign v_17531 = v_17526 | v_17530;
assign v_17533 = v_17392 | v_17532;
assign v_17535 = v_17390 | v_17534;
assign v_17537 = v_17532 | v_17536;
assign v_17540 = ~v_17389 | v_17539;
assign v_17547 = v_17437 | v_17546;
assign v_17550 = v_17548 | v_17549;
assign v_17552 = v_17434 | v_17551;
assign v_17555 = v_17553 | v_17554;
assign v_17557 = v_17431 | v_17556;
assign v_17560 = v_17558 | v_17559;
assign v_17562 = v_17428 | v_17561;
assign v_17565 = v_17563 | v_17564;
assign v_17567 = v_17425 | v_17566;
assign v_17570 = v_17568 | v_17569;
assign v_17572 = v_17422 | v_17571;
assign v_17575 = v_17573 | v_17574;
assign v_17577 = v_17419 | v_17576;
assign v_17580 = v_17578 | v_17579;
assign v_17582 = v_17416 | v_17581;
assign v_17585 = v_17583 | v_17584;
assign v_17587 = v_17413 | v_17586;
assign v_17590 = v_17588 | v_17589;
assign v_17592 = v_17410 | v_17591;
assign v_17595 = v_17593 | v_17594;
assign v_17597 = v_17407 | v_17596;
assign v_17600 = v_17598 | v_17599;
assign v_17602 = v_17404 | v_17601;
assign v_17605 = v_17603 | v_17604;
assign v_17607 = v_17401 | v_17606;
assign v_17610 = v_17608 | v_17609;
assign v_17612 = v_17398 | v_17611;
assign v_17615 = v_17613 | v_17614;
assign v_17617 = v_17395 | v_17616;
assign v_17620 = v_17618 | v_17619;
assign v_17622 = v_17392 | v_17621;
assign v_17625 = v_17623 | v_17624;
assign v_17627 = v_17389 | v_17626;
assign v_17630 = v_17388 | v_17629;
assign v_17684 = v_17681 | v_17683;
assign v_17686 = v_17680 | v_17685;
assign v_17688 = v_17678 | v_17687;
assign v_17690 = v_17685 | v_17689;
assign v_17692 = v_17677 | v_17691;
assign v_17694 = v_17675 | v_17693;
assign v_17696 = v_17691 | v_17695;
assign v_17698 = v_17674 | v_17697;
assign v_17700 = v_17672 | v_17699;
assign v_17702 = v_17697 | v_17701;
assign v_17704 = v_17671 | v_17703;
assign v_17706 = v_17669 | v_17705;
assign v_17708 = v_17703 | v_17707;
assign v_17710 = v_17668 | v_17709;
assign v_17712 = v_17666 | v_17711;
assign v_17714 = v_17709 | v_17713;
assign v_17716 = v_17665 | v_17715;
assign v_17718 = v_17663 | v_17717;
assign v_17720 = v_17715 | v_17719;
assign v_17722 = v_17662 | v_17721;
assign v_17724 = v_17660 | v_17723;
assign v_17726 = v_17721 | v_17725;
assign v_17728 = v_17659 | v_17727;
assign v_17730 = v_17657 | v_17729;
assign v_17732 = v_17727 | v_17731;
assign v_17734 = v_17656 | v_17733;
assign v_17736 = v_17654 | v_17735;
assign v_17738 = v_17733 | v_17737;
assign v_17740 = v_17653 | v_17739;
assign v_17742 = v_17651 | v_17741;
assign v_17744 = v_17739 | v_17743;
assign v_17746 = v_17650 | v_17745;
assign v_17748 = v_17648 | v_17747;
assign v_17750 = v_17745 | v_17749;
assign v_17752 = v_17647 | v_17751;
assign v_17754 = v_17645 | v_17753;
assign v_17756 = v_17751 | v_17755;
assign v_17758 = v_17644 | v_17757;
assign v_17760 = v_17642 | v_17759;
assign v_17762 = v_17757 | v_17761;
assign v_17764 = v_17641 | v_17763;
assign v_17766 = v_17639 | v_17765;
assign v_17768 = v_17763 | v_17767;
assign v_17770 = v_17638 | v_17769;
assign v_17772 = v_17636 | v_17771;
assign v_17774 = v_17769 | v_17773;
assign v_17776 = v_17635 | v_17775;
assign v_17778 = v_17633 | v_17777;
assign v_17780 = v_17775 | v_17779;
assign v_17783 = ~v_17632 | v_17782;
assign v_17790 = v_17680 | v_17789;
assign v_17793 = v_17791 | v_17792;
assign v_17795 = v_17677 | v_17794;
assign v_17798 = v_17796 | v_17797;
assign v_17800 = v_17674 | v_17799;
assign v_17803 = v_17801 | v_17802;
assign v_17805 = v_17671 | v_17804;
assign v_17808 = v_17806 | v_17807;
assign v_17810 = v_17668 | v_17809;
assign v_17813 = v_17811 | v_17812;
assign v_17815 = v_17665 | v_17814;
assign v_17818 = v_17816 | v_17817;
assign v_17820 = v_17662 | v_17819;
assign v_17823 = v_17821 | v_17822;
assign v_17825 = v_17659 | v_17824;
assign v_17828 = v_17826 | v_17827;
assign v_17830 = v_17656 | v_17829;
assign v_17833 = v_17831 | v_17832;
assign v_17835 = v_17653 | v_17834;
assign v_17838 = v_17836 | v_17837;
assign v_17840 = v_17650 | v_17839;
assign v_17843 = v_17841 | v_17842;
assign v_17845 = v_17647 | v_17844;
assign v_17848 = v_17846 | v_17847;
assign v_17850 = v_17644 | v_17849;
assign v_17853 = v_17851 | v_17852;
assign v_17855 = v_17641 | v_17854;
assign v_17858 = v_17856 | v_17857;
assign v_17860 = v_17638 | v_17859;
assign v_17863 = v_17861 | v_17862;
assign v_17865 = v_17635 | v_17864;
assign v_17868 = v_17866 | v_17867;
assign v_17870 = v_17632 | v_17869;
assign v_17873 = v_17631 | v_17872;
assign v_17927 = v_17924 | v_17926;
assign v_17929 = v_17923 | v_17928;
assign v_17931 = v_17921 | v_17930;
assign v_17933 = v_17928 | v_17932;
assign v_17935 = v_17920 | v_17934;
assign v_17937 = v_17918 | v_17936;
assign v_17939 = v_17934 | v_17938;
assign v_17941 = v_17917 | v_17940;
assign v_17943 = v_17915 | v_17942;
assign v_17945 = v_17940 | v_17944;
assign v_17947 = v_17914 | v_17946;
assign v_17949 = v_17912 | v_17948;
assign v_17951 = v_17946 | v_17950;
assign v_17953 = v_17911 | v_17952;
assign v_17955 = v_17909 | v_17954;
assign v_17957 = v_17952 | v_17956;
assign v_17959 = v_17908 | v_17958;
assign v_17961 = v_17906 | v_17960;
assign v_17963 = v_17958 | v_17962;
assign v_17965 = v_17905 | v_17964;
assign v_17967 = v_17903 | v_17966;
assign v_17969 = v_17964 | v_17968;
assign v_17971 = v_17902 | v_17970;
assign v_17973 = v_17900 | v_17972;
assign v_17975 = v_17970 | v_17974;
assign v_17977 = v_17899 | v_17976;
assign v_17979 = v_17897 | v_17978;
assign v_17981 = v_17976 | v_17980;
assign v_17983 = v_17896 | v_17982;
assign v_17985 = v_17894 | v_17984;
assign v_17987 = v_17982 | v_17986;
assign v_17989 = v_17893 | v_17988;
assign v_17991 = v_17891 | v_17990;
assign v_17993 = v_17988 | v_17992;
assign v_17995 = v_17890 | v_17994;
assign v_17997 = v_17888 | v_17996;
assign v_17999 = v_17994 | v_17998;
assign v_18001 = v_17887 | v_18000;
assign v_18003 = v_17885 | v_18002;
assign v_18005 = v_18000 | v_18004;
assign v_18007 = v_17884 | v_18006;
assign v_18009 = v_17882 | v_18008;
assign v_18011 = v_18006 | v_18010;
assign v_18013 = v_17881 | v_18012;
assign v_18015 = v_17879 | v_18014;
assign v_18017 = v_18012 | v_18016;
assign v_18019 = v_17878 | v_18018;
assign v_18021 = v_17876 | v_18020;
assign v_18023 = v_18018 | v_18022;
assign v_18026 = ~v_17875 | v_18025;
assign v_18033 = v_17923 | v_18032;
assign v_18036 = v_18034 | v_18035;
assign v_18038 = v_17920 | v_18037;
assign v_18041 = v_18039 | v_18040;
assign v_18043 = v_17917 | v_18042;
assign v_18046 = v_18044 | v_18045;
assign v_18048 = v_17914 | v_18047;
assign v_18051 = v_18049 | v_18050;
assign v_18053 = v_17911 | v_18052;
assign v_18056 = v_18054 | v_18055;
assign v_18058 = v_17908 | v_18057;
assign v_18061 = v_18059 | v_18060;
assign v_18063 = v_17905 | v_18062;
assign v_18066 = v_18064 | v_18065;
assign v_18068 = v_17902 | v_18067;
assign v_18071 = v_18069 | v_18070;
assign v_18073 = v_17899 | v_18072;
assign v_18076 = v_18074 | v_18075;
assign v_18078 = v_17896 | v_18077;
assign v_18081 = v_18079 | v_18080;
assign v_18083 = v_17893 | v_18082;
assign v_18086 = v_18084 | v_18085;
assign v_18088 = v_17890 | v_18087;
assign v_18091 = v_18089 | v_18090;
assign v_18093 = v_17887 | v_18092;
assign v_18096 = v_18094 | v_18095;
assign v_18098 = v_17884 | v_18097;
assign v_18101 = v_18099 | v_18100;
assign v_18103 = v_17881 | v_18102;
assign v_18106 = v_18104 | v_18105;
assign v_18108 = v_17878 | v_18107;
assign v_18111 = v_18109 | v_18110;
assign v_18113 = v_17875 | v_18112;
assign v_18116 = v_17874 | v_18115;
assign v_18170 = v_18167 | v_18169;
assign v_18172 = v_18166 | v_18171;
assign v_18174 = v_18164 | v_18173;
assign v_18176 = v_18171 | v_18175;
assign v_18178 = v_18163 | v_18177;
assign v_18180 = v_18161 | v_18179;
assign v_18182 = v_18177 | v_18181;
assign v_18184 = v_18160 | v_18183;
assign v_18186 = v_18158 | v_18185;
assign v_18188 = v_18183 | v_18187;
assign v_18190 = v_18157 | v_18189;
assign v_18192 = v_18155 | v_18191;
assign v_18194 = v_18189 | v_18193;
assign v_18196 = v_18154 | v_18195;
assign v_18198 = v_18152 | v_18197;
assign v_18200 = v_18195 | v_18199;
assign v_18202 = v_18151 | v_18201;
assign v_18204 = v_18149 | v_18203;
assign v_18206 = v_18201 | v_18205;
assign v_18208 = v_18148 | v_18207;
assign v_18210 = v_18146 | v_18209;
assign v_18212 = v_18207 | v_18211;
assign v_18214 = v_18145 | v_18213;
assign v_18216 = v_18143 | v_18215;
assign v_18218 = v_18213 | v_18217;
assign v_18220 = v_18142 | v_18219;
assign v_18222 = v_18140 | v_18221;
assign v_18224 = v_18219 | v_18223;
assign v_18226 = v_18139 | v_18225;
assign v_18228 = v_18137 | v_18227;
assign v_18230 = v_18225 | v_18229;
assign v_18232 = v_18136 | v_18231;
assign v_18234 = v_18134 | v_18233;
assign v_18236 = v_18231 | v_18235;
assign v_18238 = v_18133 | v_18237;
assign v_18240 = v_18131 | v_18239;
assign v_18242 = v_18237 | v_18241;
assign v_18244 = v_18130 | v_18243;
assign v_18246 = v_18128 | v_18245;
assign v_18248 = v_18243 | v_18247;
assign v_18250 = v_18127 | v_18249;
assign v_18252 = v_18125 | v_18251;
assign v_18254 = v_18249 | v_18253;
assign v_18256 = v_18124 | v_18255;
assign v_18258 = v_18122 | v_18257;
assign v_18260 = v_18255 | v_18259;
assign v_18262 = v_18121 | v_18261;
assign v_18264 = v_18119 | v_18263;
assign v_18266 = v_18261 | v_18265;
assign v_18269 = ~v_18118 | v_18268;
assign v_18276 = v_18166 | v_18275;
assign v_18279 = v_18277 | v_18278;
assign v_18281 = v_18163 | v_18280;
assign v_18284 = v_18282 | v_18283;
assign v_18286 = v_18160 | v_18285;
assign v_18289 = v_18287 | v_18288;
assign v_18291 = v_18157 | v_18290;
assign v_18294 = v_18292 | v_18293;
assign v_18296 = v_18154 | v_18295;
assign v_18299 = v_18297 | v_18298;
assign v_18301 = v_18151 | v_18300;
assign v_18304 = v_18302 | v_18303;
assign v_18306 = v_18148 | v_18305;
assign v_18309 = v_18307 | v_18308;
assign v_18311 = v_18145 | v_18310;
assign v_18314 = v_18312 | v_18313;
assign v_18316 = v_18142 | v_18315;
assign v_18319 = v_18317 | v_18318;
assign v_18321 = v_18139 | v_18320;
assign v_18324 = v_18322 | v_18323;
assign v_18326 = v_18136 | v_18325;
assign v_18329 = v_18327 | v_18328;
assign v_18331 = v_18133 | v_18330;
assign v_18334 = v_18332 | v_18333;
assign v_18336 = v_18130 | v_18335;
assign v_18339 = v_18337 | v_18338;
assign v_18341 = v_18127 | v_18340;
assign v_18344 = v_18342 | v_18343;
assign v_18346 = v_18124 | v_18345;
assign v_18349 = v_18347 | v_18348;
assign v_18351 = v_18121 | v_18350;
assign v_18354 = v_18352 | v_18353;
assign v_18356 = v_18118 | v_18355;
assign v_18359 = v_18117 | v_18358;
assign v_18413 = v_18410 | v_18412;
assign v_18415 = v_18409 | v_18414;
assign v_18417 = v_18407 | v_18416;
assign v_18419 = v_18414 | v_18418;
assign v_18421 = v_18406 | v_18420;
assign v_18423 = v_18404 | v_18422;
assign v_18425 = v_18420 | v_18424;
assign v_18427 = v_18403 | v_18426;
assign v_18429 = v_18401 | v_18428;
assign v_18431 = v_18426 | v_18430;
assign v_18433 = v_18400 | v_18432;
assign v_18435 = v_18398 | v_18434;
assign v_18437 = v_18432 | v_18436;
assign v_18439 = v_18397 | v_18438;
assign v_18441 = v_18395 | v_18440;
assign v_18443 = v_18438 | v_18442;
assign v_18445 = v_18394 | v_18444;
assign v_18447 = v_18392 | v_18446;
assign v_18449 = v_18444 | v_18448;
assign v_18451 = v_18391 | v_18450;
assign v_18453 = v_18389 | v_18452;
assign v_18455 = v_18450 | v_18454;
assign v_18457 = v_18388 | v_18456;
assign v_18459 = v_18386 | v_18458;
assign v_18461 = v_18456 | v_18460;
assign v_18463 = v_18385 | v_18462;
assign v_18465 = v_18383 | v_18464;
assign v_18467 = v_18462 | v_18466;
assign v_18469 = v_18382 | v_18468;
assign v_18471 = v_18380 | v_18470;
assign v_18473 = v_18468 | v_18472;
assign v_18475 = v_18379 | v_18474;
assign v_18477 = v_18377 | v_18476;
assign v_18479 = v_18474 | v_18478;
assign v_18481 = v_18376 | v_18480;
assign v_18483 = v_18374 | v_18482;
assign v_18485 = v_18480 | v_18484;
assign v_18487 = v_18373 | v_18486;
assign v_18489 = v_18371 | v_18488;
assign v_18491 = v_18486 | v_18490;
assign v_18493 = v_18370 | v_18492;
assign v_18495 = v_18368 | v_18494;
assign v_18497 = v_18492 | v_18496;
assign v_18499 = v_18367 | v_18498;
assign v_18501 = v_18365 | v_18500;
assign v_18503 = v_18498 | v_18502;
assign v_18505 = v_18364 | v_18504;
assign v_18507 = v_18362 | v_18506;
assign v_18509 = v_18504 | v_18508;
assign v_18512 = ~v_18361 | v_18511;
assign v_18519 = v_18409 | v_18518;
assign v_18522 = v_18520 | v_18521;
assign v_18524 = v_18406 | v_18523;
assign v_18527 = v_18525 | v_18526;
assign v_18529 = v_18403 | v_18528;
assign v_18532 = v_18530 | v_18531;
assign v_18534 = v_18400 | v_18533;
assign v_18537 = v_18535 | v_18536;
assign v_18539 = v_18397 | v_18538;
assign v_18542 = v_18540 | v_18541;
assign v_18544 = v_18394 | v_18543;
assign v_18547 = v_18545 | v_18546;
assign v_18549 = v_18391 | v_18548;
assign v_18552 = v_18550 | v_18551;
assign v_18554 = v_18388 | v_18553;
assign v_18557 = v_18555 | v_18556;
assign v_18559 = v_18385 | v_18558;
assign v_18562 = v_18560 | v_18561;
assign v_18564 = v_18382 | v_18563;
assign v_18567 = v_18565 | v_18566;
assign v_18569 = v_18379 | v_18568;
assign v_18572 = v_18570 | v_18571;
assign v_18574 = v_18376 | v_18573;
assign v_18577 = v_18575 | v_18576;
assign v_18579 = v_18373 | v_18578;
assign v_18582 = v_18580 | v_18581;
assign v_18584 = v_18370 | v_18583;
assign v_18587 = v_18585 | v_18586;
assign v_18589 = v_18367 | v_18588;
assign v_18592 = v_18590 | v_18591;
assign v_18594 = v_18364 | v_18593;
assign v_18597 = v_18595 | v_18596;
assign v_18599 = v_18361 | v_18598;
assign v_18602 = v_18360 | v_18601;
assign v_18656 = v_18653 | v_18655;
assign v_18658 = v_18652 | v_18657;
assign v_18660 = v_18650 | v_18659;
assign v_18662 = v_18657 | v_18661;
assign v_18664 = v_18649 | v_18663;
assign v_18666 = v_18647 | v_18665;
assign v_18668 = v_18663 | v_18667;
assign v_18670 = v_18646 | v_18669;
assign v_18672 = v_18644 | v_18671;
assign v_18674 = v_18669 | v_18673;
assign v_18676 = v_18643 | v_18675;
assign v_18678 = v_18641 | v_18677;
assign v_18680 = v_18675 | v_18679;
assign v_18682 = v_18640 | v_18681;
assign v_18684 = v_18638 | v_18683;
assign v_18686 = v_18681 | v_18685;
assign v_18688 = v_18637 | v_18687;
assign v_18690 = v_18635 | v_18689;
assign v_18692 = v_18687 | v_18691;
assign v_18694 = v_18634 | v_18693;
assign v_18696 = v_18632 | v_18695;
assign v_18698 = v_18693 | v_18697;
assign v_18700 = v_18631 | v_18699;
assign v_18702 = v_18629 | v_18701;
assign v_18704 = v_18699 | v_18703;
assign v_18706 = v_18628 | v_18705;
assign v_18708 = v_18626 | v_18707;
assign v_18710 = v_18705 | v_18709;
assign v_18712 = v_18625 | v_18711;
assign v_18714 = v_18623 | v_18713;
assign v_18716 = v_18711 | v_18715;
assign v_18718 = v_18622 | v_18717;
assign v_18720 = v_18620 | v_18719;
assign v_18722 = v_18717 | v_18721;
assign v_18724 = v_18619 | v_18723;
assign v_18726 = v_18617 | v_18725;
assign v_18728 = v_18723 | v_18727;
assign v_18730 = v_18616 | v_18729;
assign v_18732 = v_18614 | v_18731;
assign v_18734 = v_18729 | v_18733;
assign v_18736 = v_18613 | v_18735;
assign v_18738 = v_18611 | v_18737;
assign v_18740 = v_18735 | v_18739;
assign v_18742 = v_18610 | v_18741;
assign v_18744 = v_18608 | v_18743;
assign v_18746 = v_18741 | v_18745;
assign v_18748 = v_18607 | v_18747;
assign v_18750 = v_18605 | v_18749;
assign v_18752 = v_18747 | v_18751;
assign v_18755 = ~v_18604 | v_18754;
assign v_18762 = v_18652 | v_18761;
assign v_18765 = v_18763 | v_18764;
assign v_18767 = v_18649 | v_18766;
assign v_18770 = v_18768 | v_18769;
assign v_18772 = v_18646 | v_18771;
assign v_18775 = v_18773 | v_18774;
assign v_18777 = v_18643 | v_18776;
assign v_18780 = v_18778 | v_18779;
assign v_18782 = v_18640 | v_18781;
assign v_18785 = v_18783 | v_18784;
assign v_18787 = v_18637 | v_18786;
assign v_18790 = v_18788 | v_18789;
assign v_18792 = v_18634 | v_18791;
assign v_18795 = v_18793 | v_18794;
assign v_18797 = v_18631 | v_18796;
assign v_18800 = v_18798 | v_18799;
assign v_18802 = v_18628 | v_18801;
assign v_18805 = v_18803 | v_18804;
assign v_18807 = v_18625 | v_18806;
assign v_18810 = v_18808 | v_18809;
assign v_18812 = v_18622 | v_18811;
assign v_18815 = v_18813 | v_18814;
assign v_18817 = v_18619 | v_18816;
assign v_18820 = v_18818 | v_18819;
assign v_18822 = v_18616 | v_18821;
assign v_18825 = v_18823 | v_18824;
assign v_18827 = v_18613 | v_18826;
assign v_18830 = v_18828 | v_18829;
assign v_18832 = v_18610 | v_18831;
assign v_18835 = v_18833 | v_18834;
assign v_18837 = v_18607 | v_18836;
assign v_18840 = v_18838 | v_18839;
assign v_18842 = v_18604 | v_18841;
assign v_18845 = v_18603 | v_18844;
assign v_18899 = v_18896 | v_18898;
assign v_18901 = v_18895 | v_18900;
assign v_18903 = v_18893 | v_18902;
assign v_18905 = v_18900 | v_18904;
assign v_18907 = v_18892 | v_18906;
assign v_18909 = v_18890 | v_18908;
assign v_18911 = v_18906 | v_18910;
assign v_18913 = v_18889 | v_18912;
assign v_18915 = v_18887 | v_18914;
assign v_18917 = v_18912 | v_18916;
assign v_18919 = v_18886 | v_18918;
assign v_18921 = v_18884 | v_18920;
assign v_18923 = v_18918 | v_18922;
assign v_18925 = v_18883 | v_18924;
assign v_18927 = v_18881 | v_18926;
assign v_18929 = v_18924 | v_18928;
assign v_18931 = v_18880 | v_18930;
assign v_18933 = v_18878 | v_18932;
assign v_18935 = v_18930 | v_18934;
assign v_18937 = v_18877 | v_18936;
assign v_18939 = v_18875 | v_18938;
assign v_18941 = v_18936 | v_18940;
assign v_18943 = v_18874 | v_18942;
assign v_18945 = v_18872 | v_18944;
assign v_18947 = v_18942 | v_18946;
assign v_18949 = v_18871 | v_18948;
assign v_18951 = v_18869 | v_18950;
assign v_18953 = v_18948 | v_18952;
assign v_18955 = v_18868 | v_18954;
assign v_18957 = v_18866 | v_18956;
assign v_18959 = v_18954 | v_18958;
assign v_18961 = v_18865 | v_18960;
assign v_18963 = v_18863 | v_18962;
assign v_18965 = v_18960 | v_18964;
assign v_18967 = v_18862 | v_18966;
assign v_18969 = v_18860 | v_18968;
assign v_18971 = v_18966 | v_18970;
assign v_18973 = v_18859 | v_18972;
assign v_18975 = v_18857 | v_18974;
assign v_18977 = v_18972 | v_18976;
assign v_18979 = v_18856 | v_18978;
assign v_18981 = v_18854 | v_18980;
assign v_18983 = v_18978 | v_18982;
assign v_18985 = v_18853 | v_18984;
assign v_18987 = v_18851 | v_18986;
assign v_18989 = v_18984 | v_18988;
assign v_18991 = v_18850 | v_18990;
assign v_18993 = v_18848 | v_18992;
assign v_18995 = v_18990 | v_18994;
assign v_18998 = ~v_18847 | v_18997;
assign v_19005 = v_18895 | v_19004;
assign v_19008 = v_19006 | v_19007;
assign v_19010 = v_18892 | v_19009;
assign v_19013 = v_19011 | v_19012;
assign v_19015 = v_18889 | v_19014;
assign v_19018 = v_19016 | v_19017;
assign v_19020 = v_18886 | v_19019;
assign v_19023 = v_19021 | v_19022;
assign v_19025 = v_18883 | v_19024;
assign v_19028 = v_19026 | v_19027;
assign v_19030 = v_18880 | v_19029;
assign v_19033 = v_19031 | v_19032;
assign v_19035 = v_18877 | v_19034;
assign v_19038 = v_19036 | v_19037;
assign v_19040 = v_18874 | v_19039;
assign v_19043 = v_19041 | v_19042;
assign v_19045 = v_18871 | v_19044;
assign v_19048 = v_19046 | v_19047;
assign v_19050 = v_18868 | v_19049;
assign v_19053 = v_19051 | v_19052;
assign v_19055 = v_18865 | v_19054;
assign v_19058 = v_19056 | v_19057;
assign v_19060 = v_18862 | v_19059;
assign v_19063 = v_19061 | v_19062;
assign v_19065 = v_18859 | v_19064;
assign v_19068 = v_19066 | v_19067;
assign v_19070 = v_18856 | v_19069;
assign v_19073 = v_19071 | v_19072;
assign v_19075 = v_18853 | v_19074;
assign v_19078 = v_19076 | v_19077;
assign v_19080 = v_18850 | v_19079;
assign v_19083 = v_19081 | v_19082;
assign v_19085 = v_18847 | v_19084;
assign v_19088 = v_18846 | v_19087;
assign v_19142 = v_19139 | v_19141;
assign v_19144 = v_19138 | v_19143;
assign v_19146 = v_19136 | v_19145;
assign v_19148 = v_19143 | v_19147;
assign v_19150 = v_19135 | v_19149;
assign v_19152 = v_19133 | v_19151;
assign v_19154 = v_19149 | v_19153;
assign v_19156 = v_19132 | v_19155;
assign v_19158 = v_19130 | v_19157;
assign v_19160 = v_19155 | v_19159;
assign v_19162 = v_19129 | v_19161;
assign v_19164 = v_19127 | v_19163;
assign v_19166 = v_19161 | v_19165;
assign v_19168 = v_19126 | v_19167;
assign v_19170 = v_19124 | v_19169;
assign v_19172 = v_19167 | v_19171;
assign v_19174 = v_19123 | v_19173;
assign v_19176 = v_19121 | v_19175;
assign v_19178 = v_19173 | v_19177;
assign v_19180 = v_19120 | v_19179;
assign v_19182 = v_19118 | v_19181;
assign v_19184 = v_19179 | v_19183;
assign v_19186 = v_19117 | v_19185;
assign v_19188 = v_19115 | v_19187;
assign v_19190 = v_19185 | v_19189;
assign v_19192 = v_19114 | v_19191;
assign v_19194 = v_19112 | v_19193;
assign v_19196 = v_19191 | v_19195;
assign v_19198 = v_19111 | v_19197;
assign v_19200 = v_19109 | v_19199;
assign v_19202 = v_19197 | v_19201;
assign v_19204 = v_19108 | v_19203;
assign v_19206 = v_19106 | v_19205;
assign v_19208 = v_19203 | v_19207;
assign v_19210 = v_19105 | v_19209;
assign v_19212 = v_19103 | v_19211;
assign v_19214 = v_19209 | v_19213;
assign v_19216 = v_19102 | v_19215;
assign v_19218 = v_19100 | v_19217;
assign v_19220 = v_19215 | v_19219;
assign v_19222 = v_19099 | v_19221;
assign v_19224 = v_19097 | v_19223;
assign v_19226 = v_19221 | v_19225;
assign v_19228 = v_19096 | v_19227;
assign v_19230 = v_19094 | v_19229;
assign v_19232 = v_19227 | v_19231;
assign v_19234 = v_19093 | v_19233;
assign v_19236 = v_19091 | v_19235;
assign v_19238 = v_19233 | v_19237;
assign v_19241 = ~v_19090 | v_19240;
assign v_19248 = v_19138 | v_19247;
assign v_19251 = v_19249 | v_19250;
assign v_19253 = v_19135 | v_19252;
assign v_19256 = v_19254 | v_19255;
assign v_19258 = v_19132 | v_19257;
assign v_19261 = v_19259 | v_19260;
assign v_19263 = v_19129 | v_19262;
assign v_19266 = v_19264 | v_19265;
assign v_19268 = v_19126 | v_19267;
assign v_19271 = v_19269 | v_19270;
assign v_19273 = v_19123 | v_19272;
assign v_19276 = v_19274 | v_19275;
assign v_19278 = v_19120 | v_19277;
assign v_19281 = v_19279 | v_19280;
assign v_19283 = v_19117 | v_19282;
assign v_19286 = v_19284 | v_19285;
assign v_19288 = v_19114 | v_19287;
assign v_19291 = v_19289 | v_19290;
assign v_19293 = v_19111 | v_19292;
assign v_19296 = v_19294 | v_19295;
assign v_19298 = v_19108 | v_19297;
assign v_19301 = v_19299 | v_19300;
assign v_19303 = v_19105 | v_19302;
assign v_19306 = v_19304 | v_19305;
assign v_19308 = v_19102 | v_19307;
assign v_19311 = v_19309 | v_19310;
assign v_19313 = v_19099 | v_19312;
assign v_19316 = v_19314 | v_19315;
assign v_19318 = v_19096 | v_19317;
assign v_19321 = v_19319 | v_19320;
assign v_19323 = v_19093 | v_19322;
assign v_19326 = v_19324 | v_19325;
assign v_19328 = v_19090 | v_19327;
assign v_19331 = v_19089 | v_19330;
assign v_19385 = v_19382 | v_19384;
assign v_19387 = v_19381 | v_19386;
assign v_19389 = v_19379 | v_19388;
assign v_19391 = v_19386 | v_19390;
assign v_19393 = v_19378 | v_19392;
assign v_19395 = v_19376 | v_19394;
assign v_19397 = v_19392 | v_19396;
assign v_19399 = v_19375 | v_19398;
assign v_19401 = v_19373 | v_19400;
assign v_19403 = v_19398 | v_19402;
assign v_19405 = v_19372 | v_19404;
assign v_19407 = v_19370 | v_19406;
assign v_19409 = v_19404 | v_19408;
assign v_19411 = v_19369 | v_19410;
assign v_19413 = v_19367 | v_19412;
assign v_19415 = v_19410 | v_19414;
assign v_19417 = v_19366 | v_19416;
assign v_19419 = v_19364 | v_19418;
assign v_19421 = v_19416 | v_19420;
assign v_19423 = v_19363 | v_19422;
assign v_19425 = v_19361 | v_19424;
assign v_19427 = v_19422 | v_19426;
assign v_19429 = v_19360 | v_19428;
assign v_19431 = v_19358 | v_19430;
assign v_19433 = v_19428 | v_19432;
assign v_19435 = v_19357 | v_19434;
assign v_19437 = v_19355 | v_19436;
assign v_19439 = v_19434 | v_19438;
assign v_19441 = v_19354 | v_19440;
assign v_19443 = v_19352 | v_19442;
assign v_19445 = v_19440 | v_19444;
assign v_19447 = v_19351 | v_19446;
assign v_19449 = v_19349 | v_19448;
assign v_19451 = v_19446 | v_19450;
assign v_19453 = v_19348 | v_19452;
assign v_19455 = v_19346 | v_19454;
assign v_19457 = v_19452 | v_19456;
assign v_19459 = v_19345 | v_19458;
assign v_19461 = v_19343 | v_19460;
assign v_19463 = v_19458 | v_19462;
assign v_19465 = v_19342 | v_19464;
assign v_19467 = v_19340 | v_19466;
assign v_19469 = v_19464 | v_19468;
assign v_19471 = v_19339 | v_19470;
assign v_19473 = v_19337 | v_19472;
assign v_19475 = v_19470 | v_19474;
assign v_19477 = v_19336 | v_19476;
assign v_19479 = v_19334 | v_19478;
assign v_19481 = v_19476 | v_19480;
assign v_19484 = ~v_19333 | v_19483;
assign v_19491 = v_19381 | v_19490;
assign v_19494 = v_19492 | v_19493;
assign v_19496 = v_19378 | v_19495;
assign v_19499 = v_19497 | v_19498;
assign v_19501 = v_19375 | v_19500;
assign v_19504 = v_19502 | v_19503;
assign v_19506 = v_19372 | v_19505;
assign v_19509 = v_19507 | v_19508;
assign v_19511 = v_19369 | v_19510;
assign v_19514 = v_19512 | v_19513;
assign v_19516 = v_19366 | v_19515;
assign v_19519 = v_19517 | v_19518;
assign v_19521 = v_19363 | v_19520;
assign v_19524 = v_19522 | v_19523;
assign v_19526 = v_19360 | v_19525;
assign v_19529 = v_19527 | v_19528;
assign v_19531 = v_19357 | v_19530;
assign v_19534 = v_19532 | v_19533;
assign v_19536 = v_19354 | v_19535;
assign v_19539 = v_19537 | v_19538;
assign v_19541 = v_19351 | v_19540;
assign v_19544 = v_19542 | v_19543;
assign v_19546 = v_19348 | v_19545;
assign v_19549 = v_19547 | v_19548;
assign v_19551 = v_19345 | v_19550;
assign v_19554 = v_19552 | v_19553;
assign v_19556 = v_19342 | v_19555;
assign v_19559 = v_19557 | v_19558;
assign v_19561 = v_19339 | v_19560;
assign v_19564 = v_19562 | v_19563;
assign v_19566 = v_19336 | v_19565;
assign v_19569 = v_19567 | v_19568;
assign v_19571 = v_19333 | v_19570;
assign v_19574 = v_19332 | v_19573;
assign v_19628 = v_19625 | v_19627;
assign v_19630 = v_19624 | v_19629;
assign v_19632 = v_19622 | v_19631;
assign v_19634 = v_19629 | v_19633;
assign v_19636 = v_19621 | v_19635;
assign v_19638 = v_19619 | v_19637;
assign v_19640 = v_19635 | v_19639;
assign v_19642 = v_19618 | v_19641;
assign v_19644 = v_19616 | v_19643;
assign v_19646 = v_19641 | v_19645;
assign v_19648 = v_19615 | v_19647;
assign v_19650 = v_19613 | v_19649;
assign v_19652 = v_19647 | v_19651;
assign v_19654 = v_19612 | v_19653;
assign v_19656 = v_19610 | v_19655;
assign v_19658 = v_19653 | v_19657;
assign v_19660 = v_19609 | v_19659;
assign v_19662 = v_19607 | v_19661;
assign v_19664 = v_19659 | v_19663;
assign v_19666 = v_19606 | v_19665;
assign v_19668 = v_19604 | v_19667;
assign v_19670 = v_19665 | v_19669;
assign v_19672 = v_19603 | v_19671;
assign v_19674 = v_19601 | v_19673;
assign v_19676 = v_19671 | v_19675;
assign v_19678 = v_19600 | v_19677;
assign v_19680 = v_19598 | v_19679;
assign v_19682 = v_19677 | v_19681;
assign v_19684 = v_19597 | v_19683;
assign v_19686 = v_19595 | v_19685;
assign v_19688 = v_19683 | v_19687;
assign v_19690 = v_19594 | v_19689;
assign v_19692 = v_19592 | v_19691;
assign v_19694 = v_19689 | v_19693;
assign v_19696 = v_19591 | v_19695;
assign v_19698 = v_19589 | v_19697;
assign v_19700 = v_19695 | v_19699;
assign v_19702 = v_19588 | v_19701;
assign v_19704 = v_19586 | v_19703;
assign v_19706 = v_19701 | v_19705;
assign v_19708 = v_19585 | v_19707;
assign v_19710 = v_19583 | v_19709;
assign v_19712 = v_19707 | v_19711;
assign v_19714 = v_19582 | v_19713;
assign v_19716 = v_19580 | v_19715;
assign v_19718 = v_19713 | v_19717;
assign v_19720 = v_19579 | v_19719;
assign v_19722 = v_19577 | v_19721;
assign v_19724 = v_19719 | v_19723;
assign v_19727 = ~v_19576 | v_19726;
assign v_19734 = v_19624 | v_19733;
assign v_19737 = v_19735 | v_19736;
assign v_19739 = v_19621 | v_19738;
assign v_19742 = v_19740 | v_19741;
assign v_19744 = v_19618 | v_19743;
assign v_19747 = v_19745 | v_19746;
assign v_19749 = v_19615 | v_19748;
assign v_19752 = v_19750 | v_19751;
assign v_19754 = v_19612 | v_19753;
assign v_19757 = v_19755 | v_19756;
assign v_19759 = v_19609 | v_19758;
assign v_19762 = v_19760 | v_19761;
assign v_19764 = v_19606 | v_19763;
assign v_19767 = v_19765 | v_19766;
assign v_19769 = v_19603 | v_19768;
assign v_19772 = v_19770 | v_19771;
assign v_19774 = v_19600 | v_19773;
assign v_19777 = v_19775 | v_19776;
assign v_19779 = v_19597 | v_19778;
assign v_19782 = v_19780 | v_19781;
assign v_19784 = v_19594 | v_19783;
assign v_19787 = v_19785 | v_19786;
assign v_19789 = v_19591 | v_19788;
assign v_19792 = v_19790 | v_19791;
assign v_19794 = v_19588 | v_19793;
assign v_19797 = v_19795 | v_19796;
assign v_19799 = v_19585 | v_19798;
assign v_19802 = v_19800 | v_19801;
assign v_19804 = v_19582 | v_19803;
assign v_19807 = v_19805 | v_19806;
assign v_19809 = v_19579 | v_19808;
assign v_19812 = v_19810 | v_19811;
assign v_19814 = v_19576 | v_19813;
assign v_19817 = v_19575 | v_19816;
assign v_19871 = v_19868 | v_19870;
assign v_19873 = v_19867 | v_19872;
assign v_19875 = v_19865 | v_19874;
assign v_19877 = v_19872 | v_19876;
assign v_19879 = v_19864 | v_19878;
assign v_19881 = v_19862 | v_19880;
assign v_19883 = v_19878 | v_19882;
assign v_19885 = v_19861 | v_19884;
assign v_19887 = v_19859 | v_19886;
assign v_19889 = v_19884 | v_19888;
assign v_19891 = v_19858 | v_19890;
assign v_19893 = v_19856 | v_19892;
assign v_19895 = v_19890 | v_19894;
assign v_19897 = v_19855 | v_19896;
assign v_19899 = v_19853 | v_19898;
assign v_19901 = v_19896 | v_19900;
assign v_19903 = v_19852 | v_19902;
assign v_19905 = v_19850 | v_19904;
assign v_19907 = v_19902 | v_19906;
assign v_19909 = v_19849 | v_19908;
assign v_19911 = v_19847 | v_19910;
assign v_19913 = v_19908 | v_19912;
assign v_19915 = v_19846 | v_19914;
assign v_19917 = v_19844 | v_19916;
assign v_19919 = v_19914 | v_19918;
assign v_19921 = v_19843 | v_19920;
assign v_19923 = v_19841 | v_19922;
assign v_19925 = v_19920 | v_19924;
assign v_19927 = v_19840 | v_19926;
assign v_19929 = v_19838 | v_19928;
assign v_19931 = v_19926 | v_19930;
assign v_19933 = v_19837 | v_19932;
assign v_19935 = v_19835 | v_19934;
assign v_19937 = v_19932 | v_19936;
assign v_19939 = v_19834 | v_19938;
assign v_19941 = v_19832 | v_19940;
assign v_19943 = v_19938 | v_19942;
assign v_19945 = v_19831 | v_19944;
assign v_19947 = v_19829 | v_19946;
assign v_19949 = v_19944 | v_19948;
assign v_19951 = v_19828 | v_19950;
assign v_19953 = v_19826 | v_19952;
assign v_19955 = v_19950 | v_19954;
assign v_19957 = v_19825 | v_19956;
assign v_19959 = v_19823 | v_19958;
assign v_19961 = v_19956 | v_19960;
assign v_19963 = v_19822 | v_19962;
assign v_19965 = v_19820 | v_19964;
assign v_19967 = v_19962 | v_19966;
assign v_19970 = ~v_19819 | v_19969;
assign v_19977 = v_19867 | v_19976;
assign v_19980 = v_19978 | v_19979;
assign v_19982 = v_19864 | v_19981;
assign v_19985 = v_19983 | v_19984;
assign v_19987 = v_19861 | v_19986;
assign v_19990 = v_19988 | v_19989;
assign v_19992 = v_19858 | v_19991;
assign v_19995 = v_19993 | v_19994;
assign v_19997 = v_19855 | v_19996;
assign v_20000 = v_19998 | v_19999;
assign v_20002 = v_19852 | v_20001;
assign v_20005 = v_20003 | v_20004;
assign v_20007 = v_19849 | v_20006;
assign v_20010 = v_20008 | v_20009;
assign v_20012 = v_19846 | v_20011;
assign v_20015 = v_20013 | v_20014;
assign v_20017 = v_19843 | v_20016;
assign v_20020 = v_20018 | v_20019;
assign v_20022 = v_19840 | v_20021;
assign v_20025 = v_20023 | v_20024;
assign v_20027 = v_19837 | v_20026;
assign v_20030 = v_20028 | v_20029;
assign v_20032 = v_19834 | v_20031;
assign v_20035 = v_20033 | v_20034;
assign v_20037 = v_19831 | v_20036;
assign v_20040 = v_20038 | v_20039;
assign v_20042 = v_19828 | v_20041;
assign v_20045 = v_20043 | v_20044;
assign v_20047 = v_19825 | v_20046;
assign v_20050 = v_20048 | v_20049;
assign v_20052 = v_19822 | v_20051;
assign v_20055 = v_20053 | v_20054;
assign v_20057 = v_19819 | v_20056;
assign v_20060 = v_19818 | v_20059;
assign v_20114 = v_20111 | v_20113;
assign v_20116 = v_20110 | v_20115;
assign v_20118 = v_20108 | v_20117;
assign v_20120 = v_20115 | v_20119;
assign v_20122 = v_20107 | v_20121;
assign v_20124 = v_20105 | v_20123;
assign v_20126 = v_20121 | v_20125;
assign v_20128 = v_20104 | v_20127;
assign v_20130 = v_20102 | v_20129;
assign v_20132 = v_20127 | v_20131;
assign v_20134 = v_20101 | v_20133;
assign v_20136 = v_20099 | v_20135;
assign v_20138 = v_20133 | v_20137;
assign v_20140 = v_20098 | v_20139;
assign v_20142 = v_20096 | v_20141;
assign v_20144 = v_20139 | v_20143;
assign v_20146 = v_20095 | v_20145;
assign v_20148 = v_20093 | v_20147;
assign v_20150 = v_20145 | v_20149;
assign v_20152 = v_20092 | v_20151;
assign v_20154 = v_20090 | v_20153;
assign v_20156 = v_20151 | v_20155;
assign v_20158 = v_20089 | v_20157;
assign v_20160 = v_20087 | v_20159;
assign v_20162 = v_20157 | v_20161;
assign v_20164 = v_20086 | v_20163;
assign v_20166 = v_20084 | v_20165;
assign v_20168 = v_20163 | v_20167;
assign v_20170 = v_20083 | v_20169;
assign v_20172 = v_20081 | v_20171;
assign v_20174 = v_20169 | v_20173;
assign v_20176 = v_20080 | v_20175;
assign v_20178 = v_20078 | v_20177;
assign v_20180 = v_20175 | v_20179;
assign v_20182 = v_20077 | v_20181;
assign v_20184 = v_20075 | v_20183;
assign v_20186 = v_20181 | v_20185;
assign v_20188 = v_20074 | v_20187;
assign v_20190 = v_20072 | v_20189;
assign v_20192 = v_20187 | v_20191;
assign v_20194 = v_20071 | v_20193;
assign v_20196 = v_20069 | v_20195;
assign v_20198 = v_20193 | v_20197;
assign v_20200 = v_20068 | v_20199;
assign v_20202 = v_20066 | v_20201;
assign v_20204 = v_20199 | v_20203;
assign v_20206 = v_20065 | v_20205;
assign v_20208 = v_20063 | v_20207;
assign v_20210 = v_20205 | v_20209;
assign v_20213 = ~v_20062 | v_20212;
assign v_20220 = v_20110 | v_20219;
assign v_20223 = v_20221 | v_20222;
assign v_20225 = v_20107 | v_20224;
assign v_20228 = v_20226 | v_20227;
assign v_20230 = v_20104 | v_20229;
assign v_20233 = v_20231 | v_20232;
assign v_20235 = v_20101 | v_20234;
assign v_20238 = v_20236 | v_20237;
assign v_20240 = v_20098 | v_20239;
assign v_20243 = v_20241 | v_20242;
assign v_20245 = v_20095 | v_20244;
assign v_20248 = v_20246 | v_20247;
assign v_20250 = v_20092 | v_20249;
assign v_20253 = v_20251 | v_20252;
assign v_20255 = v_20089 | v_20254;
assign v_20258 = v_20256 | v_20257;
assign v_20260 = v_20086 | v_20259;
assign v_20263 = v_20261 | v_20262;
assign v_20265 = v_20083 | v_20264;
assign v_20268 = v_20266 | v_20267;
assign v_20270 = v_20080 | v_20269;
assign v_20273 = v_20271 | v_20272;
assign v_20275 = v_20077 | v_20274;
assign v_20278 = v_20276 | v_20277;
assign v_20280 = v_20074 | v_20279;
assign v_20283 = v_20281 | v_20282;
assign v_20285 = v_20071 | v_20284;
assign v_20288 = v_20286 | v_20287;
assign v_20290 = v_20068 | v_20289;
assign v_20293 = v_20291 | v_20292;
assign v_20295 = v_20065 | v_20294;
assign v_20298 = v_20296 | v_20297;
assign v_20300 = v_20062 | v_20299;
assign v_20303 = v_20061 | v_20302;
assign v_20357 = v_20354 | v_20356;
assign v_20359 = v_20353 | v_20358;
assign v_20361 = v_20351 | v_20360;
assign v_20363 = v_20358 | v_20362;
assign v_20365 = v_20350 | v_20364;
assign v_20367 = v_20348 | v_20366;
assign v_20369 = v_20364 | v_20368;
assign v_20371 = v_20347 | v_20370;
assign v_20373 = v_20345 | v_20372;
assign v_20375 = v_20370 | v_20374;
assign v_20377 = v_20344 | v_20376;
assign v_20379 = v_20342 | v_20378;
assign v_20381 = v_20376 | v_20380;
assign v_20383 = v_20341 | v_20382;
assign v_20385 = v_20339 | v_20384;
assign v_20387 = v_20382 | v_20386;
assign v_20389 = v_20338 | v_20388;
assign v_20391 = v_20336 | v_20390;
assign v_20393 = v_20388 | v_20392;
assign v_20395 = v_20335 | v_20394;
assign v_20397 = v_20333 | v_20396;
assign v_20399 = v_20394 | v_20398;
assign v_20401 = v_20332 | v_20400;
assign v_20403 = v_20330 | v_20402;
assign v_20405 = v_20400 | v_20404;
assign v_20407 = v_20329 | v_20406;
assign v_20409 = v_20327 | v_20408;
assign v_20411 = v_20406 | v_20410;
assign v_20413 = v_20326 | v_20412;
assign v_20415 = v_20324 | v_20414;
assign v_20417 = v_20412 | v_20416;
assign v_20419 = v_20323 | v_20418;
assign v_20421 = v_20321 | v_20420;
assign v_20423 = v_20418 | v_20422;
assign v_20425 = v_20320 | v_20424;
assign v_20427 = v_20318 | v_20426;
assign v_20429 = v_20424 | v_20428;
assign v_20431 = v_20317 | v_20430;
assign v_20433 = v_20315 | v_20432;
assign v_20435 = v_20430 | v_20434;
assign v_20437 = v_20314 | v_20436;
assign v_20439 = v_20312 | v_20438;
assign v_20441 = v_20436 | v_20440;
assign v_20443 = v_20311 | v_20442;
assign v_20445 = v_20309 | v_20444;
assign v_20447 = v_20442 | v_20446;
assign v_20449 = v_20308 | v_20448;
assign v_20451 = v_20306 | v_20450;
assign v_20453 = v_20448 | v_20452;
assign v_20456 = ~v_20305 | v_20455;
assign v_20463 = v_20353 | v_20462;
assign v_20466 = v_20464 | v_20465;
assign v_20468 = v_20350 | v_20467;
assign v_20471 = v_20469 | v_20470;
assign v_20473 = v_20347 | v_20472;
assign v_20476 = v_20474 | v_20475;
assign v_20478 = v_20344 | v_20477;
assign v_20481 = v_20479 | v_20480;
assign v_20483 = v_20341 | v_20482;
assign v_20486 = v_20484 | v_20485;
assign v_20488 = v_20338 | v_20487;
assign v_20491 = v_20489 | v_20490;
assign v_20493 = v_20335 | v_20492;
assign v_20496 = v_20494 | v_20495;
assign v_20498 = v_20332 | v_20497;
assign v_20501 = v_20499 | v_20500;
assign v_20503 = v_20329 | v_20502;
assign v_20506 = v_20504 | v_20505;
assign v_20508 = v_20326 | v_20507;
assign v_20511 = v_20509 | v_20510;
assign v_20513 = v_20323 | v_20512;
assign v_20516 = v_20514 | v_20515;
assign v_20518 = v_20320 | v_20517;
assign v_20521 = v_20519 | v_20520;
assign v_20523 = v_20317 | v_20522;
assign v_20526 = v_20524 | v_20525;
assign v_20528 = v_20314 | v_20527;
assign v_20531 = v_20529 | v_20530;
assign v_20533 = v_20311 | v_20532;
assign v_20536 = v_20534 | v_20535;
assign v_20538 = v_20308 | v_20537;
assign v_20541 = v_20539 | v_20540;
assign v_20543 = v_20305 | v_20542;
assign v_20546 = v_20304 | v_20545;
assign v_20600 = v_20597 | v_20599;
assign v_20602 = v_20596 | v_20601;
assign v_20604 = v_20594 | v_20603;
assign v_20606 = v_20601 | v_20605;
assign v_20608 = v_20593 | v_20607;
assign v_20610 = v_20591 | v_20609;
assign v_20612 = v_20607 | v_20611;
assign v_20614 = v_20590 | v_20613;
assign v_20616 = v_20588 | v_20615;
assign v_20618 = v_20613 | v_20617;
assign v_20620 = v_20587 | v_20619;
assign v_20622 = v_20585 | v_20621;
assign v_20624 = v_20619 | v_20623;
assign v_20626 = v_20584 | v_20625;
assign v_20628 = v_20582 | v_20627;
assign v_20630 = v_20625 | v_20629;
assign v_20632 = v_20581 | v_20631;
assign v_20634 = v_20579 | v_20633;
assign v_20636 = v_20631 | v_20635;
assign v_20638 = v_20578 | v_20637;
assign v_20640 = v_20576 | v_20639;
assign v_20642 = v_20637 | v_20641;
assign v_20644 = v_20575 | v_20643;
assign v_20646 = v_20573 | v_20645;
assign v_20648 = v_20643 | v_20647;
assign v_20650 = v_20572 | v_20649;
assign v_20652 = v_20570 | v_20651;
assign v_20654 = v_20649 | v_20653;
assign v_20656 = v_20569 | v_20655;
assign v_20658 = v_20567 | v_20657;
assign v_20660 = v_20655 | v_20659;
assign v_20662 = v_20566 | v_20661;
assign v_20664 = v_20564 | v_20663;
assign v_20666 = v_20661 | v_20665;
assign v_20668 = v_20563 | v_20667;
assign v_20670 = v_20561 | v_20669;
assign v_20672 = v_20667 | v_20671;
assign v_20674 = v_20560 | v_20673;
assign v_20676 = v_20558 | v_20675;
assign v_20678 = v_20673 | v_20677;
assign v_20680 = v_20557 | v_20679;
assign v_20682 = v_20555 | v_20681;
assign v_20684 = v_20679 | v_20683;
assign v_20686 = v_20554 | v_20685;
assign v_20688 = v_20552 | v_20687;
assign v_20690 = v_20685 | v_20689;
assign v_20692 = v_20551 | v_20691;
assign v_20694 = v_20549 | v_20693;
assign v_20696 = v_20691 | v_20695;
assign v_20699 = ~v_20548 | v_20698;
assign v_20706 = v_20596 | v_20705;
assign v_20709 = v_20707 | v_20708;
assign v_20711 = v_20593 | v_20710;
assign v_20714 = v_20712 | v_20713;
assign v_20716 = v_20590 | v_20715;
assign v_20719 = v_20717 | v_20718;
assign v_20721 = v_20587 | v_20720;
assign v_20724 = v_20722 | v_20723;
assign v_20726 = v_20584 | v_20725;
assign v_20729 = v_20727 | v_20728;
assign v_20731 = v_20581 | v_20730;
assign v_20734 = v_20732 | v_20733;
assign v_20736 = v_20578 | v_20735;
assign v_20739 = v_20737 | v_20738;
assign v_20741 = v_20575 | v_20740;
assign v_20744 = v_20742 | v_20743;
assign v_20746 = v_20572 | v_20745;
assign v_20749 = v_20747 | v_20748;
assign v_20751 = v_20569 | v_20750;
assign v_20754 = v_20752 | v_20753;
assign v_20756 = v_20566 | v_20755;
assign v_20759 = v_20757 | v_20758;
assign v_20761 = v_20563 | v_20760;
assign v_20764 = v_20762 | v_20763;
assign v_20766 = v_20560 | v_20765;
assign v_20769 = v_20767 | v_20768;
assign v_20771 = v_20557 | v_20770;
assign v_20774 = v_20772 | v_20773;
assign v_20776 = v_20554 | v_20775;
assign v_20779 = v_20777 | v_20778;
assign v_20781 = v_20551 | v_20780;
assign v_20784 = v_20782 | v_20783;
assign v_20786 = v_20548 | v_20785;
assign v_20789 = v_20547 | v_20788;
assign v_20842 = v_20839 | v_20841;
assign v_20844 = v_20838 | v_20843;
assign v_20846 = v_20836 | v_20845;
assign v_20848 = v_20843 | v_20847;
assign v_20850 = v_20835 | v_20849;
assign v_20852 = v_20833 | v_20851;
assign v_20854 = v_20849 | v_20853;
assign v_20856 = v_20832 | v_20855;
assign v_20858 = v_20830 | v_20857;
assign v_20860 = v_20855 | v_20859;
assign v_20862 = v_20829 | v_20861;
assign v_20864 = v_20827 | v_20863;
assign v_20866 = v_20861 | v_20865;
assign v_20868 = v_20826 | v_20867;
assign v_20870 = v_20824 | v_20869;
assign v_20872 = v_20867 | v_20871;
assign v_20874 = v_20823 | v_20873;
assign v_20876 = v_20821 | v_20875;
assign v_20878 = v_20873 | v_20877;
assign v_20880 = v_20820 | v_20879;
assign v_20882 = v_20818 | v_20881;
assign v_20884 = v_20879 | v_20883;
assign v_20886 = v_20817 | v_20885;
assign v_20888 = v_20815 | v_20887;
assign v_20890 = v_20885 | v_20889;
assign v_20892 = v_20814 | v_20891;
assign v_20894 = v_20812 | v_20893;
assign v_20896 = v_20891 | v_20895;
assign v_20898 = v_20811 | v_20897;
assign v_20900 = v_20809 | v_20899;
assign v_20902 = v_20897 | v_20901;
assign v_20904 = v_20808 | v_20903;
assign v_20906 = v_20806 | v_20905;
assign v_20908 = v_20903 | v_20907;
assign v_20910 = v_20805 | v_20909;
assign v_20912 = v_20803 | v_20911;
assign v_20914 = v_20909 | v_20913;
assign v_20916 = v_20802 | v_20915;
assign v_20918 = v_20800 | v_20917;
assign v_20920 = v_20915 | v_20919;
assign v_20922 = v_20799 | v_20921;
assign v_20924 = v_20797 | v_20923;
assign v_20926 = v_20921 | v_20925;
assign v_20928 = v_20796 | v_20927;
assign v_20930 = v_20794 | v_20929;
assign v_20932 = v_20927 | v_20931;
assign v_20934 = v_20793 | v_20933;
assign v_20936 = v_20791 | v_20935;
assign v_20938 = v_20933 | v_20937;
assign v_20942 = v_20939 | v_20941;
assign v_20949 = v_20838 | v_20948;
assign v_20952 = v_20950 | v_20951;
assign v_20954 = v_20835 | v_20953;
assign v_20957 = v_20955 | v_20956;
assign v_20959 = v_20832 | v_20958;
assign v_20962 = v_20960 | v_20961;
assign v_20964 = v_20829 | v_20963;
assign v_20967 = v_20965 | v_20966;
assign v_20969 = v_20826 | v_20968;
assign v_20972 = v_20970 | v_20971;
assign v_20974 = v_20823 | v_20973;
assign v_20977 = v_20975 | v_20976;
assign v_20979 = v_20820 | v_20978;
assign v_20982 = v_20980 | v_20981;
assign v_20984 = v_20817 | v_20983;
assign v_20987 = v_20985 | v_20986;
assign v_20989 = v_20814 | v_20988;
assign v_20992 = v_20990 | v_20991;
assign v_20994 = v_20811 | v_20993;
assign v_20997 = v_20995 | v_20996;
assign v_20999 = v_20808 | v_20998;
assign v_21002 = v_21000 | v_21001;
assign v_21004 = v_20805 | v_21003;
assign v_21007 = v_21005 | v_21006;
assign v_21009 = v_20802 | v_21008;
assign v_21012 = v_21010 | v_21011;
assign v_21014 = v_20799 | v_21013;
assign v_21017 = v_21015 | v_21016;
assign v_21019 = v_20796 | v_21018;
assign v_21022 = v_21020 | v_21021;
assign v_21024 = v_20793 | v_21023;
assign v_21027 = v_21025 | v_21026;
assign v_21029 = v_21027 | v_21028;
assign v_21032 = v_20790 | v_21031;
assign v_21103 = v_21100 | v_21102;
assign v_21105 = v_21098 | v_21104;
assign v_21107 = v_21096 | v_21106;
assign v_21109 = v_21104 | v_21108;
assign v_21111 = v_21094 | v_21110;
assign v_21113 = v_21092 | v_21112;
assign v_21115 = v_21110 | v_21114;
assign v_21117 = v_21090 | v_21116;
assign v_21119 = v_21088 | v_21118;
assign v_21121 = v_21116 | v_21120;
assign v_21123 = v_21086 | v_21122;
assign v_21125 = v_21084 | v_21124;
assign v_21127 = v_21122 | v_21126;
assign v_21129 = v_21082 | v_21128;
assign v_21131 = v_21080 | v_21130;
assign v_21133 = v_21128 | v_21132;
assign v_21135 = v_21078 | v_21134;
assign v_21137 = v_21076 | v_21136;
assign v_21139 = v_21134 | v_21138;
assign v_21141 = v_21074 | v_21140;
assign v_21143 = v_21072 | v_21142;
assign v_21145 = v_21140 | v_21144;
assign v_21147 = v_21070 | v_21146;
assign v_21149 = v_21068 | v_21148;
assign v_21151 = v_21146 | v_21150;
assign v_21153 = v_21066 | v_21152;
assign v_21155 = v_21064 | v_21154;
assign v_21157 = v_21152 | v_21156;
assign v_21159 = v_21062 | v_21158;
assign v_21161 = v_21060 | v_21160;
assign v_21163 = v_21158 | v_21162;
assign v_21165 = v_21058 | v_21164;
assign v_21167 = v_21056 | v_21166;
assign v_21169 = v_21164 | v_21168;
assign v_21171 = v_21054 | v_21170;
assign v_21173 = v_21052 | v_21172;
assign v_21175 = v_21170 | v_21174;
assign v_21177 = v_21050 | v_21176;
assign v_21179 = v_21047 | v_21178;
assign v_21181 = v_21176 | v_21180;
assign v_21183 = v_21046 | v_21182;
assign v_21185 = v_21043 | v_21184;
assign v_21187 = v_21182 | v_21186;
assign v_21189 = v_21042 | v_21188;
assign v_21191 = v_21039 | v_21190;
assign v_21193 = v_21188 | v_21192;
assign v_21195 = v_21038 | v_21194;
assign v_21197 = v_21035 | v_21196;
assign v_21199 = v_21194 | v_21198;
assign v_21202 = ~v_21034 | v_21201;
assign v_21209 = v_21098 | v_21208;
assign v_21212 = v_21210 | v_21211;
assign v_21214 = v_21094 | v_21213;
assign v_21217 = v_21215 | v_21216;
assign v_21219 = v_21090 | v_21218;
assign v_21222 = v_21220 | v_21221;
assign v_21224 = v_21086 | v_21223;
assign v_21227 = v_21225 | v_21226;
assign v_21229 = v_21082 | v_21228;
assign v_21232 = v_21230 | v_21231;
assign v_21234 = v_21078 | v_21233;
assign v_21237 = v_21235 | v_21236;
assign v_21239 = v_21074 | v_21238;
assign v_21242 = v_21240 | v_21241;
assign v_21244 = v_21070 | v_21243;
assign v_21247 = v_21245 | v_21246;
assign v_21249 = v_21066 | v_21248;
assign v_21252 = v_21250 | v_21251;
assign v_21254 = v_21062 | v_21253;
assign v_21257 = v_21255 | v_21256;
assign v_21259 = v_21058 | v_21258;
assign v_21262 = v_21260 | v_21261;
assign v_21264 = v_21054 | v_21263;
assign v_21267 = v_21265 | v_21266;
assign v_21269 = v_21050 | v_21268;
assign v_21272 = v_21270 | v_21271;
assign v_21274 = v_21046 | v_21273;
assign v_21277 = v_21275 | v_21276;
assign v_21279 = v_21042 | v_21278;
assign v_21282 = v_21280 | v_21281;
assign v_21284 = v_21038 | v_21283;
assign v_21287 = v_21285 | v_21286;
assign v_21289 = v_21034 | v_21288;
assign v_21292 = v_21033 | v_21291;
assign v_21346 = v_21343 | v_21345;
assign v_21348 = v_21342 | v_21347;
assign v_21350 = v_21340 | v_21349;
assign v_21352 = v_21347 | v_21351;
assign v_21354 = v_21339 | v_21353;
assign v_21356 = v_21337 | v_21355;
assign v_21358 = v_21353 | v_21357;
assign v_21360 = v_21336 | v_21359;
assign v_21362 = v_21334 | v_21361;
assign v_21364 = v_21359 | v_21363;
assign v_21366 = v_21333 | v_21365;
assign v_21368 = v_21331 | v_21367;
assign v_21370 = v_21365 | v_21369;
assign v_21372 = v_21330 | v_21371;
assign v_21374 = v_21328 | v_21373;
assign v_21376 = v_21371 | v_21375;
assign v_21378 = v_21327 | v_21377;
assign v_21380 = v_21325 | v_21379;
assign v_21382 = v_21377 | v_21381;
assign v_21384 = v_21324 | v_21383;
assign v_21386 = v_21322 | v_21385;
assign v_21388 = v_21383 | v_21387;
assign v_21390 = v_21321 | v_21389;
assign v_21392 = v_21319 | v_21391;
assign v_21394 = v_21389 | v_21393;
assign v_21396 = v_21318 | v_21395;
assign v_21398 = v_21316 | v_21397;
assign v_21400 = v_21395 | v_21399;
assign v_21402 = v_21315 | v_21401;
assign v_21404 = v_21313 | v_21403;
assign v_21406 = v_21401 | v_21405;
assign v_21408 = v_21312 | v_21407;
assign v_21410 = v_21310 | v_21409;
assign v_21412 = v_21407 | v_21411;
assign v_21414 = v_21309 | v_21413;
assign v_21416 = v_21307 | v_21415;
assign v_21418 = v_21413 | v_21417;
assign v_21420 = v_21306 | v_21419;
assign v_21422 = v_21304 | v_21421;
assign v_21424 = v_21419 | v_21423;
assign v_21426 = v_21303 | v_21425;
assign v_21428 = v_21301 | v_21427;
assign v_21430 = v_21425 | v_21429;
assign v_21432 = v_21300 | v_21431;
assign v_21434 = v_21298 | v_21433;
assign v_21436 = v_21431 | v_21435;
assign v_21438 = v_21297 | v_21437;
assign v_21440 = v_21295 | v_21439;
assign v_21442 = v_21437 | v_21441;
assign v_21445 = ~v_21294 | v_21444;
assign v_21452 = v_21342 | v_21451;
assign v_21455 = v_21453 | v_21454;
assign v_21457 = v_21339 | v_21456;
assign v_21460 = v_21458 | v_21459;
assign v_21462 = v_21336 | v_21461;
assign v_21465 = v_21463 | v_21464;
assign v_21467 = v_21333 | v_21466;
assign v_21470 = v_21468 | v_21469;
assign v_21472 = v_21330 | v_21471;
assign v_21475 = v_21473 | v_21474;
assign v_21477 = v_21327 | v_21476;
assign v_21480 = v_21478 | v_21479;
assign v_21482 = v_21324 | v_21481;
assign v_21485 = v_21483 | v_21484;
assign v_21487 = v_21321 | v_21486;
assign v_21490 = v_21488 | v_21489;
assign v_21492 = v_21318 | v_21491;
assign v_21495 = v_21493 | v_21494;
assign v_21497 = v_21315 | v_21496;
assign v_21500 = v_21498 | v_21499;
assign v_21502 = v_21312 | v_21501;
assign v_21505 = v_21503 | v_21504;
assign v_21507 = v_21309 | v_21506;
assign v_21510 = v_21508 | v_21509;
assign v_21512 = v_21306 | v_21511;
assign v_21515 = v_21513 | v_21514;
assign v_21517 = v_21303 | v_21516;
assign v_21520 = v_21518 | v_21519;
assign v_21522 = v_21300 | v_21521;
assign v_21525 = v_21523 | v_21524;
assign v_21527 = v_21297 | v_21526;
assign v_21530 = v_21528 | v_21529;
assign v_21532 = v_21294 | v_21531;
assign v_21535 = v_21293 | v_21534;
assign v_21589 = v_21586 | v_21588;
assign v_21591 = v_21585 | v_21590;
assign v_21593 = v_21583 | v_21592;
assign v_21595 = v_21590 | v_21594;
assign v_21597 = v_21582 | v_21596;
assign v_21599 = v_21580 | v_21598;
assign v_21601 = v_21596 | v_21600;
assign v_21603 = v_21579 | v_21602;
assign v_21605 = v_21577 | v_21604;
assign v_21607 = v_21602 | v_21606;
assign v_21609 = v_21576 | v_21608;
assign v_21611 = v_21574 | v_21610;
assign v_21613 = v_21608 | v_21612;
assign v_21615 = v_21573 | v_21614;
assign v_21617 = v_21571 | v_21616;
assign v_21619 = v_21614 | v_21618;
assign v_21621 = v_21570 | v_21620;
assign v_21623 = v_21568 | v_21622;
assign v_21625 = v_21620 | v_21624;
assign v_21627 = v_21567 | v_21626;
assign v_21629 = v_21565 | v_21628;
assign v_21631 = v_21626 | v_21630;
assign v_21633 = v_21564 | v_21632;
assign v_21635 = v_21562 | v_21634;
assign v_21637 = v_21632 | v_21636;
assign v_21639 = v_21561 | v_21638;
assign v_21641 = v_21559 | v_21640;
assign v_21643 = v_21638 | v_21642;
assign v_21645 = v_21558 | v_21644;
assign v_21647 = v_21556 | v_21646;
assign v_21649 = v_21644 | v_21648;
assign v_21651 = v_21555 | v_21650;
assign v_21653 = v_21553 | v_21652;
assign v_21655 = v_21650 | v_21654;
assign v_21657 = v_21552 | v_21656;
assign v_21659 = v_21550 | v_21658;
assign v_21661 = v_21656 | v_21660;
assign v_21663 = v_21549 | v_21662;
assign v_21665 = v_21547 | v_21664;
assign v_21667 = v_21662 | v_21666;
assign v_21669 = v_21546 | v_21668;
assign v_21671 = v_21544 | v_21670;
assign v_21673 = v_21668 | v_21672;
assign v_21675 = v_21543 | v_21674;
assign v_21677 = v_21541 | v_21676;
assign v_21679 = v_21674 | v_21678;
assign v_21681 = v_21540 | v_21680;
assign v_21683 = v_21538 | v_21682;
assign v_21685 = v_21680 | v_21684;
assign v_21688 = ~v_21537 | v_21687;
assign v_21695 = v_21585 | v_21694;
assign v_21698 = v_21696 | v_21697;
assign v_21700 = v_21582 | v_21699;
assign v_21703 = v_21701 | v_21702;
assign v_21705 = v_21579 | v_21704;
assign v_21708 = v_21706 | v_21707;
assign v_21710 = v_21576 | v_21709;
assign v_21713 = v_21711 | v_21712;
assign v_21715 = v_21573 | v_21714;
assign v_21718 = v_21716 | v_21717;
assign v_21720 = v_21570 | v_21719;
assign v_21723 = v_21721 | v_21722;
assign v_21725 = v_21567 | v_21724;
assign v_21728 = v_21726 | v_21727;
assign v_21730 = v_21564 | v_21729;
assign v_21733 = v_21731 | v_21732;
assign v_21735 = v_21561 | v_21734;
assign v_21738 = v_21736 | v_21737;
assign v_21740 = v_21558 | v_21739;
assign v_21743 = v_21741 | v_21742;
assign v_21745 = v_21555 | v_21744;
assign v_21748 = v_21746 | v_21747;
assign v_21750 = v_21552 | v_21749;
assign v_21753 = v_21751 | v_21752;
assign v_21755 = v_21549 | v_21754;
assign v_21758 = v_21756 | v_21757;
assign v_21760 = v_21546 | v_21759;
assign v_21763 = v_21761 | v_21762;
assign v_21765 = v_21543 | v_21764;
assign v_21768 = v_21766 | v_21767;
assign v_21770 = v_21540 | v_21769;
assign v_21773 = v_21771 | v_21772;
assign v_21775 = v_21537 | v_21774;
assign v_21778 = v_21536 | v_21777;
assign v_21832 = v_21829 | v_21831;
assign v_21834 = v_21828 | v_21833;
assign v_21836 = v_21826 | v_21835;
assign v_21838 = v_21833 | v_21837;
assign v_21840 = v_21825 | v_21839;
assign v_21842 = v_21823 | v_21841;
assign v_21844 = v_21839 | v_21843;
assign v_21846 = v_21822 | v_21845;
assign v_21848 = v_21820 | v_21847;
assign v_21850 = v_21845 | v_21849;
assign v_21852 = v_21819 | v_21851;
assign v_21854 = v_21817 | v_21853;
assign v_21856 = v_21851 | v_21855;
assign v_21858 = v_21816 | v_21857;
assign v_21860 = v_21814 | v_21859;
assign v_21862 = v_21857 | v_21861;
assign v_21864 = v_21813 | v_21863;
assign v_21866 = v_21811 | v_21865;
assign v_21868 = v_21863 | v_21867;
assign v_21870 = v_21810 | v_21869;
assign v_21872 = v_21808 | v_21871;
assign v_21874 = v_21869 | v_21873;
assign v_21876 = v_21807 | v_21875;
assign v_21878 = v_21805 | v_21877;
assign v_21880 = v_21875 | v_21879;
assign v_21882 = v_21804 | v_21881;
assign v_21884 = v_21802 | v_21883;
assign v_21886 = v_21881 | v_21885;
assign v_21888 = v_21801 | v_21887;
assign v_21890 = v_21799 | v_21889;
assign v_21892 = v_21887 | v_21891;
assign v_21894 = v_21798 | v_21893;
assign v_21896 = v_21796 | v_21895;
assign v_21898 = v_21893 | v_21897;
assign v_21900 = v_21795 | v_21899;
assign v_21902 = v_21793 | v_21901;
assign v_21904 = v_21899 | v_21903;
assign v_21906 = v_21792 | v_21905;
assign v_21908 = v_21790 | v_21907;
assign v_21910 = v_21905 | v_21909;
assign v_21912 = v_21789 | v_21911;
assign v_21914 = v_21787 | v_21913;
assign v_21916 = v_21911 | v_21915;
assign v_21918 = v_21786 | v_21917;
assign v_21920 = v_21784 | v_21919;
assign v_21922 = v_21917 | v_21921;
assign v_21924 = v_21783 | v_21923;
assign v_21926 = v_21781 | v_21925;
assign v_21928 = v_21923 | v_21927;
assign v_21931 = ~v_21780 | v_21930;
assign v_21938 = v_21828 | v_21937;
assign v_21941 = v_21939 | v_21940;
assign v_21943 = v_21825 | v_21942;
assign v_21946 = v_21944 | v_21945;
assign v_21948 = v_21822 | v_21947;
assign v_21951 = v_21949 | v_21950;
assign v_21953 = v_21819 | v_21952;
assign v_21956 = v_21954 | v_21955;
assign v_21958 = v_21816 | v_21957;
assign v_21961 = v_21959 | v_21960;
assign v_21963 = v_21813 | v_21962;
assign v_21966 = v_21964 | v_21965;
assign v_21968 = v_21810 | v_21967;
assign v_21971 = v_21969 | v_21970;
assign v_21973 = v_21807 | v_21972;
assign v_21976 = v_21974 | v_21975;
assign v_21978 = v_21804 | v_21977;
assign v_21981 = v_21979 | v_21980;
assign v_21983 = v_21801 | v_21982;
assign v_21986 = v_21984 | v_21985;
assign v_21988 = v_21798 | v_21987;
assign v_21991 = v_21989 | v_21990;
assign v_21993 = v_21795 | v_21992;
assign v_21996 = v_21994 | v_21995;
assign v_21998 = v_21792 | v_21997;
assign v_22001 = v_21999 | v_22000;
assign v_22003 = v_21789 | v_22002;
assign v_22006 = v_22004 | v_22005;
assign v_22008 = v_21786 | v_22007;
assign v_22011 = v_22009 | v_22010;
assign v_22013 = v_21783 | v_22012;
assign v_22016 = v_22014 | v_22015;
assign v_22018 = v_21780 | v_22017;
assign v_22021 = v_21779 | v_22020;
assign v_22075 = v_22072 | v_22074;
assign v_22077 = v_22071 | v_22076;
assign v_22079 = v_22069 | v_22078;
assign v_22081 = v_22076 | v_22080;
assign v_22083 = v_22068 | v_22082;
assign v_22085 = v_22066 | v_22084;
assign v_22087 = v_22082 | v_22086;
assign v_22089 = v_22065 | v_22088;
assign v_22091 = v_22063 | v_22090;
assign v_22093 = v_22088 | v_22092;
assign v_22095 = v_22062 | v_22094;
assign v_22097 = v_22060 | v_22096;
assign v_22099 = v_22094 | v_22098;
assign v_22101 = v_22059 | v_22100;
assign v_22103 = v_22057 | v_22102;
assign v_22105 = v_22100 | v_22104;
assign v_22107 = v_22056 | v_22106;
assign v_22109 = v_22054 | v_22108;
assign v_22111 = v_22106 | v_22110;
assign v_22113 = v_22053 | v_22112;
assign v_22115 = v_22051 | v_22114;
assign v_22117 = v_22112 | v_22116;
assign v_22119 = v_22050 | v_22118;
assign v_22121 = v_22048 | v_22120;
assign v_22123 = v_22118 | v_22122;
assign v_22125 = v_22047 | v_22124;
assign v_22127 = v_22045 | v_22126;
assign v_22129 = v_22124 | v_22128;
assign v_22131 = v_22044 | v_22130;
assign v_22133 = v_22042 | v_22132;
assign v_22135 = v_22130 | v_22134;
assign v_22137 = v_22041 | v_22136;
assign v_22139 = v_22039 | v_22138;
assign v_22141 = v_22136 | v_22140;
assign v_22143 = v_22038 | v_22142;
assign v_22145 = v_22036 | v_22144;
assign v_22147 = v_22142 | v_22146;
assign v_22149 = v_22035 | v_22148;
assign v_22151 = v_22033 | v_22150;
assign v_22153 = v_22148 | v_22152;
assign v_22155 = v_22032 | v_22154;
assign v_22157 = v_22030 | v_22156;
assign v_22159 = v_22154 | v_22158;
assign v_22161 = v_22029 | v_22160;
assign v_22163 = v_22027 | v_22162;
assign v_22165 = v_22160 | v_22164;
assign v_22167 = v_22026 | v_22166;
assign v_22169 = v_22024 | v_22168;
assign v_22171 = v_22166 | v_22170;
assign v_22174 = ~v_22023 | v_22173;
assign v_22181 = v_22071 | v_22180;
assign v_22184 = v_22182 | v_22183;
assign v_22186 = v_22068 | v_22185;
assign v_22189 = v_22187 | v_22188;
assign v_22191 = v_22065 | v_22190;
assign v_22194 = v_22192 | v_22193;
assign v_22196 = v_22062 | v_22195;
assign v_22199 = v_22197 | v_22198;
assign v_22201 = v_22059 | v_22200;
assign v_22204 = v_22202 | v_22203;
assign v_22206 = v_22056 | v_22205;
assign v_22209 = v_22207 | v_22208;
assign v_22211 = v_22053 | v_22210;
assign v_22214 = v_22212 | v_22213;
assign v_22216 = v_22050 | v_22215;
assign v_22219 = v_22217 | v_22218;
assign v_22221 = v_22047 | v_22220;
assign v_22224 = v_22222 | v_22223;
assign v_22226 = v_22044 | v_22225;
assign v_22229 = v_22227 | v_22228;
assign v_22231 = v_22041 | v_22230;
assign v_22234 = v_22232 | v_22233;
assign v_22236 = v_22038 | v_22235;
assign v_22239 = v_22237 | v_22238;
assign v_22241 = v_22035 | v_22240;
assign v_22244 = v_22242 | v_22243;
assign v_22246 = v_22032 | v_22245;
assign v_22249 = v_22247 | v_22248;
assign v_22251 = v_22029 | v_22250;
assign v_22254 = v_22252 | v_22253;
assign v_22256 = v_22026 | v_22255;
assign v_22259 = v_22257 | v_22258;
assign v_22261 = v_22023 | v_22260;
assign v_22264 = v_22022 | v_22263;
assign v_22318 = v_22315 | v_22317;
assign v_22320 = v_22314 | v_22319;
assign v_22322 = v_22312 | v_22321;
assign v_22324 = v_22319 | v_22323;
assign v_22326 = v_22311 | v_22325;
assign v_22328 = v_22309 | v_22327;
assign v_22330 = v_22325 | v_22329;
assign v_22332 = v_22308 | v_22331;
assign v_22334 = v_22306 | v_22333;
assign v_22336 = v_22331 | v_22335;
assign v_22338 = v_22305 | v_22337;
assign v_22340 = v_22303 | v_22339;
assign v_22342 = v_22337 | v_22341;
assign v_22344 = v_22302 | v_22343;
assign v_22346 = v_22300 | v_22345;
assign v_22348 = v_22343 | v_22347;
assign v_22350 = v_22299 | v_22349;
assign v_22352 = v_22297 | v_22351;
assign v_22354 = v_22349 | v_22353;
assign v_22356 = v_22296 | v_22355;
assign v_22358 = v_22294 | v_22357;
assign v_22360 = v_22355 | v_22359;
assign v_22362 = v_22293 | v_22361;
assign v_22364 = v_22291 | v_22363;
assign v_22366 = v_22361 | v_22365;
assign v_22368 = v_22290 | v_22367;
assign v_22370 = v_22288 | v_22369;
assign v_22372 = v_22367 | v_22371;
assign v_22374 = v_22287 | v_22373;
assign v_22376 = v_22285 | v_22375;
assign v_22378 = v_22373 | v_22377;
assign v_22380 = v_22284 | v_22379;
assign v_22382 = v_22282 | v_22381;
assign v_22384 = v_22379 | v_22383;
assign v_22386 = v_22281 | v_22385;
assign v_22388 = v_22279 | v_22387;
assign v_22390 = v_22385 | v_22389;
assign v_22392 = v_22278 | v_22391;
assign v_22394 = v_22276 | v_22393;
assign v_22396 = v_22391 | v_22395;
assign v_22398 = v_22275 | v_22397;
assign v_22400 = v_22273 | v_22399;
assign v_22402 = v_22397 | v_22401;
assign v_22404 = v_22272 | v_22403;
assign v_22406 = v_22270 | v_22405;
assign v_22408 = v_22403 | v_22407;
assign v_22410 = v_22269 | v_22409;
assign v_22412 = v_22267 | v_22411;
assign v_22414 = v_22409 | v_22413;
assign v_22417 = ~v_22266 | v_22416;
assign v_22424 = v_22314 | v_22423;
assign v_22427 = v_22425 | v_22426;
assign v_22429 = v_22311 | v_22428;
assign v_22432 = v_22430 | v_22431;
assign v_22434 = v_22308 | v_22433;
assign v_22437 = v_22435 | v_22436;
assign v_22439 = v_22305 | v_22438;
assign v_22442 = v_22440 | v_22441;
assign v_22444 = v_22302 | v_22443;
assign v_22447 = v_22445 | v_22446;
assign v_22449 = v_22299 | v_22448;
assign v_22452 = v_22450 | v_22451;
assign v_22454 = v_22296 | v_22453;
assign v_22457 = v_22455 | v_22456;
assign v_22459 = v_22293 | v_22458;
assign v_22462 = v_22460 | v_22461;
assign v_22464 = v_22290 | v_22463;
assign v_22467 = v_22465 | v_22466;
assign v_22469 = v_22287 | v_22468;
assign v_22472 = v_22470 | v_22471;
assign v_22474 = v_22284 | v_22473;
assign v_22477 = v_22475 | v_22476;
assign v_22479 = v_22281 | v_22478;
assign v_22482 = v_22480 | v_22481;
assign v_22484 = v_22278 | v_22483;
assign v_22487 = v_22485 | v_22486;
assign v_22489 = v_22275 | v_22488;
assign v_22492 = v_22490 | v_22491;
assign v_22494 = v_22272 | v_22493;
assign v_22497 = v_22495 | v_22496;
assign v_22499 = v_22269 | v_22498;
assign v_22502 = v_22500 | v_22501;
assign v_22504 = v_22266 | v_22503;
assign v_22507 = v_22265 | v_22506;
assign v_22561 = v_22558 | v_22560;
assign v_22563 = v_22557 | v_22562;
assign v_22565 = v_22555 | v_22564;
assign v_22567 = v_22562 | v_22566;
assign v_22569 = v_22554 | v_22568;
assign v_22571 = v_22552 | v_22570;
assign v_22573 = v_22568 | v_22572;
assign v_22575 = v_22551 | v_22574;
assign v_22577 = v_22549 | v_22576;
assign v_22579 = v_22574 | v_22578;
assign v_22581 = v_22548 | v_22580;
assign v_22583 = v_22546 | v_22582;
assign v_22585 = v_22580 | v_22584;
assign v_22587 = v_22545 | v_22586;
assign v_22589 = v_22543 | v_22588;
assign v_22591 = v_22586 | v_22590;
assign v_22593 = v_22542 | v_22592;
assign v_22595 = v_22540 | v_22594;
assign v_22597 = v_22592 | v_22596;
assign v_22599 = v_22539 | v_22598;
assign v_22601 = v_22537 | v_22600;
assign v_22603 = v_22598 | v_22602;
assign v_22605 = v_22536 | v_22604;
assign v_22607 = v_22534 | v_22606;
assign v_22609 = v_22604 | v_22608;
assign v_22611 = v_22533 | v_22610;
assign v_22613 = v_22531 | v_22612;
assign v_22615 = v_22610 | v_22614;
assign v_22617 = v_22530 | v_22616;
assign v_22619 = v_22528 | v_22618;
assign v_22621 = v_22616 | v_22620;
assign v_22623 = v_22527 | v_22622;
assign v_22625 = v_22525 | v_22624;
assign v_22627 = v_22622 | v_22626;
assign v_22629 = v_22524 | v_22628;
assign v_22631 = v_22522 | v_22630;
assign v_22633 = v_22628 | v_22632;
assign v_22635 = v_22521 | v_22634;
assign v_22637 = v_22519 | v_22636;
assign v_22639 = v_22634 | v_22638;
assign v_22641 = v_22518 | v_22640;
assign v_22643 = v_22516 | v_22642;
assign v_22645 = v_22640 | v_22644;
assign v_22647 = v_22515 | v_22646;
assign v_22649 = v_22513 | v_22648;
assign v_22651 = v_22646 | v_22650;
assign v_22653 = v_22512 | v_22652;
assign v_22655 = v_22510 | v_22654;
assign v_22657 = v_22652 | v_22656;
assign v_22660 = ~v_22509 | v_22659;
assign v_22667 = v_22557 | v_22666;
assign v_22670 = v_22668 | v_22669;
assign v_22672 = v_22554 | v_22671;
assign v_22675 = v_22673 | v_22674;
assign v_22677 = v_22551 | v_22676;
assign v_22680 = v_22678 | v_22679;
assign v_22682 = v_22548 | v_22681;
assign v_22685 = v_22683 | v_22684;
assign v_22687 = v_22545 | v_22686;
assign v_22690 = v_22688 | v_22689;
assign v_22692 = v_22542 | v_22691;
assign v_22695 = v_22693 | v_22694;
assign v_22697 = v_22539 | v_22696;
assign v_22700 = v_22698 | v_22699;
assign v_22702 = v_22536 | v_22701;
assign v_22705 = v_22703 | v_22704;
assign v_22707 = v_22533 | v_22706;
assign v_22710 = v_22708 | v_22709;
assign v_22712 = v_22530 | v_22711;
assign v_22715 = v_22713 | v_22714;
assign v_22717 = v_22527 | v_22716;
assign v_22720 = v_22718 | v_22719;
assign v_22722 = v_22524 | v_22721;
assign v_22725 = v_22723 | v_22724;
assign v_22727 = v_22521 | v_22726;
assign v_22730 = v_22728 | v_22729;
assign v_22732 = v_22518 | v_22731;
assign v_22735 = v_22733 | v_22734;
assign v_22737 = v_22515 | v_22736;
assign v_22740 = v_22738 | v_22739;
assign v_22742 = v_22512 | v_22741;
assign v_22745 = v_22743 | v_22744;
assign v_22747 = v_22509 | v_22746;
assign v_22750 = v_22508 | v_22749;
assign v_22804 = v_22801 | v_22803;
assign v_22806 = v_22800 | v_22805;
assign v_22808 = v_22798 | v_22807;
assign v_22810 = v_22805 | v_22809;
assign v_22812 = v_22797 | v_22811;
assign v_22814 = v_22795 | v_22813;
assign v_22816 = v_22811 | v_22815;
assign v_22818 = v_22794 | v_22817;
assign v_22820 = v_22792 | v_22819;
assign v_22822 = v_22817 | v_22821;
assign v_22824 = v_22791 | v_22823;
assign v_22826 = v_22789 | v_22825;
assign v_22828 = v_22823 | v_22827;
assign v_22830 = v_22788 | v_22829;
assign v_22832 = v_22786 | v_22831;
assign v_22834 = v_22829 | v_22833;
assign v_22836 = v_22785 | v_22835;
assign v_22838 = v_22783 | v_22837;
assign v_22840 = v_22835 | v_22839;
assign v_22842 = v_22782 | v_22841;
assign v_22844 = v_22780 | v_22843;
assign v_22846 = v_22841 | v_22845;
assign v_22848 = v_22779 | v_22847;
assign v_22850 = v_22777 | v_22849;
assign v_22852 = v_22847 | v_22851;
assign v_22854 = v_22776 | v_22853;
assign v_22856 = v_22774 | v_22855;
assign v_22858 = v_22853 | v_22857;
assign v_22860 = v_22773 | v_22859;
assign v_22862 = v_22771 | v_22861;
assign v_22864 = v_22859 | v_22863;
assign v_22866 = v_22770 | v_22865;
assign v_22868 = v_22768 | v_22867;
assign v_22870 = v_22865 | v_22869;
assign v_22872 = v_22767 | v_22871;
assign v_22874 = v_22765 | v_22873;
assign v_22876 = v_22871 | v_22875;
assign v_22878 = v_22764 | v_22877;
assign v_22880 = v_22762 | v_22879;
assign v_22882 = v_22877 | v_22881;
assign v_22884 = v_22761 | v_22883;
assign v_22886 = v_22759 | v_22885;
assign v_22888 = v_22883 | v_22887;
assign v_22890 = v_22758 | v_22889;
assign v_22892 = v_22756 | v_22891;
assign v_22894 = v_22889 | v_22893;
assign v_22896 = v_22755 | v_22895;
assign v_22898 = v_22753 | v_22897;
assign v_22900 = v_22895 | v_22899;
assign v_22903 = ~v_22752 | v_22902;
assign v_22910 = v_22800 | v_22909;
assign v_22913 = v_22911 | v_22912;
assign v_22915 = v_22797 | v_22914;
assign v_22918 = v_22916 | v_22917;
assign v_22920 = v_22794 | v_22919;
assign v_22923 = v_22921 | v_22922;
assign v_22925 = v_22791 | v_22924;
assign v_22928 = v_22926 | v_22927;
assign v_22930 = v_22788 | v_22929;
assign v_22933 = v_22931 | v_22932;
assign v_22935 = v_22785 | v_22934;
assign v_22938 = v_22936 | v_22937;
assign v_22940 = v_22782 | v_22939;
assign v_22943 = v_22941 | v_22942;
assign v_22945 = v_22779 | v_22944;
assign v_22948 = v_22946 | v_22947;
assign v_22950 = v_22776 | v_22949;
assign v_22953 = v_22951 | v_22952;
assign v_22955 = v_22773 | v_22954;
assign v_22958 = v_22956 | v_22957;
assign v_22960 = v_22770 | v_22959;
assign v_22963 = v_22961 | v_22962;
assign v_22965 = v_22767 | v_22964;
assign v_22968 = v_22966 | v_22967;
assign v_22970 = v_22764 | v_22969;
assign v_22973 = v_22971 | v_22972;
assign v_22975 = v_22761 | v_22974;
assign v_22978 = v_22976 | v_22977;
assign v_22980 = v_22758 | v_22979;
assign v_22983 = v_22981 | v_22982;
assign v_22985 = v_22755 | v_22984;
assign v_22988 = v_22986 | v_22987;
assign v_22990 = v_22752 | v_22989;
assign v_22993 = v_22751 | v_22992;
assign v_23047 = v_23044 | v_23046;
assign v_23049 = v_23043 | v_23048;
assign v_23051 = v_23041 | v_23050;
assign v_23053 = v_23048 | v_23052;
assign v_23055 = v_23040 | v_23054;
assign v_23057 = v_23038 | v_23056;
assign v_23059 = v_23054 | v_23058;
assign v_23061 = v_23037 | v_23060;
assign v_23063 = v_23035 | v_23062;
assign v_23065 = v_23060 | v_23064;
assign v_23067 = v_23034 | v_23066;
assign v_23069 = v_23032 | v_23068;
assign v_23071 = v_23066 | v_23070;
assign v_23073 = v_23031 | v_23072;
assign v_23075 = v_23029 | v_23074;
assign v_23077 = v_23072 | v_23076;
assign v_23079 = v_23028 | v_23078;
assign v_23081 = v_23026 | v_23080;
assign v_23083 = v_23078 | v_23082;
assign v_23085 = v_23025 | v_23084;
assign v_23087 = v_23023 | v_23086;
assign v_23089 = v_23084 | v_23088;
assign v_23091 = v_23022 | v_23090;
assign v_23093 = v_23020 | v_23092;
assign v_23095 = v_23090 | v_23094;
assign v_23097 = v_23019 | v_23096;
assign v_23099 = v_23017 | v_23098;
assign v_23101 = v_23096 | v_23100;
assign v_23103 = v_23016 | v_23102;
assign v_23105 = v_23014 | v_23104;
assign v_23107 = v_23102 | v_23106;
assign v_23109 = v_23013 | v_23108;
assign v_23111 = v_23011 | v_23110;
assign v_23113 = v_23108 | v_23112;
assign v_23115 = v_23010 | v_23114;
assign v_23117 = v_23008 | v_23116;
assign v_23119 = v_23114 | v_23118;
assign v_23121 = v_23007 | v_23120;
assign v_23123 = v_23005 | v_23122;
assign v_23125 = v_23120 | v_23124;
assign v_23127 = v_23004 | v_23126;
assign v_23129 = v_23002 | v_23128;
assign v_23131 = v_23126 | v_23130;
assign v_23133 = v_23001 | v_23132;
assign v_23135 = v_22999 | v_23134;
assign v_23137 = v_23132 | v_23136;
assign v_23139 = v_22998 | v_23138;
assign v_23141 = v_22996 | v_23140;
assign v_23143 = v_23138 | v_23142;
assign v_23146 = ~v_22995 | v_23145;
assign v_23153 = v_23043 | v_23152;
assign v_23156 = v_23154 | v_23155;
assign v_23158 = v_23040 | v_23157;
assign v_23161 = v_23159 | v_23160;
assign v_23163 = v_23037 | v_23162;
assign v_23166 = v_23164 | v_23165;
assign v_23168 = v_23034 | v_23167;
assign v_23171 = v_23169 | v_23170;
assign v_23173 = v_23031 | v_23172;
assign v_23176 = v_23174 | v_23175;
assign v_23178 = v_23028 | v_23177;
assign v_23181 = v_23179 | v_23180;
assign v_23183 = v_23025 | v_23182;
assign v_23186 = v_23184 | v_23185;
assign v_23188 = v_23022 | v_23187;
assign v_23191 = v_23189 | v_23190;
assign v_23193 = v_23019 | v_23192;
assign v_23196 = v_23194 | v_23195;
assign v_23198 = v_23016 | v_23197;
assign v_23201 = v_23199 | v_23200;
assign v_23203 = v_23013 | v_23202;
assign v_23206 = v_23204 | v_23205;
assign v_23208 = v_23010 | v_23207;
assign v_23211 = v_23209 | v_23210;
assign v_23213 = v_23007 | v_23212;
assign v_23216 = v_23214 | v_23215;
assign v_23218 = v_23004 | v_23217;
assign v_23221 = v_23219 | v_23220;
assign v_23223 = v_23001 | v_23222;
assign v_23226 = v_23224 | v_23225;
assign v_23228 = v_22998 | v_23227;
assign v_23231 = v_23229 | v_23230;
assign v_23233 = v_22995 | v_23232;
assign v_23236 = v_22994 | v_23235;
assign v_23290 = v_23287 | v_23289;
assign v_23292 = v_23286 | v_23291;
assign v_23294 = v_23284 | v_23293;
assign v_23296 = v_23291 | v_23295;
assign v_23298 = v_23283 | v_23297;
assign v_23300 = v_23281 | v_23299;
assign v_23302 = v_23297 | v_23301;
assign v_23304 = v_23280 | v_23303;
assign v_23306 = v_23278 | v_23305;
assign v_23308 = v_23303 | v_23307;
assign v_23310 = v_23277 | v_23309;
assign v_23312 = v_23275 | v_23311;
assign v_23314 = v_23309 | v_23313;
assign v_23316 = v_23274 | v_23315;
assign v_23318 = v_23272 | v_23317;
assign v_23320 = v_23315 | v_23319;
assign v_23322 = v_23271 | v_23321;
assign v_23324 = v_23269 | v_23323;
assign v_23326 = v_23321 | v_23325;
assign v_23328 = v_23268 | v_23327;
assign v_23330 = v_23266 | v_23329;
assign v_23332 = v_23327 | v_23331;
assign v_23334 = v_23265 | v_23333;
assign v_23336 = v_23263 | v_23335;
assign v_23338 = v_23333 | v_23337;
assign v_23340 = v_23262 | v_23339;
assign v_23342 = v_23260 | v_23341;
assign v_23344 = v_23339 | v_23343;
assign v_23346 = v_23259 | v_23345;
assign v_23348 = v_23257 | v_23347;
assign v_23350 = v_23345 | v_23349;
assign v_23352 = v_23256 | v_23351;
assign v_23354 = v_23254 | v_23353;
assign v_23356 = v_23351 | v_23355;
assign v_23358 = v_23253 | v_23357;
assign v_23360 = v_23251 | v_23359;
assign v_23362 = v_23357 | v_23361;
assign v_23364 = v_23250 | v_23363;
assign v_23366 = v_23248 | v_23365;
assign v_23368 = v_23363 | v_23367;
assign v_23370 = v_23247 | v_23369;
assign v_23372 = v_23245 | v_23371;
assign v_23374 = v_23369 | v_23373;
assign v_23376 = v_23244 | v_23375;
assign v_23378 = v_23242 | v_23377;
assign v_23380 = v_23375 | v_23379;
assign v_23382 = v_23241 | v_23381;
assign v_23384 = v_23239 | v_23383;
assign v_23386 = v_23381 | v_23385;
assign v_23389 = ~v_23238 | v_23388;
assign v_23396 = v_23286 | v_23395;
assign v_23399 = v_23397 | v_23398;
assign v_23401 = v_23283 | v_23400;
assign v_23404 = v_23402 | v_23403;
assign v_23406 = v_23280 | v_23405;
assign v_23409 = v_23407 | v_23408;
assign v_23411 = v_23277 | v_23410;
assign v_23414 = v_23412 | v_23413;
assign v_23416 = v_23274 | v_23415;
assign v_23419 = v_23417 | v_23418;
assign v_23421 = v_23271 | v_23420;
assign v_23424 = v_23422 | v_23423;
assign v_23426 = v_23268 | v_23425;
assign v_23429 = v_23427 | v_23428;
assign v_23431 = v_23265 | v_23430;
assign v_23434 = v_23432 | v_23433;
assign v_23436 = v_23262 | v_23435;
assign v_23439 = v_23437 | v_23438;
assign v_23441 = v_23259 | v_23440;
assign v_23444 = v_23442 | v_23443;
assign v_23446 = v_23256 | v_23445;
assign v_23449 = v_23447 | v_23448;
assign v_23451 = v_23253 | v_23450;
assign v_23454 = v_23452 | v_23453;
assign v_23456 = v_23250 | v_23455;
assign v_23459 = v_23457 | v_23458;
assign v_23461 = v_23247 | v_23460;
assign v_23464 = v_23462 | v_23463;
assign v_23466 = v_23244 | v_23465;
assign v_23469 = v_23467 | v_23468;
assign v_23471 = v_23241 | v_23470;
assign v_23474 = v_23472 | v_23473;
assign v_23476 = v_23238 | v_23475;
assign v_23479 = v_23237 | v_23478;
assign v_23533 = v_23530 | v_23532;
assign v_23535 = v_23529 | v_23534;
assign v_23537 = v_23527 | v_23536;
assign v_23539 = v_23534 | v_23538;
assign v_23541 = v_23526 | v_23540;
assign v_23543 = v_23524 | v_23542;
assign v_23545 = v_23540 | v_23544;
assign v_23547 = v_23523 | v_23546;
assign v_23549 = v_23521 | v_23548;
assign v_23551 = v_23546 | v_23550;
assign v_23553 = v_23520 | v_23552;
assign v_23555 = v_23518 | v_23554;
assign v_23557 = v_23552 | v_23556;
assign v_23559 = v_23517 | v_23558;
assign v_23561 = v_23515 | v_23560;
assign v_23563 = v_23558 | v_23562;
assign v_23565 = v_23514 | v_23564;
assign v_23567 = v_23512 | v_23566;
assign v_23569 = v_23564 | v_23568;
assign v_23571 = v_23511 | v_23570;
assign v_23573 = v_23509 | v_23572;
assign v_23575 = v_23570 | v_23574;
assign v_23577 = v_23508 | v_23576;
assign v_23579 = v_23506 | v_23578;
assign v_23581 = v_23576 | v_23580;
assign v_23583 = v_23505 | v_23582;
assign v_23585 = v_23503 | v_23584;
assign v_23587 = v_23582 | v_23586;
assign v_23589 = v_23502 | v_23588;
assign v_23591 = v_23500 | v_23590;
assign v_23593 = v_23588 | v_23592;
assign v_23595 = v_23499 | v_23594;
assign v_23597 = v_23497 | v_23596;
assign v_23599 = v_23594 | v_23598;
assign v_23601 = v_23496 | v_23600;
assign v_23603 = v_23494 | v_23602;
assign v_23605 = v_23600 | v_23604;
assign v_23607 = v_23493 | v_23606;
assign v_23609 = v_23491 | v_23608;
assign v_23611 = v_23606 | v_23610;
assign v_23613 = v_23490 | v_23612;
assign v_23615 = v_23488 | v_23614;
assign v_23617 = v_23612 | v_23616;
assign v_23619 = v_23487 | v_23618;
assign v_23621 = v_23485 | v_23620;
assign v_23623 = v_23618 | v_23622;
assign v_23625 = v_23484 | v_23624;
assign v_23627 = v_23482 | v_23626;
assign v_23629 = v_23624 | v_23628;
assign v_23632 = ~v_23481 | v_23631;
assign v_23639 = v_23529 | v_23638;
assign v_23642 = v_23640 | v_23641;
assign v_23644 = v_23526 | v_23643;
assign v_23647 = v_23645 | v_23646;
assign v_23649 = v_23523 | v_23648;
assign v_23652 = v_23650 | v_23651;
assign v_23654 = v_23520 | v_23653;
assign v_23657 = v_23655 | v_23656;
assign v_23659 = v_23517 | v_23658;
assign v_23662 = v_23660 | v_23661;
assign v_23664 = v_23514 | v_23663;
assign v_23667 = v_23665 | v_23666;
assign v_23669 = v_23511 | v_23668;
assign v_23672 = v_23670 | v_23671;
assign v_23674 = v_23508 | v_23673;
assign v_23677 = v_23675 | v_23676;
assign v_23679 = v_23505 | v_23678;
assign v_23682 = v_23680 | v_23681;
assign v_23684 = v_23502 | v_23683;
assign v_23687 = v_23685 | v_23686;
assign v_23689 = v_23499 | v_23688;
assign v_23692 = v_23690 | v_23691;
assign v_23694 = v_23496 | v_23693;
assign v_23697 = v_23695 | v_23696;
assign v_23699 = v_23493 | v_23698;
assign v_23702 = v_23700 | v_23701;
assign v_23704 = v_23490 | v_23703;
assign v_23707 = v_23705 | v_23706;
assign v_23709 = v_23487 | v_23708;
assign v_23712 = v_23710 | v_23711;
assign v_23714 = v_23484 | v_23713;
assign v_23717 = v_23715 | v_23716;
assign v_23719 = v_23481 | v_23718;
assign v_23722 = v_23480 | v_23721;
assign v_23776 = v_23773 | v_23775;
assign v_23778 = v_23772 | v_23777;
assign v_23780 = v_23770 | v_23779;
assign v_23782 = v_23777 | v_23781;
assign v_23784 = v_23769 | v_23783;
assign v_23786 = v_23767 | v_23785;
assign v_23788 = v_23783 | v_23787;
assign v_23790 = v_23766 | v_23789;
assign v_23792 = v_23764 | v_23791;
assign v_23794 = v_23789 | v_23793;
assign v_23796 = v_23763 | v_23795;
assign v_23798 = v_23761 | v_23797;
assign v_23800 = v_23795 | v_23799;
assign v_23802 = v_23760 | v_23801;
assign v_23804 = v_23758 | v_23803;
assign v_23806 = v_23801 | v_23805;
assign v_23808 = v_23757 | v_23807;
assign v_23810 = v_23755 | v_23809;
assign v_23812 = v_23807 | v_23811;
assign v_23814 = v_23754 | v_23813;
assign v_23816 = v_23752 | v_23815;
assign v_23818 = v_23813 | v_23817;
assign v_23820 = v_23751 | v_23819;
assign v_23822 = v_23749 | v_23821;
assign v_23824 = v_23819 | v_23823;
assign v_23826 = v_23748 | v_23825;
assign v_23828 = v_23746 | v_23827;
assign v_23830 = v_23825 | v_23829;
assign v_23832 = v_23745 | v_23831;
assign v_23834 = v_23743 | v_23833;
assign v_23836 = v_23831 | v_23835;
assign v_23838 = v_23742 | v_23837;
assign v_23840 = v_23740 | v_23839;
assign v_23842 = v_23837 | v_23841;
assign v_23844 = v_23739 | v_23843;
assign v_23846 = v_23737 | v_23845;
assign v_23848 = v_23843 | v_23847;
assign v_23850 = v_23736 | v_23849;
assign v_23852 = v_23734 | v_23851;
assign v_23854 = v_23849 | v_23853;
assign v_23856 = v_23733 | v_23855;
assign v_23858 = v_23731 | v_23857;
assign v_23860 = v_23855 | v_23859;
assign v_23862 = v_23730 | v_23861;
assign v_23864 = v_23728 | v_23863;
assign v_23866 = v_23861 | v_23865;
assign v_23868 = v_23727 | v_23867;
assign v_23870 = v_23725 | v_23869;
assign v_23872 = v_23867 | v_23871;
assign v_23875 = ~v_23724 | v_23874;
assign v_23882 = v_23772 | v_23881;
assign v_23885 = v_23883 | v_23884;
assign v_23887 = v_23769 | v_23886;
assign v_23890 = v_23888 | v_23889;
assign v_23892 = v_23766 | v_23891;
assign v_23895 = v_23893 | v_23894;
assign v_23897 = v_23763 | v_23896;
assign v_23900 = v_23898 | v_23899;
assign v_23902 = v_23760 | v_23901;
assign v_23905 = v_23903 | v_23904;
assign v_23907 = v_23757 | v_23906;
assign v_23910 = v_23908 | v_23909;
assign v_23912 = v_23754 | v_23911;
assign v_23915 = v_23913 | v_23914;
assign v_23917 = v_23751 | v_23916;
assign v_23920 = v_23918 | v_23919;
assign v_23922 = v_23748 | v_23921;
assign v_23925 = v_23923 | v_23924;
assign v_23927 = v_23745 | v_23926;
assign v_23930 = v_23928 | v_23929;
assign v_23932 = v_23742 | v_23931;
assign v_23935 = v_23933 | v_23934;
assign v_23937 = v_23739 | v_23936;
assign v_23940 = v_23938 | v_23939;
assign v_23942 = v_23736 | v_23941;
assign v_23945 = v_23943 | v_23944;
assign v_23947 = v_23733 | v_23946;
assign v_23950 = v_23948 | v_23949;
assign v_23952 = v_23730 | v_23951;
assign v_23955 = v_23953 | v_23954;
assign v_23957 = v_23727 | v_23956;
assign v_23960 = v_23958 | v_23959;
assign v_23962 = v_23724 | v_23961;
assign v_23965 = v_23723 | v_23964;
assign v_24019 = v_24016 | v_24018;
assign v_24021 = v_24015 | v_24020;
assign v_24023 = v_24013 | v_24022;
assign v_24025 = v_24020 | v_24024;
assign v_24027 = v_24012 | v_24026;
assign v_24029 = v_24010 | v_24028;
assign v_24031 = v_24026 | v_24030;
assign v_24033 = v_24009 | v_24032;
assign v_24035 = v_24007 | v_24034;
assign v_24037 = v_24032 | v_24036;
assign v_24039 = v_24006 | v_24038;
assign v_24041 = v_24004 | v_24040;
assign v_24043 = v_24038 | v_24042;
assign v_24045 = v_24003 | v_24044;
assign v_24047 = v_24001 | v_24046;
assign v_24049 = v_24044 | v_24048;
assign v_24051 = v_24000 | v_24050;
assign v_24053 = v_23998 | v_24052;
assign v_24055 = v_24050 | v_24054;
assign v_24057 = v_23997 | v_24056;
assign v_24059 = v_23995 | v_24058;
assign v_24061 = v_24056 | v_24060;
assign v_24063 = v_23994 | v_24062;
assign v_24065 = v_23992 | v_24064;
assign v_24067 = v_24062 | v_24066;
assign v_24069 = v_23991 | v_24068;
assign v_24071 = v_23989 | v_24070;
assign v_24073 = v_24068 | v_24072;
assign v_24075 = v_23988 | v_24074;
assign v_24077 = v_23986 | v_24076;
assign v_24079 = v_24074 | v_24078;
assign v_24081 = v_23985 | v_24080;
assign v_24083 = v_23983 | v_24082;
assign v_24085 = v_24080 | v_24084;
assign v_24087 = v_23982 | v_24086;
assign v_24089 = v_23980 | v_24088;
assign v_24091 = v_24086 | v_24090;
assign v_24093 = v_23979 | v_24092;
assign v_24095 = v_23977 | v_24094;
assign v_24097 = v_24092 | v_24096;
assign v_24099 = v_23976 | v_24098;
assign v_24101 = v_23974 | v_24100;
assign v_24103 = v_24098 | v_24102;
assign v_24105 = v_23973 | v_24104;
assign v_24107 = v_23971 | v_24106;
assign v_24109 = v_24104 | v_24108;
assign v_24111 = v_23970 | v_24110;
assign v_24113 = v_23968 | v_24112;
assign v_24115 = v_24110 | v_24114;
assign v_24118 = ~v_23967 | v_24117;
assign v_24125 = v_24015 | v_24124;
assign v_24128 = v_24126 | v_24127;
assign v_24130 = v_24012 | v_24129;
assign v_24133 = v_24131 | v_24132;
assign v_24135 = v_24009 | v_24134;
assign v_24138 = v_24136 | v_24137;
assign v_24140 = v_24006 | v_24139;
assign v_24143 = v_24141 | v_24142;
assign v_24145 = v_24003 | v_24144;
assign v_24148 = v_24146 | v_24147;
assign v_24150 = v_24000 | v_24149;
assign v_24153 = v_24151 | v_24152;
assign v_24155 = v_23997 | v_24154;
assign v_24158 = v_24156 | v_24157;
assign v_24160 = v_23994 | v_24159;
assign v_24163 = v_24161 | v_24162;
assign v_24165 = v_23991 | v_24164;
assign v_24168 = v_24166 | v_24167;
assign v_24170 = v_23988 | v_24169;
assign v_24173 = v_24171 | v_24172;
assign v_24175 = v_23985 | v_24174;
assign v_24178 = v_24176 | v_24177;
assign v_24180 = v_23982 | v_24179;
assign v_24183 = v_24181 | v_24182;
assign v_24185 = v_23979 | v_24184;
assign v_24188 = v_24186 | v_24187;
assign v_24190 = v_23976 | v_24189;
assign v_24193 = v_24191 | v_24192;
assign v_24195 = v_23973 | v_24194;
assign v_24198 = v_24196 | v_24197;
assign v_24200 = v_23970 | v_24199;
assign v_24203 = v_24201 | v_24202;
assign v_24205 = v_23967 | v_24204;
assign v_24208 = v_23966 | v_24207;
assign v_24262 = v_24259 | v_24261;
assign v_24264 = v_24258 | v_24263;
assign v_24266 = v_24256 | v_24265;
assign v_24268 = v_24263 | v_24267;
assign v_24270 = v_24255 | v_24269;
assign v_24272 = v_24253 | v_24271;
assign v_24274 = v_24269 | v_24273;
assign v_24276 = v_24252 | v_24275;
assign v_24278 = v_24250 | v_24277;
assign v_24280 = v_24275 | v_24279;
assign v_24282 = v_24249 | v_24281;
assign v_24284 = v_24247 | v_24283;
assign v_24286 = v_24281 | v_24285;
assign v_24288 = v_24246 | v_24287;
assign v_24290 = v_24244 | v_24289;
assign v_24292 = v_24287 | v_24291;
assign v_24294 = v_24243 | v_24293;
assign v_24296 = v_24241 | v_24295;
assign v_24298 = v_24293 | v_24297;
assign v_24300 = v_24240 | v_24299;
assign v_24302 = v_24238 | v_24301;
assign v_24304 = v_24299 | v_24303;
assign v_24306 = v_24237 | v_24305;
assign v_24308 = v_24235 | v_24307;
assign v_24310 = v_24305 | v_24309;
assign v_24312 = v_24234 | v_24311;
assign v_24314 = v_24232 | v_24313;
assign v_24316 = v_24311 | v_24315;
assign v_24318 = v_24231 | v_24317;
assign v_24320 = v_24229 | v_24319;
assign v_24322 = v_24317 | v_24321;
assign v_24324 = v_24228 | v_24323;
assign v_24326 = v_24226 | v_24325;
assign v_24328 = v_24323 | v_24327;
assign v_24330 = v_24225 | v_24329;
assign v_24332 = v_24223 | v_24331;
assign v_24334 = v_24329 | v_24333;
assign v_24336 = v_24222 | v_24335;
assign v_24338 = v_24220 | v_24337;
assign v_24340 = v_24335 | v_24339;
assign v_24342 = v_24219 | v_24341;
assign v_24344 = v_24217 | v_24343;
assign v_24346 = v_24341 | v_24345;
assign v_24348 = v_24216 | v_24347;
assign v_24350 = v_24214 | v_24349;
assign v_24352 = v_24347 | v_24351;
assign v_24354 = v_24213 | v_24353;
assign v_24356 = v_24211 | v_24355;
assign v_24358 = v_24353 | v_24357;
assign v_24361 = ~v_24210 | v_24360;
assign v_24368 = v_24258 | v_24367;
assign v_24371 = v_24369 | v_24370;
assign v_24373 = v_24255 | v_24372;
assign v_24376 = v_24374 | v_24375;
assign v_24378 = v_24252 | v_24377;
assign v_24381 = v_24379 | v_24380;
assign v_24383 = v_24249 | v_24382;
assign v_24386 = v_24384 | v_24385;
assign v_24388 = v_24246 | v_24387;
assign v_24391 = v_24389 | v_24390;
assign v_24393 = v_24243 | v_24392;
assign v_24396 = v_24394 | v_24395;
assign v_24398 = v_24240 | v_24397;
assign v_24401 = v_24399 | v_24400;
assign v_24403 = v_24237 | v_24402;
assign v_24406 = v_24404 | v_24405;
assign v_24408 = v_24234 | v_24407;
assign v_24411 = v_24409 | v_24410;
assign v_24413 = v_24231 | v_24412;
assign v_24416 = v_24414 | v_24415;
assign v_24418 = v_24228 | v_24417;
assign v_24421 = v_24419 | v_24420;
assign v_24423 = v_24225 | v_24422;
assign v_24426 = v_24424 | v_24425;
assign v_24428 = v_24222 | v_24427;
assign v_24431 = v_24429 | v_24430;
assign v_24433 = v_24219 | v_24432;
assign v_24436 = v_24434 | v_24435;
assign v_24438 = v_24216 | v_24437;
assign v_24441 = v_24439 | v_24440;
assign v_24443 = v_24213 | v_24442;
assign v_24446 = v_24444 | v_24445;
assign v_24448 = v_24210 | v_24447;
assign v_24451 = v_24209 | v_24450;
assign v_24505 = v_24502 | v_24504;
assign v_24507 = v_24501 | v_24506;
assign v_24509 = v_24499 | v_24508;
assign v_24511 = v_24506 | v_24510;
assign v_24513 = v_24498 | v_24512;
assign v_24515 = v_24496 | v_24514;
assign v_24517 = v_24512 | v_24516;
assign v_24519 = v_24495 | v_24518;
assign v_24521 = v_24493 | v_24520;
assign v_24523 = v_24518 | v_24522;
assign v_24525 = v_24492 | v_24524;
assign v_24527 = v_24490 | v_24526;
assign v_24529 = v_24524 | v_24528;
assign v_24531 = v_24489 | v_24530;
assign v_24533 = v_24487 | v_24532;
assign v_24535 = v_24530 | v_24534;
assign v_24537 = v_24486 | v_24536;
assign v_24539 = v_24484 | v_24538;
assign v_24541 = v_24536 | v_24540;
assign v_24543 = v_24483 | v_24542;
assign v_24545 = v_24481 | v_24544;
assign v_24547 = v_24542 | v_24546;
assign v_24549 = v_24480 | v_24548;
assign v_24551 = v_24478 | v_24550;
assign v_24553 = v_24548 | v_24552;
assign v_24555 = v_24477 | v_24554;
assign v_24557 = v_24475 | v_24556;
assign v_24559 = v_24554 | v_24558;
assign v_24561 = v_24474 | v_24560;
assign v_24563 = v_24472 | v_24562;
assign v_24565 = v_24560 | v_24564;
assign v_24567 = v_24471 | v_24566;
assign v_24569 = v_24469 | v_24568;
assign v_24571 = v_24566 | v_24570;
assign v_24573 = v_24468 | v_24572;
assign v_24575 = v_24466 | v_24574;
assign v_24577 = v_24572 | v_24576;
assign v_24579 = v_24465 | v_24578;
assign v_24581 = v_24463 | v_24580;
assign v_24583 = v_24578 | v_24582;
assign v_24585 = v_24462 | v_24584;
assign v_24587 = v_24460 | v_24586;
assign v_24589 = v_24584 | v_24588;
assign v_24591 = v_24459 | v_24590;
assign v_24593 = v_24457 | v_24592;
assign v_24595 = v_24590 | v_24594;
assign v_24597 = v_24456 | v_24596;
assign v_24599 = v_24454 | v_24598;
assign v_24601 = v_24596 | v_24600;
assign v_24604 = ~v_24453 | v_24603;
assign v_24611 = v_24501 | v_24610;
assign v_24614 = v_24612 | v_24613;
assign v_24616 = v_24498 | v_24615;
assign v_24619 = v_24617 | v_24618;
assign v_24621 = v_24495 | v_24620;
assign v_24624 = v_24622 | v_24623;
assign v_24626 = v_24492 | v_24625;
assign v_24629 = v_24627 | v_24628;
assign v_24631 = v_24489 | v_24630;
assign v_24634 = v_24632 | v_24633;
assign v_24636 = v_24486 | v_24635;
assign v_24639 = v_24637 | v_24638;
assign v_24641 = v_24483 | v_24640;
assign v_24644 = v_24642 | v_24643;
assign v_24646 = v_24480 | v_24645;
assign v_24649 = v_24647 | v_24648;
assign v_24651 = v_24477 | v_24650;
assign v_24654 = v_24652 | v_24653;
assign v_24656 = v_24474 | v_24655;
assign v_24659 = v_24657 | v_24658;
assign v_24661 = v_24471 | v_24660;
assign v_24664 = v_24662 | v_24663;
assign v_24666 = v_24468 | v_24665;
assign v_24669 = v_24667 | v_24668;
assign v_24671 = v_24465 | v_24670;
assign v_24674 = v_24672 | v_24673;
assign v_24676 = v_24462 | v_24675;
assign v_24679 = v_24677 | v_24678;
assign v_24681 = v_24459 | v_24680;
assign v_24684 = v_24682 | v_24683;
assign v_24686 = v_24456 | v_24685;
assign v_24689 = v_24687 | v_24688;
assign v_24691 = v_24453 | v_24690;
assign v_24694 = v_24452 | v_24693;
assign v_24748 = v_24745 | v_24747;
assign v_24750 = v_24744 | v_24749;
assign v_24752 = v_24742 | v_24751;
assign v_24754 = v_24749 | v_24753;
assign v_24756 = v_24741 | v_24755;
assign v_24758 = v_24739 | v_24757;
assign v_24760 = v_24755 | v_24759;
assign v_24762 = v_24738 | v_24761;
assign v_24764 = v_24736 | v_24763;
assign v_24766 = v_24761 | v_24765;
assign v_24768 = v_24735 | v_24767;
assign v_24770 = v_24733 | v_24769;
assign v_24772 = v_24767 | v_24771;
assign v_24774 = v_24732 | v_24773;
assign v_24776 = v_24730 | v_24775;
assign v_24778 = v_24773 | v_24777;
assign v_24780 = v_24729 | v_24779;
assign v_24782 = v_24727 | v_24781;
assign v_24784 = v_24779 | v_24783;
assign v_24786 = v_24726 | v_24785;
assign v_24788 = v_24724 | v_24787;
assign v_24790 = v_24785 | v_24789;
assign v_24792 = v_24723 | v_24791;
assign v_24794 = v_24721 | v_24793;
assign v_24796 = v_24791 | v_24795;
assign v_24798 = v_24720 | v_24797;
assign v_24800 = v_24718 | v_24799;
assign v_24802 = v_24797 | v_24801;
assign v_24804 = v_24717 | v_24803;
assign v_24806 = v_24715 | v_24805;
assign v_24808 = v_24803 | v_24807;
assign v_24810 = v_24714 | v_24809;
assign v_24812 = v_24712 | v_24811;
assign v_24814 = v_24809 | v_24813;
assign v_24816 = v_24711 | v_24815;
assign v_24818 = v_24709 | v_24817;
assign v_24820 = v_24815 | v_24819;
assign v_24822 = v_24708 | v_24821;
assign v_24824 = v_24706 | v_24823;
assign v_24826 = v_24821 | v_24825;
assign v_24828 = v_24705 | v_24827;
assign v_24830 = v_24703 | v_24829;
assign v_24832 = v_24827 | v_24831;
assign v_24834 = v_24702 | v_24833;
assign v_24836 = v_24700 | v_24835;
assign v_24838 = v_24833 | v_24837;
assign v_24840 = v_24699 | v_24839;
assign v_24842 = v_24697 | v_24841;
assign v_24844 = v_24839 | v_24843;
assign v_24847 = ~v_24696 | v_24846;
assign v_24854 = v_24744 | v_24853;
assign v_24857 = v_24855 | v_24856;
assign v_24859 = v_24741 | v_24858;
assign v_24862 = v_24860 | v_24861;
assign v_24864 = v_24738 | v_24863;
assign v_24867 = v_24865 | v_24866;
assign v_24869 = v_24735 | v_24868;
assign v_24872 = v_24870 | v_24871;
assign v_24874 = v_24732 | v_24873;
assign v_24877 = v_24875 | v_24876;
assign v_24879 = v_24729 | v_24878;
assign v_24882 = v_24880 | v_24881;
assign v_24884 = v_24726 | v_24883;
assign v_24887 = v_24885 | v_24886;
assign v_24889 = v_24723 | v_24888;
assign v_24892 = v_24890 | v_24891;
assign v_24894 = v_24720 | v_24893;
assign v_24897 = v_24895 | v_24896;
assign v_24899 = v_24717 | v_24898;
assign v_24902 = v_24900 | v_24901;
assign v_24904 = v_24714 | v_24903;
assign v_24907 = v_24905 | v_24906;
assign v_24909 = v_24711 | v_24908;
assign v_24912 = v_24910 | v_24911;
assign v_24914 = v_24708 | v_24913;
assign v_24917 = v_24915 | v_24916;
assign v_24919 = v_24705 | v_24918;
assign v_24922 = v_24920 | v_24921;
assign v_24924 = v_24702 | v_24923;
assign v_24927 = v_24925 | v_24926;
assign v_24929 = v_24699 | v_24928;
assign v_24932 = v_24930 | v_24931;
assign v_24934 = v_24696 | v_24933;
assign v_24937 = v_24695 | v_24936;
assign v_24990 = v_24987 | v_24989;
assign v_24992 = v_24986 | v_24991;
assign v_24994 = v_24984 | v_24993;
assign v_24996 = v_24991 | v_24995;
assign v_24998 = v_24983 | v_24997;
assign v_25000 = v_24981 | v_24999;
assign v_25002 = v_24997 | v_25001;
assign v_25004 = v_24980 | v_25003;
assign v_25006 = v_24978 | v_25005;
assign v_25008 = v_25003 | v_25007;
assign v_25010 = v_24977 | v_25009;
assign v_25012 = v_24975 | v_25011;
assign v_25014 = v_25009 | v_25013;
assign v_25016 = v_24974 | v_25015;
assign v_25018 = v_24972 | v_25017;
assign v_25020 = v_25015 | v_25019;
assign v_25022 = v_24971 | v_25021;
assign v_25024 = v_24969 | v_25023;
assign v_25026 = v_25021 | v_25025;
assign v_25028 = v_24968 | v_25027;
assign v_25030 = v_24966 | v_25029;
assign v_25032 = v_25027 | v_25031;
assign v_25034 = v_24965 | v_25033;
assign v_25036 = v_24963 | v_25035;
assign v_25038 = v_25033 | v_25037;
assign v_25040 = v_24962 | v_25039;
assign v_25042 = v_24960 | v_25041;
assign v_25044 = v_25039 | v_25043;
assign v_25046 = v_24959 | v_25045;
assign v_25048 = v_24957 | v_25047;
assign v_25050 = v_25045 | v_25049;
assign v_25052 = v_24956 | v_25051;
assign v_25054 = v_24954 | v_25053;
assign v_25056 = v_25051 | v_25055;
assign v_25058 = v_24953 | v_25057;
assign v_25060 = v_24951 | v_25059;
assign v_25062 = v_25057 | v_25061;
assign v_25064 = v_24950 | v_25063;
assign v_25066 = v_24948 | v_25065;
assign v_25068 = v_25063 | v_25067;
assign v_25070 = v_24947 | v_25069;
assign v_25072 = v_24945 | v_25071;
assign v_25074 = v_25069 | v_25073;
assign v_25076 = v_24944 | v_25075;
assign v_25078 = v_24942 | v_25077;
assign v_25080 = v_25075 | v_25079;
assign v_25082 = v_24941 | v_25081;
assign v_25084 = v_24939 | v_25083;
assign v_25086 = v_25081 | v_25085;
assign v_25090 = v_25087 | v_25089;
assign v_25097 = v_24986 | v_25096;
assign v_25100 = v_25098 | v_25099;
assign v_25102 = v_24983 | v_25101;
assign v_25105 = v_25103 | v_25104;
assign v_25107 = v_24980 | v_25106;
assign v_25110 = v_25108 | v_25109;
assign v_25112 = v_24977 | v_25111;
assign v_25115 = v_25113 | v_25114;
assign v_25117 = v_24974 | v_25116;
assign v_25120 = v_25118 | v_25119;
assign v_25122 = v_24971 | v_25121;
assign v_25125 = v_25123 | v_25124;
assign v_25127 = v_24968 | v_25126;
assign v_25130 = v_25128 | v_25129;
assign v_25132 = v_24965 | v_25131;
assign v_25135 = v_25133 | v_25134;
assign v_25137 = v_24962 | v_25136;
assign v_25140 = v_25138 | v_25139;
assign v_25142 = v_24959 | v_25141;
assign v_25145 = v_25143 | v_25144;
assign v_25147 = v_24956 | v_25146;
assign v_25150 = v_25148 | v_25149;
assign v_25152 = v_24953 | v_25151;
assign v_25155 = v_25153 | v_25154;
assign v_25157 = v_24950 | v_25156;
assign v_25160 = v_25158 | v_25159;
assign v_25162 = v_24947 | v_25161;
assign v_25165 = v_25163 | v_25164;
assign v_25167 = v_24944 | v_25166;
assign v_25170 = v_25168 | v_25169;
assign v_25172 = v_24941 | v_25171;
assign v_25175 = v_25173 | v_25174;
assign v_25177 = v_25175 | v_25176;
assign v_25180 = v_24938 | v_25179;
assign v_25251 = v_25248 | v_25250;
assign v_25253 = v_25246 | v_25252;
assign v_25255 = v_25244 | v_25254;
assign v_25257 = v_25252 | v_25256;
assign v_25259 = v_25242 | v_25258;
assign v_25261 = v_25240 | v_25260;
assign v_25263 = v_25258 | v_25262;
assign v_25265 = v_25238 | v_25264;
assign v_25267 = v_25236 | v_25266;
assign v_25269 = v_25264 | v_25268;
assign v_25271 = v_25234 | v_25270;
assign v_25273 = v_25232 | v_25272;
assign v_25275 = v_25270 | v_25274;
assign v_25277 = v_25230 | v_25276;
assign v_25279 = v_25228 | v_25278;
assign v_25281 = v_25276 | v_25280;
assign v_25283 = v_25226 | v_25282;
assign v_25285 = v_25224 | v_25284;
assign v_25287 = v_25282 | v_25286;
assign v_25289 = v_25222 | v_25288;
assign v_25291 = v_25220 | v_25290;
assign v_25293 = v_25288 | v_25292;
assign v_25295 = v_25218 | v_25294;
assign v_25297 = v_25216 | v_25296;
assign v_25299 = v_25294 | v_25298;
assign v_25301 = v_25214 | v_25300;
assign v_25303 = v_25212 | v_25302;
assign v_25305 = v_25300 | v_25304;
assign v_25307 = v_25210 | v_25306;
assign v_25309 = v_25208 | v_25308;
assign v_25311 = v_25306 | v_25310;
assign v_25313 = v_25206 | v_25312;
assign v_25315 = v_25204 | v_25314;
assign v_25317 = v_25312 | v_25316;
assign v_25319 = v_25202 | v_25318;
assign v_25321 = v_25200 | v_25320;
assign v_25323 = v_25318 | v_25322;
assign v_25325 = v_25198 | v_25324;
assign v_25327 = v_25195 | v_25326;
assign v_25329 = v_25324 | v_25328;
assign v_25331 = v_25194 | v_25330;
assign v_25333 = v_25191 | v_25332;
assign v_25335 = v_25330 | v_25334;
assign v_25337 = v_25190 | v_25336;
assign v_25339 = v_25187 | v_25338;
assign v_25341 = v_25336 | v_25340;
assign v_25343 = v_25186 | v_25342;
assign v_25345 = v_25183 | v_25344;
assign v_25347 = v_25342 | v_25346;
assign v_25350 = ~v_25182 | v_25349;
assign v_25357 = v_25246 | v_25356;
assign v_25360 = v_25358 | v_25359;
assign v_25362 = v_25242 | v_25361;
assign v_25365 = v_25363 | v_25364;
assign v_25367 = v_25238 | v_25366;
assign v_25370 = v_25368 | v_25369;
assign v_25372 = v_25234 | v_25371;
assign v_25375 = v_25373 | v_25374;
assign v_25377 = v_25230 | v_25376;
assign v_25380 = v_25378 | v_25379;
assign v_25382 = v_25226 | v_25381;
assign v_25385 = v_25383 | v_25384;
assign v_25387 = v_25222 | v_25386;
assign v_25390 = v_25388 | v_25389;
assign v_25392 = v_25218 | v_25391;
assign v_25395 = v_25393 | v_25394;
assign v_25397 = v_25214 | v_25396;
assign v_25400 = v_25398 | v_25399;
assign v_25402 = v_25210 | v_25401;
assign v_25405 = v_25403 | v_25404;
assign v_25407 = v_25206 | v_25406;
assign v_25410 = v_25408 | v_25409;
assign v_25412 = v_25202 | v_25411;
assign v_25415 = v_25413 | v_25414;
assign v_25417 = v_25198 | v_25416;
assign v_25420 = v_25418 | v_25419;
assign v_25422 = v_25194 | v_25421;
assign v_25425 = v_25423 | v_25424;
assign v_25427 = v_25190 | v_25426;
assign v_25430 = v_25428 | v_25429;
assign v_25432 = v_25186 | v_25431;
assign v_25435 = v_25433 | v_25434;
assign v_25437 = v_25182 | v_25436;
assign v_25440 = v_25181 | v_25439;
assign v_25494 = v_25491 | v_25493;
assign v_25496 = v_25490 | v_25495;
assign v_25498 = v_25488 | v_25497;
assign v_25500 = v_25495 | v_25499;
assign v_25502 = v_25487 | v_25501;
assign v_25504 = v_25485 | v_25503;
assign v_25506 = v_25501 | v_25505;
assign v_25508 = v_25484 | v_25507;
assign v_25510 = v_25482 | v_25509;
assign v_25512 = v_25507 | v_25511;
assign v_25514 = v_25481 | v_25513;
assign v_25516 = v_25479 | v_25515;
assign v_25518 = v_25513 | v_25517;
assign v_25520 = v_25478 | v_25519;
assign v_25522 = v_25476 | v_25521;
assign v_25524 = v_25519 | v_25523;
assign v_25526 = v_25475 | v_25525;
assign v_25528 = v_25473 | v_25527;
assign v_25530 = v_25525 | v_25529;
assign v_25532 = v_25472 | v_25531;
assign v_25534 = v_25470 | v_25533;
assign v_25536 = v_25531 | v_25535;
assign v_25538 = v_25469 | v_25537;
assign v_25540 = v_25467 | v_25539;
assign v_25542 = v_25537 | v_25541;
assign v_25544 = v_25466 | v_25543;
assign v_25546 = v_25464 | v_25545;
assign v_25548 = v_25543 | v_25547;
assign v_25550 = v_25463 | v_25549;
assign v_25552 = v_25461 | v_25551;
assign v_25554 = v_25549 | v_25553;
assign v_25556 = v_25460 | v_25555;
assign v_25558 = v_25458 | v_25557;
assign v_25560 = v_25555 | v_25559;
assign v_25562 = v_25457 | v_25561;
assign v_25564 = v_25455 | v_25563;
assign v_25566 = v_25561 | v_25565;
assign v_25568 = v_25454 | v_25567;
assign v_25570 = v_25452 | v_25569;
assign v_25572 = v_25567 | v_25571;
assign v_25574 = v_25451 | v_25573;
assign v_25576 = v_25449 | v_25575;
assign v_25578 = v_25573 | v_25577;
assign v_25580 = v_25448 | v_25579;
assign v_25582 = v_25446 | v_25581;
assign v_25584 = v_25579 | v_25583;
assign v_25586 = v_25445 | v_25585;
assign v_25588 = v_25443 | v_25587;
assign v_25590 = v_25585 | v_25589;
assign v_25593 = ~v_25442 | v_25592;
assign v_25600 = v_25490 | v_25599;
assign v_25603 = v_25601 | v_25602;
assign v_25605 = v_25487 | v_25604;
assign v_25608 = v_25606 | v_25607;
assign v_25610 = v_25484 | v_25609;
assign v_25613 = v_25611 | v_25612;
assign v_25615 = v_25481 | v_25614;
assign v_25618 = v_25616 | v_25617;
assign v_25620 = v_25478 | v_25619;
assign v_25623 = v_25621 | v_25622;
assign v_25625 = v_25475 | v_25624;
assign v_25628 = v_25626 | v_25627;
assign v_25630 = v_25472 | v_25629;
assign v_25633 = v_25631 | v_25632;
assign v_25635 = v_25469 | v_25634;
assign v_25638 = v_25636 | v_25637;
assign v_25640 = v_25466 | v_25639;
assign v_25643 = v_25641 | v_25642;
assign v_25645 = v_25463 | v_25644;
assign v_25648 = v_25646 | v_25647;
assign v_25650 = v_25460 | v_25649;
assign v_25653 = v_25651 | v_25652;
assign v_25655 = v_25457 | v_25654;
assign v_25658 = v_25656 | v_25657;
assign v_25660 = v_25454 | v_25659;
assign v_25663 = v_25661 | v_25662;
assign v_25665 = v_25451 | v_25664;
assign v_25668 = v_25666 | v_25667;
assign v_25670 = v_25448 | v_25669;
assign v_25673 = v_25671 | v_25672;
assign v_25675 = v_25445 | v_25674;
assign v_25678 = v_25676 | v_25677;
assign v_25680 = v_25442 | v_25679;
assign v_25683 = v_25441 | v_25682;
assign v_25737 = v_25734 | v_25736;
assign v_25739 = v_25733 | v_25738;
assign v_25741 = v_25731 | v_25740;
assign v_25743 = v_25738 | v_25742;
assign v_25745 = v_25730 | v_25744;
assign v_25747 = v_25728 | v_25746;
assign v_25749 = v_25744 | v_25748;
assign v_25751 = v_25727 | v_25750;
assign v_25753 = v_25725 | v_25752;
assign v_25755 = v_25750 | v_25754;
assign v_25757 = v_25724 | v_25756;
assign v_25759 = v_25722 | v_25758;
assign v_25761 = v_25756 | v_25760;
assign v_25763 = v_25721 | v_25762;
assign v_25765 = v_25719 | v_25764;
assign v_25767 = v_25762 | v_25766;
assign v_25769 = v_25718 | v_25768;
assign v_25771 = v_25716 | v_25770;
assign v_25773 = v_25768 | v_25772;
assign v_25775 = v_25715 | v_25774;
assign v_25777 = v_25713 | v_25776;
assign v_25779 = v_25774 | v_25778;
assign v_25781 = v_25712 | v_25780;
assign v_25783 = v_25710 | v_25782;
assign v_25785 = v_25780 | v_25784;
assign v_25787 = v_25709 | v_25786;
assign v_25789 = v_25707 | v_25788;
assign v_25791 = v_25786 | v_25790;
assign v_25793 = v_25706 | v_25792;
assign v_25795 = v_25704 | v_25794;
assign v_25797 = v_25792 | v_25796;
assign v_25799 = v_25703 | v_25798;
assign v_25801 = v_25701 | v_25800;
assign v_25803 = v_25798 | v_25802;
assign v_25805 = v_25700 | v_25804;
assign v_25807 = v_25698 | v_25806;
assign v_25809 = v_25804 | v_25808;
assign v_25811 = v_25697 | v_25810;
assign v_25813 = v_25695 | v_25812;
assign v_25815 = v_25810 | v_25814;
assign v_25817 = v_25694 | v_25816;
assign v_25819 = v_25692 | v_25818;
assign v_25821 = v_25816 | v_25820;
assign v_25823 = v_25691 | v_25822;
assign v_25825 = v_25689 | v_25824;
assign v_25827 = v_25822 | v_25826;
assign v_25829 = v_25688 | v_25828;
assign v_25831 = v_25686 | v_25830;
assign v_25833 = v_25828 | v_25832;
assign v_25836 = ~v_25685 | v_25835;
assign v_25843 = v_25733 | v_25842;
assign v_25846 = v_25844 | v_25845;
assign v_25848 = v_25730 | v_25847;
assign v_25851 = v_25849 | v_25850;
assign v_25853 = v_25727 | v_25852;
assign v_25856 = v_25854 | v_25855;
assign v_25858 = v_25724 | v_25857;
assign v_25861 = v_25859 | v_25860;
assign v_25863 = v_25721 | v_25862;
assign v_25866 = v_25864 | v_25865;
assign v_25868 = v_25718 | v_25867;
assign v_25871 = v_25869 | v_25870;
assign v_25873 = v_25715 | v_25872;
assign v_25876 = v_25874 | v_25875;
assign v_25878 = v_25712 | v_25877;
assign v_25881 = v_25879 | v_25880;
assign v_25883 = v_25709 | v_25882;
assign v_25886 = v_25884 | v_25885;
assign v_25888 = v_25706 | v_25887;
assign v_25891 = v_25889 | v_25890;
assign v_25893 = v_25703 | v_25892;
assign v_25896 = v_25894 | v_25895;
assign v_25898 = v_25700 | v_25897;
assign v_25901 = v_25899 | v_25900;
assign v_25903 = v_25697 | v_25902;
assign v_25906 = v_25904 | v_25905;
assign v_25908 = v_25694 | v_25907;
assign v_25911 = v_25909 | v_25910;
assign v_25913 = v_25691 | v_25912;
assign v_25916 = v_25914 | v_25915;
assign v_25918 = v_25688 | v_25917;
assign v_25921 = v_25919 | v_25920;
assign v_25923 = v_25685 | v_25922;
assign v_25926 = v_25684 | v_25925;
assign v_25980 = v_25977 | v_25979;
assign v_25982 = v_25976 | v_25981;
assign v_25984 = v_25974 | v_25983;
assign v_25986 = v_25981 | v_25985;
assign v_25988 = v_25973 | v_25987;
assign v_25990 = v_25971 | v_25989;
assign v_25992 = v_25987 | v_25991;
assign v_25994 = v_25970 | v_25993;
assign v_25996 = v_25968 | v_25995;
assign v_25998 = v_25993 | v_25997;
assign v_26000 = v_25967 | v_25999;
assign v_26002 = v_25965 | v_26001;
assign v_26004 = v_25999 | v_26003;
assign v_26006 = v_25964 | v_26005;
assign v_26008 = v_25962 | v_26007;
assign v_26010 = v_26005 | v_26009;
assign v_26012 = v_25961 | v_26011;
assign v_26014 = v_25959 | v_26013;
assign v_26016 = v_26011 | v_26015;
assign v_26018 = v_25958 | v_26017;
assign v_26020 = v_25956 | v_26019;
assign v_26022 = v_26017 | v_26021;
assign v_26024 = v_25955 | v_26023;
assign v_26026 = v_25953 | v_26025;
assign v_26028 = v_26023 | v_26027;
assign v_26030 = v_25952 | v_26029;
assign v_26032 = v_25950 | v_26031;
assign v_26034 = v_26029 | v_26033;
assign v_26036 = v_25949 | v_26035;
assign v_26038 = v_25947 | v_26037;
assign v_26040 = v_26035 | v_26039;
assign v_26042 = v_25946 | v_26041;
assign v_26044 = v_25944 | v_26043;
assign v_26046 = v_26041 | v_26045;
assign v_26048 = v_25943 | v_26047;
assign v_26050 = v_25941 | v_26049;
assign v_26052 = v_26047 | v_26051;
assign v_26054 = v_25940 | v_26053;
assign v_26056 = v_25938 | v_26055;
assign v_26058 = v_26053 | v_26057;
assign v_26060 = v_25937 | v_26059;
assign v_26062 = v_25935 | v_26061;
assign v_26064 = v_26059 | v_26063;
assign v_26066 = v_25934 | v_26065;
assign v_26068 = v_25932 | v_26067;
assign v_26070 = v_26065 | v_26069;
assign v_26072 = v_25931 | v_26071;
assign v_26074 = v_25929 | v_26073;
assign v_26076 = v_26071 | v_26075;
assign v_26079 = ~v_25928 | v_26078;
assign v_26086 = v_25976 | v_26085;
assign v_26089 = v_26087 | v_26088;
assign v_26091 = v_25973 | v_26090;
assign v_26094 = v_26092 | v_26093;
assign v_26096 = v_25970 | v_26095;
assign v_26099 = v_26097 | v_26098;
assign v_26101 = v_25967 | v_26100;
assign v_26104 = v_26102 | v_26103;
assign v_26106 = v_25964 | v_26105;
assign v_26109 = v_26107 | v_26108;
assign v_26111 = v_25961 | v_26110;
assign v_26114 = v_26112 | v_26113;
assign v_26116 = v_25958 | v_26115;
assign v_26119 = v_26117 | v_26118;
assign v_26121 = v_25955 | v_26120;
assign v_26124 = v_26122 | v_26123;
assign v_26126 = v_25952 | v_26125;
assign v_26129 = v_26127 | v_26128;
assign v_26131 = v_25949 | v_26130;
assign v_26134 = v_26132 | v_26133;
assign v_26136 = v_25946 | v_26135;
assign v_26139 = v_26137 | v_26138;
assign v_26141 = v_25943 | v_26140;
assign v_26144 = v_26142 | v_26143;
assign v_26146 = v_25940 | v_26145;
assign v_26149 = v_26147 | v_26148;
assign v_26151 = v_25937 | v_26150;
assign v_26154 = v_26152 | v_26153;
assign v_26156 = v_25934 | v_26155;
assign v_26159 = v_26157 | v_26158;
assign v_26161 = v_25931 | v_26160;
assign v_26164 = v_26162 | v_26163;
assign v_26166 = v_25928 | v_26165;
assign v_26169 = v_25927 | v_26168;
assign v_26223 = v_26220 | v_26222;
assign v_26225 = v_26219 | v_26224;
assign v_26227 = v_26217 | v_26226;
assign v_26229 = v_26224 | v_26228;
assign v_26231 = v_26216 | v_26230;
assign v_26233 = v_26214 | v_26232;
assign v_26235 = v_26230 | v_26234;
assign v_26237 = v_26213 | v_26236;
assign v_26239 = v_26211 | v_26238;
assign v_26241 = v_26236 | v_26240;
assign v_26243 = v_26210 | v_26242;
assign v_26245 = v_26208 | v_26244;
assign v_26247 = v_26242 | v_26246;
assign v_26249 = v_26207 | v_26248;
assign v_26251 = v_26205 | v_26250;
assign v_26253 = v_26248 | v_26252;
assign v_26255 = v_26204 | v_26254;
assign v_26257 = v_26202 | v_26256;
assign v_26259 = v_26254 | v_26258;
assign v_26261 = v_26201 | v_26260;
assign v_26263 = v_26199 | v_26262;
assign v_26265 = v_26260 | v_26264;
assign v_26267 = v_26198 | v_26266;
assign v_26269 = v_26196 | v_26268;
assign v_26271 = v_26266 | v_26270;
assign v_26273 = v_26195 | v_26272;
assign v_26275 = v_26193 | v_26274;
assign v_26277 = v_26272 | v_26276;
assign v_26279 = v_26192 | v_26278;
assign v_26281 = v_26190 | v_26280;
assign v_26283 = v_26278 | v_26282;
assign v_26285 = v_26189 | v_26284;
assign v_26287 = v_26187 | v_26286;
assign v_26289 = v_26284 | v_26288;
assign v_26291 = v_26186 | v_26290;
assign v_26293 = v_26184 | v_26292;
assign v_26295 = v_26290 | v_26294;
assign v_26297 = v_26183 | v_26296;
assign v_26299 = v_26181 | v_26298;
assign v_26301 = v_26296 | v_26300;
assign v_26303 = v_26180 | v_26302;
assign v_26305 = v_26178 | v_26304;
assign v_26307 = v_26302 | v_26306;
assign v_26309 = v_26177 | v_26308;
assign v_26311 = v_26175 | v_26310;
assign v_26313 = v_26308 | v_26312;
assign v_26315 = v_26174 | v_26314;
assign v_26317 = v_26172 | v_26316;
assign v_26319 = v_26314 | v_26318;
assign v_26322 = ~v_26171 | v_26321;
assign v_26329 = v_26219 | v_26328;
assign v_26332 = v_26330 | v_26331;
assign v_26334 = v_26216 | v_26333;
assign v_26337 = v_26335 | v_26336;
assign v_26339 = v_26213 | v_26338;
assign v_26342 = v_26340 | v_26341;
assign v_26344 = v_26210 | v_26343;
assign v_26347 = v_26345 | v_26346;
assign v_26349 = v_26207 | v_26348;
assign v_26352 = v_26350 | v_26351;
assign v_26354 = v_26204 | v_26353;
assign v_26357 = v_26355 | v_26356;
assign v_26359 = v_26201 | v_26358;
assign v_26362 = v_26360 | v_26361;
assign v_26364 = v_26198 | v_26363;
assign v_26367 = v_26365 | v_26366;
assign v_26369 = v_26195 | v_26368;
assign v_26372 = v_26370 | v_26371;
assign v_26374 = v_26192 | v_26373;
assign v_26377 = v_26375 | v_26376;
assign v_26379 = v_26189 | v_26378;
assign v_26382 = v_26380 | v_26381;
assign v_26384 = v_26186 | v_26383;
assign v_26387 = v_26385 | v_26386;
assign v_26389 = v_26183 | v_26388;
assign v_26392 = v_26390 | v_26391;
assign v_26394 = v_26180 | v_26393;
assign v_26397 = v_26395 | v_26396;
assign v_26399 = v_26177 | v_26398;
assign v_26402 = v_26400 | v_26401;
assign v_26404 = v_26174 | v_26403;
assign v_26407 = v_26405 | v_26406;
assign v_26409 = v_26171 | v_26408;
assign v_26412 = v_26170 | v_26411;
assign v_26466 = v_26463 | v_26465;
assign v_26468 = v_26462 | v_26467;
assign v_26470 = v_26460 | v_26469;
assign v_26472 = v_26467 | v_26471;
assign v_26474 = v_26459 | v_26473;
assign v_26476 = v_26457 | v_26475;
assign v_26478 = v_26473 | v_26477;
assign v_26480 = v_26456 | v_26479;
assign v_26482 = v_26454 | v_26481;
assign v_26484 = v_26479 | v_26483;
assign v_26486 = v_26453 | v_26485;
assign v_26488 = v_26451 | v_26487;
assign v_26490 = v_26485 | v_26489;
assign v_26492 = v_26450 | v_26491;
assign v_26494 = v_26448 | v_26493;
assign v_26496 = v_26491 | v_26495;
assign v_26498 = v_26447 | v_26497;
assign v_26500 = v_26445 | v_26499;
assign v_26502 = v_26497 | v_26501;
assign v_26504 = v_26444 | v_26503;
assign v_26506 = v_26442 | v_26505;
assign v_26508 = v_26503 | v_26507;
assign v_26510 = v_26441 | v_26509;
assign v_26512 = v_26439 | v_26511;
assign v_26514 = v_26509 | v_26513;
assign v_26516 = v_26438 | v_26515;
assign v_26518 = v_26436 | v_26517;
assign v_26520 = v_26515 | v_26519;
assign v_26522 = v_26435 | v_26521;
assign v_26524 = v_26433 | v_26523;
assign v_26526 = v_26521 | v_26525;
assign v_26528 = v_26432 | v_26527;
assign v_26530 = v_26430 | v_26529;
assign v_26532 = v_26527 | v_26531;
assign v_26534 = v_26429 | v_26533;
assign v_26536 = v_26427 | v_26535;
assign v_26538 = v_26533 | v_26537;
assign v_26540 = v_26426 | v_26539;
assign v_26542 = v_26424 | v_26541;
assign v_26544 = v_26539 | v_26543;
assign v_26546 = v_26423 | v_26545;
assign v_26548 = v_26421 | v_26547;
assign v_26550 = v_26545 | v_26549;
assign v_26552 = v_26420 | v_26551;
assign v_26554 = v_26418 | v_26553;
assign v_26556 = v_26551 | v_26555;
assign v_26558 = v_26417 | v_26557;
assign v_26560 = v_26415 | v_26559;
assign v_26562 = v_26557 | v_26561;
assign v_26565 = ~v_26414 | v_26564;
assign v_26572 = v_26462 | v_26571;
assign v_26575 = v_26573 | v_26574;
assign v_26577 = v_26459 | v_26576;
assign v_26580 = v_26578 | v_26579;
assign v_26582 = v_26456 | v_26581;
assign v_26585 = v_26583 | v_26584;
assign v_26587 = v_26453 | v_26586;
assign v_26590 = v_26588 | v_26589;
assign v_26592 = v_26450 | v_26591;
assign v_26595 = v_26593 | v_26594;
assign v_26597 = v_26447 | v_26596;
assign v_26600 = v_26598 | v_26599;
assign v_26602 = v_26444 | v_26601;
assign v_26605 = v_26603 | v_26604;
assign v_26607 = v_26441 | v_26606;
assign v_26610 = v_26608 | v_26609;
assign v_26612 = v_26438 | v_26611;
assign v_26615 = v_26613 | v_26614;
assign v_26617 = v_26435 | v_26616;
assign v_26620 = v_26618 | v_26619;
assign v_26622 = v_26432 | v_26621;
assign v_26625 = v_26623 | v_26624;
assign v_26627 = v_26429 | v_26626;
assign v_26630 = v_26628 | v_26629;
assign v_26632 = v_26426 | v_26631;
assign v_26635 = v_26633 | v_26634;
assign v_26637 = v_26423 | v_26636;
assign v_26640 = v_26638 | v_26639;
assign v_26642 = v_26420 | v_26641;
assign v_26645 = v_26643 | v_26644;
assign v_26647 = v_26417 | v_26646;
assign v_26650 = v_26648 | v_26649;
assign v_26652 = v_26414 | v_26651;
assign v_26655 = v_26413 | v_26654;
assign v_26709 = v_26706 | v_26708;
assign v_26711 = v_26705 | v_26710;
assign v_26713 = v_26703 | v_26712;
assign v_26715 = v_26710 | v_26714;
assign v_26717 = v_26702 | v_26716;
assign v_26719 = v_26700 | v_26718;
assign v_26721 = v_26716 | v_26720;
assign v_26723 = v_26699 | v_26722;
assign v_26725 = v_26697 | v_26724;
assign v_26727 = v_26722 | v_26726;
assign v_26729 = v_26696 | v_26728;
assign v_26731 = v_26694 | v_26730;
assign v_26733 = v_26728 | v_26732;
assign v_26735 = v_26693 | v_26734;
assign v_26737 = v_26691 | v_26736;
assign v_26739 = v_26734 | v_26738;
assign v_26741 = v_26690 | v_26740;
assign v_26743 = v_26688 | v_26742;
assign v_26745 = v_26740 | v_26744;
assign v_26747 = v_26687 | v_26746;
assign v_26749 = v_26685 | v_26748;
assign v_26751 = v_26746 | v_26750;
assign v_26753 = v_26684 | v_26752;
assign v_26755 = v_26682 | v_26754;
assign v_26757 = v_26752 | v_26756;
assign v_26759 = v_26681 | v_26758;
assign v_26761 = v_26679 | v_26760;
assign v_26763 = v_26758 | v_26762;
assign v_26765 = v_26678 | v_26764;
assign v_26767 = v_26676 | v_26766;
assign v_26769 = v_26764 | v_26768;
assign v_26771 = v_26675 | v_26770;
assign v_26773 = v_26673 | v_26772;
assign v_26775 = v_26770 | v_26774;
assign v_26777 = v_26672 | v_26776;
assign v_26779 = v_26670 | v_26778;
assign v_26781 = v_26776 | v_26780;
assign v_26783 = v_26669 | v_26782;
assign v_26785 = v_26667 | v_26784;
assign v_26787 = v_26782 | v_26786;
assign v_26789 = v_26666 | v_26788;
assign v_26791 = v_26664 | v_26790;
assign v_26793 = v_26788 | v_26792;
assign v_26795 = v_26663 | v_26794;
assign v_26797 = v_26661 | v_26796;
assign v_26799 = v_26794 | v_26798;
assign v_26801 = v_26660 | v_26800;
assign v_26803 = v_26658 | v_26802;
assign v_26805 = v_26800 | v_26804;
assign v_26808 = ~v_26657 | v_26807;
assign v_26815 = v_26705 | v_26814;
assign v_26818 = v_26816 | v_26817;
assign v_26820 = v_26702 | v_26819;
assign v_26823 = v_26821 | v_26822;
assign v_26825 = v_26699 | v_26824;
assign v_26828 = v_26826 | v_26827;
assign v_26830 = v_26696 | v_26829;
assign v_26833 = v_26831 | v_26832;
assign v_26835 = v_26693 | v_26834;
assign v_26838 = v_26836 | v_26837;
assign v_26840 = v_26690 | v_26839;
assign v_26843 = v_26841 | v_26842;
assign v_26845 = v_26687 | v_26844;
assign v_26848 = v_26846 | v_26847;
assign v_26850 = v_26684 | v_26849;
assign v_26853 = v_26851 | v_26852;
assign v_26855 = v_26681 | v_26854;
assign v_26858 = v_26856 | v_26857;
assign v_26860 = v_26678 | v_26859;
assign v_26863 = v_26861 | v_26862;
assign v_26865 = v_26675 | v_26864;
assign v_26868 = v_26866 | v_26867;
assign v_26870 = v_26672 | v_26869;
assign v_26873 = v_26871 | v_26872;
assign v_26875 = v_26669 | v_26874;
assign v_26878 = v_26876 | v_26877;
assign v_26880 = v_26666 | v_26879;
assign v_26883 = v_26881 | v_26882;
assign v_26885 = v_26663 | v_26884;
assign v_26888 = v_26886 | v_26887;
assign v_26890 = v_26660 | v_26889;
assign v_26893 = v_26891 | v_26892;
assign v_26895 = v_26657 | v_26894;
assign v_26898 = v_26656 | v_26897;
assign v_26952 = v_26949 | v_26951;
assign v_26954 = v_26948 | v_26953;
assign v_26956 = v_26946 | v_26955;
assign v_26958 = v_26953 | v_26957;
assign v_26960 = v_26945 | v_26959;
assign v_26962 = v_26943 | v_26961;
assign v_26964 = v_26959 | v_26963;
assign v_26966 = v_26942 | v_26965;
assign v_26968 = v_26940 | v_26967;
assign v_26970 = v_26965 | v_26969;
assign v_26972 = v_26939 | v_26971;
assign v_26974 = v_26937 | v_26973;
assign v_26976 = v_26971 | v_26975;
assign v_26978 = v_26936 | v_26977;
assign v_26980 = v_26934 | v_26979;
assign v_26982 = v_26977 | v_26981;
assign v_26984 = v_26933 | v_26983;
assign v_26986 = v_26931 | v_26985;
assign v_26988 = v_26983 | v_26987;
assign v_26990 = v_26930 | v_26989;
assign v_26992 = v_26928 | v_26991;
assign v_26994 = v_26989 | v_26993;
assign v_26996 = v_26927 | v_26995;
assign v_26998 = v_26925 | v_26997;
assign v_27000 = v_26995 | v_26999;
assign v_27002 = v_26924 | v_27001;
assign v_27004 = v_26922 | v_27003;
assign v_27006 = v_27001 | v_27005;
assign v_27008 = v_26921 | v_27007;
assign v_27010 = v_26919 | v_27009;
assign v_27012 = v_27007 | v_27011;
assign v_27014 = v_26918 | v_27013;
assign v_27016 = v_26916 | v_27015;
assign v_27018 = v_27013 | v_27017;
assign v_27020 = v_26915 | v_27019;
assign v_27022 = v_26913 | v_27021;
assign v_27024 = v_27019 | v_27023;
assign v_27026 = v_26912 | v_27025;
assign v_27028 = v_26910 | v_27027;
assign v_27030 = v_27025 | v_27029;
assign v_27032 = v_26909 | v_27031;
assign v_27034 = v_26907 | v_27033;
assign v_27036 = v_27031 | v_27035;
assign v_27038 = v_26906 | v_27037;
assign v_27040 = v_26904 | v_27039;
assign v_27042 = v_27037 | v_27041;
assign v_27044 = v_26903 | v_27043;
assign v_27046 = v_26901 | v_27045;
assign v_27048 = v_27043 | v_27047;
assign v_27051 = ~v_26900 | v_27050;
assign v_27058 = v_26948 | v_27057;
assign v_27061 = v_27059 | v_27060;
assign v_27063 = v_26945 | v_27062;
assign v_27066 = v_27064 | v_27065;
assign v_27068 = v_26942 | v_27067;
assign v_27071 = v_27069 | v_27070;
assign v_27073 = v_26939 | v_27072;
assign v_27076 = v_27074 | v_27075;
assign v_27078 = v_26936 | v_27077;
assign v_27081 = v_27079 | v_27080;
assign v_27083 = v_26933 | v_27082;
assign v_27086 = v_27084 | v_27085;
assign v_27088 = v_26930 | v_27087;
assign v_27091 = v_27089 | v_27090;
assign v_27093 = v_26927 | v_27092;
assign v_27096 = v_27094 | v_27095;
assign v_27098 = v_26924 | v_27097;
assign v_27101 = v_27099 | v_27100;
assign v_27103 = v_26921 | v_27102;
assign v_27106 = v_27104 | v_27105;
assign v_27108 = v_26918 | v_27107;
assign v_27111 = v_27109 | v_27110;
assign v_27113 = v_26915 | v_27112;
assign v_27116 = v_27114 | v_27115;
assign v_27118 = v_26912 | v_27117;
assign v_27121 = v_27119 | v_27120;
assign v_27123 = v_26909 | v_27122;
assign v_27126 = v_27124 | v_27125;
assign v_27128 = v_26906 | v_27127;
assign v_27131 = v_27129 | v_27130;
assign v_27133 = v_26903 | v_27132;
assign v_27136 = v_27134 | v_27135;
assign v_27138 = v_26900 | v_27137;
assign v_27141 = v_26899 | v_27140;
assign v_27195 = v_27192 | v_27194;
assign v_27197 = v_27191 | v_27196;
assign v_27199 = v_27189 | v_27198;
assign v_27201 = v_27196 | v_27200;
assign v_27203 = v_27188 | v_27202;
assign v_27205 = v_27186 | v_27204;
assign v_27207 = v_27202 | v_27206;
assign v_27209 = v_27185 | v_27208;
assign v_27211 = v_27183 | v_27210;
assign v_27213 = v_27208 | v_27212;
assign v_27215 = v_27182 | v_27214;
assign v_27217 = v_27180 | v_27216;
assign v_27219 = v_27214 | v_27218;
assign v_27221 = v_27179 | v_27220;
assign v_27223 = v_27177 | v_27222;
assign v_27225 = v_27220 | v_27224;
assign v_27227 = v_27176 | v_27226;
assign v_27229 = v_27174 | v_27228;
assign v_27231 = v_27226 | v_27230;
assign v_27233 = v_27173 | v_27232;
assign v_27235 = v_27171 | v_27234;
assign v_27237 = v_27232 | v_27236;
assign v_27239 = v_27170 | v_27238;
assign v_27241 = v_27168 | v_27240;
assign v_27243 = v_27238 | v_27242;
assign v_27245 = v_27167 | v_27244;
assign v_27247 = v_27165 | v_27246;
assign v_27249 = v_27244 | v_27248;
assign v_27251 = v_27164 | v_27250;
assign v_27253 = v_27162 | v_27252;
assign v_27255 = v_27250 | v_27254;
assign v_27257 = v_27161 | v_27256;
assign v_27259 = v_27159 | v_27258;
assign v_27261 = v_27256 | v_27260;
assign v_27263 = v_27158 | v_27262;
assign v_27265 = v_27156 | v_27264;
assign v_27267 = v_27262 | v_27266;
assign v_27269 = v_27155 | v_27268;
assign v_27271 = v_27153 | v_27270;
assign v_27273 = v_27268 | v_27272;
assign v_27275 = v_27152 | v_27274;
assign v_27277 = v_27150 | v_27276;
assign v_27279 = v_27274 | v_27278;
assign v_27281 = v_27149 | v_27280;
assign v_27283 = v_27147 | v_27282;
assign v_27285 = v_27280 | v_27284;
assign v_27287 = v_27146 | v_27286;
assign v_27289 = v_27144 | v_27288;
assign v_27291 = v_27286 | v_27290;
assign v_27294 = ~v_27143 | v_27293;
assign v_27301 = v_27191 | v_27300;
assign v_27304 = v_27302 | v_27303;
assign v_27306 = v_27188 | v_27305;
assign v_27309 = v_27307 | v_27308;
assign v_27311 = v_27185 | v_27310;
assign v_27314 = v_27312 | v_27313;
assign v_27316 = v_27182 | v_27315;
assign v_27319 = v_27317 | v_27318;
assign v_27321 = v_27179 | v_27320;
assign v_27324 = v_27322 | v_27323;
assign v_27326 = v_27176 | v_27325;
assign v_27329 = v_27327 | v_27328;
assign v_27331 = v_27173 | v_27330;
assign v_27334 = v_27332 | v_27333;
assign v_27336 = v_27170 | v_27335;
assign v_27339 = v_27337 | v_27338;
assign v_27341 = v_27167 | v_27340;
assign v_27344 = v_27342 | v_27343;
assign v_27346 = v_27164 | v_27345;
assign v_27349 = v_27347 | v_27348;
assign v_27351 = v_27161 | v_27350;
assign v_27354 = v_27352 | v_27353;
assign v_27356 = v_27158 | v_27355;
assign v_27359 = v_27357 | v_27358;
assign v_27361 = v_27155 | v_27360;
assign v_27364 = v_27362 | v_27363;
assign v_27366 = v_27152 | v_27365;
assign v_27369 = v_27367 | v_27368;
assign v_27371 = v_27149 | v_27370;
assign v_27374 = v_27372 | v_27373;
assign v_27376 = v_27146 | v_27375;
assign v_27379 = v_27377 | v_27378;
assign v_27381 = v_27143 | v_27380;
assign v_27384 = v_27142 | v_27383;
assign v_27438 = v_27435 | v_27437;
assign v_27440 = v_27434 | v_27439;
assign v_27442 = v_27432 | v_27441;
assign v_27444 = v_27439 | v_27443;
assign v_27446 = v_27431 | v_27445;
assign v_27448 = v_27429 | v_27447;
assign v_27450 = v_27445 | v_27449;
assign v_27452 = v_27428 | v_27451;
assign v_27454 = v_27426 | v_27453;
assign v_27456 = v_27451 | v_27455;
assign v_27458 = v_27425 | v_27457;
assign v_27460 = v_27423 | v_27459;
assign v_27462 = v_27457 | v_27461;
assign v_27464 = v_27422 | v_27463;
assign v_27466 = v_27420 | v_27465;
assign v_27468 = v_27463 | v_27467;
assign v_27470 = v_27419 | v_27469;
assign v_27472 = v_27417 | v_27471;
assign v_27474 = v_27469 | v_27473;
assign v_27476 = v_27416 | v_27475;
assign v_27478 = v_27414 | v_27477;
assign v_27480 = v_27475 | v_27479;
assign v_27482 = v_27413 | v_27481;
assign v_27484 = v_27411 | v_27483;
assign v_27486 = v_27481 | v_27485;
assign v_27488 = v_27410 | v_27487;
assign v_27490 = v_27408 | v_27489;
assign v_27492 = v_27487 | v_27491;
assign v_27494 = v_27407 | v_27493;
assign v_27496 = v_27405 | v_27495;
assign v_27498 = v_27493 | v_27497;
assign v_27500 = v_27404 | v_27499;
assign v_27502 = v_27402 | v_27501;
assign v_27504 = v_27499 | v_27503;
assign v_27506 = v_27401 | v_27505;
assign v_27508 = v_27399 | v_27507;
assign v_27510 = v_27505 | v_27509;
assign v_27512 = v_27398 | v_27511;
assign v_27514 = v_27396 | v_27513;
assign v_27516 = v_27511 | v_27515;
assign v_27518 = v_27395 | v_27517;
assign v_27520 = v_27393 | v_27519;
assign v_27522 = v_27517 | v_27521;
assign v_27524 = v_27392 | v_27523;
assign v_27526 = v_27390 | v_27525;
assign v_27528 = v_27523 | v_27527;
assign v_27530 = v_27389 | v_27529;
assign v_27532 = v_27387 | v_27531;
assign v_27534 = v_27529 | v_27533;
assign v_27537 = ~v_27386 | v_27536;
assign v_27544 = v_27434 | v_27543;
assign v_27547 = v_27545 | v_27546;
assign v_27549 = v_27431 | v_27548;
assign v_27552 = v_27550 | v_27551;
assign v_27554 = v_27428 | v_27553;
assign v_27557 = v_27555 | v_27556;
assign v_27559 = v_27425 | v_27558;
assign v_27562 = v_27560 | v_27561;
assign v_27564 = v_27422 | v_27563;
assign v_27567 = v_27565 | v_27566;
assign v_27569 = v_27419 | v_27568;
assign v_27572 = v_27570 | v_27571;
assign v_27574 = v_27416 | v_27573;
assign v_27577 = v_27575 | v_27576;
assign v_27579 = v_27413 | v_27578;
assign v_27582 = v_27580 | v_27581;
assign v_27584 = v_27410 | v_27583;
assign v_27587 = v_27585 | v_27586;
assign v_27589 = v_27407 | v_27588;
assign v_27592 = v_27590 | v_27591;
assign v_27594 = v_27404 | v_27593;
assign v_27597 = v_27595 | v_27596;
assign v_27599 = v_27401 | v_27598;
assign v_27602 = v_27600 | v_27601;
assign v_27604 = v_27398 | v_27603;
assign v_27607 = v_27605 | v_27606;
assign v_27609 = v_27395 | v_27608;
assign v_27612 = v_27610 | v_27611;
assign v_27614 = v_27392 | v_27613;
assign v_27617 = v_27615 | v_27616;
assign v_27619 = v_27389 | v_27618;
assign v_27622 = v_27620 | v_27621;
assign v_27624 = v_27386 | v_27623;
assign v_27627 = v_27385 | v_27626;
assign v_27681 = v_27678 | v_27680;
assign v_27683 = v_27677 | v_27682;
assign v_27685 = v_27675 | v_27684;
assign v_27687 = v_27682 | v_27686;
assign v_27689 = v_27674 | v_27688;
assign v_27691 = v_27672 | v_27690;
assign v_27693 = v_27688 | v_27692;
assign v_27695 = v_27671 | v_27694;
assign v_27697 = v_27669 | v_27696;
assign v_27699 = v_27694 | v_27698;
assign v_27701 = v_27668 | v_27700;
assign v_27703 = v_27666 | v_27702;
assign v_27705 = v_27700 | v_27704;
assign v_27707 = v_27665 | v_27706;
assign v_27709 = v_27663 | v_27708;
assign v_27711 = v_27706 | v_27710;
assign v_27713 = v_27662 | v_27712;
assign v_27715 = v_27660 | v_27714;
assign v_27717 = v_27712 | v_27716;
assign v_27719 = v_27659 | v_27718;
assign v_27721 = v_27657 | v_27720;
assign v_27723 = v_27718 | v_27722;
assign v_27725 = v_27656 | v_27724;
assign v_27727 = v_27654 | v_27726;
assign v_27729 = v_27724 | v_27728;
assign v_27731 = v_27653 | v_27730;
assign v_27733 = v_27651 | v_27732;
assign v_27735 = v_27730 | v_27734;
assign v_27737 = v_27650 | v_27736;
assign v_27739 = v_27648 | v_27738;
assign v_27741 = v_27736 | v_27740;
assign v_27743 = v_27647 | v_27742;
assign v_27745 = v_27645 | v_27744;
assign v_27747 = v_27742 | v_27746;
assign v_27749 = v_27644 | v_27748;
assign v_27751 = v_27642 | v_27750;
assign v_27753 = v_27748 | v_27752;
assign v_27755 = v_27641 | v_27754;
assign v_27757 = v_27639 | v_27756;
assign v_27759 = v_27754 | v_27758;
assign v_27761 = v_27638 | v_27760;
assign v_27763 = v_27636 | v_27762;
assign v_27765 = v_27760 | v_27764;
assign v_27767 = v_27635 | v_27766;
assign v_27769 = v_27633 | v_27768;
assign v_27771 = v_27766 | v_27770;
assign v_27773 = v_27632 | v_27772;
assign v_27775 = v_27630 | v_27774;
assign v_27777 = v_27772 | v_27776;
assign v_27780 = ~v_27629 | v_27779;
assign v_27787 = v_27677 | v_27786;
assign v_27790 = v_27788 | v_27789;
assign v_27792 = v_27674 | v_27791;
assign v_27795 = v_27793 | v_27794;
assign v_27797 = v_27671 | v_27796;
assign v_27800 = v_27798 | v_27799;
assign v_27802 = v_27668 | v_27801;
assign v_27805 = v_27803 | v_27804;
assign v_27807 = v_27665 | v_27806;
assign v_27810 = v_27808 | v_27809;
assign v_27812 = v_27662 | v_27811;
assign v_27815 = v_27813 | v_27814;
assign v_27817 = v_27659 | v_27816;
assign v_27820 = v_27818 | v_27819;
assign v_27822 = v_27656 | v_27821;
assign v_27825 = v_27823 | v_27824;
assign v_27827 = v_27653 | v_27826;
assign v_27830 = v_27828 | v_27829;
assign v_27832 = v_27650 | v_27831;
assign v_27835 = v_27833 | v_27834;
assign v_27837 = v_27647 | v_27836;
assign v_27840 = v_27838 | v_27839;
assign v_27842 = v_27644 | v_27841;
assign v_27845 = v_27843 | v_27844;
assign v_27847 = v_27641 | v_27846;
assign v_27850 = v_27848 | v_27849;
assign v_27852 = v_27638 | v_27851;
assign v_27855 = v_27853 | v_27854;
assign v_27857 = v_27635 | v_27856;
assign v_27860 = v_27858 | v_27859;
assign v_27862 = v_27632 | v_27861;
assign v_27865 = v_27863 | v_27864;
assign v_27867 = v_27629 | v_27866;
assign v_27870 = v_27628 | v_27869;
assign v_27924 = v_27921 | v_27923;
assign v_27926 = v_27920 | v_27925;
assign v_27928 = v_27918 | v_27927;
assign v_27930 = v_27925 | v_27929;
assign v_27932 = v_27917 | v_27931;
assign v_27934 = v_27915 | v_27933;
assign v_27936 = v_27931 | v_27935;
assign v_27938 = v_27914 | v_27937;
assign v_27940 = v_27912 | v_27939;
assign v_27942 = v_27937 | v_27941;
assign v_27944 = v_27911 | v_27943;
assign v_27946 = v_27909 | v_27945;
assign v_27948 = v_27943 | v_27947;
assign v_27950 = v_27908 | v_27949;
assign v_27952 = v_27906 | v_27951;
assign v_27954 = v_27949 | v_27953;
assign v_27956 = v_27905 | v_27955;
assign v_27958 = v_27903 | v_27957;
assign v_27960 = v_27955 | v_27959;
assign v_27962 = v_27902 | v_27961;
assign v_27964 = v_27900 | v_27963;
assign v_27966 = v_27961 | v_27965;
assign v_27968 = v_27899 | v_27967;
assign v_27970 = v_27897 | v_27969;
assign v_27972 = v_27967 | v_27971;
assign v_27974 = v_27896 | v_27973;
assign v_27976 = v_27894 | v_27975;
assign v_27978 = v_27973 | v_27977;
assign v_27980 = v_27893 | v_27979;
assign v_27982 = v_27891 | v_27981;
assign v_27984 = v_27979 | v_27983;
assign v_27986 = v_27890 | v_27985;
assign v_27988 = v_27888 | v_27987;
assign v_27990 = v_27985 | v_27989;
assign v_27992 = v_27887 | v_27991;
assign v_27994 = v_27885 | v_27993;
assign v_27996 = v_27991 | v_27995;
assign v_27998 = v_27884 | v_27997;
assign v_28000 = v_27882 | v_27999;
assign v_28002 = v_27997 | v_28001;
assign v_28004 = v_27881 | v_28003;
assign v_28006 = v_27879 | v_28005;
assign v_28008 = v_28003 | v_28007;
assign v_28010 = v_27878 | v_28009;
assign v_28012 = v_27876 | v_28011;
assign v_28014 = v_28009 | v_28013;
assign v_28016 = v_27875 | v_28015;
assign v_28018 = v_27873 | v_28017;
assign v_28020 = v_28015 | v_28019;
assign v_28023 = ~v_27872 | v_28022;
assign v_28030 = v_27920 | v_28029;
assign v_28033 = v_28031 | v_28032;
assign v_28035 = v_27917 | v_28034;
assign v_28038 = v_28036 | v_28037;
assign v_28040 = v_27914 | v_28039;
assign v_28043 = v_28041 | v_28042;
assign v_28045 = v_27911 | v_28044;
assign v_28048 = v_28046 | v_28047;
assign v_28050 = v_27908 | v_28049;
assign v_28053 = v_28051 | v_28052;
assign v_28055 = v_27905 | v_28054;
assign v_28058 = v_28056 | v_28057;
assign v_28060 = v_27902 | v_28059;
assign v_28063 = v_28061 | v_28062;
assign v_28065 = v_27899 | v_28064;
assign v_28068 = v_28066 | v_28067;
assign v_28070 = v_27896 | v_28069;
assign v_28073 = v_28071 | v_28072;
assign v_28075 = v_27893 | v_28074;
assign v_28078 = v_28076 | v_28077;
assign v_28080 = v_27890 | v_28079;
assign v_28083 = v_28081 | v_28082;
assign v_28085 = v_27887 | v_28084;
assign v_28088 = v_28086 | v_28087;
assign v_28090 = v_27884 | v_28089;
assign v_28093 = v_28091 | v_28092;
assign v_28095 = v_27881 | v_28094;
assign v_28098 = v_28096 | v_28097;
assign v_28100 = v_27878 | v_28099;
assign v_28103 = v_28101 | v_28102;
assign v_28105 = v_27875 | v_28104;
assign v_28108 = v_28106 | v_28107;
assign v_28110 = v_27872 | v_28109;
assign v_28113 = v_27871 | v_28112;
assign v_28167 = v_28164 | v_28166;
assign v_28169 = v_28163 | v_28168;
assign v_28171 = v_28161 | v_28170;
assign v_28173 = v_28168 | v_28172;
assign v_28175 = v_28160 | v_28174;
assign v_28177 = v_28158 | v_28176;
assign v_28179 = v_28174 | v_28178;
assign v_28181 = v_28157 | v_28180;
assign v_28183 = v_28155 | v_28182;
assign v_28185 = v_28180 | v_28184;
assign v_28187 = v_28154 | v_28186;
assign v_28189 = v_28152 | v_28188;
assign v_28191 = v_28186 | v_28190;
assign v_28193 = v_28151 | v_28192;
assign v_28195 = v_28149 | v_28194;
assign v_28197 = v_28192 | v_28196;
assign v_28199 = v_28148 | v_28198;
assign v_28201 = v_28146 | v_28200;
assign v_28203 = v_28198 | v_28202;
assign v_28205 = v_28145 | v_28204;
assign v_28207 = v_28143 | v_28206;
assign v_28209 = v_28204 | v_28208;
assign v_28211 = v_28142 | v_28210;
assign v_28213 = v_28140 | v_28212;
assign v_28215 = v_28210 | v_28214;
assign v_28217 = v_28139 | v_28216;
assign v_28219 = v_28137 | v_28218;
assign v_28221 = v_28216 | v_28220;
assign v_28223 = v_28136 | v_28222;
assign v_28225 = v_28134 | v_28224;
assign v_28227 = v_28222 | v_28226;
assign v_28229 = v_28133 | v_28228;
assign v_28231 = v_28131 | v_28230;
assign v_28233 = v_28228 | v_28232;
assign v_28235 = v_28130 | v_28234;
assign v_28237 = v_28128 | v_28236;
assign v_28239 = v_28234 | v_28238;
assign v_28241 = v_28127 | v_28240;
assign v_28243 = v_28125 | v_28242;
assign v_28245 = v_28240 | v_28244;
assign v_28247 = v_28124 | v_28246;
assign v_28249 = v_28122 | v_28248;
assign v_28251 = v_28246 | v_28250;
assign v_28253 = v_28121 | v_28252;
assign v_28255 = v_28119 | v_28254;
assign v_28257 = v_28252 | v_28256;
assign v_28259 = v_28118 | v_28258;
assign v_28261 = v_28116 | v_28260;
assign v_28263 = v_28258 | v_28262;
assign v_28266 = ~v_28115 | v_28265;
assign v_28273 = v_28163 | v_28272;
assign v_28276 = v_28274 | v_28275;
assign v_28278 = v_28160 | v_28277;
assign v_28281 = v_28279 | v_28280;
assign v_28283 = v_28157 | v_28282;
assign v_28286 = v_28284 | v_28285;
assign v_28288 = v_28154 | v_28287;
assign v_28291 = v_28289 | v_28290;
assign v_28293 = v_28151 | v_28292;
assign v_28296 = v_28294 | v_28295;
assign v_28298 = v_28148 | v_28297;
assign v_28301 = v_28299 | v_28300;
assign v_28303 = v_28145 | v_28302;
assign v_28306 = v_28304 | v_28305;
assign v_28308 = v_28142 | v_28307;
assign v_28311 = v_28309 | v_28310;
assign v_28313 = v_28139 | v_28312;
assign v_28316 = v_28314 | v_28315;
assign v_28318 = v_28136 | v_28317;
assign v_28321 = v_28319 | v_28320;
assign v_28323 = v_28133 | v_28322;
assign v_28326 = v_28324 | v_28325;
assign v_28328 = v_28130 | v_28327;
assign v_28331 = v_28329 | v_28330;
assign v_28333 = v_28127 | v_28332;
assign v_28336 = v_28334 | v_28335;
assign v_28338 = v_28124 | v_28337;
assign v_28341 = v_28339 | v_28340;
assign v_28343 = v_28121 | v_28342;
assign v_28346 = v_28344 | v_28345;
assign v_28348 = v_28118 | v_28347;
assign v_28351 = v_28349 | v_28350;
assign v_28353 = v_28115 | v_28352;
assign v_28356 = v_28114 | v_28355;
assign v_28410 = v_28407 | v_28409;
assign v_28412 = v_28406 | v_28411;
assign v_28414 = v_28404 | v_28413;
assign v_28416 = v_28411 | v_28415;
assign v_28418 = v_28403 | v_28417;
assign v_28420 = v_28401 | v_28419;
assign v_28422 = v_28417 | v_28421;
assign v_28424 = v_28400 | v_28423;
assign v_28426 = v_28398 | v_28425;
assign v_28428 = v_28423 | v_28427;
assign v_28430 = v_28397 | v_28429;
assign v_28432 = v_28395 | v_28431;
assign v_28434 = v_28429 | v_28433;
assign v_28436 = v_28394 | v_28435;
assign v_28438 = v_28392 | v_28437;
assign v_28440 = v_28435 | v_28439;
assign v_28442 = v_28391 | v_28441;
assign v_28444 = v_28389 | v_28443;
assign v_28446 = v_28441 | v_28445;
assign v_28448 = v_28388 | v_28447;
assign v_28450 = v_28386 | v_28449;
assign v_28452 = v_28447 | v_28451;
assign v_28454 = v_28385 | v_28453;
assign v_28456 = v_28383 | v_28455;
assign v_28458 = v_28453 | v_28457;
assign v_28460 = v_28382 | v_28459;
assign v_28462 = v_28380 | v_28461;
assign v_28464 = v_28459 | v_28463;
assign v_28466 = v_28379 | v_28465;
assign v_28468 = v_28377 | v_28467;
assign v_28470 = v_28465 | v_28469;
assign v_28472 = v_28376 | v_28471;
assign v_28474 = v_28374 | v_28473;
assign v_28476 = v_28471 | v_28475;
assign v_28478 = v_28373 | v_28477;
assign v_28480 = v_28371 | v_28479;
assign v_28482 = v_28477 | v_28481;
assign v_28484 = v_28370 | v_28483;
assign v_28486 = v_28368 | v_28485;
assign v_28488 = v_28483 | v_28487;
assign v_28490 = v_28367 | v_28489;
assign v_28492 = v_28365 | v_28491;
assign v_28494 = v_28489 | v_28493;
assign v_28496 = v_28364 | v_28495;
assign v_28498 = v_28362 | v_28497;
assign v_28500 = v_28495 | v_28499;
assign v_28502 = v_28361 | v_28501;
assign v_28504 = v_28359 | v_28503;
assign v_28506 = v_28501 | v_28505;
assign v_28509 = ~v_28358 | v_28508;
assign v_28516 = v_28406 | v_28515;
assign v_28519 = v_28517 | v_28518;
assign v_28521 = v_28403 | v_28520;
assign v_28524 = v_28522 | v_28523;
assign v_28526 = v_28400 | v_28525;
assign v_28529 = v_28527 | v_28528;
assign v_28531 = v_28397 | v_28530;
assign v_28534 = v_28532 | v_28533;
assign v_28536 = v_28394 | v_28535;
assign v_28539 = v_28537 | v_28538;
assign v_28541 = v_28391 | v_28540;
assign v_28544 = v_28542 | v_28543;
assign v_28546 = v_28388 | v_28545;
assign v_28549 = v_28547 | v_28548;
assign v_28551 = v_28385 | v_28550;
assign v_28554 = v_28552 | v_28553;
assign v_28556 = v_28382 | v_28555;
assign v_28559 = v_28557 | v_28558;
assign v_28561 = v_28379 | v_28560;
assign v_28564 = v_28562 | v_28563;
assign v_28566 = v_28376 | v_28565;
assign v_28569 = v_28567 | v_28568;
assign v_28571 = v_28373 | v_28570;
assign v_28574 = v_28572 | v_28573;
assign v_28576 = v_28370 | v_28575;
assign v_28579 = v_28577 | v_28578;
assign v_28581 = v_28367 | v_28580;
assign v_28584 = v_28582 | v_28583;
assign v_28586 = v_28364 | v_28585;
assign v_28589 = v_28587 | v_28588;
assign v_28591 = v_28361 | v_28590;
assign v_28594 = v_28592 | v_28593;
assign v_28596 = v_28358 | v_28595;
assign v_28599 = v_28357 | v_28598;
assign v_28653 = v_28650 | v_28652;
assign v_28655 = v_28649 | v_28654;
assign v_28657 = v_28647 | v_28656;
assign v_28659 = v_28654 | v_28658;
assign v_28661 = v_28646 | v_28660;
assign v_28663 = v_28644 | v_28662;
assign v_28665 = v_28660 | v_28664;
assign v_28667 = v_28643 | v_28666;
assign v_28669 = v_28641 | v_28668;
assign v_28671 = v_28666 | v_28670;
assign v_28673 = v_28640 | v_28672;
assign v_28675 = v_28638 | v_28674;
assign v_28677 = v_28672 | v_28676;
assign v_28679 = v_28637 | v_28678;
assign v_28681 = v_28635 | v_28680;
assign v_28683 = v_28678 | v_28682;
assign v_28685 = v_28634 | v_28684;
assign v_28687 = v_28632 | v_28686;
assign v_28689 = v_28684 | v_28688;
assign v_28691 = v_28631 | v_28690;
assign v_28693 = v_28629 | v_28692;
assign v_28695 = v_28690 | v_28694;
assign v_28697 = v_28628 | v_28696;
assign v_28699 = v_28626 | v_28698;
assign v_28701 = v_28696 | v_28700;
assign v_28703 = v_28625 | v_28702;
assign v_28705 = v_28623 | v_28704;
assign v_28707 = v_28702 | v_28706;
assign v_28709 = v_28622 | v_28708;
assign v_28711 = v_28620 | v_28710;
assign v_28713 = v_28708 | v_28712;
assign v_28715 = v_28619 | v_28714;
assign v_28717 = v_28617 | v_28716;
assign v_28719 = v_28714 | v_28718;
assign v_28721 = v_28616 | v_28720;
assign v_28723 = v_28614 | v_28722;
assign v_28725 = v_28720 | v_28724;
assign v_28727 = v_28613 | v_28726;
assign v_28729 = v_28611 | v_28728;
assign v_28731 = v_28726 | v_28730;
assign v_28733 = v_28610 | v_28732;
assign v_28735 = v_28608 | v_28734;
assign v_28737 = v_28732 | v_28736;
assign v_28739 = v_28607 | v_28738;
assign v_28741 = v_28605 | v_28740;
assign v_28743 = v_28738 | v_28742;
assign v_28745 = v_28604 | v_28744;
assign v_28747 = v_28602 | v_28746;
assign v_28749 = v_28744 | v_28748;
assign v_28752 = ~v_28601 | v_28751;
assign v_28759 = v_28649 | v_28758;
assign v_28762 = v_28760 | v_28761;
assign v_28764 = v_28646 | v_28763;
assign v_28767 = v_28765 | v_28766;
assign v_28769 = v_28643 | v_28768;
assign v_28772 = v_28770 | v_28771;
assign v_28774 = v_28640 | v_28773;
assign v_28777 = v_28775 | v_28776;
assign v_28779 = v_28637 | v_28778;
assign v_28782 = v_28780 | v_28781;
assign v_28784 = v_28634 | v_28783;
assign v_28787 = v_28785 | v_28786;
assign v_28789 = v_28631 | v_28788;
assign v_28792 = v_28790 | v_28791;
assign v_28794 = v_28628 | v_28793;
assign v_28797 = v_28795 | v_28796;
assign v_28799 = v_28625 | v_28798;
assign v_28802 = v_28800 | v_28801;
assign v_28804 = v_28622 | v_28803;
assign v_28807 = v_28805 | v_28806;
assign v_28809 = v_28619 | v_28808;
assign v_28812 = v_28810 | v_28811;
assign v_28814 = v_28616 | v_28813;
assign v_28817 = v_28815 | v_28816;
assign v_28819 = v_28613 | v_28818;
assign v_28822 = v_28820 | v_28821;
assign v_28824 = v_28610 | v_28823;
assign v_28827 = v_28825 | v_28826;
assign v_28829 = v_28607 | v_28828;
assign v_28832 = v_28830 | v_28831;
assign v_28834 = v_28604 | v_28833;
assign v_28837 = v_28835 | v_28836;
assign v_28839 = v_28601 | v_28838;
assign v_28842 = v_28600 | v_28841;
assign v_28896 = v_28893 | v_28895;
assign v_28898 = v_28892 | v_28897;
assign v_28900 = v_28890 | v_28899;
assign v_28902 = v_28897 | v_28901;
assign v_28904 = v_28889 | v_28903;
assign v_28906 = v_28887 | v_28905;
assign v_28908 = v_28903 | v_28907;
assign v_28910 = v_28886 | v_28909;
assign v_28912 = v_28884 | v_28911;
assign v_28914 = v_28909 | v_28913;
assign v_28916 = v_28883 | v_28915;
assign v_28918 = v_28881 | v_28917;
assign v_28920 = v_28915 | v_28919;
assign v_28922 = v_28880 | v_28921;
assign v_28924 = v_28878 | v_28923;
assign v_28926 = v_28921 | v_28925;
assign v_28928 = v_28877 | v_28927;
assign v_28930 = v_28875 | v_28929;
assign v_28932 = v_28927 | v_28931;
assign v_28934 = v_28874 | v_28933;
assign v_28936 = v_28872 | v_28935;
assign v_28938 = v_28933 | v_28937;
assign v_28940 = v_28871 | v_28939;
assign v_28942 = v_28869 | v_28941;
assign v_28944 = v_28939 | v_28943;
assign v_28946 = v_28868 | v_28945;
assign v_28948 = v_28866 | v_28947;
assign v_28950 = v_28945 | v_28949;
assign v_28952 = v_28865 | v_28951;
assign v_28954 = v_28863 | v_28953;
assign v_28956 = v_28951 | v_28955;
assign v_28958 = v_28862 | v_28957;
assign v_28960 = v_28860 | v_28959;
assign v_28962 = v_28957 | v_28961;
assign v_28964 = v_28859 | v_28963;
assign v_28966 = v_28857 | v_28965;
assign v_28968 = v_28963 | v_28967;
assign v_28970 = v_28856 | v_28969;
assign v_28972 = v_28854 | v_28971;
assign v_28974 = v_28969 | v_28973;
assign v_28976 = v_28853 | v_28975;
assign v_28978 = v_28851 | v_28977;
assign v_28980 = v_28975 | v_28979;
assign v_28982 = v_28850 | v_28981;
assign v_28984 = v_28848 | v_28983;
assign v_28986 = v_28981 | v_28985;
assign v_28988 = v_28847 | v_28987;
assign v_28990 = v_28845 | v_28989;
assign v_28992 = v_28987 | v_28991;
assign v_28995 = ~v_28844 | v_28994;
assign v_29002 = v_28892 | v_29001;
assign v_29005 = v_29003 | v_29004;
assign v_29007 = v_28889 | v_29006;
assign v_29010 = v_29008 | v_29009;
assign v_29012 = v_28886 | v_29011;
assign v_29015 = v_29013 | v_29014;
assign v_29017 = v_28883 | v_29016;
assign v_29020 = v_29018 | v_29019;
assign v_29022 = v_28880 | v_29021;
assign v_29025 = v_29023 | v_29024;
assign v_29027 = v_28877 | v_29026;
assign v_29030 = v_29028 | v_29029;
assign v_29032 = v_28874 | v_29031;
assign v_29035 = v_29033 | v_29034;
assign v_29037 = v_28871 | v_29036;
assign v_29040 = v_29038 | v_29039;
assign v_29042 = v_28868 | v_29041;
assign v_29045 = v_29043 | v_29044;
assign v_29047 = v_28865 | v_29046;
assign v_29050 = v_29048 | v_29049;
assign v_29052 = v_28862 | v_29051;
assign v_29055 = v_29053 | v_29054;
assign v_29057 = v_28859 | v_29056;
assign v_29060 = v_29058 | v_29059;
assign v_29062 = v_28856 | v_29061;
assign v_29065 = v_29063 | v_29064;
assign v_29067 = v_28853 | v_29066;
assign v_29070 = v_29068 | v_29069;
assign v_29072 = v_28850 | v_29071;
assign v_29075 = v_29073 | v_29074;
assign v_29077 = v_28847 | v_29076;
assign v_29080 = v_29078 | v_29079;
assign v_29082 = v_28844 | v_29081;
assign v_29085 = v_28843 | v_29084;
assign v_29138 = v_29135 | v_29137;
assign v_29140 = v_29134 | v_29139;
assign v_29142 = v_29132 | v_29141;
assign v_29144 = v_29139 | v_29143;
assign v_29146 = v_29131 | v_29145;
assign v_29148 = v_29129 | v_29147;
assign v_29150 = v_29145 | v_29149;
assign v_29152 = v_29128 | v_29151;
assign v_29154 = v_29126 | v_29153;
assign v_29156 = v_29151 | v_29155;
assign v_29158 = v_29125 | v_29157;
assign v_29160 = v_29123 | v_29159;
assign v_29162 = v_29157 | v_29161;
assign v_29164 = v_29122 | v_29163;
assign v_29166 = v_29120 | v_29165;
assign v_29168 = v_29163 | v_29167;
assign v_29170 = v_29119 | v_29169;
assign v_29172 = v_29117 | v_29171;
assign v_29174 = v_29169 | v_29173;
assign v_29176 = v_29116 | v_29175;
assign v_29178 = v_29114 | v_29177;
assign v_29180 = v_29175 | v_29179;
assign v_29182 = v_29113 | v_29181;
assign v_29184 = v_29111 | v_29183;
assign v_29186 = v_29181 | v_29185;
assign v_29188 = v_29110 | v_29187;
assign v_29190 = v_29108 | v_29189;
assign v_29192 = v_29187 | v_29191;
assign v_29194 = v_29107 | v_29193;
assign v_29196 = v_29105 | v_29195;
assign v_29198 = v_29193 | v_29197;
assign v_29200 = v_29104 | v_29199;
assign v_29202 = v_29102 | v_29201;
assign v_29204 = v_29199 | v_29203;
assign v_29206 = v_29101 | v_29205;
assign v_29208 = v_29099 | v_29207;
assign v_29210 = v_29205 | v_29209;
assign v_29212 = v_29098 | v_29211;
assign v_29214 = v_29096 | v_29213;
assign v_29216 = v_29211 | v_29215;
assign v_29218 = v_29095 | v_29217;
assign v_29220 = v_29093 | v_29219;
assign v_29222 = v_29217 | v_29221;
assign v_29224 = v_29092 | v_29223;
assign v_29226 = v_29090 | v_29225;
assign v_29228 = v_29223 | v_29227;
assign v_29230 = v_29089 | v_29229;
assign v_29232 = v_29087 | v_29231;
assign v_29234 = v_29229 | v_29233;
assign v_29238 = v_29235 | v_29237;
assign v_29245 = v_29134 | v_29244;
assign v_29248 = v_29246 | v_29247;
assign v_29250 = v_29131 | v_29249;
assign v_29253 = v_29251 | v_29252;
assign v_29255 = v_29128 | v_29254;
assign v_29258 = v_29256 | v_29257;
assign v_29260 = v_29125 | v_29259;
assign v_29263 = v_29261 | v_29262;
assign v_29265 = v_29122 | v_29264;
assign v_29268 = v_29266 | v_29267;
assign v_29270 = v_29119 | v_29269;
assign v_29273 = v_29271 | v_29272;
assign v_29275 = v_29116 | v_29274;
assign v_29278 = v_29276 | v_29277;
assign v_29280 = v_29113 | v_29279;
assign v_29283 = v_29281 | v_29282;
assign v_29285 = v_29110 | v_29284;
assign v_29288 = v_29286 | v_29287;
assign v_29290 = v_29107 | v_29289;
assign v_29293 = v_29291 | v_29292;
assign v_29295 = v_29104 | v_29294;
assign v_29298 = v_29296 | v_29297;
assign v_29300 = v_29101 | v_29299;
assign v_29303 = v_29301 | v_29302;
assign v_29305 = v_29098 | v_29304;
assign v_29308 = v_29306 | v_29307;
assign v_29310 = v_29095 | v_29309;
assign v_29313 = v_29311 | v_29312;
assign v_29315 = v_29092 | v_29314;
assign v_29318 = v_29316 | v_29317;
assign v_29320 = v_29089 | v_29319;
assign v_29323 = v_29321 | v_29322;
assign v_29325 = v_29323 | v_29324;
assign v_29328 = v_29086 | v_29327;
assign v_29399 = v_29396 | v_29398;
assign v_29401 = v_29394 | v_29400;
assign v_29403 = v_29392 | v_29402;
assign v_29405 = v_29400 | v_29404;
assign v_29407 = v_29390 | v_29406;
assign v_29409 = v_29388 | v_29408;
assign v_29411 = v_29406 | v_29410;
assign v_29413 = v_29386 | v_29412;
assign v_29415 = v_29384 | v_29414;
assign v_29417 = v_29412 | v_29416;
assign v_29419 = v_29382 | v_29418;
assign v_29421 = v_29380 | v_29420;
assign v_29423 = v_29418 | v_29422;
assign v_29425 = v_29378 | v_29424;
assign v_29427 = v_29376 | v_29426;
assign v_29429 = v_29424 | v_29428;
assign v_29431 = v_29374 | v_29430;
assign v_29433 = v_29372 | v_29432;
assign v_29435 = v_29430 | v_29434;
assign v_29437 = v_29370 | v_29436;
assign v_29439 = v_29368 | v_29438;
assign v_29441 = v_29436 | v_29440;
assign v_29443 = v_29366 | v_29442;
assign v_29445 = v_29364 | v_29444;
assign v_29447 = v_29442 | v_29446;
assign v_29449 = v_29362 | v_29448;
assign v_29451 = v_29360 | v_29450;
assign v_29453 = v_29448 | v_29452;
assign v_29455 = v_29358 | v_29454;
assign v_29457 = v_29356 | v_29456;
assign v_29459 = v_29454 | v_29458;
assign v_29461 = v_29354 | v_29460;
assign v_29463 = v_29352 | v_29462;
assign v_29465 = v_29460 | v_29464;
assign v_29467 = v_29350 | v_29466;
assign v_29469 = v_29348 | v_29468;
assign v_29471 = v_29466 | v_29470;
assign v_29473 = v_29346 | v_29472;
assign v_29475 = v_29343 | v_29474;
assign v_29477 = v_29472 | v_29476;
assign v_29479 = v_29342 | v_29478;
assign v_29481 = v_29339 | v_29480;
assign v_29483 = v_29478 | v_29482;
assign v_29485 = v_29338 | v_29484;
assign v_29487 = v_29335 | v_29486;
assign v_29489 = v_29484 | v_29488;
assign v_29491 = v_29334 | v_29490;
assign v_29493 = v_29331 | v_29492;
assign v_29495 = v_29490 | v_29494;
assign v_29498 = ~v_29330 | v_29497;
assign v_29505 = v_29394 | v_29504;
assign v_29508 = v_29506 | v_29507;
assign v_29510 = v_29390 | v_29509;
assign v_29513 = v_29511 | v_29512;
assign v_29515 = v_29386 | v_29514;
assign v_29518 = v_29516 | v_29517;
assign v_29520 = v_29382 | v_29519;
assign v_29523 = v_29521 | v_29522;
assign v_29525 = v_29378 | v_29524;
assign v_29528 = v_29526 | v_29527;
assign v_29530 = v_29374 | v_29529;
assign v_29533 = v_29531 | v_29532;
assign v_29535 = v_29370 | v_29534;
assign v_29538 = v_29536 | v_29537;
assign v_29540 = v_29366 | v_29539;
assign v_29543 = v_29541 | v_29542;
assign v_29545 = v_29362 | v_29544;
assign v_29548 = v_29546 | v_29547;
assign v_29550 = v_29358 | v_29549;
assign v_29553 = v_29551 | v_29552;
assign v_29555 = v_29354 | v_29554;
assign v_29558 = v_29556 | v_29557;
assign v_29560 = v_29350 | v_29559;
assign v_29563 = v_29561 | v_29562;
assign v_29565 = v_29346 | v_29564;
assign v_29568 = v_29566 | v_29567;
assign v_29570 = v_29342 | v_29569;
assign v_29573 = v_29571 | v_29572;
assign v_29575 = v_29338 | v_29574;
assign v_29578 = v_29576 | v_29577;
assign v_29580 = v_29334 | v_29579;
assign v_29583 = v_29581 | v_29582;
assign v_29585 = v_29330 | v_29584;
assign v_29588 = v_29329 | v_29587;
assign v_29642 = v_29639 | v_29641;
assign v_29644 = v_29638 | v_29643;
assign v_29646 = v_29636 | v_29645;
assign v_29648 = v_29643 | v_29647;
assign v_29650 = v_29635 | v_29649;
assign v_29652 = v_29633 | v_29651;
assign v_29654 = v_29649 | v_29653;
assign v_29656 = v_29632 | v_29655;
assign v_29658 = v_29630 | v_29657;
assign v_29660 = v_29655 | v_29659;
assign v_29662 = v_29629 | v_29661;
assign v_29664 = v_29627 | v_29663;
assign v_29666 = v_29661 | v_29665;
assign v_29668 = v_29626 | v_29667;
assign v_29670 = v_29624 | v_29669;
assign v_29672 = v_29667 | v_29671;
assign v_29674 = v_29623 | v_29673;
assign v_29676 = v_29621 | v_29675;
assign v_29678 = v_29673 | v_29677;
assign v_29680 = v_29620 | v_29679;
assign v_29682 = v_29618 | v_29681;
assign v_29684 = v_29679 | v_29683;
assign v_29686 = v_29617 | v_29685;
assign v_29688 = v_29615 | v_29687;
assign v_29690 = v_29685 | v_29689;
assign v_29692 = v_29614 | v_29691;
assign v_29694 = v_29612 | v_29693;
assign v_29696 = v_29691 | v_29695;
assign v_29698 = v_29611 | v_29697;
assign v_29700 = v_29609 | v_29699;
assign v_29702 = v_29697 | v_29701;
assign v_29704 = v_29608 | v_29703;
assign v_29706 = v_29606 | v_29705;
assign v_29708 = v_29703 | v_29707;
assign v_29710 = v_29605 | v_29709;
assign v_29712 = v_29603 | v_29711;
assign v_29714 = v_29709 | v_29713;
assign v_29716 = v_29602 | v_29715;
assign v_29718 = v_29600 | v_29717;
assign v_29720 = v_29715 | v_29719;
assign v_29722 = v_29599 | v_29721;
assign v_29724 = v_29597 | v_29723;
assign v_29726 = v_29721 | v_29725;
assign v_29728 = v_29596 | v_29727;
assign v_29730 = v_29594 | v_29729;
assign v_29732 = v_29727 | v_29731;
assign v_29734 = v_29593 | v_29733;
assign v_29736 = v_29591 | v_29735;
assign v_29738 = v_29733 | v_29737;
assign v_29741 = ~v_29590 | v_29740;
assign v_29748 = v_29638 | v_29747;
assign v_29751 = v_29749 | v_29750;
assign v_29753 = v_29635 | v_29752;
assign v_29756 = v_29754 | v_29755;
assign v_29758 = v_29632 | v_29757;
assign v_29761 = v_29759 | v_29760;
assign v_29763 = v_29629 | v_29762;
assign v_29766 = v_29764 | v_29765;
assign v_29768 = v_29626 | v_29767;
assign v_29771 = v_29769 | v_29770;
assign v_29773 = v_29623 | v_29772;
assign v_29776 = v_29774 | v_29775;
assign v_29778 = v_29620 | v_29777;
assign v_29781 = v_29779 | v_29780;
assign v_29783 = v_29617 | v_29782;
assign v_29786 = v_29784 | v_29785;
assign v_29788 = v_29614 | v_29787;
assign v_29791 = v_29789 | v_29790;
assign v_29793 = v_29611 | v_29792;
assign v_29796 = v_29794 | v_29795;
assign v_29798 = v_29608 | v_29797;
assign v_29801 = v_29799 | v_29800;
assign v_29803 = v_29605 | v_29802;
assign v_29806 = v_29804 | v_29805;
assign v_29808 = v_29602 | v_29807;
assign v_29811 = v_29809 | v_29810;
assign v_29813 = v_29599 | v_29812;
assign v_29816 = v_29814 | v_29815;
assign v_29818 = v_29596 | v_29817;
assign v_29821 = v_29819 | v_29820;
assign v_29823 = v_29593 | v_29822;
assign v_29826 = v_29824 | v_29825;
assign v_29828 = v_29590 | v_29827;
assign v_29831 = v_29589 | v_29830;
assign v_29885 = v_29882 | v_29884;
assign v_29887 = v_29881 | v_29886;
assign v_29889 = v_29879 | v_29888;
assign v_29891 = v_29886 | v_29890;
assign v_29893 = v_29878 | v_29892;
assign v_29895 = v_29876 | v_29894;
assign v_29897 = v_29892 | v_29896;
assign v_29899 = v_29875 | v_29898;
assign v_29901 = v_29873 | v_29900;
assign v_29903 = v_29898 | v_29902;
assign v_29905 = v_29872 | v_29904;
assign v_29907 = v_29870 | v_29906;
assign v_29909 = v_29904 | v_29908;
assign v_29911 = v_29869 | v_29910;
assign v_29913 = v_29867 | v_29912;
assign v_29915 = v_29910 | v_29914;
assign v_29917 = v_29866 | v_29916;
assign v_29919 = v_29864 | v_29918;
assign v_29921 = v_29916 | v_29920;
assign v_29923 = v_29863 | v_29922;
assign v_29925 = v_29861 | v_29924;
assign v_29927 = v_29922 | v_29926;
assign v_29929 = v_29860 | v_29928;
assign v_29931 = v_29858 | v_29930;
assign v_29933 = v_29928 | v_29932;
assign v_29935 = v_29857 | v_29934;
assign v_29937 = v_29855 | v_29936;
assign v_29939 = v_29934 | v_29938;
assign v_29941 = v_29854 | v_29940;
assign v_29943 = v_29852 | v_29942;
assign v_29945 = v_29940 | v_29944;
assign v_29947 = v_29851 | v_29946;
assign v_29949 = v_29849 | v_29948;
assign v_29951 = v_29946 | v_29950;
assign v_29953 = v_29848 | v_29952;
assign v_29955 = v_29846 | v_29954;
assign v_29957 = v_29952 | v_29956;
assign v_29959 = v_29845 | v_29958;
assign v_29961 = v_29843 | v_29960;
assign v_29963 = v_29958 | v_29962;
assign v_29965 = v_29842 | v_29964;
assign v_29967 = v_29840 | v_29966;
assign v_29969 = v_29964 | v_29968;
assign v_29971 = v_29839 | v_29970;
assign v_29973 = v_29837 | v_29972;
assign v_29975 = v_29970 | v_29974;
assign v_29977 = v_29836 | v_29976;
assign v_29979 = v_29834 | v_29978;
assign v_29981 = v_29976 | v_29980;
assign v_29984 = ~v_29833 | v_29983;
assign v_29991 = v_29881 | v_29990;
assign v_29994 = v_29992 | v_29993;
assign v_29996 = v_29878 | v_29995;
assign v_29999 = v_29997 | v_29998;
assign v_30001 = v_29875 | v_30000;
assign v_30004 = v_30002 | v_30003;
assign v_30006 = v_29872 | v_30005;
assign v_30009 = v_30007 | v_30008;
assign v_30011 = v_29869 | v_30010;
assign v_30014 = v_30012 | v_30013;
assign v_30016 = v_29866 | v_30015;
assign v_30019 = v_30017 | v_30018;
assign v_30021 = v_29863 | v_30020;
assign v_30024 = v_30022 | v_30023;
assign v_30026 = v_29860 | v_30025;
assign v_30029 = v_30027 | v_30028;
assign v_30031 = v_29857 | v_30030;
assign v_30034 = v_30032 | v_30033;
assign v_30036 = v_29854 | v_30035;
assign v_30039 = v_30037 | v_30038;
assign v_30041 = v_29851 | v_30040;
assign v_30044 = v_30042 | v_30043;
assign v_30046 = v_29848 | v_30045;
assign v_30049 = v_30047 | v_30048;
assign v_30051 = v_29845 | v_30050;
assign v_30054 = v_30052 | v_30053;
assign v_30056 = v_29842 | v_30055;
assign v_30059 = v_30057 | v_30058;
assign v_30061 = v_29839 | v_30060;
assign v_30064 = v_30062 | v_30063;
assign v_30066 = v_29836 | v_30065;
assign v_30069 = v_30067 | v_30068;
assign v_30071 = v_29833 | v_30070;
assign v_30074 = v_29832 | v_30073;
assign v_30128 = v_30125 | v_30127;
assign v_30130 = v_30124 | v_30129;
assign v_30132 = v_30122 | v_30131;
assign v_30134 = v_30129 | v_30133;
assign v_30136 = v_30121 | v_30135;
assign v_30138 = v_30119 | v_30137;
assign v_30140 = v_30135 | v_30139;
assign v_30142 = v_30118 | v_30141;
assign v_30144 = v_30116 | v_30143;
assign v_30146 = v_30141 | v_30145;
assign v_30148 = v_30115 | v_30147;
assign v_30150 = v_30113 | v_30149;
assign v_30152 = v_30147 | v_30151;
assign v_30154 = v_30112 | v_30153;
assign v_30156 = v_30110 | v_30155;
assign v_30158 = v_30153 | v_30157;
assign v_30160 = v_30109 | v_30159;
assign v_30162 = v_30107 | v_30161;
assign v_30164 = v_30159 | v_30163;
assign v_30166 = v_30106 | v_30165;
assign v_30168 = v_30104 | v_30167;
assign v_30170 = v_30165 | v_30169;
assign v_30172 = v_30103 | v_30171;
assign v_30174 = v_30101 | v_30173;
assign v_30176 = v_30171 | v_30175;
assign v_30178 = v_30100 | v_30177;
assign v_30180 = v_30098 | v_30179;
assign v_30182 = v_30177 | v_30181;
assign v_30184 = v_30097 | v_30183;
assign v_30186 = v_30095 | v_30185;
assign v_30188 = v_30183 | v_30187;
assign v_30190 = v_30094 | v_30189;
assign v_30192 = v_30092 | v_30191;
assign v_30194 = v_30189 | v_30193;
assign v_30196 = v_30091 | v_30195;
assign v_30198 = v_30089 | v_30197;
assign v_30200 = v_30195 | v_30199;
assign v_30202 = v_30088 | v_30201;
assign v_30204 = v_30086 | v_30203;
assign v_30206 = v_30201 | v_30205;
assign v_30208 = v_30085 | v_30207;
assign v_30210 = v_30083 | v_30209;
assign v_30212 = v_30207 | v_30211;
assign v_30214 = v_30082 | v_30213;
assign v_30216 = v_30080 | v_30215;
assign v_30218 = v_30213 | v_30217;
assign v_30220 = v_30079 | v_30219;
assign v_30222 = v_30077 | v_30221;
assign v_30224 = v_30219 | v_30223;
assign v_30227 = ~v_30076 | v_30226;
assign v_30234 = v_30124 | v_30233;
assign v_30237 = v_30235 | v_30236;
assign v_30239 = v_30121 | v_30238;
assign v_30242 = v_30240 | v_30241;
assign v_30244 = v_30118 | v_30243;
assign v_30247 = v_30245 | v_30246;
assign v_30249 = v_30115 | v_30248;
assign v_30252 = v_30250 | v_30251;
assign v_30254 = v_30112 | v_30253;
assign v_30257 = v_30255 | v_30256;
assign v_30259 = v_30109 | v_30258;
assign v_30262 = v_30260 | v_30261;
assign v_30264 = v_30106 | v_30263;
assign v_30267 = v_30265 | v_30266;
assign v_30269 = v_30103 | v_30268;
assign v_30272 = v_30270 | v_30271;
assign v_30274 = v_30100 | v_30273;
assign v_30277 = v_30275 | v_30276;
assign v_30279 = v_30097 | v_30278;
assign v_30282 = v_30280 | v_30281;
assign v_30284 = v_30094 | v_30283;
assign v_30287 = v_30285 | v_30286;
assign v_30289 = v_30091 | v_30288;
assign v_30292 = v_30290 | v_30291;
assign v_30294 = v_30088 | v_30293;
assign v_30297 = v_30295 | v_30296;
assign v_30299 = v_30085 | v_30298;
assign v_30302 = v_30300 | v_30301;
assign v_30304 = v_30082 | v_30303;
assign v_30307 = v_30305 | v_30306;
assign v_30309 = v_30079 | v_30308;
assign v_30312 = v_30310 | v_30311;
assign v_30314 = v_30076 | v_30313;
assign v_30317 = v_30075 | v_30316;
assign v_30371 = v_30368 | v_30370;
assign v_30373 = v_30367 | v_30372;
assign v_30375 = v_30365 | v_30374;
assign v_30377 = v_30372 | v_30376;
assign v_30379 = v_30364 | v_30378;
assign v_30381 = v_30362 | v_30380;
assign v_30383 = v_30378 | v_30382;
assign v_30385 = v_30361 | v_30384;
assign v_30387 = v_30359 | v_30386;
assign v_30389 = v_30384 | v_30388;
assign v_30391 = v_30358 | v_30390;
assign v_30393 = v_30356 | v_30392;
assign v_30395 = v_30390 | v_30394;
assign v_30397 = v_30355 | v_30396;
assign v_30399 = v_30353 | v_30398;
assign v_30401 = v_30396 | v_30400;
assign v_30403 = v_30352 | v_30402;
assign v_30405 = v_30350 | v_30404;
assign v_30407 = v_30402 | v_30406;
assign v_30409 = v_30349 | v_30408;
assign v_30411 = v_30347 | v_30410;
assign v_30413 = v_30408 | v_30412;
assign v_30415 = v_30346 | v_30414;
assign v_30417 = v_30344 | v_30416;
assign v_30419 = v_30414 | v_30418;
assign v_30421 = v_30343 | v_30420;
assign v_30423 = v_30341 | v_30422;
assign v_30425 = v_30420 | v_30424;
assign v_30427 = v_30340 | v_30426;
assign v_30429 = v_30338 | v_30428;
assign v_30431 = v_30426 | v_30430;
assign v_30433 = v_30337 | v_30432;
assign v_30435 = v_30335 | v_30434;
assign v_30437 = v_30432 | v_30436;
assign v_30439 = v_30334 | v_30438;
assign v_30441 = v_30332 | v_30440;
assign v_30443 = v_30438 | v_30442;
assign v_30445 = v_30331 | v_30444;
assign v_30447 = v_30329 | v_30446;
assign v_30449 = v_30444 | v_30448;
assign v_30451 = v_30328 | v_30450;
assign v_30453 = v_30326 | v_30452;
assign v_30455 = v_30450 | v_30454;
assign v_30457 = v_30325 | v_30456;
assign v_30459 = v_30323 | v_30458;
assign v_30461 = v_30456 | v_30460;
assign v_30463 = v_30322 | v_30462;
assign v_30465 = v_30320 | v_30464;
assign v_30467 = v_30462 | v_30466;
assign v_30470 = ~v_30319 | v_30469;
assign v_30477 = v_30367 | v_30476;
assign v_30480 = v_30478 | v_30479;
assign v_30482 = v_30364 | v_30481;
assign v_30485 = v_30483 | v_30484;
assign v_30487 = v_30361 | v_30486;
assign v_30490 = v_30488 | v_30489;
assign v_30492 = v_30358 | v_30491;
assign v_30495 = v_30493 | v_30494;
assign v_30497 = v_30355 | v_30496;
assign v_30500 = v_30498 | v_30499;
assign v_30502 = v_30352 | v_30501;
assign v_30505 = v_30503 | v_30504;
assign v_30507 = v_30349 | v_30506;
assign v_30510 = v_30508 | v_30509;
assign v_30512 = v_30346 | v_30511;
assign v_30515 = v_30513 | v_30514;
assign v_30517 = v_30343 | v_30516;
assign v_30520 = v_30518 | v_30519;
assign v_30522 = v_30340 | v_30521;
assign v_30525 = v_30523 | v_30524;
assign v_30527 = v_30337 | v_30526;
assign v_30530 = v_30528 | v_30529;
assign v_30532 = v_30334 | v_30531;
assign v_30535 = v_30533 | v_30534;
assign v_30537 = v_30331 | v_30536;
assign v_30540 = v_30538 | v_30539;
assign v_30542 = v_30328 | v_30541;
assign v_30545 = v_30543 | v_30544;
assign v_30547 = v_30325 | v_30546;
assign v_30550 = v_30548 | v_30549;
assign v_30552 = v_30322 | v_30551;
assign v_30555 = v_30553 | v_30554;
assign v_30557 = v_30319 | v_30556;
assign v_30560 = v_30318 | v_30559;
assign v_30614 = v_30611 | v_30613;
assign v_30616 = v_30610 | v_30615;
assign v_30618 = v_30608 | v_30617;
assign v_30620 = v_30615 | v_30619;
assign v_30622 = v_30607 | v_30621;
assign v_30624 = v_30605 | v_30623;
assign v_30626 = v_30621 | v_30625;
assign v_30628 = v_30604 | v_30627;
assign v_30630 = v_30602 | v_30629;
assign v_30632 = v_30627 | v_30631;
assign v_30634 = v_30601 | v_30633;
assign v_30636 = v_30599 | v_30635;
assign v_30638 = v_30633 | v_30637;
assign v_30640 = v_30598 | v_30639;
assign v_30642 = v_30596 | v_30641;
assign v_30644 = v_30639 | v_30643;
assign v_30646 = v_30595 | v_30645;
assign v_30648 = v_30593 | v_30647;
assign v_30650 = v_30645 | v_30649;
assign v_30652 = v_30592 | v_30651;
assign v_30654 = v_30590 | v_30653;
assign v_30656 = v_30651 | v_30655;
assign v_30658 = v_30589 | v_30657;
assign v_30660 = v_30587 | v_30659;
assign v_30662 = v_30657 | v_30661;
assign v_30664 = v_30586 | v_30663;
assign v_30666 = v_30584 | v_30665;
assign v_30668 = v_30663 | v_30667;
assign v_30670 = v_30583 | v_30669;
assign v_30672 = v_30581 | v_30671;
assign v_30674 = v_30669 | v_30673;
assign v_30676 = v_30580 | v_30675;
assign v_30678 = v_30578 | v_30677;
assign v_30680 = v_30675 | v_30679;
assign v_30682 = v_30577 | v_30681;
assign v_30684 = v_30575 | v_30683;
assign v_30686 = v_30681 | v_30685;
assign v_30688 = v_30574 | v_30687;
assign v_30690 = v_30572 | v_30689;
assign v_30692 = v_30687 | v_30691;
assign v_30694 = v_30571 | v_30693;
assign v_30696 = v_30569 | v_30695;
assign v_30698 = v_30693 | v_30697;
assign v_30700 = v_30568 | v_30699;
assign v_30702 = v_30566 | v_30701;
assign v_30704 = v_30699 | v_30703;
assign v_30706 = v_30565 | v_30705;
assign v_30708 = v_30563 | v_30707;
assign v_30710 = v_30705 | v_30709;
assign v_30713 = ~v_30562 | v_30712;
assign v_30720 = v_30610 | v_30719;
assign v_30723 = v_30721 | v_30722;
assign v_30725 = v_30607 | v_30724;
assign v_30728 = v_30726 | v_30727;
assign v_30730 = v_30604 | v_30729;
assign v_30733 = v_30731 | v_30732;
assign v_30735 = v_30601 | v_30734;
assign v_30738 = v_30736 | v_30737;
assign v_30740 = v_30598 | v_30739;
assign v_30743 = v_30741 | v_30742;
assign v_30745 = v_30595 | v_30744;
assign v_30748 = v_30746 | v_30747;
assign v_30750 = v_30592 | v_30749;
assign v_30753 = v_30751 | v_30752;
assign v_30755 = v_30589 | v_30754;
assign v_30758 = v_30756 | v_30757;
assign v_30760 = v_30586 | v_30759;
assign v_30763 = v_30761 | v_30762;
assign v_30765 = v_30583 | v_30764;
assign v_30768 = v_30766 | v_30767;
assign v_30770 = v_30580 | v_30769;
assign v_30773 = v_30771 | v_30772;
assign v_30775 = v_30577 | v_30774;
assign v_30778 = v_30776 | v_30777;
assign v_30780 = v_30574 | v_30779;
assign v_30783 = v_30781 | v_30782;
assign v_30785 = v_30571 | v_30784;
assign v_30788 = v_30786 | v_30787;
assign v_30790 = v_30568 | v_30789;
assign v_30793 = v_30791 | v_30792;
assign v_30795 = v_30565 | v_30794;
assign v_30798 = v_30796 | v_30797;
assign v_30800 = v_30562 | v_30799;
assign v_30803 = v_30561 | v_30802;
assign v_30857 = v_30854 | v_30856;
assign v_30859 = v_30853 | v_30858;
assign v_30861 = v_30851 | v_30860;
assign v_30863 = v_30858 | v_30862;
assign v_30865 = v_30850 | v_30864;
assign v_30867 = v_30848 | v_30866;
assign v_30869 = v_30864 | v_30868;
assign v_30871 = v_30847 | v_30870;
assign v_30873 = v_30845 | v_30872;
assign v_30875 = v_30870 | v_30874;
assign v_30877 = v_30844 | v_30876;
assign v_30879 = v_30842 | v_30878;
assign v_30881 = v_30876 | v_30880;
assign v_30883 = v_30841 | v_30882;
assign v_30885 = v_30839 | v_30884;
assign v_30887 = v_30882 | v_30886;
assign v_30889 = v_30838 | v_30888;
assign v_30891 = v_30836 | v_30890;
assign v_30893 = v_30888 | v_30892;
assign v_30895 = v_30835 | v_30894;
assign v_30897 = v_30833 | v_30896;
assign v_30899 = v_30894 | v_30898;
assign v_30901 = v_30832 | v_30900;
assign v_30903 = v_30830 | v_30902;
assign v_30905 = v_30900 | v_30904;
assign v_30907 = v_30829 | v_30906;
assign v_30909 = v_30827 | v_30908;
assign v_30911 = v_30906 | v_30910;
assign v_30913 = v_30826 | v_30912;
assign v_30915 = v_30824 | v_30914;
assign v_30917 = v_30912 | v_30916;
assign v_30919 = v_30823 | v_30918;
assign v_30921 = v_30821 | v_30920;
assign v_30923 = v_30918 | v_30922;
assign v_30925 = v_30820 | v_30924;
assign v_30927 = v_30818 | v_30926;
assign v_30929 = v_30924 | v_30928;
assign v_30931 = v_30817 | v_30930;
assign v_30933 = v_30815 | v_30932;
assign v_30935 = v_30930 | v_30934;
assign v_30937 = v_30814 | v_30936;
assign v_30939 = v_30812 | v_30938;
assign v_30941 = v_30936 | v_30940;
assign v_30943 = v_30811 | v_30942;
assign v_30945 = v_30809 | v_30944;
assign v_30947 = v_30942 | v_30946;
assign v_30949 = v_30808 | v_30948;
assign v_30951 = v_30806 | v_30950;
assign v_30953 = v_30948 | v_30952;
assign v_30956 = ~v_30805 | v_30955;
assign v_30963 = v_30853 | v_30962;
assign v_30966 = v_30964 | v_30965;
assign v_30968 = v_30850 | v_30967;
assign v_30971 = v_30969 | v_30970;
assign v_30973 = v_30847 | v_30972;
assign v_30976 = v_30974 | v_30975;
assign v_30978 = v_30844 | v_30977;
assign v_30981 = v_30979 | v_30980;
assign v_30983 = v_30841 | v_30982;
assign v_30986 = v_30984 | v_30985;
assign v_30988 = v_30838 | v_30987;
assign v_30991 = v_30989 | v_30990;
assign v_30993 = v_30835 | v_30992;
assign v_30996 = v_30994 | v_30995;
assign v_30998 = v_30832 | v_30997;
assign v_31001 = v_30999 | v_31000;
assign v_31003 = v_30829 | v_31002;
assign v_31006 = v_31004 | v_31005;
assign v_31008 = v_30826 | v_31007;
assign v_31011 = v_31009 | v_31010;
assign v_31013 = v_30823 | v_31012;
assign v_31016 = v_31014 | v_31015;
assign v_31018 = v_30820 | v_31017;
assign v_31021 = v_31019 | v_31020;
assign v_31023 = v_30817 | v_31022;
assign v_31026 = v_31024 | v_31025;
assign v_31028 = v_30814 | v_31027;
assign v_31031 = v_31029 | v_31030;
assign v_31033 = v_30811 | v_31032;
assign v_31036 = v_31034 | v_31035;
assign v_31038 = v_30808 | v_31037;
assign v_31041 = v_31039 | v_31040;
assign v_31043 = v_30805 | v_31042;
assign v_31046 = v_30804 | v_31045;
assign v_31100 = v_31097 | v_31099;
assign v_31102 = v_31096 | v_31101;
assign v_31104 = v_31094 | v_31103;
assign v_31106 = v_31101 | v_31105;
assign v_31108 = v_31093 | v_31107;
assign v_31110 = v_31091 | v_31109;
assign v_31112 = v_31107 | v_31111;
assign v_31114 = v_31090 | v_31113;
assign v_31116 = v_31088 | v_31115;
assign v_31118 = v_31113 | v_31117;
assign v_31120 = v_31087 | v_31119;
assign v_31122 = v_31085 | v_31121;
assign v_31124 = v_31119 | v_31123;
assign v_31126 = v_31084 | v_31125;
assign v_31128 = v_31082 | v_31127;
assign v_31130 = v_31125 | v_31129;
assign v_31132 = v_31081 | v_31131;
assign v_31134 = v_31079 | v_31133;
assign v_31136 = v_31131 | v_31135;
assign v_31138 = v_31078 | v_31137;
assign v_31140 = v_31076 | v_31139;
assign v_31142 = v_31137 | v_31141;
assign v_31144 = v_31075 | v_31143;
assign v_31146 = v_31073 | v_31145;
assign v_31148 = v_31143 | v_31147;
assign v_31150 = v_31072 | v_31149;
assign v_31152 = v_31070 | v_31151;
assign v_31154 = v_31149 | v_31153;
assign v_31156 = v_31069 | v_31155;
assign v_31158 = v_31067 | v_31157;
assign v_31160 = v_31155 | v_31159;
assign v_31162 = v_31066 | v_31161;
assign v_31164 = v_31064 | v_31163;
assign v_31166 = v_31161 | v_31165;
assign v_31168 = v_31063 | v_31167;
assign v_31170 = v_31061 | v_31169;
assign v_31172 = v_31167 | v_31171;
assign v_31174 = v_31060 | v_31173;
assign v_31176 = v_31058 | v_31175;
assign v_31178 = v_31173 | v_31177;
assign v_31180 = v_31057 | v_31179;
assign v_31182 = v_31055 | v_31181;
assign v_31184 = v_31179 | v_31183;
assign v_31186 = v_31054 | v_31185;
assign v_31188 = v_31052 | v_31187;
assign v_31190 = v_31185 | v_31189;
assign v_31192 = v_31051 | v_31191;
assign v_31194 = v_31049 | v_31193;
assign v_31196 = v_31191 | v_31195;
assign v_31199 = ~v_31048 | v_31198;
assign v_31206 = v_31096 | v_31205;
assign v_31209 = v_31207 | v_31208;
assign v_31211 = v_31093 | v_31210;
assign v_31214 = v_31212 | v_31213;
assign v_31216 = v_31090 | v_31215;
assign v_31219 = v_31217 | v_31218;
assign v_31221 = v_31087 | v_31220;
assign v_31224 = v_31222 | v_31223;
assign v_31226 = v_31084 | v_31225;
assign v_31229 = v_31227 | v_31228;
assign v_31231 = v_31081 | v_31230;
assign v_31234 = v_31232 | v_31233;
assign v_31236 = v_31078 | v_31235;
assign v_31239 = v_31237 | v_31238;
assign v_31241 = v_31075 | v_31240;
assign v_31244 = v_31242 | v_31243;
assign v_31246 = v_31072 | v_31245;
assign v_31249 = v_31247 | v_31248;
assign v_31251 = v_31069 | v_31250;
assign v_31254 = v_31252 | v_31253;
assign v_31256 = v_31066 | v_31255;
assign v_31259 = v_31257 | v_31258;
assign v_31261 = v_31063 | v_31260;
assign v_31264 = v_31262 | v_31263;
assign v_31266 = v_31060 | v_31265;
assign v_31269 = v_31267 | v_31268;
assign v_31271 = v_31057 | v_31270;
assign v_31274 = v_31272 | v_31273;
assign v_31276 = v_31054 | v_31275;
assign v_31279 = v_31277 | v_31278;
assign v_31281 = v_31051 | v_31280;
assign v_31284 = v_31282 | v_31283;
assign v_31286 = v_31048 | v_31285;
assign v_31289 = v_31047 | v_31288;
assign v_31343 = v_31340 | v_31342;
assign v_31345 = v_31339 | v_31344;
assign v_31347 = v_31337 | v_31346;
assign v_31349 = v_31344 | v_31348;
assign v_31351 = v_31336 | v_31350;
assign v_31353 = v_31334 | v_31352;
assign v_31355 = v_31350 | v_31354;
assign v_31357 = v_31333 | v_31356;
assign v_31359 = v_31331 | v_31358;
assign v_31361 = v_31356 | v_31360;
assign v_31363 = v_31330 | v_31362;
assign v_31365 = v_31328 | v_31364;
assign v_31367 = v_31362 | v_31366;
assign v_31369 = v_31327 | v_31368;
assign v_31371 = v_31325 | v_31370;
assign v_31373 = v_31368 | v_31372;
assign v_31375 = v_31324 | v_31374;
assign v_31377 = v_31322 | v_31376;
assign v_31379 = v_31374 | v_31378;
assign v_31381 = v_31321 | v_31380;
assign v_31383 = v_31319 | v_31382;
assign v_31385 = v_31380 | v_31384;
assign v_31387 = v_31318 | v_31386;
assign v_31389 = v_31316 | v_31388;
assign v_31391 = v_31386 | v_31390;
assign v_31393 = v_31315 | v_31392;
assign v_31395 = v_31313 | v_31394;
assign v_31397 = v_31392 | v_31396;
assign v_31399 = v_31312 | v_31398;
assign v_31401 = v_31310 | v_31400;
assign v_31403 = v_31398 | v_31402;
assign v_31405 = v_31309 | v_31404;
assign v_31407 = v_31307 | v_31406;
assign v_31409 = v_31404 | v_31408;
assign v_31411 = v_31306 | v_31410;
assign v_31413 = v_31304 | v_31412;
assign v_31415 = v_31410 | v_31414;
assign v_31417 = v_31303 | v_31416;
assign v_31419 = v_31301 | v_31418;
assign v_31421 = v_31416 | v_31420;
assign v_31423 = v_31300 | v_31422;
assign v_31425 = v_31298 | v_31424;
assign v_31427 = v_31422 | v_31426;
assign v_31429 = v_31297 | v_31428;
assign v_31431 = v_31295 | v_31430;
assign v_31433 = v_31428 | v_31432;
assign v_31435 = v_31294 | v_31434;
assign v_31437 = v_31292 | v_31436;
assign v_31439 = v_31434 | v_31438;
assign v_31442 = ~v_31291 | v_31441;
assign v_31449 = v_31339 | v_31448;
assign v_31452 = v_31450 | v_31451;
assign v_31454 = v_31336 | v_31453;
assign v_31457 = v_31455 | v_31456;
assign v_31459 = v_31333 | v_31458;
assign v_31462 = v_31460 | v_31461;
assign v_31464 = v_31330 | v_31463;
assign v_31467 = v_31465 | v_31466;
assign v_31469 = v_31327 | v_31468;
assign v_31472 = v_31470 | v_31471;
assign v_31474 = v_31324 | v_31473;
assign v_31477 = v_31475 | v_31476;
assign v_31479 = v_31321 | v_31478;
assign v_31482 = v_31480 | v_31481;
assign v_31484 = v_31318 | v_31483;
assign v_31487 = v_31485 | v_31486;
assign v_31489 = v_31315 | v_31488;
assign v_31492 = v_31490 | v_31491;
assign v_31494 = v_31312 | v_31493;
assign v_31497 = v_31495 | v_31496;
assign v_31499 = v_31309 | v_31498;
assign v_31502 = v_31500 | v_31501;
assign v_31504 = v_31306 | v_31503;
assign v_31507 = v_31505 | v_31506;
assign v_31509 = v_31303 | v_31508;
assign v_31512 = v_31510 | v_31511;
assign v_31514 = v_31300 | v_31513;
assign v_31517 = v_31515 | v_31516;
assign v_31519 = v_31297 | v_31518;
assign v_31522 = v_31520 | v_31521;
assign v_31524 = v_31294 | v_31523;
assign v_31527 = v_31525 | v_31526;
assign v_31529 = v_31291 | v_31528;
assign v_31532 = v_31290 | v_31531;
assign v_31586 = v_31583 | v_31585;
assign v_31588 = v_31582 | v_31587;
assign v_31590 = v_31580 | v_31589;
assign v_31592 = v_31587 | v_31591;
assign v_31594 = v_31579 | v_31593;
assign v_31596 = v_31577 | v_31595;
assign v_31598 = v_31593 | v_31597;
assign v_31600 = v_31576 | v_31599;
assign v_31602 = v_31574 | v_31601;
assign v_31604 = v_31599 | v_31603;
assign v_31606 = v_31573 | v_31605;
assign v_31608 = v_31571 | v_31607;
assign v_31610 = v_31605 | v_31609;
assign v_31612 = v_31570 | v_31611;
assign v_31614 = v_31568 | v_31613;
assign v_31616 = v_31611 | v_31615;
assign v_31618 = v_31567 | v_31617;
assign v_31620 = v_31565 | v_31619;
assign v_31622 = v_31617 | v_31621;
assign v_31624 = v_31564 | v_31623;
assign v_31626 = v_31562 | v_31625;
assign v_31628 = v_31623 | v_31627;
assign v_31630 = v_31561 | v_31629;
assign v_31632 = v_31559 | v_31631;
assign v_31634 = v_31629 | v_31633;
assign v_31636 = v_31558 | v_31635;
assign v_31638 = v_31556 | v_31637;
assign v_31640 = v_31635 | v_31639;
assign v_31642 = v_31555 | v_31641;
assign v_31644 = v_31553 | v_31643;
assign v_31646 = v_31641 | v_31645;
assign v_31648 = v_31552 | v_31647;
assign v_31650 = v_31550 | v_31649;
assign v_31652 = v_31647 | v_31651;
assign v_31654 = v_31549 | v_31653;
assign v_31656 = v_31547 | v_31655;
assign v_31658 = v_31653 | v_31657;
assign v_31660 = v_31546 | v_31659;
assign v_31662 = v_31544 | v_31661;
assign v_31664 = v_31659 | v_31663;
assign v_31666 = v_31543 | v_31665;
assign v_31668 = v_31541 | v_31667;
assign v_31670 = v_31665 | v_31669;
assign v_31672 = v_31540 | v_31671;
assign v_31674 = v_31538 | v_31673;
assign v_31676 = v_31671 | v_31675;
assign v_31678 = v_31537 | v_31677;
assign v_31680 = v_31535 | v_31679;
assign v_31682 = v_31677 | v_31681;
assign v_31685 = ~v_31534 | v_31684;
assign v_31692 = v_31582 | v_31691;
assign v_31695 = v_31693 | v_31694;
assign v_31697 = v_31579 | v_31696;
assign v_31700 = v_31698 | v_31699;
assign v_31702 = v_31576 | v_31701;
assign v_31705 = v_31703 | v_31704;
assign v_31707 = v_31573 | v_31706;
assign v_31710 = v_31708 | v_31709;
assign v_31712 = v_31570 | v_31711;
assign v_31715 = v_31713 | v_31714;
assign v_31717 = v_31567 | v_31716;
assign v_31720 = v_31718 | v_31719;
assign v_31722 = v_31564 | v_31721;
assign v_31725 = v_31723 | v_31724;
assign v_31727 = v_31561 | v_31726;
assign v_31730 = v_31728 | v_31729;
assign v_31732 = v_31558 | v_31731;
assign v_31735 = v_31733 | v_31734;
assign v_31737 = v_31555 | v_31736;
assign v_31740 = v_31738 | v_31739;
assign v_31742 = v_31552 | v_31741;
assign v_31745 = v_31743 | v_31744;
assign v_31747 = v_31549 | v_31746;
assign v_31750 = v_31748 | v_31749;
assign v_31752 = v_31546 | v_31751;
assign v_31755 = v_31753 | v_31754;
assign v_31757 = v_31543 | v_31756;
assign v_31760 = v_31758 | v_31759;
assign v_31762 = v_31540 | v_31761;
assign v_31765 = v_31763 | v_31764;
assign v_31767 = v_31537 | v_31766;
assign v_31770 = v_31768 | v_31769;
assign v_31772 = v_31534 | v_31771;
assign v_31775 = v_31533 | v_31774;
assign v_31829 = v_31826 | v_31828;
assign v_31831 = v_31825 | v_31830;
assign v_31833 = v_31823 | v_31832;
assign v_31835 = v_31830 | v_31834;
assign v_31837 = v_31822 | v_31836;
assign v_31839 = v_31820 | v_31838;
assign v_31841 = v_31836 | v_31840;
assign v_31843 = v_31819 | v_31842;
assign v_31845 = v_31817 | v_31844;
assign v_31847 = v_31842 | v_31846;
assign v_31849 = v_31816 | v_31848;
assign v_31851 = v_31814 | v_31850;
assign v_31853 = v_31848 | v_31852;
assign v_31855 = v_31813 | v_31854;
assign v_31857 = v_31811 | v_31856;
assign v_31859 = v_31854 | v_31858;
assign v_31861 = v_31810 | v_31860;
assign v_31863 = v_31808 | v_31862;
assign v_31865 = v_31860 | v_31864;
assign v_31867 = v_31807 | v_31866;
assign v_31869 = v_31805 | v_31868;
assign v_31871 = v_31866 | v_31870;
assign v_31873 = v_31804 | v_31872;
assign v_31875 = v_31802 | v_31874;
assign v_31877 = v_31872 | v_31876;
assign v_31879 = v_31801 | v_31878;
assign v_31881 = v_31799 | v_31880;
assign v_31883 = v_31878 | v_31882;
assign v_31885 = v_31798 | v_31884;
assign v_31887 = v_31796 | v_31886;
assign v_31889 = v_31884 | v_31888;
assign v_31891 = v_31795 | v_31890;
assign v_31893 = v_31793 | v_31892;
assign v_31895 = v_31890 | v_31894;
assign v_31897 = v_31792 | v_31896;
assign v_31899 = v_31790 | v_31898;
assign v_31901 = v_31896 | v_31900;
assign v_31903 = v_31789 | v_31902;
assign v_31905 = v_31787 | v_31904;
assign v_31907 = v_31902 | v_31906;
assign v_31909 = v_31786 | v_31908;
assign v_31911 = v_31784 | v_31910;
assign v_31913 = v_31908 | v_31912;
assign v_31915 = v_31783 | v_31914;
assign v_31917 = v_31781 | v_31916;
assign v_31919 = v_31914 | v_31918;
assign v_31921 = v_31780 | v_31920;
assign v_31923 = v_31778 | v_31922;
assign v_31925 = v_31920 | v_31924;
assign v_31928 = ~v_31777 | v_31927;
assign v_31935 = v_31825 | v_31934;
assign v_31938 = v_31936 | v_31937;
assign v_31940 = v_31822 | v_31939;
assign v_31943 = v_31941 | v_31942;
assign v_31945 = v_31819 | v_31944;
assign v_31948 = v_31946 | v_31947;
assign v_31950 = v_31816 | v_31949;
assign v_31953 = v_31951 | v_31952;
assign v_31955 = v_31813 | v_31954;
assign v_31958 = v_31956 | v_31957;
assign v_31960 = v_31810 | v_31959;
assign v_31963 = v_31961 | v_31962;
assign v_31965 = v_31807 | v_31964;
assign v_31968 = v_31966 | v_31967;
assign v_31970 = v_31804 | v_31969;
assign v_31973 = v_31971 | v_31972;
assign v_31975 = v_31801 | v_31974;
assign v_31978 = v_31976 | v_31977;
assign v_31980 = v_31798 | v_31979;
assign v_31983 = v_31981 | v_31982;
assign v_31985 = v_31795 | v_31984;
assign v_31988 = v_31986 | v_31987;
assign v_31990 = v_31792 | v_31989;
assign v_31993 = v_31991 | v_31992;
assign v_31995 = v_31789 | v_31994;
assign v_31998 = v_31996 | v_31997;
assign v_32000 = v_31786 | v_31999;
assign v_32003 = v_32001 | v_32002;
assign v_32005 = v_31783 | v_32004;
assign v_32008 = v_32006 | v_32007;
assign v_32010 = v_31780 | v_32009;
assign v_32013 = v_32011 | v_32012;
assign v_32015 = v_31777 | v_32014;
assign v_32018 = v_31776 | v_32017;
assign v_32072 = v_32069 | v_32071;
assign v_32074 = v_32068 | v_32073;
assign v_32076 = v_32066 | v_32075;
assign v_32078 = v_32073 | v_32077;
assign v_32080 = v_32065 | v_32079;
assign v_32082 = v_32063 | v_32081;
assign v_32084 = v_32079 | v_32083;
assign v_32086 = v_32062 | v_32085;
assign v_32088 = v_32060 | v_32087;
assign v_32090 = v_32085 | v_32089;
assign v_32092 = v_32059 | v_32091;
assign v_32094 = v_32057 | v_32093;
assign v_32096 = v_32091 | v_32095;
assign v_32098 = v_32056 | v_32097;
assign v_32100 = v_32054 | v_32099;
assign v_32102 = v_32097 | v_32101;
assign v_32104 = v_32053 | v_32103;
assign v_32106 = v_32051 | v_32105;
assign v_32108 = v_32103 | v_32107;
assign v_32110 = v_32050 | v_32109;
assign v_32112 = v_32048 | v_32111;
assign v_32114 = v_32109 | v_32113;
assign v_32116 = v_32047 | v_32115;
assign v_32118 = v_32045 | v_32117;
assign v_32120 = v_32115 | v_32119;
assign v_32122 = v_32044 | v_32121;
assign v_32124 = v_32042 | v_32123;
assign v_32126 = v_32121 | v_32125;
assign v_32128 = v_32041 | v_32127;
assign v_32130 = v_32039 | v_32129;
assign v_32132 = v_32127 | v_32131;
assign v_32134 = v_32038 | v_32133;
assign v_32136 = v_32036 | v_32135;
assign v_32138 = v_32133 | v_32137;
assign v_32140 = v_32035 | v_32139;
assign v_32142 = v_32033 | v_32141;
assign v_32144 = v_32139 | v_32143;
assign v_32146 = v_32032 | v_32145;
assign v_32148 = v_32030 | v_32147;
assign v_32150 = v_32145 | v_32149;
assign v_32152 = v_32029 | v_32151;
assign v_32154 = v_32027 | v_32153;
assign v_32156 = v_32151 | v_32155;
assign v_32158 = v_32026 | v_32157;
assign v_32160 = v_32024 | v_32159;
assign v_32162 = v_32157 | v_32161;
assign v_32164 = v_32023 | v_32163;
assign v_32166 = v_32021 | v_32165;
assign v_32168 = v_32163 | v_32167;
assign v_32171 = ~v_32020 | v_32170;
assign v_32178 = v_32068 | v_32177;
assign v_32181 = v_32179 | v_32180;
assign v_32183 = v_32065 | v_32182;
assign v_32186 = v_32184 | v_32185;
assign v_32188 = v_32062 | v_32187;
assign v_32191 = v_32189 | v_32190;
assign v_32193 = v_32059 | v_32192;
assign v_32196 = v_32194 | v_32195;
assign v_32198 = v_32056 | v_32197;
assign v_32201 = v_32199 | v_32200;
assign v_32203 = v_32053 | v_32202;
assign v_32206 = v_32204 | v_32205;
assign v_32208 = v_32050 | v_32207;
assign v_32211 = v_32209 | v_32210;
assign v_32213 = v_32047 | v_32212;
assign v_32216 = v_32214 | v_32215;
assign v_32218 = v_32044 | v_32217;
assign v_32221 = v_32219 | v_32220;
assign v_32223 = v_32041 | v_32222;
assign v_32226 = v_32224 | v_32225;
assign v_32228 = v_32038 | v_32227;
assign v_32231 = v_32229 | v_32230;
assign v_32233 = v_32035 | v_32232;
assign v_32236 = v_32234 | v_32235;
assign v_32238 = v_32032 | v_32237;
assign v_32241 = v_32239 | v_32240;
assign v_32243 = v_32029 | v_32242;
assign v_32246 = v_32244 | v_32245;
assign v_32248 = v_32026 | v_32247;
assign v_32251 = v_32249 | v_32250;
assign v_32253 = v_32023 | v_32252;
assign v_32256 = v_32254 | v_32255;
assign v_32258 = v_32020 | v_32257;
assign v_32261 = v_32019 | v_32260;
assign v_32315 = v_32312 | v_32314;
assign v_32317 = v_32311 | v_32316;
assign v_32319 = v_32309 | v_32318;
assign v_32321 = v_32316 | v_32320;
assign v_32323 = v_32308 | v_32322;
assign v_32325 = v_32306 | v_32324;
assign v_32327 = v_32322 | v_32326;
assign v_32329 = v_32305 | v_32328;
assign v_32331 = v_32303 | v_32330;
assign v_32333 = v_32328 | v_32332;
assign v_32335 = v_32302 | v_32334;
assign v_32337 = v_32300 | v_32336;
assign v_32339 = v_32334 | v_32338;
assign v_32341 = v_32299 | v_32340;
assign v_32343 = v_32297 | v_32342;
assign v_32345 = v_32340 | v_32344;
assign v_32347 = v_32296 | v_32346;
assign v_32349 = v_32294 | v_32348;
assign v_32351 = v_32346 | v_32350;
assign v_32353 = v_32293 | v_32352;
assign v_32355 = v_32291 | v_32354;
assign v_32357 = v_32352 | v_32356;
assign v_32359 = v_32290 | v_32358;
assign v_32361 = v_32288 | v_32360;
assign v_32363 = v_32358 | v_32362;
assign v_32365 = v_32287 | v_32364;
assign v_32367 = v_32285 | v_32366;
assign v_32369 = v_32364 | v_32368;
assign v_32371 = v_32284 | v_32370;
assign v_32373 = v_32282 | v_32372;
assign v_32375 = v_32370 | v_32374;
assign v_32377 = v_32281 | v_32376;
assign v_32379 = v_32279 | v_32378;
assign v_32381 = v_32376 | v_32380;
assign v_32383 = v_32278 | v_32382;
assign v_32385 = v_32276 | v_32384;
assign v_32387 = v_32382 | v_32386;
assign v_32389 = v_32275 | v_32388;
assign v_32391 = v_32273 | v_32390;
assign v_32393 = v_32388 | v_32392;
assign v_32395 = v_32272 | v_32394;
assign v_32397 = v_32270 | v_32396;
assign v_32399 = v_32394 | v_32398;
assign v_32401 = v_32269 | v_32400;
assign v_32403 = v_32267 | v_32402;
assign v_32405 = v_32400 | v_32404;
assign v_32407 = v_32266 | v_32406;
assign v_32409 = v_32264 | v_32408;
assign v_32411 = v_32406 | v_32410;
assign v_32414 = ~v_32263 | v_32413;
assign v_32421 = v_32311 | v_32420;
assign v_32424 = v_32422 | v_32423;
assign v_32426 = v_32308 | v_32425;
assign v_32429 = v_32427 | v_32428;
assign v_32431 = v_32305 | v_32430;
assign v_32434 = v_32432 | v_32433;
assign v_32436 = v_32302 | v_32435;
assign v_32439 = v_32437 | v_32438;
assign v_32441 = v_32299 | v_32440;
assign v_32444 = v_32442 | v_32443;
assign v_32446 = v_32296 | v_32445;
assign v_32449 = v_32447 | v_32448;
assign v_32451 = v_32293 | v_32450;
assign v_32454 = v_32452 | v_32453;
assign v_32456 = v_32290 | v_32455;
assign v_32459 = v_32457 | v_32458;
assign v_32461 = v_32287 | v_32460;
assign v_32464 = v_32462 | v_32463;
assign v_32466 = v_32284 | v_32465;
assign v_32469 = v_32467 | v_32468;
assign v_32471 = v_32281 | v_32470;
assign v_32474 = v_32472 | v_32473;
assign v_32476 = v_32278 | v_32475;
assign v_32479 = v_32477 | v_32478;
assign v_32481 = v_32275 | v_32480;
assign v_32484 = v_32482 | v_32483;
assign v_32486 = v_32272 | v_32485;
assign v_32489 = v_32487 | v_32488;
assign v_32491 = v_32269 | v_32490;
assign v_32494 = v_32492 | v_32493;
assign v_32496 = v_32266 | v_32495;
assign v_32499 = v_32497 | v_32498;
assign v_32501 = v_32263 | v_32500;
assign v_32504 = v_32262 | v_32503;
assign v_32558 = v_32555 | v_32557;
assign v_32560 = v_32554 | v_32559;
assign v_32562 = v_32552 | v_32561;
assign v_32564 = v_32559 | v_32563;
assign v_32566 = v_32551 | v_32565;
assign v_32568 = v_32549 | v_32567;
assign v_32570 = v_32565 | v_32569;
assign v_32572 = v_32548 | v_32571;
assign v_32574 = v_32546 | v_32573;
assign v_32576 = v_32571 | v_32575;
assign v_32578 = v_32545 | v_32577;
assign v_32580 = v_32543 | v_32579;
assign v_32582 = v_32577 | v_32581;
assign v_32584 = v_32542 | v_32583;
assign v_32586 = v_32540 | v_32585;
assign v_32588 = v_32583 | v_32587;
assign v_32590 = v_32539 | v_32589;
assign v_32592 = v_32537 | v_32591;
assign v_32594 = v_32589 | v_32593;
assign v_32596 = v_32536 | v_32595;
assign v_32598 = v_32534 | v_32597;
assign v_32600 = v_32595 | v_32599;
assign v_32602 = v_32533 | v_32601;
assign v_32604 = v_32531 | v_32603;
assign v_32606 = v_32601 | v_32605;
assign v_32608 = v_32530 | v_32607;
assign v_32610 = v_32528 | v_32609;
assign v_32612 = v_32607 | v_32611;
assign v_32614 = v_32527 | v_32613;
assign v_32616 = v_32525 | v_32615;
assign v_32618 = v_32613 | v_32617;
assign v_32620 = v_32524 | v_32619;
assign v_32622 = v_32522 | v_32621;
assign v_32624 = v_32619 | v_32623;
assign v_32626 = v_32521 | v_32625;
assign v_32628 = v_32519 | v_32627;
assign v_32630 = v_32625 | v_32629;
assign v_32632 = v_32518 | v_32631;
assign v_32634 = v_32516 | v_32633;
assign v_32636 = v_32631 | v_32635;
assign v_32638 = v_32515 | v_32637;
assign v_32640 = v_32513 | v_32639;
assign v_32642 = v_32637 | v_32641;
assign v_32644 = v_32512 | v_32643;
assign v_32646 = v_32510 | v_32645;
assign v_32648 = v_32643 | v_32647;
assign v_32650 = v_32509 | v_32649;
assign v_32652 = v_32507 | v_32651;
assign v_32654 = v_32649 | v_32653;
assign v_32657 = ~v_32506 | v_32656;
assign v_32664 = v_32554 | v_32663;
assign v_32667 = v_32665 | v_32666;
assign v_32669 = v_32551 | v_32668;
assign v_32672 = v_32670 | v_32671;
assign v_32674 = v_32548 | v_32673;
assign v_32677 = v_32675 | v_32676;
assign v_32679 = v_32545 | v_32678;
assign v_32682 = v_32680 | v_32681;
assign v_32684 = v_32542 | v_32683;
assign v_32687 = v_32685 | v_32686;
assign v_32689 = v_32539 | v_32688;
assign v_32692 = v_32690 | v_32691;
assign v_32694 = v_32536 | v_32693;
assign v_32697 = v_32695 | v_32696;
assign v_32699 = v_32533 | v_32698;
assign v_32702 = v_32700 | v_32701;
assign v_32704 = v_32530 | v_32703;
assign v_32707 = v_32705 | v_32706;
assign v_32709 = v_32527 | v_32708;
assign v_32712 = v_32710 | v_32711;
assign v_32714 = v_32524 | v_32713;
assign v_32717 = v_32715 | v_32716;
assign v_32719 = v_32521 | v_32718;
assign v_32722 = v_32720 | v_32721;
assign v_32724 = v_32518 | v_32723;
assign v_32727 = v_32725 | v_32726;
assign v_32729 = v_32515 | v_32728;
assign v_32732 = v_32730 | v_32731;
assign v_32734 = v_32512 | v_32733;
assign v_32737 = v_32735 | v_32736;
assign v_32739 = v_32509 | v_32738;
assign v_32742 = v_32740 | v_32741;
assign v_32744 = v_32506 | v_32743;
assign v_32747 = v_32505 | v_32746;
assign v_32801 = v_32798 | v_32800;
assign v_32803 = v_32797 | v_32802;
assign v_32805 = v_32795 | v_32804;
assign v_32807 = v_32802 | v_32806;
assign v_32809 = v_32794 | v_32808;
assign v_32811 = v_32792 | v_32810;
assign v_32813 = v_32808 | v_32812;
assign v_32815 = v_32791 | v_32814;
assign v_32817 = v_32789 | v_32816;
assign v_32819 = v_32814 | v_32818;
assign v_32821 = v_32788 | v_32820;
assign v_32823 = v_32786 | v_32822;
assign v_32825 = v_32820 | v_32824;
assign v_32827 = v_32785 | v_32826;
assign v_32829 = v_32783 | v_32828;
assign v_32831 = v_32826 | v_32830;
assign v_32833 = v_32782 | v_32832;
assign v_32835 = v_32780 | v_32834;
assign v_32837 = v_32832 | v_32836;
assign v_32839 = v_32779 | v_32838;
assign v_32841 = v_32777 | v_32840;
assign v_32843 = v_32838 | v_32842;
assign v_32845 = v_32776 | v_32844;
assign v_32847 = v_32774 | v_32846;
assign v_32849 = v_32844 | v_32848;
assign v_32851 = v_32773 | v_32850;
assign v_32853 = v_32771 | v_32852;
assign v_32855 = v_32850 | v_32854;
assign v_32857 = v_32770 | v_32856;
assign v_32859 = v_32768 | v_32858;
assign v_32861 = v_32856 | v_32860;
assign v_32863 = v_32767 | v_32862;
assign v_32865 = v_32765 | v_32864;
assign v_32867 = v_32862 | v_32866;
assign v_32869 = v_32764 | v_32868;
assign v_32871 = v_32762 | v_32870;
assign v_32873 = v_32868 | v_32872;
assign v_32875 = v_32761 | v_32874;
assign v_32877 = v_32759 | v_32876;
assign v_32879 = v_32874 | v_32878;
assign v_32881 = v_32758 | v_32880;
assign v_32883 = v_32756 | v_32882;
assign v_32885 = v_32880 | v_32884;
assign v_32887 = v_32755 | v_32886;
assign v_32889 = v_32753 | v_32888;
assign v_32891 = v_32886 | v_32890;
assign v_32893 = v_32752 | v_32892;
assign v_32895 = v_32750 | v_32894;
assign v_32897 = v_32892 | v_32896;
assign v_32900 = ~v_32749 | v_32899;
assign v_32907 = v_32797 | v_32906;
assign v_32910 = v_32908 | v_32909;
assign v_32912 = v_32794 | v_32911;
assign v_32915 = v_32913 | v_32914;
assign v_32917 = v_32791 | v_32916;
assign v_32920 = v_32918 | v_32919;
assign v_32922 = v_32788 | v_32921;
assign v_32925 = v_32923 | v_32924;
assign v_32927 = v_32785 | v_32926;
assign v_32930 = v_32928 | v_32929;
assign v_32932 = v_32782 | v_32931;
assign v_32935 = v_32933 | v_32934;
assign v_32937 = v_32779 | v_32936;
assign v_32940 = v_32938 | v_32939;
assign v_32942 = v_32776 | v_32941;
assign v_32945 = v_32943 | v_32944;
assign v_32947 = v_32773 | v_32946;
assign v_32950 = v_32948 | v_32949;
assign v_32952 = v_32770 | v_32951;
assign v_32955 = v_32953 | v_32954;
assign v_32957 = v_32767 | v_32956;
assign v_32960 = v_32958 | v_32959;
assign v_32962 = v_32764 | v_32961;
assign v_32965 = v_32963 | v_32964;
assign v_32967 = v_32761 | v_32966;
assign v_32970 = v_32968 | v_32969;
assign v_32972 = v_32758 | v_32971;
assign v_32975 = v_32973 | v_32974;
assign v_32977 = v_32755 | v_32976;
assign v_32980 = v_32978 | v_32979;
assign v_32982 = v_32752 | v_32981;
assign v_32985 = v_32983 | v_32984;
assign v_32987 = v_32749 | v_32986;
assign v_32990 = v_32748 | v_32989;
assign v_33044 = v_33041 | v_33043;
assign v_33046 = v_33040 | v_33045;
assign v_33048 = v_33038 | v_33047;
assign v_33050 = v_33045 | v_33049;
assign v_33052 = v_33037 | v_33051;
assign v_33054 = v_33035 | v_33053;
assign v_33056 = v_33051 | v_33055;
assign v_33058 = v_33034 | v_33057;
assign v_33060 = v_33032 | v_33059;
assign v_33062 = v_33057 | v_33061;
assign v_33064 = v_33031 | v_33063;
assign v_33066 = v_33029 | v_33065;
assign v_33068 = v_33063 | v_33067;
assign v_33070 = v_33028 | v_33069;
assign v_33072 = v_33026 | v_33071;
assign v_33074 = v_33069 | v_33073;
assign v_33076 = v_33025 | v_33075;
assign v_33078 = v_33023 | v_33077;
assign v_33080 = v_33075 | v_33079;
assign v_33082 = v_33022 | v_33081;
assign v_33084 = v_33020 | v_33083;
assign v_33086 = v_33081 | v_33085;
assign v_33088 = v_33019 | v_33087;
assign v_33090 = v_33017 | v_33089;
assign v_33092 = v_33087 | v_33091;
assign v_33094 = v_33016 | v_33093;
assign v_33096 = v_33014 | v_33095;
assign v_33098 = v_33093 | v_33097;
assign v_33100 = v_33013 | v_33099;
assign v_33102 = v_33011 | v_33101;
assign v_33104 = v_33099 | v_33103;
assign v_33106 = v_33010 | v_33105;
assign v_33108 = v_33008 | v_33107;
assign v_33110 = v_33105 | v_33109;
assign v_33112 = v_33007 | v_33111;
assign v_33114 = v_33005 | v_33113;
assign v_33116 = v_33111 | v_33115;
assign v_33118 = v_33004 | v_33117;
assign v_33120 = v_33002 | v_33119;
assign v_33122 = v_33117 | v_33121;
assign v_33124 = v_33001 | v_33123;
assign v_33126 = v_32999 | v_33125;
assign v_33128 = v_33123 | v_33127;
assign v_33130 = v_32998 | v_33129;
assign v_33132 = v_32996 | v_33131;
assign v_33134 = v_33129 | v_33133;
assign v_33136 = v_32995 | v_33135;
assign v_33138 = v_32993 | v_33137;
assign v_33140 = v_33135 | v_33139;
assign v_33143 = ~v_32992 | v_33142;
assign v_33150 = v_33040 | v_33149;
assign v_33153 = v_33151 | v_33152;
assign v_33155 = v_33037 | v_33154;
assign v_33158 = v_33156 | v_33157;
assign v_33160 = v_33034 | v_33159;
assign v_33163 = v_33161 | v_33162;
assign v_33165 = v_33031 | v_33164;
assign v_33168 = v_33166 | v_33167;
assign v_33170 = v_33028 | v_33169;
assign v_33173 = v_33171 | v_33172;
assign v_33175 = v_33025 | v_33174;
assign v_33178 = v_33176 | v_33177;
assign v_33180 = v_33022 | v_33179;
assign v_33183 = v_33181 | v_33182;
assign v_33185 = v_33019 | v_33184;
assign v_33188 = v_33186 | v_33187;
assign v_33190 = v_33016 | v_33189;
assign v_33193 = v_33191 | v_33192;
assign v_33195 = v_33013 | v_33194;
assign v_33198 = v_33196 | v_33197;
assign v_33200 = v_33010 | v_33199;
assign v_33203 = v_33201 | v_33202;
assign v_33205 = v_33007 | v_33204;
assign v_33208 = v_33206 | v_33207;
assign v_33210 = v_33004 | v_33209;
assign v_33213 = v_33211 | v_33212;
assign v_33215 = v_33001 | v_33214;
assign v_33218 = v_33216 | v_33217;
assign v_33220 = v_32998 | v_33219;
assign v_33223 = v_33221 | v_33222;
assign v_33225 = v_32995 | v_33224;
assign v_33228 = v_33226 | v_33227;
assign v_33230 = v_32992 | v_33229;
assign v_33233 = v_32991 | v_33232;
assign v_33286 = v_33283 | v_33285;
assign v_33288 = v_33282 | v_33287;
assign v_33290 = v_33280 | v_33289;
assign v_33292 = v_33287 | v_33291;
assign v_33294 = v_33279 | v_33293;
assign v_33296 = v_33277 | v_33295;
assign v_33298 = v_33293 | v_33297;
assign v_33300 = v_33276 | v_33299;
assign v_33302 = v_33274 | v_33301;
assign v_33304 = v_33299 | v_33303;
assign v_33306 = v_33273 | v_33305;
assign v_33308 = v_33271 | v_33307;
assign v_33310 = v_33305 | v_33309;
assign v_33312 = v_33270 | v_33311;
assign v_33314 = v_33268 | v_33313;
assign v_33316 = v_33311 | v_33315;
assign v_33318 = v_33267 | v_33317;
assign v_33320 = v_33265 | v_33319;
assign v_33322 = v_33317 | v_33321;
assign v_33324 = v_33264 | v_33323;
assign v_33326 = v_33262 | v_33325;
assign v_33328 = v_33323 | v_33327;
assign v_33330 = v_33261 | v_33329;
assign v_33332 = v_33259 | v_33331;
assign v_33334 = v_33329 | v_33333;
assign v_33336 = v_33258 | v_33335;
assign v_33338 = v_33256 | v_33337;
assign v_33340 = v_33335 | v_33339;
assign v_33342 = v_33255 | v_33341;
assign v_33344 = v_33253 | v_33343;
assign v_33346 = v_33341 | v_33345;
assign v_33348 = v_33252 | v_33347;
assign v_33350 = v_33250 | v_33349;
assign v_33352 = v_33347 | v_33351;
assign v_33354 = v_33249 | v_33353;
assign v_33356 = v_33247 | v_33355;
assign v_33358 = v_33353 | v_33357;
assign v_33360 = v_33246 | v_33359;
assign v_33362 = v_33244 | v_33361;
assign v_33364 = v_33359 | v_33363;
assign v_33366 = v_33243 | v_33365;
assign v_33368 = v_33241 | v_33367;
assign v_33370 = v_33365 | v_33369;
assign v_33372 = v_33240 | v_33371;
assign v_33374 = v_33238 | v_33373;
assign v_33376 = v_33371 | v_33375;
assign v_33378 = v_33237 | v_33377;
assign v_33380 = v_33235 | v_33379;
assign v_33382 = v_33377 | v_33381;
assign v_33386 = v_33383 | v_33385;
assign v_33393 = v_33282 | v_33392;
assign v_33396 = v_33394 | v_33395;
assign v_33398 = v_33279 | v_33397;
assign v_33401 = v_33399 | v_33400;
assign v_33403 = v_33276 | v_33402;
assign v_33406 = v_33404 | v_33405;
assign v_33408 = v_33273 | v_33407;
assign v_33411 = v_33409 | v_33410;
assign v_33413 = v_33270 | v_33412;
assign v_33416 = v_33414 | v_33415;
assign v_33418 = v_33267 | v_33417;
assign v_33421 = v_33419 | v_33420;
assign v_33423 = v_33264 | v_33422;
assign v_33426 = v_33424 | v_33425;
assign v_33428 = v_33261 | v_33427;
assign v_33431 = v_33429 | v_33430;
assign v_33433 = v_33258 | v_33432;
assign v_33436 = v_33434 | v_33435;
assign v_33438 = v_33255 | v_33437;
assign v_33441 = v_33439 | v_33440;
assign v_33443 = v_33252 | v_33442;
assign v_33446 = v_33444 | v_33445;
assign v_33448 = v_33249 | v_33447;
assign v_33451 = v_33449 | v_33450;
assign v_33453 = v_33246 | v_33452;
assign v_33456 = v_33454 | v_33455;
assign v_33458 = v_33243 | v_33457;
assign v_33461 = v_33459 | v_33460;
assign v_33463 = v_33240 | v_33462;
assign v_33466 = v_33464 | v_33465;
assign v_33468 = v_33237 | v_33467;
assign v_33471 = v_33469 | v_33470;
assign v_33473 = v_33471 | v_33472;
assign v_33476 = v_33234 | v_33475;
assign v_33547 = v_33544 | v_33546;
assign v_33549 = v_33542 | v_33548;
assign v_33551 = v_33540 | v_33550;
assign v_33553 = v_33548 | v_33552;
assign v_33555 = v_33538 | v_33554;
assign v_33557 = v_33536 | v_33556;
assign v_33559 = v_33554 | v_33558;
assign v_33561 = v_33534 | v_33560;
assign v_33563 = v_33532 | v_33562;
assign v_33565 = v_33560 | v_33564;
assign v_33567 = v_33530 | v_33566;
assign v_33569 = v_33528 | v_33568;
assign v_33571 = v_33566 | v_33570;
assign v_33573 = v_33526 | v_33572;
assign v_33575 = v_33524 | v_33574;
assign v_33577 = v_33572 | v_33576;
assign v_33579 = v_33522 | v_33578;
assign v_33581 = v_33520 | v_33580;
assign v_33583 = v_33578 | v_33582;
assign v_33585 = v_33518 | v_33584;
assign v_33587 = v_33516 | v_33586;
assign v_33589 = v_33584 | v_33588;
assign v_33591 = v_33514 | v_33590;
assign v_33593 = v_33512 | v_33592;
assign v_33595 = v_33590 | v_33594;
assign v_33597 = v_33510 | v_33596;
assign v_33599 = v_33508 | v_33598;
assign v_33601 = v_33596 | v_33600;
assign v_33603 = v_33506 | v_33602;
assign v_33605 = v_33504 | v_33604;
assign v_33607 = v_33602 | v_33606;
assign v_33609 = v_33502 | v_33608;
assign v_33611 = v_33500 | v_33610;
assign v_33613 = v_33608 | v_33612;
assign v_33615 = v_33498 | v_33614;
assign v_33617 = v_33496 | v_33616;
assign v_33619 = v_33614 | v_33618;
assign v_33621 = v_33494 | v_33620;
assign v_33623 = v_33491 | v_33622;
assign v_33625 = v_33620 | v_33624;
assign v_33627 = v_33490 | v_33626;
assign v_33629 = v_33487 | v_33628;
assign v_33631 = v_33626 | v_33630;
assign v_33633 = v_33486 | v_33632;
assign v_33635 = v_33483 | v_33634;
assign v_33637 = v_33632 | v_33636;
assign v_33639 = v_33482 | v_33638;
assign v_33641 = v_33479 | v_33640;
assign v_33643 = v_33638 | v_33642;
assign v_33646 = ~v_33478 | v_33645;
assign v_33653 = v_33542 | v_33652;
assign v_33656 = v_33654 | v_33655;
assign v_33658 = v_33538 | v_33657;
assign v_33661 = v_33659 | v_33660;
assign v_33663 = v_33534 | v_33662;
assign v_33666 = v_33664 | v_33665;
assign v_33668 = v_33530 | v_33667;
assign v_33671 = v_33669 | v_33670;
assign v_33673 = v_33526 | v_33672;
assign v_33676 = v_33674 | v_33675;
assign v_33678 = v_33522 | v_33677;
assign v_33681 = v_33679 | v_33680;
assign v_33683 = v_33518 | v_33682;
assign v_33686 = v_33684 | v_33685;
assign v_33688 = v_33514 | v_33687;
assign v_33691 = v_33689 | v_33690;
assign v_33693 = v_33510 | v_33692;
assign v_33696 = v_33694 | v_33695;
assign v_33698 = v_33506 | v_33697;
assign v_33701 = v_33699 | v_33700;
assign v_33703 = v_33502 | v_33702;
assign v_33706 = v_33704 | v_33705;
assign v_33708 = v_33498 | v_33707;
assign v_33711 = v_33709 | v_33710;
assign v_33713 = v_33494 | v_33712;
assign v_33716 = v_33714 | v_33715;
assign v_33718 = v_33490 | v_33717;
assign v_33721 = v_33719 | v_33720;
assign v_33723 = v_33486 | v_33722;
assign v_33726 = v_33724 | v_33725;
assign v_33728 = v_33482 | v_33727;
assign v_33731 = v_33729 | v_33730;
assign v_33733 = v_33478 | v_33732;
assign v_33736 = v_33477 | v_33735;
assign v_33790 = v_33787 | v_33789;
assign v_33792 = v_33786 | v_33791;
assign v_33794 = v_33784 | v_33793;
assign v_33796 = v_33791 | v_33795;
assign v_33798 = v_33783 | v_33797;
assign v_33800 = v_33781 | v_33799;
assign v_33802 = v_33797 | v_33801;
assign v_33804 = v_33780 | v_33803;
assign v_33806 = v_33778 | v_33805;
assign v_33808 = v_33803 | v_33807;
assign v_33810 = v_33777 | v_33809;
assign v_33812 = v_33775 | v_33811;
assign v_33814 = v_33809 | v_33813;
assign v_33816 = v_33774 | v_33815;
assign v_33818 = v_33772 | v_33817;
assign v_33820 = v_33815 | v_33819;
assign v_33822 = v_33771 | v_33821;
assign v_33824 = v_33769 | v_33823;
assign v_33826 = v_33821 | v_33825;
assign v_33828 = v_33768 | v_33827;
assign v_33830 = v_33766 | v_33829;
assign v_33832 = v_33827 | v_33831;
assign v_33834 = v_33765 | v_33833;
assign v_33836 = v_33763 | v_33835;
assign v_33838 = v_33833 | v_33837;
assign v_33840 = v_33762 | v_33839;
assign v_33842 = v_33760 | v_33841;
assign v_33844 = v_33839 | v_33843;
assign v_33846 = v_33759 | v_33845;
assign v_33848 = v_33757 | v_33847;
assign v_33850 = v_33845 | v_33849;
assign v_33852 = v_33756 | v_33851;
assign v_33854 = v_33754 | v_33853;
assign v_33856 = v_33851 | v_33855;
assign v_33858 = v_33753 | v_33857;
assign v_33860 = v_33751 | v_33859;
assign v_33862 = v_33857 | v_33861;
assign v_33864 = v_33750 | v_33863;
assign v_33866 = v_33748 | v_33865;
assign v_33868 = v_33863 | v_33867;
assign v_33870 = v_33747 | v_33869;
assign v_33872 = v_33745 | v_33871;
assign v_33874 = v_33869 | v_33873;
assign v_33876 = v_33744 | v_33875;
assign v_33878 = v_33742 | v_33877;
assign v_33880 = v_33875 | v_33879;
assign v_33882 = v_33741 | v_33881;
assign v_33884 = v_33739 | v_33883;
assign v_33886 = v_33881 | v_33885;
assign v_33889 = ~v_33738 | v_33888;
assign v_33896 = v_33786 | v_33895;
assign v_33899 = v_33897 | v_33898;
assign v_33901 = v_33783 | v_33900;
assign v_33904 = v_33902 | v_33903;
assign v_33906 = v_33780 | v_33905;
assign v_33909 = v_33907 | v_33908;
assign v_33911 = v_33777 | v_33910;
assign v_33914 = v_33912 | v_33913;
assign v_33916 = v_33774 | v_33915;
assign v_33919 = v_33917 | v_33918;
assign v_33921 = v_33771 | v_33920;
assign v_33924 = v_33922 | v_33923;
assign v_33926 = v_33768 | v_33925;
assign v_33929 = v_33927 | v_33928;
assign v_33931 = v_33765 | v_33930;
assign v_33934 = v_33932 | v_33933;
assign v_33936 = v_33762 | v_33935;
assign v_33939 = v_33937 | v_33938;
assign v_33941 = v_33759 | v_33940;
assign v_33944 = v_33942 | v_33943;
assign v_33946 = v_33756 | v_33945;
assign v_33949 = v_33947 | v_33948;
assign v_33951 = v_33753 | v_33950;
assign v_33954 = v_33952 | v_33953;
assign v_33956 = v_33750 | v_33955;
assign v_33959 = v_33957 | v_33958;
assign v_33961 = v_33747 | v_33960;
assign v_33964 = v_33962 | v_33963;
assign v_33966 = v_33744 | v_33965;
assign v_33969 = v_33967 | v_33968;
assign v_33971 = v_33741 | v_33970;
assign v_33974 = v_33972 | v_33973;
assign v_33976 = v_33738 | v_33975;
assign v_33979 = v_33737 | v_33978;
assign v_34033 = v_34030 | v_34032;
assign v_34035 = v_34029 | v_34034;
assign v_34037 = v_34027 | v_34036;
assign v_34039 = v_34034 | v_34038;
assign v_34041 = v_34026 | v_34040;
assign v_34043 = v_34024 | v_34042;
assign v_34045 = v_34040 | v_34044;
assign v_34047 = v_34023 | v_34046;
assign v_34049 = v_34021 | v_34048;
assign v_34051 = v_34046 | v_34050;
assign v_34053 = v_34020 | v_34052;
assign v_34055 = v_34018 | v_34054;
assign v_34057 = v_34052 | v_34056;
assign v_34059 = v_34017 | v_34058;
assign v_34061 = v_34015 | v_34060;
assign v_34063 = v_34058 | v_34062;
assign v_34065 = v_34014 | v_34064;
assign v_34067 = v_34012 | v_34066;
assign v_34069 = v_34064 | v_34068;
assign v_34071 = v_34011 | v_34070;
assign v_34073 = v_34009 | v_34072;
assign v_34075 = v_34070 | v_34074;
assign v_34077 = v_34008 | v_34076;
assign v_34079 = v_34006 | v_34078;
assign v_34081 = v_34076 | v_34080;
assign v_34083 = v_34005 | v_34082;
assign v_34085 = v_34003 | v_34084;
assign v_34087 = v_34082 | v_34086;
assign v_34089 = v_34002 | v_34088;
assign v_34091 = v_34000 | v_34090;
assign v_34093 = v_34088 | v_34092;
assign v_34095 = v_33999 | v_34094;
assign v_34097 = v_33997 | v_34096;
assign v_34099 = v_34094 | v_34098;
assign v_34101 = v_33996 | v_34100;
assign v_34103 = v_33994 | v_34102;
assign v_34105 = v_34100 | v_34104;
assign v_34107 = v_33993 | v_34106;
assign v_34109 = v_33991 | v_34108;
assign v_34111 = v_34106 | v_34110;
assign v_34113 = v_33990 | v_34112;
assign v_34115 = v_33988 | v_34114;
assign v_34117 = v_34112 | v_34116;
assign v_34119 = v_33987 | v_34118;
assign v_34121 = v_33985 | v_34120;
assign v_34123 = v_34118 | v_34122;
assign v_34125 = v_33984 | v_34124;
assign v_34127 = v_33982 | v_34126;
assign v_34129 = v_34124 | v_34128;
assign v_34132 = ~v_33981 | v_34131;
assign v_34139 = v_34029 | v_34138;
assign v_34142 = v_34140 | v_34141;
assign v_34144 = v_34026 | v_34143;
assign v_34147 = v_34145 | v_34146;
assign v_34149 = v_34023 | v_34148;
assign v_34152 = v_34150 | v_34151;
assign v_34154 = v_34020 | v_34153;
assign v_34157 = v_34155 | v_34156;
assign v_34159 = v_34017 | v_34158;
assign v_34162 = v_34160 | v_34161;
assign v_34164 = v_34014 | v_34163;
assign v_34167 = v_34165 | v_34166;
assign v_34169 = v_34011 | v_34168;
assign v_34172 = v_34170 | v_34171;
assign v_34174 = v_34008 | v_34173;
assign v_34177 = v_34175 | v_34176;
assign v_34179 = v_34005 | v_34178;
assign v_34182 = v_34180 | v_34181;
assign v_34184 = v_34002 | v_34183;
assign v_34187 = v_34185 | v_34186;
assign v_34189 = v_33999 | v_34188;
assign v_34192 = v_34190 | v_34191;
assign v_34194 = v_33996 | v_34193;
assign v_34197 = v_34195 | v_34196;
assign v_34199 = v_33993 | v_34198;
assign v_34202 = v_34200 | v_34201;
assign v_34204 = v_33990 | v_34203;
assign v_34207 = v_34205 | v_34206;
assign v_34209 = v_33987 | v_34208;
assign v_34212 = v_34210 | v_34211;
assign v_34214 = v_33984 | v_34213;
assign v_34217 = v_34215 | v_34216;
assign v_34219 = v_33981 | v_34218;
assign v_34222 = v_33980 | v_34221;
assign v_34276 = v_34273 | v_34275;
assign v_34278 = v_34272 | v_34277;
assign v_34280 = v_34270 | v_34279;
assign v_34282 = v_34277 | v_34281;
assign v_34284 = v_34269 | v_34283;
assign v_34286 = v_34267 | v_34285;
assign v_34288 = v_34283 | v_34287;
assign v_34290 = v_34266 | v_34289;
assign v_34292 = v_34264 | v_34291;
assign v_34294 = v_34289 | v_34293;
assign v_34296 = v_34263 | v_34295;
assign v_34298 = v_34261 | v_34297;
assign v_34300 = v_34295 | v_34299;
assign v_34302 = v_34260 | v_34301;
assign v_34304 = v_34258 | v_34303;
assign v_34306 = v_34301 | v_34305;
assign v_34308 = v_34257 | v_34307;
assign v_34310 = v_34255 | v_34309;
assign v_34312 = v_34307 | v_34311;
assign v_34314 = v_34254 | v_34313;
assign v_34316 = v_34252 | v_34315;
assign v_34318 = v_34313 | v_34317;
assign v_34320 = v_34251 | v_34319;
assign v_34322 = v_34249 | v_34321;
assign v_34324 = v_34319 | v_34323;
assign v_34326 = v_34248 | v_34325;
assign v_34328 = v_34246 | v_34327;
assign v_34330 = v_34325 | v_34329;
assign v_34332 = v_34245 | v_34331;
assign v_34334 = v_34243 | v_34333;
assign v_34336 = v_34331 | v_34335;
assign v_34338 = v_34242 | v_34337;
assign v_34340 = v_34240 | v_34339;
assign v_34342 = v_34337 | v_34341;
assign v_34344 = v_34239 | v_34343;
assign v_34346 = v_34237 | v_34345;
assign v_34348 = v_34343 | v_34347;
assign v_34350 = v_34236 | v_34349;
assign v_34352 = v_34234 | v_34351;
assign v_34354 = v_34349 | v_34353;
assign v_34356 = v_34233 | v_34355;
assign v_34358 = v_34231 | v_34357;
assign v_34360 = v_34355 | v_34359;
assign v_34362 = v_34230 | v_34361;
assign v_34364 = v_34228 | v_34363;
assign v_34366 = v_34361 | v_34365;
assign v_34368 = v_34227 | v_34367;
assign v_34370 = v_34225 | v_34369;
assign v_34372 = v_34367 | v_34371;
assign v_34375 = ~v_34224 | v_34374;
assign v_34382 = v_34272 | v_34381;
assign v_34385 = v_34383 | v_34384;
assign v_34387 = v_34269 | v_34386;
assign v_34390 = v_34388 | v_34389;
assign v_34392 = v_34266 | v_34391;
assign v_34395 = v_34393 | v_34394;
assign v_34397 = v_34263 | v_34396;
assign v_34400 = v_34398 | v_34399;
assign v_34402 = v_34260 | v_34401;
assign v_34405 = v_34403 | v_34404;
assign v_34407 = v_34257 | v_34406;
assign v_34410 = v_34408 | v_34409;
assign v_34412 = v_34254 | v_34411;
assign v_34415 = v_34413 | v_34414;
assign v_34417 = v_34251 | v_34416;
assign v_34420 = v_34418 | v_34419;
assign v_34422 = v_34248 | v_34421;
assign v_34425 = v_34423 | v_34424;
assign v_34427 = v_34245 | v_34426;
assign v_34430 = v_34428 | v_34429;
assign v_34432 = v_34242 | v_34431;
assign v_34435 = v_34433 | v_34434;
assign v_34437 = v_34239 | v_34436;
assign v_34440 = v_34438 | v_34439;
assign v_34442 = v_34236 | v_34441;
assign v_34445 = v_34443 | v_34444;
assign v_34447 = v_34233 | v_34446;
assign v_34450 = v_34448 | v_34449;
assign v_34452 = v_34230 | v_34451;
assign v_34455 = v_34453 | v_34454;
assign v_34457 = v_34227 | v_34456;
assign v_34460 = v_34458 | v_34459;
assign v_34462 = v_34224 | v_34461;
assign v_34465 = v_34223 | v_34464;
assign v_34519 = v_34516 | v_34518;
assign v_34521 = v_34515 | v_34520;
assign v_34523 = v_34513 | v_34522;
assign v_34525 = v_34520 | v_34524;
assign v_34527 = v_34512 | v_34526;
assign v_34529 = v_34510 | v_34528;
assign v_34531 = v_34526 | v_34530;
assign v_34533 = v_34509 | v_34532;
assign v_34535 = v_34507 | v_34534;
assign v_34537 = v_34532 | v_34536;
assign v_34539 = v_34506 | v_34538;
assign v_34541 = v_34504 | v_34540;
assign v_34543 = v_34538 | v_34542;
assign v_34545 = v_34503 | v_34544;
assign v_34547 = v_34501 | v_34546;
assign v_34549 = v_34544 | v_34548;
assign v_34551 = v_34500 | v_34550;
assign v_34553 = v_34498 | v_34552;
assign v_34555 = v_34550 | v_34554;
assign v_34557 = v_34497 | v_34556;
assign v_34559 = v_34495 | v_34558;
assign v_34561 = v_34556 | v_34560;
assign v_34563 = v_34494 | v_34562;
assign v_34565 = v_34492 | v_34564;
assign v_34567 = v_34562 | v_34566;
assign v_34569 = v_34491 | v_34568;
assign v_34571 = v_34489 | v_34570;
assign v_34573 = v_34568 | v_34572;
assign v_34575 = v_34488 | v_34574;
assign v_34577 = v_34486 | v_34576;
assign v_34579 = v_34574 | v_34578;
assign v_34581 = v_34485 | v_34580;
assign v_34583 = v_34483 | v_34582;
assign v_34585 = v_34580 | v_34584;
assign v_34587 = v_34482 | v_34586;
assign v_34589 = v_34480 | v_34588;
assign v_34591 = v_34586 | v_34590;
assign v_34593 = v_34479 | v_34592;
assign v_34595 = v_34477 | v_34594;
assign v_34597 = v_34592 | v_34596;
assign v_34599 = v_34476 | v_34598;
assign v_34601 = v_34474 | v_34600;
assign v_34603 = v_34598 | v_34602;
assign v_34605 = v_34473 | v_34604;
assign v_34607 = v_34471 | v_34606;
assign v_34609 = v_34604 | v_34608;
assign v_34611 = v_34470 | v_34610;
assign v_34613 = v_34468 | v_34612;
assign v_34615 = v_34610 | v_34614;
assign v_34618 = ~v_34467 | v_34617;
assign v_34625 = v_34515 | v_34624;
assign v_34628 = v_34626 | v_34627;
assign v_34630 = v_34512 | v_34629;
assign v_34633 = v_34631 | v_34632;
assign v_34635 = v_34509 | v_34634;
assign v_34638 = v_34636 | v_34637;
assign v_34640 = v_34506 | v_34639;
assign v_34643 = v_34641 | v_34642;
assign v_34645 = v_34503 | v_34644;
assign v_34648 = v_34646 | v_34647;
assign v_34650 = v_34500 | v_34649;
assign v_34653 = v_34651 | v_34652;
assign v_34655 = v_34497 | v_34654;
assign v_34658 = v_34656 | v_34657;
assign v_34660 = v_34494 | v_34659;
assign v_34663 = v_34661 | v_34662;
assign v_34665 = v_34491 | v_34664;
assign v_34668 = v_34666 | v_34667;
assign v_34670 = v_34488 | v_34669;
assign v_34673 = v_34671 | v_34672;
assign v_34675 = v_34485 | v_34674;
assign v_34678 = v_34676 | v_34677;
assign v_34680 = v_34482 | v_34679;
assign v_34683 = v_34681 | v_34682;
assign v_34685 = v_34479 | v_34684;
assign v_34688 = v_34686 | v_34687;
assign v_34690 = v_34476 | v_34689;
assign v_34693 = v_34691 | v_34692;
assign v_34695 = v_34473 | v_34694;
assign v_34698 = v_34696 | v_34697;
assign v_34700 = v_34470 | v_34699;
assign v_34703 = v_34701 | v_34702;
assign v_34705 = v_34467 | v_34704;
assign v_34708 = v_34466 | v_34707;
assign v_34762 = v_34759 | v_34761;
assign v_34764 = v_34758 | v_34763;
assign v_34766 = v_34756 | v_34765;
assign v_34768 = v_34763 | v_34767;
assign v_34770 = v_34755 | v_34769;
assign v_34772 = v_34753 | v_34771;
assign v_34774 = v_34769 | v_34773;
assign v_34776 = v_34752 | v_34775;
assign v_34778 = v_34750 | v_34777;
assign v_34780 = v_34775 | v_34779;
assign v_34782 = v_34749 | v_34781;
assign v_34784 = v_34747 | v_34783;
assign v_34786 = v_34781 | v_34785;
assign v_34788 = v_34746 | v_34787;
assign v_34790 = v_34744 | v_34789;
assign v_34792 = v_34787 | v_34791;
assign v_34794 = v_34743 | v_34793;
assign v_34796 = v_34741 | v_34795;
assign v_34798 = v_34793 | v_34797;
assign v_34800 = v_34740 | v_34799;
assign v_34802 = v_34738 | v_34801;
assign v_34804 = v_34799 | v_34803;
assign v_34806 = v_34737 | v_34805;
assign v_34808 = v_34735 | v_34807;
assign v_34810 = v_34805 | v_34809;
assign v_34812 = v_34734 | v_34811;
assign v_34814 = v_34732 | v_34813;
assign v_34816 = v_34811 | v_34815;
assign v_34818 = v_34731 | v_34817;
assign v_34820 = v_34729 | v_34819;
assign v_34822 = v_34817 | v_34821;
assign v_34824 = v_34728 | v_34823;
assign v_34826 = v_34726 | v_34825;
assign v_34828 = v_34823 | v_34827;
assign v_34830 = v_34725 | v_34829;
assign v_34832 = v_34723 | v_34831;
assign v_34834 = v_34829 | v_34833;
assign v_34836 = v_34722 | v_34835;
assign v_34838 = v_34720 | v_34837;
assign v_34840 = v_34835 | v_34839;
assign v_34842 = v_34719 | v_34841;
assign v_34844 = v_34717 | v_34843;
assign v_34846 = v_34841 | v_34845;
assign v_34848 = v_34716 | v_34847;
assign v_34850 = v_34714 | v_34849;
assign v_34852 = v_34847 | v_34851;
assign v_34854 = v_34713 | v_34853;
assign v_34856 = v_34711 | v_34855;
assign v_34858 = v_34853 | v_34857;
assign v_34861 = ~v_34710 | v_34860;
assign v_34868 = v_34758 | v_34867;
assign v_34871 = v_34869 | v_34870;
assign v_34873 = v_34755 | v_34872;
assign v_34876 = v_34874 | v_34875;
assign v_34878 = v_34752 | v_34877;
assign v_34881 = v_34879 | v_34880;
assign v_34883 = v_34749 | v_34882;
assign v_34886 = v_34884 | v_34885;
assign v_34888 = v_34746 | v_34887;
assign v_34891 = v_34889 | v_34890;
assign v_34893 = v_34743 | v_34892;
assign v_34896 = v_34894 | v_34895;
assign v_34898 = v_34740 | v_34897;
assign v_34901 = v_34899 | v_34900;
assign v_34903 = v_34737 | v_34902;
assign v_34906 = v_34904 | v_34905;
assign v_34908 = v_34734 | v_34907;
assign v_34911 = v_34909 | v_34910;
assign v_34913 = v_34731 | v_34912;
assign v_34916 = v_34914 | v_34915;
assign v_34918 = v_34728 | v_34917;
assign v_34921 = v_34919 | v_34920;
assign v_34923 = v_34725 | v_34922;
assign v_34926 = v_34924 | v_34925;
assign v_34928 = v_34722 | v_34927;
assign v_34931 = v_34929 | v_34930;
assign v_34933 = v_34719 | v_34932;
assign v_34936 = v_34934 | v_34935;
assign v_34938 = v_34716 | v_34937;
assign v_34941 = v_34939 | v_34940;
assign v_34943 = v_34713 | v_34942;
assign v_34946 = v_34944 | v_34945;
assign v_34948 = v_34710 | v_34947;
assign v_34951 = v_34709 | v_34950;
assign v_35005 = v_35002 | v_35004;
assign v_35007 = v_35001 | v_35006;
assign v_35009 = v_34999 | v_35008;
assign v_35011 = v_35006 | v_35010;
assign v_35013 = v_34998 | v_35012;
assign v_35015 = v_34996 | v_35014;
assign v_35017 = v_35012 | v_35016;
assign v_35019 = v_34995 | v_35018;
assign v_35021 = v_34993 | v_35020;
assign v_35023 = v_35018 | v_35022;
assign v_35025 = v_34992 | v_35024;
assign v_35027 = v_34990 | v_35026;
assign v_35029 = v_35024 | v_35028;
assign v_35031 = v_34989 | v_35030;
assign v_35033 = v_34987 | v_35032;
assign v_35035 = v_35030 | v_35034;
assign v_35037 = v_34986 | v_35036;
assign v_35039 = v_34984 | v_35038;
assign v_35041 = v_35036 | v_35040;
assign v_35043 = v_34983 | v_35042;
assign v_35045 = v_34981 | v_35044;
assign v_35047 = v_35042 | v_35046;
assign v_35049 = v_34980 | v_35048;
assign v_35051 = v_34978 | v_35050;
assign v_35053 = v_35048 | v_35052;
assign v_35055 = v_34977 | v_35054;
assign v_35057 = v_34975 | v_35056;
assign v_35059 = v_35054 | v_35058;
assign v_35061 = v_34974 | v_35060;
assign v_35063 = v_34972 | v_35062;
assign v_35065 = v_35060 | v_35064;
assign v_35067 = v_34971 | v_35066;
assign v_35069 = v_34969 | v_35068;
assign v_35071 = v_35066 | v_35070;
assign v_35073 = v_34968 | v_35072;
assign v_35075 = v_34966 | v_35074;
assign v_35077 = v_35072 | v_35076;
assign v_35079 = v_34965 | v_35078;
assign v_35081 = v_34963 | v_35080;
assign v_35083 = v_35078 | v_35082;
assign v_35085 = v_34962 | v_35084;
assign v_35087 = v_34960 | v_35086;
assign v_35089 = v_35084 | v_35088;
assign v_35091 = v_34959 | v_35090;
assign v_35093 = v_34957 | v_35092;
assign v_35095 = v_35090 | v_35094;
assign v_35097 = v_34956 | v_35096;
assign v_35099 = v_34954 | v_35098;
assign v_35101 = v_35096 | v_35100;
assign v_35104 = ~v_34953 | v_35103;
assign v_35111 = v_35001 | v_35110;
assign v_35114 = v_35112 | v_35113;
assign v_35116 = v_34998 | v_35115;
assign v_35119 = v_35117 | v_35118;
assign v_35121 = v_34995 | v_35120;
assign v_35124 = v_35122 | v_35123;
assign v_35126 = v_34992 | v_35125;
assign v_35129 = v_35127 | v_35128;
assign v_35131 = v_34989 | v_35130;
assign v_35134 = v_35132 | v_35133;
assign v_35136 = v_34986 | v_35135;
assign v_35139 = v_35137 | v_35138;
assign v_35141 = v_34983 | v_35140;
assign v_35144 = v_35142 | v_35143;
assign v_35146 = v_34980 | v_35145;
assign v_35149 = v_35147 | v_35148;
assign v_35151 = v_34977 | v_35150;
assign v_35154 = v_35152 | v_35153;
assign v_35156 = v_34974 | v_35155;
assign v_35159 = v_35157 | v_35158;
assign v_35161 = v_34971 | v_35160;
assign v_35164 = v_35162 | v_35163;
assign v_35166 = v_34968 | v_35165;
assign v_35169 = v_35167 | v_35168;
assign v_35171 = v_34965 | v_35170;
assign v_35174 = v_35172 | v_35173;
assign v_35176 = v_34962 | v_35175;
assign v_35179 = v_35177 | v_35178;
assign v_35181 = v_34959 | v_35180;
assign v_35184 = v_35182 | v_35183;
assign v_35186 = v_34956 | v_35185;
assign v_35189 = v_35187 | v_35188;
assign v_35191 = v_34953 | v_35190;
assign v_35194 = v_34952 | v_35193;
assign v_35248 = v_35245 | v_35247;
assign v_35250 = v_35244 | v_35249;
assign v_35252 = v_35242 | v_35251;
assign v_35254 = v_35249 | v_35253;
assign v_35256 = v_35241 | v_35255;
assign v_35258 = v_35239 | v_35257;
assign v_35260 = v_35255 | v_35259;
assign v_35262 = v_35238 | v_35261;
assign v_35264 = v_35236 | v_35263;
assign v_35266 = v_35261 | v_35265;
assign v_35268 = v_35235 | v_35267;
assign v_35270 = v_35233 | v_35269;
assign v_35272 = v_35267 | v_35271;
assign v_35274 = v_35232 | v_35273;
assign v_35276 = v_35230 | v_35275;
assign v_35278 = v_35273 | v_35277;
assign v_35280 = v_35229 | v_35279;
assign v_35282 = v_35227 | v_35281;
assign v_35284 = v_35279 | v_35283;
assign v_35286 = v_35226 | v_35285;
assign v_35288 = v_35224 | v_35287;
assign v_35290 = v_35285 | v_35289;
assign v_35292 = v_35223 | v_35291;
assign v_35294 = v_35221 | v_35293;
assign v_35296 = v_35291 | v_35295;
assign v_35298 = v_35220 | v_35297;
assign v_35300 = v_35218 | v_35299;
assign v_35302 = v_35297 | v_35301;
assign v_35304 = v_35217 | v_35303;
assign v_35306 = v_35215 | v_35305;
assign v_35308 = v_35303 | v_35307;
assign v_35310 = v_35214 | v_35309;
assign v_35312 = v_35212 | v_35311;
assign v_35314 = v_35309 | v_35313;
assign v_35316 = v_35211 | v_35315;
assign v_35318 = v_35209 | v_35317;
assign v_35320 = v_35315 | v_35319;
assign v_35322 = v_35208 | v_35321;
assign v_35324 = v_35206 | v_35323;
assign v_35326 = v_35321 | v_35325;
assign v_35328 = v_35205 | v_35327;
assign v_35330 = v_35203 | v_35329;
assign v_35332 = v_35327 | v_35331;
assign v_35334 = v_35202 | v_35333;
assign v_35336 = v_35200 | v_35335;
assign v_35338 = v_35333 | v_35337;
assign v_35340 = v_35199 | v_35339;
assign v_35342 = v_35197 | v_35341;
assign v_35344 = v_35339 | v_35343;
assign v_35347 = ~v_35196 | v_35346;
assign v_35354 = v_35244 | v_35353;
assign v_35357 = v_35355 | v_35356;
assign v_35359 = v_35241 | v_35358;
assign v_35362 = v_35360 | v_35361;
assign v_35364 = v_35238 | v_35363;
assign v_35367 = v_35365 | v_35366;
assign v_35369 = v_35235 | v_35368;
assign v_35372 = v_35370 | v_35371;
assign v_35374 = v_35232 | v_35373;
assign v_35377 = v_35375 | v_35376;
assign v_35379 = v_35229 | v_35378;
assign v_35382 = v_35380 | v_35381;
assign v_35384 = v_35226 | v_35383;
assign v_35387 = v_35385 | v_35386;
assign v_35389 = v_35223 | v_35388;
assign v_35392 = v_35390 | v_35391;
assign v_35394 = v_35220 | v_35393;
assign v_35397 = v_35395 | v_35396;
assign v_35399 = v_35217 | v_35398;
assign v_35402 = v_35400 | v_35401;
assign v_35404 = v_35214 | v_35403;
assign v_35407 = v_35405 | v_35406;
assign v_35409 = v_35211 | v_35408;
assign v_35412 = v_35410 | v_35411;
assign v_35414 = v_35208 | v_35413;
assign v_35417 = v_35415 | v_35416;
assign v_35419 = v_35205 | v_35418;
assign v_35422 = v_35420 | v_35421;
assign v_35424 = v_35202 | v_35423;
assign v_35427 = v_35425 | v_35426;
assign v_35429 = v_35199 | v_35428;
assign v_35432 = v_35430 | v_35431;
assign v_35434 = v_35196 | v_35433;
assign v_35437 = v_35195 | v_35436;
assign v_35491 = v_35488 | v_35490;
assign v_35493 = v_35487 | v_35492;
assign v_35495 = v_35485 | v_35494;
assign v_35497 = v_35492 | v_35496;
assign v_35499 = v_35484 | v_35498;
assign v_35501 = v_35482 | v_35500;
assign v_35503 = v_35498 | v_35502;
assign v_35505 = v_35481 | v_35504;
assign v_35507 = v_35479 | v_35506;
assign v_35509 = v_35504 | v_35508;
assign v_35511 = v_35478 | v_35510;
assign v_35513 = v_35476 | v_35512;
assign v_35515 = v_35510 | v_35514;
assign v_35517 = v_35475 | v_35516;
assign v_35519 = v_35473 | v_35518;
assign v_35521 = v_35516 | v_35520;
assign v_35523 = v_35472 | v_35522;
assign v_35525 = v_35470 | v_35524;
assign v_35527 = v_35522 | v_35526;
assign v_35529 = v_35469 | v_35528;
assign v_35531 = v_35467 | v_35530;
assign v_35533 = v_35528 | v_35532;
assign v_35535 = v_35466 | v_35534;
assign v_35537 = v_35464 | v_35536;
assign v_35539 = v_35534 | v_35538;
assign v_35541 = v_35463 | v_35540;
assign v_35543 = v_35461 | v_35542;
assign v_35545 = v_35540 | v_35544;
assign v_35547 = v_35460 | v_35546;
assign v_35549 = v_35458 | v_35548;
assign v_35551 = v_35546 | v_35550;
assign v_35553 = v_35457 | v_35552;
assign v_35555 = v_35455 | v_35554;
assign v_35557 = v_35552 | v_35556;
assign v_35559 = v_35454 | v_35558;
assign v_35561 = v_35452 | v_35560;
assign v_35563 = v_35558 | v_35562;
assign v_35565 = v_35451 | v_35564;
assign v_35567 = v_35449 | v_35566;
assign v_35569 = v_35564 | v_35568;
assign v_35571 = v_35448 | v_35570;
assign v_35573 = v_35446 | v_35572;
assign v_35575 = v_35570 | v_35574;
assign v_35577 = v_35445 | v_35576;
assign v_35579 = v_35443 | v_35578;
assign v_35581 = v_35576 | v_35580;
assign v_35583 = v_35442 | v_35582;
assign v_35585 = v_35440 | v_35584;
assign v_35587 = v_35582 | v_35586;
assign v_35590 = ~v_35439 | v_35589;
assign v_35597 = v_35487 | v_35596;
assign v_35600 = v_35598 | v_35599;
assign v_35602 = v_35484 | v_35601;
assign v_35605 = v_35603 | v_35604;
assign v_35607 = v_35481 | v_35606;
assign v_35610 = v_35608 | v_35609;
assign v_35612 = v_35478 | v_35611;
assign v_35615 = v_35613 | v_35614;
assign v_35617 = v_35475 | v_35616;
assign v_35620 = v_35618 | v_35619;
assign v_35622 = v_35472 | v_35621;
assign v_35625 = v_35623 | v_35624;
assign v_35627 = v_35469 | v_35626;
assign v_35630 = v_35628 | v_35629;
assign v_35632 = v_35466 | v_35631;
assign v_35635 = v_35633 | v_35634;
assign v_35637 = v_35463 | v_35636;
assign v_35640 = v_35638 | v_35639;
assign v_35642 = v_35460 | v_35641;
assign v_35645 = v_35643 | v_35644;
assign v_35647 = v_35457 | v_35646;
assign v_35650 = v_35648 | v_35649;
assign v_35652 = v_35454 | v_35651;
assign v_35655 = v_35653 | v_35654;
assign v_35657 = v_35451 | v_35656;
assign v_35660 = v_35658 | v_35659;
assign v_35662 = v_35448 | v_35661;
assign v_35665 = v_35663 | v_35664;
assign v_35667 = v_35445 | v_35666;
assign v_35670 = v_35668 | v_35669;
assign v_35672 = v_35442 | v_35671;
assign v_35675 = v_35673 | v_35674;
assign v_35677 = v_35439 | v_35676;
assign v_35680 = v_35438 | v_35679;
assign v_35734 = v_35731 | v_35733;
assign v_35736 = v_35730 | v_35735;
assign v_35738 = v_35728 | v_35737;
assign v_35740 = v_35735 | v_35739;
assign v_35742 = v_35727 | v_35741;
assign v_35744 = v_35725 | v_35743;
assign v_35746 = v_35741 | v_35745;
assign v_35748 = v_35724 | v_35747;
assign v_35750 = v_35722 | v_35749;
assign v_35752 = v_35747 | v_35751;
assign v_35754 = v_35721 | v_35753;
assign v_35756 = v_35719 | v_35755;
assign v_35758 = v_35753 | v_35757;
assign v_35760 = v_35718 | v_35759;
assign v_35762 = v_35716 | v_35761;
assign v_35764 = v_35759 | v_35763;
assign v_35766 = v_35715 | v_35765;
assign v_35768 = v_35713 | v_35767;
assign v_35770 = v_35765 | v_35769;
assign v_35772 = v_35712 | v_35771;
assign v_35774 = v_35710 | v_35773;
assign v_35776 = v_35771 | v_35775;
assign v_35778 = v_35709 | v_35777;
assign v_35780 = v_35707 | v_35779;
assign v_35782 = v_35777 | v_35781;
assign v_35784 = v_35706 | v_35783;
assign v_35786 = v_35704 | v_35785;
assign v_35788 = v_35783 | v_35787;
assign v_35790 = v_35703 | v_35789;
assign v_35792 = v_35701 | v_35791;
assign v_35794 = v_35789 | v_35793;
assign v_35796 = v_35700 | v_35795;
assign v_35798 = v_35698 | v_35797;
assign v_35800 = v_35795 | v_35799;
assign v_35802 = v_35697 | v_35801;
assign v_35804 = v_35695 | v_35803;
assign v_35806 = v_35801 | v_35805;
assign v_35808 = v_35694 | v_35807;
assign v_35810 = v_35692 | v_35809;
assign v_35812 = v_35807 | v_35811;
assign v_35814 = v_35691 | v_35813;
assign v_35816 = v_35689 | v_35815;
assign v_35818 = v_35813 | v_35817;
assign v_35820 = v_35688 | v_35819;
assign v_35822 = v_35686 | v_35821;
assign v_35824 = v_35819 | v_35823;
assign v_35826 = v_35685 | v_35825;
assign v_35828 = v_35683 | v_35827;
assign v_35830 = v_35825 | v_35829;
assign v_35833 = ~v_35682 | v_35832;
assign v_35840 = v_35730 | v_35839;
assign v_35843 = v_35841 | v_35842;
assign v_35845 = v_35727 | v_35844;
assign v_35848 = v_35846 | v_35847;
assign v_35850 = v_35724 | v_35849;
assign v_35853 = v_35851 | v_35852;
assign v_35855 = v_35721 | v_35854;
assign v_35858 = v_35856 | v_35857;
assign v_35860 = v_35718 | v_35859;
assign v_35863 = v_35861 | v_35862;
assign v_35865 = v_35715 | v_35864;
assign v_35868 = v_35866 | v_35867;
assign v_35870 = v_35712 | v_35869;
assign v_35873 = v_35871 | v_35872;
assign v_35875 = v_35709 | v_35874;
assign v_35878 = v_35876 | v_35877;
assign v_35880 = v_35706 | v_35879;
assign v_35883 = v_35881 | v_35882;
assign v_35885 = v_35703 | v_35884;
assign v_35888 = v_35886 | v_35887;
assign v_35890 = v_35700 | v_35889;
assign v_35893 = v_35891 | v_35892;
assign v_35895 = v_35697 | v_35894;
assign v_35898 = v_35896 | v_35897;
assign v_35900 = v_35694 | v_35899;
assign v_35903 = v_35901 | v_35902;
assign v_35905 = v_35691 | v_35904;
assign v_35908 = v_35906 | v_35907;
assign v_35910 = v_35688 | v_35909;
assign v_35913 = v_35911 | v_35912;
assign v_35915 = v_35685 | v_35914;
assign v_35918 = v_35916 | v_35917;
assign v_35920 = v_35682 | v_35919;
assign v_35923 = v_35681 | v_35922;
assign v_35977 = v_35974 | v_35976;
assign v_35979 = v_35973 | v_35978;
assign v_35981 = v_35971 | v_35980;
assign v_35983 = v_35978 | v_35982;
assign v_35985 = v_35970 | v_35984;
assign v_35987 = v_35968 | v_35986;
assign v_35989 = v_35984 | v_35988;
assign v_35991 = v_35967 | v_35990;
assign v_35993 = v_35965 | v_35992;
assign v_35995 = v_35990 | v_35994;
assign v_35997 = v_35964 | v_35996;
assign v_35999 = v_35962 | v_35998;
assign v_36001 = v_35996 | v_36000;
assign v_36003 = v_35961 | v_36002;
assign v_36005 = v_35959 | v_36004;
assign v_36007 = v_36002 | v_36006;
assign v_36009 = v_35958 | v_36008;
assign v_36011 = v_35956 | v_36010;
assign v_36013 = v_36008 | v_36012;
assign v_36015 = v_35955 | v_36014;
assign v_36017 = v_35953 | v_36016;
assign v_36019 = v_36014 | v_36018;
assign v_36021 = v_35952 | v_36020;
assign v_36023 = v_35950 | v_36022;
assign v_36025 = v_36020 | v_36024;
assign v_36027 = v_35949 | v_36026;
assign v_36029 = v_35947 | v_36028;
assign v_36031 = v_36026 | v_36030;
assign v_36033 = v_35946 | v_36032;
assign v_36035 = v_35944 | v_36034;
assign v_36037 = v_36032 | v_36036;
assign v_36039 = v_35943 | v_36038;
assign v_36041 = v_35941 | v_36040;
assign v_36043 = v_36038 | v_36042;
assign v_36045 = v_35940 | v_36044;
assign v_36047 = v_35938 | v_36046;
assign v_36049 = v_36044 | v_36048;
assign v_36051 = v_35937 | v_36050;
assign v_36053 = v_35935 | v_36052;
assign v_36055 = v_36050 | v_36054;
assign v_36057 = v_35934 | v_36056;
assign v_36059 = v_35932 | v_36058;
assign v_36061 = v_36056 | v_36060;
assign v_36063 = v_35931 | v_36062;
assign v_36065 = v_35929 | v_36064;
assign v_36067 = v_36062 | v_36066;
assign v_36069 = v_35928 | v_36068;
assign v_36071 = v_35926 | v_36070;
assign v_36073 = v_36068 | v_36072;
assign v_36076 = ~v_35925 | v_36075;
assign v_36083 = v_35973 | v_36082;
assign v_36086 = v_36084 | v_36085;
assign v_36088 = v_35970 | v_36087;
assign v_36091 = v_36089 | v_36090;
assign v_36093 = v_35967 | v_36092;
assign v_36096 = v_36094 | v_36095;
assign v_36098 = v_35964 | v_36097;
assign v_36101 = v_36099 | v_36100;
assign v_36103 = v_35961 | v_36102;
assign v_36106 = v_36104 | v_36105;
assign v_36108 = v_35958 | v_36107;
assign v_36111 = v_36109 | v_36110;
assign v_36113 = v_35955 | v_36112;
assign v_36116 = v_36114 | v_36115;
assign v_36118 = v_35952 | v_36117;
assign v_36121 = v_36119 | v_36120;
assign v_36123 = v_35949 | v_36122;
assign v_36126 = v_36124 | v_36125;
assign v_36128 = v_35946 | v_36127;
assign v_36131 = v_36129 | v_36130;
assign v_36133 = v_35943 | v_36132;
assign v_36136 = v_36134 | v_36135;
assign v_36138 = v_35940 | v_36137;
assign v_36141 = v_36139 | v_36140;
assign v_36143 = v_35937 | v_36142;
assign v_36146 = v_36144 | v_36145;
assign v_36148 = v_35934 | v_36147;
assign v_36151 = v_36149 | v_36150;
assign v_36153 = v_35931 | v_36152;
assign v_36156 = v_36154 | v_36155;
assign v_36158 = v_35928 | v_36157;
assign v_36161 = v_36159 | v_36160;
assign v_36163 = v_35925 | v_36162;
assign v_36166 = v_35924 | v_36165;
assign v_36220 = v_36217 | v_36219;
assign v_36222 = v_36216 | v_36221;
assign v_36224 = v_36214 | v_36223;
assign v_36226 = v_36221 | v_36225;
assign v_36228 = v_36213 | v_36227;
assign v_36230 = v_36211 | v_36229;
assign v_36232 = v_36227 | v_36231;
assign v_36234 = v_36210 | v_36233;
assign v_36236 = v_36208 | v_36235;
assign v_36238 = v_36233 | v_36237;
assign v_36240 = v_36207 | v_36239;
assign v_36242 = v_36205 | v_36241;
assign v_36244 = v_36239 | v_36243;
assign v_36246 = v_36204 | v_36245;
assign v_36248 = v_36202 | v_36247;
assign v_36250 = v_36245 | v_36249;
assign v_36252 = v_36201 | v_36251;
assign v_36254 = v_36199 | v_36253;
assign v_36256 = v_36251 | v_36255;
assign v_36258 = v_36198 | v_36257;
assign v_36260 = v_36196 | v_36259;
assign v_36262 = v_36257 | v_36261;
assign v_36264 = v_36195 | v_36263;
assign v_36266 = v_36193 | v_36265;
assign v_36268 = v_36263 | v_36267;
assign v_36270 = v_36192 | v_36269;
assign v_36272 = v_36190 | v_36271;
assign v_36274 = v_36269 | v_36273;
assign v_36276 = v_36189 | v_36275;
assign v_36278 = v_36187 | v_36277;
assign v_36280 = v_36275 | v_36279;
assign v_36282 = v_36186 | v_36281;
assign v_36284 = v_36184 | v_36283;
assign v_36286 = v_36281 | v_36285;
assign v_36288 = v_36183 | v_36287;
assign v_36290 = v_36181 | v_36289;
assign v_36292 = v_36287 | v_36291;
assign v_36294 = v_36180 | v_36293;
assign v_36296 = v_36178 | v_36295;
assign v_36298 = v_36293 | v_36297;
assign v_36300 = v_36177 | v_36299;
assign v_36302 = v_36175 | v_36301;
assign v_36304 = v_36299 | v_36303;
assign v_36306 = v_36174 | v_36305;
assign v_36308 = v_36172 | v_36307;
assign v_36310 = v_36305 | v_36309;
assign v_36312 = v_36171 | v_36311;
assign v_36314 = v_36169 | v_36313;
assign v_36316 = v_36311 | v_36315;
assign v_36319 = ~v_36168 | v_36318;
assign v_36326 = v_36216 | v_36325;
assign v_36329 = v_36327 | v_36328;
assign v_36331 = v_36213 | v_36330;
assign v_36334 = v_36332 | v_36333;
assign v_36336 = v_36210 | v_36335;
assign v_36339 = v_36337 | v_36338;
assign v_36341 = v_36207 | v_36340;
assign v_36344 = v_36342 | v_36343;
assign v_36346 = v_36204 | v_36345;
assign v_36349 = v_36347 | v_36348;
assign v_36351 = v_36201 | v_36350;
assign v_36354 = v_36352 | v_36353;
assign v_36356 = v_36198 | v_36355;
assign v_36359 = v_36357 | v_36358;
assign v_36361 = v_36195 | v_36360;
assign v_36364 = v_36362 | v_36363;
assign v_36366 = v_36192 | v_36365;
assign v_36369 = v_36367 | v_36368;
assign v_36371 = v_36189 | v_36370;
assign v_36374 = v_36372 | v_36373;
assign v_36376 = v_36186 | v_36375;
assign v_36379 = v_36377 | v_36378;
assign v_36381 = v_36183 | v_36380;
assign v_36384 = v_36382 | v_36383;
assign v_36386 = v_36180 | v_36385;
assign v_36389 = v_36387 | v_36388;
assign v_36391 = v_36177 | v_36390;
assign v_36394 = v_36392 | v_36393;
assign v_36396 = v_36174 | v_36395;
assign v_36399 = v_36397 | v_36398;
assign v_36401 = v_36171 | v_36400;
assign v_36404 = v_36402 | v_36403;
assign v_36406 = v_36168 | v_36405;
assign v_36409 = v_36167 | v_36408;
assign v_36463 = v_36460 | v_36462;
assign v_36465 = v_36459 | v_36464;
assign v_36467 = v_36457 | v_36466;
assign v_36469 = v_36464 | v_36468;
assign v_36471 = v_36456 | v_36470;
assign v_36473 = v_36454 | v_36472;
assign v_36475 = v_36470 | v_36474;
assign v_36477 = v_36453 | v_36476;
assign v_36479 = v_36451 | v_36478;
assign v_36481 = v_36476 | v_36480;
assign v_36483 = v_36450 | v_36482;
assign v_36485 = v_36448 | v_36484;
assign v_36487 = v_36482 | v_36486;
assign v_36489 = v_36447 | v_36488;
assign v_36491 = v_36445 | v_36490;
assign v_36493 = v_36488 | v_36492;
assign v_36495 = v_36444 | v_36494;
assign v_36497 = v_36442 | v_36496;
assign v_36499 = v_36494 | v_36498;
assign v_36501 = v_36441 | v_36500;
assign v_36503 = v_36439 | v_36502;
assign v_36505 = v_36500 | v_36504;
assign v_36507 = v_36438 | v_36506;
assign v_36509 = v_36436 | v_36508;
assign v_36511 = v_36506 | v_36510;
assign v_36513 = v_36435 | v_36512;
assign v_36515 = v_36433 | v_36514;
assign v_36517 = v_36512 | v_36516;
assign v_36519 = v_36432 | v_36518;
assign v_36521 = v_36430 | v_36520;
assign v_36523 = v_36518 | v_36522;
assign v_36525 = v_36429 | v_36524;
assign v_36527 = v_36427 | v_36526;
assign v_36529 = v_36524 | v_36528;
assign v_36531 = v_36426 | v_36530;
assign v_36533 = v_36424 | v_36532;
assign v_36535 = v_36530 | v_36534;
assign v_36537 = v_36423 | v_36536;
assign v_36539 = v_36421 | v_36538;
assign v_36541 = v_36536 | v_36540;
assign v_36543 = v_36420 | v_36542;
assign v_36545 = v_36418 | v_36544;
assign v_36547 = v_36542 | v_36546;
assign v_36549 = v_36417 | v_36548;
assign v_36551 = v_36415 | v_36550;
assign v_36553 = v_36548 | v_36552;
assign v_36555 = v_36414 | v_36554;
assign v_36557 = v_36412 | v_36556;
assign v_36559 = v_36554 | v_36558;
assign v_36562 = ~v_36411 | v_36561;
assign v_36569 = v_36459 | v_36568;
assign v_36572 = v_36570 | v_36571;
assign v_36574 = v_36456 | v_36573;
assign v_36577 = v_36575 | v_36576;
assign v_36579 = v_36453 | v_36578;
assign v_36582 = v_36580 | v_36581;
assign v_36584 = v_36450 | v_36583;
assign v_36587 = v_36585 | v_36586;
assign v_36589 = v_36447 | v_36588;
assign v_36592 = v_36590 | v_36591;
assign v_36594 = v_36444 | v_36593;
assign v_36597 = v_36595 | v_36596;
assign v_36599 = v_36441 | v_36598;
assign v_36602 = v_36600 | v_36601;
assign v_36604 = v_36438 | v_36603;
assign v_36607 = v_36605 | v_36606;
assign v_36609 = v_36435 | v_36608;
assign v_36612 = v_36610 | v_36611;
assign v_36614 = v_36432 | v_36613;
assign v_36617 = v_36615 | v_36616;
assign v_36619 = v_36429 | v_36618;
assign v_36622 = v_36620 | v_36621;
assign v_36624 = v_36426 | v_36623;
assign v_36627 = v_36625 | v_36626;
assign v_36629 = v_36423 | v_36628;
assign v_36632 = v_36630 | v_36631;
assign v_36634 = v_36420 | v_36633;
assign v_36637 = v_36635 | v_36636;
assign v_36639 = v_36417 | v_36638;
assign v_36642 = v_36640 | v_36641;
assign v_36644 = v_36414 | v_36643;
assign v_36647 = v_36645 | v_36646;
assign v_36649 = v_36411 | v_36648;
assign v_36652 = v_36410 | v_36651;
assign v_36706 = v_36703 | v_36705;
assign v_36708 = v_36702 | v_36707;
assign v_36710 = v_36700 | v_36709;
assign v_36712 = v_36707 | v_36711;
assign v_36714 = v_36699 | v_36713;
assign v_36716 = v_36697 | v_36715;
assign v_36718 = v_36713 | v_36717;
assign v_36720 = v_36696 | v_36719;
assign v_36722 = v_36694 | v_36721;
assign v_36724 = v_36719 | v_36723;
assign v_36726 = v_36693 | v_36725;
assign v_36728 = v_36691 | v_36727;
assign v_36730 = v_36725 | v_36729;
assign v_36732 = v_36690 | v_36731;
assign v_36734 = v_36688 | v_36733;
assign v_36736 = v_36731 | v_36735;
assign v_36738 = v_36687 | v_36737;
assign v_36740 = v_36685 | v_36739;
assign v_36742 = v_36737 | v_36741;
assign v_36744 = v_36684 | v_36743;
assign v_36746 = v_36682 | v_36745;
assign v_36748 = v_36743 | v_36747;
assign v_36750 = v_36681 | v_36749;
assign v_36752 = v_36679 | v_36751;
assign v_36754 = v_36749 | v_36753;
assign v_36756 = v_36678 | v_36755;
assign v_36758 = v_36676 | v_36757;
assign v_36760 = v_36755 | v_36759;
assign v_36762 = v_36675 | v_36761;
assign v_36764 = v_36673 | v_36763;
assign v_36766 = v_36761 | v_36765;
assign v_36768 = v_36672 | v_36767;
assign v_36770 = v_36670 | v_36769;
assign v_36772 = v_36767 | v_36771;
assign v_36774 = v_36669 | v_36773;
assign v_36776 = v_36667 | v_36775;
assign v_36778 = v_36773 | v_36777;
assign v_36780 = v_36666 | v_36779;
assign v_36782 = v_36664 | v_36781;
assign v_36784 = v_36779 | v_36783;
assign v_36786 = v_36663 | v_36785;
assign v_36788 = v_36661 | v_36787;
assign v_36790 = v_36785 | v_36789;
assign v_36792 = v_36660 | v_36791;
assign v_36794 = v_36658 | v_36793;
assign v_36796 = v_36791 | v_36795;
assign v_36798 = v_36657 | v_36797;
assign v_36800 = v_36655 | v_36799;
assign v_36802 = v_36797 | v_36801;
assign v_36805 = ~v_36654 | v_36804;
assign v_36812 = v_36702 | v_36811;
assign v_36815 = v_36813 | v_36814;
assign v_36817 = v_36699 | v_36816;
assign v_36820 = v_36818 | v_36819;
assign v_36822 = v_36696 | v_36821;
assign v_36825 = v_36823 | v_36824;
assign v_36827 = v_36693 | v_36826;
assign v_36830 = v_36828 | v_36829;
assign v_36832 = v_36690 | v_36831;
assign v_36835 = v_36833 | v_36834;
assign v_36837 = v_36687 | v_36836;
assign v_36840 = v_36838 | v_36839;
assign v_36842 = v_36684 | v_36841;
assign v_36845 = v_36843 | v_36844;
assign v_36847 = v_36681 | v_36846;
assign v_36850 = v_36848 | v_36849;
assign v_36852 = v_36678 | v_36851;
assign v_36855 = v_36853 | v_36854;
assign v_36857 = v_36675 | v_36856;
assign v_36860 = v_36858 | v_36859;
assign v_36862 = v_36672 | v_36861;
assign v_36865 = v_36863 | v_36864;
assign v_36867 = v_36669 | v_36866;
assign v_36870 = v_36868 | v_36869;
assign v_36872 = v_36666 | v_36871;
assign v_36875 = v_36873 | v_36874;
assign v_36877 = v_36663 | v_36876;
assign v_36880 = v_36878 | v_36879;
assign v_36882 = v_36660 | v_36881;
assign v_36885 = v_36883 | v_36884;
assign v_36887 = v_36657 | v_36886;
assign v_36890 = v_36888 | v_36889;
assign v_36892 = v_36654 | v_36891;
assign v_36895 = v_36653 | v_36894;
assign v_36949 = v_36946 | v_36948;
assign v_36951 = v_36945 | v_36950;
assign v_36953 = v_36943 | v_36952;
assign v_36955 = v_36950 | v_36954;
assign v_36957 = v_36942 | v_36956;
assign v_36959 = v_36940 | v_36958;
assign v_36961 = v_36956 | v_36960;
assign v_36963 = v_36939 | v_36962;
assign v_36965 = v_36937 | v_36964;
assign v_36967 = v_36962 | v_36966;
assign v_36969 = v_36936 | v_36968;
assign v_36971 = v_36934 | v_36970;
assign v_36973 = v_36968 | v_36972;
assign v_36975 = v_36933 | v_36974;
assign v_36977 = v_36931 | v_36976;
assign v_36979 = v_36974 | v_36978;
assign v_36981 = v_36930 | v_36980;
assign v_36983 = v_36928 | v_36982;
assign v_36985 = v_36980 | v_36984;
assign v_36987 = v_36927 | v_36986;
assign v_36989 = v_36925 | v_36988;
assign v_36991 = v_36986 | v_36990;
assign v_36993 = v_36924 | v_36992;
assign v_36995 = v_36922 | v_36994;
assign v_36997 = v_36992 | v_36996;
assign v_36999 = v_36921 | v_36998;
assign v_37001 = v_36919 | v_37000;
assign v_37003 = v_36998 | v_37002;
assign v_37005 = v_36918 | v_37004;
assign v_37007 = v_36916 | v_37006;
assign v_37009 = v_37004 | v_37008;
assign v_37011 = v_36915 | v_37010;
assign v_37013 = v_36913 | v_37012;
assign v_37015 = v_37010 | v_37014;
assign v_37017 = v_36912 | v_37016;
assign v_37019 = v_36910 | v_37018;
assign v_37021 = v_37016 | v_37020;
assign v_37023 = v_36909 | v_37022;
assign v_37025 = v_36907 | v_37024;
assign v_37027 = v_37022 | v_37026;
assign v_37029 = v_36906 | v_37028;
assign v_37031 = v_36904 | v_37030;
assign v_37033 = v_37028 | v_37032;
assign v_37035 = v_36903 | v_37034;
assign v_37037 = v_36901 | v_37036;
assign v_37039 = v_37034 | v_37038;
assign v_37041 = v_36900 | v_37040;
assign v_37043 = v_36898 | v_37042;
assign v_37045 = v_37040 | v_37044;
assign v_37048 = ~v_36897 | v_37047;
assign v_37055 = v_36945 | v_37054;
assign v_37058 = v_37056 | v_37057;
assign v_37060 = v_36942 | v_37059;
assign v_37063 = v_37061 | v_37062;
assign v_37065 = v_36939 | v_37064;
assign v_37068 = v_37066 | v_37067;
assign v_37070 = v_36936 | v_37069;
assign v_37073 = v_37071 | v_37072;
assign v_37075 = v_36933 | v_37074;
assign v_37078 = v_37076 | v_37077;
assign v_37080 = v_36930 | v_37079;
assign v_37083 = v_37081 | v_37082;
assign v_37085 = v_36927 | v_37084;
assign v_37088 = v_37086 | v_37087;
assign v_37090 = v_36924 | v_37089;
assign v_37093 = v_37091 | v_37092;
assign v_37095 = v_36921 | v_37094;
assign v_37098 = v_37096 | v_37097;
assign v_37100 = v_36918 | v_37099;
assign v_37103 = v_37101 | v_37102;
assign v_37105 = v_36915 | v_37104;
assign v_37108 = v_37106 | v_37107;
assign v_37110 = v_36912 | v_37109;
assign v_37113 = v_37111 | v_37112;
assign v_37115 = v_36909 | v_37114;
assign v_37118 = v_37116 | v_37117;
assign v_37120 = v_36906 | v_37119;
assign v_37123 = v_37121 | v_37122;
assign v_37125 = v_36903 | v_37124;
assign v_37128 = v_37126 | v_37127;
assign v_37130 = v_36900 | v_37129;
assign v_37133 = v_37131 | v_37132;
assign v_37135 = v_36897 | v_37134;
assign v_37138 = v_36896 | v_37137;
assign v_37192 = v_37189 | v_37191;
assign v_37194 = v_37188 | v_37193;
assign v_37196 = v_37186 | v_37195;
assign v_37198 = v_37193 | v_37197;
assign v_37200 = v_37185 | v_37199;
assign v_37202 = v_37183 | v_37201;
assign v_37204 = v_37199 | v_37203;
assign v_37206 = v_37182 | v_37205;
assign v_37208 = v_37180 | v_37207;
assign v_37210 = v_37205 | v_37209;
assign v_37212 = v_37179 | v_37211;
assign v_37214 = v_37177 | v_37213;
assign v_37216 = v_37211 | v_37215;
assign v_37218 = v_37176 | v_37217;
assign v_37220 = v_37174 | v_37219;
assign v_37222 = v_37217 | v_37221;
assign v_37224 = v_37173 | v_37223;
assign v_37226 = v_37171 | v_37225;
assign v_37228 = v_37223 | v_37227;
assign v_37230 = v_37170 | v_37229;
assign v_37232 = v_37168 | v_37231;
assign v_37234 = v_37229 | v_37233;
assign v_37236 = v_37167 | v_37235;
assign v_37238 = v_37165 | v_37237;
assign v_37240 = v_37235 | v_37239;
assign v_37242 = v_37164 | v_37241;
assign v_37244 = v_37162 | v_37243;
assign v_37246 = v_37241 | v_37245;
assign v_37248 = v_37161 | v_37247;
assign v_37250 = v_37159 | v_37249;
assign v_37252 = v_37247 | v_37251;
assign v_37254 = v_37158 | v_37253;
assign v_37256 = v_37156 | v_37255;
assign v_37258 = v_37253 | v_37257;
assign v_37260 = v_37155 | v_37259;
assign v_37262 = v_37153 | v_37261;
assign v_37264 = v_37259 | v_37263;
assign v_37266 = v_37152 | v_37265;
assign v_37268 = v_37150 | v_37267;
assign v_37270 = v_37265 | v_37269;
assign v_37272 = v_37149 | v_37271;
assign v_37274 = v_37147 | v_37273;
assign v_37276 = v_37271 | v_37275;
assign v_37278 = v_37146 | v_37277;
assign v_37280 = v_37144 | v_37279;
assign v_37282 = v_37277 | v_37281;
assign v_37284 = v_37143 | v_37283;
assign v_37286 = v_37141 | v_37285;
assign v_37288 = v_37283 | v_37287;
assign v_37291 = ~v_37140 | v_37290;
assign v_37298 = v_37188 | v_37297;
assign v_37301 = v_37299 | v_37300;
assign v_37303 = v_37185 | v_37302;
assign v_37306 = v_37304 | v_37305;
assign v_37308 = v_37182 | v_37307;
assign v_37311 = v_37309 | v_37310;
assign v_37313 = v_37179 | v_37312;
assign v_37316 = v_37314 | v_37315;
assign v_37318 = v_37176 | v_37317;
assign v_37321 = v_37319 | v_37320;
assign v_37323 = v_37173 | v_37322;
assign v_37326 = v_37324 | v_37325;
assign v_37328 = v_37170 | v_37327;
assign v_37331 = v_37329 | v_37330;
assign v_37333 = v_37167 | v_37332;
assign v_37336 = v_37334 | v_37335;
assign v_37338 = v_37164 | v_37337;
assign v_37341 = v_37339 | v_37340;
assign v_37343 = v_37161 | v_37342;
assign v_37346 = v_37344 | v_37345;
assign v_37348 = v_37158 | v_37347;
assign v_37351 = v_37349 | v_37350;
assign v_37353 = v_37155 | v_37352;
assign v_37356 = v_37354 | v_37355;
assign v_37358 = v_37152 | v_37357;
assign v_37361 = v_37359 | v_37360;
assign v_37363 = v_37149 | v_37362;
assign v_37366 = v_37364 | v_37365;
assign v_37368 = v_37146 | v_37367;
assign v_37371 = v_37369 | v_37370;
assign v_37373 = v_37143 | v_37372;
assign v_37376 = v_37374 | v_37375;
assign v_37378 = v_37140 | v_37377;
assign v_37381 = v_37139 | v_37380;
assign v_37434 = v_37431 | v_37433;
assign v_37436 = v_37430 | v_37435;
assign v_37438 = v_37428 | v_37437;
assign v_37440 = v_37435 | v_37439;
assign v_37442 = v_37427 | v_37441;
assign v_37444 = v_37425 | v_37443;
assign v_37446 = v_37441 | v_37445;
assign v_37448 = v_37424 | v_37447;
assign v_37450 = v_37422 | v_37449;
assign v_37452 = v_37447 | v_37451;
assign v_37454 = v_37421 | v_37453;
assign v_37456 = v_37419 | v_37455;
assign v_37458 = v_37453 | v_37457;
assign v_37460 = v_37418 | v_37459;
assign v_37462 = v_37416 | v_37461;
assign v_37464 = v_37459 | v_37463;
assign v_37466 = v_37415 | v_37465;
assign v_37468 = v_37413 | v_37467;
assign v_37470 = v_37465 | v_37469;
assign v_37472 = v_37412 | v_37471;
assign v_37474 = v_37410 | v_37473;
assign v_37476 = v_37471 | v_37475;
assign v_37478 = v_37409 | v_37477;
assign v_37480 = v_37407 | v_37479;
assign v_37482 = v_37477 | v_37481;
assign v_37484 = v_37406 | v_37483;
assign v_37486 = v_37404 | v_37485;
assign v_37488 = v_37483 | v_37487;
assign v_37490 = v_37403 | v_37489;
assign v_37492 = v_37401 | v_37491;
assign v_37494 = v_37489 | v_37493;
assign v_37496 = v_37400 | v_37495;
assign v_37498 = v_37398 | v_37497;
assign v_37500 = v_37495 | v_37499;
assign v_37502 = v_37397 | v_37501;
assign v_37504 = v_37395 | v_37503;
assign v_37506 = v_37501 | v_37505;
assign v_37508 = v_37394 | v_37507;
assign v_37510 = v_37392 | v_37509;
assign v_37512 = v_37507 | v_37511;
assign v_37514 = v_37391 | v_37513;
assign v_37516 = v_37389 | v_37515;
assign v_37518 = v_37513 | v_37517;
assign v_37520 = v_37388 | v_37519;
assign v_37522 = v_37386 | v_37521;
assign v_37524 = v_37519 | v_37523;
assign v_37526 = v_37385 | v_37525;
assign v_37528 = v_37383 | v_37527;
assign v_37530 = v_37525 | v_37529;
assign v_37534 = v_37531 | v_37533;
assign v_37541 = v_37430 | v_37540;
assign v_37544 = v_37542 | v_37543;
assign v_37546 = v_37427 | v_37545;
assign v_37549 = v_37547 | v_37548;
assign v_37551 = v_37424 | v_37550;
assign v_37554 = v_37552 | v_37553;
assign v_37556 = v_37421 | v_37555;
assign v_37559 = v_37557 | v_37558;
assign v_37561 = v_37418 | v_37560;
assign v_37564 = v_37562 | v_37563;
assign v_37566 = v_37415 | v_37565;
assign v_37569 = v_37567 | v_37568;
assign v_37571 = v_37412 | v_37570;
assign v_37574 = v_37572 | v_37573;
assign v_37576 = v_37409 | v_37575;
assign v_37579 = v_37577 | v_37578;
assign v_37581 = v_37406 | v_37580;
assign v_37584 = v_37582 | v_37583;
assign v_37586 = v_37403 | v_37585;
assign v_37589 = v_37587 | v_37588;
assign v_37591 = v_37400 | v_37590;
assign v_37594 = v_37592 | v_37593;
assign v_37596 = v_37397 | v_37595;
assign v_37599 = v_37597 | v_37598;
assign v_37601 = v_37394 | v_37600;
assign v_37604 = v_37602 | v_37603;
assign v_37606 = v_37391 | v_37605;
assign v_37609 = v_37607 | v_37608;
assign v_37611 = v_37388 | v_37610;
assign v_37614 = v_37612 | v_37613;
assign v_37616 = v_37385 | v_37615;
assign v_37619 = v_37617 | v_37618;
assign v_37621 = v_37619 | v_37620;
assign v_37624 = v_37382 | v_37623;
assign v_37695 = v_37692 | v_37694;
assign v_37697 = v_37690 | v_37696;
assign v_37699 = v_37688 | v_37698;
assign v_37701 = v_37696 | v_37700;
assign v_37703 = v_37686 | v_37702;
assign v_37705 = v_37684 | v_37704;
assign v_37707 = v_37702 | v_37706;
assign v_37709 = v_37682 | v_37708;
assign v_37711 = v_37680 | v_37710;
assign v_37713 = v_37708 | v_37712;
assign v_37715 = v_37678 | v_37714;
assign v_37717 = v_37676 | v_37716;
assign v_37719 = v_37714 | v_37718;
assign v_37721 = v_37674 | v_37720;
assign v_37723 = v_37672 | v_37722;
assign v_37725 = v_37720 | v_37724;
assign v_37727 = v_37670 | v_37726;
assign v_37729 = v_37668 | v_37728;
assign v_37731 = v_37726 | v_37730;
assign v_37733 = v_37666 | v_37732;
assign v_37735 = v_37664 | v_37734;
assign v_37737 = v_37732 | v_37736;
assign v_37739 = v_37662 | v_37738;
assign v_37741 = v_37660 | v_37740;
assign v_37743 = v_37738 | v_37742;
assign v_37745 = v_37658 | v_37744;
assign v_37747 = v_37656 | v_37746;
assign v_37749 = v_37744 | v_37748;
assign v_37751 = v_37654 | v_37750;
assign v_37753 = v_37652 | v_37752;
assign v_37755 = v_37750 | v_37754;
assign v_37757 = v_37650 | v_37756;
assign v_37759 = v_37648 | v_37758;
assign v_37761 = v_37756 | v_37760;
assign v_37763 = v_37646 | v_37762;
assign v_37765 = v_37644 | v_37764;
assign v_37767 = v_37762 | v_37766;
assign v_37769 = v_37642 | v_37768;
assign v_37771 = v_37639 | v_37770;
assign v_37773 = v_37768 | v_37772;
assign v_37775 = v_37638 | v_37774;
assign v_37777 = v_37635 | v_37776;
assign v_37779 = v_37774 | v_37778;
assign v_37781 = v_37634 | v_37780;
assign v_37783 = v_37631 | v_37782;
assign v_37785 = v_37780 | v_37784;
assign v_37787 = v_37630 | v_37786;
assign v_37789 = v_37627 | v_37788;
assign v_37791 = v_37786 | v_37790;
assign v_37794 = ~v_37626 | v_37793;
assign v_37801 = v_37690 | v_37800;
assign v_37804 = v_37802 | v_37803;
assign v_37806 = v_37686 | v_37805;
assign v_37809 = v_37807 | v_37808;
assign v_37811 = v_37682 | v_37810;
assign v_37814 = v_37812 | v_37813;
assign v_37816 = v_37678 | v_37815;
assign v_37819 = v_37817 | v_37818;
assign v_37821 = v_37674 | v_37820;
assign v_37824 = v_37822 | v_37823;
assign v_37826 = v_37670 | v_37825;
assign v_37829 = v_37827 | v_37828;
assign v_37831 = v_37666 | v_37830;
assign v_37834 = v_37832 | v_37833;
assign v_37836 = v_37662 | v_37835;
assign v_37839 = v_37837 | v_37838;
assign v_37841 = v_37658 | v_37840;
assign v_37844 = v_37842 | v_37843;
assign v_37846 = v_37654 | v_37845;
assign v_37849 = v_37847 | v_37848;
assign v_37851 = v_37650 | v_37850;
assign v_37854 = v_37852 | v_37853;
assign v_37856 = v_37646 | v_37855;
assign v_37859 = v_37857 | v_37858;
assign v_37861 = v_37642 | v_37860;
assign v_37864 = v_37862 | v_37863;
assign v_37866 = v_37638 | v_37865;
assign v_37869 = v_37867 | v_37868;
assign v_37871 = v_37634 | v_37870;
assign v_37874 = v_37872 | v_37873;
assign v_37876 = v_37630 | v_37875;
assign v_37879 = v_37877 | v_37878;
assign v_37881 = v_37626 | v_37880;
assign v_37884 = v_37625 | v_37883;
assign v_37938 = v_37935 | v_37937;
assign v_37940 = v_37934 | v_37939;
assign v_37942 = v_37932 | v_37941;
assign v_37944 = v_37939 | v_37943;
assign v_37946 = v_37931 | v_37945;
assign v_37948 = v_37929 | v_37947;
assign v_37950 = v_37945 | v_37949;
assign v_37952 = v_37928 | v_37951;
assign v_37954 = v_37926 | v_37953;
assign v_37956 = v_37951 | v_37955;
assign v_37958 = v_37925 | v_37957;
assign v_37960 = v_37923 | v_37959;
assign v_37962 = v_37957 | v_37961;
assign v_37964 = v_37922 | v_37963;
assign v_37966 = v_37920 | v_37965;
assign v_37968 = v_37963 | v_37967;
assign v_37970 = v_37919 | v_37969;
assign v_37972 = v_37917 | v_37971;
assign v_37974 = v_37969 | v_37973;
assign v_37976 = v_37916 | v_37975;
assign v_37978 = v_37914 | v_37977;
assign v_37980 = v_37975 | v_37979;
assign v_37982 = v_37913 | v_37981;
assign v_37984 = v_37911 | v_37983;
assign v_37986 = v_37981 | v_37985;
assign v_37988 = v_37910 | v_37987;
assign v_37990 = v_37908 | v_37989;
assign v_37992 = v_37987 | v_37991;
assign v_37994 = v_37907 | v_37993;
assign v_37996 = v_37905 | v_37995;
assign v_37998 = v_37993 | v_37997;
assign v_38000 = v_37904 | v_37999;
assign v_38002 = v_37902 | v_38001;
assign v_38004 = v_37999 | v_38003;
assign v_38006 = v_37901 | v_38005;
assign v_38008 = v_37899 | v_38007;
assign v_38010 = v_38005 | v_38009;
assign v_38012 = v_37898 | v_38011;
assign v_38014 = v_37896 | v_38013;
assign v_38016 = v_38011 | v_38015;
assign v_38018 = v_37895 | v_38017;
assign v_38020 = v_37893 | v_38019;
assign v_38022 = v_38017 | v_38021;
assign v_38024 = v_37892 | v_38023;
assign v_38026 = v_37890 | v_38025;
assign v_38028 = v_38023 | v_38027;
assign v_38030 = v_37889 | v_38029;
assign v_38032 = v_37887 | v_38031;
assign v_38034 = v_38029 | v_38033;
assign v_38037 = ~v_37886 | v_38036;
assign v_38044 = v_37934 | v_38043;
assign v_38047 = v_38045 | v_38046;
assign v_38049 = v_37931 | v_38048;
assign v_38052 = v_38050 | v_38051;
assign v_38054 = v_37928 | v_38053;
assign v_38057 = v_38055 | v_38056;
assign v_38059 = v_37925 | v_38058;
assign v_38062 = v_38060 | v_38061;
assign v_38064 = v_37922 | v_38063;
assign v_38067 = v_38065 | v_38066;
assign v_38069 = v_37919 | v_38068;
assign v_38072 = v_38070 | v_38071;
assign v_38074 = v_37916 | v_38073;
assign v_38077 = v_38075 | v_38076;
assign v_38079 = v_37913 | v_38078;
assign v_38082 = v_38080 | v_38081;
assign v_38084 = v_37910 | v_38083;
assign v_38087 = v_38085 | v_38086;
assign v_38089 = v_37907 | v_38088;
assign v_38092 = v_38090 | v_38091;
assign v_38094 = v_37904 | v_38093;
assign v_38097 = v_38095 | v_38096;
assign v_38099 = v_37901 | v_38098;
assign v_38102 = v_38100 | v_38101;
assign v_38104 = v_37898 | v_38103;
assign v_38107 = v_38105 | v_38106;
assign v_38109 = v_37895 | v_38108;
assign v_38112 = v_38110 | v_38111;
assign v_38114 = v_37892 | v_38113;
assign v_38117 = v_38115 | v_38116;
assign v_38119 = v_37889 | v_38118;
assign v_38122 = v_38120 | v_38121;
assign v_38124 = v_37886 | v_38123;
assign v_38127 = v_37885 | v_38126;
assign v_38181 = v_38178 | v_38180;
assign v_38183 = v_38177 | v_38182;
assign v_38185 = v_38175 | v_38184;
assign v_38187 = v_38182 | v_38186;
assign v_38189 = v_38174 | v_38188;
assign v_38191 = v_38172 | v_38190;
assign v_38193 = v_38188 | v_38192;
assign v_38195 = v_38171 | v_38194;
assign v_38197 = v_38169 | v_38196;
assign v_38199 = v_38194 | v_38198;
assign v_38201 = v_38168 | v_38200;
assign v_38203 = v_38166 | v_38202;
assign v_38205 = v_38200 | v_38204;
assign v_38207 = v_38165 | v_38206;
assign v_38209 = v_38163 | v_38208;
assign v_38211 = v_38206 | v_38210;
assign v_38213 = v_38162 | v_38212;
assign v_38215 = v_38160 | v_38214;
assign v_38217 = v_38212 | v_38216;
assign v_38219 = v_38159 | v_38218;
assign v_38221 = v_38157 | v_38220;
assign v_38223 = v_38218 | v_38222;
assign v_38225 = v_38156 | v_38224;
assign v_38227 = v_38154 | v_38226;
assign v_38229 = v_38224 | v_38228;
assign v_38231 = v_38153 | v_38230;
assign v_38233 = v_38151 | v_38232;
assign v_38235 = v_38230 | v_38234;
assign v_38237 = v_38150 | v_38236;
assign v_38239 = v_38148 | v_38238;
assign v_38241 = v_38236 | v_38240;
assign v_38243 = v_38147 | v_38242;
assign v_38245 = v_38145 | v_38244;
assign v_38247 = v_38242 | v_38246;
assign v_38249 = v_38144 | v_38248;
assign v_38251 = v_38142 | v_38250;
assign v_38253 = v_38248 | v_38252;
assign v_38255 = v_38141 | v_38254;
assign v_38257 = v_38139 | v_38256;
assign v_38259 = v_38254 | v_38258;
assign v_38261 = v_38138 | v_38260;
assign v_38263 = v_38136 | v_38262;
assign v_38265 = v_38260 | v_38264;
assign v_38267 = v_38135 | v_38266;
assign v_38269 = v_38133 | v_38268;
assign v_38271 = v_38266 | v_38270;
assign v_38273 = v_38132 | v_38272;
assign v_38275 = v_38130 | v_38274;
assign v_38277 = v_38272 | v_38276;
assign v_38280 = ~v_38129 | v_38279;
assign v_38287 = v_38177 | v_38286;
assign v_38290 = v_38288 | v_38289;
assign v_38292 = v_38174 | v_38291;
assign v_38295 = v_38293 | v_38294;
assign v_38297 = v_38171 | v_38296;
assign v_38300 = v_38298 | v_38299;
assign v_38302 = v_38168 | v_38301;
assign v_38305 = v_38303 | v_38304;
assign v_38307 = v_38165 | v_38306;
assign v_38310 = v_38308 | v_38309;
assign v_38312 = v_38162 | v_38311;
assign v_38315 = v_38313 | v_38314;
assign v_38317 = v_38159 | v_38316;
assign v_38320 = v_38318 | v_38319;
assign v_38322 = v_38156 | v_38321;
assign v_38325 = v_38323 | v_38324;
assign v_38327 = v_38153 | v_38326;
assign v_38330 = v_38328 | v_38329;
assign v_38332 = v_38150 | v_38331;
assign v_38335 = v_38333 | v_38334;
assign v_38337 = v_38147 | v_38336;
assign v_38340 = v_38338 | v_38339;
assign v_38342 = v_38144 | v_38341;
assign v_38345 = v_38343 | v_38344;
assign v_38347 = v_38141 | v_38346;
assign v_38350 = v_38348 | v_38349;
assign v_38352 = v_38138 | v_38351;
assign v_38355 = v_38353 | v_38354;
assign v_38357 = v_38135 | v_38356;
assign v_38360 = v_38358 | v_38359;
assign v_38362 = v_38132 | v_38361;
assign v_38365 = v_38363 | v_38364;
assign v_38367 = v_38129 | v_38366;
assign v_38370 = v_38128 | v_38369;
assign v_38424 = v_38421 | v_38423;
assign v_38426 = v_38420 | v_38425;
assign v_38428 = v_38418 | v_38427;
assign v_38430 = v_38425 | v_38429;
assign v_38432 = v_38417 | v_38431;
assign v_38434 = v_38415 | v_38433;
assign v_38436 = v_38431 | v_38435;
assign v_38438 = v_38414 | v_38437;
assign v_38440 = v_38412 | v_38439;
assign v_38442 = v_38437 | v_38441;
assign v_38444 = v_38411 | v_38443;
assign v_38446 = v_38409 | v_38445;
assign v_38448 = v_38443 | v_38447;
assign v_38450 = v_38408 | v_38449;
assign v_38452 = v_38406 | v_38451;
assign v_38454 = v_38449 | v_38453;
assign v_38456 = v_38405 | v_38455;
assign v_38458 = v_38403 | v_38457;
assign v_38460 = v_38455 | v_38459;
assign v_38462 = v_38402 | v_38461;
assign v_38464 = v_38400 | v_38463;
assign v_38466 = v_38461 | v_38465;
assign v_38468 = v_38399 | v_38467;
assign v_38470 = v_38397 | v_38469;
assign v_38472 = v_38467 | v_38471;
assign v_38474 = v_38396 | v_38473;
assign v_38476 = v_38394 | v_38475;
assign v_38478 = v_38473 | v_38477;
assign v_38480 = v_38393 | v_38479;
assign v_38482 = v_38391 | v_38481;
assign v_38484 = v_38479 | v_38483;
assign v_38486 = v_38390 | v_38485;
assign v_38488 = v_38388 | v_38487;
assign v_38490 = v_38485 | v_38489;
assign v_38492 = v_38387 | v_38491;
assign v_38494 = v_38385 | v_38493;
assign v_38496 = v_38491 | v_38495;
assign v_38498 = v_38384 | v_38497;
assign v_38500 = v_38382 | v_38499;
assign v_38502 = v_38497 | v_38501;
assign v_38504 = v_38381 | v_38503;
assign v_38506 = v_38379 | v_38505;
assign v_38508 = v_38503 | v_38507;
assign v_38510 = v_38378 | v_38509;
assign v_38512 = v_38376 | v_38511;
assign v_38514 = v_38509 | v_38513;
assign v_38516 = v_38375 | v_38515;
assign v_38518 = v_38373 | v_38517;
assign v_38520 = v_38515 | v_38519;
assign v_38523 = ~v_38372 | v_38522;
assign v_38530 = v_38420 | v_38529;
assign v_38533 = v_38531 | v_38532;
assign v_38535 = v_38417 | v_38534;
assign v_38538 = v_38536 | v_38537;
assign v_38540 = v_38414 | v_38539;
assign v_38543 = v_38541 | v_38542;
assign v_38545 = v_38411 | v_38544;
assign v_38548 = v_38546 | v_38547;
assign v_38550 = v_38408 | v_38549;
assign v_38553 = v_38551 | v_38552;
assign v_38555 = v_38405 | v_38554;
assign v_38558 = v_38556 | v_38557;
assign v_38560 = v_38402 | v_38559;
assign v_38563 = v_38561 | v_38562;
assign v_38565 = v_38399 | v_38564;
assign v_38568 = v_38566 | v_38567;
assign v_38570 = v_38396 | v_38569;
assign v_38573 = v_38571 | v_38572;
assign v_38575 = v_38393 | v_38574;
assign v_38578 = v_38576 | v_38577;
assign v_38580 = v_38390 | v_38579;
assign v_38583 = v_38581 | v_38582;
assign v_38585 = v_38387 | v_38584;
assign v_38588 = v_38586 | v_38587;
assign v_38590 = v_38384 | v_38589;
assign v_38593 = v_38591 | v_38592;
assign v_38595 = v_38381 | v_38594;
assign v_38598 = v_38596 | v_38597;
assign v_38600 = v_38378 | v_38599;
assign v_38603 = v_38601 | v_38602;
assign v_38605 = v_38375 | v_38604;
assign v_38608 = v_38606 | v_38607;
assign v_38610 = v_38372 | v_38609;
assign v_38613 = v_38371 | v_38612;
assign v_38667 = v_38664 | v_38666;
assign v_38669 = v_38663 | v_38668;
assign v_38671 = v_38661 | v_38670;
assign v_38673 = v_38668 | v_38672;
assign v_38675 = v_38660 | v_38674;
assign v_38677 = v_38658 | v_38676;
assign v_38679 = v_38674 | v_38678;
assign v_38681 = v_38657 | v_38680;
assign v_38683 = v_38655 | v_38682;
assign v_38685 = v_38680 | v_38684;
assign v_38687 = v_38654 | v_38686;
assign v_38689 = v_38652 | v_38688;
assign v_38691 = v_38686 | v_38690;
assign v_38693 = v_38651 | v_38692;
assign v_38695 = v_38649 | v_38694;
assign v_38697 = v_38692 | v_38696;
assign v_38699 = v_38648 | v_38698;
assign v_38701 = v_38646 | v_38700;
assign v_38703 = v_38698 | v_38702;
assign v_38705 = v_38645 | v_38704;
assign v_38707 = v_38643 | v_38706;
assign v_38709 = v_38704 | v_38708;
assign v_38711 = v_38642 | v_38710;
assign v_38713 = v_38640 | v_38712;
assign v_38715 = v_38710 | v_38714;
assign v_38717 = v_38639 | v_38716;
assign v_38719 = v_38637 | v_38718;
assign v_38721 = v_38716 | v_38720;
assign v_38723 = v_38636 | v_38722;
assign v_38725 = v_38634 | v_38724;
assign v_38727 = v_38722 | v_38726;
assign v_38729 = v_38633 | v_38728;
assign v_38731 = v_38631 | v_38730;
assign v_38733 = v_38728 | v_38732;
assign v_38735 = v_38630 | v_38734;
assign v_38737 = v_38628 | v_38736;
assign v_38739 = v_38734 | v_38738;
assign v_38741 = v_38627 | v_38740;
assign v_38743 = v_38625 | v_38742;
assign v_38745 = v_38740 | v_38744;
assign v_38747 = v_38624 | v_38746;
assign v_38749 = v_38622 | v_38748;
assign v_38751 = v_38746 | v_38750;
assign v_38753 = v_38621 | v_38752;
assign v_38755 = v_38619 | v_38754;
assign v_38757 = v_38752 | v_38756;
assign v_38759 = v_38618 | v_38758;
assign v_38761 = v_38616 | v_38760;
assign v_38763 = v_38758 | v_38762;
assign v_38766 = ~v_38615 | v_38765;
assign v_38773 = v_38663 | v_38772;
assign v_38776 = v_38774 | v_38775;
assign v_38778 = v_38660 | v_38777;
assign v_38781 = v_38779 | v_38780;
assign v_38783 = v_38657 | v_38782;
assign v_38786 = v_38784 | v_38785;
assign v_38788 = v_38654 | v_38787;
assign v_38791 = v_38789 | v_38790;
assign v_38793 = v_38651 | v_38792;
assign v_38796 = v_38794 | v_38795;
assign v_38798 = v_38648 | v_38797;
assign v_38801 = v_38799 | v_38800;
assign v_38803 = v_38645 | v_38802;
assign v_38806 = v_38804 | v_38805;
assign v_38808 = v_38642 | v_38807;
assign v_38811 = v_38809 | v_38810;
assign v_38813 = v_38639 | v_38812;
assign v_38816 = v_38814 | v_38815;
assign v_38818 = v_38636 | v_38817;
assign v_38821 = v_38819 | v_38820;
assign v_38823 = v_38633 | v_38822;
assign v_38826 = v_38824 | v_38825;
assign v_38828 = v_38630 | v_38827;
assign v_38831 = v_38829 | v_38830;
assign v_38833 = v_38627 | v_38832;
assign v_38836 = v_38834 | v_38835;
assign v_38838 = v_38624 | v_38837;
assign v_38841 = v_38839 | v_38840;
assign v_38843 = v_38621 | v_38842;
assign v_38846 = v_38844 | v_38845;
assign v_38848 = v_38618 | v_38847;
assign v_38851 = v_38849 | v_38850;
assign v_38853 = v_38615 | v_38852;
assign v_38856 = v_38614 | v_38855;
assign v_38910 = v_38907 | v_38909;
assign v_38912 = v_38906 | v_38911;
assign v_38914 = v_38904 | v_38913;
assign v_38916 = v_38911 | v_38915;
assign v_38918 = v_38903 | v_38917;
assign v_38920 = v_38901 | v_38919;
assign v_38922 = v_38917 | v_38921;
assign v_38924 = v_38900 | v_38923;
assign v_38926 = v_38898 | v_38925;
assign v_38928 = v_38923 | v_38927;
assign v_38930 = v_38897 | v_38929;
assign v_38932 = v_38895 | v_38931;
assign v_38934 = v_38929 | v_38933;
assign v_38936 = v_38894 | v_38935;
assign v_38938 = v_38892 | v_38937;
assign v_38940 = v_38935 | v_38939;
assign v_38942 = v_38891 | v_38941;
assign v_38944 = v_38889 | v_38943;
assign v_38946 = v_38941 | v_38945;
assign v_38948 = v_38888 | v_38947;
assign v_38950 = v_38886 | v_38949;
assign v_38952 = v_38947 | v_38951;
assign v_38954 = v_38885 | v_38953;
assign v_38956 = v_38883 | v_38955;
assign v_38958 = v_38953 | v_38957;
assign v_38960 = v_38882 | v_38959;
assign v_38962 = v_38880 | v_38961;
assign v_38964 = v_38959 | v_38963;
assign v_38966 = v_38879 | v_38965;
assign v_38968 = v_38877 | v_38967;
assign v_38970 = v_38965 | v_38969;
assign v_38972 = v_38876 | v_38971;
assign v_38974 = v_38874 | v_38973;
assign v_38976 = v_38971 | v_38975;
assign v_38978 = v_38873 | v_38977;
assign v_38980 = v_38871 | v_38979;
assign v_38982 = v_38977 | v_38981;
assign v_38984 = v_38870 | v_38983;
assign v_38986 = v_38868 | v_38985;
assign v_38988 = v_38983 | v_38987;
assign v_38990 = v_38867 | v_38989;
assign v_38992 = v_38865 | v_38991;
assign v_38994 = v_38989 | v_38993;
assign v_38996 = v_38864 | v_38995;
assign v_38998 = v_38862 | v_38997;
assign v_39000 = v_38995 | v_38999;
assign v_39002 = v_38861 | v_39001;
assign v_39004 = v_38859 | v_39003;
assign v_39006 = v_39001 | v_39005;
assign v_39009 = ~v_38858 | v_39008;
assign v_39016 = v_38906 | v_39015;
assign v_39019 = v_39017 | v_39018;
assign v_39021 = v_38903 | v_39020;
assign v_39024 = v_39022 | v_39023;
assign v_39026 = v_38900 | v_39025;
assign v_39029 = v_39027 | v_39028;
assign v_39031 = v_38897 | v_39030;
assign v_39034 = v_39032 | v_39033;
assign v_39036 = v_38894 | v_39035;
assign v_39039 = v_39037 | v_39038;
assign v_39041 = v_38891 | v_39040;
assign v_39044 = v_39042 | v_39043;
assign v_39046 = v_38888 | v_39045;
assign v_39049 = v_39047 | v_39048;
assign v_39051 = v_38885 | v_39050;
assign v_39054 = v_39052 | v_39053;
assign v_39056 = v_38882 | v_39055;
assign v_39059 = v_39057 | v_39058;
assign v_39061 = v_38879 | v_39060;
assign v_39064 = v_39062 | v_39063;
assign v_39066 = v_38876 | v_39065;
assign v_39069 = v_39067 | v_39068;
assign v_39071 = v_38873 | v_39070;
assign v_39074 = v_39072 | v_39073;
assign v_39076 = v_38870 | v_39075;
assign v_39079 = v_39077 | v_39078;
assign v_39081 = v_38867 | v_39080;
assign v_39084 = v_39082 | v_39083;
assign v_39086 = v_38864 | v_39085;
assign v_39089 = v_39087 | v_39088;
assign v_39091 = v_38861 | v_39090;
assign v_39094 = v_39092 | v_39093;
assign v_39096 = v_38858 | v_39095;
assign v_39099 = v_38857 | v_39098;
assign v_39153 = v_39150 | v_39152;
assign v_39155 = v_39149 | v_39154;
assign v_39157 = v_39147 | v_39156;
assign v_39159 = v_39154 | v_39158;
assign v_39161 = v_39146 | v_39160;
assign v_39163 = v_39144 | v_39162;
assign v_39165 = v_39160 | v_39164;
assign v_39167 = v_39143 | v_39166;
assign v_39169 = v_39141 | v_39168;
assign v_39171 = v_39166 | v_39170;
assign v_39173 = v_39140 | v_39172;
assign v_39175 = v_39138 | v_39174;
assign v_39177 = v_39172 | v_39176;
assign v_39179 = v_39137 | v_39178;
assign v_39181 = v_39135 | v_39180;
assign v_39183 = v_39178 | v_39182;
assign v_39185 = v_39134 | v_39184;
assign v_39187 = v_39132 | v_39186;
assign v_39189 = v_39184 | v_39188;
assign v_39191 = v_39131 | v_39190;
assign v_39193 = v_39129 | v_39192;
assign v_39195 = v_39190 | v_39194;
assign v_39197 = v_39128 | v_39196;
assign v_39199 = v_39126 | v_39198;
assign v_39201 = v_39196 | v_39200;
assign v_39203 = v_39125 | v_39202;
assign v_39205 = v_39123 | v_39204;
assign v_39207 = v_39202 | v_39206;
assign v_39209 = v_39122 | v_39208;
assign v_39211 = v_39120 | v_39210;
assign v_39213 = v_39208 | v_39212;
assign v_39215 = v_39119 | v_39214;
assign v_39217 = v_39117 | v_39216;
assign v_39219 = v_39214 | v_39218;
assign v_39221 = v_39116 | v_39220;
assign v_39223 = v_39114 | v_39222;
assign v_39225 = v_39220 | v_39224;
assign v_39227 = v_39113 | v_39226;
assign v_39229 = v_39111 | v_39228;
assign v_39231 = v_39226 | v_39230;
assign v_39233 = v_39110 | v_39232;
assign v_39235 = v_39108 | v_39234;
assign v_39237 = v_39232 | v_39236;
assign v_39239 = v_39107 | v_39238;
assign v_39241 = v_39105 | v_39240;
assign v_39243 = v_39238 | v_39242;
assign v_39245 = v_39104 | v_39244;
assign v_39247 = v_39102 | v_39246;
assign v_39249 = v_39244 | v_39248;
assign v_39252 = ~v_39101 | v_39251;
assign v_39259 = v_39149 | v_39258;
assign v_39262 = v_39260 | v_39261;
assign v_39264 = v_39146 | v_39263;
assign v_39267 = v_39265 | v_39266;
assign v_39269 = v_39143 | v_39268;
assign v_39272 = v_39270 | v_39271;
assign v_39274 = v_39140 | v_39273;
assign v_39277 = v_39275 | v_39276;
assign v_39279 = v_39137 | v_39278;
assign v_39282 = v_39280 | v_39281;
assign v_39284 = v_39134 | v_39283;
assign v_39287 = v_39285 | v_39286;
assign v_39289 = v_39131 | v_39288;
assign v_39292 = v_39290 | v_39291;
assign v_39294 = v_39128 | v_39293;
assign v_39297 = v_39295 | v_39296;
assign v_39299 = v_39125 | v_39298;
assign v_39302 = v_39300 | v_39301;
assign v_39304 = v_39122 | v_39303;
assign v_39307 = v_39305 | v_39306;
assign v_39309 = v_39119 | v_39308;
assign v_39312 = v_39310 | v_39311;
assign v_39314 = v_39116 | v_39313;
assign v_39317 = v_39315 | v_39316;
assign v_39319 = v_39113 | v_39318;
assign v_39322 = v_39320 | v_39321;
assign v_39324 = v_39110 | v_39323;
assign v_39327 = v_39325 | v_39326;
assign v_39329 = v_39107 | v_39328;
assign v_39332 = v_39330 | v_39331;
assign v_39334 = v_39104 | v_39333;
assign v_39337 = v_39335 | v_39336;
assign v_39339 = v_39101 | v_39338;
assign v_39342 = v_39100 | v_39341;
assign v_39396 = v_39393 | v_39395;
assign v_39398 = v_39392 | v_39397;
assign v_39400 = v_39390 | v_39399;
assign v_39402 = v_39397 | v_39401;
assign v_39404 = v_39389 | v_39403;
assign v_39406 = v_39387 | v_39405;
assign v_39408 = v_39403 | v_39407;
assign v_39410 = v_39386 | v_39409;
assign v_39412 = v_39384 | v_39411;
assign v_39414 = v_39409 | v_39413;
assign v_39416 = v_39383 | v_39415;
assign v_39418 = v_39381 | v_39417;
assign v_39420 = v_39415 | v_39419;
assign v_39422 = v_39380 | v_39421;
assign v_39424 = v_39378 | v_39423;
assign v_39426 = v_39421 | v_39425;
assign v_39428 = v_39377 | v_39427;
assign v_39430 = v_39375 | v_39429;
assign v_39432 = v_39427 | v_39431;
assign v_39434 = v_39374 | v_39433;
assign v_39436 = v_39372 | v_39435;
assign v_39438 = v_39433 | v_39437;
assign v_39440 = v_39371 | v_39439;
assign v_39442 = v_39369 | v_39441;
assign v_39444 = v_39439 | v_39443;
assign v_39446 = v_39368 | v_39445;
assign v_39448 = v_39366 | v_39447;
assign v_39450 = v_39445 | v_39449;
assign v_39452 = v_39365 | v_39451;
assign v_39454 = v_39363 | v_39453;
assign v_39456 = v_39451 | v_39455;
assign v_39458 = v_39362 | v_39457;
assign v_39460 = v_39360 | v_39459;
assign v_39462 = v_39457 | v_39461;
assign v_39464 = v_39359 | v_39463;
assign v_39466 = v_39357 | v_39465;
assign v_39468 = v_39463 | v_39467;
assign v_39470 = v_39356 | v_39469;
assign v_39472 = v_39354 | v_39471;
assign v_39474 = v_39469 | v_39473;
assign v_39476 = v_39353 | v_39475;
assign v_39478 = v_39351 | v_39477;
assign v_39480 = v_39475 | v_39479;
assign v_39482 = v_39350 | v_39481;
assign v_39484 = v_39348 | v_39483;
assign v_39486 = v_39481 | v_39485;
assign v_39488 = v_39347 | v_39487;
assign v_39490 = v_39345 | v_39489;
assign v_39492 = v_39487 | v_39491;
assign v_39495 = ~v_39344 | v_39494;
assign v_39502 = v_39392 | v_39501;
assign v_39505 = v_39503 | v_39504;
assign v_39507 = v_39389 | v_39506;
assign v_39510 = v_39508 | v_39509;
assign v_39512 = v_39386 | v_39511;
assign v_39515 = v_39513 | v_39514;
assign v_39517 = v_39383 | v_39516;
assign v_39520 = v_39518 | v_39519;
assign v_39522 = v_39380 | v_39521;
assign v_39525 = v_39523 | v_39524;
assign v_39527 = v_39377 | v_39526;
assign v_39530 = v_39528 | v_39529;
assign v_39532 = v_39374 | v_39531;
assign v_39535 = v_39533 | v_39534;
assign v_39537 = v_39371 | v_39536;
assign v_39540 = v_39538 | v_39539;
assign v_39542 = v_39368 | v_39541;
assign v_39545 = v_39543 | v_39544;
assign v_39547 = v_39365 | v_39546;
assign v_39550 = v_39548 | v_39549;
assign v_39552 = v_39362 | v_39551;
assign v_39555 = v_39553 | v_39554;
assign v_39557 = v_39359 | v_39556;
assign v_39560 = v_39558 | v_39559;
assign v_39562 = v_39356 | v_39561;
assign v_39565 = v_39563 | v_39564;
assign v_39567 = v_39353 | v_39566;
assign v_39570 = v_39568 | v_39569;
assign v_39572 = v_39350 | v_39571;
assign v_39575 = v_39573 | v_39574;
assign v_39577 = v_39347 | v_39576;
assign v_39580 = v_39578 | v_39579;
assign v_39582 = v_39344 | v_39581;
assign v_39585 = v_39343 | v_39584;
assign v_39639 = v_39636 | v_39638;
assign v_39641 = v_39635 | v_39640;
assign v_39643 = v_39633 | v_39642;
assign v_39645 = v_39640 | v_39644;
assign v_39647 = v_39632 | v_39646;
assign v_39649 = v_39630 | v_39648;
assign v_39651 = v_39646 | v_39650;
assign v_39653 = v_39629 | v_39652;
assign v_39655 = v_39627 | v_39654;
assign v_39657 = v_39652 | v_39656;
assign v_39659 = v_39626 | v_39658;
assign v_39661 = v_39624 | v_39660;
assign v_39663 = v_39658 | v_39662;
assign v_39665 = v_39623 | v_39664;
assign v_39667 = v_39621 | v_39666;
assign v_39669 = v_39664 | v_39668;
assign v_39671 = v_39620 | v_39670;
assign v_39673 = v_39618 | v_39672;
assign v_39675 = v_39670 | v_39674;
assign v_39677 = v_39617 | v_39676;
assign v_39679 = v_39615 | v_39678;
assign v_39681 = v_39676 | v_39680;
assign v_39683 = v_39614 | v_39682;
assign v_39685 = v_39612 | v_39684;
assign v_39687 = v_39682 | v_39686;
assign v_39689 = v_39611 | v_39688;
assign v_39691 = v_39609 | v_39690;
assign v_39693 = v_39688 | v_39692;
assign v_39695 = v_39608 | v_39694;
assign v_39697 = v_39606 | v_39696;
assign v_39699 = v_39694 | v_39698;
assign v_39701 = v_39605 | v_39700;
assign v_39703 = v_39603 | v_39702;
assign v_39705 = v_39700 | v_39704;
assign v_39707 = v_39602 | v_39706;
assign v_39709 = v_39600 | v_39708;
assign v_39711 = v_39706 | v_39710;
assign v_39713 = v_39599 | v_39712;
assign v_39715 = v_39597 | v_39714;
assign v_39717 = v_39712 | v_39716;
assign v_39719 = v_39596 | v_39718;
assign v_39721 = v_39594 | v_39720;
assign v_39723 = v_39718 | v_39722;
assign v_39725 = v_39593 | v_39724;
assign v_39727 = v_39591 | v_39726;
assign v_39729 = v_39724 | v_39728;
assign v_39731 = v_39590 | v_39730;
assign v_39733 = v_39588 | v_39732;
assign v_39735 = v_39730 | v_39734;
assign v_39738 = ~v_39587 | v_39737;
assign v_39745 = v_39635 | v_39744;
assign v_39748 = v_39746 | v_39747;
assign v_39750 = v_39632 | v_39749;
assign v_39753 = v_39751 | v_39752;
assign v_39755 = v_39629 | v_39754;
assign v_39758 = v_39756 | v_39757;
assign v_39760 = v_39626 | v_39759;
assign v_39763 = v_39761 | v_39762;
assign v_39765 = v_39623 | v_39764;
assign v_39768 = v_39766 | v_39767;
assign v_39770 = v_39620 | v_39769;
assign v_39773 = v_39771 | v_39772;
assign v_39775 = v_39617 | v_39774;
assign v_39778 = v_39776 | v_39777;
assign v_39780 = v_39614 | v_39779;
assign v_39783 = v_39781 | v_39782;
assign v_39785 = v_39611 | v_39784;
assign v_39788 = v_39786 | v_39787;
assign v_39790 = v_39608 | v_39789;
assign v_39793 = v_39791 | v_39792;
assign v_39795 = v_39605 | v_39794;
assign v_39798 = v_39796 | v_39797;
assign v_39800 = v_39602 | v_39799;
assign v_39803 = v_39801 | v_39802;
assign v_39805 = v_39599 | v_39804;
assign v_39808 = v_39806 | v_39807;
assign v_39810 = v_39596 | v_39809;
assign v_39813 = v_39811 | v_39812;
assign v_39815 = v_39593 | v_39814;
assign v_39818 = v_39816 | v_39817;
assign v_39820 = v_39590 | v_39819;
assign v_39823 = v_39821 | v_39822;
assign v_39825 = v_39587 | v_39824;
assign v_39828 = v_39586 | v_39827;
assign v_39882 = v_39879 | v_39881;
assign v_39884 = v_39878 | v_39883;
assign v_39886 = v_39876 | v_39885;
assign v_39888 = v_39883 | v_39887;
assign v_39890 = v_39875 | v_39889;
assign v_39892 = v_39873 | v_39891;
assign v_39894 = v_39889 | v_39893;
assign v_39896 = v_39872 | v_39895;
assign v_39898 = v_39870 | v_39897;
assign v_39900 = v_39895 | v_39899;
assign v_39902 = v_39869 | v_39901;
assign v_39904 = v_39867 | v_39903;
assign v_39906 = v_39901 | v_39905;
assign v_39908 = v_39866 | v_39907;
assign v_39910 = v_39864 | v_39909;
assign v_39912 = v_39907 | v_39911;
assign v_39914 = v_39863 | v_39913;
assign v_39916 = v_39861 | v_39915;
assign v_39918 = v_39913 | v_39917;
assign v_39920 = v_39860 | v_39919;
assign v_39922 = v_39858 | v_39921;
assign v_39924 = v_39919 | v_39923;
assign v_39926 = v_39857 | v_39925;
assign v_39928 = v_39855 | v_39927;
assign v_39930 = v_39925 | v_39929;
assign v_39932 = v_39854 | v_39931;
assign v_39934 = v_39852 | v_39933;
assign v_39936 = v_39931 | v_39935;
assign v_39938 = v_39851 | v_39937;
assign v_39940 = v_39849 | v_39939;
assign v_39942 = v_39937 | v_39941;
assign v_39944 = v_39848 | v_39943;
assign v_39946 = v_39846 | v_39945;
assign v_39948 = v_39943 | v_39947;
assign v_39950 = v_39845 | v_39949;
assign v_39952 = v_39843 | v_39951;
assign v_39954 = v_39949 | v_39953;
assign v_39956 = v_39842 | v_39955;
assign v_39958 = v_39840 | v_39957;
assign v_39960 = v_39955 | v_39959;
assign v_39962 = v_39839 | v_39961;
assign v_39964 = v_39837 | v_39963;
assign v_39966 = v_39961 | v_39965;
assign v_39968 = v_39836 | v_39967;
assign v_39970 = v_39834 | v_39969;
assign v_39972 = v_39967 | v_39971;
assign v_39974 = v_39833 | v_39973;
assign v_39976 = v_39831 | v_39975;
assign v_39978 = v_39973 | v_39977;
assign v_39981 = ~v_39830 | v_39980;
assign v_39988 = v_39878 | v_39987;
assign v_39991 = v_39989 | v_39990;
assign v_39993 = v_39875 | v_39992;
assign v_39996 = v_39994 | v_39995;
assign v_39998 = v_39872 | v_39997;
assign v_40001 = v_39999 | v_40000;
assign v_40003 = v_39869 | v_40002;
assign v_40006 = v_40004 | v_40005;
assign v_40008 = v_39866 | v_40007;
assign v_40011 = v_40009 | v_40010;
assign v_40013 = v_39863 | v_40012;
assign v_40016 = v_40014 | v_40015;
assign v_40018 = v_39860 | v_40017;
assign v_40021 = v_40019 | v_40020;
assign v_40023 = v_39857 | v_40022;
assign v_40026 = v_40024 | v_40025;
assign v_40028 = v_39854 | v_40027;
assign v_40031 = v_40029 | v_40030;
assign v_40033 = v_39851 | v_40032;
assign v_40036 = v_40034 | v_40035;
assign v_40038 = v_39848 | v_40037;
assign v_40041 = v_40039 | v_40040;
assign v_40043 = v_39845 | v_40042;
assign v_40046 = v_40044 | v_40045;
assign v_40048 = v_39842 | v_40047;
assign v_40051 = v_40049 | v_40050;
assign v_40053 = v_39839 | v_40052;
assign v_40056 = v_40054 | v_40055;
assign v_40058 = v_39836 | v_40057;
assign v_40061 = v_40059 | v_40060;
assign v_40063 = v_39833 | v_40062;
assign v_40066 = v_40064 | v_40065;
assign v_40068 = v_39830 | v_40067;
assign v_40071 = v_39829 | v_40070;
assign v_40125 = v_40122 | v_40124;
assign v_40127 = v_40121 | v_40126;
assign v_40129 = v_40119 | v_40128;
assign v_40131 = v_40126 | v_40130;
assign v_40133 = v_40118 | v_40132;
assign v_40135 = v_40116 | v_40134;
assign v_40137 = v_40132 | v_40136;
assign v_40139 = v_40115 | v_40138;
assign v_40141 = v_40113 | v_40140;
assign v_40143 = v_40138 | v_40142;
assign v_40145 = v_40112 | v_40144;
assign v_40147 = v_40110 | v_40146;
assign v_40149 = v_40144 | v_40148;
assign v_40151 = v_40109 | v_40150;
assign v_40153 = v_40107 | v_40152;
assign v_40155 = v_40150 | v_40154;
assign v_40157 = v_40106 | v_40156;
assign v_40159 = v_40104 | v_40158;
assign v_40161 = v_40156 | v_40160;
assign v_40163 = v_40103 | v_40162;
assign v_40165 = v_40101 | v_40164;
assign v_40167 = v_40162 | v_40166;
assign v_40169 = v_40100 | v_40168;
assign v_40171 = v_40098 | v_40170;
assign v_40173 = v_40168 | v_40172;
assign v_40175 = v_40097 | v_40174;
assign v_40177 = v_40095 | v_40176;
assign v_40179 = v_40174 | v_40178;
assign v_40181 = v_40094 | v_40180;
assign v_40183 = v_40092 | v_40182;
assign v_40185 = v_40180 | v_40184;
assign v_40187 = v_40091 | v_40186;
assign v_40189 = v_40089 | v_40188;
assign v_40191 = v_40186 | v_40190;
assign v_40193 = v_40088 | v_40192;
assign v_40195 = v_40086 | v_40194;
assign v_40197 = v_40192 | v_40196;
assign v_40199 = v_40085 | v_40198;
assign v_40201 = v_40083 | v_40200;
assign v_40203 = v_40198 | v_40202;
assign v_40205 = v_40082 | v_40204;
assign v_40207 = v_40080 | v_40206;
assign v_40209 = v_40204 | v_40208;
assign v_40211 = v_40079 | v_40210;
assign v_40213 = v_40077 | v_40212;
assign v_40215 = v_40210 | v_40214;
assign v_40217 = v_40076 | v_40216;
assign v_40219 = v_40074 | v_40218;
assign v_40221 = v_40216 | v_40220;
assign v_40224 = ~v_40073 | v_40223;
assign v_40231 = v_40121 | v_40230;
assign v_40234 = v_40232 | v_40233;
assign v_40236 = v_40118 | v_40235;
assign v_40239 = v_40237 | v_40238;
assign v_40241 = v_40115 | v_40240;
assign v_40244 = v_40242 | v_40243;
assign v_40246 = v_40112 | v_40245;
assign v_40249 = v_40247 | v_40248;
assign v_40251 = v_40109 | v_40250;
assign v_40254 = v_40252 | v_40253;
assign v_40256 = v_40106 | v_40255;
assign v_40259 = v_40257 | v_40258;
assign v_40261 = v_40103 | v_40260;
assign v_40264 = v_40262 | v_40263;
assign v_40266 = v_40100 | v_40265;
assign v_40269 = v_40267 | v_40268;
assign v_40271 = v_40097 | v_40270;
assign v_40274 = v_40272 | v_40273;
assign v_40276 = v_40094 | v_40275;
assign v_40279 = v_40277 | v_40278;
assign v_40281 = v_40091 | v_40280;
assign v_40284 = v_40282 | v_40283;
assign v_40286 = v_40088 | v_40285;
assign v_40289 = v_40287 | v_40288;
assign v_40291 = v_40085 | v_40290;
assign v_40294 = v_40292 | v_40293;
assign v_40296 = v_40082 | v_40295;
assign v_40299 = v_40297 | v_40298;
assign v_40301 = v_40079 | v_40300;
assign v_40304 = v_40302 | v_40303;
assign v_40306 = v_40076 | v_40305;
assign v_40309 = v_40307 | v_40308;
assign v_40311 = v_40073 | v_40310;
assign v_40314 = v_40072 | v_40313;
assign v_40368 = v_40365 | v_40367;
assign v_40370 = v_40364 | v_40369;
assign v_40372 = v_40362 | v_40371;
assign v_40374 = v_40369 | v_40373;
assign v_40376 = v_40361 | v_40375;
assign v_40378 = v_40359 | v_40377;
assign v_40380 = v_40375 | v_40379;
assign v_40382 = v_40358 | v_40381;
assign v_40384 = v_40356 | v_40383;
assign v_40386 = v_40381 | v_40385;
assign v_40388 = v_40355 | v_40387;
assign v_40390 = v_40353 | v_40389;
assign v_40392 = v_40387 | v_40391;
assign v_40394 = v_40352 | v_40393;
assign v_40396 = v_40350 | v_40395;
assign v_40398 = v_40393 | v_40397;
assign v_40400 = v_40349 | v_40399;
assign v_40402 = v_40347 | v_40401;
assign v_40404 = v_40399 | v_40403;
assign v_40406 = v_40346 | v_40405;
assign v_40408 = v_40344 | v_40407;
assign v_40410 = v_40405 | v_40409;
assign v_40412 = v_40343 | v_40411;
assign v_40414 = v_40341 | v_40413;
assign v_40416 = v_40411 | v_40415;
assign v_40418 = v_40340 | v_40417;
assign v_40420 = v_40338 | v_40419;
assign v_40422 = v_40417 | v_40421;
assign v_40424 = v_40337 | v_40423;
assign v_40426 = v_40335 | v_40425;
assign v_40428 = v_40423 | v_40427;
assign v_40430 = v_40334 | v_40429;
assign v_40432 = v_40332 | v_40431;
assign v_40434 = v_40429 | v_40433;
assign v_40436 = v_40331 | v_40435;
assign v_40438 = v_40329 | v_40437;
assign v_40440 = v_40435 | v_40439;
assign v_40442 = v_40328 | v_40441;
assign v_40444 = v_40326 | v_40443;
assign v_40446 = v_40441 | v_40445;
assign v_40448 = v_40325 | v_40447;
assign v_40450 = v_40323 | v_40449;
assign v_40452 = v_40447 | v_40451;
assign v_40454 = v_40322 | v_40453;
assign v_40456 = v_40320 | v_40455;
assign v_40458 = v_40453 | v_40457;
assign v_40460 = v_40319 | v_40459;
assign v_40462 = v_40317 | v_40461;
assign v_40464 = v_40459 | v_40463;
assign v_40467 = ~v_40316 | v_40466;
assign v_40474 = v_40364 | v_40473;
assign v_40477 = v_40475 | v_40476;
assign v_40479 = v_40361 | v_40478;
assign v_40482 = v_40480 | v_40481;
assign v_40484 = v_40358 | v_40483;
assign v_40487 = v_40485 | v_40486;
assign v_40489 = v_40355 | v_40488;
assign v_40492 = v_40490 | v_40491;
assign v_40494 = v_40352 | v_40493;
assign v_40497 = v_40495 | v_40496;
assign v_40499 = v_40349 | v_40498;
assign v_40502 = v_40500 | v_40501;
assign v_40504 = v_40346 | v_40503;
assign v_40507 = v_40505 | v_40506;
assign v_40509 = v_40343 | v_40508;
assign v_40512 = v_40510 | v_40511;
assign v_40514 = v_40340 | v_40513;
assign v_40517 = v_40515 | v_40516;
assign v_40519 = v_40337 | v_40518;
assign v_40522 = v_40520 | v_40521;
assign v_40524 = v_40334 | v_40523;
assign v_40527 = v_40525 | v_40526;
assign v_40529 = v_40331 | v_40528;
assign v_40532 = v_40530 | v_40531;
assign v_40534 = v_40328 | v_40533;
assign v_40537 = v_40535 | v_40536;
assign v_40539 = v_40325 | v_40538;
assign v_40542 = v_40540 | v_40541;
assign v_40544 = v_40322 | v_40543;
assign v_40547 = v_40545 | v_40546;
assign v_40549 = v_40319 | v_40548;
assign v_40552 = v_40550 | v_40551;
assign v_40554 = v_40316 | v_40553;
assign v_40557 = v_40315 | v_40556;
assign v_40611 = v_40608 | v_40610;
assign v_40613 = v_40607 | v_40612;
assign v_40615 = v_40605 | v_40614;
assign v_40617 = v_40612 | v_40616;
assign v_40619 = v_40604 | v_40618;
assign v_40621 = v_40602 | v_40620;
assign v_40623 = v_40618 | v_40622;
assign v_40625 = v_40601 | v_40624;
assign v_40627 = v_40599 | v_40626;
assign v_40629 = v_40624 | v_40628;
assign v_40631 = v_40598 | v_40630;
assign v_40633 = v_40596 | v_40632;
assign v_40635 = v_40630 | v_40634;
assign v_40637 = v_40595 | v_40636;
assign v_40639 = v_40593 | v_40638;
assign v_40641 = v_40636 | v_40640;
assign v_40643 = v_40592 | v_40642;
assign v_40645 = v_40590 | v_40644;
assign v_40647 = v_40642 | v_40646;
assign v_40649 = v_40589 | v_40648;
assign v_40651 = v_40587 | v_40650;
assign v_40653 = v_40648 | v_40652;
assign v_40655 = v_40586 | v_40654;
assign v_40657 = v_40584 | v_40656;
assign v_40659 = v_40654 | v_40658;
assign v_40661 = v_40583 | v_40660;
assign v_40663 = v_40581 | v_40662;
assign v_40665 = v_40660 | v_40664;
assign v_40667 = v_40580 | v_40666;
assign v_40669 = v_40578 | v_40668;
assign v_40671 = v_40666 | v_40670;
assign v_40673 = v_40577 | v_40672;
assign v_40675 = v_40575 | v_40674;
assign v_40677 = v_40672 | v_40676;
assign v_40679 = v_40574 | v_40678;
assign v_40681 = v_40572 | v_40680;
assign v_40683 = v_40678 | v_40682;
assign v_40685 = v_40571 | v_40684;
assign v_40687 = v_40569 | v_40686;
assign v_40689 = v_40684 | v_40688;
assign v_40691 = v_40568 | v_40690;
assign v_40693 = v_40566 | v_40692;
assign v_40695 = v_40690 | v_40694;
assign v_40697 = v_40565 | v_40696;
assign v_40699 = v_40563 | v_40698;
assign v_40701 = v_40696 | v_40700;
assign v_40703 = v_40562 | v_40702;
assign v_40705 = v_40560 | v_40704;
assign v_40707 = v_40702 | v_40706;
assign v_40710 = ~v_40559 | v_40709;
assign v_40717 = v_40607 | v_40716;
assign v_40720 = v_40718 | v_40719;
assign v_40722 = v_40604 | v_40721;
assign v_40725 = v_40723 | v_40724;
assign v_40727 = v_40601 | v_40726;
assign v_40730 = v_40728 | v_40729;
assign v_40732 = v_40598 | v_40731;
assign v_40735 = v_40733 | v_40734;
assign v_40737 = v_40595 | v_40736;
assign v_40740 = v_40738 | v_40739;
assign v_40742 = v_40592 | v_40741;
assign v_40745 = v_40743 | v_40744;
assign v_40747 = v_40589 | v_40746;
assign v_40750 = v_40748 | v_40749;
assign v_40752 = v_40586 | v_40751;
assign v_40755 = v_40753 | v_40754;
assign v_40757 = v_40583 | v_40756;
assign v_40760 = v_40758 | v_40759;
assign v_40762 = v_40580 | v_40761;
assign v_40765 = v_40763 | v_40764;
assign v_40767 = v_40577 | v_40766;
assign v_40770 = v_40768 | v_40769;
assign v_40772 = v_40574 | v_40771;
assign v_40775 = v_40773 | v_40774;
assign v_40777 = v_40571 | v_40776;
assign v_40780 = v_40778 | v_40779;
assign v_40782 = v_40568 | v_40781;
assign v_40785 = v_40783 | v_40784;
assign v_40787 = v_40565 | v_40786;
assign v_40790 = v_40788 | v_40789;
assign v_40792 = v_40562 | v_40791;
assign v_40795 = v_40793 | v_40794;
assign v_40797 = v_40559 | v_40796;
assign v_40800 = v_40558 | v_40799;
assign v_40854 = v_40851 | v_40853;
assign v_40856 = v_40850 | v_40855;
assign v_40858 = v_40848 | v_40857;
assign v_40860 = v_40855 | v_40859;
assign v_40862 = v_40847 | v_40861;
assign v_40864 = v_40845 | v_40863;
assign v_40866 = v_40861 | v_40865;
assign v_40868 = v_40844 | v_40867;
assign v_40870 = v_40842 | v_40869;
assign v_40872 = v_40867 | v_40871;
assign v_40874 = v_40841 | v_40873;
assign v_40876 = v_40839 | v_40875;
assign v_40878 = v_40873 | v_40877;
assign v_40880 = v_40838 | v_40879;
assign v_40882 = v_40836 | v_40881;
assign v_40884 = v_40879 | v_40883;
assign v_40886 = v_40835 | v_40885;
assign v_40888 = v_40833 | v_40887;
assign v_40890 = v_40885 | v_40889;
assign v_40892 = v_40832 | v_40891;
assign v_40894 = v_40830 | v_40893;
assign v_40896 = v_40891 | v_40895;
assign v_40898 = v_40829 | v_40897;
assign v_40900 = v_40827 | v_40899;
assign v_40902 = v_40897 | v_40901;
assign v_40904 = v_40826 | v_40903;
assign v_40906 = v_40824 | v_40905;
assign v_40908 = v_40903 | v_40907;
assign v_40910 = v_40823 | v_40909;
assign v_40912 = v_40821 | v_40911;
assign v_40914 = v_40909 | v_40913;
assign v_40916 = v_40820 | v_40915;
assign v_40918 = v_40818 | v_40917;
assign v_40920 = v_40915 | v_40919;
assign v_40922 = v_40817 | v_40921;
assign v_40924 = v_40815 | v_40923;
assign v_40926 = v_40921 | v_40925;
assign v_40928 = v_40814 | v_40927;
assign v_40930 = v_40812 | v_40929;
assign v_40932 = v_40927 | v_40931;
assign v_40934 = v_40811 | v_40933;
assign v_40936 = v_40809 | v_40935;
assign v_40938 = v_40933 | v_40937;
assign v_40940 = v_40808 | v_40939;
assign v_40942 = v_40806 | v_40941;
assign v_40944 = v_40939 | v_40943;
assign v_40946 = v_40805 | v_40945;
assign v_40948 = v_40803 | v_40947;
assign v_40950 = v_40945 | v_40949;
assign v_40953 = ~v_40802 | v_40952;
assign v_40960 = v_40850 | v_40959;
assign v_40963 = v_40961 | v_40962;
assign v_40965 = v_40847 | v_40964;
assign v_40968 = v_40966 | v_40967;
assign v_40970 = v_40844 | v_40969;
assign v_40973 = v_40971 | v_40972;
assign v_40975 = v_40841 | v_40974;
assign v_40978 = v_40976 | v_40977;
assign v_40980 = v_40838 | v_40979;
assign v_40983 = v_40981 | v_40982;
assign v_40985 = v_40835 | v_40984;
assign v_40988 = v_40986 | v_40987;
assign v_40990 = v_40832 | v_40989;
assign v_40993 = v_40991 | v_40992;
assign v_40995 = v_40829 | v_40994;
assign v_40998 = v_40996 | v_40997;
assign v_41000 = v_40826 | v_40999;
assign v_41003 = v_41001 | v_41002;
assign v_41005 = v_40823 | v_41004;
assign v_41008 = v_41006 | v_41007;
assign v_41010 = v_40820 | v_41009;
assign v_41013 = v_41011 | v_41012;
assign v_41015 = v_40817 | v_41014;
assign v_41018 = v_41016 | v_41017;
assign v_41020 = v_40814 | v_41019;
assign v_41023 = v_41021 | v_41022;
assign v_41025 = v_40811 | v_41024;
assign v_41028 = v_41026 | v_41027;
assign v_41030 = v_40808 | v_41029;
assign v_41033 = v_41031 | v_41032;
assign v_41035 = v_40805 | v_41034;
assign v_41038 = v_41036 | v_41037;
assign v_41040 = v_40802 | v_41039;
assign v_41043 = v_40801 | v_41042;
assign v_41097 = v_41094 | v_41096;
assign v_41099 = v_41093 | v_41098;
assign v_41101 = v_41091 | v_41100;
assign v_41103 = v_41098 | v_41102;
assign v_41105 = v_41090 | v_41104;
assign v_41107 = v_41088 | v_41106;
assign v_41109 = v_41104 | v_41108;
assign v_41111 = v_41087 | v_41110;
assign v_41113 = v_41085 | v_41112;
assign v_41115 = v_41110 | v_41114;
assign v_41117 = v_41084 | v_41116;
assign v_41119 = v_41082 | v_41118;
assign v_41121 = v_41116 | v_41120;
assign v_41123 = v_41081 | v_41122;
assign v_41125 = v_41079 | v_41124;
assign v_41127 = v_41122 | v_41126;
assign v_41129 = v_41078 | v_41128;
assign v_41131 = v_41076 | v_41130;
assign v_41133 = v_41128 | v_41132;
assign v_41135 = v_41075 | v_41134;
assign v_41137 = v_41073 | v_41136;
assign v_41139 = v_41134 | v_41138;
assign v_41141 = v_41072 | v_41140;
assign v_41143 = v_41070 | v_41142;
assign v_41145 = v_41140 | v_41144;
assign v_41147 = v_41069 | v_41146;
assign v_41149 = v_41067 | v_41148;
assign v_41151 = v_41146 | v_41150;
assign v_41153 = v_41066 | v_41152;
assign v_41155 = v_41064 | v_41154;
assign v_41157 = v_41152 | v_41156;
assign v_41159 = v_41063 | v_41158;
assign v_41161 = v_41061 | v_41160;
assign v_41163 = v_41158 | v_41162;
assign v_41165 = v_41060 | v_41164;
assign v_41167 = v_41058 | v_41166;
assign v_41169 = v_41164 | v_41168;
assign v_41171 = v_41057 | v_41170;
assign v_41173 = v_41055 | v_41172;
assign v_41175 = v_41170 | v_41174;
assign v_41177 = v_41054 | v_41176;
assign v_41179 = v_41052 | v_41178;
assign v_41181 = v_41176 | v_41180;
assign v_41183 = v_41051 | v_41182;
assign v_41185 = v_41049 | v_41184;
assign v_41187 = v_41182 | v_41186;
assign v_41189 = v_41048 | v_41188;
assign v_41191 = v_41046 | v_41190;
assign v_41193 = v_41188 | v_41192;
assign v_41196 = ~v_41045 | v_41195;
assign v_41203 = v_41093 | v_41202;
assign v_41206 = v_41204 | v_41205;
assign v_41208 = v_41090 | v_41207;
assign v_41211 = v_41209 | v_41210;
assign v_41213 = v_41087 | v_41212;
assign v_41216 = v_41214 | v_41215;
assign v_41218 = v_41084 | v_41217;
assign v_41221 = v_41219 | v_41220;
assign v_41223 = v_41081 | v_41222;
assign v_41226 = v_41224 | v_41225;
assign v_41228 = v_41078 | v_41227;
assign v_41231 = v_41229 | v_41230;
assign v_41233 = v_41075 | v_41232;
assign v_41236 = v_41234 | v_41235;
assign v_41238 = v_41072 | v_41237;
assign v_41241 = v_41239 | v_41240;
assign v_41243 = v_41069 | v_41242;
assign v_41246 = v_41244 | v_41245;
assign v_41248 = v_41066 | v_41247;
assign v_41251 = v_41249 | v_41250;
assign v_41253 = v_41063 | v_41252;
assign v_41256 = v_41254 | v_41255;
assign v_41258 = v_41060 | v_41257;
assign v_41261 = v_41259 | v_41260;
assign v_41263 = v_41057 | v_41262;
assign v_41266 = v_41264 | v_41265;
assign v_41268 = v_41054 | v_41267;
assign v_41271 = v_41269 | v_41270;
assign v_41273 = v_41051 | v_41272;
assign v_41276 = v_41274 | v_41275;
assign v_41278 = v_41048 | v_41277;
assign v_41281 = v_41279 | v_41280;
assign v_41283 = v_41045 | v_41282;
assign v_41286 = v_41044 | v_41285;
assign v_41340 = v_41337 | v_41339;
assign v_41342 = v_41336 | v_41341;
assign v_41344 = v_41334 | v_41343;
assign v_41346 = v_41341 | v_41345;
assign v_41348 = v_41333 | v_41347;
assign v_41350 = v_41331 | v_41349;
assign v_41352 = v_41347 | v_41351;
assign v_41354 = v_41330 | v_41353;
assign v_41356 = v_41328 | v_41355;
assign v_41358 = v_41353 | v_41357;
assign v_41360 = v_41327 | v_41359;
assign v_41362 = v_41325 | v_41361;
assign v_41364 = v_41359 | v_41363;
assign v_41366 = v_41324 | v_41365;
assign v_41368 = v_41322 | v_41367;
assign v_41370 = v_41365 | v_41369;
assign v_41372 = v_41321 | v_41371;
assign v_41374 = v_41319 | v_41373;
assign v_41376 = v_41371 | v_41375;
assign v_41378 = v_41318 | v_41377;
assign v_41380 = v_41316 | v_41379;
assign v_41382 = v_41377 | v_41381;
assign v_41384 = v_41315 | v_41383;
assign v_41386 = v_41313 | v_41385;
assign v_41388 = v_41383 | v_41387;
assign v_41390 = v_41312 | v_41389;
assign v_41392 = v_41310 | v_41391;
assign v_41394 = v_41389 | v_41393;
assign v_41396 = v_41309 | v_41395;
assign v_41398 = v_41307 | v_41397;
assign v_41400 = v_41395 | v_41399;
assign v_41402 = v_41306 | v_41401;
assign v_41404 = v_41304 | v_41403;
assign v_41406 = v_41401 | v_41405;
assign v_41408 = v_41303 | v_41407;
assign v_41410 = v_41301 | v_41409;
assign v_41412 = v_41407 | v_41411;
assign v_41414 = v_41300 | v_41413;
assign v_41416 = v_41298 | v_41415;
assign v_41418 = v_41413 | v_41417;
assign v_41420 = v_41297 | v_41419;
assign v_41422 = v_41295 | v_41421;
assign v_41424 = v_41419 | v_41423;
assign v_41426 = v_41294 | v_41425;
assign v_41428 = v_41292 | v_41427;
assign v_41430 = v_41425 | v_41429;
assign v_41432 = v_41291 | v_41431;
assign v_41434 = v_41289 | v_41433;
assign v_41436 = v_41431 | v_41435;
assign v_41439 = ~v_41288 | v_41438;
assign v_41446 = v_41336 | v_41445;
assign v_41449 = v_41447 | v_41448;
assign v_41451 = v_41333 | v_41450;
assign v_41454 = v_41452 | v_41453;
assign v_41456 = v_41330 | v_41455;
assign v_41459 = v_41457 | v_41458;
assign v_41461 = v_41327 | v_41460;
assign v_41464 = v_41462 | v_41463;
assign v_41466 = v_41324 | v_41465;
assign v_41469 = v_41467 | v_41468;
assign v_41471 = v_41321 | v_41470;
assign v_41474 = v_41472 | v_41473;
assign v_41476 = v_41318 | v_41475;
assign v_41479 = v_41477 | v_41478;
assign v_41481 = v_41315 | v_41480;
assign v_41484 = v_41482 | v_41483;
assign v_41486 = v_41312 | v_41485;
assign v_41489 = v_41487 | v_41488;
assign v_41491 = v_41309 | v_41490;
assign v_41494 = v_41492 | v_41493;
assign v_41496 = v_41306 | v_41495;
assign v_41499 = v_41497 | v_41498;
assign v_41501 = v_41303 | v_41500;
assign v_41504 = v_41502 | v_41503;
assign v_41506 = v_41300 | v_41505;
assign v_41509 = v_41507 | v_41508;
assign v_41511 = v_41297 | v_41510;
assign v_41514 = v_41512 | v_41513;
assign v_41516 = v_41294 | v_41515;
assign v_41519 = v_41517 | v_41518;
assign v_41521 = v_41291 | v_41520;
assign v_41524 = v_41522 | v_41523;
assign v_41526 = v_41288 | v_41525;
assign v_41529 = v_41287 | v_41528;
assign v_41582 = v_41579 | v_41581;
assign v_41584 = v_41578 | v_41583;
assign v_41586 = v_41576 | v_41585;
assign v_41588 = v_41583 | v_41587;
assign v_41590 = v_41575 | v_41589;
assign v_41592 = v_41573 | v_41591;
assign v_41594 = v_41589 | v_41593;
assign v_41596 = v_41572 | v_41595;
assign v_41598 = v_41570 | v_41597;
assign v_41600 = v_41595 | v_41599;
assign v_41602 = v_41569 | v_41601;
assign v_41604 = v_41567 | v_41603;
assign v_41606 = v_41601 | v_41605;
assign v_41608 = v_41566 | v_41607;
assign v_41610 = v_41564 | v_41609;
assign v_41612 = v_41607 | v_41611;
assign v_41614 = v_41563 | v_41613;
assign v_41616 = v_41561 | v_41615;
assign v_41618 = v_41613 | v_41617;
assign v_41620 = v_41560 | v_41619;
assign v_41622 = v_41558 | v_41621;
assign v_41624 = v_41619 | v_41623;
assign v_41626 = v_41557 | v_41625;
assign v_41628 = v_41555 | v_41627;
assign v_41630 = v_41625 | v_41629;
assign v_41632 = v_41554 | v_41631;
assign v_41634 = v_41552 | v_41633;
assign v_41636 = v_41631 | v_41635;
assign v_41638 = v_41551 | v_41637;
assign v_41640 = v_41549 | v_41639;
assign v_41642 = v_41637 | v_41641;
assign v_41644 = v_41548 | v_41643;
assign v_41646 = v_41546 | v_41645;
assign v_41648 = v_41643 | v_41647;
assign v_41650 = v_41545 | v_41649;
assign v_41652 = v_41543 | v_41651;
assign v_41654 = v_41649 | v_41653;
assign v_41656 = v_41542 | v_41655;
assign v_41658 = v_41540 | v_41657;
assign v_41660 = v_41655 | v_41659;
assign v_41662 = v_41539 | v_41661;
assign v_41664 = v_41537 | v_41663;
assign v_41666 = v_41661 | v_41665;
assign v_41668 = v_41536 | v_41667;
assign v_41670 = v_41534 | v_41669;
assign v_41672 = v_41667 | v_41671;
assign v_41674 = v_41533 | v_41673;
assign v_41676 = v_41531 | v_41675;
assign v_41678 = v_41673 | v_41677;
assign v_41682 = v_41679 | v_41681;
assign v_41689 = v_41578 | v_41688;
assign v_41692 = v_41690 | v_41691;
assign v_41694 = v_41575 | v_41693;
assign v_41697 = v_41695 | v_41696;
assign v_41699 = v_41572 | v_41698;
assign v_41702 = v_41700 | v_41701;
assign v_41704 = v_41569 | v_41703;
assign v_41707 = v_41705 | v_41706;
assign v_41709 = v_41566 | v_41708;
assign v_41712 = v_41710 | v_41711;
assign v_41714 = v_41563 | v_41713;
assign v_41717 = v_41715 | v_41716;
assign v_41719 = v_41560 | v_41718;
assign v_41722 = v_41720 | v_41721;
assign v_41724 = v_41557 | v_41723;
assign v_41727 = v_41725 | v_41726;
assign v_41729 = v_41554 | v_41728;
assign v_41732 = v_41730 | v_41731;
assign v_41734 = v_41551 | v_41733;
assign v_41737 = v_41735 | v_41736;
assign v_41739 = v_41548 | v_41738;
assign v_41742 = v_41740 | v_41741;
assign v_41744 = v_41545 | v_41743;
assign v_41747 = v_41745 | v_41746;
assign v_41749 = v_41542 | v_41748;
assign v_41752 = v_41750 | v_41751;
assign v_41754 = v_41539 | v_41753;
assign v_41757 = v_41755 | v_41756;
assign v_41759 = v_41536 | v_41758;
assign v_41762 = v_41760 | v_41761;
assign v_41764 = v_41533 | v_41763;
assign v_41767 = v_41765 | v_41766;
assign v_41769 = v_41767 | v_41768;
assign v_41772 = v_41530 | v_41771;
assign v_41843 = v_41840 | v_41842;
assign v_41845 = v_41838 | v_41844;
assign v_41847 = v_41836 | v_41846;
assign v_41849 = v_41844 | v_41848;
assign v_41851 = v_41834 | v_41850;
assign v_41853 = v_41832 | v_41852;
assign v_41855 = v_41850 | v_41854;
assign v_41857 = v_41830 | v_41856;
assign v_41859 = v_41828 | v_41858;
assign v_41861 = v_41856 | v_41860;
assign v_41863 = v_41826 | v_41862;
assign v_41865 = v_41824 | v_41864;
assign v_41867 = v_41862 | v_41866;
assign v_41869 = v_41822 | v_41868;
assign v_41871 = v_41820 | v_41870;
assign v_41873 = v_41868 | v_41872;
assign v_41875 = v_41818 | v_41874;
assign v_41877 = v_41816 | v_41876;
assign v_41879 = v_41874 | v_41878;
assign v_41881 = v_41814 | v_41880;
assign v_41883 = v_41812 | v_41882;
assign v_41885 = v_41880 | v_41884;
assign v_41887 = v_41810 | v_41886;
assign v_41889 = v_41808 | v_41888;
assign v_41891 = v_41886 | v_41890;
assign v_41893 = v_41806 | v_41892;
assign v_41895 = v_41804 | v_41894;
assign v_41897 = v_41892 | v_41896;
assign v_41899 = v_41802 | v_41898;
assign v_41901 = v_41800 | v_41900;
assign v_41903 = v_41898 | v_41902;
assign v_41905 = v_41798 | v_41904;
assign v_41907 = v_41796 | v_41906;
assign v_41909 = v_41904 | v_41908;
assign v_41911 = v_41794 | v_41910;
assign v_41913 = v_41792 | v_41912;
assign v_41915 = v_41910 | v_41914;
assign v_41917 = v_41790 | v_41916;
assign v_41919 = v_41787 | v_41918;
assign v_41921 = v_41916 | v_41920;
assign v_41923 = v_41786 | v_41922;
assign v_41925 = v_41783 | v_41924;
assign v_41927 = v_41922 | v_41926;
assign v_41929 = v_41782 | v_41928;
assign v_41931 = v_41779 | v_41930;
assign v_41933 = v_41928 | v_41932;
assign v_41935 = v_41778 | v_41934;
assign v_41937 = v_41775 | v_41936;
assign v_41939 = v_41934 | v_41938;
assign v_41942 = ~v_41774 | v_41941;
assign v_41949 = v_41838 | v_41948;
assign v_41952 = v_41950 | v_41951;
assign v_41954 = v_41834 | v_41953;
assign v_41957 = v_41955 | v_41956;
assign v_41959 = v_41830 | v_41958;
assign v_41962 = v_41960 | v_41961;
assign v_41964 = v_41826 | v_41963;
assign v_41967 = v_41965 | v_41966;
assign v_41969 = v_41822 | v_41968;
assign v_41972 = v_41970 | v_41971;
assign v_41974 = v_41818 | v_41973;
assign v_41977 = v_41975 | v_41976;
assign v_41979 = v_41814 | v_41978;
assign v_41982 = v_41980 | v_41981;
assign v_41984 = v_41810 | v_41983;
assign v_41987 = v_41985 | v_41986;
assign v_41989 = v_41806 | v_41988;
assign v_41992 = v_41990 | v_41991;
assign v_41994 = v_41802 | v_41993;
assign v_41997 = v_41995 | v_41996;
assign v_41999 = v_41798 | v_41998;
assign v_42002 = v_42000 | v_42001;
assign v_42004 = v_41794 | v_42003;
assign v_42007 = v_42005 | v_42006;
assign v_42009 = v_41790 | v_42008;
assign v_42012 = v_42010 | v_42011;
assign v_42014 = v_41786 | v_42013;
assign v_42017 = v_42015 | v_42016;
assign v_42019 = v_41782 | v_42018;
assign v_42022 = v_42020 | v_42021;
assign v_42024 = v_41778 | v_42023;
assign v_42027 = v_42025 | v_42026;
assign v_42029 = v_41774 | v_42028;
assign v_42032 = v_41773 | v_42031;
assign v_42086 = v_42083 | v_42085;
assign v_42088 = v_42082 | v_42087;
assign v_42090 = v_42080 | v_42089;
assign v_42092 = v_42087 | v_42091;
assign v_42094 = v_42079 | v_42093;
assign v_42096 = v_42077 | v_42095;
assign v_42098 = v_42093 | v_42097;
assign v_42100 = v_42076 | v_42099;
assign v_42102 = v_42074 | v_42101;
assign v_42104 = v_42099 | v_42103;
assign v_42106 = v_42073 | v_42105;
assign v_42108 = v_42071 | v_42107;
assign v_42110 = v_42105 | v_42109;
assign v_42112 = v_42070 | v_42111;
assign v_42114 = v_42068 | v_42113;
assign v_42116 = v_42111 | v_42115;
assign v_42118 = v_42067 | v_42117;
assign v_42120 = v_42065 | v_42119;
assign v_42122 = v_42117 | v_42121;
assign v_42124 = v_42064 | v_42123;
assign v_42126 = v_42062 | v_42125;
assign v_42128 = v_42123 | v_42127;
assign v_42130 = v_42061 | v_42129;
assign v_42132 = v_42059 | v_42131;
assign v_42134 = v_42129 | v_42133;
assign v_42136 = v_42058 | v_42135;
assign v_42138 = v_42056 | v_42137;
assign v_42140 = v_42135 | v_42139;
assign v_42142 = v_42055 | v_42141;
assign v_42144 = v_42053 | v_42143;
assign v_42146 = v_42141 | v_42145;
assign v_42148 = v_42052 | v_42147;
assign v_42150 = v_42050 | v_42149;
assign v_42152 = v_42147 | v_42151;
assign v_42154 = v_42049 | v_42153;
assign v_42156 = v_42047 | v_42155;
assign v_42158 = v_42153 | v_42157;
assign v_42160 = v_42046 | v_42159;
assign v_42162 = v_42044 | v_42161;
assign v_42164 = v_42159 | v_42163;
assign v_42166 = v_42043 | v_42165;
assign v_42168 = v_42041 | v_42167;
assign v_42170 = v_42165 | v_42169;
assign v_42172 = v_42040 | v_42171;
assign v_42174 = v_42038 | v_42173;
assign v_42176 = v_42171 | v_42175;
assign v_42178 = v_42037 | v_42177;
assign v_42180 = v_42035 | v_42179;
assign v_42182 = v_42177 | v_42181;
assign v_42185 = ~v_42034 | v_42184;
assign v_42192 = v_42082 | v_42191;
assign v_42195 = v_42193 | v_42194;
assign v_42197 = v_42079 | v_42196;
assign v_42200 = v_42198 | v_42199;
assign v_42202 = v_42076 | v_42201;
assign v_42205 = v_42203 | v_42204;
assign v_42207 = v_42073 | v_42206;
assign v_42210 = v_42208 | v_42209;
assign v_42212 = v_42070 | v_42211;
assign v_42215 = v_42213 | v_42214;
assign v_42217 = v_42067 | v_42216;
assign v_42220 = v_42218 | v_42219;
assign v_42222 = v_42064 | v_42221;
assign v_42225 = v_42223 | v_42224;
assign v_42227 = v_42061 | v_42226;
assign v_42230 = v_42228 | v_42229;
assign v_42232 = v_42058 | v_42231;
assign v_42235 = v_42233 | v_42234;
assign v_42237 = v_42055 | v_42236;
assign v_42240 = v_42238 | v_42239;
assign v_42242 = v_42052 | v_42241;
assign v_42245 = v_42243 | v_42244;
assign v_42247 = v_42049 | v_42246;
assign v_42250 = v_42248 | v_42249;
assign v_42252 = v_42046 | v_42251;
assign v_42255 = v_42253 | v_42254;
assign v_42257 = v_42043 | v_42256;
assign v_42260 = v_42258 | v_42259;
assign v_42262 = v_42040 | v_42261;
assign v_42265 = v_42263 | v_42264;
assign v_42267 = v_42037 | v_42266;
assign v_42270 = v_42268 | v_42269;
assign v_42272 = v_42034 | v_42271;
assign v_42275 = v_42033 | v_42274;
assign v_42329 = v_42326 | v_42328;
assign v_42331 = v_42325 | v_42330;
assign v_42333 = v_42323 | v_42332;
assign v_42335 = v_42330 | v_42334;
assign v_42337 = v_42322 | v_42336;
assign v_42339 = v_42320 | v_42338;
assign v_42341 = v_42336 | v_42340;
assign v_42343 = v_42319 | v_42342;
assign v_42345 = v_42317 | v_42344;
assign v_42347 = v_42342 | v_42346;
assign v_42349 = v_42316 | v_42348;
assign v_42351 = v_42314 | v_42350;
assign v_42353 = v_42348 | v_42352;
assign v_42355 = v_42313 | v_42354;
assign v_42357 = v_42311 | v_42356;
assign v_42359 = v_42354 | v_42358;
assign v_42361 = v_42310 | v_42360;
assign v_42363 = v_42308 | v_42362;
assign v_42365 = v_42360 | v_42364;
assign v_42367 = v_42307 | v_42366;
assign v_42369 = v_42305 | v_42368;
assign v_42371 = v_42366 | v_42370;
assign v_42373 = v_42304 | v_42372;
assign v_42375 = v_42302 | v_42374;
assign v_42377 = v_42372 | v_42376;
assign v_42379 = v_42301 | v_42378;
assign v_42381 = v_42299 | v_42380;
assign v_42383 = v_42378 | v_42382;
assign v_42385 = v_42298 | v_42384;
assign v_42387 = v_42296 | v_42386;
assign v_42389 = v_42384 | v_42388;
assign v_42391 = v_42295 | v_42390;
assign v_42393 = v_42293 | v_42392;
assign v_42395 = v_42390 | v_42394;
assign v_42397 = v_42292 | v_42396;
assign v_42399 = v_42290 | v_42398;
assign v_42401 = v_42396 | v_42400;
assign v_42403 = v_42289 | v_42402;
assign v_42405 = v_42287 | v_42404;
assign v_42407 = v_42402 | v_42406;
assign v_42409 = v_42286 | v_42408;
assign v_42411 = v_42284 | v_42410;
assign v_42413 = v_42408 | v_42412;
assign v_42415 = v_42283 | v_42414;
assign v_42417 = v_42281 | v_42416;
assign v_42419 = v_42414 | v_42418;
assign v_42421 = v_42280 | v_42420;
assign v_42423 = v_42278 | v_42422;
assign v_42425 = v_42420 | v_42424;
assign v_42428 = ~v_42277 | v_42427;
assign v_42435 = v_42325 | v_42434;
assign v_42438 = v_42436 | v_42437;
assign v_42440 = v_42322 | v_42439;
assign v_42443 = v_42441 | v_42442;
assign v_42445 = v_42319 | v_42444;
assign v_42448 = v_42446 | v_42447;
assign v_42450 = v_42316 | v_42449;
assign v_42453 = v_42451 | v_42452;
assign v_42455 = v_42313 | v_42454;
assign v_42458 = v_42456 | v_42457;
assign v_42460 = v_42310 | v_42459;
assign v_42463 = v_42461 | v_42462;
assign v_42465 = v_42307 | v_42464;
assign v_42468 = v_42466 | v_42467;
assign v_42470 = v_42304 | v_42469;
assign v_42473 = v_42471 | v_42472;
assign v_42475 = v_42301 | v_42474;
assign v_42478 = v_42476 | v_42477;
assign v_42480 = v_42298 | v_42479;
assign v_42483 = v_42481 | v_42482;
assign v_42485 = v_42295 | v_42484;
assign v_42488 = v_42486 | v_42487;
assign v_42490 = v_42292 | v_42489;
assign v_42493 = v_42491 | v_42492;
assign v_42495 = v_42289 | v_42494;
assign v_42498 = v_42496 | v_42497;
assign v_42500 = v_42286 | v_42499;
assign v_42503 = v_42501 | v_42502;
assign v_42505 = v_42283 | v_42504;
assign v_42508 = v_42506 | v_42507;
assign v_42510 = v_42280 | v_42509;
assign v_42513 = v_42511 | v_42512;
assign v_42515 = v_42277 | v_42514;
assign v_42518 = v_42276 | v_42517;
assign v_42572 = v_42569 | v_42571;
assign v_42574 = v_42568 | v_42573;
assign v_42576 = v_42566 | v_42575;
assign v_42578 = v_42573 | v_42577;
assign v_42580 = v_42565 | v_42579;
assign v_42582 = v_42563 | v_42581;
assign v_42584 = v_42579 | v_42583;
assign v_42586 = v_42562 | v_42585;
assign v_42588 = v_42560 | v_42587;
assign v_42590 = v_42585 | v_42589;
assign v_42592 = v_42559 | v_42591;
assign v_42594 = v_42557 | v_42593;
assign v_42596 = v_42591 | v_42595;
assign v_42598 = v_42556 | v_42597;
assign v_42600 = v_42554 | v_42599;
assign v_42602 = v_42597 | v_42601;
assign v_42604 = v_42553 | v_42603;
assign v_42606 = v_42551 | v_42605;
assign v_42608 = v_42603 | v_42607;
assign v_42610 = v_42550 | v_42609;
assign v_42612 = v_42548 | v_42611;
assign v_42614 = v_42609 | v_42613;
assign v_42616 = v_42547 | v_42615;
assign v_42618 = v_42545 | v_42617;
assign v_42620 = v_42615 | v_42619;
assign v_42622 = v_42544 | v_42621;
assign v_42624 = v_42542 | v_42623;
assign v_42626 = v_42621 | v_42625;
assign v_42628 = v_42541 | v_42627;
assign v_42630 = v_42539 | v_42629;
assign v_42632 = v_42627 | v_42631;
assign v_42634 = v_42538 | v_42633;
assign v_42636 = v_42536 | v_42635;
assign v_42638 = v_42633 | v_42637;
assign v_42640 = v_42535 | v_42639;
assign v_42642 = v_42533 | v_42641;
assign v_42644 = v_42639 | v_42643;
assign v_42646 = v_42532 | v_42645;
assign v_42648 = v_42530 | v_42647;
assign v_42650 = v_42645 | v_42649;
assign v_42652 = v_42529 | v_42651;
assign v_42654 = v_42527 | v_42653;
assign v_42656 = v_42651 | v_42655;
assign v_42658 = v_42526 | v_42657;
assign v_42660 = v_42524 | v_42659;
assign v_42662 = v_42657 | v_42661;
assign v_42664 = v_42523 | v_42663;
assign v_42666 = v_42521 | v_42665;
assign v_42668 = v_42663 | v_42667;
assign v_42671 = ~v_42520 | v_42670;
assign v_42678 = v_42568 | v_42677;
assign v_42681 = v_42679 | v_42680;
assign v_42683 = v_42565 | v_42682;
assign v_42686 = v_42684 | v_42685;
assign v_42688 = v_42562 | v_42687;
assign v_42691 = v_42689 | v_42690;
assign v_42693 = v_42559 | v_42692;
assign v_42696 = v_42694 | v_42695;
assign v_42698 = v_42556 | v_42697;
assign v_42701 = v_42699 | v_42700;
assign v_42703 = v_42553 | v_42702;
assign v_42706 = v_42704 | v_42705;
assign v_42708 = v_42550 | v_42707;
assign v_42711 = v_42709 | v_42710;
assign v_42713 = v_42547 | v_42712;
assign v_42716 = v_42714 | v_42715;
assign v_42718 = v_42544 | v_42717;
assign v_42721 = v_42719 | v_42720;
assign v_42723 = v_42541 | v_42722;
assign v_42726 = v_42724 | v_42725;
assign v_42728 = v_42538 | v_42727;
assign v_42731 = v_42729 | v_42730;
assign v_42733 = v_42535 | v_42732;
assign v_42736 = v_42734 | v_42735;
assign v_42738 = v_42532 | v_42737;
assign v_42741 = v_42739 | v_42740;
assign v_42743 = v_42529 | v_42742;
assign v_42746 = v_42744 | v_42745;
assign v_42748 = v_42526 | v_42747;
assign v_42751 = v_42749 | v_42750;
assign v_42753 = v_42523 | v_42752;
assign v_42756 = v_42754 | v_42755;
assign v_42758 = v_42520 | v_42757;
assign v_42761 = v_42519 | v_42760;
assign v_42815 = v_42812 | v_42814;
assign v_42817 = v_42811 | v_42816;
assign v_42819 = v_42809 | v_42818;
assign v_42821 = v_42816 | v_42820;
assign v_42823 = v_42808 | v_42822;
assign v_42825 = v_42806 | v_42824;
assign v_42827 = v_42822 | v_42826;
assign v_42829 = v_42805 | v_42828;
assign v_42831 = v_42803 | v_42830;
assign v_42833 = v_42828 | v_42832;
assign v_42835 = v_42802 | v_42834;
assign v_42837 = v_42800 | v_42836;
assign v_42839 = v_42834 | v_42838;
assign v_42841 = v_42799 | v_42840;
assign v_42843 = v_42797 | v_42842;
assign v_42845 = v_42840 | v_42844;
assign v_42847 = v_42796 | v_42846;
assign v_42849 = v_42794 | v_42848;
assign v_42851 = v_42846 | v_42850;
assign v_42853 = v_42793 | v_42852;
assign v_42855 = v_42791 | v_42854;
assign v_42857 = v_42852 | v_42856;
assign v_42859 = v_42790 | v_42858;
assign v_42861 = v_42788 | v_42860;
assign v_42863 = v_42858 | v_42862;
assign v_42865 = v_42787 | v_42864;
assign v_42867 = v_42785 | v_42866;
assign v_42869 = v_42864 | v_42868;
assign v_42871 = v_42784 | v_42870;
assign v_42873 = v_42782 | v_42872;
assign v_42875 = v_42870 | v_42874;
assign v_42877 = v_42781 | v_42876;
assign v_42879 = v_42779 | v_42878;
assign v_42881 = v_42876 | v_42880;
assign v_42883 = v_42778 | v_42882;
assign v_42885 = v_42776 | v_42884;
assign v_42887 = v_42882 | v_42886;
assign v_42889 = v_42775 | v_42888;
assign v_42891 = v_42773 | v_42890;
assign v_42893 = v_42888 | v_42892;
assign v_42895 = v_42772 | v_42894;
assign v_42897 = v_42770 | v_42896;
assign v_42899 = v_42894 | v_42898;
assign v_42901 = v_42769 | v_42900;
assign v_42903 = v_42767 | v_42902;
assign v_42905 = v_42900 | v_42904;
assign v_42907 = v_42766 | v_42906;
assign v_42909 = v_42764 | v_42908;
assign v_42911 = v_42906 | v_42910;
assign v_42914 = ~v_42763 | v_42913;
assign v_42921 = v_42811 | v_42920;
assign v_42924 = v_42922 | v_42923;
assign v_42926 = v_42808 | v_42925;
assign v_42929 = v_42927 | v_42928;
assign v_42931 = v_42805 | v_42930;
assign v_42934 = v_42932 | v_42933;
assign v_42936 = v_42802 | v_42935;
assign v_42939 = v_42937 | v_42938;
assign v_42941 = v_42799 | v_42940;
assign v_42944 = v_42942 | v_42943;
assign v_42946 = v_42796 | v_42945;
assign v_42949 = v_42947 | v_42948;
assign v_42951 = v_42793 | v_42950;
assign v_42954 = v_42952 | v_42953;
assign v_42956 = v_42790 | v_42955;
assign v_42959 = v_42957 | v_42958;
assign v_42961 = v_42787 | v_42960;
assign v_42964 = v_42962 | v_42963;
assign v_42966 = v_42784 | v_42965;
assign v_42969 = v_42967 | v_42968;
assign v_42971 = v_42781 | v_42970;
assign v_42974 = v_42972 | v_42973;
assign v_42976 = v_42778 | v_42975;
assign v_42979 = v_42977 | v_42978;
assign v_42981 = v_42775 | v_42980;
assign v_42984 = v_42982 | v_42983;
assign v_42986 = v_42772 | v_42985;
assign v_42989 = v_42987 | v_42988;
assign v_42991 = v_42769 | v_42990;
assign v_42994 = v_42992 | v_42993;
assign v_42996 = v_42766 | v_42995;
assign v_42999 = v_42997 | v_42998;
assign v_43001 = v_42763 | v_43000;
assign v_43004 = v_42762 | v_43003;
assign v_43058 = v_43055 | v_43057;
assign v_43060 = v_43054 | v_43059;
assign v_43062 = v_43052 | v_43061;
assign v_43064 = v_43059 | v_43063;
assign v_43066 = v_43051 | v_43065;
assign v_43068 = v_43049 | v_43067;
assign v_43070 = v_43065 | v_43069;
assign v_43072 = v_43048 | v_43071;
assign v_43074 = v_43046 | v_43073;
assign v_43076 = v_43071 | v_43075;
assign v_43078 = v_43045 | v_43077;
assign v_43080 = v_43043 | v_43079;
assign v_43082 = v_43077 | v_43081;
assign v_43084 = v_43042 | v_43083;
assign v_43086 = v_43040 | v_43085;
assign v_43088 = v_43083 | v_43087;
assign v_43090 = v_43039 | v_43089;
assign v_43092 = v_43037 | v_43091;
assign v_43094 = v_43089 | v_43093;
assign v_43096 = v_43036 | v_43095;
assign v_43098 = v_43034 | v_43097;
assign v_43100 = v_43095 | v_43099;
assign v_43102 = v_43033 | v_43101;
assign v_43104 = v_43031 | v_43103;
assign v_43106 = v_43101 | v_43105;
assign v_43108 = v_43030 | v_43107;
assign v_43110 = v_43028 | v_43109;
assign v_43112 = v_43107 | v_43111;
assign v_43114 = v_43027 | v_43113;
assign v_43116 = v_43025 | v_43115;
assign v_43118 = v_43113 | v_43117;
assign v_43120 = v_43024 | v_43119;
assign v_43122 = v_43022 | v_43121;
assign v_43124 = v_43119 | v_43123;
assign v_43126 = v_43021 | v_43125;
assign v_43128 = v_43019 | v_43127;
assign v_43130 = v_43125 | v_43129;
assign v_43132 = v_43018 | v_43131;
assign v_43134 = v_43016 | v_43133;
assign v_43136 = v_43131 | v_43135;
assign v_43138 = v_43015 | v_43137;
assign v_43140 = v_43013 | v_43139;
assign v_43142 = v_43137 | v_43141;
assign v_43144 = v_43012 | v_43143;
assign v_43146 = v_43010 | v_43145;
assign v_43148 = v_43143 | v_43147;
assign v_43150 = v_43009 | v_43149;
assign v_43152 = v_43007 | v_43151;
assign v_43154 = v_43149 | v_43153;
assign v_43157 = ~v_43006 | v_43156;
assign v_43164 = v_43054 | v_43163;
assign v_43167 = v_43165 | v_43166;
assign v_43169 = v_43051 | v_43168;
assign v_43172 = v_43170 | v_43171;
assign v_43174 = v_43048 | v_43173;
assign v_43177 = v_43175 | v_43176;
assign v_43179 = v_43045 | v_43178;
assign v_43182 = v_43180 | v_43181;
assign v_43184 = v_43042 | v_43183;
assign v_43187 = v_43185 | v_43186;
assign v_43189 = v_43039 | v_43188;
assign v_43192 = v_43190 | v_43191;
assign v_43194 = v_43036 | v_43193;
assign v_43197 = v_43195 | v_43196;
assign v_43199 = v_43033 | v_43198;
assign v_43202 = v_43200 | v_43201;
assign v_43204 = v_43030 | v_43203;
assign v_43207 = v_43205 | v_43206;
assign v_43209 = v_43027 | v_43208;
assign v_43212 = v_43210 | v_43211;
assign v_43214 = v_43024 | v_43213;
assign v_43217 = v_43215 | v_43216;
assign v_43219 = v_43021 | v_43218;
assign v_43222 = v_43220 | v_43221;
assign v_43224 = v_43018 | v_43223;
assign v_43227 = v_43225 | v_43226;
assign v_43229 = v_43015 | v_43228;
assign v_43232 = v_43230 | v_43231;
assign v_43234 = v_43012 | v_43233;
assign v_43237 = v_43235 | v_43236;
assign v_43239 = v_43009 | v_43238;
assign v_43242 = v_43240 | v_43241;
assign v_43244 = v_43006 | v_43243;
assign v_43247 = v_43005 | v_43246;
assign v_43301 = v_43298 | v_43300;
assign v_43303 = v_43297 | v_43302;
assign v_43305 = v_43295 | v_43304;
assign v_43307 = v_43302 | v_43306;
assign v_43309 = v_43294 | v_43308;
assign v_43311 = v_43292 | v_43310;
assign v_43313 = v_43308 | v_43312;
assign v_43315 = v_43291 | v_43314;
assign v_43317 = v_43289 | v_43316;
assign v_43319 = v_43314 | v_43318;
assign v_43321 = v_43288 | v_43320;
assign v_43323 = v_43286 | v_43322;
assign v_43325 = v_43320 | v_43324;
assign v_43327 = v_43285 | v_43326;
assign v_43329 = v_43283 | v_43328;
assign v_43331 = v_43326 | v_43330;
assign v_43333 = v_43282 | v_43332;
assign v_43335 = v_43280 | v_43334;
assign v_43337 = v_43332 | v_43336;
assign v_43339 = v_43279 | v_43338;
assign v_43341 = v_43277 | v_43340;
assign v_43343 = v_43338 | v_43342;
assign v_43345 = v_43276 | v_43344;
assign v_43347 = v_43274 | v_43346;
assign v_43349 = v_43344 | v_43348;
assign v_43351 = v_43273 | v_43350;
assign v_43353 = v_43271 | v_43352;
assign v_43355 = v_43350 | v_43354;
assign v_43357 = v_43270 | v_43356;
assign v_43359 = v_43268 | v_43358;
assign v_43361 = v_43356 | v_43360;
assign v_43363 = v_43267 | v_43362;
assign v_43365 = v_43265 | v_43364;
assign v_43367 = v_43362 | v_43366;
assign v_43369 = v_43264 | v_43368;
assign v_43371 = v_43262 | v_43370;
assign v_43373 = v_43368 | v_43372;
assign v_43375 = v_43261 | v_43374;
assign v_43377 = v_43259 | v_43376;
assign v_43379 = v_43374 | v_43378;
assign v_43381 = v_43258 | v_43380;
assign v_43383 = v_43256 | v_43382;
assign v_43385 = v_43380 | v_43384;
assign v_43387 = v_43255 | v_43386;
assign v_43389 = v_43253 | v_43388;
assign v_43391 = v_43386 | v_43390;
assign v_43393 = v_43252 | v_43392;
assign v_43395 = v_43250 | v_43394;
assign v_43397 = v_43392 | v_43396;
assign v_43400 = ~v_43249 | v_43399;
assign v_43407 = v_43297 | v_43406;
assign v_43410 = v_43408 | v_43409;
assign v_43412 = v_43294 | v_43411;
assign v_43415 = v_43413 | v_43414;
assign v_43417 = v_43291 | v_43416;
assign v_43420 = v_43418 | v_43419;
assign v_43422 = v_43288 | v_43421;
assign v_43425 = v_43423 | v_43424;
assign v_43427 = v_43285 | v_43426;
assign v_43430 = v_43428 | v_43429;
assign v_43432 = v_43282 | v_43431;
assign v_43435 = v_43433 | v_43434;
assign v_43437 = v_43279 | v_43436;
assign v_43440 = v_43438 | v_43439;
assign v_43442 = v_43276 | v_43441;
assign v_43445 = v_43443 | v_43444;
assign v_43447 = v_43273 | v_43446;
assign v_43450 = v_43448 | v_43449;
assign v_43452 = v_43270 | v_43451;
assign v_43455 = v_43453 | v_43454;
assign v_43457 = v_43267 | v_43456;
assign v_43460 = v_43458 | v_43459;
assign v_43462 = v_43264 | v_43461;
assign v_43465 = v_43463 | v_43464;
assign v_43467 = v_43261 | v_43466;
assign v_43470 = v_43468 | v_43469;
assign v_43472 = v_43258 | v_43471;
assign v_43475 = v_43473 | v_43474;
assign v_43477 = v_43255 | v_43476;
assign v_43480 = v_43478 | v_43479;
assign v_43482 = v_43252 | v_43481;
assign v_43485 = v_43483 | v_43484;
assign v_43487 = v_43249 | v_43486;
assign v_43490 = v_43248 | v_43489;
assign v_43544 = v_43541 | v_43543;
assign v_43546 = v_43540 | v_43545;
assign v_43548 = v_43538 | v_43547;
assign v_43550 = v_43545 | v_43549;
assign v_43552 = v_43537 | v_43551;
assign v_43554 = v_43535 | v_43553;
assign v_43556 = v_43551 | v_43555;
assign v_43558 = v_43534 | v_43557;
assign v_43560 = v_43532 | v_43559;
assign v_43562 = v_43557 | v_43561;
assign v_43564 = v_43531 | v_43563;
assign v_43566 = v_43529 | v_43565;
assign v_43568 = v_43563 | v_43567;
assign v_43570 = v_43528 | v_43569;
assign v_43572 = v_43526 | v_43571;
assign v_43574 = v_43569 | v_43573;
assign v_43576 = v_43525 | v_43575;
assign v_43578 = v_43523 | v_43577;
assign v_43580 = v_43575 | v_43579;
assign v_43582 = v_43522 | v_43581;
assign v_43584 = v_43520 | v_43583;
assign v_43586 = v_43581 | v_43585;
assign v_43588 = v_43519 | v_43587;
assign v_43590 = v_43517 | v_43589;
assign v_43592 = v_43587 | v_43591;
assign v_43594 = v_43516 | v_43593;
assign v_43596 = v_43514 | v_43595;
assign v_43598 = v_43593 | v_43597;
assign v_43600 = v_43513 | v_43599;
assign v_43602 = v_43511 | v_43601;
assign v_43604 = v_43599 | v_43603;
assign v_43606 = v_43510 | v_43605;
assign v_43608 = v_43508 | v_43607;
assign v_43610 = v_43605 | v_43609;
assign v_43612 = v_43507 | v_43611;
assign v_43614 = v_43505 | v_43613;
assign v_43616 = v_43611 | v_43615;
assign v_43618 = v_43504 | v_43617;
assign v_43620 = v_43502 | v_43619;
assign v_43622 = v_43617 | v_43621;
assign v_43624 = v_43501 | v_43623;
assign v_43626 = v_43499 | v_43625;
assign v_43628 = v_43623 | v_43627;
assign v_43630 = v_43498 | v_43629;
assign v_43632 = v_43496 | v_43631;
assign v_43634 = v_43629 | v_43633;
assign v_43636 = v_43495 | v_43635;
assign v_43638 = v_43493 | v_43637;
assign v_43640 = v_43635 | v_43639;
assign v_43643 = ~v_43492 | v_43642;
assign v_43650 = v_43540 | v_43649;
assign v_43653 = v_43651 | v_43652;
assign v_43655 = v_43537 | v_43654;
assign v_43658 = v_43656 | v_43657;
assign v_43660 = v_43534 | v_43659;
assign v_43663 = v_43661 | v_43662;
assign v_43665 = v_43531 | v_43664;
assign v_43668 = v_43666 | v_43667;
assign v_43670 = v_43528 | v_43669;
assign v_43673 = v_43671 | v_43672;
assign v_43675 = v_43525 | v_43674;
assign v_43678 = v_43676 | v_43677;
assign v_43680 = v_43522 | v_43679;
assign v_43683 = v_43681 | v_43682;
assign v_43685 = v_43519 | v_43684;
assign v_43688 = v_43686 | v_43687;
assign v_43690 = v_43516 | v_43689;
assign v_43693 = v_43691 | v_43692;
assign v_43695 = v_43513 | v_43694;
assign v_43698 = v_43696 | v_43697;
assign v_43700 = v_43510 | v_43699;
assign v_43703 = v_43701 | v_43702;
assign v_43705 = v_43507 | v_43704;
assign v_43708 = v_43706 | v_43707;
assign v_43710 = v_43504 | v_43709;
assign v_43713 = v_43711 | v_43712;
assign v_43715 = v_43501 | v_43714;
assign v_43718 = v_43716 | v_43717;
assign v_43720 = v_43498 | v_43719;
assign v_43723 = v_43721 | v_43722;
assign v_43725 = v_43495 | v_43724;
assign v_43728 = v_43726 | v_43727;
assign v_43730 = v_43492 | v_43729;
assign v_43733 = v_43491 | v_43732;
assign v_43787 = v_43784 | v_43786;
assign v_43789 = v_43783 | v_43788;
assign v_43791 = v_43781 | v_43790;
assign v_43793 = v_43788 | v_43792;
assign v_43795 = v_43780 | v_43794;
assign v_43797 = v_43778 | v_43796;
assign v_43799 = v_43794 | v_43798;
assign v_43801 = v_43777 | v_43800;
assign v_43803 = v_43775 | v_43802;
assign v_43805 = v_43800 | v_43804;
assign v_43807 = v_43774 | v_43806;
assign v_43809 = v_43772 | v_43808;
assign v_43811 = v_43806 | v_43810;
assign v_43813 = v_43771 | v_43812;
assign v_43815 = v_43769 | v_43814;
assign v_43817 = v_43812 | v_43816;
assign v_43819 = v_43768 | v_43818;
assign v_43821 = v_43766 | v_43820;
assign v_43823 = v_43818 | v_43822;
assign v_43825 = v_43765 | v_43824;
assign v_43827 = v_43763 | v_43826;
assign v_43829 = v_43824 | v_43828;
assign v_43831 = v_43762 | v_43830;
assign v_43833 = v_43760 | v_43832;
assign v_43835 = v_43830 | v_43834;
assign v_43837 = v_43759 | v_43836;
assign v_43839 = v_43757 | v_43838;
assign v_43841 = v_43836 | v_43840;
assign v_43843 = v_43756 | v_43842;
assign v_43845 = v_43754 | v_43844;
assign v_43847 = v_43842 | v_43846;
assign v_43849 = v_43753 | v_43848;
assign v_43851 = v_43751 | v_43850;
assign v_43853 = v_43848 | v_43852;
assign v_43855 = v_43750 | v_43854;
assign v_43857 = v_43748 | v_43856;
assign v_43859 = v_43854 | v_43858;
assign v_43861 = v_43747 | v_43860;
assign v_43863 = v_43745 | v_43862;
assign v_43865 = v_43860 | v_43864;
assign v_43867 = v_43744 | v_43866;
assign v_43869 = v_43742 | v_43868;
assign v_43871 = v_43866 | v_43870;
assign v_43873 = v_43741 | v_43872;
assign v_43875 = v_43739 | v_43874;
assign v_43877 = v_43872 | v_43876;
assign v_43879 = v_43738 | v_43878;
assign v_43881 = v_43736 | v_43880;
assign v_43883 = v_43878 | v_43882;
assign v_43886 = ~v_43735 | v_43885;
assign v_43893 = v_43783 | v_43892;
assign v_43896 = v_43894 | v_43895;
assign v_43898 = v_43780 | v_43897;
assign v_43901 = v_43899 | v_43900;
assign v_43903 = v_43777 | v_43902;
assign v_43906 = v_43904 | v_43905;
assign v_43908 = v_43774 | v_43907;
assign v_43911 = v_43909 | v_43910;
assign v_43913 = v_43771 | v_43912;
assign v_43916 = v_43914 | v_43915;
assign v_43918 = v_43768 | v_43917;
assign v_43921 = v_43919 | v_43920;
assign v_43923 = v_43765 | v_43922;
assign v_43926 = v_43924 | v_43925;
assign v_43928 = v_43762 | v_43927;
assign v_43931 = v_43929 | v_43930;
assign v_43933 = v_43759 | v_43932;
assign v_43936 = v_43934 | v_43935;
assign v_43938 = v_43756 | v_43937;
assign v_43941 = v_43939 | v_43940;
assign v_43943 = v_43753 | v_43942;
assign v_43946 = v_43944 | v_43945;
assign v_43948 = v_43750 | v_43947;
assign v_43951 = v_43949 | v_43950;
assign v_43953 = v_43747 | v_43952;
assign v_43956 = v_43954 | v_43955;
assign v_43958 = v_43744 | v_43957;
assign v_43961 = v_43959 | v_43960;
assign v_43963 = v_43741 | v_43962;
assign v_43966 = v_43964 | v_43965;
assign v_43968 = v_43738 | v_43967;
assign v_43971 = v_43969 | v_43970;
assign v_43973 = v_43735 | v_43972;
assign v_43976 = v_43734 | v_43975;
assign v_44030 = v_44027 | v_44029;
assign v_44032 = v_44026 | v_44031;
assign v_44034 = v_44024 | v_44033;
assign v_44036 = v_44031 | v_44035;
assign v_44038 = v_44023 | v_44037;
assign v_44040 = v_44021 | v_44039;
assign v_44042 = v_44037 | v_44041;
assign v_44044 = v_44020 | v_44043;
assign v_44046 = v_44018 | v_44045;
assign v_44048 = v_44043 | v_44047;
assign v_44050 = v_44017 | v_44049;
assign v_44052 = v_44015 | v_44051;
assign v_44054 = v_44049 | v_44053;
assign v_44056 = v_44014 | v_44055;
assign v_44058 = v_44012 | v_44057;
assign v_44060 = v_44055 | v_44059;
assign v_44062 = v_44011 | v_44061;
assign v_44064 = v_44009 | v_44063;
assign v_44066 = v_44061 | v_44065;
assign v_44068 = v_44008 | v_44067;
assign v_44070 = v_44006 | v_44069;
assign v_44072 = v_44067 | v_44071;
assign v_44074 = v_44005 | v_44073;
assign v_44076 = v_44003 | v_44075;
assign v_44078 = v_44073 | v_44077;
assign v_44080 = v_44002 | v_44079;
assign v_44082 = v_44000 | v_44081;
assign v_44084 = v_44079 | v_44083;
assign v_44086 = v_43999 | v_44085;
assign v_44088 = v_43997 | v_44087;
assign v_44090 = v_44085 | v_44089;
assign v_44092 = v_43996 | v_44091;
assign v_44094 = v_43994 | v_44093;
assign v_44096 = v_44091 | v_44095;
assign v_44098 = v_43993 | v_44097;
assign v_44100 = v_43991 | v_44099;
assign v_44102 = v_44097 | v_44101;
assign v_44104 = v_43990 | v_44103;
assign v_44106 = v_43988 | v_44105;
assign v_44108 = v_44103 | v_44107;
assign v_44110 = v_43987 | v_44109;
assign v_44112 = v_43985 | v_44111;
assign v_44114 = v_44109 | v_44113;
assign v_44116 = v_43984 | v_44115;
assign v_44118 = v_43982 | v_44117;
assign v_44120 = v_44115 | v_44119;
assign v_44122 = v_43981 | v_44121;
assign v_44124 = v_43979 | v_44123;
assign v_44126 = v_44121 | v_44125;
assign v_44129 = ~v_43978 | v_44128;
assign v_44136 = v_44026 | v_44135;
assign v_44139 = v_44137 | v_44138;
assign v_44141 = v_44023 | v_44140;
assign v_44144 = v_44142 | v_44143;
assign v_44146 = v_44020 | v_44145;
assign v_44149 = v_44147 | v_44148;
assign v_44151 = v_44017 | v_44150;
assign v_44154 = v_44152 | v_44153;
assign v_44156 = v_44014 | v_44155;
assign v_44159 = v_44157 | v_44158;
assign v_44161 = v_44011 | v_44160;
assign v_44164 = v_44162 | v_44163;
assign v_44166 = v_44008 | v_44165;
assign v_44169 = v_44167 | v_44168;
assign v_44171 = v_44005 | v_44170;
assign v_44174 = v_44172 | v_44173;
assign v_44176 = v_44002 | v_44175;
assign v_44179 = v_44177 | v_44178;
assign v_44181 = v_43999 | v_44180;
assign v_44184 = v_44182 | v_44183;
assign v_44186 = v_43996 | v_44185;
assign v_44189 = v_44187 | v_44188;
assign v_44191 = v_43993 | v_44190;
assign v_44194 = v_44192 | v_44193;
assign v_44196 = v_43990 | v_44195;
assign v_44199 = v_44197 | v_44198;
assign v_44201 = v_43987 | v_44200;
assign v_44204 = v_44202 | v_44203;
assign v_44206 = v_43984 | v_44205;
assign v_44209 = v_44207 | v_44208;
assign v_44211 = v_43981 | v_44210;
assign v_44214 = v_44212 | v_44213;
assign v_44216 = v_43978 | v_44215;
assign v_44219 = v_43977 | v_44218;
assign v_44273 = v_44270 | v_44272;
assign v_44275 = v_44269 | v_44274;
assign v_44277 = v_44267 | v_44276;
assign v_44279 = v_44274 | v_44278;
assign v_44281 = v_44266 | v_44280;
assign v_44283 = v_44264 | v_44282;
assign v_44285 = v_44280 | v_44284;
assign v_44287 = v_44263 | v_44286;
assign v_44289 = v_44261 | v_44288;
assign v_44291 = v_44286 | v_44290;
assign v_44293 = v_44260 | v_44292;
assign v_44295 = v_44258 | v_44294;
assign v_44297 = v_44292 | v_44296;
assign v_44299 = v_44257 | v_44298;
assign v_44301 = v_44255 | v_44300;
assign v_44303 = v_44298 | v_44302;
assign v_44305 = v_44254 | v_44304;
assign v_44307 = v_44252 | v_44306;
assign v_44309 = v_44304 | v_44308;
assign v_44311 = v_44251 | v_44310;
assign v_44313 = v_44249 | v_44312;
assign v_44315 = v_44310 | v_44314;
assign v_44317 = v_44248 | v_44316;
assign v_44319 = v_44246 | v_44318;
assign v_44321 = v_44316 | v_44320;
assign v_44323 = v_44245 | v_44322;
assign v_44325 = v_44243 | v_44324;
assign v_44327 = v_44322 | v_44326;
assign v_44329 = v_44242 | v_44328;
assign v_44331 = v_44240 | v_44330;
assign v_44333 = v_44328 | v_44332;
assign v_44335 = v_44239 | v_44334;
assign v_44337 = v_44237 | v_44336;
assign v_44339 = v_44334 | v_44338;
assign v_44341 = v_44236 | v_44340;
assign v_44343 = v_44234 | v_44342;
assign v_44345 = v_44340 | v_44344;
assign v_44347 = v_44233 | v_44346;
assign v_44349 = v_44231 | v_44348;
assign v_44351 = v_44346 | v_44350;
assign v_44353 = v_44230 | v_44352;
assign v_44355 = v_44228 | v_44354;
assign v_44357 = v_44352 | v_44356;
assign v_44359 = v_44227 | v_44358;
assign v_44361 = v_44225 | v_44360;
assign v_44363 = v_44358 | v_44362;
assign v_44365 = v_44224 | v_44364;
assign v_44367 = v_44222 | v_44366;
assign v_44369 = v_44364 | v_44368;
assign v_44372 = ~v_44221 | v_44371;
assign v_44379 = v_44269 | v_44378;
assign v_44382 = v_44380 | v_44381;
assign v_44384 = v_44266 | v_44383;
assign v_44387 = v_44385 | v_44386;
assign v_44389 = v_44263 | v_44388;
assign v_44392 = v_44390 | v_44391;
assign v_44394 = v_44260 | v_44393;
assign v_44397 = v_44395 | v_44396;
assign v_44399 = v_44257 | v_44398;
assign v_44402 = v_44400 | v_44401;
assign v_44404 = v_44254 | v_44403;
assign v_44407 = v_44405 | v_44406;
assign v_44409 = v_44251 | v_44408;
assign v_44412 = v_44410 | v_44411;
assign v_44414 = v_44248 | v_44413;
assign v_44417 = v_44415 | v_44416;
assign v_44419 = v_44245 | v_44418;
assign v_44422 = v_44420 | v_44421;
assign v_44424 = v_44242 | v_44423;
assign v_44427 = v_44425 | v_44426;
assign v_44429 = v_44239 | v_44428;
assign v_44432 = v_44430 | v_44431;
assign v_44434 = v_44236 | v_44433;
assign v_44437 = v_44435 | v_44436;
assign v_44439 = v_44233 | v_44438;
assign v_44442 = v_44440 | v_44441;
assign v_44444 = v_44230 | v_44443;
assign v_44447 = v_44445 | v_44446;
assign v_44449 = v_44227 | v_44448;
assign v_44452 = v_44450 | v_44451;
assign v_44454 = v_44224 | v_44453;
assign v_44457 = v_44455 | v_44456;
assign v_44459 = v_44221 | v_44458;
assign v_44462 = v_44220 | v_44461;
assign v_44516 = v_44513 | v_44515;
assign v_44518 = v_44512 | v_44517;
assign v_44520 = v_44510 | v_44519;
assign v_44522 = v_44517 | v_44521;
assign v_44524 = v_44509 | v_44523;
assign v_44526 = v_44507 | v_44525;
assign v_44528 = v_44523 | v_44527;
assign v_44530 = v_44506 | v_44529;
assign v_44532 = v_44504 | v_44531;
assign v_44534 = v_44529 | v_44533;
assign v_44536 = v_44503 | v_44535;
assign v_44538 = v_44501 | v_44537;
assign v_44540 = v_44535 | v_44539;
assign v_44542 = v_44500 | v_44541;
assign v_44544 = v_44498 | v_44543;
assign v_44546 = v_44541 | v_44545;
assign v_44548 = v_44497 | v_44547;
assign v_44550 = v_44495 | v_44549;
assign v_44552 = v_44547 | v_44551;
assign v_44554 = v_44494 | v_44553;
assign v_44556 = v_44492 | v_44555;
assign v_44558 = v_44553 | v_44557;
assign v_44560 = v_44491 | v_44559;
assign v_44562 = v_44489 | v_44561;
assign v_44564 = v_44559 | v_44563;
assign v_44566 = v_44488 | v_44565;
assign v_44568 = v_44486 | v_44567;
assign v_44570 = v_44565 | v_44569;
assign v_44572 = v_44485 | v_44571;
assign v_44574 = v_44483 | v_44573;
assign v_44576 = v_44571 | v_44575;
assign v_44578 = v_44482 | v_44577;
assign v_44580 = v_44480 | v_44579;
assign v_44582 = v_44577 | v_44581;
assign v_44584 = v_44479 | v_44583;
assign v_44586 = v_44477 | v_44585;
assign v_44588 = v_44583 | v_44587;
assign v_44590 = v_44476 | v_44589;
assign v_44592 = v_44474 | v_44591;
assign v_44594 = v_44589 | v_44593;
assign v_44596 = v_44473 | v_44595;
assign v_44598 = v_44471 | v_44597;
assign v_44600 = v_44595 | v_44599;
assign v_44602 = v_44470 | v_44601;
assign v_44604 = v_44468 | v_44603;
assign v_44606 = v_44601 | v_44605;
assign v_44608 = v_44467 | v_44607;
assign v_44610 = v_44465 | v_44609;
assign v_44612 = v_44607 | v_44611;
assign v_44615 = ~v_44464 | v_44614;
assign v_44622 = v_44512 | v_44621;
assign v_44625 = v_44623 | v_44624;
assign v_44627 = v_44509 | v_44626;
assign v_44630 = v_44628 | v_44629;
assign v_44632 = v_44506 | v_44631;
assign v_44635 = v_44633 | v_44634;
assign v_44637 = v_44503 | v_44636;
assign v_44640 = v_44638 | v_44639;
assign v_44642 = v_44500 | v_44641;
assign v_44645 = v_44643 | v_44644;
assign v_44647 = v_44497 | v_44646;
assign v_44650 = v_44648 | v_44649;
assign v_44652 = v_44494 | v_44651;
assign v_44655 = v_44653 | v_44654;
assign v_44657 = v_44491 | v_44656;
assign v_44660 = v_44658 | v_44659;
assign v_44662 = v_44488 | v_44661;
assign v_44665 = v_44663 | v_44664;
assign v_44667 = v_44485 | v_44666;
assign v_44670 = v_44668 | v_44669;
assign v_44672 = v_44482 | v_44671;
assign v_44675 = v_44673 | v_44674;
assign v_44677 = v_44479 | v_44676;
assign v_44680 = v_44678 | v_44679;
assign v_44682 = v_44476 | v_44681;
assign v_44685 = v_44683 | v_44684;
assign v_44687 = v_44473 | v_44686;
assign v_44690 = v_44688 | v_44689;
assign v_44692 = v_44470 | v_44691;
assign v_44695 = v_44693 | v_44694;
assign v_44697 = v_44467 | v_44696;
assign v_44700 = v_44698 | v_44699;
assign v_44702 = v_44464 | v_44701;
assign v_44705 = v_44463 | v_44704;
assign v_44759 = v_44756 | v_44758;
assign v_44761 = v_44755 | v_44760;
assign v_44763 = v_44753 | v_44762;
assign v_44765 = v_44760 | v_44764;
assign v_44767 = v_44752 | v_44766;
assign v_44769 = v_44750 | v_44768;
assign v_44771 = v_44766 | v_44770;
assign v_44773 = v_44749 | v_44772;
assign v_44775 = v_44747 | v_44774;
assign v_44777 = v_44772 | v_44776;
assign v_44779 = v_44746 | v_44778;
assign v_44781 = v_44744 | v_44780;
assign v_44783 = v_44778 | v_44782;
assign v_44785 = v_44743 | v_44784;
assign v_44787 = v_44741 | v_44786;
assign v_44789 = v_44784 | v_44788;
assign v_44791 = v_44740 | v_44790;
assign v_44793 = v_44738 | v_44792;
assign v_44795 = v_44790 | v_44794;
assign v_44797 = v_44737 | v_44796;
assign v_44799 = v_44735 | v_44798;
assign v_44801 = v_44796 | v_44800;
assign v_44803 = v_44734 | v_44802;
assign v_44805 = v_44732 | v_44804;
assign v_44807 = v_44802 | v_44806;
assign v_44809 = v_44731 | v_44808;
assign v_44811 = v_44729 | v_44810;
assign v_44813 = v_44808 | v_44812;
assign v_44815 = v_44728 | v_44814;
assign v_44817 = v_44726 | v_44816;
assign v_44819 = v_44814 | v_44818;
assign v_44821 = v_44725 | v_44820;
assign v_44823 = v_44723 | v_44822;
assign v_44825 = v_44820 | v_44824;
assign v_44827 = v_44722 | v_44826;
assign v_44829 = v_44720 | v_44828;
assign v_44831 = v_44826 | v_44830;
assign v_44833 = v_44719 | v_44832;
assign v_44835 = v_44717 | v_44834;
assign v_44837 = v_44832 | v_44836;
assign v_44839 = v_44716 | v_44838;
assign v_44841 = v_44714 | v_44840;
assign v_44843 = v_44838 | v_44842;
assign v_44845 = v_44713 | v_44844;
assign v_44847 = v_44711 | v_44846;
assign v_44849 = v_44844 | v_44848;
assign v_44851 = v_44710 | v_44850;
assign v_44853 = v_44708 | v_44852;
assign v_44855 = v_44850 | v_44854;
assign v_44858 = ~v_44707 | v_44857;
assign v_44865 = v_44755 | v_44864;
assign v_44868 = v_44866 | v_44867;
assign v_44870 = v_44752 | v_44869;
assign v_44873 = v_44871 | v_44872;
assign v_44875 = v_44749 | v_44874;
assign v_44878 = v_44876 | v_44877;
assign v_44880 = v_44746 | v_44879;
assign v_44883 = v_44881 | v_44882;
assign v_44885 = v_44743 | v_44884;
assign v_44888 = v_44886 | v_44887;
assign v_44890 = v_44740 | v_44889;
assign v_44893 = v_44891 | v_44892;
assign v_44895 = v_44737 | v_44894;
assign v_44898 = v_44896 | v_44897;
assign v_44900 = v_44734 | v_44899;
assign v_44903 = v_44901 | v_44902;
assign v_44905 = v_44731 | v_44904;
assign v_44908 = v_44906 | v_44907;
assign v_44910 = v_44728 | v_44909;
assign v_44913 = v_44911 | v_44912;
assign v_44915 = v_44725 | v_44914;
assign v_44918 = v_44916 | v_44917;
assign v_44920 = v_44722 | v_44919;
assign v_44923 = v_44921 | v_44922;
assign v_44925 = v_44719 | v_44924;
assign v_44928 = v_44926 | v_44927;
assign v_44930 = v_44716 | v_44929;
assign v_44933 = v_44931 | v_44932;
assign v_44935 = v_44713 | v_44934;
assign v_44938 = v_44936 | v_44937;
assign v_44940 = v_44710 | v_44939;
assign v_44943 = v_44941 | v_44942;
assign v_44945 = v_44707 | v_44944;
assign v_44948 = v_44706 | v_44947;
assign v_45002 = v_44999 | v_45001;
assign v_45004 = v_44998 | v_45003;
assign v_45006 = v_44996 | v_45005;
assign v_45008 = v_45003 | v_45007;
assign v_45010 = v_44995 | v_45009;
assign v_45012 = v_44993 | v_45011;
assign v_45014 = v_45009 | v_45013;
assign v_45016 = v_44992 | v_45015;
assign v_45018 = v_44990 | v_45017;
assign v_45020 = v_45015 | v_45019;
assign v_45022 = v_44989 | v_45021;
assign v_45024 = v_44987 | v_45023;
assign v_45026 = v_45021 | v_45025;
assign v_45028 = v_44986 | v_45027;
assign v_45030 = v_44984 | v_45029;
assign v_45032 = v_45027 | v_45031;
assign v_45034 = v_44983 | v_45033;
assign v_45036 = v_44981 | v_45035;
assign v_45038 = v_45033 | v_45037;
assign v_45040 = v_44980 | v_45039;
assign v_45042 = v_44978 | v_45041;
assign v_45044 = v_45039 | v_45043;
assign v_45046 = v_44977 | v_45045;
assign v_45048 = v_44975 | v_45047;
assign v_45050 = v_45045 | v_45049;
assign v_45052 = v_44974 | v_45051;
assign v_45054 = v_44972 | v_45053;
assign v_45056 = v_45051 | v_45055;
assign v_45058 = v_44971 | v_45057;
assign v_45060 = v_44969 | v_45059;
assign v_45062 = v_45057 | v_45061;
assign v_45064 = v_44968 | v_45063;
assign v_45066 = v_44966 | v_45065;
assign v_45068 = v_45063 | v_45067;
assign v_45070 = v_44965 | v_45069;
assign v_45072 = v_44963 | v_45071;
assign v_45074 = v_45069 | v_45073;
assign v_45076 = v_44962 | v_45075;
assign v_45078 = v_44960 | v_45077;
assign v_45080 = v_45075 | v_45079;
assign v_45082 = v_44959 | v_45081;
assign v_45084 = v_44957 | v_45083;
assign v_45086 = v_45081 | v_45085;
assign v_45088 = v_44956 | v_45087;
assign v_45090 = v_44954 | v_45089;
assign v_45092 = v_45087 | v_45091;
assign v_45094 = v_44953 | v_45093;
assign v_45096 = v_44951 | v_45095;
assign v_45098 = v_45093 | v_45097;
assign v_45101 = ~v_44950 | v_45100;
assign v_45108 = v_44998 | v_45107;
assign v_45111 = v_45109 | v_45110;
assign v_45113 = v_44995 | v_45112;
assign v_45116 = v_45114 | v_45115;
assign v_45118 = v_44992 | v_45117;
assign v_45121 = v_45119 | v_45120;
assign v_45123 = v_44989 | v_45122;
assign v_45126 = v_45124 | v_45125;
assign v_45128 = v_44986 | v_45127;
assign v_45131 = v_45129 | v_45130;
assign v_45133 = v_44983 | v_45132;
assign v_45136 = v_45134 | v_45135;
assign v_45138 = v_44980 | v_45137;
assign v_45141 = v_45139 | v_45140;
assign v_45143 = v_44977 | v_45142;
assign v_45146 = v_45144 | v_45145;
assign v_45148 = v_44974 | v_45147;
assign v_45151 = v_45149 | v_45150;
assign v_45153 = v_44971 | v_45152;
assign v_45156 = v_45154 | v_45155;
assign v_45158 = v_44968 | v_45157;
assign v_45161 = v_45159 | v_45160;
assign v_45163 = v_44965 | v_45162;
assign v_45166 = v_45164 | v_45165;
assign v_45168 = v_44962 | v_45167;
assign v_45171 = v_45169 | v_45170;
assign v_45173 = v_44959 | v_45172;
assign v_45176 = v_45174 | v_45175;
assign v_45178 = v_44956 | v_45177;
assign v_45181 = v_45179 | v_45180;
assign v_45183 = v_44953 | v_45182;
assign v_45186 = v_45184 | v_45185;
assign v_45188 = v_44950 | v_45187;
assign v_45191 = v_44949 | v_45190;
assign v_45245 = v_45242 | v_45244;
assign v_45247 = v_45241 | v_45246;
assign v_45249 = v_45239 | v_45248;
assign v_45251 = v_45246 | v_45250;
assign v_45253 = v_45238 | v_45252;
assign v_45255 = v_45236 | v_45254;
assign v_45257 = v_45252 | v_45256;
assign v_45259 = v_45235 | v_45258;
assign v_45261 = v_45233 | v_45260;
assign v_45263 = v_45258 | v_45262;
assign v_45265 = v_45232 | v_45264;
assign v_45267 = v_45230 | v_45266;
assign v_45269 = v_45264 | v_45268;
assign v_45271 = v_45229 | v_45270;
assign v_45273 = v_45227 | v_45272;
assign v_45275 = v_45270 | v_45274;
assign v_45277 = v_45226 | v_45276;
assign v_45279 = v_45224 | v_45278;
assign v_45281 = v_45276 | v_45280;
assign v_45283 = v_45223 | v_45282;
assign v_45285 = v_45221 | v_45284;
assign v_45287 = v_45282 | v_45286;
assign v_45289 = v_45220 | v_45288;
assign v_45291 = v_45218 | v_45290;
assign v_45293 = v_45288 | v_45292;
assign v_45295 = v_45217 | v_45294;
assign v_45297 = v_45215 | v_45296;
assign v_45299 = v_45294 | v_45298;
assign v_45301 = v_45214 | v_45300;
assign v_45303 = v_45212 | v_45302;
assign v_45305 = v_45300 | v_45304;
assign v_45307 = v_45211 | v_45306;
assign v_45309 = v_45209 | v_45308;
assign v_45311 = v_45306 | v_45310;
assign v_45313 = v_45208 | v_45312;
assign v_45315 = v_45206 | v_45314;
assign v_45317 = v_45312 | v_45316;
assign v_45319 = v_45205 | v_45318;
assign v_45321 = v_45203 | v_45320;
assign v_45323 = v_45318 | v_45322;
assign v_45325 = v_45202 | v_45324;
assign v_45327 = v_45200 | v_45326;
assign v_45329 = v_45324 | v_45328;
assign v_45331 = v_45199 | v_45330;
assign v_45333 = v_45197 | v_45332;
assign v_45335 = v_45330 | v_45334;
assign v_45337 = v_45196 | v_45336;
assign v_45339 = v_45194 | v_45338;
assign v_45341 = v_45336 | v_45340;
assign v_45344 = ~v_45193 | v_45343;
assign v_45351 = v_45241 | v_45350;
assign v_45354 = v_45352 | v_45353;
assign v_45356 = v_45238 | v_45355;
assign v_45359 = v_45357 | v_45358;
assign v_45361 = v_45235 | v_45360;
assign v_45364 = v_45362 | v_45363;
assign v_45366 = v_45232 | v_45365;
assign v_45369 = v_45367 | v_45368;
assign v_45371 = v_45229 | v_45370;
assign v_45374 = v_45372 | v_45373;
assign v_45376 = v_45226 | v_45375;
assign v_45379 = v_45377 | v_45378;
assign v_45381 = v_45223 | v_45380;
assign v_45384 = v_45382 | v_45383;
assign v_45386 = v_45220 | v_45385;
assign v_45389 = v_45387 | v_45388;
assign v_45391 = v_45217 | v_45390;
assign v_45394 = v_45392 | v_45393;
assign v_45396 = v_45214 | v_45395;
assign v_45399 = v_45397 | v_45398;
assign v_45401 = v_45211 | v_45400;
assign v_45404 = v_45402 | v_45403;
assign v_45406 = v_45208 | v_45405;
assign v_45409 = v_45407 | v_45408;
assign v_45411 = v_45205 | v_45410;
assign v_45414 = v_45412 | v_45413;
assign v_45416 = v_45202 | v_45415;
assign v_45419 = v_45417 | v_45418;
assign v_45421 = v_45199 | v_45420;
assign v_45424 = v_45422 | v_45423;
assign v_45426 = v_45196 | v_45425;
assign v_45429 = v_45427 | v_45428;
assign v_45431 = v_45193 | v_45430;
assign v_45434 = v_45192 | v_45433;
assign v_45488 = v_45485 | v_45487;
assign v_45490 = v_45484 | v_45489;
assign v_45492 = v_45482 | v_45491;
assign v_45494 = v_45489 | v_45493;
assign v_45496 = v_45481 | v_45495;
assign v_45498 = v_45479 | v_45497;
assign v_45500 = v_45495 | v_45499;
assign v_45502 = v_45478 | v_45501;
assign v_45504 = v_45476 | v_45503;
assign v_45506 = v_45501 | v_45505;
assign v_45508 = v_45475 | v_45507;
assign v_45510 = v_45473 | v_45509;
assign v_45512 = v_45507 | v_45511;
assign v_45514 = v_45472 | v_45513;
assign v_45516 = v_45470 | v_45515;
assign v_45518 = v_45513 | v_45517;
assign v_45520 = v_45469 | v_45519;
assign v_45522 = v_45467 | v_45521;
assign v_45524 = v_45519 | v_45523;
assign v_45526 = v_45466 | v_45525;
assign v_45528 = v_45464 | v_45527;
assign v_45530 = v_45525 | v_45529;
assign v_45532 = v_45463 | v_45531;
assign v_45534 = v_45461 | v_45533;
assign v_45536 = v_45531 | v_45535;
assign v_45538 = v_45460 | v_45537;
assign v_45540 = v_45458 | v_45539;
assign v_45542 = v_45537 | v_45541;
assign v_45544 = v_45457 | v_45543;
assign v_45546 = v_45455 | v_45545;
assign v_45548 = v_45543 | v_45547;
assign v_45550 = v_45454 | v_45549;
assign v_45552 = v_45452 | v_45551;
assign v_45554 = v_45549 | v_45553;
assign v_45556 = v_45451 | v_45555;
assign v_45558 = v_45449 | v_45557;
assign v_45560 = v_45555 | v_45559;
assign v_45562 = v_45448 | v_45561;
assign v_45564 = v_45446 | v_45563;
assign v_45566 = v_45561 | v_45565;
assign v_45568 = v_45445 | v_45567;
assign v_45570 = v_45443 | v_45569;
assign v_45572 = v_45567 | v_45571;
assign v_45574 = v_45442 | v_45573;
assign v_45576 = v_45440 | v_45575;
assign v_45578 = v_45573 | v_45577;
assign v_45580 = v_45439 | v_45579;
assign v_45582 = v_45437 | v_45581;
assign v_45584 = v_45579 | v_45583;
assign v_45587 = ~v_45436 | v_45586;
assign v_45594 = v_45484 | v_45593;
assign v_45597 = v_45595 | v_45596;
assign v_45599 = v_45481 | v_45598;
assign v_45602 = v_45600 | v_45601;
assign v_45604 = v_45478 | v_45603;
assign v_45607 = v_45605 | v_45606;
assign v_45609 = v_45475 | v_45608;
assign v_45612 = v_45610 | v_45611;
assign v_45614 = v_45472 | v_45613;
assign v_45617 = v_45615 | v_45616;
assign v_45619 = v_45469 | v_45618;
assign v_45622 = v_45620 | v_45621;
assign v_45624 = v_45466 | v_45623;
assign v_45627 = v_45625 | v_45626;
assign v_45629 = v_45463 | v_45628;
assign v_45632 = v_45630 | v_45631;
assign v_45634 = v_45460 | v_45633;
assign v_45637 = v_45635 | v_45636;
assign v_45639 = v_45457 | v_45638;
assign v_45642 = v_45640 | v_45641;
assign v_45644 = v_45454 | v_45643;
assign v_45647 = v_45645 | v_45646;
assign v_45649 = v_45451 | v_45648;
assign v_45652 = v_45650 | v_45651;
assign v_45654 = v_45448 | v_45653;
assign v_45657 = v_45655 | v_45656;
assign v_45659 = v_45445 | v_45658;
assign v_45662 = v_45660 | v_45661;
assign v_45664 = v_45442 | v_45663;
assign v_45667 = v_45665 | v_45666;
assign v_45669 = v_45439 | v_45668;
assign v_45672 = v_45670 | v_45671;
assign v_45674 = v_45436 | v_45673;
assign v_45677 = v_45435 | v_45676;
assign v_45730 = v_45727 | v_45729;
assign v_45732 = v_45726 | v_45731;
assign v_45734 = v_45724 | v_45733;
assign v_45736 = v_45731 | v_45735;
assign v_45738 = v_45723 | v_45737;
assign v_45740 = v_45721 | v_45739;
assign v_45742 = v_45737 | v_45741;
assign v_45744 = v_45720 | v_45743;
assign v_45746 = v_45718 | v_45745;
assign v_45748 = v_45743 | v_45747;
assign v_45750 = v_45717 | v_45749;
assign v_45752 = v_45715 | v_45751;
assign v_45754 = v_45749 | v_45753;
assign v_45756 = v_45714 | v_45755;
assign v_45758 = v_45712 | v_45757;
assign v_45760 = v_45755 | v_45759;
assign v_45762 = v_45711 | v_45761;
assign v_45764 = v_45709 | v_45763;
assign v_45766 = v_45761 | v_45765;
assign v_45768 = v_45708 | v_45767;
assign v_45770 = v_45706 | v_45769;
assign v_45772 = v_45767 | v_45771;
assign v_45774 = v_45705 | v_45773;
assign v_45776 = v_45703 | v_45775;
assign v_45778 = v_45773 | v_45777;
assign v_45780 = v_45702 | v_45779;
assign v_45782 = v_45700 | v_45781;
assign v_45784 = v_45779 | v_45783;
assign v_45786 = v_45699 | v_45785;
assign v_45788 = v_45697 | v_45787;
assign v_45790 = v_45785 | v_45789;
assign v_45792 = v_45696 | v_45791;
assign v_45794 = v_45694 | v_45793;
assign v_45796 = v_45791 | v_45795;
assign v_45798 = v_45693 | v_45797;
assign v_45800 = v_45691 | v_45799;
assign v_45802 = v_45797 | v_45801;
assign v_45804 = v_45690 | v_45803;
assign v_45806 = v_45688 | v_45805;
assign v_45808 = v_45803 | v_45807;
assign v_45810 = v_45687 | v_45809;
assign v_45812 = v_45685 | v_45811;
assign v_45814 = v_45809 | v_45813;
assign v_45816 = v_45684 | v_45815;
assign v_45818 = v_45682 | v_45817;
assign v_45820 = v_45815 | v_45819;
assign v_45822 = v_45681 | v_45821;
assign v_45824 = v_45679 | v_45823;
assign v_45826 = v_45821 | v_45825;
assign v_45830 = v_45827 | v_45829;
assign v_45837 = v_45726 | v_45836;
assign v_45840 = v_45838 | v_45839;
assign v_45842 = v_45723 | v_45841;
assign v_45845 = v_45843 | v_45844;
assign v_45847 = v_45720 | v_45846;
assign v_45850 = v_45848 | v_45849;
assign v_45852 = v_45717 | v_45851;
assign v_45855 = v_45853 | v_45854;
assign v_45857 = v_45714 | v_45856;
assign v_45860 = v_45858 | v_45859;
assign v_45862 = v_45711 | v_45861;
assign v_45865 = v_45863 | v_45864;
assign v_45867 = v_45708 | v_45866;
assign v_45870 = v_45868 | v_45869;
assign v_45872 = v_45705 | v_45871;
assign v_45875 = v_45873 | v_45874;
assign v_45877 = v_45702 | v_45876;
assign v_45880 = v_45878 | v_45879;
assign v_45882 = v_45699 | v_45881;
assign v_45885 = v_45883 | v_45884;
assign v_45887 = v_45696 | v_45886;
assign v_45890 = v_45888 | v_45889;
assign v_45892 = v_45693 | v_45891;
assign v_45895 = v_45893 | v_45894;
assign v_45897 = v_45690 | v_45896;
assign v_45900 = v_45898 | v_45899;
assign v_45902 = v_45687 | v_45901;
assign v_45905 = v_45903 | v_45904;
assign v_45907 = v_45684 | v_45906;
assign v_45910 = v_45908 | v_45909;
assign v_45912 = v_45681 | v_45911;
assign v_45915 = v_45913 | v_45914;
assign v_45917 = v_45915 | v_45916;
assign v_45920 = v_45678 | v_45919;
assign v_45991 = v_45988 | v_45990;
assign v_45993 = v_45986 | v_45992;
assign v_45995 = v_45984 | v_45994;
assign v_45997 = v_45992 | v_45996;
assign v_45999 = v_45982 | v_45998;
assign v_46001 = v_45980 | v_46000;
assign v_46003 = v_45998 | v_46002;
assign v_46005 = v_45978 | v_46004;
assign v_46007 = v_45976 | v_46006;
assign v_46009 = v_46004 | v_46008;
assign v_46011 = v_45974 | v_46010;
assign v_46013 = v_45972 | v_46012;
assign v_46015 = v_46010 | v_46014;
assign v_46017 = v_45970 | v_46016;
assign v_46019 = v_45968 | v_46018;
assign v_46021 = v_46016 | v_46020;
assign v_46023 = v_45966 | v_46022;
assign v_46025 = v_45964 | v_46024;
assign v_46027 = v_46022 | v_46026;
assign v_46029 = v_45962 | v_46028;
assign v_46031 = v_45960 | v_46030;
assign v_46033 = v_46028 | v_46032;
assign v_46035 = v_45958 | v_46034;
assign v_46037 = v_45956 | v_46036;
assign v_46039 = v_46034 | v_46038;
assign v_46041 = v_45954 | v_46040;
assign v_46043 = v_45952 | v_46042;
assign v_46045 = v_46040 | v_46044;
assign v_46047 = v_45950 | v_46046;
assign v_46049 = v_45948 | v_46048;
assign v_46051 = v_46046 | v_46050;
assign v_46053 = v_45946 | v_46052;
assign v_46055 = v_45944 | v_46054;
assign v_46057 = v_46052 | v_46056;
assign v_46059 = v_45942 | v_46058;
assign v_46061 = v_45940 | v_46060;
assign v_46063 = v_46058 | v_46062;
assign v_46065 = v_45938 | v_46064;
assign v_46067 = v_45935 | v_46066;
assign v_46069 = v_46064 | v_46068;
assign v_46071 = v_45934 | v_46070;
assign v_46073 = v_45931 | v_46072;
assign v_46075 = v_46070 | v_46074;
assign v_46077 = v_45930 | v_46076;
assign v_46079 = v_45927 | v_46078;
assign v_46081 = v_46076 | v_46080;
assign v_46083 = v_45926 | v_46082;
assign v_46085 = v_45923 | v_46084;
assign v_46087 = v_46082 | v_46086;
assign v_46090 = ~v_45922 | v_46089;
assign v_46097 = v_45986 | v_46096;
assign v_46100 = v_46098 | v_46099;
assign v_46102 = v_45982 | v_46101;
assign v_46105 = v_46103 | v_46104;
assign v_46107 = v_45978 | v_46106;
assign v_46110 = v_46108 | v_46109;
assign v_46112 = v_45974 | v_46111;
assign v_46115 = v_46113 | v_46114;
assign v_46117 = v_45970 | v_46116;
assign v_46120 = v_46118 | v_46119;
assign v_46122 = v_45966 | v_46121;
assign v_46125 = v_46123 | v_46124;
assign v_46127 = v_45962 | v_46126;
assign v_46130 = v_46128 | v_46129;
assign v_46132 = v_45958 | v_46131;
assign v_46135 = v_46133 | v_46134;
assign v_46137 = v_45954 | v_46136;
assign v_46140 = v_46138 | v_46139;
assign v_46142 = v_45950 | v_46141;
assign v_46145 = v_46143 | v_46144;
assign v_46147 = v_45946 | v_46146;
assign v_46150 = v_46148 | v_46149;
assign v_46152 = v_45942 | v_46151;
assign v_46155 = v_46153 | v_46154;
assign v_46157 = v_45938 | v_46156;
assign v_46160 = v_46158 | v_46159;
assign v_46162 = v_45934 | v_46161;
assign v_46165 = v_46163 | v_46164;
assign v_46167 = v_45930 | v_46166;
assign v_46170 = v_46168 | v_46169;
assign v_46172 = v_45926 | v_46171;
assign v_46175 = v_46173 | v_46174;
assign v_46177 = v_45922 | v_46176;
assign v_46180 = v_45921 | v_46179;
assign v_46234 = v_46231 | v_46233;
assign v_46236 = v_46230 | v_46235;
assign v_46238 = v_46228 | v_46237;
assign v_46240 = v_46235 | v_46239;
assign v_46242 = v_46227 | v_46241;
assign v_46244 = v_46225 | v_46243;
assign v_46246 = v_46241 | v_46245;
assign v_46248 = v_46224 | v_46247;
assign v_46250 = v_46222 | v_46249;
assign v_46252 = v_46247 | v_46251;
assign v_46254 = v_46221 | v_46253;
assign v_46256 = v_46219 | v_46255;
assign v_46258 = v_46253 | v_46257;
assign v_46260 = v_46218 | v_46259;
assign v_46262 = v_46216 | v_46261;
assign v_46264 = v_46259 | v_46263;
assign v_46266 = v_46215 | v_46265;
assign v_46268 = v_46213 | v_46267;
assign v_46270 = v_46265 | v_46269;
assign v_46272 = v_46212 | v_46271;
assign v_46274 = v_46210 | v_46273;
assign v_46276 = v_46271 | v_46275;
assign v_46278 = v_46209 | v_46277;
assign v_46280 = v_46207 | v_46279;
assign v_46282 = v_46277 | v_46281;
assign v_46284 = v_46206 | v_46283;
assign v_46286 = v_46204 | v_46285;
assign v_46288 = v_46283 | v_46287;
assign v_46290 = v_46203 | v_46289;
assign v_46292 = v_46201 | v_46291;
assign v_46294 = v_46289 | v_46293;
assign v_46296 = v_46200 | v_46295;
assign v_46298 = v_46198 | v_46297;
assign v_46300 = v_46295 | v_46299;
assign v_46302 = v_46197 | v_46301;
assign v_46304 = v_46195 | v_46303;
assign v_46306 = v_46301 | v_46305;
assign v_46308 = v_46194 | v_46307;
assign v_46310 = v_46192 | v_46309;
assign v_46312 = v_46307 | v_46311;
assign v_46314 = v_46191 | v_46313;
assign v_46316 = v_46189 | v_46315;
assign v_46318 = v_46313 | v_46317;
assign v_46320 = v_46188 | v_46319;
assign v_46322 = v_46186 | v_46321;
assign v_46324 = v_46319 | v_46323;
assign v_46326 = v_46185 | v_46325;
assign v_46328 = v_46183 | v_46327;
assign v_46330 = v_46325 | v_46329;
assign v_46333 = ~v_46182 | v_46332;
assign v_46340 = v_46230 | v_46339;
assign v_46343 = v_46341 | v_46342;
assign v_46345 = v_46227 | v_46344;
assign v_46348 = v_46346 | v_46347;
assign v_46350 = v_46224 | v_46349;
assign v_46353 = v_46351 | v_46352;
assign v_46355 = v_46221 | v_46354;
assign v_46358 = v_46356 | v_46357;
assign v_46360 = v_46218 | v_46359;
assign v_46363 = v_46361 | v_46362;
assign v_46365 = v_46215 | v_46364;
assign v_46368 = v_46366 | v_46367;
assign v_46370 = v_46212 | v_46369;
assign v_46373 = v_46371 | v_46372;
assign v_46375 = v_46209 | v_46374;
assign v_46378 = v_46376 | v_46377;
assign v_46380 = v_46206 | v_46379;
assign v_46383 = v_46381 | v_46382;
assign v_46385 = v_46203 | v_46384;
assign v_46388 = v_46386 | v_46387;
assign v_46390 = v_46200 | v_46389;
assign v_46393 = v_46391 | v_46392;
assign v_46395 = v_46197 | v_46394;
assign v_46398 = v_46396 | v_46397;
assign v_46400 = v_46194 | v_46399;
assign v_46403 = v_46401 | v_46402;
assign v_46405 = v_46191 | v_46404;
assign v_46408 = v_46406 | v_46407;
assign v_46410 = v_46188 | v_46409;
assign v_46413 = v_46411 | v_46412;
assign v_46415 = v_46185 | v_46414;
assign v_46418 = v_46416 | v_46417;
assign v_46420 = v_46182 | v_46419;
assign v_46423 = v_46181 | v_46422;
assign v_46477 = v_46474 | v_46476;
assign v_46479 = v_46473 | v_46478;
assign v_46481 = v_46471 | v_46480;
assign v_46483 = v_46478 | v_46482;
assign v_46485 = v_46470 | v_46484;
assign v_46487 = v_46468 | v_46486;
assign v_46489 = v_46484 | v_46488;
assign v_46491 = v_46467 | v_46490;
assign v_46493 = v_46465 | v_46492;
assign v_46495 = v_46490 | v_46494;
assign v_46497 = v_46464 | v_46496;
assign v_46499 = v_46462 | v_46498;
assign v_46501 = v_46496 | v_46500;
assign v_46503 = v_46461 | v_46502;
assign v_46505 = v_46459 | v_46504;
assign v_46507 = v_46502 | v_46506;
assign v_46509 = v_46458 | v_46508;
assign v_46511 = v_46456 | v_46510;
assign v_46513 = v_46508 | v_46512;
assign v_46515 = v_46455 | v_46514;
assign v_46517 = v_46453 | v_46516;
assign v_46519 = v_46514 | v_46518;
assign v_46521 = v_46452 | v_46520;
assign v_46523 = v_46450 | v_46522;
assign v_46525 = v_46520 | v_46524;
assign v_46527 = v_46449 | v_46526;
assign v_46529 = v_46447 | v_46528;
assign v_46531 = v_46526 | v_46530;
assign v_46533 = v_46446 | v_46532;
assign v_46535 = v_46444 | v_46534;
assign v_46537 = v_46532 | v_46536;
assign v_46539 = v_46443 | v_46538;
assign v_46541 = v_46441 | v_46540;
assign v_46543 = v_46538 | v_46542;
assign v_46545 = v_46440 | v_46544;
assign v_46547 = v_46438 | v_46546;
assign v_46549 = v_46544 | v_46548;
assign v_46551 = v_46437 | v_46550;
assign v_46553 = v_46435 | v_46552;
assign v_46555 = v_46550 | v_46554;
assign v_46557 = v_46434 | v_46556;
assign v_46559 = v_46432 | v_46558;
assign v_46561 = v_46556 | v_46560;
assign v_46563 = v_46431 | v_46562;
assign v_46565 = v_46429 | v_46564;
assign v_46567 = v_46562 | v_46566;
assign v_46569 = v_46428 | v_46568;
assign v_46571 = v_46426 | v_46570;
assign v_46573 = v_46568 | v_46572;
assign v_46576 = ~v_46425 | v_46575;
assign v_46583 = v_46473 | v_46582;
assign v_46586 = v_46584 | v_46585;
assign v_46588 = v_46470 | v_46587;
assign v_46591 = v_46589 | v_46590;
assign v_46593 = v_46467 | v_46592;
assign v_46596 = v_46594 | v_46595;
assign v_46598 = v_46464 | v_46597;
assign v_46601 = v_46599 | v_46600;
assign v_46603 = v_46461 | v_46602;
assign v_46606 = v_46604 | v_46605;
assign v_46608 = v_46458 | v_46607;
assign v_46611 = v_46609 | v_46610;
assign v_46613 = v_46455 | v_46612;
assign v_46616 = v_46614 | v_46615;
assign v_46618 = v_46452 | v_46617;
assign v_46621 = v_46619 | v_46620;
assign v_46623 = v_46449 | v_46622;
assign v_46626 = v_46624 | v_46625;
assign v_46628 = v_46446 | v_46627;
assign v_46631 = v_46629 | v_46630;
assign v_46633 = v_46443 | v_46632;
assign v_46636 = v_46634 | v_46635;
assign v_46638 = v_46440 | v_46637;
assign v_46641 = v_46639 | v_46640;
assign v_46643 = v_46437 | v_46642;
assign v_46646 = v_46644 | v_46645;
assign v_46648 = v_46434 | v_46647;
assign v_46651 = v_46649 | v_46650;
assign v_46653 = v_46431 | v_46652;
assign v_46656 = v_46654 | v_46655;
assign v_46658 = v_46428 | v_46657;
assign v_46661 = v_46659 | v_46660;
assign v_46663 = v_46425 | v_46662;
assign v_46666 = v_46424 | v_46665;
assign v_46720 = v_46717 | v_46719;
assign v_46722 = v_46716 | v_46721;
assign v_46724 = v_46714 | v_46723;
assign v_46726 = v_46721 | v_46725;
assign v_46728 = v_46713 | v_46727;
assign v_46730 = v_46711 | v_46729;
assign v_46732 = v_46727 | v_46731;
assign v_46734 = v_46710 | v_46733;
assign v_46736 = v_46708 | v_46735;
assign v_46738 = v_46733 | v_46737;
assign v_46740 = v_46707 | v_46739;
assign v_46742 = v_46705 | v_46741;
assign v_46744 = v_46739 | v_46743;
assign v_46746 = v_46704 | v_46745;
assign v_46748 = v_46702 | v_46747;
assign v_46750 = v_46745 | v_46749;
assign v_46752 = v_46701 | v_46751;
assign v_46754 = v_46699 | v_46753;
assign v_46756 = v_46751 | v_46755;
assign v_46758 = v_46698 | v_46757;
assign v_46760 = v_46696 | v_46759;
assign v_46762 = v_46757 | v_46761;
assign v_46764 = v_46695 | v_46763;
assign v_46766 = v_46693 | v_46765;
assign v_46768 = v_46763 | v_46767;
assign v_46770 = v_46692 | v_46769;
assign v_46772 = v_46690 | v_46771;
assign v_46774 = v_46769 | v_46773;
assign v_46776 = v_46689 | v_46775;
assign v_46778 = v_46687 | v_46777;
assign v_46780 = v_46775 | v_46779;
assign v_46782 = v_46686 | v_46781;
assign v_46784 = v_46684 | v_46783;
assign v_46786 = v_46781 | v_46785;
assign v_46788 = v_46683 | v_46787;
assign v_46790 = v_46681 | v_46789;
assign v_46792 = v_46787 | v_46791;
assign v_46794 = v_46680 | v_46793;
assign v_46796 = v_46678 | v_46795;
assign v_46798 = v_46793 | v_46797;
assign v_46800 = v_46677 | v_46799;
assign v_46802 = v_46675 | v_46801;
assign v_46804 = v_46799 | v_46803;
assign v_46806 = v_46674 | v_46805;
assign v_46808 = v_46672 | v_46807;
assign v_46810 = v_46805 | v_46809;
assign v_46812 = v_46671 | v_46811;
assign v_46814 = v_46669 | v_46813;
assign v_46816 = v_46811 | v_46815;
assign v_46819 = ~v_46668 | v_46818;
assign v_46826 = v_46716 | v_46825;
assign v_46829 = v_46827 | v_46828;
assign v_46831 = v_46713 | v_46830;
assign v_46834 = v_46832 | v_46833;
assign v_46836 = v_46710 | v_46835;
assign v_46839 = v_46837 | v_46838;
assign v_46841 = v_46707 | v_46840;
assign v_46844 = v_46842 | v_46843;
assign v_46846 = v_46704 | v_46845;
assign v_46849 = v_46847 | v_46848;
assign v_46851 = v_46701 | v_46850;
assign v_46854 = v_46852 | v_46853;
assign v_46856 = v_46698 | v_46855;
assign v_46859 = v_46857 | v_46858;
assign v_46861 = v_46695 | v_46860;
assign v_46864 = v_46862 | v_46863;
assign v_46866 = v_46692 | v_46865;
assign v_46869 = v_46867 | v_46868;
assign v_46871 = v_46689 | v_46870;
assign v_46874 = v_46872 | v_46873;
assign v_46876 = v_46686 | v_46875;
assign v_46879 = v_46877 | v_46878;
assign v_46881 = v_46683 | v_46880;
assign v_46884 = v_46882 | v_46883;
assign v_46886 = v_46680 | v_46885;
assign v_46889 = v_46887 | v_46888;
assign v_46891 = v_46677 | v_46890;
assign v_46894 = v_46892 | v_46893;
assign v_46896 = v_46674 | v_46895;
assign v_46899 = v_46897 | v_46898;
assign v_46901 = v_46671 | v_46900;
assign v_46904 = v_46902 | v_46903;
assign v_46906 = v_46668 | v_46905;
assign v_46909 = v_46667 | v_46908;
assign v_46963 = v_46960 | v_46962;
assign v_46965 = v_46959 | v_46964;
assign v_46967 = v_46957 | v_46966;
assign v_46969 = v_46964 | v_46968;
assign v_46971 = v_46956 | v_46970;
assign v_46973 = v_46954 | v_46972;
assign v_46975 = v_46970 | v_46974;
assign v_46977 = v_46953 | v_46976;
assign v_46979 = v_46951 | v_46978;
assign v_46981 = v_46976 | v_46980;
assign v_46983 = v_46950 | v_46982;
assign v_46985 = v_46948 | v_46984;
assign v_46987 = v_46982 | v_46986;
assign v_46989 = v_46947 | v_46988;
assign v_46991 = v_46945 | v_46990;
assign v_46993 = v_46988 | v_46992;
assign v_46995 = v_46944 | v_46994;
assign v_46997 = v_46942 | v_46996;
assign v_46999 = v_46994 | v_46998;
assign v_47001 = v_46941 | v_47000;
assign v_47003 = v_46939 | v_47002;
assign v_47005 = v_47000 | v_47004;
assign v_47007 = v_46938 | v_47006;
assign v_47009 = v_46936 | v_47008;
assign v_47011 = v_47006 | v_47010;
assign v_47013 = v_46935 | v_47012;
assign v_47015 = v_46933 | v_47014;
assign v_47017 = v_47012 | v_47016;
assign v_47019 = v_46932 | v_47018;
assign v_47021 = v_46930 | v_47020;
assign v_47023 = v_47018 | v_47022;
assign v_47025 = v_46929 | v_47024;
assign v_47027 = v_46927 | v_47026;
assign v_47029 = v_47024 | v_47028;
assign v_47031 = v_46926 | v_47030;
assign v_47033 = v_46924 | v_47032;
assign v_47035 = v_47030 | v_47034;
assign v_47037 = v_46923 | v_47036;
assign v_47039 = v_46921 | v_47038;
assign v_47041 = v_47036 | v_47040;
assign v_47043 = v_46920 | v_47042;
assign v_47045 = v_46918 | v_47044;
assign v_47047 = v_47042 | v_47046;
assign v_47049 = v_46917 | v_47048;
assign v_47051 = v_46915 | v_47050;
assign v_47053 = v_47048 | v_47052;
assign v_47055 = v_46914 | v_47054;
assign v_47057 = v_46912 | v_47056;
assign v_47059 = v_47054 | v_47058;
assign v_47062 = ~v_46911 | v_47061;
assign v_47069 = v_46959 | v_47068;
assign v_47072 = v_47070 | v_47071;
assign v_47074 = v_46956 | v_47073;
assign v_47077 = v_47075 | v_47076;
assign v_47079 = v_46953 | v_47078;
assign v_47082 = v_47080 | v_47081;
assign v_47084 = v_46950 | v_47083;
assign v_47087 = v_47085 | v_47086;
assign v_47089 = v_46947 | v_47088;
assign v_47092 = v_47090 | v_47091;
assign v_47094 = v_46944 | v_47093;
assign v_47097 = v_47095 | v_47096;
assign v_47099 = v_46941 | v_47098;
assign v_47102 = v_47100 | v_47101;
assign v_47104 = v_46938 | v_47103;
assign v_47107 = v_47105 | v_47106;
assign v_47109 = v_46935 | v_47108;
assign v_47112 = v_47110 | v_47111;
assign v_47114 = v_46932 | v_47113;
assign v_47117 = v_47115 | v_47116;
assign v_47119 = v_46929 | v_47118;
assign v_47122 = v_47120 | v_47121;
assign v_47124 = v_46926 | v_47123;
assign v_47127 = v_47125 | v_47126;
assign v_47129 = v_46923 | v_47128;
assign v_47132 = v_47130 | v_47131;
assign v_47134 = v_46920 | v_47133;
assign v_47137 = v_47135 | v_47136;
assign v_47139 = v_46917 | v_47138;
assign v_47142 = v_47140 | v_47141;
assign v_47144 = v_46914 | v_47143;
assign v_47147 = v_47145 | v_47146;
assign v_47149 = v_46911 | v_47148;
assign v_47152 = v_46910 | v_47151;
assign v_47206 = v_47203 | v_47205;
assign v_47208 = v_47202 | v_47207;
assign v_47210 = v_47200 | v_47209;
assign v_47212 = v_47207 | v_47211;
assign v_47214 = v_47199 | v_47213;
assign v_47216 = v_47197 | v_47215;
assign v_47218 = v_47213 | v_47217;
assign v_47220 = v_47196 | v_47219;
assign v_47222 = v_47194 | v_47221;
assign v_47224 = v_47219 | v_47223;
assign v_47226 = v_47193 | v_47225;
assign v_47228 = v_47191 | v_47227;
assign v_47230 = v_47225 | v_47229;
assign v_47232 = v_47190 | v_47231;
assign v_47234 = v_47188 | v_47233;
assign v_47236 = v_47231 | v_47235;
assign v_47238 = v_47187 | v_47237;
assign v_47240 = v_47185 | v_47239;
assign v_47242 = v_47237 | v_47241;
assign v_47244 = v_47184 | v_47243;
assign v_47246 = v_47182 | v_47245;
assign v_47248 = v_47243 | v_47247;
assign v_47250 = v_47181 | v_47249;
assign v_47252 = v_47179 | v_47251;
assign v_47254 = v_47249 | v_47253;
assign v_47256 = v_47178 | v_47255;
assign v_47258 = v_47176 | v_47257;
assign v_47260 = v_47255 | v_47259;
assign v_47262 = v_47175 | v_47261;
assign v_47264 = v_47173 | v_47263;
assign v_47266 = v_47261 | v_47265;
assign v_47268 = v_47172 | v_47267;
assign v_47270 = v_47170 | v_47269;
assign v_47272 = v_47267 | v_47271;
assign v_47274 = v_47169 | v_47273;
assign v_47276 = v_47167 | v_47275;
assign v_47278 = v_47273 | v_47277;
assign v_47280 = v_47166 | v_47279;
assign v_47282 = v_47164 | v_47281;
assign v_47284 = v_47279 | v_47283;
assign v_47286 = v_47163 | v_47285;
assign v_47288 = v_47161 | v_47287;
assign v_47290 = v_47285 | v_47289;
assign v_47292 = v_47160 | v_47291;
assign v_47294 = v_47158 | v_47293;
assign v_47296 = v_47291 | v_47295;
assign v_47298 = v_47157 | v_47297;
assign v_47300 = v_47155 | v_47299;
assign v_47302 = v_47297 | v_47301;
assign v_47305 = ~v_47154 | v_47304;
assign v_47312 = v_47202 | v_47311;
assign v_47315 = v_47313 | v_47314;
assign v_47317 = v_47199 | v_47316;
assign v_47320 = v_47318 | v_47319;
assign v_47322 = v_47196 | v_47321;
assign v_47325 = v_47323 | v_47324;
assign v_47327 = v_47193 | v_47326;
assign v_47330 = v_47328 | v_47329;
assign v_47332 = v_47190 | v_47331;
assign v_47335 = v_47333 | v_47334;
assign v_47337 = v_47187 | v_47336;
assign v_47340 = v_47338 | v_47339;
assign v_47342 = v_47184 | v_47341;
assign v_47345 = v_47343 | v_47344;
assign v_47347 = v_47181 | v_47346;
assign v_47350 = v_47348 | v_47349;
assign v_47352 = v_47178 | v_47351;
assign v_47355 = v_47353 | v_47354;
assign v_47357 = v_47175 | v_47356;
assign v_47360 = v_47358 | v_47359;
assign v_47362 = v_47172 | v_47361;
assign v_47365 = v_47363 | v_47364;
assign v_47367 = v_47169 | v_47366;
assign v_47370 = v_47368 | v_47369;
assign v_47372 = v_47166 | v_47371;
assign v_47375 = v_47373 | v_47374;
assign v_47377 = v_47163 | v_47376;
assign v_47380 = v_47378 | v_47379;
assign v_47382 = v_47160 | v_47381;
assign v_47385 = v_47383 | v_47384;
assign v_47387 = v_47157 | v_47386;
assign v_47390 = v_47388 | v_47389;
assign v_47392 = v_47154 | v_47391;
assign v_47395 = v_47153 | v_47394;
assign v_47449 = v_47446 | v_47448;
assign v_47451 = v_47445 | v_47450;
assign v_47453 = v_47443 | v_47452;
assign v_47455 = v_47450 | v_47454;
assign v_47457 = v_47442 | v_47456;
assign v_47459 = v_47440 | v_47458;
assign v_47461 = v_47456 | v_47460;
assign v_47463 = v_47439 | v_47462;
assign v_47465 = v_47437 | v_47464;
assign v_47467 = v_47462 | v_47466;
assign v_47469 = v_47436 | v_47468;
assign v_47471 = v_47434 | v_47470;
assign v_47473 = v_47468 | v_47472;
assign v_47475 = v_47433 | v_47474;
assign v_47477 = v_47431 | v_47476;
assign v_47479 = v_47474 | v_47478;
assign v_47481 = v_47430 | v_47480;
assign v_47483 = v_47428 | v_47482;
assign v_47485 = v_47480 | v_47484;
assign v_47487 = v_47427 | v_47486;
assign v_47489 = v_47425 | v_47488;
assign v_47491 = v_47486 | v_47490;
assign v_47493 = v_47424 | v_47492;
assign v_47495 = v_47422 | v_47494;
assign v_47497 = v_47492 | v_47496;
assign v_47499 = v_47421 | v_47498;
assign v_47501 = v_47419 | v_47500;
assign v_47503 = v_47498 | v_47502;
assign v_47505 = v_47418 | v_47504;
assign v_47507 = v_47416 | v_47506;
assign v_47509 = v_47504 | v_47508;
assign v_47511 = v_47415 | v_47510;
assign v_47513 = v_47413 | v_47512;
assign v_47515 = v_47510 | v_47514;
assign v_47517 = v_47412 | v_47516;
assign v_47519 = v_47410 | v_47518;
assign v_47521 = v_47516 | v_47520;
assign v_47523 = v_47409 | v_47522;
assign v_47525 = v_47407 | v_47524;
assign v_47527 = v_47522 | v_47526;
assign v_47529 = v_47406 | v_47528;
assign v_47531 = v_47404 | v_47530;
assign v_47533 = v_47528 | v_47532;
assign v_47535 = v_47403 | v_47534;
assign v_47537 = v_47401 | v_47536;
assign v_47539 = v_47534 | v_47538;
assign v_47541 = v_47400 | v_47540;
assign v_47543 = v_47398 | v_47542;
assign v_47545 = v_47540 | v_47544;
assign v_47548 = ~v_47397 | v_47547;
assign v_47555 = v_47445 | v_47554;
assign v_47558 = v_47556 | v_47557;
assign v_47560 = v_47442 | v_47559;
assign v_47563 = v_47561 | v_47562;
assign v_47565 = v_47439 | v_47564;
assign v_47568 = v_47566 | v_47567;
assign v_47570 = v_47436 | v_47569;
assign v_47573 = v_47571 | v_47572;
assign v_47575 = v_47433 | v_47574;
assign v_47578 = v_47576 | v_47577;
assign v_47580 = v_47430 | v_47579;
assign v_47583 = v_47581 | v_47582;
assign v_47585 = v_47427 | v_47584;
assign v_47588 = v_47586 | v_47587;
assign v_47590 = v_47424 | v_47589;
assign v_47593 = v_47591 | v_47592;
assign v_47595 = v_47421 | v_47594;
assign v_47598 = v_47596 | v_47597;
assign v_47600 = v_47418 | v_47599;
assign v_47603 = v_47601 | v_47602;
assign v_47605 = v_47415 | v_47604;
assign v_47608 = v_47606 | v_47607;
assign v_47610 = v_47412 | v_47609;
assign v_47613 = v_47611 | v_47612;
assign v_47615 = v_47409 | v_47614;
assign v_47618 = v_47616 | v_47617;
assign v_47620 = v_47406 | v_47619;
assign v_47623 = v_47621 | v_47622;
assign v_47625 = v_47403 | v_47624;
assign v_47628 = v_47626 | v_47627;
assign v_47630 = v_47400 | v_47629;
assign v_47633 = v_47631 | v_47632;
assign v_47635 = v_47397 | v_47634;
assign v_47638 = v_47396 | v_47637;
assign v_47692 = v_47689 | v_47691;
assign v_47694 = v_47688 | v_47693;
assign v_47696 = v_47686 | v_47695;
assign v_47698 = v_47693 | v_47697;
assign v_47700 = v_47685 | v_47699;
assign v_47702 = v_47683 | v_47701;
assign v_47704 = v_47699 | v_47703;
assign v_47706 = v_47682 | v_47705;
assign v_47708 = v_47680 | v_47707;
assign v_47710 = v_47705 | v_47709;
assign v_47712 = v_47679 | v_47711;
assign v_47714 = v_47677 | v_47713;
assign v_47716 = v_47711 | v_47715;
assign v_47718 = v_47676 | v_47717;
assign v_47720 = v_47674 | v_47719;
assign v_47722 = v_47717 | v_47721;
assign v_47724 = v_47673 | v_47723;
assign v_47726 = v_47671 | v_47725;
assign v_47728 = v_47723 | v_47727;
assign v_47730 = v_47670 | v_47729;
assign v_47732 = v_47668 | v_47731;
assign v_47734 = v_47729 | v_47733;
assign v_47736 = v_47667 | v_47735;
assign v_47738 = v_47665 | v_47737;
assign v_47740 = v_47735 | v_47739;
assign v_47742 = v_47664 | v_47741;
assign v_47744 = v_47662 | v_47743;
assign v_47746 = v_47741 | v_47745;
assign v_47748 = v_47661 | v_47747;
assign v_47750 = v_47659 | v_47749;
assign v_47752 = v_47747 | v_47751;
assign v_47754 = v_47658 | v_47753;
assign v_47756 = v_47656 | v_47755;
assign v_47758 = v_47753 | v_47757;
assign v_47760 = v_47655 | v_47759;
assign v_47762 = v_47653 | v_47761;
assign v_47764 = v_47759 | v_47763;
assign v_47766 = v_47652 | v_47765;
assign v_47768 = v_47650 | v_47767;
assign v_47770 = v_47765 | v_47769;
assign v_47772 = v_47649 | v_47771;
assign v_47774 = v_47647 | v_47773;
assign v_47776 = v_47771 | v_47775;
assign v_47778 = v_47646 | v_47777;
assign v_47780 = v_47644 | v_47779;
assign v_47782 = v_47777 | v_47781;
assign v_47784 = v_47643 | v_47783;
assign v_47786 = v_47641 | v_47785;
assign v_47788 = v_47783 | v_47787;
assign v_47791 = ~v_47640 | v_47790;
assign v_47798 = v_47688 | v_47797;
assign v_47801 = v_47799 | v_47800;
assign v_47803 = v_47685 | v_47802;
assign v_47806 = v_47804 | v_47805;
assign v_47808 = v_47682 | v_47807;
assign v_47811 = v_47809 | v_47810;
assign v_47813 = v_47679 | v_47812;
assign v_47816 = v_47814 | v_47815;
assign v_47818 = v_47676 | v_47817;
assign v_47821 = v_47819 | v_47820;
assign v_47823 = v_47673 | v_47822;
assign v_47826 = v_47824 | v_47825;
assign v_47828 = v_47670 | v_47827;
assign v_47831 = v_47829 | v_47830;
assign v_47833 = v_47667 | v_47832;
assign v_47836 = v_47834 | v_47835;
assign v_47838 = v_47664 | v_47837;
assign v_47841 = v_47839 | v_47840;
assign v_47843 = v_47661 | v_47842;
assign v_47846 = v_47844 | v_47845;
assign v_47848 = v_47658 | v_47847;
assign v_47851 = v_47849 | v_47850;
assign v_47853 = v_47655 | v_47852;
assign v_47856 = v_47854 | v_47855;
assign v_47858 = v_47652 | v_47857;
assign v_47861 = v_47859 | v_47860;
assign v_47863 = v_47649 | v_47862;
assign v_47866 = v_47864 | v_47865;
assign v_47868 = v_47646 | v_47867;
assign v_47871 = v_47869 | v_47870;
assign v_47873 = v_47643 | v_47872;
assign v_47876 = v_47874 | v_47875;
assign v_47878 = v_47640 | v_47877;
assign v_47881 = v_47639 | v_47880;
assign v_47935 = v_47932 | v_47934;
assign v_47937 = v_47931 | v_47936;
assign v_47939 = v_47929 | v_47938;
assign v_47941 = v_47936 | v_47940;
assign v_47943 = v_47928 | v_47942;
assign v_47945 = v_47926 | v_47944;
assign v_47947 = v_47942 | v_47946;
assign v_47949 = v_47925 | v_47948;
assign v_47951 = v_47923 | v_47950;
assign v_47953 = v_47948 | v_47952;
assign v_47955 = v_47922 | v_47954;
assign v_47957 = v_47920 | v_47956;
assign v_47959 = v_47954 | v_47958;
assign v_47961 = v_47919 | v_47960;
assign v_47963 = v_47917 | v_47962;
assign v_47965 = v_47960 | v_47964;
assign v_47967 = v_47916 | v_47966;
assign v_47969 = v_47914 | v_47968;
assign v_47971 = v_47966 | v_47970;
assign v_47973 = v_47913 | v_47972;
assign v_47975 = v_47911 | v_47974;
assign v_47977 = v_47972 | v_47976;
assign v_47979 = v_47910 | v_47978;
assign v_47981 = v_47908 | v_47980;
assign v_47983 = v_47978 | v_47982;
assign v_47985 = v_47907 | v_47984;
assign v_47987 = v_47905 | v_47986;
assign v_47989 = v_47984 | v_47988;
assign v_47991 = v_47904 | v_47990;
assign v_47993 = v_47902 | v_47992;
assign v_47995 = v_47990 | v_47994;
assign v_47997 = v_47901 | v_47996;
assign v_47999 = v_47899 | v_47998;
assign v_48001 = v_47996 | v_48000;
assign v_48003 = v_47898 | v_48002;
assign v_48005 = v_47896 | v_48004;
assign v_48007 = v_48002 | v_48006;
assign v_48009 = v_47895 | v_48008;
assign v_48011 = v_47893 | v_48010;
assign v_48013 = v_48008 | v_48012;
assign v_48015 = v_47892 | v_48014;
assign v_48017 = v_47890 | v_48016;
assign v_48019 = v_48014 | v_48018;
assign v_48021 = v_47889 | v_48020;
assign v_48023 = v_47887 | v_48022;
assign v_48025 = v_48020 | v_48024;
assign v_48027 = v_47886 | v_48026;
assign v_48029 = v_47884 | v_48028;
assign v_48031 = v_48026 | v_48030;
assign v_48034 = ~v_47883 | v_48033;
assign v_48041 = v_47931 | v_48040;
assign v_48044 = v_48042 | v_48043;
assign v_48046 = v_47928 | v_48045;
assign v_48049 = v_48047 | v_48048;
assign v_48051 = v_47925 | v_48050;
assign v_48054 = v_48052 | v_48053;
assign v_48056 = v_47922 | v_48055;
assign v_48059 = v_48057 | v_48058;
assign v_48061 = v_47919 | v_48060;
assign v_48064 = v_48062 | v_48063;
assign v_48066 = v_47916 | v_48065;
assign v_48069 = v_48067 | v_48068;
assign v_48071 = v_47913 | v_48070;
assign v_48074 = v_48072 | v_48073;
assign v_48076 = v_47910 | v_48075;
assign v_48079 = v_48077 | v_48078;
assign v_48081 = v_47907 | v_48080;
assign v_48084 = v_48082 | v_48083;
assign v_48086 = v_47904 | v_48085;
assign v_48089 = v_48087 | v_48088;
assign v_48091 = v_47901 | v_48090;
assign v_48094 = v_48092 | v_48093;
assign v_48096 = v_47898 | v_48095;
assign v_48099 = v_48097 | v_48098;
assign v_48101 = v_47895 | v_48100;
assign v_48104 = v_48102 | v_48103;
assign v_48106 = v_47892 | v_48105;
assign v_48109 = v_48107 | v_48108;
assign v_48111 = v_47889 | v_48110;
assign v_48114 = v_48112 | v_48113;
assign v_48116 = v_47886 | v_48115;
assign v_48119 = v_48117 | v_48118;
assign v_48121 = v_47883 | v_48120;
assign v_48124 = v_47882 | v_48123;
assign v_48178 = v_48175 | v_48177;
assign v_48180 = v_48174 | v_48179;
assign v_48182 = v_48172 | v_48181;
assign v_48184 = v_48179 | v_48183;
assign v_48186 = v_48171 | v_48185;
assign v_48188 = v_48169 | v_48187;
assign v_48190 = v_48185 | v_48189;
assign v_48192 = v_48168 | v_48191;
assign v_48194 = v_48166 | v_48193;
assign v_48196 = v_48191 | v_48195;
assign v_48198 = v_48165 | v_48197;
assign v_48200 = v_48163 | v_48199;
assign v_48202 = v_48197 | v_48201;
assign v_48204 = v_48162 | v_48203;
assign v_48206 = v_48160 | v_48205;
assign v_48208 = v_48203 | v_48207;
assign v_48210 = v_48159 | v_48209;
assign v_48212 = v_48157 | v_48211;
assign v_48214 = v_48209 | v_48213;
assign v_48216 = v_48156 | v_48215;
assign v_48218 = v_48154 | v_48217;
assign v_48220 = v_48215 | v_48219;
assign v_48222 = v_48153 | v_48221;
assign v_48224 = v_48151 | v_48223;
assign v_48226 = v_48221 | v_48225;
assign v_48228 = v_48150 | v_48227;
assign v_48230 = v_48148 | v_48229;
assign v_48232 = v_48227 | v_48231;
assign v_48234 = v_48147 | v_48233;
assign v_48236 = v_48145 | v_48235;
assign v_48238 = v_48233 | v_48237;
assign v_48240 = v_48144 | v_48239;
assign v_48242 = v_48142 | v_48241;
assign v_48244 = v_48239 | v_48243;
assign v_48246 = v_48141 | v_48245;
assign v_48248 = v_48139 | v_48247;
assign v_48250 = v_48245 | v_48249;
assign v_48252 = v_48138 | v_48251;
assign v_48254 = v_48136 | v_48253;
assign v_48256 = v_48251 | v_48255;
assign v_48258 = v_48135 | v_48257;
assign v_48260 = v_48133 | v_48259;
assign v_48262 = v_48257 | v_48261;
assign v_48264 = v_48132 | v_48263;
assign v_48266 = v_48130 | v_48265;
assign v_48268 = v_48263 | v_48267;
assign v_48270 = v_48129 | v_48269;
assign v_48272 = v_48127 | v_48271;
assign v_48274 = v_48269 | v_48273;
assign v_48277 = ~v_48126 | v_48276;
assign v_48284 = v_48174 | v_48283;
assign v_48287 = v_48285 | v_48286;
assign v_48289 = v_48171 | v_48288;
assign v_48292 = v_48290 | v_48291;
assign v_48294 = v_48168 | v_48293;
assign v_48297 = v_48295 | v_48296;
assign v_48299 = v_48165 | v_48298;
assign v_48302 = v_48300 | v_48301;
assign v_48304 = v_48162 | v_48303;
assign v_48307 = v_48305 | v_48306;
assign v_48309 = v_48159 | v_48308;
assign v_48312 = v_48310 | v_48311;
assign v_48314 = v_48156 | v_48313;
assign v_48317 = v_48315 | v_48316;
assign v_48319 = v_48153 | v_48318;
assign v_48322 = v_48320 | v_48321;
assign v_48324 = v_48150 | v_48323;
assign v_48327 = v_48325 | v_48326;
assign v_48329 = v_48147 | v_48328;
assign v_48332 = v_48330 | v_48331;
assign v_48334 = v_48144 | v_48333;
assign v_48337 = v_48335 | v_48336;
assign v_48339 = v_48141 | v_48338;
assign v_48342 = v_48340 | v_48341;
assign v_48344 = v_48138 | v_48343;
assign v_48347 = v_48345 | v_48346;
assign v_48349 = v_48135 | v_48348;
assign v_48352 = v_48350 | v_48351;
assign v_48354 = v_48132 | v_48353;
assign v_48357 = v_48355 | v_48356;
assign v_48359 = v_48129 | v_48358;
assign v_48362 = v_48360 | v_48361;
assign v_48364 = v_48126 | v_48363;
assign v_48367 = v_48125 | v_48366;
assign v_48421 = v_48418 | v_48420;
assign v_48423 = v_48417 | v_48422;
assign v_48425 = v_48415 | v_48424;
assign v_48427 = v_48422 | v_48426;
assign v_48429 = v_48414 | v_48428;
assign v_48431 = v_48412 | v_48430;
assign v_48433 = v_48428 | v_48432;
assign v_48435 = v_48411 | v_48434;
assign v_48437 = v_48409 | v_48436;
assign v_48439 = v_48434 | v_48438;
assign v_48441 = v_48408 | v_48440;
assign v_48443 = v_48406 | v_48442;
assign v_48445 = v_48440 | v_48444;
assign v_48447 = v_48405 | v_48446;
assign v_48449 = v_48403 | v_48448;
assign v_48451 = v_48446 | v_48450;
assign v_48453 = v_48402 | v_48452;
assign v_48455 = v_48400 | v_48454;
assign v_48457 = v_48452 | v_48456;
assign v_48459 = v_48399 | v_48458;
assign v_48461 = v_48397 | v_48460;
assign v_48463 = v_48458 | v_48462;
assign v_48465 = v_48396 | v_48464;
assign v_48467 = v_48394 | v_48466;
assign v_48469 = v_48464 | v_48468;
assign v_48471 = v_48393 | v_48470;
assign v_48473 = v_48391 | v_48472;
assign v_48475 = v_48470 | v_48474;
assign v_48477 = v_48390 | v_48476;
assign v_48479 = v_48388 | v_48478;
assign v_48481 = v_48476 | v_48480;
assign v_48483 = v_48387 | v_48482;
assign v_48485 = v_48385 | v_48484;
assign v_48487 = v_48482 | v_48486;
assign v_48489 = v_48384 | v_48488;
assign v_48491 = v_48382 | v_48490;
assign v_48493 = v_48488 | v_48492;
assign v_48495 = v_48381 | v_48494;
assign v_48497 = v_48379 | v_48496;
assign v_48499 = v_48494 | v_48498;
assign v_48501 = v_48378 | v_48500;
assign v_48503 = v_48376 | v_48502;
assign v_48505 = v_48500 | v_48504;
assign v_48507 = v_48375 | v_48506;
assign v_48509 = v_48373 | v_48508;
assign v_48511 = v_48506 | v_48510;
assign v_48513 = v_48372 | v_48512;
assign v_48515 = v_48370 | v_48514;
assign v_48517 = v_48512 | v_48516;
assign v_48520 = ~v_48369 | v_48519;
assign v_48527 = v_48417 | v_48526;
assign v_48530 = v_48528 | v_48529;
assign v_48532 = v_48414 | v_48531;
assign v_48535 = v_48533 | v_48534;
assign v_48537 = v_48411 | v_48536;
assign v_48540 = v_48538 | v_48539;
assign v_48542 = v_48408 | v_48541;
assign v_48545 = v_48543 | v_48544;
assign v_48547 = v_48405 | v_48546;
assign v_48550 = v_48548 | v_48549;
assign v_48552 = v_48402 | v_48551;
assign v_48555 = v_48553 | v_48554;
assign v_48557 = v_48399 | v_48556;
assign v_48560 = v_48558 | v_48559;
assign v_48562 = v_48396 | v_48561;
assign v_48565 = v_48563 | v_48564;
assign v_48567 = v_48393 | v_48566;
assign v_48570 = v_48568 | v_48569;
assign v_48572 = v_48390 | v_48571;
assign v_48575 = v_48573 | v_48574;
assign v_48577 = v_48387 | v_48576;
assign v_48580 = v_48578 | v_48579;
assign v_48582 = v_48384 | v_48581;
assign v_48585 = v_48583 | v_48584;
assign v_48587 = v_48381 | v_48586;
assign v_48590 = v_48588 | v_48589;
assign v_48592 = v_48378 | v_48591;
assign v_48595 = v_48593 | v_48594;
assign v_48597 = v_48375 | v_48596;
assign v_48600 = v_48598 | v_48599;
assign v_48602 = v_48372 | v_48601;
assign v_48605 = v_48603 | v_48604;
assign v_48607 = v_48369 | v_48606;
assign v_48610 = v_48368 | v_48609;
assign v_48664 = v_48661 | v_48663;
assign v_48666 = v_48660 | v_48665;
assign v_48668 = v_48658 | v_48667;
assign v_48670 = v_48665 | v_48669;
assign v_48672 = v_48657 | v_48671;
assign v_48674 = v_48655 | v_48673;
assign v_48676 = v_48671 | v_48675;
assign v_48678 = v_48654 | v_48677;
assign v_48680 = v_48652 | v_48679;
assign v_48682 = v_48677 | v_48681;
assign v_48684 = v_48651 | v_48683;
assign v_48686 = v_48649 | v_48685;
assign v_48688 = v_48683 | v_48687;
assign v_48690 = v_48648 | v_48689;
assign v_48692 = v_48646 | v_48691;
assign v_48694 = v_48689 | v_48693;
assign v_48696 = v_48645 | v_48695;
assign v_48698 = v_48643 | v_48697;
assign v_48700 = v_48695 | v_48699;
assign v_48702 = v_48642 | v_48701;
assign v_48704 = v_48640 | v_48703;
assign v_48706 = v_48701 | v_48705;
assign v_48708 = v_48639 | v_48707;
assign v_48710 = v_48637 | v_48709;
assign v_48712 = v_48707 | v_48711;
assign v_48714 = v_48636 | v_48713;
assign v_48716 = v_48634 | v_48715;
assign v_48718 = v_48713 | v_48717;
assign v_48720 = v_48633 | v_48719;
assign v_48722 = v_48631 | v_48721;
assign v_48724 = v_48719 | v_48723;
assign v_48726 = v_48630 | v_48725;
assign v_48728 = v_48628 | v_48727;
assign v_48730 = v_48725 | v_48729;
assign v_48732 = v_48627 | v_48731;
assign v_48734 = v_48625 | v_48733;
assign v_48736 = v_48731 | v_48735;
assign v_48738 = v_48624 | v_48737;
assign v_48740 = v_48622 | v_48739;
assign v_48742 = v_48737 | v_48741;
assign v_48744 = v_48621 | v_48743;
assign v_48746 = v_48619 | v_48745;
assign v_48748 = v_48743 | v_48747;
assign v_48750 = v_48618 | v_48749;
assign v_48752 = v_48616 | v_48751;
assign v_48754 = v_48749 | v_48753;
assign v_48756 = v_48615 | v_48755;
assign v_48758 = v_48613 | v_48757;
assign v_48760 = v_48755 | v_48759;
assign v_48763 = ~v_48612 | v_48762;
assign v_48770 = v_48660 | v_48769;
assign v_48773 = v_48771 | v_48772;
assign v_48775 = v_48657 | v_48774;
assign v_48778 = v_48776 | v_48777;
assign v_48780 = v_48654 | v_48779;
assign v_48783 = v_48781 | v_48782;
assign v_48785 = v_48651 | v_48784;
assign v_48788 = v_48786 | v_48787;
assign v_48790 = v_48648 | v_48789;
assign v_48793 = v_48791 | v_48792;
assign v_48795 = v_48645 | v_48794;
assign v_48798 = v_48796 | v_48797;
assign v_48800 = v_48642 | v_48799;
assign v_48803 = v_48801 | v_48802;
assign v_48805 = v_48639 | v_48804;
assign v_48808 = v_48806 | v_48807;
assign v_48810 = v_48636 | v_48809;
assign v_48813 = v_48811 | v_48812;
assign v_48815 = v_48633 | v_48814;
assign v_48818 = v_48816 | v_48817;
assign v_48820 = v_48630 | v_48819;
assign v_48823 = v_48821 | v_48822;
assign v_48825 = v_48627 | v_48824;
assign v_48828 = v_48826 | v_48827;
assign v_48830 = v_48624 | v_48829;
assign v_48833 = v_48831 | v_48832;
assign v_48835 = v_48621 | v_48834;
assign v_48838 = v_48836 | v_48837;
assign v_48840 = v_48618 | v_48839;
assign v_48843 = v_48841 | v_48842;
assign v_48845 = v_48615 | v_48844;
assign v_48848 = v_48846 | v_48847;
assign v_48850 = v_48612 | v_48849;
assign v_48853 = v_48611 | v_48852;
assign v_48907 = v_48904 | v_48906;
assign v_48909 = v_48903 | v_48908;
assign v_48911 = v_48901 | v_48910;
assign v_48913 = v_48908 | v_48912;
assign v_48915 = v_48900 | v_48914;
assign v_48917 = v_48898 | v_48916;
assign v_48919 = v_48914 | v_48918;
assign v_48921 = v_48897 | v_48920;
assign v_48923 = v_48895 | v_48922;
assign v_48925 = v_48920 | v_48924;
assign v_48927 = v_48894 | v_48926;
assign v_48929 = v_48892 | v_48928;
assign v_48931 = v_48926 | v_48930;
assign v_48933 = v_48891 | v_48932;
assign v_48935 = v_48889 | v_48934;
assign v_48937 = v_48932 | v_48936;
assign v_48939 = v_48888 | v_48938;
assign v_48941 = v_48886 | v_48940;
assign v_48943 = v_48938 | v_48942;
assign v_48945 = v_48885 | v_48944;
assign v_48947 = v_48883 | v_48946;
assign v_48949 = v_48944 | v_48948;
assign v_48951 = v_48882 | v_48950;
assign v_48953 = v_48880 | v_48952;
assign v_48955 = v_48950 | v_48954;
assign v_48957 = v_48879 | v_48956;
assign v_48959 = v_48877 | v_48958;
assign v_48961 = v_48956 | v_48960;
assign v_48963 = v_48876 | v_48962;
assign v_48965 = v_48874 | v_48964;
assign v_48967 = v_48962 | v_48966;
assign v_48969 = v_48873 | v_48968;
assign v_48971 = v_48871 | v_48970;
assign v_48973 = v_48968 | v_48972;
assign v_48975 = v_48870 | v_48974;
assign v_48977 = v_48868 | v_48976;
assign v_48979 = v_48974 | v_48978;
assign v_48981 = v_48867 | v_48980;
assign v_48983 = v_48865 | v_48982;
assign v_48985 = v_48980 | v_48984;
assign v_48987 = v_48864 | v_48986;
assign v_48989 = v_48862 | v_48988;
assign v_48991 = v_48986 | v_48990;
assign v_48993 = v_48861 | v_48992;
assign v_48995 = v_48859 | v_48994;
assign v_48997 = v_48992 | v_48996;
assign v_48999 = v_48858 | v_48998;
assign v_49001 = v_48856 | v_49000;
assign v_49003 = v_48998 | v_49002;
assign v_49006 = ~v_48855 | v_49005;
assign v_49013 = v_48903 | v_49012;
assign v_49016 = v_49014 | v_49015;
assign v_49018 = v_48900 | v_49017;
assign v_49021 = v_49019 | v_49020;
assign v_49023 = v_48897 | v_49022;
assign v_49026 = v_49024 | v_49025;
assign v_49028 = v_48894 | v_49027;
assign v_49031 = v_49029 | v_49030;
assign v_49033 = v_48891 | v_49032;
assign v_49036 = v_49034 | v_49035;
assign v_49038 = v_48888 | v_49037;
assign v_49041 = v_49039 | v_49040;
assign v_49043 = v_48885 | v_49042;
assign v_49046 = v_49044 | v_49045;
assign v_49048 = v_48882 | v_49047;
assign v_49051 = v_49049 | v_49050;
assign v_49053 = v_48879 | v_49052;
assign v_49056 = v_49054 | v_49055;
assign v_49058 = v_48876 | v_49057;
assign v_49061 = v_49059 | v_49060;
assign v_49063 = v_48873 | v_49062;
assign v_49066 = v_49064 | v_49065;
assign v_49068 = v_48870 | v_49067;
assign v_49071 = v_49069 | v_49070;
assign v_49073 = v_48867 | v_49072;
assign v_49076 = v_49074 | v_49075;
assign v_49078 = v_48864 | v_49077;
assign v_49081 = v_49079 | v_49080;
assign v_49083 = v_48861 | v_49082;
assign v_49086 = v_49084 | v_49085;
assign v_49088 = v_48858 | v_49087;
assign v_49091 = v_49089 | v_49090;
assign v_49093 = v_48855 | v_49092;
assign v_49096 = v_48854 | v_49095;
assign v_49150 = v_49147 | v_49149;
assign v_49152 = v_49146 | v_49151;
assign v_49154 = v_49144 | v_49153;
assign v_49156 = v_49151 | v_49155;
assign v_49158 = v_49143 | v_49157;
assign v_49160 = v_49141 | v_49159;
assign v_49162 = v_49157 | v_49161;
assign v_49164 = v_49140 | v_49163;
assign v_49166 = v_49138 | v_49165;
assign v_49168 = v_49163 | v_49167;
assign v_49170 = v_49137 | v_49169;
assign v_49172 = v_49135 | v_49171;
assign v_49174 = v_49169 | v_49173;
assign v_49176 = v_49134 | v_49175;
assign v_49178 = v_49132 | v_49177;
assign v_49180 = v_49175 | v_49179;
assign v_49182 = v_49131 | v_49181;
assign v_49184 = v_49129 | v_49183;
assign v_49186 = v_49181 | v_49185;
assign v_49188 = v_49128 | v_49187;
assign v_49190 = v_49126 | v_49189;
assign v_49192 = v_49187 | v_49191;
assign v_49194 = v_49125 | v_49193;
assign v_49196 = v_49123 | v_49195;
assign v_49198 = v_49193 | v_49197;
assign v_49200 = v_49122 | v_49199;
assign v_49202 = v_49120 | v_49201;
assign v_49204 = v_49199 | v_49203;
assign v_49206 = v_49119 | v_49205;
assign v_49208 = v_49117 | v_49207;
assign v_49210 = v_49205 | v_49209;
assign v_49212 = v_49116 | v_49211;
assign v_49214 = v_49114 | v_49213;
assign v_49216 = v_49211 | v_49215;
assign v_49218 = v_49113 | v_49217;
assign v_49220 = v_49111 | v_49219;
assign v_49222 = v_49217 | v_49221;
assign v_49224 = v_49110 | v_49223;
assign v_49226 = v_49108 | v_49225;
assign v_49228 = v_49223 | v_49227;
assign v_49230 = v_49107 | v_49229;
assign v_49232 = v_49105 | v_49231;
assign v_49234 = v_49229 | v_49233;
assign v_49236 = v_49104 | v_49235;
assign v_49238 = v_49102 | v_49237;
assign v_49240 = v_49235 | v_49239;
assign v_49242 = v_49101 | v_49241;
assign v_49244 = v_49099 | v_49243;
assign v_49246 = v_49241 | v_49245;
assign v_49249 = ~v_49098 | v_49248;
assign v_49256 = v_49146 | v_49255;
assign v_49259 = v_49257 | v_49258;
assign v_49261 = v_49143 | v_49260;
assign v_49264 = v_49262 | v_49263;
assign v_49266 = v_49140 | v_49265;
assign v_49269 = v_49267 | v_49268;
assign v_49271 = v_49137 | v_49270;
assign v_49274 = v_49272 | v_49273;
assign v_49276 = v_49134 | v_49275;
assign v_49279 = v_49277 | v_49278;
assign v_49281 = v_49131 | v_49280;
assign v_49284 = v_49282 | v_49283;
assign v_49286 = v_49128 | v_49285;
assign v_49289 = v_49287 | v_49288;
assign v_49291 = v_49125 | v_49290;
assign v_49294 = v_49292 | v_49293;
assign v_49296 = v_49122 | v_49295;
assign v_49299 = v_49297 | v_49298;
assign v_49301 = v_49119 | v_49300;
assign v_49304 = v_49302 | v_49303;
assign v_49306 = v_49116 | v_49305;
assign v_49309 = v_49307 | v_49308;
assign v_49311 = v_49113 | v_49310;
assign v_49314 = v_49312 | v_49313;
assign v_49316 = v_49110 | v_49315;
assign v_49319 = v_49317 | v_49318;
assign v_49321 = v_49107 | v_49320;
assign v_49324 = v_49322 | v_49323;
assign v_49326 = v_49104 | v_49325;
assign v_49329 = v_49327 | v_49328;
assign v_49331 = v_49101 | v_49330;
assign v_49334 = v_49332 | v_49333;
assign v_49336 = v_49098 | v_49335;
assign v_49339 = v_49097 | v_49338;
assign v_49393 = v_49390 | v_49392;
assign v_49395 = v_49389 | v_49394;
assign v_49397 = v_49387 | v_49396;
assign v_49399 = v_49394 | v_49398;
assign v_49401 = v_49386 | v_49400;
assign v_49403 = v_49384 | v_49402;
assign v_49405 = v_49400 | v_49404;
assign v_49407 = v_49383 | v_49406;
assign v_49409 = v_49381 | v_49408;
assign v_49411 = v_49406 | v_49410;
assign v_49413 = v_49380 | v_49412;
assign v_49415 = v_49378 | v_49414;
assign v_49417 = v_49412 | v_49416;
assign v_49419 = v_49377 | v_49418;
assign v_49421 = v_49375 | v_49420;
assign v_49423 = v_49418 | v_49422;
assign v_49425 = v_49374 | v_49424;
assign v_49427 = v_49372 | v_49426;
assign v_49429 = v_49424 | v_49428;
assign v_49431 = v_49371 | v_49430;
assign v_49433 = v_49369 | v_49432;
assign v_49435 = v_49430 | v_49434;
assign v_49437 = v_49368 | v_49436;
assign v_49439 = v_49366 | v_49438;
assign v_49441 = v_49436 | v_49440;
assign v_49443 = v_49365 | v_49442;
assign v_49445 = v_49363 | v_49444;
assign v_49447 = v_49442 | v_49446;
assign v_49449 = v_49362 | v_49448;
assign v_49451 = v_49360 | v_49450;
assign v_49453 = v_49448 | v_49452;
assign v_49455 = v_49359 | v_49454;
assign v_49457 = v_49357 | v_49456;
assign v_49459 = v_49454 | v_49458;
assign v_49461 = v_49356 | v_49460;
assign v_49463 = v_49354 | v_49462;
assign v_49465 = v_49460 | v_49464;
assign v_49467 = v_49353 | v_49466;
assign v_49469 = v_49351 | v_49468;
assign v_49471 = v_49466 | v_49470;
assign v_49473 = v_49350 | v_49472;
assign v_49475 = v_49348 | v_49474;
assign v_49477 = v_49472 | v_49476;
assign v_49479 = v_49347 | v_49478;
assign v_49481 = v_49345 | v_49480;
assign v_49483 = v_49478 | v_49482;
assign v_49485 = v_49344 | v_49484;
assign v_49487 = v_49342 | v_49486;
assign v_49489 = v_49484 | v_49488;
assign v_49492 = ~v_49341 | v_49491;
assign v_49499 = v_49389 | v_49498;
assign v_49502 = v_49500 | v_49501;
assign v_49504 = v_49386 | v_49503;
assign v_49507 = v_49505 | v_49506;
assign v_49509 = v_49383 | v_49508;
assign v_49512 = v_49510 | v_49511;
assign v_49514 = v_49380 | v_49513;
assign v_49517 = v_49515 | v_49516;
assign v_49519 = v_49377 | v_49518;
assign v_49522 = v_49520 | v_49521;
assign v_49524 = v_49374 | v_49523;
assign v_49527 = v_49525 | v_49526;
assign v_49529 = v_49371 | v_49528;
assign v_49532 = v_49530 | v_49531;
assign v_49534 = v_49368 | v_49533;
assign v_49537 = v_49535 | v_49536;
assign v_49539 = v_49365 | v_49538;
assign v_49542 = v_49540 | v_49541;
assign v_49544 = v_49362 | v_49543;
assign v_49547 = v_49545 | v_49546;
assign v_49549 = v_49359 | v_49548;
assign v_49552 = v_49550 | v_49551;
assign v_49554 = v_49356 | v_49553;
assign v_49557 = v_49555 | v_49556;
assign v_49559 = v_49353 | v_49558;
assign v_49562 = v_49560 | v_49561;
assign v_49564 = v_49350 | v_49563;
assign v_49567 = v_49565 | v_49566;
assign v_49569 = v_49347 | v_49568;
assign v_49572 = v_49570 | v_49571;
assign v_49574 = v_49344 | v_49573;
assign v_49577 = v_49575 | v_49576;
assign v_49579 = v_49341 | v_49578;
assign v_49582 = v_49340 | v_49581;
assign v_49636 = v_49633 | v_49635;
assign v_49638 = v_49632 | v_49637;
assign v_49640 = v_49630 | v_49639;
assign v_49642 = v_49637 | v_49641;
assign v_49644 = v_49629 | v_49643;
assign v_49646 = v_49627 | v_49645;
assign v_49648 = v_49643 | v_49647;
assign v_49650 = v_49626 | v_49649;
assign v_49652 = v_49624 | v_49651;
assign v_49654 = v_49649 | v_49653;
assign v_49656 = v_49623 | v_49655;
assign v_49658 = v_49621 | v_49657;
assign v_49660 = v_49655 | v_49659;
assign v_49662 = v_49620 | v_49661;
assign v_49664 = v_49618 | v_49663;
assign v_49666 = v_49661 | v_49665;
assign v_49668 = v_49617 | v_49667;
assign v_49670 = v_49615 | v_49669;
assign v_49672 = v_49667 | v_49671;
assign v_49674 = v_49614 | v_49673;
assign v_49676 = v_49612 | v_49675;
assign v_49678 = v_49673 | v_49677;
assign v_49680 = v_49611 | v_49679;
assign v_49682 = v_49609 | v_49681;
assign v_49684 = v_49679 | v_49683;
assign v_49686 = v_49608 | v_49685;
assign v_49688 = v_49606 | v_49687;
assign v_49690 = v_49685 | v_49689;
assign v_49692 = v_49605 | v_49691;
assign v_49694 = v_49603 | v_49693;
assign v_49696 = v_49691 | v_49695;
assign v_49698 = v_49602 | v_49697;
assign v_49700 = v_49600 | v_49699;
assign v_49702 = v_49697 | v_49701;
assign v_49704 = v_49599 | v_49703;
assign v_49706 = v_49597 | v_49705;
assign v_49708 = v_49703 | v_49707;
assign v_49710 = v_49596 | v_49709;
assign v_49712 = v_49594 | v_49711;
assign v_49714 = v_49709 | v_49713;
assign v_49716 = v_49593 | v_49715;
assign v_49718 = v_49591 | v_49717;
assign v_49720 = v_49715 | v_49719;
assign v_49722 = v_49590 | v_49721;
assign v_49724 = v_49588 | v_49723;
assign v_49726 = v_49721 | v_49725;
assign v_49728 = v_49587 | v_49727;
assign v_49730 = v_49585 | v_49729;
assign v_49732 = v_49727 | v_49731;
assign v_49735 = ~v_49584 | v_49734;
assign v_49742 = v_49632 | v_49741;
assign v_49745 = v_49743 | v_49744;
assign v_49747 = v_49629 | v_49746;
assign v_49750 = v_49748 | v_49749;
assign v_49752 = v_49626 | v_49751;
assign v_49755 = v_49753 | v_49754;
assign v_49757 = v_49623 | v_49756;
assign v_49760 = v_49758 | v_49759;
assign v_49762 = v_49620 | v_49761;
assign v_49765 = v_49763 | v_49764;
assign v_49767 = v_49617 | v_49766;
assign v_49770 = v_49768 | v_49769;
assign v_49772 = v_49614 | v_49771;
assign v_49775 = v_49773 | v_49774;
assign v_49777 = v_49611 | v_49776;
assign v_49780 = v_49778 | v_49779;
assign v_49782 = v_49608 | v_49781;
assign v_49785 = v_49783 | v_49784;
assign v_49787 = v_49605 | v_49786;
assign v_49790 = v_49788 | v_49789;
assign v_49792 = v_49602 | v_49791;
assign v_49795 = v_49793 | v_49794;
assign v_49797 = v_49599 | v_49796;
assign v_49800 = v_49798 | v_49799;
assign v_49802 = v_49596 | v_49801;
assign v_49805 = v_49803 | v_49804;
assign v_49807 = v_49593 | v_49806;
assign v_49810 = v_49808 | v_49809;
assign v_49812 = v_49590 | v_49811;
assign v_49815 = v_49813 | v_49814;
assign v_49817 = v_49587 | v_49816;
assign v_49820 = v_49818 | v_49819;
assign v_49822 = v_49584 | v_49821;
assign v_49825 = v_49583 | v_49824;
assign v_49878 = v_49875 | v_49877;
assign v_49880 = v_49874 | v_49879;
assign v_49882 = v_49872 | v_49881;
assign v_49884 = v_49879 | v_49883;
assign v_49886 = v_49871 | v_49885;
assign v_49888 = v_49869 | v_49887;
assign v_49890 = v_49885 | v_49889;
assign v_49892 = v_49868 | v_49891;
assign v_49894 = v_49866 | v_49893;
assign v_49896 = v_49891 | v_49895;
assign v_49898 = v_49865 | v_49897;
assign v_49900 = v_49863 | v_49899;
assign v_49902 = v_49897 | v_49901;
assign v_49904 = v_49862 | v_49903;
assign v_49906 = v_49860 | v_49905;
assign v_49908 = v_49903 | v_49907;
assign v_49910 = v_49859 | v_49909;
assign v_49912 = v_49857 | v_49911;
assign v_49914 = v_49909 | v_49913;
assign v_49916 = v_49856 | v_49915;
assign v_49918 = v_49854 | v_49917;
assign v_49920 = v_49915 | v_49919;
assign v_49922 = v_49853 | v_49921;
assign v_49924 = v_49851 | v_49923;
assign v_49926 = v_49921 | v_49925;
assign v_49928 = v_49850 | v_49927;
assign v_49930 = v_49848 | v_49929;
assign v_49932 = v_49927 | v_49931;
assign v_49934 = v_49847 | v_49933;
assign v_49936 = v_49845 | v_49935;
assign v_49938 = v_49933 | v_49937;
assign v_49940 = v_49844 | v_49939;
assign v_49942 = v_49842 | v_49941;
assign v_49944 = v_49939 | v_49943;
assign v_49946 = v_49841 | v_49945;
assign v_49948 = v_49839 | v_49947;
assign v_49950 = v_49945 | v_49949;
assign v_49952 = v_49838 | v_49951;
assign v_49954 = v_49836 | v_49953;
assign v_49956 = v_49951 | v_49955;
assign v_49958 = v_49835 | v_49957;
assign v_49960 = v_49833 | v_49959;
assign v_49962 = v_49957 | v_49961;
assign v_49964 = v_49832 | v_49963;
assign v_49966 = v_49830 | v_49965;
assign v_49968 = v_49963 | v_49967;
assign v_49970 = v_49829 | v_49969;
assign v_49972 = v_49827 | v_49971;
assign v_49974 = v_49969 | v_49973;
assign v_49978 = v_49975 | v_49977;
assign v_49985 = v_49874 | v_49984;
assign v_49988 = v_49986 | v_49987;
assign v_49990 = v_49871 | v_49989;
assign v_49993 = v_49991 | v_49992;
assign v_49995 = v_49868 | v_49994;
assign v_49998 = v_49996 | v_49997;
assign v_50000 = v_49865 | v_49999;
assign v_50003 = v_50001 | v_50002;
assign v_50005 = v_49862 | v_50004;
assign v_50008 = v_50006 | v_50007;
assign v_50010 = v_49859 | v_50009;
assign v_50013 = v_50011 | v_50012;
assign v_50015 = v_49856 | v_50014;
assign v_50018 = v_50016 | v_50017;
assign v_50020 = v_49853 | v_50019;
assign v_50023 = v_50021 | v_50022;
assign v_50025 = v_49850 | v_50024;
assign v_50028 = v_50026 | v_50027;
assign v_50030 = v_49847 | v_50029;
assign v_50033 = v_50031 | v_50032;
assign v_50035 = v_49844 | v_50034;
assign v_50038 = v_50036 | v_50037;
assign v_50040 = v_49841 | v_50039;
assign v_50043 = v_50041 | v_50042;
assign v_50045 = v_49838 | v_50044;
assign v_50048 = v_50046 | v_50047;
assign v_50050 = v_49835 | v_50049;
assign v_50053 = v_50051 | v_50052;
assign v_50055 = v_49832 | v_50054;
assign v_50058 = v_50056 | v_50057;
assign v_50060 = v_49829 | v_50059;
assign v_50063 = v_50061 | v_50062;
assign v_50065 = v_50063 | v_50064;
assign v_50068 = v_49826 | v_50067;
assign v_50139 = v_50136 | v_50138;
assign v_50141 = v_50134 | v_50140;
assign v_50143 = v_50132 | v_50142;
assign v_50145 = v_50140 | v_50144;
assign v_50147 = v_50130 | v_50146;
assign v_50149 = v_50128 | v_50148;
assign v_50151 = v_50146 | v_50150;
assign v_50153 = v_50126 | v_50152;
assign v_50155 = v_50124 | v_50154;
assign v_50157 = v_50152 | v_50156;
assign v_50159 = v_50122 | v_50158;
assign v_50161 = v_50120 | v_50160;
assign v_50163 = v_50158 | v_50162;
assign v_50165 = v_50118 | v_50164;
assign v_50167 = v_50116 | v_50166;
assign v_50169 = v_50164 | v_50168;
assign v_50171 = v_50114 | v_50170;
assign v_50173 = v_50112 | v_50172;
assign v_50175 = v_50170 | v_50174;
assign v_50177 = v_50110 | v_50176;
assign v_50179 = v_50108 | v_50178;
assign v_50181 = v_50176 | v_50180;
assign v_50183 = v_50106 | v_50182;
assign v_50185 = v_50104 | v_50184;
assign v_50187 = v_50182 | v_50186;
assign v_50189 = v_50102 | v_50188;
assign v_50191 = v_50100 | v_50190;
assign v_50193 = v_50188 | v_50192;
assign v_50195 = v_50098 | v_50194;
assign v_50197 = v_50096 | v_50196;
assign v_50199 = v_50194 | v_50198;
assign v_50201 = v_50094 | v_50200;
assign v_50203 = v_50092 | v_50202;
assign v_50205 = v_50200 | v_50204;
assign v_50207 = v_50090 | v_50206;
assign v_50209 = v_50088 | v_50208;
assign v_50211 = v_50206 | v_50210;
assign v_50213 = v_50086 | v_50212;
assign v_50215 = v_50083 | v_50214;
assign v_50217 = v_50212 | v_50216;
assign v_50219 = v_50082 | v_50218;
assign v_50221 = v_50079 | v_50220;
assign v_50223 = v_50218 | v_50222;
assign v_50225 = v_50078 | v_50224;
assign v_50227 = v_50075 | v_50226;
assign v_50229 = v_50224 | v_50228;
assign v_50231 = v_50074 | v_50230;
assign v_50233 = v_50071 | v_50232;
assign v_50235 = v_50230 | v_50234;
assign v_50238 = ~v_50070 | v_50237;
assign v_50245 = v_50134 | v_50244;
assign v_50248 = v_50246 | v_50247;
assign v_50250 = v_50130 | v_50249;
assign v_50253 = v_50251 | v_50252;
assign v_50255 = v_50126 | v_50254;
assign v_50258 = v_50256 | v_50257;
assign v_50260 = v_50122 | v_50259;
assign v_50263 = v_50261 | v_50262;
assign v_50265 = v_50118 | v_50264;
assign v_50268 = v_50266 | v_50267;
assign v_50270 = v_50114 | v_50269;
assign v_50273 = v_50271 | v_50272;
assign v_50275 = v_50110 | v_50274;
assign v_50278 = v_50276 | v_50277;
assign v_50280 = v_50106 | v_50279;
assign v_50283 = v_50281 | v_50282;
assign v_50285 = v_50102 | v_50284;
assign v_50288 = v_50286 | v_50287;
assign v_50290 = v_50098 | v_50289;
assign v_50293 = v_50291 | v_50292;
assign v_50295 = v_50094 | v_50294;
assign v_50298 = v_50296 | v_50297;
assign v_50300 = v_50090 | v_50299;
assign v_50303 = v_50301 | v_50302;
assign v_50305 = v_50086 | v_50304;
assign v_50308 = v_50306 | v_50307;
assign v_50310 = v_50082 | v_50309;
assign v_50313 = v_50311 | v_50312;
assign v_50315 = v_50078 | v_50314;
assign v_50318 = v_50316 | v_50317;
assign v_50320 = v_50074 | v_50319;
assign v_50323 = v_50321 | v_50322;
assign v_50325 = v_50070 | v_50324;
assign v_50328 = v_50069 | v_50327;
assign v_50382 = v_50379 | v_50381;
assign v_50384 = v_50378 | v_50383;
assign v_50386 = v_50376 | v_50385;
assign v_50388 = v_50383 | v_50387;
assign v_50390 = v_50375 | v_50389;
assign v_50392 = v_50373 | v_50391;
assign v_50394 = v_50389 | v_50393;
assign v_50396 = v_50372 | v_50395;
assign v_50398 = v_50370 | v_50397;
assign v_50400 = v_50395 | v_50399;
assign v_50402 = v_50369 | v_50401;
assign v_50404 = v_50367 | v_50403;
assign v_50406 = v_50401 | v_50405;
assign v_50408 = v_50366 | v_50407;
assign v_50410 = v_50364 | v_50409;
assign v_50412 = v_50407 | v_50411;
assign v_50414 = v_50363 | v_50413;
assign v_50416 = v_50361 | v_50415;
assign v_50418 = v_50413 | v_50417;
assign v_50420 = v_50360 | v_50419;
assign v_50422 = v_50358 | v_50421;
assign v_50424 = v_50419 | v_50423;
assign v_50426 = v_50357 | v_50425;
assign v_50428 = v_50355 | v_50427;
assign v_50430 = v_50425 | v_50429;
assign v_50432 = v_50354 | v_50431;
assign v_50434 = v_50352 | v_50433;
assign v_50436 = v_50431 | v_50435;
assign v_50438 = v_50351 | v_50437;
assign v_50440 = v_50349 | v_50439;
assign v_50442 = v_50437 | v_50441;
assign v_50444 = v_50348 | v_50443;
assign v_50446 = v_50346 | v_50445;
assign v_50448 = v_50443 | v_50447;
assign v_50450 = v_50345 | v_50449;
assign v_50452 = v_50343 | v_50451;
assign v_50454 = v_50449 | v_50453;
assign v_50456 = v_50342 | v_50455;
assign v_50458 = v_50340 | v_50457;
assign v_50460 = v_50455 | v_50459;
assign v_50462 = v_50339 | v_50461;
assign v_50464 = v_50337 | v_50463;
assign v_50466 = v_50461 | v_50465;
assign v_50468 = v_50336 | v_50467;
assign v_50470 = v_50334 | v_50469;
assign v_50472 = v_50467 | v_50471;
assign v_50474 = v_50333 | v_50473;
assign v_50476 = v_50331 | v_50475;
assign v_50478 = v_50473 | v_50477;
assign v_50481 = ~v_50330 | v_50480;
assign v_50488 = v_50378 | v_50487;
assign v_50491 = v_50489 | v_50490;
assign v_50493 = v_50375 | v_50492;
assign v_50496 = v_50494 | v_50495;
assign v_50498 = v_50372 | v_50497;
assign v_50501 = v_50499 | v_50500;
assign v_50503 = v_50369 | v_50502;
assign v_50506 = v_50504 | v_50505;
assign v_50508 = v_50366 | v_50507;
assign v_50511 = v_50509 | v_50510;
assign v_50513 = v_50363 | v_50512;
assign v_50516 = v_50514 | v_50515;
assign v_50518 = v_50360 | v_50517;
assign v_50521 = v_50519 | v_50520;
assign v_50523 = v_50357 | v_50522;
assign v_50526 = v_50524 | v_50525;
assign v_50528 = v_50354 | v_50527;
assign v_50531 = v_50529 | v_50530;
assign v_50533 = v_50351 | v_50532;
assign v_50536 = v_50534 | v_50535;
assign v_50538 = v_50348 | v_50537;
assign v_50541 = v_50539 | v_50540;
assign v_50543 = v_50345 | v_50542;
assign v_50546 = v_50544 | v_50545;
assign v_50548 = v_50342 | v_50547;
assign v_50551 = v_50549 | v_50550;
assign v_50553 = v_50339 | v_50552;
assign v_50556 = v_50554 | v_50555;
assign v_50558 = v_50336 | v_50557;
assign v_50561 = v_50559 | v_50560;
assign v_50563 = v_50333 | v_50562;
assign v_50566 = v_50564 | v_50565;
assign v_50568 = v_50330 | v_50567;
assign v_50571 = v_50329 | v_50570;
assign v_50625 = v_50622 | v_50624;
assign v_50627 = v_50621 | v_50626;
assign v_50629 = v_50619 | v_50628;
assign v_50631 = v_50626 | v_50630;
assign v_50633 = v_50618 | v_50632;
assign v_50635 = v_50616 | v_50634;
assign v_50637 = v_50632 | v_50636;
assign v_50639 = v_50615 | v_50638;
assign v_50641 = v_50613 | v_50640;
assign v_50643 = v_50638 | v_50642;
assign v_50645 = v_50612 | v_50644;
assign v_50647 = v_50610 | v_50646;
assign v_50649 = v_50644 | v_50648;
assign v_50651 = v_50609 | v_50650;
assign v_50653 = v_50607 | v_50652;
assign v_50655 = v_50650 | v_50654;
assign v_50657 = v_50606 | v_50656;
assign v_50659 = v_50604 | v_50658;
assign v_50661 = v_50656 | v_50660;
assign v_50663 = v_50603 | v_50662;
assign v_50665 = v_50601 | v_50664;
assign v_50667 = v_50662 | v_50666;
assign v_50669 = v_50600 | v_50668;
assign v_50671 = v_50598 | v_50670;
assign v_50673 = v_50668 | v_50672;
assign v_50675 = v_50597 | v_50674;
assign v_50677 = v_50595 | v_50676;
assign v_50679 = v_50674 | v_50678;
assign v_50681 = v_50594 | v_50680;
assign v_50683 = v_50592 | v_50682;
assign v_50685 = v_50680 | v_50684;
assign v_50687 = v_50591 | v_50686;
assign v_50689 = v_50589 | v_50688;
assign v_50691 = v_50686 | v_50690;
assign v_50693 = v_50588 | v_50692;
assign v_50695 = v_50586 | v_50694;
assign v_50697 = v_50692 | v_50696;
assign v_50699 = v_50585 | v_50698;
assign v_50701 = v_50583 | v_50700;
assign v_50703 = v_50698 | v_50702;
assign v_50705 = v_50582 | v_50704;
assign v_50707 = v_50580 | v_50706;
assign v_50709 = v_50704 | v_50708;
assign v_50711 = v_50579 | v_50710;
assign v_50713 = v_50577 | v_50712;
assign v_50715 = v_50710 | v_50714;
assign v_50717 = v_50576 | v_50716;
assign v_50719 = v_50574 | v_50718;
assign v_50721 = v_50716 | v_50720;
assign v_50724 = ~v_50573 | v_50723;
assign v_50731 = v_50621 | v_50730;
assign v_50734 = v_50732 | v_50733;
assign v_50736 = v_50618 | v_50735;
assign v_50739 = v_50737 | v_50738;
assign v_50741 = v_50615 | v_50740;
assign v_50744 = v_50742 | v_50743;
assign v_50746 = v_50612 | v_50745;
assign v_50749 = v_50747 | v_50748;
assign v_50751 = v_50609 | v_50750;
assign v_50754 = v_50752 | v_50753;
assign v_50756 = v_50606 | v_50755;
assign v_50759 = v_50757 | v_50758;
assign v_50761 = v_50603 | v_50760;
assign v_50764 = v_50762 | v_50763;
assign v_50766 = v_50600 | v_50765;
assign v_50769 = v_50767 | v_50768;
assign v_50771 = v_50597 | v_50770;
assign v_50774 = v_50772 | v_50773;
assign v_50776 = v_50594 | v_50775;
assign v_50779 = v_50777 | v_50778;
assign v_50781 = v_50591 | v_50780;
assign v_50784 = v_50782 | v_50783;
assign v_50786 = v_50588 | v_50785;
assign v_50789 = v_50787 | v_50788;
assign v_50791 = v_50585 | v_50790;
assign v_50794 = v_50792 | v_50793;
assign v_50796 = v_50582 | v_50795;
assign v_50799 = v_50797 | v_50798;
assign v_50801 = v_50579 | v_50800;
assign v_50804 = v_50802 | v_50803;
assign v_50806 = v_50576 | v_50805;
assign v_50809 = v_50807 | v_50808;
assign v_50811 = v_50573 | v_50810;
assign v_50814 = v_50572 | v_50813;
assign v_50868 = v_50865 | v_50867;
assign v_50870 = v_50864 | v_50869;
assign v_50872 = v_50862 | v_50871;
assign v_50874 = v_50869 | v_50873;
assign v_50876 = v_50861 | v_50875;
assign v_50878 = v_50859 | v_50877;
assign v_50880 = v_50875 | v_50879;
assign v_50882 = v_50858 | v_50881;
assign v_50884 = v_50856 | v_50883;
assign v_50886 = v_50881 | v_50885;
assign v_50888 = v_50855 | v_50887;
assign v_50890 = v_50853 | v_50889;
assign v_50892 = v_50887 | v_50891;
assign v_50894 = v_50852 | v_50893;
assign v_50896 = v_50850 | v_50895;
assign v_50898 = v_50893 | v_50897;
assign v_50900 = v_50849 | v_50899;
assign v_50902 = v_50847 | v_50901;
assign v_50904 = v_50899 | v_50903;
assign v_50906 = v_50846 | v_50905;
assign v_50908 = v_50844 | v_50907;
assign v_50910 = v_50905 | v_50909;
assign v_50912 = v_50843 | v_50911;
assign v_50914 = v_50841 | v_50913;
assign v_50916 = v_50911 | v_50915;
assign v_50918 = v_50840 | v_50917;
assign v_50920 = v_50838 | v_50919;
assign v_50922 = v_50917 | v_50921;
assign v_50924 = v_50837 | v_50923;
assign v_50926 = v_50835 | v_50925;
assign v_50928 = v_50923 | v_50927;
assign v_50930 = v_50834 | v_50929;
assign v_50932 = v_50832 | v_50931;
assign v_50934 = v_50929 | v_50933;
assign v_50936 = v_50831 | v_50935;
assign v_50938 = v_50829 | v_50937;
assign v_50940 = v_50935 | v_50939;
assign v_50942 = v_50828 | v_50941;
assign v_50944 = v_50826 | v_50943;
assign v_50946 = v_50941 | v_50945;
assign v_50948 = v_50825 | v_50947;
assign v_50950 = v_50823 | v_50949;
assign v_50952 = v_50947 | v_50951;
assign v_50954 = v_50822 | v_50953;
assign v_50956 = v_50820 | v_50955;
assign v_50958 = v_50953 | v_50957;
assign v_50960 = v_50819 | v_50959;
assign v_50962 = v_50817 | v_50961;
assign v_50964 = v_50959 | v_50963;
assign v_50967 = ~v_50816 | v_50966;
assign v_50974 = v_50864 | v_50973;
assign v_50977 = v_50975 | v_50976;
assign v_50979 = v_50861 | v_50978;
assign v_50982 = v_50980 | v_50981;
assign v_50984 = v_50858 | v_50983;
assign v_50987 = v_50985 | v_50986;
assign v_50989 = v_50855 | v_50988;
assign v_50992 = v_50990 | v_50991;
assign v_50994 = v_50852 | v_50993;
assign v_50997 = v_50995 | v_50996;
assign v_50999 = v_50849 | v_50998;
assign v_51002 = v_51000 | v_51001;
assign v_51004 = v_50846 | v_51003;
assign v_51007 = v_51005 | v_51006;
assign v_51009 = v_50843 | v_51008;
assign v_51012 = v_51010 | v_51011;
assign v_51014 = v_50840 | v_51013;
assign v_51017 = v_51015 | v_51016;
assign v_51019 = v_50837 | v_51018;
assign v_51022 = v_51020 | v_51021;
assign v_51024 = v_50834 | v_51023;
assign v_51027 = v_51025 | v_51026;
assign v_51029 = v_50831 | v_51028;
assign v_51032 = v_51030 | v_51031;
assign v_51034 = v_50828 | v_51033;
assign v_51037 = v_51035 | v_51036;
assign v_51039 = v_50825 | v_51038;
assign v_51042 = v_51040 | v_51041;
assign v_51044 = v_50822 | v_51043;
assign v_51047 = v_51045 | v_51046;
assign v_51049 = v_50819 | v_51048;
assign v_51052 = v_51050 | v_51051;
assign v_51054 = v_50816 | v_51053;
assign v_51057 = v_50815 | v_51056;
assign v_51111 = v_51108 | v_51110;
assign v_51113 = v_51107 | v_51112;
assign v_51115 = v_51105 | v_51114;
assign v_51117 = v_51112 | v_51116;
assign v_51119 = v_51104 | v_51118;
assign v_51121 = v_51102 | v_51120;
assign v_51123 = v_51118 | v_51122;
assign v_51125 = v_51101 | v_51124;
assign v_51127 = v_51099 | v_51126;
assign v_51129 = v_51124 | v_51128;
assign v_51131 = v_51098 | v_51130;
assign v_51133 = v_51096 | v_51132;
assign v_51135 = v_51130 | v_51134;
assign v_51137 = v_51095 | v_51136;
assign v_51139 = v_51093 | v_51138;
assign v_51141 = v_51136 | v_51140;
assign v_51143 = v_51092 | v_51142;
assign v_51145 = v_51090 | v_51144;
assign v_51147 = v_51142 | v_51146;
assign v_51149 = v_51089 | v_51148;
assign v_51151 = v_51087 | v_51150;
assign v_51153 = v_51148 | v_51152;
assign v_51155 = v_51086 | v_51154;
assign v_51157 = v_51084 | v_51156;
assign v_51159 = v_51154 | v_51158;
assign v_51161 = v_51083 | v_51160;
assign v_51163 = v_51081 | v_51162;
assign v_51165 = v_51160 | v_51164;
assign v_51167 = v_51080 | v_51166;
assign v_51169 = v_51078 | v_51168;
assign v_51171 = v_51166 | v_51170;
assign v_51173 = v_51077 | v_51172;
assign v_51175 = v_51075 | v_51174;
assign v_51177 = v_51172 | v_51176;
assign v_51179 = v_51074 | v_51178;
assign v_51181 = v_51072 | v_51180;
assign v_51183 = v_51178 | v_51182;
assign v_51185 = v_51071 | v_51184;
assign v_51187 = v_51069 | v_51186;
assign v_51189 = v_51184 | v_51188;
assign v_51191 = v_51068 | v_51190;
assign v_51193 = v_51066 | v_51192;
assign v_51195 = v_51190 | v_51194;
assign v_51197 = v_51065 | v_51196;
assign v_51199 = v_51063 | v_51198;
assign v_51201 = v_51196 | v_51200;
assign v_51203 = v_51062 | v_51202;
assign v_51205 = v_51060 | v_51204;
assign v_51207 = v_51202 | v_51206;
assign v_51210 = ~v_51059 | v_51209;
assign v_51217 = v_51107 | v_51216;
assign v_51220 = v_51218 | v_51219;
assign v_51222 = v_51104 | v_51221;
assign v_51225 = v_51223 | v_51224;
assign v_51227 = v_51101 | v_51226;
assign v_51230 = v_51228 | v_51229;
assign v_51232 = v_51098 | v_51231;
assign v_51235 = v_51233 | v_51234;
assign v_51237 = v_51095 | v_51236;
assign v_51240 = v_51238 | v_51239;
assign v_51242 = v_51092 | v_51241;
assign v_51245 = v_51243 | v_51244;
assign v_51247 = v_51089 | v_51246;
assign v_51250 = v_51248 | v_51249;
assign v_51252 = v_51086 | v_51251;
assign v_51255 = v_51253 | v_51254;
assign v_51257 = v_51083 | v_51256;
assign v_51260 = v_51258 | v_51259;
assign v_51262 = v_51080 | v_51261;
assign v_51265 = v_51263 | v_51264;
assign v_51267 = v_51077 | v_51266;
assign v_51270 = v_51268 | v_51269;
assign v_51272 = v_51074 | v_51271;
assign v_51275 = v_51273 | v_51274;
assign v_51277 = v_51071 | v_51276;
assign v_51280 = v_51278 | v_51279;
assign v_51282 = v_51068 | v_51281;
assign v_51285 = v_51283 | v_51284;
assign v_51287 = v_51065 | v_51286;
assign v_51290 = v_51288 | v_51289;
assign v_51292 = v_51062 | v_51291;
assign v_51295 = v_51293 | v_51294;
assign v_51297 = v_51059 | v_51296;
assign v_51300 = v_51058 | v_51299;
assign v_51354 = v_51351 | v_51353;
assign v_51356 = v_51350 | v_51355;
assign v_51358 = v_51348 | v_51357;
assign v_51360 = v_51355 | v_51359;
assign v_51362 = v_51347 | v_51361;
assign v_51364 = v_51345 | v_51363;
assign v_51366 = v_51361 | v_51365;
assign v_51368 = v_51344 | v_51367;
assign v_51370 = v_51342 | v_51369;
assign v_51372 = v_51367 | v_51371;
assign v_51374 = v_51341 | v_51373;
assign v_51376 = v_51339 | v_51375;
assign v_51378 = v_51373 | v_51377;
assign v_51380 = v_51338 | v_51379;
assign v_51382 = v_51336 | v_51381;
assign v_51384 = v_51379 | v_51383;
assign v_51386 = v_51335 | v_51385;
assign v_51388 = v_51333 | v_51387;
assign v_51390 = v_51385 | v_51389;
assign v_51392 = v_51332 | v_51391;
assign v_51394 = v_51330 | v_51393;
assign v_51396 = v_51391 | v_51395;
assign v_51398 = v_51329 | v_51397;
assign v_51400 = v_51327 | v_51399;
assign v_51402 = v_51397 | v_51401;
assign v_51404 = v_51326 | v_51403;
assign v_51406 = v_51324 | v_51405;
assign v_51408 = v_51403 | v_51407;
assign v_51410 = v_51323 | v_51409;
assign v_51412 = v_51321 | v_51411;
assign v_51414 = v_51409 | v_51413;
assign v_51416 = v_51320 | v_51415;
assign v_51418 = v_51318 | v_51417;
assign v_51420 = v_51415 | v_51419;
assign v_51422 = v_51317 | v_51421;
assign v_51424 = v_51315 | v_51423;
assign v_51426 = v_51421 | v_51425;
assign v_51428 = v_51314 | v_51427;
assign v_51430 = v_51312 | v_51429;
assign v_51432 = v_51427 | v_51431;
assign v_51434 = v_51311 | v_51433;
assign v_51436 = v_51309 | v_51435;
assign v_51438 = v_51433 | v_51437;
assign v_51440 = v_51308 | v_51439;
assign v_51442 = v_51306 | v_51441;
assign v_51444 = v_51439 | v_51443;
assign v_51446 = v_51305 | v_51445;
assign v_51448 = v_51303 | v_51447;
assign v_51450 = v_51445 | v_51449;
assign v_51453 = ~v_51302 | v_51452;
assign v_51460 = v_51350 | v_51459;
assign v_51463 = v_51461 | v_51462;
assign v_51465 = v_51347 | v_51464;
assign v_51468 = v_51466 | v_51467;
assign v_51470 = v_51344 | v_51469;
assign v_51473 = v_51471 | v_51472;
assign v_51475 = v_51341 | v_51474;
assign v_51478 = v_51476 | v_51477;
assign v_51480 = v_51338 | v_51479;
assign v_51483 = v_51481 | v_51482;
assign v_51485 = v_51335 | v_51484;
assign v_51488 = v_51486 | v_51487;
assign v_51490 = v_51332 | v_51489;
assign v_51493 = v_51491 | v_51492;
assign v_51495 = v_51329 | v_51494;
assign v_51498 = v_51496 | v_51497;
assign v_51500 = v_51326 | v_51499;
assign v_51503 = v_51501 | v_51502;
assign v_51505 = v_51323 | v_51504;
assign v_51508 = v_51506 | v_51507;
assign v_51510 = v_51320 | v_51509;
assign v_51513 = v_51511 | v_51512;
assign v_51515 = v_51317 | v_51514;
assign v_51518 = v_51516 | v_51517;
assign v_51520 = v_51314 | v_51519;
assign v_51523 = v_51521 | v_51522;
assign v_51525 = v_51311 | v_51524;
assign v_51528 = v_51526 | v_51527;
assign v_51530 = v_51308 | v_51529;
assign v_51533 = v_51531 | v_51532;
assign v_51535 = v_51305 | v_51534;
assign v_51538 = v_51536 | v_51537;
assign v_51540 = v_51302 | v_51539;
assign v_51543 = v_51301 | v_51542;
assign v_51597 = v_51594 | v_51596;
assign v_51599 = v_51593 | v_51598;
assign v_51601 = v_51591 | v_51600;
assign v_51603 = v_51598 | v_51602;
assign v_51605 = v_51590 | v_51604;
assign v_51607 = v_51588 | v_51606;
assign v_51609 = v_51604 | v_51608;
assign v_51611 = v_51587 | v_51610;
assign v_51613 = v_51585 | v_51612;
assign v_51615 = v_51610 | v_51614;
assign v_51617 = v_51584 | v_51616;
assign v_51619 = v_51582 | v_51618;
assign v_51621 = v_51616 | v_51620;
assign v_51623 = v_51581 | v_51622;
assign v_51625 = v_51579 | v_51624;
assign v_51627 = v_51622 | v_51626;
assign v_51629 = v_51578 | v_51628;
assign v_51631 = v_51576 | v_51630;
assign v_51633 = v_51628 | v_51632;
assign v_51635 = v_51575 | v_51634;
assign v_51637 = v_51573 | v_51636;
assign v_51639 = v_51634 | v_51638;
assign v_51641 = v_51572 | v_51640;
assign v_51643 = v_51570 | v_51642;
assign v_51645 = v_51640 | v_51644;
assign v_51647 = v_51569 | v_51646;
assign v_51649 = v_51567 | v_51648;
assign v_51651 = v_51646 | v_51650;
assign v_51653 = v_51566 | v_51652;
assign v_51655 = v_51564 | v_51654;
assign v_51657 = v_51652 | v_51656;
assign v_51659 = v_51563 | v_51658;
assign v_51661 = v_51561 | v_51660;
assign v_51663 = v_51658 | v_51662;
assign v_51665 = v_51560 | v_51664;
assign v_51667 = v_51558 | v_51666;
assign v_51669 = v_51664 | v_51668;
assign v_51671 = v_51557 | v_51670;
assign v_51673 = v_51555 | v_51672;
assign v_51675 = v_51670 | v_51674;
assign v_51677 = v_51554 | v_51676;
assign v_51679 = v_51552 | v_51678;
assign v_51681 = v_51676 | v_51680;
assign v_51683 = v_51551 | v_51682;
assign v_51685 = v_51549 | v_51684;
assign v_51687 = v_51682 | v_51686;
assign v_51689 = v_51548 | v_51688;
assign v_51691 = v_51546 | v_51690;
assign v_51693 = v_51688 | v_51692;
assign v_51696 = ~v_51545 | v_51695;
assign v_51703 = v_51593 | v_51702;
assign v_51706 = v_51704 | v_51705;
assign v_51708 = v_51590 | v_51707;
assign v_51711 = v_51709 | v_51710;
assign v_51713 = v_51587 | v_51712;
assign v_51716 = v_51714 | v_51715;
assign v_51718 = v_51584 | v_51717;
assign v_51721 = v_51719 | v_51720;
assign v_51723 = v_51581 | v_51722;
assign v_51726 = v_51724 | v_51725;
assign v_51728 = v_51578 | v_51727;
assign v_51731 = v_51729 | v_51730;
assign v_51733 = v_51575 | v_51732;
assign v_51736 = v_51734 | v_51735;
assign v_51738 = v_51572 | v_51737;
assign v_51741 = v_51739 | v_51740;
assign v_51743 = v_51569 | v_51742;
assign v_51746 = v_51744 | v_51745;
assign v_51748 = v_51566 | v_51747;
assign v_51751 = v_51749 | v_51750;
assign v_51753 = v_51563 | v_51752;
assign v_51756 = v_51754 | v_51755;
assign v_51758 = v_51560 | v_51757;
assign v_51761 = v_51759 | v_51760;
assign v_51763 = v_51557 | v_51762;
assign v_51766 = v_51764 | v_51765;
assign v_51768 = v_51554 | v_51767;
assign v_51771 = v_51769 | v_51770;
assign v_51773 = v_51551 | v_51772;
assign v_51776 = v_51774 | v_51775;
assign v_51778 = v_51548 | v_51777;
assign v_51781 = v_51779 | v_51780;
assign v_51783 = v_51545 | v_51782;
assign v_51786 = v_51544 | v_51785;
assign v_51840 = v_51837 | v_51839;
assign v_51842 = v_51836 | v_51841;
assign v_51844 = v_51834 | v_51843;
assign v_51846 = v_51841 | v_51845;
assign v_51848 = v_51833 | v_51847;
assign v_51850 = v_51831 | v_51849;
assign v_51852 = v_51847 | v_51851;
assign v_51854 = v_51830 | v_51853;
assign v_51856 = v_51828 | v_51855;
assign v_51858 = v_51853 | v_51857;
assign v_51860 = v_51827 | v_51859;
assign v_51862 = v_51825 | v_51861;
assign v_51864 = v_51859 | v_51863;
assign v_51866 = v_51824 | v_51865;
assign v_51868 = v_51822 | v_51867;
assign v_51870 = v_51865 | v_51869;
assign v_51872 = v_51821 | v_51871;
assign v_51874 = v_51819 | v_51873;
assign v_51876 = v_51871 | v_51875;
assign v_51878 = v_51818 | v_51877;
assign v_51880 = v_51816 | v_51879;
assign v_51882 = v_51877 | v_51881;
assign v_51884 = v_51815 | v_51883;
assign v_51886 = v_51813 | v_51885;
assign v_51888 = v_51883 | v_51887;
assign v_51890 = v_51812 | v_51889;
assign v_51892 = v_51810 | v_51891;
assign v_51894 = v_51889 | v_51893;
assign v_51896 = v_51809 | v_51895;
assign v_51898 = v_51807 | v_51897;
assign v_51900 = v_51895 | v_51899;
assign v_51902 = v_51806 | v_51901;
assign v_51904 = v_51804 | v_51903;
assign v_51906 = v_51901 | v_51905;
assign v_51908 = v_51803 | v_51907;
assign v_51910 = v_51801 | v_51909;
assign v_51912 = v_51907 | v_51911;
assign v_51914 = v_51800 | v_51913;
assign v_51916 = v_51798 | v_51915;
assign v_51918 = v_51913 | v_51917;
assign v_51920 = v_51797 | v_51919;
assign v_51922 = v_51795 | v_51921;
assign v_51924 = v_51919 | v_51923;
assign v_51926 = v_51794 | v_51925;
assign v_51928 = v_51792 | v_51927;
assign v_51930 = v_51925 | v_51929;
assign v_51932 = v_51791 | v_51931;
assign v_51934 = v_51789 | v_51933;
assign v_51936 = v_51931 | v_51935;
assign v_51939 = ~v_51788 | v_51938;
assign v_51946 = v_51836 | v_51945;
assign v_51949 = v_51947 | v_51948;
assign v_51951 = v_51833 | v_51950;
assign v_51954 = v_51952 | v_51953;
assign v_51956 = v_51830 | v_51955;
assign v_51959 = v_51957 | v_51958;
assign v_51961 = v_51827 | v_51960;
assign v_51964 = v_51962 | v_51963;
assign v_51966 = v_51824 | v_51965;
assign v_51969 = v_51967 | v_51968;
assign v_51971 = v_51821 | v_51970;
assign v_51974 = v_51972 | v_51973;
assign v_51976 = v_51818 | v_51975;
assign v_51979 = v_51977 | v_51978;
assign v_51981 = v_51815 | v_51980;
assign v_51984 = v_51982 | v_51983;
assign v_51986 = v_51812 | v_51985;
assign v_51989 = v_51987 | v_51988;
assign v_51991 = v_51809 | v_51990;
assign v_51994 = v_51992 | v_51993;
assign v_51996 = v_51806 | v_51995;
assign v_51999 = v_51997 | v_51998;
assign v_52001 = v_51803 | v_52000;
assign v_52004 = v_52002 | v_52003;
assign v_52006 = v_51800 | v_52005;
assign v_52009 = v_52007 | v_52008;
assign v_52011 = v_51797 | v_52010;
assign v_52014 = v_52012 | v_52013;
assign v_52016 = v_51794 | v_52015;
assign v_52019 = v_52017 | v_52018;
assign v_52021 = v_51791 | v_52020;
assign v_52024 = v_52022 | v_52023;
assign v_52026 = v_51788 | v_52025;
assign v_52029 = v_51787 | v_52028;
assign v_52083 = v_52080 | v_52082;
assign v_52085 = v_52079 | v_52084;
assign v_52087 = v_52077 | v_52086;
assign v_52089 = v_52084 | v_52088;
assign v_52091 = v_52076 | v_52090;
assign v_52093 = v_52074 | v_52092;
assign v_52095 = v_52090 | v_52094;
assign v_52097 = v_52073 | v_52096;
assign v_52099 = v_52071 | v_52098;
assign v_52101 = v_52096 | v_52100;
assign v_52103 = v_52070 | v_52102;
assign v_52105 = v_52068 | v_52104;
assign v_52107 = v_52102 | v_52106;
assign v_52109 = v_52067 | v_52108;
assign v_52111 = v_52065 | v_52110;
assign v_52113 = v_52108 | v_52112;
assign v_52115 = v_52064 | v_52114;
assign v_52117 = v_52062 | v_52116;
assign v_52119 = v_52114 | v_52118;
assign v_52121 = v_52061 | v_52120;
assign v_52123 = v_52059 | v_52122;
assign v_52125 = v_52120 | v_52124;
assign v_52127 = v_52058 | v_52126;
assign v_52129 = v_52056 | v_52128;
assign v_52131 = v_52126 | v_52130;
assign v_52133 = v_52055 | v_52132;
assign v_52135 = v_52053 | v_52134;
assign v_52137 = v_52132 | v_52136;
assign v_52139 = v_52052 | v_52138;
assign v_52141 = v_52050 | v_52140;
assign v_52143 = v_52138 | v_52142;
assign v_52145 = v_52049 | v_52144;
assign v_52147 = v_52047 | v_52146;
assign v_52149 = v_52144 | v_52148;
assign v_52151 = v_52046 | v_52150;
assign v_52153 = v_52044 | v_52152;
assign v_52155 = v_52150 | v_52154;
assign v_52157 = v_52043 | v_52156;
assign v_52159 = v_52041 | v_52158;
assign v_52161 = v_52156 | v_52160;
assign v_52163 = v_52040 | v_52162;
assign v_52165 = v_52038 | v_52164;
assign v_52167 = v_52162 | v_52166;
assign v_52169 = v_52037 | v_52168;
assign v_52171 = v_52035 | v_52170;
assign v_52173 = v_52168 | v_52172;
assign v_52175 = v_52034 | v_52174;
assign v_52177 = v_52032 | v_52176;
assign v_52179 = v_52174 | v_52178;
assign v_52182 = ~v_52031 | v_52181;
assign v_52189 = v_52079 | v_52188;
assign v_52192 = v_52190 | v_52191;
assign v_52194 = v_52076 | v_52193;
assign v_52197 = v_52195 | v_52196;
assign v_52199 = v_52073 | v_52198;
assign v_52202 = v_52200 | v_52201;
assign v_52204 = v_52070 | v_52203;
assign v_52207 = v_52205 | v_52206;
assign v_52209 = v_52067 | v_52208;
assign v_52212 = v_52210 | v_52211;
assign v_52214 = v_52064 | v_52213;
assign v_52217 = v_52215 | v_52216;
assign v_52219 = v_52061 | v_52218;
assign v_52222 = v_52220 | v_52221;
assign v_52224 = v_52058 | v_52223;
assign v_52227 = v_52225 | v_52226;
assign v_52229 = v_52055 | v_52228;
assign v_52232 = v_52230 | v_52231;
assign v_52234 = v_52052 | v_52233;
assign v_52237 = v_52235 | v_52236;
assign v_52239 = v_52049 | v_52238;
assign v_52242 = v_52240 | v_52241;
assign v_52244 = v_52046 | v_52243;
assign v_52247 = v_52245 | v_52246;
assign v_52249 = v_52043 | v_52248;
assign v_52252 = v_52250 | v_52251;
assign v_52254 = v_52040 | v_52253;
assign v_52257 = v_52255 | v_52256;
assign v_52259 = v_52037 | v_52258;
assign v_52262 = v_52260 | v_52261;
assign v_52264 = v_52034 | v_52263;
assign v_52267 = v_52265 | v_52266;
assign v_52269 = v_52031 | v_52268;
assign v_52272 = v_52030 | v_52271;
assign v_52326 = v_52323 | v_52325;
assign v_52328 = v_52322 | v_52327;
assign v_52330 = v_52320 | v_52329;
assign v_52332 = v_52327 | v_52331;
assign v_52334 = v_52319 | v_52333;
assign v_52336 = v_52317 | v_52335;
assign v_52338 = v_52333 | v_52337;
assign v_52340 = v_52316 | v_52339;
assign v_52342 = v_52314 | v_52341;
assign v_52344 = v_52339 | v_52343;
assign v_52346 = v_52313 | v_52345;
assign v_52348 = v_52311 | v_52347;
assign v_52350 = v_52345 | v_52349;
assign v_52352 = v_52310 | v_52351;
assign v_52354 = v_52308 | v_52353;
assign v_52356 = v_52351 | v_52355;
assign v_52358 = v_52307 | v_52357;
assign v_52360 = v_52305 | v_52359;
assign v_52362 = v_52357 | v_52361;
assign v_52364 = v_52304 | v_52363;
assign v_52366 = v_52302 | v_52365;
assign v_52368 = v_52363 | v_52367;
assign v_52370 = v_52301 | v_52369;
assign v_52372 = v_52299 | v_52371;
assign v_52374 = v_52369 | v_52373;
assign v_52376 = v_52298 | v_52375;
assign v_52378 = v_52296 | v_52377;
assign v_52380 = v_52375 | v_52379;
assign v_52382 = v_52295 | v_52381;
assign v_52384 = v_52293 | v_52383;
assign v_52386 = v_52381 | v_52385;
assign v_52388 = v_52292 | v_52387;
assign v_52390 = v_52290 | v_52389;
assign v_52392 = v_52387 | v_52391;
assign v_52394 = v_52289 | v_52393;
assign v_52396 = v_52287 | v_52395;
assign v_52398 = v_52393 | v_52397;
assign v_52400 = v_52286 | v_52399;
assign v_52402 = v_52284 | v_52401;
assign v_52404 = v_52399 | v_52403;
assign v_52406 = v_52283 | v_52405;
assign v_52408 = v_52281 | v_52407;
assign v_52410 = v_52405 | v_52409;
assign v_52412 = v_52280 | v_52411;
assign v_52414 = v_52278 | v_52413;
assign v_52416 = v_52411 | v_52415;
assign v_52418 = v_52277 | v_52417;
assign v_52420 = v_52275 | v_52419;
assign v_52422 = v_52417 | v_52421;
assign v_52425 = ~v_52274 | v_52424;
assign v_52432 = v_52322 | v_52431;
assign v_52435 = v_52433 | v_52434;
assign v_52437 = v_52319 | v_52436;
assign v_52440 = v_52438 | v_52439;
assign v_52442 = v_52316 | v_52441;
assign v_52445 = v_52443 | v_52444;
assign v_52447 = v_52313 | v_52446;
assign v_52450 = v_52448 | v_52449;
assign v_52452 = v_52310 | v_52451;
assign v_52455 = v_52453 | v_52454;
assign v_52457 = v_52307 | v_52456;
assign v_52460 = v_52458 | v_52459;
assign v_52462 = v_52304 | v_52461;
assign v_52465 = v_52463 | v_52464;
assign v_52467 = v_52301 | v_52466;
assign v_52470 = v_52468 | v_52469;
assign v_52472 = v_52298 | v_52471;
assign v_52475 = v_52473 | v_52474;
assign v_52477 = v_52295 | v_52476;
assign v_52480 = v_52478 | v_52479;
assign v_52482 = v_52292 | v_52481;
assign v_52485 = v_52483 | v_52484;
assign v_52487 = v_52289 | v_52486;
assign v_52490 = v_52488 | v_52489;
assign v_52492 = v_52286 | v_52491;
assign v_52495 = v_52493 | v_52494;
assign v_52497 = v_52283 | v_52496;
assign v_52500 = v_52498 | v_52499;
assign v_52502 = v_52280 | v_52501;
assign v_52505 = v_52503 | v_52504;
assign v_52507 = v_52277 | v_52506;
assign v_52510 = v_52508 | v_52509;
assign v_52512 = v_52274 | v_52511;
assign v_52515 = v_52273 | v_52514;
assign v_52569 = v_52566 | v_52568;
assign v_52571 = v_52565 | v_52570;
assign v_52573 = v_52563 | v_52572;
assign v_52575 = v_52570 | v_52574;
assign v_52577 = v_52562 | v_52576;
assign v_52579 = v_52560 | v_52578;
assign v_52581 = v_52576 | v_52580;
assign v_52583 = v_52559 | v_52582;
assign v_52585 = v_52557 | v_52584;
assign v_52587 = v_52582 | v_52586;
assign v_52589 = v_52556 | v_52588;
assign v_52591 = v_52554 | v_52590;
assign v_52593 = v_52588 | v_52592;
assign v_52595 = v_52553 | v_52594;
assign v_52597 = v_52551 | v_52596;
assign v_52599 = v_52594 | v_52598;
assign v_52601 = v_52550 | v_52600;
assign v_52603 = v_52548 | v_52602;
assign v_52605 = v_52600 | v_52604;
assign v_52607 = v_52547 | v_52606;
assign v_52609 = v_52545 | v_52608;
assign v_52611 = v_52606 | v_52610;
assign v_52613 = v_52544 | v_52612;
assign v_52615 = v_52542 | v_52614;
assign v_52617 = v_52612 | v_52616;
assign v_52619 = v_52541 | v_52618;
assign v_52621 = v_52539 | v_52620;
assign v_52623 = v_52618 | v_52622;
assign v_52625 = v_52538 | v_52624;
assign v_52627 = v_52536 | v_52626;
assign v_52629 = v_52624 | v_52628;
assign v_52631 = v_52535 | v_52630;
assign v_52633 = v_52533 | v_52632;
assign v_52635 = v_52630 | v_52634;
assign v_52637 = v_52532 | v_52636;
assign v_52639 = v_52530 | v_52638;
assign v_52641 = v_52636 | v_52640;
assign v_52643 = v_52529 | v_52642;
assign v_52645 = v_52527 | v_52644;
assign v_52647 = v_52642 | v_52646;
assign v_52649 = v_52526 | v_52648;
assign v_52651 = v_52524 | v_52650;
assign v_52653 = v_52648 | v_52652;
assign v_52655 = v_52523 | v_52654;
assign v_52657 = v_52521 | v_52656;
assign v_52659 = v_52654 | v_52658;
assign v_52661 = v_52520 | v_52660;
assign v_52663 = v_52518 | v_52662;
assign v_52665 = v_52660 | v_52664;
assign v_52668 = ~v_52517 | v_52667;
assign v_52675 = v_52565 | v_52674;
assign v_52678 = v_52676 | v_52677;
assign v_52680 = v_52562 | v_52679;
assign v_52683 = v_52681 | v_52682;
assign v_52685 = v_52559 | v_52684;
assign v_52688 = v_52686 | v_52687;
assign v_52690 = v_52556 | v_52689;
assign v_52693 = v_52691 | v_52692;
assign v_52695 = v_52553 | v_52694;
assign v_52698 = v_52696 | v_52697;
assign v_52700 = v_52550 | v_52699;
assign v_52703 = v_52701 | v_52702;
assign v_52705 = v_52547 | v_52704;
assign v_52708 = v_52706 | v_52707;
assign v_52710 = v_52544 | v_52709;
assign v_52713 = v_52711 | v_52712;
assign v_52715 = v_52541 | v_52714;
assign v_52718 = v_52716 | v_52717;
assign v_52720 = v_52538 | v_52719;
assign v_52723 = v_52721 | v_52722;
assign v_52725 = v_52535 | v_52724;
assign v_52728 = v_52726 | v_52727;
assign v_52730 = v_52532 | v_52729;
assign v_52733 = v_52731 | v_52732;
assign v_52735 = v_52529 | v_52734;
assign v_52738 = v_52736 | v_52737;
assign v_52740 = v_52526 | v_52739;
assign v_52743 = v_52741 | v_52742;
assign v_52745 = v_52523 | v_52744;
assign v_52748 = v_52746 | v_52747;
assign v_52750 = v_52520 | v_52749;
assign v_52753 = v_52751 | v_52752;
assign v_52755 = v_52517 | v_52754;
assign v_52758 = v_52516 | v_52757;
assign v_52812 = v_52809 | v_52811;
assign v_52814 = v_52808 | v_52813;
assign v_52816 = v_52806 | v_52815;
assign v_52818 = v_52813 | v_52817;
assign v_52820 = v_52805 | v_52819;
assign v_52822 = v_52803 | v_52821;
assign v_52824 = v_52819 | v_52823;
assign v_52826 = v_52802 | v_52825;
assign v_52828 = v_52800 | v_52827;
assign v_52830 = v_52825 | v_52829;
assign v_52832 = v_52799 | v_52831;
assign v_52834 = v_52797 | v_52833;
assign v_52836 = v_52831 | v_52835;
assign v_52838 = v_52796 | v_52837;
assign v_52840 = v_52794 | v_52839;
assign v_52842 = v_52837 | v_52841;
assign v_52844 = v_52793 | v_52843;
assign v_52846 = v_52791 | v_52845;
assign v_52848 = v_52843 | v_52847;
assign v_52850 = v_52790 | v_52849;
assign v_52852 = v_52788 | v_52851;
assign v_52854 = v_52849 | v_52853;
assign v_52856 = v_52787 | v_52855;
assign v_52858 = v_52785 | v_52857;
assign v_52860 = v_52855 | v_52859;
assign v_52862 = v_52784 | v_52861;
assign v_52864 = v_52782 | v_52863;
assign v_52866 = v_52861 | v_52865;
assign v_52868 = v_52781 | v_52867;
assign v_52870 = v_52779 | v_52869;
assign v_52872 = v_52867 | v_52871;
assign v_52874 = v_52778 | v_52873;
assign v_52876 = v_52776 | v_52875;
assign v_52878 = v_52873 | v_52877;
assign v_52880 = v_52775 | v_52879;
assign v_52882 = v_52773 | v_52881;
assign v_52884 = v_52879 | v_52883;
assign v_52886 = v_52772 | v_52885;
assign v_52888 = v_52770 | v_52887;
assign v_52890 = v_52885 | v_52889;
assign v_52892 = v_52769 | v_52891;
assign v_52894 = v_52767 | v_52893;
assign v_52896 = v_52891 | v_52895;
assign v_52898 = v_52766 | v_52897;
assign v_52900 = v_52764 | v_52899;
assign v_52902 = v_52897 | v_52901;
assign v_52904 = v_52763 | v_52903;
assign v_52906 = v_52761 | v_52905;
assign v_52908 = v_52903 | v_52907;
assign v_52911 = ~v_52760 | v_52910;
assign v_52918 = v_52808 | v_52917;
assign v_52921 = v_52919 | v_52920;
assign v_52923 = v_52805 | v_52922;
assign v_52926 = v_52924 | v_52925;
assign v_52928 = v_52802 | v_52927;
assign v_52931 = v_52929 | v_52930;
assign v_52933 = v_52799 | v_52932;
assign v_52936 = v_52934 | v_52935;
assign v_52938 = v_52796 | v_52937;
assign v_52941 = v_52939 | v_52940;
assign v_52943 = v_52793 | v_52942;
assign v_52946 = v_52944 | v_52945;
assign v_52948 = v_52790 | v_52947;
assign v_52951 = v_52949 | v_52950;
assign v_52953 = v_52787 | v_52952;
assign v_52956 = v_52954 | v_52955;
assign v_52958 = v_52784 | v_52957;
assign v_52961 = v_52959 | v_52960;
assign v_52963 = v_52781 | v_52962;
assign v_52966 = v_52964 | v_52965;
assign v_52968 = v_52778 | v_52967;
assign v_52971 = v_52969 | v_52970;
assign v_52973 = v_52775 | v_52972;
assign v_52976 = v_52974 | v_52975;
assign v_52978 = v_52772 | v_52977;
assign v_52981 = v_52979 | v_52980;
assign v_52983 = v_52769 | v_52982;
assign v_52986 = v_52984 | v_52985;
assign v_52988 = v_52766 | v_52987;
assign v_52991 = v_52989 | v_52990;
assign v_52993 = v_52763 | v_52992;
assign v_52996 = v_52994 | v_52995;
assign v_52998 = v_52760 | v_52997;
assign v_53001 = v_52759 | v_53000;
assign v_53055 = v_53052 | v_53054;
assign v_53057 = v_53051 | v_53056;
assign v_53059 = v_53049 | v_53058;
assign v_53061 = v_53056 | v_53060;
assign v_53063 = v_53048 | v_53062;
assign v_53065 = v_53046 | v_53064;
assign v_53067 = v_53062 | v_53066;
assign v_53069 = v_53045 | v_53068;
assign v_53071 = v_53043 | v_53070;
assign v_53073 = v_53068 | v_53072;
assign v_53075 = v_53042 | v_53074;
assign v_53077 = v_53040 | v_53076;
assign v_53079 = v_53074 | v_53078;
assign v_53081 = v_53039 | v_53080;
assign v_53083 = v_53037 | v_53082;
assign v_53085 = v_53080 | v_53084;
assign v_53087 = v_53036 | v_53086;
assign v_53089 = v_53034 | v_53088;
assign v_53091 = v_53086 | v_53090;
assign v_53093 = v_53033 | v_53092;
assign v_53095 = v_53031 | v_53094;
assign v_53097 = v_53092 | v_53096;
assign v_53099 = v_53030 | v_53098;
assign v_53101 = v_53028 | v_53100;
assign v_53103 = v_53098 | v_53102;
assign v_53105 = v_53027 | v_53104;
assign v_53107 = v_53025 | v_53106;
assign v_53109 = v_53104 | v_53108;
assign v_53111 = v_53024 | v_53110;
assign v_53113 = v_53022 | v_53112;
assign v_53115 = v_53110 | v_53114;
assign v_53117 = v_53021 | v_53116;
assign v_53119 = v_53019 | v_53118;
assign v_53121 = v_53116 | v_53120;
assign v_53123 = v_53018 | v_53122;
assign v_53125 = v_53016 | v_53124;
assign v_53127 = v_53122 | v_53126;
assign v_53129 = v_53015 | v_53128;
assign v_53131 = v_53013 | v_53130;
assign v_53133 = v_53128 | v_53132;
assign v_53135 = v_53012 | v_53134;
assign v_53137 = v_53010 | v_53136;
assign v_53139 = v_53134 | v_53138;
assign v_53141 = v_53009 | v_53140;
assign v_53143 = v_53007 | v_53142;
assign v_53145 = v_53140 | v_53144;
assign v_53147 = v_53006 | v_53146;
assign v_53149 = v_53004 | v_53148;
assign v_53151 = v_53146 | v_53150;
assign v_53154 = ~v_53003 | v_53153;
assign v_53161 = v_53051 | v_53160;
assign v_53164 = v_53162 | v_53163;
assign v_53166 = v_53048 | v_53165;
assign v_53169 = v_53167 | v_53168;
assign v_53171 = v_53045 | v_53170;
assign v_53174 = v_53172 | v_53173;
assign v_53176 = v_53042 | v_53175;
assign v_53179 = v_53177 | v_53178;
assign v_53181 = v_53039 | v_53180;
assign v_53184 = v_53182 | v_53183;
assign v_53186 = v_53036 | v_53185;
assign v_53189 = v_53187 | v_53188;
assign v_53191 = v_53033 | v_53190;
assign v_53194 = v_53192 | v_53193;
assign v_53196 = v_53030 | v_53195;
assign v_53199 = v_53197 | v_53198;
assign v_53201 = v_53027 | v_53200;
assign v_53204 = v_53202 | v_53203;
assign v_53206 = v_53024 | v_53205;
assign v_53209 = v_53207 | v_53208;
assign v_53211 = v_53021 | v_53210;
assign v_53214 = v_53212 | v_53213;
assign v_53216 = v_53018 | v_53215;
assign v_53219 = v_53217 | v_53218;
assign v_53221 = v_53015 | v_53220;
assign v_53224 = v_53222 | v_53223;
assign v_53226 = v_53012 | v_53225;
assign v_53229 = v_53227 | v_53228;
assign v_53231 = v_53009 | v_53230;
assign v_53234 = v_53232 | v_53233;
assign v_53236 = v_53006 | v_53235;
assign v_53239 = v_53237 | v_53238;
assign v_53241 = v_53003 | v_53240;
assign v_53244 = v_53002 | v_53243;
assign v_53298 = v_53295 | v_53297;
assign v_53300 = v_53294 | v_53299;
assign v_53302 = v_53292 | v_53301;
assign v_53304 = v_53299 | v_53303;
assign v_53306 = v_53291 | v_53305;
assign v_53308 = v_53289 | v_53307;
assign v_53310 = v_53305 | v_53309;
assign v_53312 = v_53288 | v_53311;
assign v_53314 = v_53286 | v_53313;
assign v_53316 = v_53311 | v_53315;
assign v_53318 = v_53285 | v_53317;
assign v_53320 = v_53283 | v_53319;
assign v_53322 = v_53317 | v_53321;
assign v_53324 = v_53282 | v_53323;
assign v_53326 = v_53280 | v_53325;
assign v_53328 = v_53323 | v_53327;
assign v_53330 = v_53279 | v_53329;
assign v_53332 = v_53277 | v_53331;
assign v_53334 = v_53329 | v_53333;
assign v_53336 = v_53276 | v_53335;
assign v_53338 = v_53274 | v_53337;
assign v_53340 = v_53335 | v_53339;
assign v_53342 = v_53273 | v_53341;
assign v_53344 = v_53271 | v_53343;
assign v_53346 = v_53341 | v_53345;
assign v_53348 = v_53270 | v_53347;
assign v_53350 = v_53268 | v_53349;
assign v_53352 = v_53347 | v_53351;
assign v_53354 = v_53267 | v_53353;
assign v_53356 = v_53265 | v_53355;
assign v_53358 = v_53353 | v_53357;
assign v_53360 = v_53264 | v_53359;
assign v_53362 = v_53262 | v_53361;
assign v_53364 = v_53359 | v_53363;
assign v_53366 = v_53261 | v_53365;
assign v_53368 = v_53259 | v_53367;
assign v_53370 = v_53365 | v_53369;
assign v_53372 = v_53258 | v_53371;
assign v_53374 = v_53256 | v_53373;
assign v_53376 = v_53371 | v_53375;
assign v_53378 = v_53255 | v_53377;
assign v_53380 = v_53253 | v_53379;
assign v_53382 = v_53377 | v_53381;
assign v_53384 = v_53252 | v_53383;
assign v_53386 = v_53250 | v_53385;
assign v_53388 = v_53383 | v_53387;
assign v_53390 = v_53249 | v_53389;
assign v_53392 = v_53247 | v_53391;
assign v_53394 = v_53389 | v_53393;
assign v_53397 = ~v_53246 | v_53396;
assign v_53404 = v_53294 | v_53403;
assign v_53407 = v_53405 | v_53406;
assign v_53409 = v_53291 | v_53408;
assign v_53412 = v_53410 | v_53411;
assign v_53414 = v_53288 | v_53413;
assign v_53417 = v_53415 | v_53416;
assign v_53419 = v_53285 | v_53418;
assign v_53422 = v_53420 | v_53421;
assign v_53424 = v_53282 | v_53423;
assign v_53427 = v_53425 | v_53426;
assign v_53429 = v_53279 | v_53428;
assign v_53432 = v_53430 | v_53431;
assign v_53434 = v_53276 | v_53433;
assign v_53437 = v_53435 | v_53436;
assign v_53439 = v_53273 | v_53438;
assign v_53442 = v_53440 | v_53441;
assign v_53444 = v_53270 | v_53443;
assign v_53447 = v_53445 | v_53446;
assign v_53449 = v_53267 | v_53448;
assign v_53452 = v_53450 | v_53451;
assign v_53454 = v_53264 | v_53453;
assign v_53457 = v_53455 | v_53456;
assign v_53459 = v_53261 | v_53458;
assign v_53462 = v_53460 | v_53461;
assign v_53464 = v_53258 | v_53463;
assign v_53467 = v_53465 | v_53466;
assign v_53469 = v_53255 | v_53468;
assign v_53472 = v_53470 | v_53471;
assign v_53474 = v_53252 | v_53473;
assign v_53477 = v_53475 | v_53476;
assign v_53479 = v_53249 | v_53478;
assign v_53482 = v_53480 | v_53481;
assign v_53484 = v_53246 | v_53483;
assign v_53487 = v_53245 | v_53486;
assign v_53541 = v_53538 | v_53540;
assign v_53543 = v_53537 | v_53542;
assign v_53545 = v_53535 | v_53544;
assign v_53547 = v_53542 | v_53546;
assign v_53549 = v_53534 | v_53548;
assign v_53551 = v_53532 | v_53550;
assign v_53553 = v_53548 | v_53552;
assign v_53555 = v_53531 | v_53554;
assign v_53557 = v_53529 | v_53556;
assign v_53559 = v_53554 | v_53558;
assign v_53561 = v_53528 | v_53560;
assign v_53563 = v_53526 | v_53562;
assign v_53565 = v_53560 | v_53564;
assign v_53567 = v_53525 | v_53566;
assign v_53569 = v_53523 | v_53568;
assign v_53571 = v_53566 | v_53570;
assign v_53573 = v_53522 | v_53572;
assign v_53575 = v_53520 | v_53574;
assign v_53577 = v_53572 | v_53576;
assign v_53579 = v_53519 | v_53578;
assign v_53581 = v_53517 | v_53580;
assign v_53583 = v_53578 | v_53582;
assign v_53585 = v_53516 | v_53584;
assign v_53587 = v_53514 | v_53586;
assign v_53589 = v_53584 | v_53588;
assign v_53591 = v_53513 | v_53590;
assign v_53593 = v_53511 | v_53592;
assign v_53595 = v_53590 | v_53594;
assign v_53597 = v_53510 | v_53596;
assign v_53599 = v_53508 | v_53598;
assign v_53601 = v_53596 | v_53600;
assign v_53603 = v_53507 | v_53602;
assign v_53605 = v_53505 | v_53604;
assign v_53607 = v_53602 | v_53606;
assign v_53609 = v_53504 | v_53608;
assign v_53611 = v_53502 | v_53610;
assign v_53613 = v_53608 | v_53612;
assign v_53615 = v_53501 | v_53614;
assign v_53617 = v_53499 | v_53616;
assign v_53619 = v_53614 | v_53618;
assign v_53621 = v_53498 | v_53620;
assign v_53623 = v_53496 | v_53622;
assign v_53625 = v_53620 | v_53624;
assign v_53627 = v_53495 | v_53626;
assign v_53629 = v_53493 | v_53628;
assign v_53631 = v_53626 | v_53630;
assign v_53633 = v_53492 | v_53632;
assign v_53635 = v_53490 | v_53634;
assign v_53637 = v_53632 | v_53636;
assign v_53640 = ~v_53489 | v_53639;
assign v_53647 = v_53537 | v_53646;
assign v_53650 = v_53648 | v_53649;
assign v_53652 = v_53534 | v_53651;
assign v_53655 = v_53653 | v_53654;
assign v_53657 = v_53531 | v_53656;
assign v_53660 = v_53658 | v_53659;
assign v_53662 = v_53528 | v_53661;
assign v_53665 = v_53663 | v_53664;
assign v_53667 = v_53525 | v_53666;
assign v_53670 = v_53668 | v_53669;
assign v_53672 = v_53522 | v_53671;
assign v_53675 = v_53673 | v_53674;
assign v_53677 = v_53519 | v_53676;
assign v_53680 = v_53678 | v_53679;
assign v_53682 = v_53516 | v_53681;
assign v_53685 = v_53683 | v_53684;
assign v_53687 = v_53513 | v_53686;
assign v_53690 = v_53688 | v_53689;
assign v_53692 = v_53510 | v_53691;
assign v_53695 = v_53693 | v_53694;
assign v_53697 = v_53507 | v_53696;
assign v_53700 = v_53698 | v_53699;
assign v_53702 = v_53504 | v_53701;
assign v_53705 = v_53703 | v_53704;
assign v_53707 = v_53501 | v_53706;
assign v_53710 = v_53708 | v_53709;
assign v_53712 = v_53498 | v_53711;
assign v_53715 = v_53713 | v_53714;
assign v_53717 = v_53495 | v_53716;
assign v_53720 = v_53718 | v_53719;
assign v_53722 = v_53492 | v_53721;
assign v_53725 = v_53723 | v_53724;
assign v_53727 = v_53489 | v_53726;
assign v_53730 = v_53488 | v_53729;
assign v_53784 = v_53781 | v_53783;
assign v_53786 = v_53780 | v_53785;
assign v_53788 = v_53778 | v_53787;
assign v_53790 = v_53785 | v_53789;
assign v_53792 = v_53777 | v_53791;
assign v_53794 = v_53775 | v_53793;
assign v_53796 = v_53791 | v_53795;
assign v_53798 = v_53774 | v_53797;
assign v_53800 = v_53772 | v_53799;
assign v_53802 = v_53797 | v_53801;
assign v_53804 = v_53771 | v_53803;
assign v_53806 = v_53769 | v_53805;
assign v_53808 = v_53803 | v_53807;
assign v_53810 = v_53768 | v_53809;
assign v_53812 = v_53766 | v_53811;
assign v_53814 = v_53809 | v_53813;
assign v_53816 = v_53765 | v_53815;
assign v_53818 = v_53763 | v_53817;
assign v_53820 = v_53815 | v_53819;
assign v_53822 = v_53762 | v_53821;
assign v_53824 = v_53760 | v_53823;
assign v_53826 = v_53821 | v_53825;
assign v_53828 = v_53759 | v_53827;
assign v_53830 = v_53757 | v_53829;
assign v_53832 = v_53827 | v_53831;
assign v_53834 = v_53756 | v_53833;
assign v_53836 = v_53754 | v_53835;
assign v_53838 = v_53833 | v_53837;
assign v_53840 = v_53753 | v_53839;
assign v_53842 = v_53751 | v_53841;
assign v_53844 = v_53839 | v_53843;
assign v_53846 = v_53750 | v_53845;
assign v_53848 = v_53748 | v_53847;
assign v_53850 = v_53845 | v_53849;
assign v_53852 = v_53747 | v_53851;
assign v_53854 = v_53745 | v_53853;
assign v_53856 = v_53851 | v_53855;
assign v_53858 = v_53744 | v_53857;
assign v_53860 = v_53742 | v_53859;
assign v_53862 = v_53857 | v_53861;
assign v_53864 = v_53741 | v_53863;
assign v_53866 = v_53739 | v_53865;
assign v_53868 = v_53863 | v_53867;
assign v_53870 = v_53738 | v_53869;
assign v_53872 = v_53736 | v_53871;
assign v_53874 = v_53869 | v_53873;
assign v_53876 = v_53735 | v_53875;
assign v_53878 = v_53733 | v_53877;
assign v_53880 = v_53875 | v_53879;
assign v_53883 = ~v_53732 | v_53882;
assign v_53890 = v_53780 | v_53889;
assign v_53893 = v_53891 | v_53892;
assign v_53895 = v_53777 | v_53894;
assign v_53898 = v_53896 | v_53897;
assign v_53900 = v_53774 | v_53899;
assign v_53903 = v_53901 | v_53902;
assign v_53905 = v_53771 | v_53904;
assign v_53908 = v_53906 | v_53907;
assign v_53910 = v_53768 | v_53909;
assign v_53913 = v_53911 | v_53912;
assign v_53915 = v_53765 | v_53914;
assign v_53918 = v_53916 | v_53917;
assign v_53920 = v_53762 | v_53919;
assign v_53923 = v_53921 | v_53922;
assign v_53925 = v_53759 | v_53924;
assign v_53928 = v_53926 | v_53927;
assign v_53930 = v_53756 | v_53929;
assign v_53933 = v_53931 | v_53932;
assign v_53935 = v_53753 | v_53934;
assign v_53938 = v_53936 | v_53937;
assign v_53940 = v_53750 | v_53939;
assign v_53943 = v_53941 | v_53942;
assign v_53945 = v_53747 | v_53944;
assign v_53948 = v_53946 | v_53947;
assign v_53950 = v_53744 | v_53949;
assign v_53953 = v_53951 | v_53952;
assign v_53955 = v_53741 | v_53954;
assign v_53958 = v_53956 | v_53957;
assign v_53960 = v_53738 | v_53959;
assign v_53963 = v_53961 | v_53962;
assign v_53965 = v_53735 | v_53964;
assign v_53968 = v_53966 | v_53967;
assign v_53970 = v_53732 | v_53969;
assign v_53973 = v_53731 | v_53972;
assign v_54026 = v_54023 | v_54025;
assign v_54028 = v_54022 | v_54027;
assign v_54030 = v_54020 | v_54029;
assign v_54032 = v_54027 | v_54031;
assign v_54034 = v_54019 | v_54033;
assign v_54036 = v_54017 | v_54035;
assign v_54038 = v_54033 | v_54037;
assign v_54040 = v_54016 | v_54039;
assign v_54042 = v_54014 | v_54041;
assign v_54044 = v_54039 | v_54043;
assign v_54046 = v_54013 | v_54045;
assign v_54048 = v_54011 | v_54047;
assign v_54050 = v_54045 | v_54049;
assign v_54052 = v_54010 | v_54051;
assign v_54054 = v_54008 | v_54053;
assign v_54056 = v_54051 | v_54055;
assign v_54058 = v_54007 | v_54057;
assign v_54060 = v_54005 | v_54059;
assign v_54062 = v_54057 | v_54061;
assign v_54064 = v_54004 | v_54063;
assign v_54066 = v_54002 | v_54065;
assign v_54068 = v_54063 | v_54067;
assign v_54070 = v_54001 | v_54069;
assign v_54072 = v_53999 | v_54071;
assign v_54074 = v_54069 | v_54073;
assign v_54076 = v_53998 | v_54075;
assign v_54078 = v_53996 | v_54077;
assign v_54080 = v_54075 | v_54079;
assign v_54082 = v_53995 | v_54081;
assign v_54084 = v_53993 | v_54083;
assign v_54086 = v_54081 | v_54085;
assign v_54088 = v_53992 | v_54087;
assign v_54090 = v_53990 | v_54089;
assign v_54092 = v_54087 | v_54091;
assign v_54094 = v_53989 | v_54093;
assign v_54096 = v_53987 | v_54095;
assign v_54098 = v_54093 | v_54097;
assign v_54100 = v_53986 | v_54099;
assign v_54102 = v_53984 | v_54101;
assign v_54104 = v_54099 | v_54103;
assign v_54106 = v_53983 | v_54105;
assign v_54108 = v_53981 | v_54107;
assign v_54110 = v_54105 | v_54109;
assign v_54112 = v_53980 | v_54111;
assign v_54114 = v_53978 | v_54113;
assign v_54116 = v_54111 | v_54115;
assign v_54118 = v_53977 | v_54117;
assign v_54120 = v_53975 | v_54119;
assign v_54122 = v_54117 | v_54121;
assign v_54126 = v_54123 | v_54125;
assign v_54133 = v_54022 | v_54132;
assign v_54136 = v_54134 | v_54135;
assign v_54138 = v_54019 | v_54137;
assign v_54141 = v_54139 | v_54140;
assign v_54143 = v_54016 | v_54142;
assign v_54146 = v_54144 | v_54145;
assign v_54148 = v_54013 | v_54147;
assign v_54151 = v_54149 | v_54150;
assign v_54153 = v_54010 | v_54152;
assign v_54156 = v_54154 | v_54155;
assign v_54158 = v_54007 | v_54157;
assign v_54161 = v_54159 | v_54160;
assign v_54163 = v_54004 | v_54162;
assign v_54166 = v_54164 | v_54165;
assign v_54168 = v_54001 | v_54167;
assign v_54171 = v_54169 | v_54170;
assign v_54173 = v_53998 | v_54172;
assign v_54176 = v_54174 | v_54175;
assign v_54178 = v_53995 | v_54177;
assign v_54181 = v_54179 | v_54180;
assign v_54183 = v_53992 | v_54182;
assign v_54186 = v_54184 | v_54185;
assign v_54188 = v_53989 | v_54187;
assign v_54191 = v_54189 | v_54190;
assign v_54193 = v_53986 | v_54192;
assign v_54196 = v_54194 | v_54195;
assign v_54198 = v_53983 | v_54197;
assign v_54201 = v_54199 | v_54200;
assign v_54203 = v_53980 | v_54202;
assign v_54206 = v_54204 | v_54205;
assign v_54208 = v_53977 | v_54207;
assign v_54211 = v_54209 | v_54210;
assign v_54213 = v_54211 | v_54212;
assign v_54216 = v_53974 | v_54215;
assign v_54287 = v_54284 | v_54286;
assign v_54289 = v_54282 | v_54288;
assign v_54291 = v_54280 | v_54290;
assign v_54293 = v_54288 | v_54292;
assign v_54295 = v_54278 | v_54294;
assign v_54297 = v_54276 | v_54296;
assign v_54299 = v_54294 | v_54298;
assign v_54301 = v_54274 | v_54300;
assign v_54303 = v_54272 | v_54302;
assign v_54305 = v_54300 | v_54304;
assign v_54307 = v_54270 | v_54306;
assign v_54309 = v_54268 | v_54308;
assign v_54311 = v_54306 | v_54310;
assign v_54313 = v_54266 | v_54312;
assign v_54315 = v_54264 | v_54314;
assign v_54317 = v_54312 | v_54316;
assign v_54319 = v_54262 | v_54318;
assign v_54321 = v_54260 | v_54320;
assign v_54323 = v_54318 | v_54322;
assign v_54325 = v_54258 | v_54324;
assign v_54327 = v_54256 | v_54326;
assign v_54329 = v_54324 | v_54328;
assign v_54331 = v_54254 | v_54330;
assign v_54333 = v_54252 | v_54332;
assign v_54335 = v_54330 | v_54334;
assign v_54337 = v_54250 | v_54336;
assign v_54339 = v_54248 | v_54338;
assign v_54341 = v_54336 | v_54340;
assign v_54343 = v_54246 | v_54342;
assign v_54345 = v_54244 | v_54344;
assign v_54347 = v_54342 | v_54346;
assign v_54349 = v_54242 | v_54348;
assign v_54351 = v_54240 | v_54350;
assign v_54353 = v_54348 | v_54352;
assign v_54355 = v_54238 | v_54354;
assign v_54357 = v_54236 | v_54356;
assign v_54359 = v_54354 | v_54358;
assign v_54361 = v_54234 | v_54360;
assign v_54363 = v_54231 | v_54362;
assign v_54365 = v_54360 | v_54364;
assign v_54367 = v_54230 | v_54366;
assign v_54369 = v_54227 | v_54368;
assign v_54371 = v_54366 | v_54370;
assign v_54373 = v_54226 | v_54372;
assign v_54375 = v_54223 | v_54374;
assign v_54377 = v_54372 | v_54376;
assign v_54379 = v_54222 | v_54378;
assign v_54381 = v_54219 | v_54380;
assign v_54383 = v_54378 | v_54382;
assign v_54386 = ~v_54218 | v_54385;
assign v_54393 = v_54282 | v_54392;
assign v_54396 = v_54394 | v_54395;
assign v_54398 = v_54278 | v_54397;
assign v_54401 = v_54399 | v_54400;
assign v_54403 = v_54274 | v_54402;
assign v_54406 = v_54404 | v_54405;
assign v_54408 = v_54270 | v_54407;
assign v_54411 = v_54409 | v_54410;
assign v_54413 = v_54266 | v_54412;
assign v_54416 = v_54414 | v_54415;
assign v_54418 = v_54262 | v_54417;
assign v_54421 = v_54419 | v_54420;
assign v_54423 = v_54258 | v_54422;
assign v_54426 = v_54424 | v_54425;
assign v_54428 = v_54254 | v_54427;
assign v_54431 = v_54429 | v_54430;
assign v_54433 = v_54250 | v_54432;
assign v_54436 = v_54434 | v_54435;
assign v_54438 = v_54246 | v_54437;
assign v_54441 = v_54439 | v_54440;
assign v_54443 = v_54242 | v_54442;
assign v_54446 = v_54444 | v_54445;
assign v_54448 = v_54238 | v_54447;
assign v_54451 = v_54449 | v_54450;
assign v_54453 = v_54234 | v_54452;
assign v_54456 = v_54454 | v_54455;
assign v_54458 = v_54230 | v_54457;
assign v_54461 = v_54459 | v_54460;
assign v_54463 = v_54226 | v_54462;
assign v_54466 = v_54464 | v_54465;
assign v_54468 = v_54222 | v_54467;
assign v_54471 = v_54469 | v_54470;
assign v_54473 = v_54218 | v_54472;
assign v_54476 = v_54217 | v_54475;
assign v_54530 = v_54527 | v_54529;
assign v_54532 = v_54526 | v_54531;
assign v_54534 = v_54524 | v_54533;
assign v_54536 = v_54531 | v_54535;
assign v_54538 = v_54523 | v_54537;
assign v_54540 = v_54521 | v_54539;
assign v_54542 = v_54537 | v_54541;
assign v_54544 = v_54520 | v_54543;
assign v_54546 = v_54518 | v_54545;
assign v_54548 = v_54543 | v_54547;
assign v_54550 = v_54517 | v_54549;
assign v_54552 = v_54515 | v_54551;
assign v_54554 = v_54549 | v_54553;
assign v_54556 = v_54514 | v_54555;
assign v_54558 = v_54512 | v_54557;
assign v_54560 = v_54555 | v_54559;
assign v_54562 = v_54511 | v_54561;
assign v_54564 = v_54509 | v_54563;
assign v_54566 = v_54561 | v_54565;
assign v_54568 = v_54508 | v_54567;
assign v_54570 = v_54506 | v_54569;
assign v_54572 = v_54567 | v_54571;
assign v_54574 = v_54505 | v_54573;
assign v_54576 = v_54503 | v_54575;
assign v_54578 = v_54573 | v_54577;
assign v_54580 = v_54502 | v_54579;
assign v_54582 = v_54500 | v_54581;
assign v_54584 = v_54579 | v_54583;
assign v_54586 = v_54499 | v_54585;
assign v_54588 = v_54497 | v_54587;
assign v_54590 = v_54585 | v_54589;
assign v_54592 = v_54496 | v_54591;
assign v_54594 = v_54494 | v_54593;
assign v_54596 = v_54591 | v_54595;
assign v_54598 = v_54493 | v_54597;
assign v_54600 = v_54491 | v_54599;
assign v_54602 = v_54597 | v_54601;
assign v_54604 = v_54490 | v_54603;
assign v_54606 = v_54488 | v_54605;
assign v_54608 = v_54603 | v_54607;
assign v_54610 = v_54487 | v_54609;
assign v_54612 = v_54485 | v_54611;
assign v_54614 = v_54609 | v_54613;
assign v_54616 = v_54484 | v_54615;
assign v_54618 = v_54482 | v_54617;
assign v_54620 = v_54615 | v_54619;
assign v_54622 = v_54481 | v_54621;
assign v_54624 = v_54479 | v_54623;
assign v_54626 = v_54621 | v_54625;
assign v_54629 = ~v_54478 | v_54628;
assign v_54636 = v_54526 | v_54635;
assign v_54639 = v_54637 | v_54638;
assign v_54641 = v_54523 | v_54640;
assign v_54644 = v_54642 | v_54643;
assign v_54646 = v_54520 | v_54645;
assign v_54649 = v_54647 | v_54648;
assign v_54651 = v_54517 | v_54650;
assign v_54654 = v_54652 | v_54653;
assign v_54656 = v_54514 | v_54655;
assign v_54659 = v_54657 | v_54658;
assign v_54661 = v_54511 | v_54660;
assign v_54664 = v_54662 | v_54663;
assign v_54666 = v_54508 | v_54665;
assign v_54669 = v_54667 | v_54668;
assign v_54671 = v_54505 | v_54670;
assign v_54674 = v_54672 | v_54673;
assign v_54676 = v_54502 | v_54675;
assign v_54679 = v_54677 | v_54678;
assign v_54681 = v_54499 | v_54680;
assign v_54684 = v_54682 | v_54683;
assign v_54686 = v_54496 | v_54685;
assign v_54689 = v_54687 | v_54688;
assign v_54691 = v_54493 | v_54690;
assign v_54694 = v_54692 | v_54693;
assign v_54696 = v_54490 | v_54695;
assign v_54699 = v_54697 | v_54698;
assign v_54701 = v_54487 | v_54700;
assign v_54704 = v_54702 | v_54703;
assign v_54706 = v_54484 | v_54705;
assign v_54709 = v_54707 | v_54708;
assign v_54711 = v_54481 | v_54710;
assign v_54714 = v_54712 | v_54713;
assign v_54716 = v_54478 | v_54715;
assign v_54719 = v_54477 | v_54718;
assign v_54773 = v_54770 | v_54772;
assign v_54775 = v_54769 | v_54774;
assign v_54777 = v_54767 | v_54776;
assign v_54779 = v_54774 | v_54778;
assign v_54781 = v_54766 | v_54780;
assign v_54783 = v_54764 | v_54782;
assign v_54785 = v_54780 | v_54784;
assign v_54787 = v_54763 | v_54786;
assign v_54789 = v_54761 | v_54788;
assign v_54791 = v_54786 | v_54790;
assign v_54793 = v_54760 | v_54792;
assign v_54795 = v_54758 | v_54794;
assign v_54797 = v_54792 | v_54796;
assign v_54799 = v_54757 | v_54798;
assign v_54801 = v_54755 | v_54800;
assign v_54803 = v_54798 | v_54802;
assign v_54805 = v_54754 | v_54804;
assign v_54807 = v_54752 | v_54806;
assign v_54809 = v_54804 | v_54808;
assign v_54811 = v_54751 | v_54810;
assign v_54813 = v_54749 | v_54812;
assign v_54815 = v_54810 | v_54814;
assign v_54817 = v_54748 | v_54816;
assign v_54819 = v_54746 | v_54818;
assign v_54821 = v_54816 | v_54820;
assign v_54823 = v_54745 | v_54822;
assign v_54825 = v_54743 | v_54824;
assign v_54827 = v_54822 | v_54826;
assign v_54829 = v_54742 | v_54828;
assign v_54831 = v_54740 | v_54830;
assign v_54833 = v_54828 | v_54832;
assign v_54835 = v_54739 | v_54834;
assign v_54837 = v_54737 | v_54836;
assign v_54839 = v_54834 | v_54838;
assign v_54841 = v_54736 | v_54840;
assign v_54843 = v_54734 | v_54842;
assign v_54845 = v_54840 | v_54844;
assign v_54847 = v_54733 | v_54846;
assign v_54849 = v_54731 | v_54848;
assign v_54851 = v_54846 | v_54850;
assign v_54853 = v_54730 | v_54852;
assign v_54855 = v_54728 | v_54854;
assign v_54857 = v_54852 | v_54856;
assign v_54859 = v_54727 | v_54858;
assign v_54861 = v_54725 | v_54860;
assign v_54863 = v_54858 | v_54862;
assign v_54865 = v_54724 | v_54864;
assign v_54867 = v_54722 | v_54866;
assign v_54869 = v_54864 | v_54868;
assign v_54872 = ~v_54721 | v_54871;
assign v_54879 = v_54769 | v_54878;
assign v_54882 = v_54880 | v_54881;
assign v_54884 = v_54766 | v_54883;
assign v_54887 = v_54885 | v_54886;
assign v_54889 = v_54763 | v_54888;
assign v_54892 = v_54890 | v_54891;
assign v_54894 = v_54760 | v_54893;
assign v_54897 = v_54895 | v_54896;
assign v_54899 = v_54757 | v_54898;
assign v_54902 = v_54900 | v_54901;
assign v_54904 = v_54754 | v_54903;
assign v_54907 = v_54905 | v_54906;
assign v_54909 = v_54751 | v_54908;
assign v_54912 = v_54910 | v_54911;
assign v_54914 = v_54748 | v_54913;
assign v_54917 = v_54915 | v_54916;
assign v_54919 = v_54745 | v_54918;
assign v_54922 = v_54920 | v_54921;
assign v_54924 = v_54742 | v_54923;
assign v_54927 = v_54925 | v_54926;
assign v_54929 = v_54739 | v_54928;
assign v_54932 = v_54930 | v_54931;
assign v_54934 = v_54736 | v_54933;
assign v_54937 = v_54935 | v_54936;
assign v_54939 = v_54733 | v_54938;
assign v_54942 = v_54940 | v_54941;
assign v_54944 = v_54730 | v_54943;
assign v_54947 = v_54945 | v_54946;
assign v_54949 = v_54727 | v_54948;
assign v_54952 = v_54950 | v_54951;
assign v_54954 = v_54724 | v_54953;
assign v_54957 = v_54955 | v_54956;
assign v_54959 = v_54721 | v_54958;
assign v_54962 = v_54720 | v_54961;
assign v_55016 = v_55013 | v_55015;
assign v_55018 = v_55012 | v_55017;
assign v_55020 = v_55010 | v_55019;
assign v_55022 = v_55017 | v_55021;
assign v_55024 = v_55009 | v_55023;
assign v_55026 = v_55007 | v_55025;
assign v_55028 = v_55023 | v_55027;
assign v_55030 = v_55006 | v_55029;
assign v_55032 = v_55004 | v_55031;
assign v_55034 = v_55029 | v_55033;
assign v_55036 = v_55003 | v_55035;
assign v_55038 = v_55001 | v_55037;
assign v_55040 = v_55035 | v_55039;
assign v_55042 = v_55000 | v_55041;
assign v_55044 = v_54998 | v_55043;
assign v_55046 = v_55041 | v_55045;
assign v_55048 = v_54997 | v_55047;
assign v_55050 = v_54995 | v_55049;
assign v_55052 = v_55047 | v_55051;
assign v_55054 = v_54994 | v_55053;
assign v_55056 = v_54992 | v_55055;
assign v_55058 = v_55053 | v_55057;
assign v_55060 = v_54991 | v_55059;
assign v_55062 = v_54989 | v_55061;
assign v_55064 = v_55059 | v_55063;
assign v_55066 = v_54988 | v_55065;
assign v_55068 = v_54986 | v_55067;
assign v_55070 = v_55065 | v_55069;
assign v_55072 = v_54985 | v_55071;
assign v_55074 = v_54983 | v_55073;
assign v_55076 = v_55071 | v_55075;
assign v_55078 = v_54982 | v_55077;
assign v_55080 = v_54980 | v_55079;
assign v_55082 = v_55077 | v_55081;
assign v_55084 = v_54979 | v_55083;
assign v_55086 = v_54977 | v_55085;
assign v_55088 = v_55083 | v_55087;
assign v_55090 = v_54976 | v_55089;
assign v_55092 = v_54974 | v_55091;
assign v_55094 = v_55089 | v_55093;
assign v_55096 = v_54973 | v_55095;
assign v_55098 = v_54971 | v_55097;
assign v_55100 = v_55095 | v_55099;
assign v_55102 = v_54970 | v_55101;
assign v_55104 = v_54968 | v_55103;
assign v_55106 = v_55101 | v_55105;
assign v_55108 = v_54967 | v_55107;
assign v_55110 = v_54965 | v_55109;
assign v_55112 = v_55107 | v_55111;
assign v_55115 = ~v_54964 | v_55114;
assign v_55122 = v_55012 | v_55121;
assign v_55125 = v_55123 | v_55124;
assign v_55127 = v_55009 | v_55126;
assign v_55130 = v_55128 | v_55129;
assign v_55132 = v_55006 | v_55131;
assign v_55135 = v_55133 | v_55134;
assign v_55137 = v_55003 | v_55136;
assign v_55140 = v_55138 | v_55139;
assign v_55142 = v_55000 | v_55141;
assign v_55145 = v_55143 | v_55144;
assign v_55147 = v_54997 | v_55146;
assign v_55150 = v_55148 | v_55149;
assign v_55152 = v_54994 | v_55151;
assign v_55155 = v_55153 | v_55154;
assign v_55157 = v_54991 | v_55156;
assign v_55160 = v_55158 | v_55159;
assign v_55162 = v_54988 | v_55161;
assign v_55165 = v_55163 | v_55164;
assign v_55167 = v_54985 | v_55166;
assign v_55170 = v_55168 | v_55169;
assign v_55172 = v_54982 | v_55171;
assign v_55175 = v_55173 | v_55174;
assign v_55177 = v_54979 | v_55176;
assign v_55180 = v_55178 | v_55179;
assign v_55182 = v_54976 | v_55181;
assign v_55185 = v_55183 | v_55184;
assign v_55187 = v_54973 | v_55186;
assign v_55190 = v_55188 | v_55189;
assign v_55192 = v_54970 | v_55191;
assign v_55195 = v_55193 | v_55194;
assign v_55197 = v_54967 | v_55196;
assign v_55200 = v_55198 | v_55199;
assign v_55202 = v_54964 | v_55201;
assign v_55205 = v_54963 | v_55204;
assign v_55259 = v_55256 | v_55258;
assign v_55261 = v_55255 | v_55260;
assign v_55263 = v_55253 | v_55262;
assign v_55265 = v_55260 | v_55264;
assign v_55267 = v_55252 | v_55266;
assign v_55269 = v_55250 | v_55268;
assign v_55271 = v_55266 | v_55270;
assign v_55273 = v_55249 | v_55272;
assign v_55275 = v_55247 | v_55274;
assign v_55277 = v_55272 | v_55276;
assign v_55279 = v_55246 | v_55278;
assign v_55281 = v_55244 | v_55280;
assign v_55283 = v_55278 | v_55282;
assign v_55285 = v_55243 | v_55284;
assign v_55287 = v_55241 | v_55286;
assign v_55289 = v_55284 | v_55288;
assign v_55291 = v_55240 | v_55290;
assign v_55293 = v_55238 | v_55292;
assign v_55295 = v_55290 | v_55294;
assign v_55297 = v_55237 | v_55296;
assign v_55299 = v_55235 | v_55298;
assign v_55301 = v_55296 | v_55300;
assign v_55303 = v_55234 | v_55302;
assign v_55305 = v_55232 | v_55304;
assign v_55307 = v_55302 | v_55306;
assign v_55309 = v_55231 | v_55308;
assign v_55311 = v_55229 | v_55310;
assign v_55313 = v_55308 | v_55312;
assign v_55315 = v_55228 | v_55314;
assign v_55317 = v_55226 | v_55316;
assign v_55319 = v_55314 | v_55318;
assign v_55321 = v_55225 | v_55320;
assign v_55323 = v_55223 | v_55322;
assign v_55325 = v_55320 | v_55324;
assign v_55327 = v_55222 | v_55326;
assign v_55329 = v_55220 | v_55328;
assign v_55331 = v_55326 | v_55330;
assign v_55333 = v_55219 | v_55332;
assign v_55335 = v_55217 | v_55334;
assign v_55337 = v_55332 | v_55336;
assign v_55339 = v_55216 | v_55338;
assign v_55341 = v_55214 | v_55340;
assign v_55343 = v_55338 | v_55342;
assign v_55345 = v_55213 | v_55344;
assign v_55347 = v_55211 | v_55346;
assign v_55349 = v_55344 | v_55348;
assign v_55351 = v_55210 | v_55350;
assign v_55353 = v_55208 | v_55352;
assign v_55355 = v_55350 | v_55354;
assign v_55358 = ~v_55207 | v_55357;
assign v_55365 = v_55255 | v_55364;
assign v_55368 = v_55366 | v_55367;
assign v_55370 = v_55252 | v_55369;
assign v_55373 = v_55371 | v_55372;
assign v_55375 = v_55249 | v_55374;
assign v_55378 = v_55376 | v_55377;
assign v_55380 = v_55246 | v_55379;
assign v_55383 = v_55381 | v_55382;
assign v_55385 = v_55243 | v_55384;
assign v_55388 = v_55386 | v_55387;
assign v_55390 = v_55240 | v_55389;
assign v_55393 = v_55391 | v_55392;
assign v_55395 = v_55237 | v_55394;
assign v_55398 = v_55396 | v_55397;
assign v_55400 = v_55234 | v_55399;
assign v_55403 = v_55401 | v_55402;
assign v_55405 = v_55231 | v_55404;
assign v_55408 = v_55406 | v_55407;
assign v_55410 = v_55228 | v_55409;
assign v_55413 = v_55411 | v_55412;
assign v_55415 = v_55225 | v_55414;
assign v_55418 = v_55416 | v_55417;
assign v_55420 = v_55222 | v_55419;
assign v_55423 = v_55421 | v_55422;
assign v_55425 = v_55219 | v_55424;
assign v_55428 = v_55426 | v_55427;
assign v_55430 = v_55216 | v_55429;
assign v_55433 = v_55431 | v_55432;
assign v_55435 = v_55213 | v_55434;
assign v_55438 = v_55436 | v_55437;
assign v_55440 = v_55210 | v_55439;
assign v_55443 = v_55441 | v_55442;
assign v_55445 = v_55207 | v_55444;
assign v_55448 = v_55206 | v_55447;
assign v_55502 = v_55499 | v_55501;
assign v_55504 = v_55498 | v_55503;
assign v_55506 = v_55496 | v_55505;
assign v_55508 = v_55503 | v_55507;
assign v_55510 = v_55495 | v_55509;
assign v_55512 = v_55493 | v_55511;
assign v_55514 = v_55509 | v_55513;
assign v_55516 = v_55492 | v_55515;
assign v_55518 = v_55490 | v_55517;
assign v_55520 = v_55515 | v_55519;
assign v_55522 = v_55489 | v_55521;
assign v_55524 = v_55487 | v_55523;
assign v_55526 = v_55521 | v_55525;
assign v_55528 = v_55486 | v_55527;
assign v_55530 = v_55484 | v_55529;
assign v_55532 = v_55527 | v_55531;
assign v_55534 = v_55483 | v_55533;
assign v_55536 = v_55481 | v_55535;
assign v_55538 = v_55533 | v_55537;
assign v_55540 = v_55480 | v_55539;
assign v_55542 = v_55478 | v_55541;
assign v_55544 = v_55539 | v_55543;
assign v_55546 = v_55477 | v_55545;
assign v_55548 = v_55475 | v_55547;
assign v_55550 = v_55545 | v_55549;
assign v_55552 = v_55474 | v_55551;
assign v_55554 = v_55472 | v_55553;
assign v_55556 = v_55551 | v_55555;
assign v_55558 = v_55471 | v_55557;
assign v_55560 = v_55469 | v_55559;
assign v_55562 = v_55557 | v_55561;
assign v_55564 = v_55468 | v_55563;
assign v_55566 = v_55466 | v_55565;
assign v_55568 = v_55563 | v_55567;
assign v_55570 = v_55465 | v_55569;
assign v_55572 = v_55463 | v_55571;
assign v_55574 = v_55569 | v_55573;
assign v_55576 = v_55462 | v_55575;
assign v_55578 = v_55460 | v_55577;
assign v_55580 = v_55575 | v_55579;
assign v_55582 = v_55459 | v_55581;
assign v_55584 = v_55457 | v_55583;
assign v_55586 = v_55581 | v_55585;
assign v_55588 = v_55456 | v_55587;
assign v_55590 = v_55454 | v_55589;
assign v_55592 = v_55587 | v_55591;
assign v_55594 = v_55453 | v_55593;
assign v_55596 = v_55451 | v_55595;
assign v_55598 = v_55593 | v_55597;
assign v_55601 = ~v_55450 | v_55600;
assign v_55608 = v_55498 | v_55607;
assign v_55611 = v_55609 | v_55610;
assign v_55613 = v_55495 | v_55612;
assign v_55616 = v_55614 | v_55615;
assign v_55618 = v_55492 | v_55617;
assign v_55621 = v_55619 | v_55620;
assign v_55623 = v_55489 | v_55622;
assign v_55626 = v_55624 | v_55625;
assign v_55628 = v_55486 | v_55627;
assign v_55631 = v_55629 | v_55630;
assign v_55633 = v_55483 | v_55632;
assign v_55636 = v_55634 | v_55635;
assign v_55638 = v_55480 | v_55637;
assign v_55641 = v_55639 | v_55640;
assign v_55643 = v_55477 | v_55642;
assign v_55646 = v_55644 | v_55645;
assign v_55648 = v_55474 | v_55647;
assign v_55651 = v_55649 | v_55650;
assign v_55653 = v_55471 | v_55652;
assign v_55656 = v_55654 | v_55655;
assign v_55658 = v_55468 | v_55657;
assign v_55661 = v_55659 | v_55660;
assign v_55663 = v_55465 | v_55662;
assign v_55666 = v_55664 | v_55665;
assign v_55668 = v_55462 | v_55667;
assign v_55671 = v_55669 | v_55670;
assign v_55673 = v_55459 | v_55672;
assign v_55676 = v_55674 | v_55675;
assign v_55678 = v_55456 | v_55677;
assign v_55681 = v_55679 | v_55680;
assign v_55683 = v_55453 | v_55682;
assign v_55686 = v_55684 | v_55685;
assign v_55688 = v_55450 | v_55687;
assign v_55691 = v_55449 | v_55690;
assign v_55745 = v_55742 | v_55744;
assign v_55747 = v_55741 | v_55746;
assign v_55749 = v_55739 | v_55748;
assign v_55751 = v_55746 | v_55750;
assign v_55753 = v_55738 | v_55752;
assign v_55755 = v_55736 | v_55754;
assign v_55757 = v_55752 | v_55756;
assign v_55759 = v_55735 | v_55758;
assign v_55761 = v_55733 | v_55760;
assign v_55763 = v_55758 | v_55762;
assign v_55765 = v_55732 | v_55764;
assign v_55767 = v_55730 | v_55766;
assign v_55769 = v_55764 | v_55768;
assign v_55771 = v_55729 | v_55770;
assign v_55773 = v_55727 | v_55772;
assign v_55775 = v_55770 | v_55774;
assign v_55777 = v_55726 | v_55776;
assign v_55779 = v_55724 | v_55778;
assign v_55781 = v_55776 | v_55780;
assign v_55783 = v_55723 | v_55782;
assign v_55785 = v_55721 | v_55784;
assign v_55787 = v_55782 | v_55786;
assign v_55789 = v_55720 | v_55788;
assign v_55791 = v_55718 | v_55790;
assign v_55793 = v_55788 | v_55792;
assign v_55795 = v_55717 | v_55794;
assign v_55797 = v_55715 | v_55796;
assign v_55799 = v_55794 | v_55798;
assign v_55801 = v_55714 | v_55800;
assign v_55803 = v_55712 | v_55802;
assign v_55805 = v_55800 | v_55804;
assign v_55807 = v_55711 | v_55806;
assign v_55809 = v_55709 | v_55808;
assign v_55811 = v_55806 | v_55810;
assign v_55813 = v_55708 | v_55812;
assign v_55815 = v_55706 | v_55814;
assign v_55817 = v_55812 | v_55816;
assign v_55819 = v_55705 | v_55818;
assign v_55821 = v_55703 | v_55820;
assign v_55823 = v_55818 | v_55822;
assign v_55825 = v_55702 | v_55824;
assign v_55827 = v_55700 | v_55826;
assign v_55829 = v_55824 | v_55828;
assign v_55831 = v_55699 | v_55830;
assign v_55833 = v_55697 | v_55832;
assign v_55835 = v_55830 | v_55834;
assign v_55837 = v_55696 | v_55836;
assign v_55839 = v_55694 | v_55838;
assign v_55841 = v_55836 | v_55840;
assign v_55844 = ~v_55693 | v_55843;
assign v_55851 = v_55741 | v_55850;
assign v_55854 = v_55852 | v_55853;
assign v_55856 = v_55738 | v_55855;
assign v_55859 = v_55857 | v_55858;
assign v_55861 = v_55735 | v_55860;
assign v_55864 = v_55862 | v_55863;
assign v_55866 = v_55732 | v_55865;
assign v_55869 = v_55867 | v_55868;
assign v_55871 = v_55729 | v_55870;
assign v_55874 = v_55872 | v_55873;
assign v_55876 = v_55726 | v_55875;
assign v_55879 = v_55877 | v_55878;
assign v_55881 = v_55723 | v_55880;
assign v_55884 = v_55882 | v_55883;
assign v_55886 = v_55720 | v_55885;
assign v_55889 = v_55887 | v_55888;
assign v_55891 = v_55717 | v_55890;
assign v_55894 = v_55892 | v_55893;
assign v_55896 = v_55714 | v_55895;
assign v_55899 = v_55897 | v_55898;
assign v_55901 = v_55711 | v_55900;
assign v_55904 = v_55902 | v_55903;
assign v_55906 = v_55708 | v_55905;
assign v_55909 = v_55907 | v_55908;
assign v_55911 = v_55705 | v_55910;
assign v_55914 = v_55912 | v_55913;
assign v_55916 = v_55702 | v_55915;
assign v_55919 = v_55917 | v_55918;
assign v_55921 = v_55699 | v_55920;
assign v_55924 = v_55922 | v_55923;
assign v_55926 = v_55696 | v_55925;
assign v_55929 = v_55927 | v_55928;
assign v_55931 = v_55693 | v_55930;
assign v_55934 = v_55692 | v_55933;
assign v_55988 = v_55985 | v_55987;
assign v_55990 = v_55984 | v_55989;
assign v_55992 = v_55982 | v_55991;
assign v_55994 = v_55989 | v_55993;
assign v_55996 = v_55981 | v_55995;
assign v_55998 = v_55979 | v_55997;
assign v_56000 = v_55995 | v_55999;
assign v_56002 = v_55978 | v_56001;
assign v_56004 = v_55976 | v_56003;
assign v_56006 = v_56001 | v_56005;
assign v_56008 = v_55975 | v_56007;
assign v_56010 = v_55973 | v_56009;
assign v_56012 = v_56007 | v_56011;
assign v_56014 = v_55972 | v_56013;
assign v_56016 = v_55970 | v_56015;
assign v_56018 = v_56013 | v_56017;
assign v_56020 = v_55969 | v_56019;
assign v_56022 = v_55967 | v_56021;
assign v_56024 = v_56019 | v_56023;
assign v_56026 = v_55966 | v_56025;
assign v_56028 = v_55964 | v_56027;
assign v_56030 = v_56025 | v_56029;
assign v_56032 = v_55963 | v_56031;
assign v_56034 = v_55961 | v_56033;
assign v_56036 = v_56031 | v_56035;
assign v_56038 = v_55960 | v_56037;
assign v_56040 = v_55958 | v_56039;
assign v_56042 = v_56037 | v_56041;
assign v_56044 = v_55957 | v_56043;
assign v_56046 = v_55955 | v_56045;
assign v_56048 = v_56043 | v_56047;
assign v_56050 = v_55954 | v_56049;
assign v_56052 = v_55952 | v_56051;
assign v_56054 = v_56049 | v_56053;
assign v_56056 = v_55951 | v_56055;
assign v_56058 = v_55949 | v_56057;
assign v_56060 = v_56055 | v_56059;
assign v_56062 = v_55948 | v_56061;
assign v_56064 = v_55946 | v_56063;
assign v_56066 = v_56061 | v_56065;
assign v_56068 = v_55945 | v_56067;
assign v_56070 = v_55943 | v_56069;
assign v_56072 = v_56067 | v_56071;
assign v_56074 = v_55942 | v_56073;
assign v_56076 = v_55940 | v_56075;
assign v_56078 = v_56073 | v_56077;
assign v_56080 = v_55939 | v_56079;
assign v_56082 = v_55937 | v_56081;
assign v_56084 = v_56079 | v_56083;
assign v_56087 = ~v_55936 | v_56086;
assign v_56094 = v_55984 | v_56093;
assign v_56097 = v_56095 | v_56096;
assign v_56099 = v_55981 | v_56098;
assign v_56102 = v_56100 | v_56101;
assign v_56104 = v_55978 | v_56103;
assign v_56107 = v_56105 | v_56106;
assign v_56109 = v_55975 | v_56108;
assign v_56112 = v_56110 | v_56111;
assign v_56114 = v_55972 | v_56113;
assign v_56117 = v_56115 | v_56116;
assign v_56119 = v_55969 | v_56118;
assign v_56122 = v_56120 | v_56121;
assign v_56124 = v_55966 | v_56123;
assign v_56127 = v_56125 | v_56126;
assign v_56129 = v_55963 | v_56128;
assign v_56132 = v_56130 | v_56131;
assign v_56134 = v_55960 | v_56133;
assign v_56137 = v_56135 | v_56136;
assign v_56139 = v_55957 | v_56138;
assign v_56142 = v_56140 | v_56141;
assign v_56144 = v_55954 | v_56143;
assign v_56147 = v_56145 | v_56146;
assign v_56149 = v_55951 | v_56148;
assign v_56152 = v_56150 | v_56151;
assign v_56154 = v_55948 | v_56153;
assign v_56157 = v_56155 | v_56156;
assign v_56159 = v_55945 | v_56158;
assign v_56162 = v_56160 | v_56161;
assign v_56164 = v_55942 | v_56163;
assign v_56167 = v_56165 | v_56166;
assign v_56169 = v_55939 | v_56168;
assign v_56172 = v_56170 | v_56171;
assign v_56174 = v_55936 | v_56173;
assign v_56177 = v_55935 | v_56176;
assign v_56231 = v_56228 | v_56230;
assign v_56233 = v_56227 | v_56232;
assign v_56235 = v_56225 | v_56234;
assign v_56237 = v_56232 | v_56236;
assign v_56239 = v_56224 | v_56238;
assign v_56241 = v_56222 | v_56240;
assign v_56243 = v_56238 | v_56242;
assign v_56245 = v_56221 | v_56244;
assign v_56247 = v_56219 | v_56246;
assign v_56249 = v_56244 | v_56248;
assign v_56251 = v_56218 | v_56250;
assign v_56253 = v_56216 | v_56252;
assign v_56255 = v_56250 | v_56254;
assign v_56257 = v_56215 | v_56256;
assign v_56259 = v_56213 | v_56258;
assign v_56261 = v_56256 | v_56260;
assign v_56263 = v_56212 | v_56262;
assign v_56265 = v_56210 | v_56264;
assign v_56267 = v_56262 | v_56266;
assign v_56269 = v_56209 | v_56268;
assign v_56271 = v_56207 | v_56270;
assign v_56273 = v_56268 | v_56272;
assign v_56275 = v_56206 | v_56274;
assign v_56277 = v_56204 | v_56276;
assign v_56279 = v_56274 | v_56278;
assign v_56281 = v_56203 | v_56280;
assign v_56283 = v_56201 | v_56282;
assign v_56285 = v_56280 | v_56284;
assign v_56287 = v_56200 | v_56286;
assign v_56289 = v_56198 | v_56288;
assign v_56291 = v_56286 | v_56290;
assign v_56293 = v_56197 | v_56292;
assign v_56295 = v_56195 | v_56294;
assign v_56297 = v_56292 | v_56296;
assign v_56299 = v_56194 | v_56298;
assign v_56301 = v_56192 | v_56300;
assign v_56303 = v_56298 | v_56302;
assign v_56305 = v_56191 | v_56304;
assign v_56307 = v_56189 | v_56306;
assign v_56309 = v_56304 | v_56308;
assign v_56311 = v_56188 | v_56310;
assign v_56313 = v_56186 | v_56312;
assign v_56315 = v_56310 | v_56314;
assign v_56317 = v_56185 | v_56316;
assign v_56319 = v_56183 | v_56318;
assign v_56321 = v_56316 | v_56320;
assign v_56323 = v_56182 | v_56322;
assign v_56325 = v_56180 | v_56324;
assign v_56327 = v_56322 | v_56326;
assign v_56330 = ~v_56179 | v_56329;
assign v_56337 = v_56227 | v_56336;
assign v_56340 = v_56338 | v_56339;
assign v_56342 = v_56224 | v_56341;
assign v_56345 = v_56343 | v_56344;
assign v_56347 = v_56221 | v_56346;
assign v_56350 = v_56348 | v_56349;
assign v_56352 = v_56218 | v_56351;
assign v_56355 = v_56353 | v_56354;
assign v_56357 = v_56215 | v_56356;
assign v_56360 = v_56358 | v_56359;
assign v_56362 = v_56212 | v_56361;
assign v_56365 = v_56363 | v_56364;
assign v_56367 = v_56209 | v_56366;
assign v_56370 = v_56368 | v_56369;
assign v_56372 = v_56206 | v_56371;
assign v_56375 = v_56373 | v_56374;
assign v_56377 = v_56203 | v_56376;
assign v_56380 = v_56378 | v_56379;
assign v_56382 = v_56200 | v_56381;
assign v_56385 = v_56383 | v_56384;
assign v_56387 = v_56197 | v_56386;
assign v_56390 = v_56388 | v_56389;
assign v_56392 = v_56194 | v_56391;
assign v_56395 = v_56393 | v_56394;
assign v_56397 = v_56191 | v_56396;
assign v_56400 = v_56398 | v_56399;
assign v_56402 = v_56188 | v_56401;
assign v_56405 = v_56403 | v_56404;
assign v_56407 = v_56185 | v_56406;
assign v_56410 = v_56408 | v_56409;
assign v_56412 = v_56182 | v_56411;
assign v_56415 = v_56413 | v_56414;
assign v_56417 = v_56179 | v_56416;
assign v_56420 = v_56178 | v_56419;
assign v_56474 = v_56471 | v_56473;
assign v_56476 = v_56470 | v_56475;
assign v_56478 = v_56468 | v_56477;
assign v_56480 = v_56475 | v_56479;
assign v_56482 = v_56467 | v_56481;
assign v_56484 = v_56465 | v_56483;
assign v_56486 = v_56481 | v_56485;
assign v_56488 = v_56464 | v_56487;
assign v_56490 = v_56462 | v_56489;
assign v_56492 = v_56487 | v_56491;
assign v_56494 = v_56461 | v_56493;
assign v_56496 = v_56459 | v_56495;
assign v_56498 = v_56493 | v_56497;
assign v_56500 = v_56458 | v_56499;
assign v_56502 = v_56456 | v_56501;
assign v_56504 = v_56499 | v_56503;
assign v_56506 = v_56455 | v_56505;
assign v_56508 = v_56453 | v_56507;
assign v_56510 = v_56505 | v_56509;
assign v_56512 = v_56452 | v_56511;
assign v_56514 = v_56450 | v_56513;
assign v_56516 = v_56511 | v_56515;
assign v_56518 = v_56449 | v_56517;
assign v_56520 = v_56447 | v_56519;
assign v_56522 = v_56517 | v_56521;
assign v_56524 = v_56446 | v_56523;
assign v_56526 = v_56444 | v_56525;
assign v_56528 = v_56523 | v_56527;
assign v_56530 = v_56443 | v_56529;
assign v_56532 = v_56441 | v_56531;
assign v_56534 = v_56529 | v_56533;
assign v_56536 = v_56440 | v_56535;
assign v_56538 = v_56438 | v_56537;
assign v_56540 = v_56535 | v_56539;
assign v_56542 = v_56437 | v_56541;
assign v_56544 = v_56435 | v_56543;
assign v_56546 = v_56541 | v_56545;
assign v_56548 = v_56434 | v_56547;
assign v_56550 = v_56432 | v_56549;
assign v_56552 = v_56547 | v_56551;
assign v_56554 = v_56431 | v_56553;
assign v_56556 = v_56429 | v_56555;
assign v_56558 = v_56553 | v_56557;
assign v_56560 = v_56428 | v_56559;
assign v_56562 = v_56426 | v_56561;
assign v_56564 = v_56559 | v_56563;
assign v_56566 = v_56425 | v_56565;
assign v_56568 = v_56423 | v_56567;
assign v_56570 = v_56565 | v_56569;
assign v_56573 = ~v_56422 | v_56572;
assign v_56580 = v_56470 | v_56579;
assign v_56583 = v_56581 | v_56582;
assign v_56585 = v_56467 | v_56584;
assign v_56588 = v_56586 | v_56587;
assign v_56590 = v_56464 | v_56589;
assign v_56593 = v_56591 | v_56592;
assign v_56595 = v_56461 | v_56594;
assign v_56598 = v_56596 | v_56597;
assign v_56600 = v_56458 | v_56599;
assign v_56603 = v_56601 | v_56602;
assign v_56605 = v_56455 | v_56604;
assign v_56608 = v_56606 | v_56607;
assign v_56610 = v_56452 | v_56609;
assign v_56613 = v_56611 | v_56612;
assign v_56615 = v_56449 | v_56614;
assign v_56618 = v_56616 | v_56617;
assign v_56620 = v_56446 | v_56619;
assign v_56623 = v_56621 | v_56622;
assign v_56625 = v_56443 | v_56624;
assign v_56628 = v_56626 | v_56627;
assign v_56630 = v_56440 | v_56629;
assign v_56633 = v_56631 | v_56632;
assign v_56635 = v_56437 | v_56634;
assign v_56638 = v_56636 | v_56637;
assign v_56640 = v_56434 | v_56639;
assign v_56643 = v_56641 | v_56642;
assign v_56645 = v_56431 | v_56644;
assign v_56648 = v_56646 | v_56647;
assign v_56650 = v_56428 | v_56649;
assign v_56653 = v_56651 | v_56652;
assign v_56655 = v_56425 | v_56654;
assign v_56658 = v_56656 | v_56657;
assign v_56660 = v_56422 | v_56659;
assign v_56663 = v_56421 | v_56662;
assign v_56717 = v_56714 | v_56716;
assign v_56719 = v_56713 | v_56718;
assign v_56721 = v_56711 | v_56720;
assign v_56723 = v_56718 | v_56722;
assign v_56725 = v_56710 | v_56724;
assign v_56727 = v_56708 | v_56726;
assign v_56729 = v_56724 | v_56728;
assign v_56731 = v_56707 | v_56730;
assign v_56733 = v_56705 | v_56732;
assign v_56735 = v_56730 | v_56734;
assign v_56737 = v_56704 | v_56736;
assign v_56739 = v_56702 | v_56738;
assign v_56741 = v_56736 | v_56740;
assign v_56743 = v_56701 | v_56742;
assign v_56745 = v_56699 | v_56744;
assign v_56747 = v_56742 | v_56746;
assign v_56749 = v_56698 | v_56748;
assign v_56751 = v_56696 | v_56750;
assign v_56753 = v_56748 | v_56752;
assign v_56755 = v_56695 | v_56754;
assign v_56757 = v_56693 | v_56756;
assign v_56759 = v_56754 | v_56758;
assign v_56761 = v_56692 | v_56760;
assign v_56763 = v_56690 | v_56762;
assign v_56765 = v_56760 | v_56764;
assign v_56767 = v_56689 | v_56766;
assign v_56769 = v_56687 | v_56768;
assign v_56771 = v_56766 | v_56770;
assign v_56773 = v_56686 | v_56772;
assign v_56775 = v_56684 | v_56774;
assign v_56777 = v_56772 | v_56776;
assign v_56779 = v_56683 | v_56778;
assign v_56781 = v_56681 | v_56780;
assign v_56783 = v_56778 | v_56782;
assign v_56785 = v_56680 | v_56784;
assign v_56787 = v_56678 | v_56786;
assign v_56789 = v_56784 | v_56788;
assign v_56791 = v_56677 | v_56790;
assign v_56793 = v_56675 | v_56792;
assign v_56795 = v_56790 | v_56794;
assign v_56797 = v_56674 | v_56796;
assign v_56799 = v_56672 | v_56798;
assign v_56801 = v_56796 | v_56800;
assign v_56803 = v_56671 | v_56802;
assign v_56805 = v_56669 | v_56804;
assign v_56807 = v_56802 | v_56806;
assign v_56809 = v_56668 | v_56808;
assign v_56811 = v_56666 | v_56810;
assign v_56813 = v_56808 | v_56812;
assign v_56816 = ~v_56665 | v_56815;
assign v_56823 = v_56713 | v_56822;
assign v_56826 = v_56824 | v_56825;
assign v_56828 = v_56710 | v_56827;
assign v_56831 = v_56829 | v_56830;
assign v_56833 = v_56707 | v_56832;
assign v_56836 = v_56834 | v_56835;
assign v_56838 = v_56704 | v_56837;
assign v_56841 = v_56839 | v_56840;
assign v_56843 = v_56701 | v_56842;
assign v_56846 = v_56844 | v_56845;
assign v_56848 = v_56698 | v_56847;
assign v_56851 = v_56849 | v_56850;
assign v_56853 = v_56695 | v_56852;
assign v_56856 = v_56854 | v_56855;
assign v_56858 = v_56692 | v_56857;
assign v_56861 = v_56859 | v_56860;
assign v_56863 = v_56689 | v_56862;
assign v_56866 = v_56864 | v_56865;
assign v_56868 = v_56686 | v_56867;
assign v_56871 = v_56869 | v_56870;
assign v_56873 = v_56683 | v_56872;
assign v_56876 = v_56874 | v_56875;
assign v_56878 = v_56680 | v_56877;
assign v_56881 = v_56879 | v_56880;
assign v_56883 = v_56677 | v_56882;
assign v_56886 = v_56884 | v_56885;
assign v_56888 = v_56674 | v_56887;
assign v_56891 = v_56889 | v_56890;
assign v_56893 = v_56671 | v_56892;
assign v_56896 = v_56894 | v_56895;
assign v_56898 = v_56668 | v_56897;
assign v_56901 = v_56899 | v_56900;
assign v_56903 = v_56665 | v_56902;
assign v_56906 = v_56664 | v_56905;
assign v_56960 = v_56957 | v_56959;
assign v_56962 = v_56956 | v_56961;
assign v_56964 = v_56954 | v_56963;
assign v_56966 = v_56961 | v_56965;
assign v_56968 = v_56953 | v_56967;
assign v_56970 = v_56951 | v_56969;
assign v_56972 = v_56967 | v_56971;
assign v_56974 = v_56950 | v_56973;
assign v_56976 = v_56948 | v_56975;
assign v_56978 = v_56973 | v_56977;
assign v_56980 = v_56947 | v_56979;
assign v_56982 = v_56945 | v_56981;
assign v_56984 = v_56979 | v_56983;
assign v_56986 = v_56944 | v_56985;
assign v_56988 = v_56942 | v_56987;
assign v_56990 = v_56985 | v_56989;
assign v_56992 = v_56941 | v_56991;
assign v_56994 = v_56939 | v_56993;
assign v_56996 = v_56991 | v_56995;
assign v_56998 = v_56938 | v_56997;
assign v_57000 = v_56936 | v_56999;
assign v_57002 = v_56997 | v_57001;
assign v_57004 = v_56935 | v_57003;
assign v_57006 = v_56933 | v_57005;
assign v_57008 = v_57003 | v_57007;
assign v_57010 = v_56932 | v_57009;
assign v_57012 = v_56930 | v_57011;
assign v_57014 = v_57009 | v_57013;
assign v_57016 = v_56929 | v_57015;
assign v_57018 = v_56927 | v_57017;
assign v_57020 = v_57015 | v_57019;
assign v_57022 = v_56926 | v_57021;
assign v_57024 = v_56924 | v_57023;
assign v_57026 = v_57021 | v_57025;
assign v_57028 = v_56923 | v_57027;
assign v_57030 = v_56921 | v_57029;
assign v_57032 = v_57027 | v_57031;
assign v_57034 = v_56920 | v_57033;
assign v_57036 = v_56918 | v_57035;
assign v_57038 = v_57033 | v_57037;
assign v_57040 = v_56917 | v_57039;
assign v_57042 = v_56915 | v_57041;
assign v_57044 = v_57039 | v_57043;
assign v_57046 = v_56914 | v_57045;
assign v_57048 = v_56912 | v_57047;
assign v_57050 = v_57045 | v_57049;
assign v_57052 = v_56911 | v_57051;
assign v_57054 = v_56909 | v_57053;
assign v_57056 = v_57051 | v_57055;
assign v_57059 = ~v_56908 | v_57058;
assign v_57066 = v_56956 | v_57065;
assign v_57069 = v_57067 | v_57068;
assign v_57071 = v_56953 | v_57070;
assign v_57074 = v_57072 | v_57073;
assign v_57076 = v_56950 | v_57075;
assign v_57079 = v_57077 | v_57078;
assign v_57081 = v_56947 | v_57080;
assign v_57084 = v_57082 | v_57083;
assign v_57086 = v_56944 | v_57085;
assign v_57089 = v_57087 | v_57088;
assign v_57091 = v_56941 | v_57090;
assign v_57094 = v_57092 | v_57093;
assign v_57096 = v_56938 | v_57095;
assign v_57099 = v_57097 | v_57098;
assign v_57101 = v_56935 | v_57100;
assign v_57104 = v_57102 | v_57103;
assign v_57106 = v_56932 | v_57105;
assign v_57109 = v_57107 | v_57108;
assign v_57111 = v_56929 | v_57110;
assign v_57114 = v_57112 | v_57113;
assign v_57116 = v_56926 | v_57115;
assign v_57119 = v_57117 | v_57118;
assign v_57121 = v_56923 | v_57120;
assign v_57124 = v_57122 | v_57123;
assign v_57126 = v_56920 | v_57125;
assign v_57129 = v_57127 | v_57128;
assign v_57131 = v_56917 | v_57130;
assign v_57134 = v_57132 | v_57133;
assign v_57136 = v_56914 | v_57135;
assign v_57139 = v_57137 | v_57138;
assign v_57141 = v_56911 | v_57140;
assign v_57144 = v_57142 | v_57143;
assign v_57146 = v_56908 | v_57145;
assign v_57149 = v_56907 | v_57148;
assign v_57203 = v_57200 | v_57202;
assign v_57205 = v_57199 | v_57204;
assign v_57207 = v_57197 | v_57206;
assign v_57209 = v_57204 | v_57208;
assign v_57211 = v_57196 | v_57210;
assign v_57213 = v_57194 | v_57212;
assign v_57215 = v_57210 | v_57214;
assign v_57217 = v_57193 | v_57216;
assign v_57219 = v_57191 | v_57218;
assign v_57221 = v_57216 | v_57220;
assign v_57223 = v_57190 | v_57222;
assign v_57225 = v_57188 | v_57224;
assign v_57227 = v_57222 | v_57226;
assign v_57229 = v_57187 | v_57228;
assign v_57231 = v_57185 | v_57230;
assign v_57233 = v_57228 | v_57232;
assign v_57235 = v_57184 | v_57234;
assign v_57237 = v_57182 | v_57236;
assign v_57239 = v_57234 | v_57238;
assign v_57241 = v_57181 | v_57240;
assign v_57243 = v_57179 | v_57242;
assign v_57245 = v_57240 | v_57244;
assign v_57247 = v_57178 | v_57246;
assign v_57249 = v_57176 | v_57248;
assign v_57251 = v_57246 | v_57250;
assign v_57253 = v_57175 | v_57252;
assign v_57255 = v_57173 | v_57254;
assign v_57257 = v_57252 | v_57256;
assign v_57259 = v_57172 | v_57258;
assign v_57261 = v_57170 | v_57260;
assign v_57263 = v_57258 | v_57262;
assign v_57265 = v_57169 | v_57264;
assign v_57267 = v_57167 | v_57266;
assign v_57269 = v_57264 | v_57268;
assign v_57271 = v_57166 | v_57270;
assign v_57273 = v_57164 | v_57272;
assign v_57275 = v_57270 | v_57274;
assign v_57277 = v_57163 | v_57276;
assign v_57279 = v_57161 | v_57278;
assign v_57281 = v_57276 | v_57280;
assign v_57283 = v_57160 | v_57282;
assign v_57285 = v_57158 | v_57284;
assign v_57287 = v_57282 | v_57286;
assign v_57289 = v_57157 | v_57288;
assign v_57291 = v_57155 | v_57290;
assign v_57293 = v_57288 | v_57292;
assign v_57295 = v_57154 | v_57294;
assign v_57297 = v_57152 | v_57296;
assign v_57299 = v_57294 | v_57298;
assign v_57302 = ~v_57151 | v_57301;
assign v_57309 = v_57199 | v_57308;
assign v_57312 = v_57310 | v_57311;
assign v_57314 = v_57196 | v_57313;
assign v_57317 = v_57315 | v_57316;
assign v_57319 = v_57193 | v_57318;
assign v_57322 = v_57320 | v_57321;
assign v_57324 = v_57190 | v_57323;
assign v_57327 = v_57325 | v_57326;
assign v_57329 = v_57187 | v_57328;
assign v_57332 = v_57330 | v_57331;
assign v_57334 = v_57184 | v_57333;
assign v_57337 = v_57335 | v_57336;
assign v_57339 = v_57181 | v_57338;
assign v_57342 = v_57340 | v_57341;
assign v_57344 = v_57178 | v_57343;
assign v_57347 = v_57345 | v_57346;
assign v_57349 = v_57175 | v_57348;
assign v_57352 = v_57350 | v_57351;
assign v_57354 = v_57172 | v_57353;
assign v_57357 = v_57355 | v_57356;
assign v_57359 = v_57169 | v_57358;
assign v_57362 = v_57360 | v_57361;
assign v_57364 = v_57166 | v_57363;
assign v_57367 = v_57365 | v_57366;
assign v_57369 = v_57163 | v_57368;
assign v_57372 = v_57370 | v_57371;
assign v_57374 = v_57160 | v_57373;
assign v_57377 = v_57375 | v_57376;
assign v_57379 = v_57157 | v_57378;
assign v_57382 = v_57380 | v_57381;
assign v_57384 = v_57154 | v_57383;
assign v_57387 = v_57385 | v_57386;
assign v_57389 = v_57151 | v_57388;
assign v_57392 = v_57150 | v_57391;
assign v_57446 = v_57443 | v_57445;
assign v_57448 = v_57442 | v_57447;
assign v_57450 = v_57440 | v_57449;
assign v_57452 = v_57447 | v_57451;
assign v_57454 = v_57439 | v_57453;
assign v_57456 = v_57437 | v_57455;
assign v_57458 = v_57453 | v_57457;
assign v_57460 = v_57436 | v_57459;
assign v_57462 = v_57434 | v_57461;
assign v_57464 = v_57459 | v_57463;
assign v_57466 = v_57433 | v_57465;
assign v_57468 = v_57431 | v_57467;
assign v_57470 = v_57465 | v_57469;
assign v_57472 = v_57430 | v_57471;
assign v_57474 = v_57428 | v_57473;
assign v_57476 = v_57471 | v_57475;
assign v_57478 = v_57427 | v_57477;
assign v_57480 = v_57425 | v_57479;
assign v_57482 = v_57477 | v_57481;
assign v_57484 = v_57424 | v_57483;
assign v_57486 = v_57422 | v_57485;
assign v_57488 = v_57483 | v_57487;
assign v_57490 = v_57421 | v_57489;
assign v_57492 = v_57419 | v_57491;
assign v_57494 = v_57489 | v_57493;
assign v_57496 = v_57418 | v_57495;
assign v_57498 = v_57416 | v_57497;
assign v_57500 = v_57495 | v_57499;
assign v_57502 = v_57415 | v_57501;
assign v_57504 = v_57413 | v_57503;
assign v_57506 = v_57501 | v_57505;
assign v_57508 = v_57412 | v_57507;
assign v_57510 = v_57410 | v_57509;
assign v_57512 = v_57507 | v_57511;
assign v_57514 = v_57409 | v_57513;
assign v_57516 = v_57407 | v_57515;
assign v_57518 = v_57513 | v_57517;
assign v_57520 = v_57406 | v_57519;
assign v_57522 = v_57404 | v_57521;
assign v_57524 = v_57519 | v_57523;
assign v_57526 = v_57403 | v_57525;
assign v_57528 = v_57401 | v_57527;
assign v_57530 = v_57525 | v_57529;
assign v_57532 = v_57400 | v_57531;
assign v_57534 = v_57398 | v_57533;
assign v_57536 = v_57531 | v_57535;
assign v_57538 = v_57397 | v_57537;
assign v_57540 = v_57395 | v_57539;
assign v_57542 = v_57537 | v_57541;
assign v_57545 = ~v_57394 | v_57544;
assign v_57552 = v_57442 | v_57551;
assign v_57555 = v_57553 | v_57554;
assign v_57557 = v_57439 | v_57556;
assign v_57560 = v_57558 | v_57559;
assign v_57562 = v_57436 | v_57561;
assign v_57565 = v_57563 | v_57564;
assign v_57567 = v_57433 | v_57566;
assign v_57570 = v_57568 | v_57569;
assign v_57572 = v_57430 | v_57571;
assign v_57575 = v_57573 | v_57574;
assign v_57577 = v_57427 | v_57576;
assign v_57580 = v_57578 | v_57579;
assign v_57582 = v_57424 | v_57581;
assign v_57585 = v_57583 | v_57584;
assign v_57587 = v_57421 | v_57586;
assign v_57590 = v_57588 | v_57589;
assign v_57592 = v_57418 | v_57591;
assign v_57595 = v_57593 | v_57594;
assign v_57597 = v_57415 | v_57596;
assign v_57600 = v_57598 | v_57599;
assign v_57602 = v_57412 | v_57601;
assign v_57605 = v_57603 | v_57604;
assign v_57607 = v_57409 | v_57606;
assign v_57610 = v_57608 | v_57609;
assign v_57612 = v_57406 | v_57611;
assign v_57615 = v_57613 | v_57614;
assign v_57617 = v_57403 | v_57616;
assign v_57620 = v_57618 | v_57619;
assign v_57622 = v_57400 | v_57621;
assign v_57625 = v_57623 | v_57624;
assign v_57627 = v_57397 | v_57626;
assign v_57630 = v_57628 | v_57629;
assign v_57632 = v_57394 | v_57631;
assign v_57635 = v_57393 | v_57634;
assign v_57689 = v_57686 | v_57688;
assign v_57691 = v_57685 | v_57690;
assign v_57693 = v_57683 | v_57692;
assign v_57695 = v_57690 | v_57694;
assign v_57697 = v_57682 | v_57696;
assign v_57699 = v_57680 | v_57698;
assign v_57701 = v_57696 | v_57700;
assign v_57703 = v_57679 | v_57702;
assign v_57705 = v_57677 | v_57704;
assign v_57707 = v_57702 | v_57706;
assign v_57709 = v_57676 | v_57708;
assign v_57711 = v_57674 | v_57710;
assign v_57713 = v_57708 | v_57712;
assign v_57715 = v_57673 | v_57714;
assign v_57717 = v_57671 | v_57716;
assign v_57719 = v_57714 | v_57718;
assign v_57721 = v_57670 | v_57720;
assign v_57723 = v_57668 | v_57722;
assign v_57725 = v_57720 | v_57724;
assign v_57727 = v_57667 | v_57726;
assign v_57729 = v_57665 | v_57728;
assign v_57731 = v_57726 | v_57730;
assign v_57733 = v_57664 | v_57732;
assign v_57735 = v_57662 | v_57734;
assign v_57737 = v_57732 | v_57736;
assign v_57739 = v_57661 | v_57738;
assign v_57741 = v_57659 | v_57740;
assign v_57743 = v_57738 | v_57742;
assign v_57745 = v_57658 | v_57744;
assign v_57747 = v_57656 | v_57746;
assign v_57749 = v_57744 | v_57748;
assign v_57751 = v_57655 | v_57750;
assign v_57753 = v_57653 | v_57752;
assign v_57755 = v_57750 | v_57754;
assign v_57757 = v_57652 | v_57756;
assign v_57759 = v_57650 | v_57758;
assign v_57761 = v_57756 | v_57760;
assign v_57763 = v_57649 | v_57762;
assign v_57765 = v_57647 | v_57764;
assign v_57767 = v_57762 | v_57766;
assign v_57769 = v_57646 | v_57768;
assign v_57771 = v_57644 | v_57770;
assign v_57773 = v_57768 | v_57772;
assign v_57775 = v_57643 | v_57774;
assign v_57777 = v_57641 | v_57776;
assign v_57779 = v_57774 | v_57778;
assign v_57781 = v_57640 | v_57780;
assign v_57783 = v_57638 | v_57782;
assign v_57785 = v_57780 | v_57784;
assign v_57788 = ~v_57637 | v_57787;
assign v_57795 = v_57685 | v_57794;
assign v_57798 = v_57796 | v_57797;
assign v_57800 = v_57682 | v_57799;
assign v_57803 = v_57801 | v_57802;
assign v_57805 = v_57679 | v_57804;
assign v_57808 = v_57806 | v_57807;
assign v_57810 = v_57676 | v_57809;
assign v_57813 = v_57811 | v_57812;
assign v_57815 = v_57673 | v_57814;
assign v_57818 = v_57816 | v_57817;
assign v_57820 = v_57670 | v_57819;
assign v_57823 = v_57821 | v_57822;
assign v_57825 = v_57667 | v_57824;
assign v_57828 = v_57826 | v_57827;
assign v_57830 = v_57664 | v_57829;
assign v_57833 = v_57831 | v_57832;
assign v_57835 = v_57661 | v_57834;
assign v_57838 = v_57836 | v_57837;
assign v_57840 = v_57658 | v_57839;
assign v_57843 = v_57841 | v_57842;
assign v_57845 = v_57655 | v_57844;
assign v_57848 = v_57846 | v_57847;
assign v_57850 = v_57652 | v_57849;
assign v_57853 = v_57851 | v_57852;
assign v_57855 = v_57649 | v_57854;
assign v_57858 = v_57856 | v_57857;
assign v_57860 = v_57646 | v_57859;
assign v_57863 = v_57861 | v_57862;
assign v_57865 = v_57643 | v_57864;
assign v_57868 = v_57866 | v_57867;
assign v_57870 = v_57640 | v_57869;
assign v_57873 = v_57871 | v_57872;
assign v_57875 = v_57637 | v_57874;
assign v_57878 = v_57636 | v_57877;
assign v_57932 = v_57929 | v_57931;
assign v_57934 = v_57928 | v_57933;
assign v_57936 = v_57926 | v_57935;
assign v_57938 = v_57933 | v_57937;
assign v_57940 = v_57925 | v_57939;
assign v_57942 = v_57923 | v_57941;
assign v_57944 = v_57939 | v_57943;
assign v_57946 = v_57922 | v_57945;
assign v_57948 = v_57920 | v_57947;
assign v_57950 = v_57945 | v_57949;
assign v_57952 = v_57919 | v_57951;
assign v_57954 = v_57917 | v_57953;
assign v_57956 = v_57951 | v_57955;
assign v_57958 = v_57916 | v_57957;
assign v_57960 = v_57914 | v_57959;
assign v_57962 = v_57957 | v_57961;
assign v_57964 = v_57913 | v_57963;
assign v_57966 = v_57911 | v_57965;
assign v_57968 = v_57963 | v_57967;
assign v_57970 = v_57910 | v_57969;
assign v_57972 = v_57908 | v_57971;
assign v_57974 = v_57969 | v_57973;
assign v_57976 = v_57907 | v_57975;
assign v_57978 = v_57905 | v_57977;
assign v_57980 = v_57975 | v_57979;
assign v_57982 = v_57904 | v_57981;
assign v_57984 = v_57902 | v_57983;
assign v_57986 = v_57981 | v_57985;
assign v_57988 = v_57901 | v_57987;
assign v_57990 = v_57899 | v_57989;
assign v_57992 = v_57987 | v_57991;
assign v_57994 = v_57898 | v_57993;
assign v_57996 = v_57896 | v_57995;
assign v_57998 = v_57993 | v_57997;
assign v_58000 = v_57895 | v_57999;
assign v_58002 = v_57893 | v_58001;
assign v_58004 = v_57999 | v_58003;
assign v_58006 = v_57892 | v_58005;
assign v_58008 = v_57890 | v_58007;
assign v_58010 = v_58005 | v_58009;
assign v_58012 = v_57889 | v_58011;
assign v_58014 = v_57887 | v_58013;
assign v_58016 = v_58011 | v_58015;
assign v_58018 = v_57886 | v_58017;
assign v_58020 = v_57884 | v_58019;
assign v_58022 = v_58017 | v_58021;
assign v_58024 = v_57883 | v_58023;
assign v_58026 = v_57881 | v_58025;
assign v_58028 = v_58023 | v_58027;
assign v_58031 = ~v_57880 | v_58030;
assign v_58038 = v_57928 | v_58037;
assign v_58041 = v_58039 | v_58040;
assign v_58043 = v_57925 | v_58042;
assign v_58046 = v_58044 | v_58045;
assign v_58048 = v_57922 | v_58047;
assign v_58051 = v_58049 | v_58050;
assign v_58053 = v_57919 | v_58052;
assign v_58056 = v_58054 | v_58055;
assign v_58058 = v_57916 | v_58057;
assign v_58061 = v_58059 | v_58060;
assign v_58063 = v_57913 | v_58062;
assign v_58066 = v_58064 | v_58065;
assign v_58068 = v_57910 | v_58067;
assign v_58071 = v_58069 | v_58070;
assign v_58073 = v_57907 | v_58072;
assign v_58076 = v_58074 | v_58075;
assign v_58078 = v_57904 | v_58077;
assign v_58081 = v_58079 | v_58080;
assign v_58083 = v_57901 | v_58082;
assign v_58086 = v_58084 | v_58085;
assign v_58088 = v_57898 | v_58087;
assign v_58091 = v_58089 | v_58090;
assign v_58093 = v_57895 | v_58092;
assign v_58096 = v_58094 | v_58095;
assign v_58098 = v_57892 | v_58097;
assign v_58101 = v_58099 | v_58100;
assign v_58103 = v_57889 | v_58102;
assign v_58106 = v_58104 | v_58105;
assign v_58108 = v_57886 | v_58107;
assign v_58111 = v_58109 | v_58110;
assign v_58113 = v_57883 | v_58112;
assign v_58116 = v_58114 | v_58115;
assign v_58118 = v_57880 | v_58117;
assign v_58121 = v_57879 | v_58120;
assign v_58174 = v_58171 | v_58173;
assign v_58176 = v_58170 | v_58175;
assign v_58178 = v_58168 | v_58177;
assign v_58180 = v_58175 | v_58179;
assign v_58182 = v_58167 | v_58181;
assign v_58184 = v_58165 | v_58183;
assign v_58186 = v_58181 | v_58185;
assign v_58188 = v_58164 | v_58187;
assign v_58190 = v_58162 | v_58189;
assign v_58192 = v_58187 | v_58191;
assign v_58194 = v_58161 | v_58193;
assign v_58196 = v_58159 | v_58195;
assign v_58198 = v_58193 | v_58197;
assign v_58200 = v_58158 | v_58199;
assign v_58202 = v_58156 | v_58201;
assign v_58204 = v_58199 | v_58203;
assign v_58206 = v_58155 | v_58205;
assign v_58208 = v_58153 | v_58207;
assign v_58210 = v_58205 | v_58209;
assign v_58212 = v_58152 | v_58211;
assign v_58214 = v_58150 | v_58213;
assign v_58216 = v_58211 | v_58215;
assign v_58218 = v_58149 | v_58217;
assign v_58220 = v_58147 | v_58219;
assign v_58222 = v_58217 | v_58221;
assign v_58224 = v_58146 | v_58223;
assign v_58226 = v_58144 | v_58225;
assign v_58228 = v_58223 | v_58227;
assign v_58230 = v_58143 | v_58229;
assign v_58232 = v_58141 | v_58231;
assign v_58234 = v_58229 | v_58233;
assign v_58236 = v_58140 | v_58235;
assign v_58238 = v_58138 | v_58237;
assign v_58240 = v_58235 | v_58239;
assign v_58242 = v_58137 | v_58241;
assign v_58244 = v_58135 | v_58243;
assign v_58246 = v_58241 | v_58245;
assign v_58248 = v_58134 | v_58247;
assign v_58250 = v_58132 | v_58249;
assign v_58252 = v_58247 | v_58251;
assign v_58254 = v_58131 | v_58253;
assign v_58256 = v_58129 | v_58255;
assign v_58258 = v_58253 | v_58257;
assign v_58260 = v_58128 | v_58259;
assign v_58262 = v_58126 | v_58261;
assign v_58264 = v_58259 | v_58263;
assign v_58266 = v_58125 | v_58265;
assign v_58268 = v_58123 | v_58267;
assign v_58270 = v_58265 | v_58269;
assign v_58274 = v_58271 | v_58273;
assign v_58281 = v_58170 | v_58280;
assign v_58284 = v_58282 | v_58283;
assign v_58286 = v_58167 | v_58285;
assign v_58289 = v_58287 | v_58288;
assign v_58291 = v_58164 | v_58290;
assign v_58294 = v_58292 | v_58293;
assign v_58296 = v_58161 | v_58295;
assign v_58299 = v_58297 | v_58298;
assign v_58301 = v_58158 | v_58300;
assign v_58304 = v_58302 | v_58303;
assign v_58306 = v_58155 | v_58305;
assign v_58309 = v_58307 | v_58308;
assign v_58311 = v_58152 | v_58310;
assign v_58314 = v_58312 | v_58313;
assign v_58316 = v_58149 | v_58315;
assign v_58319 = v_58317 | v_58318;
assign v_58321 = v_58146 | v_58320;
assign v_58324 = v_58322 | v_58323;
assign v_58326 = v_58143 | v_58325;
assign v_58329 = v_58327 | v_58328;
assign v_58331 = v_58140 | v_58330;
assign v_58334 = v_58332 | v_58333;
assign v_58336 = v_58137 | v_58335;
assign v_58339 = v_58337 | v_58338;
assign v_58341 = v_58134 | v_58340;
assign v_58344 = v_58342 | v_58343;
assign v_58346 = v_58131 | v_58345;
assign v_58349 = v_58347 | v_58348;
assign v_58351 = v_58128 | v_58350;
assign v_58354 = v_58352 | v_58353;
assign v_58356 = v_58125 | v_58355;
assign v_58359 = v_58357 | v_58358;
assign v_58361 = v_58359 | v_58360;
assign v_58364 = v_58122 | v_58363;
assign v_58435 = v_58432 | v_58434;
assign v_58437 = v_58430 | v_58436;
assign v_58439 = v_58428 | v_58438;
assign v_58441 = v_58436 | v_58440;
assign v_58443 = v_58426 | v_58442;
assign v_58445 = v_58424 | v_58444;
assign v_58447 = v_58442 | v_58446;
assign v_58449 = v_58422 | v_58448;
assign v_58451 = v_58420 | v_58450;
assign v_58453 = v_58448 | v_58452;
assign v_58455 = v_58418 | v_58454;
assign v_58457 = v_58416 | v_58456;
assign v_58459 = v_58454 | v_58458;
assign v_58461 = v_58414 | v_58460;
assign v_58463 = v_58412 | v_58462;
assign v_58465 = v_58460 | v_58464;
assign v_58467 = v_58410 | v_58466;
assign v_58469 = v_58408 | v_58468;
assign v_58471 = v_58466 | v_58470;
assign v_58473 = v_58406 | v_58472;
assign v_58475 = v_58404 | v_58474;
assign v_58477 = v_58472 | v_58476;
assign v_58479 = v_58402 | v_58478;
assign v_58481 = v_58400 | v_58480;
assign v_58483 = v_58478 | v_58482;
assign v_58485 = v_58398 | v_58484;
assign v_58487 = v_58396 | v_58486;
assign v_58489 = v_58484 | v_58488;
assign v_58491 = v_58394 | v_58490;
assign v_58493 = v_58392 | v_58492;
assign v_58495 = v_58490 | v_58494;
assign v_58497 = v_58390 | v_58496;
assign v_58499 = v_58388 | v_58498;
assign v_58501 = v_58496 | v_58500;
assign v_58503 = v_58386 | v_58502;
assign v_58505 = v_58384 | v_58504;
assign v_58507 = v_58502 | v_58506;
assign v_58509 = v_58382 | v_58508;
assign v_58511 = v_58379 | v_58510;
assign v_58513 = v_58508 | v_58512;
assign v_58515 = v_58378 | v_58514;
assign v_58517 = v_58375 | v_58516;
assign v_58519 = v_58514 | v_58518;
assign v_58521 = v_58374 | v_58520;
assign v_58523 = v_58371 | v_58522;
assign v_58525 = v_58520 | v_58524;
assign v_58527 = v_58370 | v_58526;
assign v_58529 = v_58367 | v_58528;
assign v_58531 = v_58526 | v_58530;
assign v_58534 = ~v_58366 | v_58533;
assign v_58541 = v_58430 | v_58540;
assign v_58544 = v_58542 | v_58543;
assign v_58546 = v_58426 | v_58545;
assign v_58549 = v_58547 | v_58548;
assign v_58551 = v_58422 | v_58550;
assign v_58554 = v_58552 | v_58553;
assign v_58556 = v_58418 | v_58555;
assign v_58559 = v_58557 | v_58558;
assign v_58561 = v_58414 | v_58560;
assign v_58564 = v_58562 | v_58563;
assign v_58566 = v_58410 | v_58565;
assign v_58569 = v_58567 | v_58568;
assign v_58571 = v_58406 | v_58570;
assign v_58574 = v_58572 | v_58573;
assign v_58576 = v_58402 | v_58575;
assign v_58579 = v_58577 | v_58578;
assign v_58581 = v_58398 | v_58580;
assign v_58584 = v_58582 | v_58583;
assign v_58586 = v_58394 | v_58585;
assign v_58589 = v_58587 | v_58588;
assign v_58591 = v_58390 | v_58590;
assign v_58594 = v_58592 | v_58593;
assign v_58596 = v_58386 | v_58595;
assign v_58599 = v_58597 | v_58598;
assign v_58601 = v_58382 | v_58600;
assign v_58604 = v_58602 | v_58603;
assign v_58606 = v_58378 | v_58605;
assign v_58609 = v_58607 | v_58608;
assign v_58611 = v_58374 | v_58610;
assign v_58614 = v_58612 | v_58613;
assign v_58616 = v_58370 | v_58615;
assign v_58619 = v_58617 | v_58618;
assign v_58621 = v_58366 | v_58620;
assign v_58624 = v_58365 | v_58623;
assign v_58678 = v_58675 | v_58677;
assign v_58680 = v_58674 | v_58679;
assign v_58682 = v_58672 | v_58681;
assign v_58684 = v_58679 | v_58683;
assign v_58686 = v_58671 | v_58685;
assign v_58688 = v_58669 | v_58687;
assign v_58690 = v_58685 | v_58689;
assign v_58692 = v_58668 | v_58691;
assign v_58694 = v_58666 | v_58693;
assign v_58696 = v_58691 | v_58695;
assign v_58698 = v_58665 | v_58697;
assign v_58700 = v_58663 | v_58699;
assign v_58702 = v_58697 | v_58701;
assign v_58704 = v_58662 | v_58703;
assign v_58706 = v_58660 | v_58705;
assign v_58708 = v_58703 | v_58707;
assign v_58710 = v_58659 | v_58709;
assign v_58712 = v_58657 | v_58711;
assign v_58714 = v_58709 | v_58713;
assign v_58716 = v_58656 | v_58715;
assign v_58718 = v_58654 | v_58717;
assign v_58720 = v_58715 | v_58719;
assign v_58722 = v_58653 | v_58721;
assign v_58724 = v_58651 | v_58723;
assign v_58726 = v_58721 | v_58725;
assign v_58728 = v_58650 | v_58727;
assign v_58730 = v_58648 | v_58729;
assign v_58732 = v_58727 | v_58731;
assign v_58734 = v_58647 | v_58733;
assign v_58736 = v_58645 | v_58735;
assign v_58738 = v_58733 | v_58737;
assign v_58740 = v_58644 | v_58739;
assign v_58742 = v_58642 | v_58741;
assign v_58744 = v_58739 | v_58743;
assign v_58746 = v_58641 | v_58745;
assign v_58748 = v_58639 | v_58747;
assign v_58750 = v_58745 | v_58749;
assign v_58752 = v_58638 | v_58751;
assign v_58754 = v_58636 | v_58753;
assign v_58756 = v_58751 | v_58755;
assign v_58758 = v_58635 | v_58757;
assign v_58760 = v_58633 | v_58759;
assign v_58762 = v_58757 | v_58761;
assign v_58764 = v_58632 | v_58763;
assign v_58766 = v_58630 | v_58765;
assign v_58768 = v_58763 | v_58767;
assign v_58770 = v_58629 | v_58769;
assign v_58772 = v_58627 | v_58771;
assign v_58774 = v_58769 | v_58773;
assign v_58777 = ~v_58626 | v_58776;
assign v_58784 = v_58674 | v_58783;
assign v_58787 = v_58785 | v_58786;
assign v_58789 = v_58671 | v_58788;
assign v_58792 = v_58790 | v_58791;
assign v_58794 = v_58668 | v_58793;
assign v_58797 = v_58795 | v_58796;
assign v_58799 = v_58665 | v_58798;
assign v_58802 = v_58800 | v_58801;
assign v_58804 = v_58662 | v_58803;
assign v_58807 = v_58805 | v_58806;
assign v_58809 = v_58659 | v_58808;
assign v_58812 = v_58810 | v_58811;
assign v_58814 = v_58656 | v_58813;
assign v_58817 = v_58815 | v_58816;
assign v_58819 = v_58653 | v_58818;
assign v_58822 = v_58820 | v_58821;
assign v_58824 = v_58650 | v_58823;
assign v_58827 = v_58825 | v_58826;
assign v_58829 = v_58647 | v_58828;
assign v_58832 = v_58830 | v_58831;
assign v_58834 = v_58644 | v_58833;
assign v_58837 = v_58835 | v_58836;
assign v_58839 = v_58641 | v_58838;
assign v_58842 = v_58840 | v_58841;
assign v_58844 = v_58638 | v_58843;
assign v_58847 = v_58845 | v_58846;
assign v_58849 = v_58635 | v_58848;
assign v_58852 = v_58850 | v_58851;
assign v_58854 = v_58632 | v_58853;
assign v_58857 = v_58855 | v_58856;
assign v_58859 = v_58629 | v_58858;
assign v_58862 = v_58860 | v_58861;
assign v_58864 = v_58626 | v_58863;
assign v_58867 = v_58625 | v_58866;
assign v_58921 = v_58918 | v_58920;
assign v_58923 = v_58917 | v_58922;
assign v_58925 = v_58915 | v_58924;
assign v_58927 = v_58922 | v_58926;
assign v_58929 = v_58914 | v_58928;
assign v_58931 = v_58912 | v_58930;
assign v_58933 = v_58928 | v_58932;
assign v_58935 = v_58911 | v_58934;
assign v_58937 = v_58909 | v_58936;
assign v_58939 = v_58934 | v_58938;
assign v_58941 = v_58908 | v_58940;
assign v_58943 = v_58906 | v_58942;
assign v_58945 = v_58940 | v_58944;
assign v_58947 = v_58905 | v_58946;
assign v_58949 = v_58903 | v_58948;
assign v_58951 = v_58946 | v_58950;
assign v_58953 = v_58902 | v_58952;
assign v_58955 = v_58900 | v_58954;
assign v_58957 = v_58952 | v_58956;
assign v_58959 = v_58899 | v_58958;
assign v_58961 = v_58897 | v_58960;
assign v_58963 = v_58958 | v_58962;
assign v_58965 = v_58896 | v_58964;
assign v_58967 = v_58894 | v_58966;
assign v_58969 = v_58964 | v_58968;
assign v_58971 = v_58893 | v_58970;
assign v_58973 = v_58891 | v_58972;
assign v_58975 = v_58970 | v_58974;
assign v_58977 = v_58890 | v_58976;
assign v_58979 = v_58888 | v_58978;
assign v_58981 = v_58976 | v_58980;
assign v_58983 = v_58887 | v_58982;
assign v_58985 = v_58885 | v_58984;
assign v_58987 = v_58982 | v_58986;
assign v_58989 = v_58884 | v_58988;
assign v_58991 = v_58882 | v_58990;
assign v_58993 = v_58988 | v_58992;
assign v_58995 = v_58881 | v_58994;
assign v_58997 = v_58879 | v_58996;
assign v_58999 = v_58994 | v_58998;
assign v_59001 = v_58878 | v_59000;
assign v_59003 = v_58876 | v_59002;
assign v_59005 = v_59000 | v_59004;
assign v_59007 = v_58875 | v_59006;
assign v_59009 = v_58873 | v_59008;
assign v_59011 = v_59006 | v_59010;
assign v_59013 = v_58872 | v_59012;
assign v_59015 = v_58870 | v_59014;
assign v_59017 = v_59012 | v_59016;
assign v_59020 = ~v_58869 | v_59019;
assign v_59027 = v_58917 | v_59026;
assign v_59030 = v_59028 | v_59029;
assign v_59032 = v_58914 | v_59031;
assign v_59035 = v_59033 | v_59034;
assign v_59037 = v_58911 | v_59036;
assign v_59040 = v_59038 | v_59039;
assign v_59042 = v_58908 | v_59041;
assign v_59045 = v_59043 | v_59044;
assign v_59047 = v_58905 | v_59046;
assign v_59050 = v_59048 | v_59049;
assign v_59052 = v_58902 | v_59051;
assign v_59055 = v_59053 | v_59054;
assign v_59057 = v_58899 | v_59056;
assign v_59060 = v_59058 | v_59059;
assign v_59062 = v_58896 | v_59061;
assign v_59065 = v_59063 | v_59064;
assign v_59067 = v_58893 | v_59066;
assign v_59070 = v_59068 | v_59069;
assign v_59072 = v_58890 | v_59071;
assign v_59075 = v_59073 | v_59074;
assign v_59077 = v_58887 | v_59076;
assign v_59080 = v_59078 | v_59079;
assign v_59082 = v_58884 | v_59081;
assign v_59085 = v_59083 | v_59084;
assign v_59087 = v_58881 | v_59086;
assign v_59090 = v_59088 | v_59089;
assign v_59092 = v_58878 | v_59091;
assign v_59095 = v_59093 | v_59094;
assign v_59097 = v_58875 | v_59096;
assign v_59100 = v_59098 | v_59099;
assign v_59102 = v_58872 | v_59101;
assign v_59105 = v_59103 | v_59104;
assign v_59107 = v_58869 | v_59106;
assign v_59110 = v_58868 | v_59109;
assign v_59164 = v_59161 | v_59163;
assign v_59166 = v_59160 | v_59165;
assign v_59168 = v_59158 | v_59167;
assign v_59170 = v_59165 | v_59169;
assign v_59172 = v_59157 | v_59171;
assign v_59174 = v_59155 | v_59173;
assign v_59176 = v_59171 | v_59175;
assign v_59178 = v_59154 | v_59177;
assign v_59180 = v_59152 | v_59179;
assign v_59182 = v_59177 | v_59181;
assign v_59184 = v_59151 | v_59183;
assign v_59186 = v_59149 | v_59185;
assign v_59188 = v_59183 | v_59187;
assign v_59190 = v_59148 | v_59189;
assign v_59192 = v_59146 | v_59191;
assign v_59194 = v_59189 | v_59193;
assign v_59196 = v_59145 | v_59195;
assign v_59198 = v_59143 | v_59197;
assign v_59200 = v_59195 | v_59199;
assign v_59202 = v_59142 | v_59201;
assign v_59204 = v_59140 | v_59203;
assign v_59206 = v_59201 | v_59205;
assign v_59208 = v_59139 | v_59207;
assign v_59210 = v_59137 | v_59209;
assign v_59212 = v_59207 | v_59211;
assign v_59214 = v_59136 | v_59213;
assign v_59216 = v_59134 | v_59215;
assign v_59218 = v_59213 | v_59217;
assign v_59220 = v_59133 | v_59219;
assign v_59222 = v_59131 | v_59221;
assign v_59224 = v_59219 | v_59223;
assign v_59226 = v_59130 | v_59225;
assign v_59228 = v_59128 | v_59227;
assign v_59230 = v_59225 | v_59229;
assign v_59232 = v_59127 | v_59231;
assign v_59234 = v_59125 | v_59233;
assign v_59236 = v_59231 | v_59235;
assign v_59238 = v_59124 | v_59237;
assign v_59240 = v_59122 | v_59239;
assign v_59242 = v_59237 | v_59241;
assign v_59244 = v_59121 | v_59243;
assign v_59246 = v_59119 | v_59245;
assign v_59248 = v_59243 | v_59247;
assign v_59250 = v_59118 | v_59249;
assign v_59252 = v_59116 | v_59251;
assign v_59254 = v_59249 | v_59253;
assign v_59256 = v_59115 | v_59255;
assign v_59258 = v_59113 | v_59257;
assign v_59260 = v_59255 | v_59259;
assign v_59263 = ~v_59112 | v_59262;
assign v_59270 = v_59160 | v_59269;
assign v_59273 = v_59271 | v_59272;
assign v_59275 = v_59157 | v_59274;
assign v_59278 = v_59276 | v_59277;
assign v_59280 = v_59154 | v_59279;
assign v_59283 = v_59281 | v_59282;
assign v_59285 = v_59151 | v_59284;
assign v_59288 = v_59286 | v_59287;
assign v_59290 = v_59148 | v_59289;
assign v_59293 = v_59291 | v_59292;
assign v_59295 = v_59145 | v_59294;
assign v_59298 = v_59296 | v_59297;
assign v_59300 = v_59142 | v_59299;
assign v_59303 = v_59301 | v_59302;
assign v_59305 = v_59139 | v_59304;
assign v_59308 = v_59306 | v_59307;
assign v_59310 = v_59136 | v_59309;
assign v_59313 = v_59311 | v_59312;
assign v_59315 = v_59133 | v_59314;
assign v_59318 = v_59316 | v_59317;
assign v_59320 = v_59130 | v_59319;
assign v_59323 = v_59321 | v_59322;
assign v_59325 = v_59127 | v_59324;
assign v_59328 = v_59326 | v_59327;
assign v_59330 = v_59124 | v_59329;
assign v_59333 = v_59331 | v_59332;
assign v_59335 = v_59121 | v_59334;
assign v_59338 = v_59336 | v_59337;
assign v_59340 = v_59118 | v_59339;
assign v_59343 = v_59341 | v_59342;
assign v_59345 = v_59115 | v_59344;
assign v_59348 = v_59346 | v_59347;
assign v_59350 = v_59112 | v_59349;
assign v_59353 = v_59111 | v_59352;
assign v_59407 = v_59404 | v_59406;
assign v_59409 = v_59403 | v_59408;
assign v_59411 = v_59401 | v_59410;
assign v_59413 = v_59408 | v_59412;
assign v_59415 = v_59400 | v_59414;
assign v_59417 = v_59398 | v_59416;
assign v_59419 = v_59414 | v_59418;
assign v_59421 = v_59397 | v_59420;
assign v_59423 = v_59395 | v_59422;
assign v_59425 = v_59420 | v_59424;
assign v_59427 = v_59394 | v_59426;
assign v_59429 = v_59392 | v_59428;
assign v_59431 = v_59426 | v_59430;
assign v_59433 = v_59391 | v_59432;
assign v_59435 = v_59389 | v_59434;
assign v_59437 = v_59432 | v_59436;
assign v_59439 = v_59388 | v_59438;
assign v_59441 = v_59386 | v_59440;
assign v_59443 = v_59438 | v_59442;
assign v_59445 = v_59385 | v_59444;
assign v_59447 = v_59383 | v_59446;
assign v_59449 = v_59444 | v_59448;
assign v_59451 = v_59382 | v_59450;
assign v_59453 = v_59380 | v_59452;
assign v_59455 = v_59450 | v_59454;
assign v_59457 = v_59379 | v_59456;
assign v_59459 = v_59377 | v_59458;
assign v_59461 = v_59456 | v_59460;
assign v_59463 = v_59376 | v_59462;
assign v_59465 = v_59374 | v_59464;
assign v_59467 = v_59462 | v_59466;
assign v_59469 = v_59373 | v_59468;
assign v_59471 = v_59371 | v_59470;
assign v_59473 = v_59468 | v_59472;
assign v_59475 = v_59370 | v_59474;
assign v_59477 = v_59368 | v_59476;
assign v_59479 = v_59474 | v_59478;
assign v_59481 = v_59367 | v_59480;
assign v_59483 = v_59365 | v_59482;
assign v_59485 = v_59480 | v_59484;
assign v_59487 = v_59364 | v_59486;
assign v_59489 = v_59362 | v_59488;
assign v_59491 = v_59486 | v_59490;
assign v_59493 = v_59361 | v_59492;
assign v_59495 = v_59359 | v_59494;
assign v_59497 = v_59492 | v_59496;
assign v_59499 = v_59358 | v_59498;
assign v_59501 = v_59356 | v_59500;
assign v_59503 = v_59498 | v_59502;
assign v_59506 = ~v_59355 | v_59505;
assign v_59513 = v_59403 | v_59512;
assign v_59516 = v_59514 | v_59515;
assign v_59518 = v_59400 | v_59517;
assign v_59521 = v_59519 | v_59520;
assign v_59523 = v_59397 | v_59522;
assign v_59526 = v_59524 | v_59525;
assign v_59528 = v_59394 | v_59527;
assign v_59531 = v_59529 | v_59530;
assign v_59533 = v_59391 | v_59532;
assign v_59536 = v_59534 | v_59535;
assign v_59538 = v_59388 | v_59537;
assign v_59541 = v_59539 | v_59540;
assign v_59543 = v_59385 | v_59542;
assign v_59546 = v_59544 | v_59545;
assign v_59548 = v_59382 | v_59547;
assign v_59551 = v_59549 | v_59550;
assign v_59553 = v_59379 | v_59552;
assign v_59556 = v_59554 | v_59555;
assign v_59558 = v_59376 | v_59557;
assign v_59561 = v_59559 | v_59560;
assign v_59563 = v_59373 | v_59562;
assign v_59566 = v_59564 | v_59565;
assign v_59568 = v_59370 | v_59567;
assign v_59571 = v_59569 | v_59570;
assign v_59573 = v_59367 | v_59572;
assign v_59576 = v_59574 | v_59575;
assign v_59578 = v_59364 | v_59577;
assign v_59581 = v_59579 | v_59580;
assign v_59583 = v_59361 | v_59582;
assign v_59586 = v_59584 | v_59585;
assign v_59588 = v_59358 | v_59587;
assign v_59591 = v_59589 | v_59590;
assign v_59593 = v_59355 | v_59592;
assign v_59596 = v_59354 | v_59595;
assign v_59650 = v_59647 | v_59649;
assign v_59652 = v_59646 | v_59651;
assign v_59654 = v_59644 | v_59653;
assign v_59656 = v_59651 | v_59655;
assign v_59658 = v_59643 | v_59657;
assign v_59660 = v_59641 | v_59659;
assign v_59662 = v_59657 | v_59661;
assign v_59664 = v_59640 | v_59663;
assign v_59666 = v_59638 | v_59665;
assign v_59668 = v_59663 | v_59667;
assign v_59670 = v_59637 | v_59669;
assign v_59672 = v_59635 | v_59671;
assign v_59674 = v_59669 | v_59673;
assign v_59676 = v_59634 | v_59675;
assign v_59678 = v_59632 | v_59677;
assign v_59680 = v_59675 | v_59679;
assign v_59682 = v_59631 | v_59681;
assign v_59684 = v_59629 | v_59683;
assign v_59686 = v_59681 | v_59685;
assign v_59688 = v_59628 | v_59687;
assign v_59690 = v_59626 | v_59689;
assign v_59692 = v_59687 | v_59691;
assign v_59694 = v_59625 | v_59693;
assign v_59696 = v_59623 | v_59695;
assign v_59698 = v_59693 | v_59697;
assign v_59700 = v_59622 | v_59699;
assign v_59702 = v_59620 | v_59701;
assign v_59704 = v_59699 | v_59703;
assign v_59706 = v_59619 | v_59705;
assign v_59708 = v_59617 | v_59707;
assign v_59710 = v_59705 | v_59709;
assign v_59712 = v_59616 | v_59711;
assign v_59714 = v_59614 | v_59713;
assign v_59716 = v_59711 | v_59715;
assign v_59718 = v_59613 | v_59717;
assign v_59720 = v_59611 | v_59719;
assign v_59722 = v_59717 | v_59721;
assign v_59724 = v_59610 | v_59723;
assign v_59726 = v_59608 | v_59725;
assign v_59728 = v_59723 | v_59727;
assign v_59730 = v_59607 | v_59729;
assign v_59732 = v_59605 | v_59731;
assign v_59734 = v_59729 | v_59733;
assign v_59736 = v_59604 | v_59735;
assign v_59738 = v_59602 | v_59737;
assign v_59740 = v_59735 | v_59739;
assign v_59742 = v_59601 | v_59741;
assign v_59744 = v_59599 | v_59743;
assign v_59746 = v_59741 | v_59745;
assign v_59749 = ~v_59598 | v_59748;
assign v_59756 = v_59646 | v_59755;
assign v_59759 = v_59757 | v_59758;
assign v_59761 = v_59643 | v_59760;
assign v_59764 = v_59762 | v_59763;
assign v_59766 = v_59640 | v_59765;
assign v_59769 = v_59767 | v_59768;
assign v_59771 = v_59637 | v_59770;
assign v_59774 = v_59772 | v_59773;
assign v_59776 = v_59634 | v_59775;
assign v_59779 = v_59777 | v_59778;
assign v_59781 = v_59631 | v_59780;
assign v_59784 = v_59782 | v_59783;
assign v_59786 = v_59628 | v_59785;
assign v_59789 = v_59787 | v_59788;
assign v_59791 = v_59625 | v_59790;
assign v_59794 = v_59792 | v_59793;
assign v_59796 = v_59622 | v_59795;
assign v_59799 = v_59797 | v_59798;
assign v_59801 = v_59619 | v_59800;
assign v_59804 = v_59802 | v_59803;
assign v_59806 = v_59616 | v_59805;
assign v_59809 = v_59807 | v_59808;
assign v_59811 = v_59613 | v_59810;
assign v_59814 = v_59812 | v_59813;
assign v_59816 = v_59610 | v_59815;
assign v_59819 = v_59817 | v_59818;
assign v_59821 = v_59607 | v_59820;
assign v_59824 = v_59822 | v_59823;
assign v_59826 = v_59604 | v_59825;
assign v_59829 = v_59827 | v_59828;
assign v_59831 = v_59601 | v_59830;
assign v_59834 = v_59832 | v_59833;
assign v_59836 = v_59598 | v_59835;
assign v_59839 = v_59597 | v_59838;
assign v_59893 = v_59890 | v_59892;
assign v_59895 = v_59889 | v_59894;
assign v_59897 = v_59887 | v_59896;
assign v_59899 = v_59894 | v_59898;
assign v_59901 = v_59886 | v_59900;
assign v_59903 = v_59884 | v_59902;
assign v_59905 = v_59900 | v_59904;
assign v_59907 = v_59883 | v_59906;
assign v_59909 = v_59881 | v_59908;
assign v_59911 = v_59906 | v_59910;
assign v_59913 = v_59880 | v_59912;
assign v_59915 = v_59878 | v_59914;
assign v_59917 = v_59912 | v_59916;
assign v_59919 = v_59877 | v_59918;
assign v_59921 = v_59875 | v_59920;
assign v_59923 = v_59918 | v_59922;
assign v_59925 = v_59874 | v_59924;
assign v_59927 = v_59872 | v_59926;
assign v_59929 = v_59924 | v_59928;
assign v_59931 = v_59871 | v_59930;
assign v_59933 = v_59869 | v_59932;
assign v_59935 = v_59930 | v_59934;
assign v_59937 = v_59868 | v_59936;
assign v_59939 = v_59866 | v_59938;
assign v_59941 = v_59936 | v_59940;
assign v_59943 = v_59865 | v_59942;
assign v_59945 = v_59863 | v_59944;
assign v_59947 = v_59942 | v_59946;
assign v_59949 = v_59862 | v_59948;
assign v_59951 = v_59860 | v_59950;
assign v_59953 = v_59948 | v_59952;
assign v_59955 = v_59859 | v_59954;
assign v_59957 = v_59857 | v_59956;
assign v_59959 = v_59954 | v_59958;
assign v_59961 = v_59856 | v_59960;
assign v_59963 = v_59854 | v_59962;
assign v_59965 = v_59960 | v_59964;
assign v_59967 = v_59853 | v_59966;
assign v_59969 = v_59851 | v_59968;
assign v_59971 = v_59966 | v_59970;
assign v_59973 = v_59850 | v_59972;
assign v_59975 = v_59848 | v_59974;
assign v_59977 = v_59972 | v_59976;
assign v_59979 = v_59847 | v_59978;
assign v_59981 = v_59845 | v_59980;
assign v_59983 = v_59978 | v_59982;
assign v_59985 = v_59844 | v_59984;
assign v_59987 = v_59842 | v_59986;
assign v_59989 = v_59984 | v_59988;
assign v_59992 = ~v_59841 | v_59991;
assign v_59999 = v_59889 | v_59998;
assign v_60002 = v_60000 | v_60001;
assign v_60004 = v_59886 | v_60003;
assign v_60007 = v_60005 | v_60006;
assign v_60009 = v_59883 | v_60008;
assign v_60012 = v_60010 | v_60011;
assign v_60014 = v_59880 | v_60013;
assign v_60017 = v_60015 | v_60016;
assign v_60019 = v_59877 | v_60018;
assign v_60022 = v_60020 | v_60021;
assign v_60024 = v_59874 | v_60023;
assign v_60027 = v_60025 | v_60026;
assign v_60029 = v_59871 | v_60028;
assign v_60032 = v_60030 | v_60031;
assign v_60034 = v_59868 | v_60033;
assign v_60037 = v_60035 | v_60036;
assign v_60039 = v_59865 | v_60038;
assign v_60042 = v_60040 | v_60041;
assign v_60044 = v_59862 | v_60043;
assign v_60047 = v_60045 | v_60046;
assign v_60049 = v_59859 | v_60048;
assign v_60052 = v_60050 | v_60051;
assign v_60054 = v_59856 | v_60053;
assign v_60057 = v_60055 | v_60056;
assign v_60059 = v_59853 | v_60058;
assign v_60062 = v_60060 | v_60061;
assign v_60064 = v_59850 | v_60063;
assign v_60067 = v_60065 | v_60066;
assign v_60069 = v_59847 | v_60068;
assign v_60072 = v_60070 | v_60071;
assign v_60074 = v_59844 | v_60073;
assign v_60077 = v_60075 | v_60076;
assign v_60079 = v_59841 | v_60078;
assign v_60082 = v_59840 | v_60081;
assign v_60136 = v_60133 | v_60135;
assign v_60138 = v_60132 | v_60137;
assign v_60140 = v_60130 | v_60139;
assign v_60142 = v_60137 | v_60141;
assign v_60144 = v_60129 | v_60143;
assign v_60146 = v_60127 | v_60145;
assign v_60148 = v_60143 | v_60147;
assign v_60150 = v_60126 | v_60149;
assign v_60152 = v_60124 | v_60151;
assign v_60154 = v_60149 | v_60153;
assign v_60156 = v_60123 | v_60155;
assign v_60158 = v_60121 | v_60157;
assign v_60160 = v_60155 | v_60159;
assign v_60162 = v_60120 | v_60161;
assign v_60164 = v_60118 | v_60163;
assign v_60166 = v_60161 | v_60165;
assign v_60168 = v_60117 | v_60167;
assign v_60170 = v_60115 | v_60169;
assign v_60172 = v_60167 | v_60171;
assign v_60174 = v_60114 | v_60173;
assign v_60176 = v_60112 | v_60175;
assign v_60178 = v_60173 | v_60177;
assign v_60180 = v_60111 | v_60179;
assign v_60182 = v_60109 | v_60181;
assign v_60184 = v_60179 | v_60183;
assign v_60186 = v_60108 | v_60185;
assign v_60188 = v_60106 | v_60187;
assign v_60190 = v_60185 | v_60189;
assign v_60192 = v_60105 | v_60191;
assign v_60194 = v_60103 | v_60193;
assign v_60196 = v_60191 | v_60195;
assign v_60198 = v_60102 | v_60197;
assign v_60200 = v_60100 | v_60199;
assign v_60202 = v_60197 | v_60201;
assign v_60204 = v_60099 | v_60203;
assign v_60206 = v_60097 | v_60205;
assign v_60208 = v_60203 | v_60207;
assign v_60210 = v_60096 | v_60209;
assign v_60212 = v_60094 | v_60211;
assign v_60214 = v_60209 | v_60213;
assign v_60216 = v_60093 | v_60215;
assign v_60218 = v_60091 | v_60217;
assign v_60220 = v_60215 | v_60219;
assign v_60222 = v_60090 | v_60221;
assign v_60224 = v_60088 | v_60223;
assign v_60226 = v_60221 | v_60225;
assign v_60228 = v_60087 | v_60227;
assign v_60230 = v_60085 | v_60229;
assign v_60232 = v_60227 | v_60231;
assign v_60235 = ~v_60084 | v_60234;
assign v_60242 = v_60132 | v_60241;
assign v_60245 = v_60243 | v_60244;
assign v_60247 = v_60129 | v_60246;
assign v_60250 = v_60248 | v_60249;
assign v_60252 = v_60126 | v_60251;
assign v_60255 = v_60253 | v_60254;
assign v_60257 = v_60123 | v_60256;
assign v_60260 = v_60258 | v_60259;
assign v_60262 = v_60120 | v_60261;
assign v_60265 = v_60263 | v_60264;
assign v_60267 = v_60117 | v_60266;
assign v_60270 = v_60268 | v_60269;
assign v_60272 = v_60114 | v_60271;
assign v_60275 = v_60273 | v_60274;
assign v_60277 = v_60111 | v_60276;
assign v_60280 = v_60278 | v_60279;
assign v_60282 = v_60108 | v_60281;
assign v_60285 = v_60283 | v_60284;
assign v_60287 = v_60105 | v_60286;
assign v_60290 = v_60288 | v_60289;
assign v_60292 = v_60102 | v_60291;
assign v_60295 = v_60293 | v_60294;
assign v_60297 = v_60099 | v_60296;
assign v_60300 = v_60298 | v_60299;
assign v_60302 = v_60096 | v_60301;
assign v_60305 = v_60303 | v_60304;
assign v_60307 = v_60093 | v_60306;
assign v_60310 = v_60308 | v_60309;
assign v_60312 = v_60090 | v_60311;
assign v_60315 = v_60313 | v_60314;
assign v_60317 = v_60087 | v_60316;
assign v_60320 = v_60318 | v_60319;
assign v_60322 = v_60084 | v_60321;
assign v_60325 = v_60083 | v_60324;
assign v_60379 = v_60376 | v_60378;
assign v_60381 = v_60375 | v_60380;
assign v_60383 = v_60373 | v_60382;
assign v_60385 = v_60380 | v_60384;
assign v_60387 = v_60372 | v_60386;
assign v_60389 = v_60370 | v_60388;
assign v_60391 = v_60386 | v_60390;
assign v_60393 = v_60369 | v_60392;
assign v_60395 = v_60367 | v_60394;
assign v_60397 = v_60392 | v_60396;
assign v_60399 = v_60366 | v_60398;
assign v_60401 = v_60364 | v_60400;
assign v_60403 = v_60398 | v_60402;
assign v_60405 = v_60363 | v_60404;
assign v_60407 = v_60361 | v_60406;
assign v_60409 = v_60404 | v_60408;
assign v_60411 = v_60360 | v_60410;
assign v_60413 = v_60358 | v_60412;
assign v_60415 = v_60410 | v_60414;
assign v_60417 = v_60357 | v_60416;
assign v_60419 = v_60355 | v_60418;
assign v_60421 = v_60416 | v_60420;
assign v_60423 = v_60354 | v_60422;
assign v_60425 = v_60352 | v_60424;
assign v_60427 = v_60422 | v_60426;
assign v_60429 = v_60351 | v_60428;
assign v_60431 = v_60349 | v_60430;
assign v_60433 = v_60428 | v_60432;
assign v_60435 = v_60348 | v_60434;
assign v_60437 = v_60346 | v_60436;
assign v_60439 = v_60434 | v_60438;
assign v_60441 = v_60345 | v_60440;
assign v_60443 = v_60343 | v_60442;
assign v_60445 = v_60440 | v_60444;
assign v_60447 = v_60342 | v_60446;
assign v_60449 = v_60340 | v_60448;
assign v_60451 = v_60446 | v_60450;
assign v_60453 = v_60339 | v_60452;
assign v_60455 = v_60337 | v_60454;
assign v_60457 = v_60452 | v_60456;
assign v_60459 = v_60336 | v_60458;
assign v_60461 = v_60334 | v_60460;
assign v_60463 = v_60458 | v_60462;
assign v_60465 = v_60333 | v_60464;
assign v_60467 = v_60331 | v_60466;
assign v_60469 = v_60464 | v_60468;
assign v_60471 = v_60330 | v_60470;
assign v_60473 = v_60328 | v_60472;
assign v_60475 = v_60470 | v_60474;
assign v_60478 = ~v_60327 | v_60477;
assign v_60485 = v_60375 | v_60484;
assign v_60488 = v_60486 | v_60487;
assign v_60490 = v_60372 | v_60489;
assign v_60493 = v_60491 | v_60492;
assign v_60495 = v_60369 | v_60494;
assign v_60498 = v_60496 | v_60497;
assign v_60500 = v_60366 | v_60499;
assign v_60503 = v_60501 | v_60502;
assign v_60505 = v_60363 | v_60504;
assign v_60508 = v_60506 | v_60507;
assign v_60510 = v_60360 | v_60509;
assign v_60513 = v_60511 | v_60512;
assign v_60515 = v_60357 | v_60514;
assign v_60518 = v_60516 | v_60517;
assign v_60520 = v_60354 | v_60519;
assign v_60523 = v_60521 | v_60522;
assign v_60525 = v_60351 | v_60524;
assign v_60528 = v_60526 | v_60527;
assign v_60530 = v_60348 | v_60529;
assign v_60533 = v_60531 | v_60532;
assign v_60535 = v_60345 | v_60534;
assign v_60538 = v_60536 | v_60537;
assign v_60540 = v_60342 | v_60539;
assign v_60543 = v_60541 | v_60542;
assign v_60545 = v_60339 | v_60544;
assign v_60548 = v_60546 | v_60547;
assign v_60550 = v_60336 | v_60549;
assign v_60553 = v_60551 | v_60552;
assign v_60555 = v_60333 | v_60554;
assign v_60558 = v_60556 | v_60557;
assign v_60560 = v_60330 | v_60559;
assign v_60563 = v_60561 | v_60562;
assign v_60565 = v_60327 | v_60564;
assign v_60568 = v_60326 | v_60567;
assign v_60622 = v_60619 | v_60621;
assign v_60624 = v_60618 | v_60623;
assign v_60626 = v_60616 | v_60625;
assign v_60628 = v_60623 | v_60627;
assign v_60630 = v_60615 | v_60629;
assign v_60632 = v_60613 | v_60631;
assign v_60634 = v_60629 | v_60633;
assign v_60636 = v_60612 | v_60635;
assign v_60638 = v_60610 | v_60637;
assign v_60640 = v_60635 | v_60639;
assign v_60642 = v_60609 | v_60641;
assign v_60644 = v_60607 | v_60643;
assign v_60646 = v_60641 | v_60645;
assign v_60648 = v_60606 | v_60647;
assign v_60650 = v_60604 | v_60649;
assign v_60652 = v_60647 | v_60651;
assign v_60654 = v_60603 | v_60653;
assign v_60656 = v_60601 | v_60655;
assign v_60658 = v_60653 | v_60657;
assign v_60660 = v_60600 | v_60659;
assign v_60662 = v_60598 | v_60661;
assign v_60664 = v_60659 | v_60663;
assign v_60666 = v_60597 | v_60665;
assign v_60668 = v_60595 | v_60667;
assign v_60670 = v_60665 | v_60669;
assign v_60672 = v_60594 | v_60671;
assign v_60674 = v_60592 | v_60673;
assign v_60676 = v_60671 | v_60675;
assign v_60678 = v_60591 | v_60677;
assign v_60680 = v_60589 | v_60679;
assign v_60682 = v_60677 | v_60681;
assign v_60684 = v_60588 | v_60683;
assign v_60686 = v_60586 | v_60685;
assign v_60688 = v_60683 | v_60687;
assign v_60690 = v_60585 | v_60689;
assign v_60692 = v_60583 | v_60691;
assign v_60694 = v_60689 | v_60693;
assign v_60696 = v_60582 | v_60695;
assign v_60698 = v_60580 | v_60697;
assign v_60700 = v_60695 | v_60699;
assign v_60702 = v_60579 | v_60701;
assign v_60704 = v_60577 | v_60703;
assign v_60706 = v_60701 | v_60705;
assign v_60708 = v_60576 | v_60707;
assign v_60710 = v_60574 | v_60709;
assign v_60712 = v_60707 | v_60711;
assign v_60714 = v_60573 | v_60713;
assign v_60716 = v_60571 | v_60715;
assign v_60718 = v_60713 | v_60717;
assign v_60721 = ~v_60570 | v_60720;
assign v_60728 = v_60618 | v_60727;
assign v_60731 = v_60729 | v_60730;
assign v_60733 = v_60615 | v_60732;
assign v_60736 = v_60734 | v_60735;
assign v_60738 = v_60612 | v_60737;
assign v_60741 = v_60739 | v_60740;
assign v_60743 = v_60609 | v_60742;
assign v_60746 = v_60744 | v_60745;
assign v_60748 = v_60606 | v_60747;
assign v_60751 = v_60749 | v_60750;
assign v_60753 = v_60603 | v_60752;
assign v_60756 = v_60754 | v_60755;
assign v_60758 = v_60600 | v_60757;
assign v_60761 = v_60759 | v_60760;
assign v_60763 = v_60597 | v_60762;
assign v_60766 = v_60764 | v_60765;
assign v_60768 = v_60594 | v_60767;
assign v_60771 = v_60769 | v_60770;
assign v_60773 = v_60591 | v_60772;
assign v_60776 = v_60774 | v_60775;
assign v_60778 = v_60588 | v_60777;
assign v_60781 = v_60779 | v_60780;
assign v_60783 = v_60585 | v_60782;
assign v_60786 = v_60784 | v_60785;
assign v_60788 = v_60582 | v_60787;
assign v_60791 = v_60789 | v_60790;
assign v_60793 = v_60579 | v_60792;
assign v_60796 = v_60794 | v_60795;
assign v_60798 = v_60576 | v_60797;
assign v_60801 = v_60799 | v_60800;
assign v_60803 = v_60573 | v_60802;
assign v_60806 = v_60804 | v_60805;
assign v_60808 = v_60570 | v_60807;
assign v_60811 = v_60569 | v_60810;
assign v_60865 = v_60862 | v_60864;
assign v_60867 = v_60861 | v_60866;
assign v_60869 = v_60859 | v_60868;
assign v_60871 = v_60866 | v_60870;
assign v_60873 = v_60858 | v_60872;
assign v_60875 = v_60856 | v_60874;
assign v_60877 = v_60872 | v_60876;
assign v_60879 = v_60855 | v_60878;
assign v_60881 = v_60853 | v_60880;
assign v_60883 = v_60878 | v_60882;
assign v_60885 = v_60852 | v_60884;
assign v_60887 = v_60850 | v_60886;
assign v_60889 = v_60884 | v_60888;
assign v_60891 = v_60849 | v_60890;
assign v_60893 = v_60847 | v_60892;
assign v_60895 = v_60890 | v_60894;
assign v_60897 = v_60846 | v_60896;
assign v_60899 = v_60844 | v_60898;
assign v_60901 = v_60896 | v_60900;
assign v_60903 = v_60843 | v_60902;
assign v_60905 = v_60841 | v_60904;
assign v_60907 = v_60902 | v_60906;
assign v_60909 = v_60840 | v_60908;
assign v_60911 = v_60838 | v_60910;
assign v_60913 = v_60908 | v_60912;
assign v_60915 = v_60837 | v_60914;
assign v_60917 = v_60835 | v_60916;
assign v_60919 = v_60914 | v_60918;
assign v_60921 = v_60834 | v_60920;
assign v_60923 = v_60832 | v_60922;
assign v_60925 = v_60920 | v_60924;
assign v_60927 = v_60831 | v_60926;
assign v_60929 = v_60829 | v_60928;
assign v_60931 = v_60926 | v_60930;
assign v_60933 = v_60828 | v_60932;
assign v_60935 = v_60826 | v_60934;
assign v_60937 = v_60932 | v_60936;
assign v_60939 = v_60825 | v_60938;
assign v_60941 = v_60823 | v_60940;
assign v_60943 = v_60938 | v_60942;
assign v_60945 = v_60822 | v_60944;
assign v_60947 = v_60820 | v_60946;
assign v_60949 = v_60944 | v_60948;
assign v_60951 = v_60819 | v_60950;
assign v_60953 = v_60817 | v_60952;
assign v_60955 = v_60950 | v_60954;
assign v_60957 = v_60816 | v_60956;
assign v_60959 = v_60814 | v_60958;
assign v_60961 = v_60956 | v_60960;
assign v_60964 = ~v_60813 | v_60963;
assign v_60971 = v_60861 | v_60970;
assign v_60974 = v_60972 | v_60973;
assign v_60976 = v_60858 | v_60975;
assign v_60979 = v_60977 | v_60978;
assign v_60981 = v_60855 | v_60980;
assign v_60984 = v_60982 | v_60983;
assign v_60986 = v_60852 | v_60985;
assign v_60989 = v_60987 | v_60988;
assign v_60991 = v_60849 | v_60990;
assign v_60994 = v_60992 | v_60993;
assign v_60996 = v_60846 | v_60995;
assign v_60999 = v_60997 | v_60998;
assign v_61001 = v_60843 | v_61000;
assign v_61004 = v_61002 | v_61003;
assign v_61006 = v_60840 | v_61005;
assign v_61009 = v_61007 | v_61008;
assign v_61011 = v_60837 | v_61010;
assign v_61014 = v_61012 | v_61013;
assign v_61016 = v_60834 | v_61015;
assign v_61019 = v_61017 | v_61018;
assign v_61021 = v_60831 | v_61020;
assign v_61024 = v_61022 | v_61023;
assign v_61026 = v_60828 | v_61025;
assign v_61029 = v_61027 | v_61028;
assign v_61031 = v_60825 | v_61030;
assign v_61034 = v_61032 | v_61033;
assign v_61036 = v_60822 | v_61035;
assign v_61039 = v_61037 | v_61038;
assign v_61041 = v_60819 | v_61040;
assign v_61044 = v_61042 | v_61043;
assign v_61046 = v_60816 | v_61045;
assign v_61049 = v_61047 | v_61048;
assign v_61051 = v_60813 | v_61050;
assign v_61054 = v_60812 | v_61053;
assign v_61108 = v_61105 | v_61107;
assign v_61110 = v_61104 | v_61109;
assign v_61112 = v_61102 | v_61111;
assign v_61114 = v_61109 | v_61113;
assign v_61116 = v_61101 | v_61115;
assign v_61118 = v_61099 | v_61117;
assign v_61120 = v_61115 | v_61119;
assign v_61122 = v_61098 | v_61121;
assign v_61124 = v_61096 | v_61123;
assign v_61126 = v_61121 | v_61125;
assign v_61128 = v_61095 | v_61127;
assign v_61130 = v_61093 | v_61129;
assign v_61132 = v_61127 | v_61131;
assign v_61134 = v_61092 | v_61133;
assign v_61136 = v_61090 | v_61135;
assign v_61138 = v_61133 | v_61137;
assign v_61140 = v_61089 | v_61139;
assign v_61142 = v_61087 | v_61141;
assign v_61144 = v_61139 | v_61143;
assign v_61146 = v_61086 | v_61145;
assign v_61148 = v_61084 | v_61147;
assign v_61150 = v_61145 | v_61149;
assign v_61152 = v_61083 | v_61151;
assign v_61154 = v_61081 | v_61153;
assign v_61156 = v_61151 | v_61155;
assign v_61158 = v_61080 | v_61157;
assign v_61160 = v_61078 | v_61159;
assign v_61162 = v_61157 | v_61161;
assign v_61164 = v_61077 | v_61163;
assign v_61166 = v_61075 | v_61165;
assign v_61168 = v_61163 | v_61167;
assign v_61170 = v_61074 | v_61169;
assign v_61172 = v_61072 | v_61171;
assign v_61174 = v_61169 | v_61173;
assign v_61176 = v_61071 | v_61175;
assign v_61178 = v_61069 | v_61177;
assign v_61180 = v_61175 | v_61179;
assign v_61182 = v_61068 | v_61181;
assign v_61184 = v_61066 | v_61183;
assign v_61186 = v_61181 | v_61185;
assign v_61188 = v_61065 | v_61187;
assign v_61190 = v_61063 | v_61189;
assign v_61192 = v_61187 | v_61191;
assign v_61194 = v_61062 | v_61193;
assign v_61196 = v_61060 | v_61195;
assign v_61198 = v_61193 | v_61197;
assign v_61200 = v_61059 | v_61199;
assign v_61202 = v_61057 | v_61201;
assign v_61204 = v_61199 | v_61203;
assign v_61207 = ~v_61056 | v_61206;
assign v_61214 = v_61104 | v_61213;
assign v_61217 = v_61215 | v_61216;
assign v_61219 = v_61101 | v_61218;
assign v_61222 = v_61220 | v_61221;
assign v_61224 = v_61098 | v_61223;
assign v_61227 = v_61225 | v_61226;
assign v_61229 = v_61095 | v_61228;
assign v_61232 = v_61230 | v_61231;
assign v_61234 = v_61092 | v_61233;
assign v_61237 = v_61235 | v_61236;
assign v_61239 = v_61089 | v_61238;
assign v_61242 = v_61240 | v_61241;
assign v_61244 = v_61086 | v_61243;
assign v_61247 = v_61245 | v_61246;
assign v_61249 = v_61083 | v_61248;
assign v_61252 = v_61250 | v_61251;
assign v_61254 = v_61080 | v_61253;
assign v_61257 = v_61255 | v_61256;
assign v_61259 = v_61077 | v_61258;
assign v_61262 = v_61260 | v_61261;
assign v_61264 = v_61074 | v_61263;
assign v_61267 = v_61265 | v_61266;
assign v_61269 = v_61071 | v_61268;
assign v_61272 = v_61270 | v_61271;
assign v_61274 = v_61068 | v_61273;
assign v_61277 = v_61275 | v_61276;
assign v_61279 = v_61065 | v_61278;
assign v_61282 = v_61280 | v_61281;
assign v_61284 = v_61062 | v_61283;
assign v_61287 = v_61285 | v_61286;
assign v_61289 = v_61059 | v_61288;
assign v_61292 = v_61290 | v_61291;
assign v_61294 = v_61056 | v_61293;
assign v_61297 = v_61055 | v_61296;
assign v_61351 = v_61348 | v_61350;
assign v_61353 = v_61347 | v_61352;
assign v_61355 = v_61345 | v_61354;
assign v_61357 = v_61352 | v_61356;
assign v_61359 = v_61344 | v_61358;
assign v_61361 = v_61342 | v_61360;
assign v_61363 = v_61358 | v_61362;
assign v_61365 = v_61341 | v_61364;
assign v_61367 = v_61339 | v_61366;
assign v_61369 = v_61364 | v_61368;
assign v_61371 = v_61338 | v_61370;
assign v_61373 = v_61336 | v_61372;
assign v_61375 = v_61370 | v_61374;
assign v_61377 = v_61335 | v_61376;
assign v_61379 = v_61333 | v_61378;
assign v_61381 = v_61376 | v_61380;
assign v_61383 = v_61332 | v_61382;
assign v_61385 = v_61330 | v_61384;
assign v_61387 = v_61382 | v_61386;
assign v_61389 = v_61329 | v_61388;
assign v_61391 = v_61327 | v_61390;
assign v_61393 = v_61388 | v_61392;
assign v_61395 = v_61326 | v_61394;
assign v_61397 = v_61324 | v_61396;
assign v_61399 = v_61394 | v_61398;
assign v_61401 = v_61323 | v_61400;
assign v_61403 = v_61321 | v_61402;
assign v_61405 = v_61400 | v_61404;
assign v_61407 = v_61320 | v_61406;
assign v_61409 = v_61318 | v_61408;
assign v_61411 = v_61406 | v_61410;
assign v_61413 = v_61317 | v_61412;
assign v_61415 = v_61315 | v_61414;
assign v_61417 = v_61412 | v_61416;
assign v_61419 = v_61314 | v_61418;
assign v_61421 = v_61312 | v_61420;
assign v_61423 = v_61418 | v_61422;
assign v_61425 = v_61311 | v_61424;
assign v_61427 = v_61309 | v_61426;
assign v_61429 = v_61424 | v_61428;
assign v_61431 = v_61308 | v_61430;
assign v_61433 = v_61306 | v_61432;
assign v_61435 = v_61430 | v_61434;
assign v_61437 = v_61305 | v_61436;
assign v_61439 = v_61303 | v_61438;
assign v_61441 = v_61436 | v_61440;
assign v_61443 = v_61302 | v_61442;
assign v_61445 = v_61300 | v_61444;
assign v_61447 = v_61442 | v_61446;
assign v_61450 = ~v_61299 | v_61449;
assign v_61457 = v_61347 | v_61456;
assign v_61460 = v_61458 | v_61459;
assign v_61462 = v_61344 | v_61461;
assign v_61465 = v_61463 | v_61464;
assign v_61467 = v_61341 | v_61466;
assign v_61470 = v_61468 | v_61469;
assign v_61472 = v_61338 | v_61471;
assign v_61475 = v_61473 | v_61474;
assign v_61477 = v_61335 | v_61476;
assign v_61480 = v_61478 | v_61479;
assign v_61482 = v_61332 | v_61481;
assign v_61485 = v_61483 | v_61484;
assign v_61487 = v_61329 | v_61486;
assign v_61490 = v_61488 | v_61489;
assign v_61492 = v_61326 | v_61491;
assign v_61495 = v_61493 | v_61494;
assign v_61497 = v_61323 | v_61496;
assign v_61500 = v_61498 | v_61499;
assign v_61502 = v_61320 | v_61501;
assign v_61505 = v_61503 | v_61504;
assign v_61507 = v_61317 | v_61506;
assign v_61510 = v_61508 | v_61509;
assign v_61512 = v_61314 | v_61511;
assign v_61515 = v_61513 | v_61514;
assign v_61517 = v_61311 | v_61516;
assign v_61520 = v_61518 | v_61519;
assign v_61522 = v_61308 | v_61521;
assign v_61525 = v_61523 | v_61524;
assign v_61527 = v_61305 | v_61526;
assign v_61530 = v_61528 | v_61529;
assign v_61532 = v_61302 | v_61531;
assign v_61535 = v_61533 | v_61534;
assign v_61537 = v_61299 | v_61536;
assign v_61540 = v_61298 | v_61539;
assign v_61594 = v_61591 | v_61593;
assign v_61596 = v_61590 | v_61595;
assign v_61598 = v_61588 | v_61597;
assign v_61600 = v_61595 | v_61599;
assign v_61602 = v_61587 | v_61601;
assign v_61604 = v_61585 | v_61603;
assign v_61606 = v_61601 | v_61605;
assign v_61608 = v_61584 | v_61607;
assign v_61610 = v_61582 | v_61609;
assign v_61612 = v_61607 | v_61611;
assign v_61614 = v_61581 | v_61613;
assign v_61616 = v_61579 | v_61615;
assign v_61618 = v_61613 | v_61617;
assign v_61620 = v_61578 | v_61619;
assign v_61622 = v_61576 | v_61621;
assign v_61624 = v_61619 | v_61623;
assign v_61626 = v_61575 | v_61625;
assign v_61628 = v_61573 | v_61627;
assign v_61630 = v_61625 | v_61629;
assign v_61632 = v_61572 | v_61631;
assign v_61634 = v_61570 | v_61633;
assign v_61636 = v_61631 | v_61635;
assign v_61638 = v_61569 | v_61637;
assign v_61640 = v_61567 | v_61639;
assign v_61642 = v_61637 | v_61641;
assign v_61644 = v_61566 | v_61643;
assign v_61646 = v_61564 | v_61645;
assign v_61648 = v_61643 | v_61647;
assign v_61650 = v_61563 | v_61649;
assign v_61652 = v_61561 | v_61651;
assign v_61654 = v_61649 | v_61653;
assign v_61656 = v_61560 | v_61655;
assign v_61658 = v_61558 | v_61657;
assign v_61660 = v_61655 | v_61659;
assign v_61662 = v_61557 | v_61661;
assign v_61664 = v_61555 | v_61663;
assign v_61666 = v_61661 | v_61665;
assign v_61668 = v_61554 | v_61667;
assign v_61670 = v_61552 | v_61669;
assign v_61672 = v_61667 | v_61671;
assign v_61674 = v_61551 | v_61673;
assign v_61676 = v_61549 | v_61675;
assign v_61678 = v_61673 | v_61677;
assign v_61680 = v_61548 | v_61679;
assign v_61682 = v_61546 | v_61681;
assign v_61684 = v_61679 | v_61683;
assign v_61686 = v_61545 | v_61685;
assign v_61688 = v_61543 | v_61687;
assign v_61690 = v_61685 | v_61689;
assign v_61693 = ~v_61542 | v_61692;
assign v_61700 = v_61590 | v_61699;
assign v_61703 = v_61701 | v_61702;
assign v_61705 = v_61587 | v_61704;
assign v_61708 = v_61706 | v_61707;
assign v_61710 = v_61584 | v_61709;
assign v_61713 = v_61711 | v_61712;
assign v_61715 = v_61581 | v_61714;
assign v_61718 = v_61716 | v_61717;
assign v_61720 = v_61578 | v_61719;
assign v_61723 = v_61721 | v_61722;
assign v_61725 = v_61575 | v_61724;
assign v_61728 = v_61726 | v_61727;
assign v_61730 = v_61572 | v_61729;
assign v_61733 = v_61731 | v_61732;
assign v_61735 = v_61569 | v_61734;
assign v_61738 = v_61736 | v_61737;
assign v_61740 = v_61566 | v_61739;
assign v_61743 = v_61741 | v_61742;
assign v_61745 = v_61563 | v_61744;
assign v_61748 = v_61746 | v_61747;
assign v_61750 = v_61560 | v_61749;
assign v_61753 = v_61751 | v_61752;
assign v_61755 = v_61557 | v_61754;
assign v_61758 = v_61756 | v_61757;
assign v_61760 = v_61554 | v_61759;
assign v_61763 = v_61761 | v_61762;
assign v_61765 = v_61551 | v_61764;
assign v_61768 = v_61766 | v_61767;
assign v_61770 = v_61548 | v_61769;
assign v_61773 = v_61771 | v_61772;
assign v_61775 = v_61545 | v_61774;
assign v_61778 = v_61776 | v_61777;
assign v_61780 = v_61542 | v_61779;
assign v_61783 = v_61541 | v_61782;
assign v_61837 = v_61834 | v_61836;
assign v_61839 = v_61833 | v_61838;
assign v_61841 = v_61831 | v_61840;
assign v_61843 = v_61838 | v_61842;
assign v_61845 = v_61830 | v_61844;
assign v_61847 = v_61828 | v_61846;
assign v_61849 = v_61844 | v_61848;
assign v_61851 = v_61827 | v_61850;
assign v_61853 = v_61825 | v_61852;
assign v_61855 = v_61850 | v_61854;
assign v_61857 = v_61824 | v_61856;
assign v_61859 = v_61822 | v_61858;
assign v_61861 = v_61856 | v_61860;
assign v_61863 = v_61821 | v_61862;
assign v_61865 = v_61819 | v_61864;
assign v_61867 = v_61862 | v_61866;
assign v_61869 = v_61818 | v_61868;
assign v_61871 = v_61816 | v_61870;
assign v_61873 = v_61868 | v_61872;
assign v_61875 = v_61815 | v_61874;
assign v_61877 = v_61813 | v_61876;
assign v_61879 = v_61874 | v_61878;
assign v_61881 = v_61812 | v_61880;
assign v_61883 = v_61810 | v_61882;
assign v_61885 = v_61880 | v_61884;
assign v_61887 = v_61809 | v_61886;
assign v_61889 = v_61807 | v_61888;
assign v_61891 = v_61886 | v_61890;
assign v_61893 = v_61806 | v_61892;
assign v_61895 = v_61804 | v_61894;
assign v_61897 = v_61892 | v_61896;
assign v_61899 = v_61803 | v_61898;
assign v_61901 = v_61801 | v_61900;
assign v_61903 = v_61898 | v_61902;
assign v_61905 = v_61800 | v_61904;
assign v_61907 = v_61798 | v_61906;
assign v_61909 = v_61904 | v_61908;
assign v_61911 = v_61797 | v_61910;
assign v_61913 = v_61795 | v_61912;
assign v_61915 = v_61910 | v_61914;
assign v_61917 = v_61794 | v_61916;
assign v_61919 = v_61792 | v_61918;
assign v_61921 = v_61916 | v_61920;
assign v_61923 = v_61791 | v_61922;
assign v_61925 = v_61789 | v_61924;
assign v_61927 = v_61922 | v_61926;
assign v_61929 = v_61788 | v_61928;
assign v_61931 = v_61786 | v_61930;
assign v_61933 = v_61928 | v_61932;
assign v_61936 = ~v_61785 | v_61935;
assign v_61943 = v_61833 | v_61942;
assign v_61946 = v_61944 | v_61945;
assign v_61948 = v_61830 | v_61947;
assign v_61951 = v_61949 | v_61950;
assign v_61953 = v_61827 | v_61952;
assign v_61956 = v_61954 | v_61955;
assign v_61958 = v_61824 | v_61957;
assign v_61961 = v_61959 | v_61960;
assign v_61963 = v_61821 | v_61962;
assign v_61966 = v_61964 | v_61965;
assign v_61968 = v_61818 | v_61967;
assign v_61971 = v_61969 | v_61970;
assign v_61973 = v_61815 | v_61972;
assign v_61976 = v_61974 | v_61975;
assign v_61978 = v_61812 | v_61977;
assign v_61981 = v_61979 | v_61980;
assign v_61983 = v_61809 | v_61982;
assign v_61986 = v_61984 | v_61985;
assign v_61988 = v_61806 | v_61987;
assign v_61991 = v_61989 | v_61990;
assign v_61993 = v_61803 | v_61992;
assign v_61996 = v_61994 | v_61995;
assign v_61998 = v_61800 | v_61997;
assign v_62001 = v_61999 | v_62000;
assign v_62003 = v_61797 | v_62002;
assign v_62006 = v_62004 | v_62005;
assign v_62008 = v_61794 | v_62007;
assign v_62011 = v_62009 | v_62010;
assign v_62013 = v_61791 | v_62012;
assign v_62016 = v_62014 | v_62015;
assign v_62018 = v_61788 | v_62017;
assign v_62021 = v_62019 | v_62020;
assign v_62023 = v_61785 | v_62022;
assign v_62026 = v_61784 | v_62025;
assign v_62080 = v_62077 | v_62079;
assign v_62082 = v_62076 | v_62081;
assign v_62084 = v_62074 | v_62083;
assign v_62086 = v_62081 | v_62085;
assign v_62088 = v_62073 | v_62087;
assign v_62090 = v_62071 | v_62089;
assign v_62092 = v_62087 | v_62091;
assign v_62094 = v_62070 | v_62093;
assign v_62096 = v_62068 | v_62095;
assign v_62098 = v_62093 | v_62097;
assign v_62100 = v_62067 | v_62099;
assign v_62102 = v_62065 | v_62101;
assign v_62104 = v_62099 | v_62103;
assign v_62106 = v_62064 | v_62105;
assign v_62108 = v_62062 | v_62107;
assign v_62110 = v_62105 | v_62109;
assign v_62112 = v_62061 | v_62111;
assign v_62114 = v_62059 | v_62113;
assign v_62116 = v_62111 | v_62115;
assign v_62118 = v_62058 | v_62117;
assign v_62120 = v_62056 | v_62119;
assign v_62122 = v_62117 | v_62121;
assign v_62124 = v_62055 | v_62123;
assign v_62126 = v_62053 | v_62125;
assign v_62128 = v_62123 | v_62127;
assign v_62130 = v_62052 | v_62129;
assign v_62132 = v_62050 | v_62131;
assign v_62134 = v_62129 | v_62133;
assign v_62136 = v_62049 | v_62135;
assign v_62138 = v_62047 | v_62137;
assign v_62140 = v_62135 | v_62139;
assign v_62142 = v_62046 | v_62141;
assign v_62144 = v_62044 | v_62143;
assign v_62146 = v_62141 | v_62145;
assign v_62148 = v_62043 | v_62147;
assign v_62150 = v_62041 | v_62149;
assign v_62152 = v_62147 | v_62151;
assign v_62154 = v_62040 | v_62153;
assign v_62156 = v_62038 | v_62155;
assign v_62158 = v_62153 | v_62157;
assign v_62160 = v_62037 | v_62159;
assign v_62162 = v_62035 | v_62161;
assign v_62164 = v_62159 | v_62163;
assign v_62166 = v_62034 | v_62165;
assign v_62168 = v_62032 | v_62167;
assign v_62170 = v_62165 | v_62169;
assign v_62172 = v_62031 | v_62171;
assign v_62174 = v_62029 | v_62173;
assign v_62176 = v_62171 | v_62175;
assign v_62179 = ~v_62028 | v_62178;
assign v_62186 = v_62076 | v_62185;
assign v_62189 = v_62187 | v_62188;
assign v_62191 = v_62073 | v_62190;
assign v_62194 = v_62192 | v_62193;
assign v_62196 = v_62070 | v_62195;
assign v_62199 = v_62197 | v_62198;
assign v_62201 = v_62067 | v_62200;
assign v_62204 = v_62202 | v_62203;
assign v_62206 = v_62064 | v_62205;
assign v_62209 = v_62207 | v_62208;
assign v_62211 = v_62061 | v_62210;
assign v_62214 = v_62212 | v_62213;
assign v_62216 = v_62058 | v_62215;
assign v_62219 = v_62217 | v_62218;
assign v_62221 = v_62055 | v_62220;
assign v_62224 = v_62222 | v_62223;
assign v_62226 = v_62052 | v_62225;
assign v_62229 = v_62227 | v_62228;
assign v_62231 = v_62049 | v_62230;
assign v_62234 = v_62232 | v_62233;
assign v_62236 = v_62046 | v_62235;
assign v_62239 = v_62237 | v_62238;
assign v_62241 = v_62043 | v_62240;
assign v_62244 = v_62242 | v_62243;
assign v_62246 = v_62040 | v_62245;
assign v_62249 = v_62247 | v_62248;
assign v_62251 = v_62037 | v_62250;
assign v_62254 = v_62252 | v_62253;
assign v_62256 = v_62034 | v_62255;
assign v_62259 = v_62257 | v_62258;
assign v_62261 = v_62031 | v_62260;
assign v_62264 = v_62262 | v_62263;
assign v_62266 = v_62028 | v_62265;
assign v_62269 = v_62027 | v_62268;
assign v_62322 = v_62319 | v_62321;
assign v_62324 = v_62318 | v_62323;
assign v_62326 = v_62316 | v_62325;
assign v_62328 = v_62323 | v_62327;
assign v_62330 = v_62315 | v_62329;
assign v_62332 = v_62313 | v_62331;
assign v_62334 = v_62329 | v_62333;
assign v_62336 = v_62312 | v_62335;
assign v_62338 = v_62310 | v_62337;
assign v_62340 = v_62335 | v_62339;
assign v_62342 = v_62309 | v_62341;
assign v_62344 = v_62307 | v_62343;
assign v_62346 = v_62341 | v_62345;
assign v_62348 = v_62306 | v_62347;
assign v_62350 = v_62304 | v_62349;
assign v_62352 = v_62347 | v_62351;
assign v_62354 = v_62303 | v_62353;
assign v_62356 = v_62301 | v_62355;
assign v_62358 = v_62353 | v_62357;
assign v_62360 = v_62300 | v_62359;
assign v_62362 = v_62298 | v_62361;
assign v_62364 = v_62359 | v_62363;
assign v_62366 = v_62297 | v_62365;
assign v_62368 = v_62295 | v_62367;
assign v_62370 = v_62365 | v_62369;
assign v_62372 = v_62294 | v_62371;
assign v_62374 = v_62292 | v_62373;
assign v_62376 = v_62371 | v_62375;
assign v_62378 = v_62291 | v_62377;
assign v_62380 = v_62289 | v_62379;
assign v_62382 = v_62377 | v_62381;
assign v_62384 = v_62288 | v_62383;
assign v_62386 = v_62286 | v_62385;
assign v_62388 = v_62383 | v_62387;
assign v_62390 = v_62285 | v_62389;
assign v_62392 = v_62283 | v_62391;
assign v_62394 = v_62389 | v_62393;
assign v_62396 = v_62282 | v_62395;
assign v_62398 = v_62280 | v_62397;
assign v_62400 = v_62395 | v_62399;
assign v_62402 = v_62279 | v_62401;
assign v_62404 = v_62277 | v_62403;
assign v_62406 = v_62401 | v_62405;
assign v_62408 = v_62276 | v_62407;
assign v_62410 = v_62274 | v_62409;
assign v_62412 = v_62407 | v_62411;
assign v_62414 = v_62273 | v_62413;
assign v_62416 = v_62271 | v_62415;
assign v_62418 = v_62413 | v_62417;
assign v_62422 = v_62419 | v_62421;
assign v_62429 = v_62318 | v_62428;
assign v_62432 = v_62430 | v_62431;
assign v_62434 = v_62315 | v_62433;
assign v_62437 = v_62435 | v_62436;
assign v_62439 = v_62312 | v_62438;
assign v_62442 = v_62440 | v_62441;
assign v_62444 = v_62309 | v_62443;
assign v_62447 = v_62445 | v_62446;
assign v_62449 = v_62306 | v_62448;
assign v_62452 = v_62450 | v_62451;
assign v_62454 = v_62303 | v_62453;
assign v_62457 = v_62455 | v_62456;
assign v_62459 = v_62300 | v_62458;
assign v_62462 = v_62460 | v_62461;
assign v_62464 = v_62297 | v_62463;
assign v_62467 = v_62465 | v_62466;
assign v_62469 = v_62294 | v_62468;
assign v_62472 = v_62470 | v_62471;
assign v_62474 = v_62291 | v_62473;
assign v_62477 = v_62475 | v_62476;
assign v_62479 = v_62288 | v_62478;
assign v_62482 = v_62480 | v_62481;
assign v_62484 = v_62285 | v_62483;
assign v_62487 = v_62485 | v_62486;
assign v_62489 = v_62282 | v_62488;
assign v_62492 = v_62490 | v_62491;
assign v_62494 = v_62279 | v_62493;
assign v_62497 = v_62495 | v_62496;
assign v_62499 = v_62276 | v_62498;
assign v_62502 = v_62500 | v_62501;
assign v_62504 = v_62273 | v_62503;
assign v_62507 = v_62505 | v_62506;
assign v_62509 = v_62507 | v_62508;
assign v_62512 = v_62270 | v_62511;
assign v_62583 = v_62580 | v_62582;
assign v_62585 = v_62578 | v_62584;
assign v_62587 = v_62576 | v_62586;
assign v_62589 = v_62584 | v_62588;
assign v_62591 = v_62574 | v_62590;
assign v_62593 = v_62572 | v_62592;
assign v_62595 = v_62590 | v_62594;
assign v_62597 = v_62570 | v_62596;
assign v_62599 = v_62568 | v_62598;
assign v_62601 = v_62596 | v_62600;
assign v_62603 = v_62566 | v_62602;
assign v_62605 = v_62564 | v_62604;
assign v_62607 = v_62602 | v_62606;
assign v_62609 = v_62562 | v_62608;
assign v_62611 = v_62560 | v_62610;
assign v_62613 = v_62608 | v_62612;
assign v_62615 = v_62558 | v_62614;
assign v_62617 = v_62556 | v_62616;
assign v_62619 = v_62614 | v_62618;
assign v_62621 = v_62554 | v_62620;
assign v_62623 = v_62552 | v_62622;
assign v_62625 = v_62620 | v_62624;
assign v_62627 = v_62550 | v_62626;
assign v_62629 = v_62548 | v_62628;
assign v_62631 = v_62626 | v_62630;
assign v_62633 = v_62546 | v_62632;
assign v_62635 = v_62544 | v_62634;
assign v_62637 = v_62632 | v_62636;
assign v_62639 = v_62542 | v_62638;
assign v_62641 = v_62540 | v_62640;
assign v_62643 = v_62638 | v_62642;
assign v_62645 = v_62538 | v_62644;
assign v_62647 = v_62536 | v_62646;
assign v_62649 = v_62644 | v_62648;
assign v_62651 = v_62534 | v_62650;
assign v_62653 = v_62532 | v_62652;
assign v_62655 = v_62650 | v_62654;
assign v_62657 = v_62530 | v_62656;
assign v_62659 = v_62527 | v_62658;
assign v_62661 = v_62656 | v_62660;
assign v_62663 = v_62526 | v_62662;
assign v_62665 = v_62523 | v_62664;
assign v_62667 = v_62662 | v_62666;
assign v_62669 = v_62522 | v_62668;
assign v_62671 = v_62519 | v_62670;
assign v_62673 = v_62668 | v_62672;
assign v_62675 = v_62518 | v_62674;
assign v_62677 = v_62515 | v_62676;
assign v_62679 = v_62674 | v_62678;
assign v_62682 = ~v_62514 | v_62681;
assign v_62689 = v_62578 | v_62688;
assign v_62692 = v_62690 | v_62691;
assign v_62694 = v_62574 | v_62693;
assign v_62697 = v_62695 | v_62696;
assign v_62699 = v_62570 | v_62698;
assign v_62702 = v_62700 | v_62701;
assign v_62704 = v_62566 | v_62703;
assign v_62707 = v_62705 | v_62706;
assign v_62709 = v_62562 | v_62708;
assign v_62712 = v_62710 | v_62711;
assign v_62714 = v_62558 | v_62713;
assign v_62717 = v_62715 | v_62716;
assign v_62719 = v_62554 | v_62718;
assign v_62722 = v_62720 | v_62721;
assign v_62724 = v_62550 | v_62723;
assign v_62727 = v_62725 | v_62726;
assign v_62729 = v_62546 | v_62728;
assign v_62732 = v_62730 | v_62731;
assign v_62734 = v_62542 | v_62733;
assign v_62737 = v_62735 | v_62736;
assign v_62739 = v_62538 | v_62738;
assign v_62742 = v_62740 | v_62741;
assign v_62744 = v_62534 | v_62743;
assign v_62747 = v_62745 | v_62746;
assign v_62749 = v_62530 | v_62748;
assign v_62752 = v_62750 | v_62751;
assign v_62754 = v_62526 | v_62753;
assign v_62757 = v_62755 | v_62756;
assign v_62759 = v_62522 | v_62758;
assign v_62762 = v_62760 | v_62761;
assign v_62764 = v_62518 | v_62763;
assign v_62767 = v_62765 | v_62766;
assign v_62769 = v_62514 | v_62768;
assign v_62772 = v_62513 | v_62771;
assign v_62826 = v_62823 | v_62825;
assign v_62828 = v_62822 | v_62827;
assign v_62830 = v_62820 | v_62829;
assign v_62832 = v_62827 | v_62831;
assign v_62834 = v_62819 | v_62833;
assign v_62836 = v_62817 | v_62835;
assign v_62838 = v_62833 | v_62837;
assign v_62840 = v_62816 | v_62839;
assign v_62842 = v_62814 | v_62841;
assign v_62844 = v_62839 | v_62843;
assign v_62846 = v_62813 | v_62845;
assign v_62848 = v_62811 | v_62847;
assign v_62850 = v_62845 | v_62849;
assign v_62852 = v_62810 | v_62851;
assign v_62854 = v_62808 | v_62853;
assign v_62856 = v_62851 | v_62855;
assign v_62858 = v_62807 | v_62857;
assign v_62860 = v_62805 | v_62859;
assign v_62862 = v_62857 | v_62861;
assign v_62864 = v_62804 | v_62863;
assign v_62866 = v_62802 | v_62865;
assign v_62868 = v_62863 | v_62867;
assign v_62870 = v_62801 | v_62869;
assign v_62872 = v_62799 | v_62871;
assign v_62874 = v_62869 | v_62873;
assign v_62876 = v_62798 | v_62875;
assign v_62878 = v_62796 | v_62877;
assign v_62880 = v_62875 | v_62879;
assign v_62882 = v_62795 | v_62881;
assign v_62884 = v_62793 | v_62883;
assign v_62886 = v_62881 | v_62885;
assign v_62888 = v_62792 | v_62887;
assign v_62890 = v_62790 | v_62889;
assign v_62892 = v_62887 | v_62891;
assign v_62894 = v_62789 | v_62893;
assign v_62896 = v_62787 | v_62895;
assign v_62898 = v_62893 | v_62897;
assign v_62900 = v_62786 | v_62899;
assign v_62902 = v_62784 | v_62901;
assign v_62904 = v_62899 | v_62903;
assign v_62906 = v_62783 | v_62905;
assign v_62908 = v_62781 | v_62907;
assign v_62910 = v_62905 | v_62909;
assign v_62912 = v_62780 | v_62911;
assign v_62914 = v_62778 | v_62913;
assign v_62916 = v_62911 | v_62915;
assign v_62918 = v_62777 | v_62917;
assign v_62920 = v_62775 | v_62919;
assign v_62922 = v_62917 | v_62921;
assign v_62925 = ~v_62774 | v_62924;
assign v_62932 = v_62822 | v_62931;
assign v_62935 = v_62933 | v_62934;
assign v_62937 = v_62819 | v_62936;
assign v_62940 = v_62938 | v_62939;
assign v_62942 = v_62816 | v_62941;
assign v_62945 = v_62943 | v_62944;
assign v_62947 = v_62813 | v_62946;
assign v_62950 = v_62948 | v_62949;
assign v_62952 = v_62810 | v_62951;
assign v_62955 = v_62953 | v_62954;
assign v_62957 = v_62807 | v_62956;
assign v_62960 = v_62958 | v_62959;
assign v_62962 = v_62804 | v_62961;
assign v_62965 = v_62963 | v_62964;
assign v_62967 = v_62801 | v_62966;
assign v_62970 = v_62968 | v_62969;
assign v_62972 = v_62798 | v_62971;
assign v_62975 = v_62973 | v_62974;
assign v_62977 = v_62795 | v_62976;
assign v_62980 = v_62978 | v_62979;
assign v_62982 = v_62792 | v_62981;
assign v_62985 = v_62983 | v_62984;
assign v_62987 = v_62789 | v_62986;
assign v_62990 = v_62988 | v_62989;
assign v_62992 = v_62786 | v_62991;
assign v_62995 = v_62993 | v_62994;
assign v_62997 = v_62783 | v_62996;
assign v_63000 = v_62998 | v_62999;
assign v_63002 = v_62780 | v_63001;
assign v_63005 = v_63003 | v_63004;
assign v_63007 = v_62777 | v_63006;
assign v_63010 = v_63008 | v_63009;
assign v_63012 = v_62774 | v_63011;
assign v_63015 = v_62773 | v_63014;
assign v_63069 = v_63066 | v_63068;
assign v_63071 = v_63065 | v_63070;
assign v_63073 = v_63063 | v_63072;
assign v_63075 = v_63070 | v_63074;
assign v_63077 = v_63062 | v_63076;
assign v_63079 = v_63060 | v_63078;
assign v_63081 = v_63076 | v_63080;
assign v_63083 = v_63059 | v_63082;
assign v_63085 = v_63057 | v_63084;
assign v_63087 = v_63082 | v_63086;
assign v_63089 = v_63056 | v_63088;
assign v_63091 = v_63054 | v_63090;
assign v_63093 = v_63088 | v_63092;
assign v_63095 = v_63053 | v_63094;
assign v_63097 = v_63051 | v_63096;
assign v_63099 = v_63094 | v_63098;
assign v_63101 = v_63050 | v_63100;
assign v_63103 = v_63048 | v_63102;
assign v_63105 = v_63100 | v_63104;
assign v_63107 = v_63047 | v_63106;
assign v_63109 = v_63045 | v_63108;
assign v_63111 = v_63106 | v_63110;
assign v_63113 = v_63044 | v_63112;
assign v_63115 = v_63042 | v_63114;
assign v_63117 = v_63112 | v_63116;
assign v_63119 = v_63041 | v_63118;
assign v_63121 = v_63039 | v_63120;
assign v_63123 = v_63118 | v_63122;
assign v_63125 = v_63038 | v_63124;
assign v_63127 = v_63036 | v_63126;
assign v_63129 = v_63124 | v_63128;
assign v_63131 = v_63035 | v_63130;
assign v_63133 = v_63033 | v_63132;
assign v_63135 = v_63130 | v_63134;
assign v_63137 = v_63032 | v_63136;
assign v_63139 = v_63030 | v_63138;
assign v_63141 = v_63136 | v_63140;
assign v_63143 = v_63029 | v_63142;
assign v_63145 = v_63027 | v_63144;
assign v_63147 = v_63142 | v_63146;
assign v_63149 = v_63026 | v_63148;
assign v_63151 = v_63024 | v_63150;
assign v_63153 = v_63148 | v_63152;
assign v_63155 = v_63023 | v_63154;
assign v_63157 = v_63021 | v_63156;
assign v_63159 = v_63154 | v_63158;
assign v_63161 = v_63020 | v_63160;
assign v_63163 = v_63018 | v_63162;
assign v_63165 = v_63160 | v_63164;
assign v_63168 = ~v_63017 | v_63167;
assign v_63175 = v_63065 | v_63174;
assign v_63178 = v_63176 | v_63177;
assign v_63180 = v_63062 | v_63179;
assign v_63183 = v_63181 | v_63182;
assign v_63185 = v_63059 | v_63184;
assign v_63188 = v_63186 | v_63187;
assign v_63190 = v_63056 | v_63189;
assign v_63193 = v_63191 | v_63192;
assign v_63195 = v_63053 | v_63194;
assign v_63198 = v_63196 | v_63197;
assign v_63200 = v_63050 | v_63199;
assign v_63203 = v_63201 | v_63202;
assign v_63205 = v_63047 | v_63204;
assign v_63208 = v_63206 | v_63207;
assign v_63210 = v_63044 | v_63209;
assign v_63213 = v_63211 | v_63212;
assign v_63215 = v_63041 | v_63214;
assign v_63218 = v_63216 | v_63217;
assign v_63220 = v_63038 | v_63219;
assign v_63223 = v_63221 | v_63222;
assign v_63225 = v_63035 | v_63224;
assign v_63228 = v_63226 | v_63227;
assign v_63230 = v_63032 | v_63229;
assign v_63233 = v_63231 | v_63232;
assign v_63235 = v_63029 | v_63234;
assign v_63238 = v_63236 | v_63237;
assign v_63240 = v_63026 | v_63239;
assign v_63243 = v_63241 | v_63242;
assign v_63245 = v_63023 | v_63244;
assign v_63248 = v_63246 | v_63247;
assign v_63250 = v_63020 | v_63249;
assign v_63253 = v_63251 | v_63252;
assign v_63255 = v_63017 | v_63254;
assign v_63258 = v_63016 | v_63257;
assign v_63312 = v_63309 | v_63311;
assign v_63314 = v_63308 | v_63313;
assign v_63316 = v_63306 | v_63315;
assign v_63318 = v_63313 | v_63317;
assign v_63320 = v_63305 | v_63319;
assign v_63322 = v_63303 | v_63321;
assign v_63324 = v_63319 | v_63323;
assign v_63326 = v_63302 | v_63325;
assign v_63328 = v_63300 | v_63327;
assign v_63330 = v_63325 | v_63329;
assign v_63332 = v_63299 | v_63331;
assign v_63334 = v_63297 | v_63333;
assign v_63336 = v_63331 | v_63335;
assign v_63338 = v_63296 | v_63337;
assign v_63340 = v_63294 | v_63339;
assign v_63342 = v_63337 | v_63341;
assign v_63344 = v_63293 | v_63343;
assign v_63346 = v_63291 | v_63345;
assign v_63348 = v_63343 | v_63347;
assign v_63350 = v_63290 | v_63349;
assign v_63352 = v_63288 | v_63351;
assign v_63354 = v_63349 | v_63353;
assign v_63356 = v_63287 | v_63355;
assign v_63358 = v_63285 | v_63357;
assign v_63360 = v_63355 | v_63359;
assign v_63362 = v_63284 | v_63361;
assign v_63364 = v_63282 | v_63363;
assign v_63366 = v_63361 | v_63365;
assign v_63368 = v_63281 | v_63367;
assign v_63370 = v_63279 | v_63369;
assign v_63372 = v_63367 | v_63371;
assign v_63374 = v_63278 | v_63373;
assign v_63376 = v_63276 | v_63375;
assign v_63378 = v_63373 | v_63377;
assign v_63380 = v_63275 | v_63379;
assign v_63382 = v_63273 | v_63381;
assign v_63384 = v_63379 | v_63383;
assign v_63386 = v_63272 | v_63385;
assign v_63388 = v_63270 | v_63387;
assign v_63390 = v_63385 | v_63389;
assign v_63392 = v_63269 | v_63391;
assign v_63394 = v_63267 | v_63393;
assign v_63396 = v_63391 | v_63395;
assign v_63398 = v_63266 | v_63397;
assign v_63400 = v_63264 | v_63399;
assign v_63402 = v_63397 | v_63401;
assign v_63404 = v_63263 | v_63403;
assign v_63406 = v_63261 | v_63405;
assign v_63408 = v_63403 | v_63407;
assign v_63411 = ~v_63260 | v_63410;
assign v_63418 = v_63308 | v_63417;
assign v_63421 = v_63419 | v_63420;
assign v_63423 = v_63305 | v_63422;
assign v_63426 = v_63424 | v_63425;
assign v_63428 = v_63302 | v_63427;
assign v_63431 = v_63429 | v_63430;
assign v_63433 = v_63299 | v_63432;
assign v_63436 = v_63434 | v_63435;
assign v_63438 = v_63296 | v_63437;
assign v_63441 = v_63439 | v_63440;
assign v_63443 = v_63293 | v_63442;
assign v_63446 = v_63444 | v_63445;
assign v_63448 = v_63290 | v_63447;
assign v_63451 = v_63449 | v_63450;
assign v_63453 = v_63287 | v_63452;
assign v_63456 = v_63454 | v_63455;
assign v_63458 = v_63284 | v_63457;
assign v_63461 = v_63459 | v_63460;
assign v_63463 = v_63281 | v_63462;
assign v_63466 = v_63464 | v_63465;
assign v_63468 = v_63278 | v_63467;
assign v_63471 = v_63469 | v_63470;
assign v_63473 = v_63275 | v_63472;
assign v_63476 = v_63474 | v_63475;
assign v_63478 = v_63272 | v_63477;
assign v_63481 = v_63479 | v_63480;
assign v_63483 = v_63269 | v_63482;
assign v_63486 = v_63484 | v_63485;
assign v_63488 = v_63266 | v_63487;
assign v_63491 = v_63489 | v_63490;
assign v_63493 = v_63263 | v_63492;
assign v_63496 = v_63494 | v_63495;
assign v_63498 = v_63260 | v_63497;
assign v_63501 = v_63259 | v_63500;
assign v_63555 = v_63552 | v_63554;
assign v_63557 = v_63551 | v_63556;
assign v_63559 = v_63549 | v_63558;
assign v_63561 = v_63556 | v_63560;
assign v_63563 = v_63548 | v_63562;
assign v_63565 = v_63546 | v_63564;
assign v_63567 = v_63562 | v_63566;
assign v_63569 = v_63545 | v_63568;
assign v_63571 = v_63543 | v_63570;
assign v_63573 = v_63568 | v_63572;
assign v_63575 = v_63542 | v_63574;
assign v_63577 = v_63540 | v_63576;
assign v_63579 = v_63574 | v_63578;
assign v_63581 = v_63539 | v_63580;
assign v_63583 = v_63537 | v_63582;
assign v_63585 = v_63580 | v_63584;
assign v_63587 = v_63536 | v_63586;
assign v_63589 = v_63534 | v_63588;
assign v_63591 = v_63586 | v_63590;
assign v_63593 = v_63533 | v_63592;
assign v_63595 = v_63531 | v_63594;
assign v_63597 = v_63592 | v_63596;
assign v_63599 = v_63530 | v_63598;
assign v_63601 = v_63528 | v_63600;
assign v_63603 = v_63598 | v_63602;
assign v_63605 = v_63527 | v_63604;
assign v_63607 = v_63525 | v_63606;
assign v_63609 = v_63604 | v_63608;
assign v_63611 = v_63524 | v_63610;
assign v_63613 = v_63522 | v_63612;
assign v_63615 = v_63610 | v_63614;
assign v_63617 = v_63521 | v_63616;
assign v_63619 = v_63519 | v_63618;
assign v_63621 = v_63616 | v_63620;
assign v_63623 = v_63518 | v_63622;
assign v_63625 = v_63516 | v_63624;
assign v_63627 = v_63622 | v_63626;
assign v_63629 = v_63515 | v_63628;
assign v_63631 = v_63513 | v_63630;
assign v_63633 = v_63628 | v_63632;
assign v_63635 = v_63512 | v_63634;
assign v_63637 = v_63510 | v_63636;
assign v_63639 = v_63634 | v_63638;
assign v_63641 = v_63509 | v_63640;
assign v_63643 = v_63507 | v_63642;
assign v_63645 = v_63640 | v_63644;
assign v_63647 = v_63506 | v_63646;
assign v_63649 = v_63504 | v_63648;
assign v_63651 = v_63646 | v_63650;
assign v_63654 = ~v_63503 | v_63653;
assign v_63661 = v_63551 | v_63660;
assign v_63664 = v_63662 | v_63663;
assign v_63666 = v_63548 | v_63665;
assign v_63669 = v_63667 | v_63668;
assign v_63671 = v_63545 | v_63670;
assign v_63674 = v_63672 | v_63673;
assign v_63676 = v_63542 | v_63675;
assign v_63679 = v_63677 | v_63678;
assign v_63681 = v_63539 | v_63680;
assign v_63684 = v_63682 | v_63683;
assign v_63686 = v_63536 | v_63685;
assign v_63689 = v_63687 | v_63688;
assign v_63691 = v_63533 | v_63690;
assign v_63694 = v_63692 | v_63693;
assign v_63696 = v_63530 | v_63695;
assign v_63699 = v_63697 | v_63698;
assign v_63701 = v_63527 | v_63700;
assign v_63704 = v_63702 | v_63703;
assign v_63706 = v_63524 | v_63705;
assign v_63709 = v_63707 | v_63708;
assign v_63711 = v_63521 | v_63710;
assign v_63714 = v_63712 | v_63713;
assign v_63716 = v_63518 | v_63715;
assign v_63719 = v_63717 | v_63718;
assign v_63721 = v_63515 | v_63720;
assign v_63724 = v_63722 | v_63723;
assign v_63726 = v_63512 | v_63725;
assign v_63729 = v_63727 | v_63728;
assign v_63731 = v_63509 | v_63730;
assign v_63734 = v_63732 | v_63733;
assign v_63736 = v_63506 | v_63735;
assign v_63739 = v_63737 | v_63738;
assign v_63741 = v_63503 | v_63740;
assign v_63744 = v_63502 | v_63743;
assign v_63798 = v_63795 | v_63797;
assign v_63800 = v_63794 | v_63799;
assign v_63802 = v_63792 | v_63801;
assign v_63804 = v_63799 | v_63803;
assign v_63806 = v_63791 | v_63805;
assign v_63808 = v_63789 | v_63807;
assign v_63810 = v_63805 | v_63809;
assign v_63812 = v_63788 | v_63811;
assign v_63814 = v_63786 | v_63813;
assign v_63816 = v_63811 | v_63815;
assign v_63818 = v_63785 | v_63817;
assign v_63820 = v_63783 | v_63819;
assign v_63822 = v_63817 | v_63821;
assign v_63824 = v_63782 | v_63823;
assign v_63826 = v_63780 | v_63825;
assign v_63828 = v_63823 | v_63827;
assign v_63830 = v_63779 | v_63829;
assign v_63832 = v_63777 | v_63831;
assign v_63834 = v_63829 | v_63833;
assign v_63836 = v_63776 | v_63835;
assign v_63838 = v_63774 | v_63837;
assign v_63840 = v_63835 | v_63839;
assign v_63842 = v_63773 | v_63841;
assign v_63844 = v_63771 | v_63843;
assign v_63846 = v_63841 | v_63845;
assign v_63848 = v_63770 | v_63847;
assign v_63850 = v_63768 | v_63849;
assign v_63852 = v_63847 | v_63851;
assign v_63854 = v_63767 | v_63853;
assign v_63856 = v_63765 | v_63855;
assign v_63858 = v_63853 | v_63857;
assign v_63860 = v_63764 | v_63859;
assign v_63862 = v_63762 | v_63861;
assign v_63864 = v_63859 | v_63863;
assign v_63866 = v_63761 | v_63865;
assign v_63868 = v_63759 | v_63867;
assign v_63870 = v_63865 | v_63869;
assign v_63872 = v_63758 | v_63871;
assign v_63874 = v_63756 | v_63873;
assign v_63876 = v_63871 | v_63875;
assign v_63878 = v_63755 | v_63877;
assign v_63880 = v_63753 | v_63879;
assign v_63882 = v_63877 | v_63881;
assign v_63884 = v_63752 | v_63883;
assign v_63886 = v_63750 | v_63885;
assign v_63888 = v_63883 | v_63887;
assign v_63890 = v_63749 | v_63889;
assign v_63892 = v_63747 | v_63891;
assign v_63894 = v_63889 | v_63893;
assign v_63897 = ~v_63746 | v_63896;
assign v_63904 = v_63794 | v_63903;
assign v_63907 = v_63905 | v_63906;
assign v_63909 = v_63791 | v_63908;
assign v_63912 = v_63910 | v_63911;
assign v_63914 = v_63788 | v_63913;
assign v_63917 = v_63915 | v_63916;
assign v_63919 = v_63785 | v_63918;
assign v_63922 = v_63920 | v_63921;
assign v_63924 = v_63782 | v_63923;
assign v_63927 = v_63925 | v_63926;
assign v_63929 = v_63779 | v_63928;
assign v_63932 = v_63930 | v_63931;
assign v_63934 = v_63776 | v_63933;
assign v_63937 = v_63935 | v_63936;
assign v_63939 = v_63773 | v_63938;
assign v_63942 = v_63940 | v_63941;
assign v_63944 = v_63770 | v_63943;
assign v_63947 = v_63945 | v_63946;
assign v_63949 = v_63767 | v_63948;
assign v_63952 = v_63950 | v_63951;
assign v_63954 = v_63764 | v_63953;
assign v_63957 = v_63955 | v_63956;
assign v_63959 = v_63761 | v_63958;
assign v_63962 = v_63960 | v_63961;
assign v_63964 = v_63758 | v_63963;
assign v_63967 = v_63965 | v_63966;
assign v_63969 = v_63755 | v_63968;
assign v_63972 = v_63970 | v_63971;
assign v_63974 = v_63752 | v_63973;
assign v_63977 = v_63975 | v_63976;
assign v_63979 = v_63749 | v_63978;
assign v_63982 = v_63980 | v_63981;
assign v_63984 = v_63746 | v_63983;
assign v_63987 = v_63745 | v_63986;
assign v_64041 = v_64038 | v_64040;
assign v_64043 = v_64037 | v_64042;
assign v_64045 = v_64035 | v_64044;
assign v_64047 = v_64042 | v_64046;
assign v_64049 = v_64034 | v_64048;
assign v_64051 = v_64032 | v_64050;
assign v_64053 = v_64048 | v_64052;
assign v_64055 = v_64031 | v_64054;
assign v_64057 = v_64029 | v_64056;
assign v_64059 = v_64054 | v_64058;
assign v_64061 = v_64028 | v_64060;
assign v_64063 = v_64026 | v_64062;
assign v_64065 = v_64060 | v_64064;
assign v_64067 = v_64025 | v_64066;
assign v_64069 = v_64023 | v_64068;
assign v_64071 = v_64066 | v_64070;
assign v_64073 = v_64022 | v_64072;
assign v_64075 = v_64020 | v_64074;
assign v_64077 = v_64072 | v_64076;
assign v_64079 = v_64019 | v_64078;
assign v_64081 = v_64017 | v_64080;
assign v_64083 = v_64078 | v_64082;
assign v_64085 = v_64016 | v_64084;
assign v_64087 = v_64014 | v_64086;
assign v_64089 = v_64084 | v_64088;
assign v_64091 = v_64013 | v_64090;
assign v_64093 = v_64011 | v_64092;
assign v_64095 = v_64090 | v_64094;
assign v_64097 = v_64010 | v_64096;
assign v_64099 = v_64008 | v_64098;
assign v_64101 = v_64096 | v_64100;
assign v_64103 = v_64007 | v_64102;
assign v_64105 = v_64005 | v_64104;
assign v_64107 = v_64102 | v_64106;
assign v_64109 = v_64004 | v_64108;
assign v_64111 = v_64002 | v_64110;
assign v_64113 = v_64108 | v_64112;
assign v_64115 = v_64001 | v_64114;
assign v_64117 = v_63999 | v_64116;
assign v_64119 = v_64114 | v_64118;
assign v_64121 = v_63998 | v_64120;
assign v_64123 = v_63996 | v_64122;
assign v_64125 = v_64120 | v_64124;
assign v_64127 = v_63995 | v_64126;
assign v_64129 = v_63993 | v_64128;
assign v_64131 = v_64126 | v_64130;
assign v_64133 = v_63992 | v_64132;
assign v_64135 = v_63990 | v_64134;
assign v_64137 = v_64132 | v_64136;
assign v_64140 = ~v_63989 | v_64139;
assign v_64147 = v_64037 | v_64146;
assign v_64150 = v_64148 | v_64149;
assign v_64152 = v_64034 | v_64151;
assign v_64155 = v_64153 | v_64154;
assign v_64157 = v_64031 | v_64156;
assign v_64160 = v_64158 | v_64159;
assign v_64162 = v_64028 | v_64161;
assign v_64165 = v_64163 | v_64164;
assign v_64167 = v_64025 | v_64166;
assign v_64170 = v_64168 | v_64169;
assign v_64172 = v_64022 | v_64171;
assign v_64175 = v_64173 | v_64174;
assign v_64177 = v_64019 | v_64176;
assign v_64180 = v_64178 | v_64179;
assign v_64182 = v_64016 | v_64181;
assign v_64185 = v_64183 | v_64184;
assign v_64187 = v_64013 | v_64186;
assign v_64190 = v_64188 | v_64189;
assign v_64192 = v_64010 | v_64191;
assign v_64195 = v_64193 | v_64194;
assign v_64197 = v_64007 | v_64196;
assign v_64200 = v_64198 | v_64199;
assign v_64202 = v_64004 | v_64201;
assign v_64205 = v_64203 | v_64204;
assign v_64207 = v_64001 | v_64206;
assign v_64210 = v_64208 | v_64209;
assign v_64212 = v_63998 | v_64211;
assign v_64215 = v_64213 | v_64214;
assign v_64217 = v_63995 | v_64216;
assign v_64220 = v_64218 | v_64219;
assign v_64222 = v_63992 | v_64221;
assign v_64225 = v_64223 | v_64224;
assign v_64227 = v_63989 | v_64226;
assign v_64230 = v_63988 | v_64229;
assign v_64284 = v_64281 | v_64283;
assign v_64286 = v_64280 | v_64285;
assign v_64288 = v_64278 | v_64287;
assign v_64290 = v_64285 | v_64289;
assign v_64292 = v_64277 | v_64291;
assign v_64294 = v_64275 | v_64293;
assign v_64296 = v_64291 | v_64295;
assign v_64298 = v_64274 | v_64297;
assign v_64300 = v_64272 | v_64299;
assign v_64302 = v_64297 | v_64301;
assign v_64304 = v_64271 | v_64303;
assign v_64306 = v_64269 | v_64305;
assign v_64308 = v_64303 | v_64307;
assign v_64310 = v_64268 | v_64309;
assign v_64312 = v_64266 | v_64311;
assign v_64314 = v_64309 | v_64313;
assign v_64316 = v_64265 | v_64315;
assign v_64318 = v_64263 | v_64317;
assign v_64320 = v_64315 | v_64319;
assign v_64322 = v_64262 | v_64321;
assign v_64324 = v_64260 | v_64323;
assign v_64326 = v_64321 | v_64325;
assign v_64328 = v_64259 | v_64327;
assign v_64330 = v_64257 | v_64329;
assign v_64332 = v_64327 | v_64331;
assign v_64334 = v_64256 | v_64333;
assign v_64336 = v_64254 | v_64335;
assign v_64338 = v_64333 | v_64337;
assign v_64340 = v_64253 | v_64339;
assign v_64342 = v_64251 | v_64341;
assign v_64344 = v_64339 | v_64343;
assign v_64346 = v_64250 | v_64345;
assign v_64348 = v_64248 | v_64347;
assign v_64350 = v_64345 | v_64349;
assign v_64352 = v_64247 | v_64351;
assign v_64354 = v_64245 | v_64353;
assign v_64356 = v_64351 | v_64355;
assign v_64358 = v_64244 | v_64357;
assign v_64360 = v_64242 | v_64359;
assign v_64362 = v_64357 | v_64361;
assign v_64364 = v_64241 | v_64363;
assign v_64366 = v_64239 | v_64365;
assign v_64368 = v_64363 | v_64367;
assign v_64370 = v_64238 | v_64369;
assign v_64372 = v_64236 | v_64371;
assign v_64374 = v_64369 | v_64373;
assign v_64376 = v_64235 | v_64375;
assign v_64378 = v_64233 | v_64377;
assign v_64380 = v_64375 | v_64379;
assign v_64383 = ~v_64232 | v_64382;
assign v_64390 = v_64280 | v_64389;
assign v_64393 = v_64391 | v_64392;
assign v_64395 = v_64277 | v_64394;
assign v_64398 = v_64396 | v_64397;
assign v_64400 = v_64274 | v_64399;
assign v_64403 = v_64401 | v_64402;
assign v_64405 = v_64271 | v_64404;
assign v_64408 = v_64406 | v_64407;
assign v_64410 = v_64268 | v_64409;
assign v_64413 = v_64411 | v_64412;
assign v_64415 = v_64265 | v_64414;
assign v_64418 = v_64416 | v_64417;
assign v_64420 = v_64262 | v_64419;
assign v_64423 = v_64421 | v_64422;
assign v_64425 = v_64259 | v_64424;
assign v_64428 = v_64426 | v_64427;
assign v_64430 = v_64256 | v_64429;
assign v_64433 = v_64431 | v_64432;
assign v_64435 = v_64253 | v_64434;
assign v_64438 = v_64436 | v_64437;
assign v_64440 = v_64250 | v_64439;
assign v_64443 = v_64441 | v_64442;
assign v_64445 = v_64247 | v_64444;
assign v_64448 = v_64446 | v_64447;
assign v_64450 = v_64244 | v_64449;
assign v_64453 = v_64451 | v_64452;
assign v_64455 = v_64241 | v_64454;
assign v_64458 = v_64456 | v_64457;
assign v_64460 = v_64238 | v_64459;
assign v_64463 = v_64461 | v_64462;
assign v_64465 = v_64235 | v_64464;
assign v_64468 = v_64466 | v_64467;
assign v_64470 = v_64232 | v_64469;
assign v_64473 = v_64231 | v_64472;
assign v_64527 = v_64524 | v_64526;
assign v_64529 = v_64523 | v_64528;
assign v_64531 = v_64521 | v_64530;
assign v_64533 = v_64528 | v_64532;
assign v_64535 = v_64520 | v_64534;
assign v_64537 = v_64518 | v_64536;
assign v_64539 = v_64534 | v_64538;
assign v_64541 = v_64517 | v_64540;
assign v_64543 = v_64515 | v_64542;
assign v_64545 = v_64540 | v_64544;
assign v_64547 = v_64514 | v_64546;
assign v_64549 = v_64512 | v_64548;
assign v_64551 = v_64546 | v_64550;
assign v_64553 = v_64511 | v_64552;
assign v_64555 = v_64509 | v_64554;
assign v_64557 = v_64552 | v_64556;
assign v_64559 = v_64508 | v_64558;
assign v_64561 = v_64506 | v_64560;
assign v_64563 = v_64558 | v_64562;
assign v_64565 = v_64505 | v_64564;
assign v_64567 = v_64503 | v_64566;
assign v_64569 = v_64564 | v_64568;
assign v_64571 = v_64502 | v_64570;
assign v_64573 = v_64500 | v_64572;
assign v_64575 = v_64570 | v_64574;
assign v_64577 = v_64499 | v_64576;
assign v_64579 = v_64497 | v_64578;
assign v_64581 = v_64576 | v_64580;
assign v_64583 = v_64496 | v_64582;
assign v_64585 = v_64494 | v_64584;
assign v_64587 = v_64582 | v_64586;
assign v_64589 = v_64493 | v_64588;
assign v_64591 = v_64491 | v_64590;
assign v_64593 = v_64588 | v_64592;
assign v_64595 = v_64490 | v_64594;
assign v_64597 = v_64488 | v_64596;
assign v_64599 = v_64594 | v_64598;
assign v_64601 = v_64487 | v_64600;
assign v_64603 = v_64485 | v_64602;
assign v_64605 = v_64600 | v_64604;
assign v_64607 = v_64484 | v_64606;
assign v_64609 = v_64482 | v_64608;
assign v_64611 = v_64606 | v_64610;
assign v_64613 = v_64481 | v_64612;
assign v_64615 = v_64479 | v_64614;
assign v_64617 = v_64612 | v_64616;
assign v_64619 = v_64478 | v_64618;
assign v_64621 = v_64476 | v_64620;
assign v_64623 = v_64618 | v_64622;
assign v_64626 = ~v_64475 | v_64625;
assign v_64633 = v_64523 | v_64632;
assign v_64636 = v_64634 | v_64635;
assign v_64638 = v_64520 | v_64637;
assign v_64641 = v_64639 | v_64640;
assign v_64643 = v_64517 | v_64642;
assign v_64646 = v_64644 | v_64645;
assign v_64648 = v_64514 | v_64647;
assign v_64651 = v_64649 | v_64650;
assign v_64653 = v_64511 | v_64652;
assign v_64656 = v_64654 | v_64655;
assign v_64658 = v_64508 | v_64657;
assign v_64661 = v_64659 | v_64660;
assign v_64663 = v_64505 | v_64662;
assign v_64666 = v_64664 | v_64665;
assign v_64668 = v_64502 | v_64667;
assign v_64671 = v_64669 | v_64670;
assign v_64673 = v_64499 | v_64672;
assign v_64676 = v_64674 | v_64675;
assign v_64678 = v_64496 | v_64677;
assign v_64681 = v_64679 | v_64680;
assign v_64683 = v_64493 | v_64682;
assign v_64686 = v_64684 | v_64685;
assign v_64688 = v_64490 | v_64687;
assign v_64691 = v_64689 | v_64690;
assign v_64693 = v_64487 | v_64692;
assign v_64696 = v_64694 | v_64695;
assign v_64698 = v_64484 | v_64697;
assign v_64701 = v_64699 | v_64700;
assign v_64703 = v_64481 | v_64702;
assign v_64706 = v_64704 | v_64705;
assign v_64708 = v_64478 | v_64707;
assign v_64711 = v_64709 | v_64710;
assign v_64713 = v_64475 | v_64712;
assign v_64716 = v_64474 | v_64715;
assign v_64770 = v_64767 | v_64769;
assign v_64772 = v_64766 | v_64771;
assign v_64774 = v_64764 | v_64773;
assign v_64776 = v_64771 | v_64775;
assign v_64778 = v_64763 | v_64777;
assign v_64780 = v_64761 | v_64779;
assign v_64782 = v_64777 | v_64781;
assign v_64784 = v_64760 | v_64783;
assign v_64786 = v_64758 | v_64785;
assign v_64788 = v_64783 | v_64787;
assign v_64790 = v_64757 | v_64789;
assign v_64792 = v_64755 | v_64791;
assign v_64794 = v_64789 | v_64793;
assign v_64796 = v_64754 | v_64795;
assign v_64798 = v_64752 | v_64797;
assign v_64800 = v_64795 | v_64799;
assign v_64802 = v_64751 | v_64801;
assign v_64804 = v_64749 | v_64803;
assign v_64806 = v_64801 | v_64805;
assign v_64808 = v_64748 | v_64807;
assign v_64810 = v_64746 | v_64809;
assign v_64812 = v_64807 | v_64811;
assign v_64814 = v_64745 | v_64813;
assign v_64816 = v_64743 | v_64815;
assign v_64818 = v_64813 | v_64817;
assign v_64820 = v_64742 | v_64819;
assign v_64822 = v_64740 | v_64821;
assign v_64824 = v_64819 | v_64823;
assign v_64826 = v_64739 | v_64825;
assign v_64828 = v_64737 | v_64827;
assign v_64830 = v_64825 | v_64829;
assign v_64832 = v_64736 | v_64831;
assign v_64834 = v_64734 | v_64833;
assign v_64836 = v_64831 | v_64835;
assign v_64838 = v_64733 | v_64837;
assign v_64840 = v_64731 | v_64839;
assign v_64842 = v_64837 | v_64841;
assign v_64844 = v_64730 | v_64843;
assign v_64846 = v_64728 | v_64845;
assign v_64848 = v_64843 | v_64847;
assign v_64850 = v_64727 | v_64849;
assign v_64852 = v_64725 | v_64851;
assign v_64854 = v_64849 | v_64853;
assign v_64856 = v_64724 | v_64855;
assign v_64858 = v_64722 | v_64857;
assign v_64860 = v_64855 | v_64859;
assign v_64862 = v_64721 | v_64861;
assign v_64864 = v_64719 | v_64863;
assign v_64866 = v_64861 | v_64865;
assign v_64869 = ~v_64718 | v_64868;
assign v_64876 = v_64766 | v_64875;
assign v_64879 = v_64877 | v_64878;
assign v_64881 = v_64763 | v_64880;
assign v_64884 = v_64882 | v_64883;
assign v_64886 = v_64760 | v_64885;
assign v_64889 = v_64887 | v_64888;
assign v_64891 = v_64757 | v_64890;
assign v_64894 = v_64892 | v_64893;
assign v_64896 = v_64754 | v_64895;
assign v_64899 = v_64897 | v_64898;
assign v_64901 = v_64751 | v_64900;
assign v_64904 = v_64902 | v_64903;
assign v_64906 = v_64748 | v_64905;
assign v_64909 = v_64907 | v_64908;
assign v_64911 = v_64745 | v_64910;
assign v_64914 = v_64912 | v_64913;
assign v_64916 = v_64742 | v_64915;
assign v_64919 = v_64917 | v_64918;
assign v_64921 = v_64739 | v_64920;
assign v_64924 = v_64922 | v_64923;
assign v_64926 = v_64736 | v_64925;
assign v_64929 = v_64927 | v_64928;
assign v_64931 = v_64733 | v_64930;
assign v_64934 = v_64932 | v_64933;
assign v_64936 = v_64730 | v_64935;
assign v_64939 = v_64937 | v_64938;
assign v_64941 = v_64727 | v_64940;
assign v_64944 = v_64942 | v_64943;
assign v_64946 = v_64724 | v_64945;
assign v_64949 = v_64947 | v_64948;
assign v_64951 = v_64721 | v_64950;
assign v_64954 = v_64952 | v_64953;
assign v_64956 = v_64718 | v_64955;
assign v_64959 = v_64717 | v_64958;
assign v_65013 = v_65010 | v_65012;
assign v_65015 = v_65009 | v_65014;
assign v_65017 = v_65007 | v_65016;
assign v_65019 = v_65014 | v_65018;
assign v_65021 = v_65006 | v_65020;
assign v_65023 = v_65004 | v_65022;
assign v_65025 = v_65020 | v_65024;
assign v_65027 = v_65003 | v_65026;
assign v_65029 = v_65001 | v_65028;
assign v_65031 = v_65026 | v_65030;
assign v_65033 = v_65000 | v_65032;
assign v_65035 = v_64998 | v_65034;
assign v_65037 = v_65032 | v_65036;
assign v_65039 = v_64997 | v_65038;
assign v_65041 = v_64995 | v_65040;
assign v_65043 = v_65038 | v_65042;
assign v_65045 = v_64994 | v_65044;
assign v_65047 = v_64992 | v_65046;
assign v_65049 = v_65044 | v_65048;
assign v_65051 = v_64991 | v_65050;
assign v_65053 = v_64989 | v_65052;
assign v_65055 = v_65050 | v_65054;
assign v_65057 = v_64988 | v_65056;
assign v_65059 = v_64986 | v_65058;
assign v_65061 = v_65056 | v_65060;
assign v_65063 = v_64985 | v_65062;
assign v_65065 = v_64983 | v_65064;
assign v_65067 = v_65062 | v_65066;
assign v_65069 = v_64982 | v_65068;
assign v_65071 = v_64980 | v_65070;
assign v_65073 = v_65068 | v_65072;
assign v_65075 = v_64979 | v_65074;
assign v_65077 = v_64977 | v_65076;
assign v_65079 = v_65074 | v_65078;
assign v_65081 = v_64976 | v_65080;
assign v_65083 = v_64974 | v_65082;
assign v_65085 = v_65080 | v_65084;
assign v_65087 = v_64973 | v_65086;
assign v_65089 = v_64971 | v_65088;
assign v_65091 = v_65086 | v_65090;
assign v_65093 = v_64970 | v_65092;
assign v_65095 = v_64968 | v_65094;
assign v_65097 = v_65092 | v_65096;
assign v_65099 = v_64967 | v_65098;
assign v_65101 = v_64965 | v_65100;
assign v_65103 = v_65098 | v_65102;
assign v_65105 = v_64964 | v_65104;
assign v_65107 = v_64962 | v_65106;
assign v_65109 = v_65104 | v_65108;
assign v_65112 = ~v_64961 | v_65111;
assign v_65119 = v_65009 | v_65118;
assign v_65122 = v_65120 | v_65121;
assign v_65124 = v_65006 | v_65123;
assign v_65127 = v_65125 | v_65126;
assign v_65129 = v_65003 | v_65128;
assign v_65132 = v_65130 | v_65131;
assign v_65134 = v_65000 | v_65133;
assign v_65137 = v_65135 | v_65136;
assign v_65139 = v_64997 | v_65138;
assign v_65142 = v_65140 | v_65141;
assign v_65144 = v_64994 | v_65143;
assign v_65147 = v_65145 | v_65146;
assign v_65149 = v_64991 | v_65148;
assign v_65152 = v_65150 | v_65151;
assign v_65154 = v_64988 | v_65153;
assign v_65157 = v_65155 | v_65156;
assign v_65159 = v_64985 | v_65158;
assign v_65162 = v_65160 | v_65161;
assign v_65164 = v_64982 | v_65163;
assign v_65167 = v_65165 | v_65166;
assign v_65169 = v_64979 | v_65168;
assign v_65172 = v_65170 | v_65171;
assign v_65174 = v_64976 | v_65173;
assign v_65177 = v_65175 | v_65176;
assign v_65179 = v_64973 | v_65178;
assign v_65182 = v_65180 | v_65181;
assign v_65184 = v_64970 | v_65183;
assign v_65187 = v_65185 | v_65186;
assign v_65189 = v_64967 | v_65188;
assign v_65192 = v_65190 | v_65191;
assign v_65194 = v_64964 | v_65193;
assign v_65197 = v_65195 | v_65196;
assign v_65199 = v_64961 | v_65198;
assign v_65202 = v_64960 | v_65201;
assign v_65256 = v_65253 | v_65255;
assign v_65258 = v_65252 | v_65257;
assign v_65260 = v_65250 | v_65259;
assign v_65262 = v_65257 | v_65261;
assign v_65264 = v_65249 | v_65263;
assign v_65266 = v_65247 | v_65265;
assign v_65268 = v_65263 | v_65267;
assign v_65270 = v_65246 | v_65269;
assign v_65272 = v_65244 | v_65271;
assign v_65274 = v_65269 | v_65273;
assign v_65276 = v_65243 | v_65275;
assign v_65278 = v_65241 | v_65277;
assign v_65280 = v_65275 | v_65279;
assign v_65282 = v_65240 | v_65281;
assign v_65284 = v_65238 | v_65283;
assign v_65286 = v_65281 | v_65285;
assign v_65288 = v_65237 | v_65287;
assign v_65290 = v_65235 | v_65289;
assign v_65292 = v_65287 | v_65291;
assign v_65294 = v_65234 | v_65293;
assign v_65296 = v_65232 | v_65295;
assign v_65298 = v_65293 | v_65297;
assign v_65300 = v_65231 | v_65299;
assign v_65302 = v_65229 | v_65301;
assign v_65304 = v_65299 | v_65303;
assign v_65306 = v_65228 | v_65305;
assign v_65308 = v_65226 | v_65307;
assign v_65310 = v_65305 | v_65309;
assign v_65312 = v_65225 | v_65311;
assign v_65314 = v_65223 | v_65313;
assign v_65316 = v_65311 | v_65315;
assign v_65318 = v_65222 | v_65317;
assign v_65320 = v_65220 | v_65319;
assign v_65322 = v_65317 | v_65321;
assign v_65324 = v_65219 | v_65323;
assign v_65326 = v_65217 | v_65325;
assign v_65328 = v_65323 | v_65327;
assign v_65330 = v_65216 | v_65329;
assign v_65332 = v_65214 | v_65331;
assign v_65334 = v_65329 | v_65333;
assign v_65336 = v_65213 | v_65335;
assign v_65338 = v_65211 | v_65337;
assign v_65340 = v_65335 | v_65339;
assign v_65342 = v_65210 | v_65341;
assign v_65344 = v_65208 | v_65343;
assign v_65346 = v_65341 | v_65345;
assign v_65348 = v_65207 | v_65347;
assign v_65350 = v_65205 | v_65349;
assign v_65352 = v_65347 | v_65351;
assign v_65355 = ~v_65204 | v_65354;
assign v_65362 = v_65252 | v_65361;
assign v_65365 = v_65363 | v_65364;
assign v_65367 = v_65249 | v_65366;
assign v_65370 = v_65368 | v_65369;
assign v_65372 = v_65246 | v_65371;
assign v_65375 = v_65373 | v_65374;
assign v_65377 = v_65243 | v_65376;
assign v_65380 = v_65378 | v_65379;
assign v_65382 = v_65240 | v_65381;
assign v_65385 = v_65383 | v_65384;
assign v_65387 = v_65237 | v_65386;
assign v_65390 = v_65388 | v_65389;
assign v_65392 = v_65234 | v_65391;
assign v_65395 = v_65393 | v_65394;
assign v_65397 = v_65231 | v_65396;
assign v_65400 = v_65398 | v_65399;
assign v_65402 = v_65228 | v_65401;
assign v_65405 = v_65403 | v_65404;
assign v_65407 = v_65225 | v_65406;
assign v_65410 = v_65408 | v_65409;
assign v_65412 = v_65222 | v_65411;
assign v_65415 = v_65413 | v_65414;
assign v_65417 = v_65219 | v_65416;
assign v_65420 = v_65418 | v_65419;
assign v_65422 = v_65216 | v_65421;
assign v_65425 = v_65423 | v_65424;
assign v_65427 = v_65213 | v_65426;
assign v_65430 = v_65428 | v_65429;
assign v_65432 = v_65210 | v_65431;
assign v_65435 = v_65433 | v_65434;
assign v_65437 = v_65207 | v_65436;
assign v_65440 = v_65438 | v_65439;
assign v_65442 = v_65204 | v_65441;
assign v_65445 = v_65203 | v_65444;
assign v_65499 = v_65496 | v_65498;
assign v_65501 = v_65495 | v_65500;
assign v_65503 = v_65493 | v_65502;
assign v_65505 = v_65500 | v_65504;
assign v_65507 = v_65492 | v_65506;
assign v_65509 = v_65490 | v_65508;
assign v_65511 = v_65506 | v_65510;
assign v_65513 = v_65489 | v_65512;
assign v_65515 = v_65487 | v_65514;
assign v_65517 = v_65512 | v_65516;
assign v_65519 = v_65486 | v_65518;
assign v_65521 = v_65484 | v_65520;
assign v_65523 = v_65518 | v_65522;
assign v_65525 = v_65483 | v_65524;
assign v_65527 = v_65481 | v_65526;
assign v_65529 = v_65524 | v_65528;
assign v_65531 = v_65480 | v_65530;
assign v_65533 = v_65478 | v_65532;
assign v_65535 = v_65530 | v_65534;
assign v_65537 = v_65477 | v_65536;
assign v_65539 = v_65475 | v_65538;
assign v_65541 = v_65536 | v_65540;
assign v_65543 = v_65474 | v_65542;
assign v_65545 = v_65472 | v_65544;
assign v_65547 = v_65542 | v_65546;
assign v_65549 = v_65471 | v_65548;
assign v_65551 = v_65469 | v_65550;
assign v_65553 = v_65548 | v_65552;
assign v_65555 = v_65468 | v_65554;
assign v_65557 = v_65466 | v_65556;
assign v_65559 = v_65554 | v_65558;
assign v_65561 = v_65465 | v_65560;
assign v_65563 = v_65463 | v_65562;
assign v_65565 = v_65560 | v_65564;
assign v_65567 = v_65462 | v_65566;
assign v_65569 = v_65460 | v_65568;
assign v_65571 = v_65566 | v_65570;
assign v_65573 = v_65459 | v_65572;
assign v_65575 = v_65457 | v_65574;
assign v_65577 = v_65572 | v_65576;
assign v_65579 = v_65456 | v_65578;
assign v_65581 = v_65454 | v_65580;
assign v_65583 = v_65578 | v_65582;
assign v_65585 = v_65453 | v_65584;
assign v_65587 = v_65451 | v_65586;
assign v_65589 = v_65584 | v_65588;
assign v_65591 = v_65450 | v_65590;
assign v_65593 = v_65448 | v_65592;
assign v_65595 = v_65590 | v_65594;
assign v_65598 = ~v_65447 | v_65597;
assign v_65605 = v_65495 | v_65604;
assign v_65608 = v_65606 | v_65607;
assign v_65610 = v_65492 | v_65609;
assign v_65613 = v_65611 | v_65612;
assign v_65615 = v_65489 | v_65614;
assign v_65618 = v_65616 | v_65617;
assign v_65620 = v_65486 | v_65619;
assign v_65623 = v_65621 | v_65622;
assign v_65625 = v_65483 | v_65624;
assign v_65628 = v_65626 | v_65627;
assign v_65630 = v_65480 | v_65629;
assign v_65633 = v_65631 | v_65632;
assign v_65635 = v_65477 | v_65634;
assign v_65638 = v_65636 | v_65637;
assign v_65640 = v_65474 | v_65639;
assign v_65643 = v_65641 | v_65642;
assign v_65645 = v_65471 | v_65644;
assign v_65648 = v_65646 | v_65647;
assign v_65650 = v_65468 | v_65649;
assign v_65653 = v_65651 | v_65652;
assign v_65655 = v_65465 | v_65654;
assign v_65658 = v_65656 | v_65657;
assign v_65660 = v_65462 | v_65659;
assign v_65663 = v_65661 | v_65662;
assign v_65665 = v_65459 | v_65664;
assign v_65668 = v_65666 | v_65667;
assign v_65670 = v_65456 | v_65669;
assign v_65673 = v_65671 | v_65672;
assign v_65675 = v_65453 | v_65674;
assign v_65678 = v_65676 | v_65677;
assign v_65680 = v_65450 | v_65679;
assign v_65683 = v_65681 | v_65682;
assign v_65685 = v_65447 | v_65684;
assign v_65688 = v_65446 | v_65687;
assign v_65742 = v_65739 | v_65741;
assign v_65744 = v_65738 | v_65743;
assign v_65746 = v_65736 | v_65745;
assign v_65748 = v_65743 | v_65747;
assign v_65750 = v_65735 | v_65749;
assign v_65752 = v_65733 | v_65751;
assign v_65754 = v_65749 | v_65753;
assign v_65756 = v_65732 | v_65755;
assign v_65758 = v_65730 | v_65757;
assign v_65760 = v_65755 | v_65759;
assign v_65762 = v_65729 | v_65761;
assign v_65764 = v_65727 | v_65763;
assign v_65766 = v_65761 | v_65765;
assign v_65768 = v_65726 | v_65767;
assign v_65770 = v_65724 | v_65769;
assign v_65772 = v_65767 | v_65771;
assign v_65774 = v_65723 | v_65773;
assign v_65776 = v_65721 | v_65775;
assign v_65778 = v_65773 | v_65777;
assign v_65780 = v_65720 | v_65779;
assign v_65782 = v_65718 | v_65781;
assign v_65784 = v_65779 | v_65783;
assign v_65786 = v_65717 | v_65785;
assign v_65788 = v_65715 | v_65787;
assign v_65790 = v_65785 | v_65789;
assign v_65792 = v_65714 | v_65791;
assign v_65794 = v_65712 | v_65793;
assign v_65796 = v_65791 | v_65795;
assign v_65798 = v_65711 | v_65797;
assign v_65800 = v_65709 | v_65799;
assign v_65802 = v_65797 | v_65801;
assign v_65804 = v_65708 | v_65803;
assign v_65806 = v_65706 | v_65805;
assign v_65808 = v_65803 | v_65807;
assign v_65810 = v_65705 | v_65809;
assign v_65812 = v_65703 | v_65811;
assign v_65814 = v_65809 | v_65813;
assign v_65816 = v_65702 | v_65815;
assign v_65818 = v_65700 | v_65817;
assign v_65820 = v_65815 | v_65819;
assign v_65822 = v_65699 | v_65821;
assign v_65824 = v_65697 | v_65823;
assign v_65826 = v_65821 | v_65825;
assign v_65828 = v_65696 | v_65827;
assign v_65830 = v_65694 | v_65829;
assign v_65832 = v_65827 | v_65831;
assign v_65834 = v_65693 | v_65833;
assign v_65836 = v_65691 | v_65835;
assign v_65838 = v_65833 | v_65837;
assign v_65841 = ~v_65690 | v_65840;
assign v_65848 = v_65738 | v_65847;
assign v_65851 = v_65849 | v_65850;
assign v_65853 = v_65735 | v_65852;
assign v_65856 = v_65854 | v_65855;
assign v_65858 = v_65732 | v_65857;
assign v_65861 = v_65859 | v_65860;
assign v_65863 = v_65729 | v_65862;
assign v_65866 = v_65864 | v_65865;
assign v_65868 = v_65726 | v_65867;
assign v_65871 = v_65869 | v_65870;
assign v_65873 = v_65723 | v_65872;
assign v_65876 = v_65874 | v_65875;
assign v_65878 = v_65720 | v_65877;
assign v_65881 = v_65879 | v_65880;
assign v_65883 = v_65717 | v_65882;
assign v_65886 = v_65884 | v_65885;
assign v_65888 = v_65714 | v_65887;
assign v_65891 = v_65889 | v_65890;
assign v_65893 = v_65711 | v_65892;
assign v_65896 = v_65894 | v_65895;
assign v_65898 = v_65708 | v_65897;
assign v_65901 = v_65899 | v_65900;
assign v_65903 = v_65705 | v_65902;
assign v_65906 = v_65904 | v_65905;
assign v_65908 = v_65702 | v_65907;
assign v_65911 = v_65909 | v_65910;
assign v_65913 = v_65699 | v_65912;
assign v_65916 = v_65914 | v_65915;
assign v_65918 = v_65696 | v_65917;
assign v_65921 = v_65919 | v_65920;
assign v_65923 = v_65693 | v_65922;
assign v_65926 = v_65924 | v_65925;
assign v_65928 = v_65690 | v_65927;
assign v_65931 = v_65689 | v_65930;
assign v_65985 = v_65982 | v_65984;
assign v_65987 = v_65981 | v_65986;
assign v_65989 = v_65979 | v_65988;
assign v_65991 = v_65986 | v_65990;
assign v_65993 = v_65978 | v_65992;
assign v_65995 = v_65976 | v_65994;
assign v_65997 = v_65992 | v_65996;
assign v_65999 = v_65975 | v_65998;
assign v_66001 = v_65973 | v_66000;
assign v_66003 = v_65998 | v_66002;
assign v_66005 = v_65972 | v_66004;
assign v_66007 = v_65970 | v_66006;
assign v_66009 = v_66004 | v_66008;
assign v_66011 = v_65969 | v_66010;
assign v_66013 = v_65967 | v_66012;
assign v_66015 = v_66010 | v_66014;
assign v_66017 = v_65966 | v_66016;
assign v_66019 = v_65964 | v_66018;
assign v_66021 = v_66016 | v_66020;
assign v_66023 = v_65963 | v_66022;
assign v_66025 = v_65961 | v_66024;
assign v_66027 = v_66022 | v_66026;
assign v_66029 = v_65960 | v_66028;
assign v_66031 = v_65958 | v_66030;
assign v_66033 = v_66028 | v_66032;
assign v_66035 = v_65957 | v_66034;
assign v_66037 = v_65955 | v_66036;
assign v_66039 = v_66034 | v_66038;
assign v_66041 = v_65954 | v_66040;
assign v_66043 = v_65952 | v_66042;
assign v_66045 = v_66040 | v_66044;
assign v_66047 = v_65951 | v_66046;
assign v_66049 = v_65949 | v_66048;
assign v_66051 = v_66046 | v_66050;
assign v_66053 = v_65948 | v_66052;
assign v_66055 = v_65946 | v_66054;
assign v_66057 = v_66052 | v_66056;
assign v_66059 = v_65945 | v_66058;
assign v_66061 = v_65943 | v_66060;
assign v_66063 = v_66058 | v_66062;
assign v_66065 = v_65942 | v_66064;
assign v_66067 = v_65940 | v_66066;
assign v_66069 = v_66064 | v_66068;
assign v_66071 = v_65939 | v_66070;
assign v_66073 = v_65937 | v_66072;
assign v_66075 = v_66070 | v_66074;
assign v_66077 = v_65936 | v_66076;
assign v_66079 = v_65934 | v_66078;
assign v_66081 = v_66076 | v_66080;
assign v_66084 = ~v_65933 | v_66083;
assign v_66091 = v_65981 | v_66090;
assign v_66094 = v_66092 | v_66093;
assign v_66096 = v_65978 | v_66095;
assign v_66099 = v_66097 | v_66098;
assign v_66101 = v_65975 | v_66100;
assign v_66104 = v_66102 | v_66103;
assign v_66106 = v_65972 | v_66105;
assign v_66109 = v_66107 | v_66108;
assign v_66111 = v_65969 | v_66110;
assign v_66114 = v_66112 | v_66113;
assign v_66116 = v_65966 | v_66115;
assign v_66119 = v_66117 | v_66118;
assign v_66121 = v_65963 | v_66120;
assign v_66124 = v_66122 | v_66123;
assign v_66126 = v_65960 | v_66125;
assign v_66129 = v_66127 | v_66128;
assign v_66131 = v_65957 | v_66130;
assign v_66134 = v_66132 | v_66133;
assign v_66136 = v_65954 | v_66135;
assign v_66139 = v_66137 | v_66138;
assign v_66141 = v_65951 | v_66140;
assign v_66144 = v_66142 | v_66143;
assign v_66146 = v_65948 | v_66145;
assign v_66149 = v_66147 | v_66148;
assign v_66151 = v_65945 | v_66150;
assign v_66154 = v_66152 | v_66153;
assign v_66156 = v_65942 | v_66155;
assign v_66159 = v_66157 | v_66158;
assign v_66161 = v_65939 | v_66160;
assign v_66164 = v_66162 | v_66163;
assign v_66166 = v_65936 | v_66165;
assign v_66169 = v_66167 | v_66168;
assign v_66171 = v_65933 | v_66170;
assign v_66174 = v_65932 | v_66173;
assign v_66228 = v_66225 | v_66227;
assign v_66230 = v_66224 | v_66229;
assign v_66232 = v_66222 | v_66231;
assign v_66234 = v_66229 | v_66233;
assign v_66236 = v_66221 | v_66235;
assign v_66238 = v_66219 | v_66237;
assign v_66240 = v_66235 | v_66239;
assign v_66242 = v_66218 | v_66241;
assign v_66244 = v_66216 | v_66243;
assign v_66246 = v_66241 | v_66245;
assign v_66248 = v_66215 | v_66247;
assign v_66250 = v_66213 | v_66249;
assign v_66252 = v_66247 | v_66251;
assign v_66254 = v_66212 | v_66253;
assign v_66256 = v_66210 | v_66255;
assign v_66258 = v_66253 | v_66257;
assign v_66260 = v_66209 | v_66259;
assign v_66262 = v_66207 | v_66261;
assign v_66264 = v_66259 | v_66263;
assign v_66266 = v_66206 | v_66265;
assign v_66268 = v_66204 | v_66267;
assign v_66270 = v_66265 | v_66269;
assign v_66272 = v_66203 | v_66271;
assign v_66274 = v_66201 | v_66273;
assign v_66276 = v_66271 | v_66275;
assign v_66278 = v_66200 | v_66277;
assign v_66280 = v_66198 | v_66279;
assign v_66282 = v_66277 | v_66281;
assign v_66284 = v_66197 | v_66283;
assign v_66286 = v_66195 | v_66285;
assign v_66288 = v_66283 | v_66287;
assign v_66290 = v_66194 | v_66289;
assign v_66292 = v_66192 | v_66291;
assign v_66294 = v_66289 | v_66293;
assign v_66296 = v_66191 | v_66295;
assign v_66298 = v_66189 | v_66297;
assign v_66300 = v_66295 | v_66299;
assign v_66302 = v_66188 | v_66301;
assign v_66304 = v_66186 | v_66303;
assign v_66306 = v_66301 | v_66305;
assign v_66308 = v_66185 | v_66307;
assign v_66310 = v_66183 | v_66309;
assign v_66312 = v_66307 | v_66311;
assign v_66314 = v_66182 | v_66313;
assign v_66316 = v_66180 | v_66315;
assign v_66318 = v_66313 | v_66317;
assign v_66320 = v_66179 | v_66319;
assign v_66322 = v_66177 | v_66321;
assign v_66324 = v_66319 | v_66323;
assign v_66327 = ~v_66176 | v_66326;
assign v_66334 = v_66224 | v_66333;
assign v_66337 = v_66335 | v_66336;
assign v_66339 = v_66221 | v_66338;
assign v_66342 = v_66340 | v_66341;
assign v_66344 = v_66218 | v_66343;
assign v_66347 = v_66345 | v_66346;
assign v_66349 = v_66215 | v_66348;
assign v_66352 = v_66350 | v_66351;
assign v_66354 = v_66212 | v_66353;
assign v_66357 = v_66355 | v_66356;
assign v_66359 = v_66209 | v_66358;
assign v_66362 = v_66360 | v_66361;
assign v_66364 = v_66206 | v_66363;
assign v_66367 = v_66365 | v_66366;
assign v_66369 = v_66203 | v_66368;
assign v_66372 = v_66370 | v_66371;
assign v_66374 = v_66200 | v_66373;
assign v_66377 = v_66375 | v_66376;
assign v_66379 = v_66197 | v_66378;
assign v_66382 = v_66380 | v_66381;
assign v_66384 = v_66194 | v_66383;
assign v_66387 = v_66385 | v_66386;
assign v_66389 = v_66191 | v_66388;
assign v_66392 = v_66390 | v_66391;
assign v_66394 = v_66188 | v_66393;
assign v_66397 = v_66395 | v_66396;
assign v_66399 = v_66185 | v_66398;
assign v_66402 = v_66400 | v_66401;
assign v_66404 = v_66182 | v_66403;
assign v_66407 = v_66405 | v_66406;
assign v_66409 = v_66179 | v_66408;
assign v_66412 = v_66410 | v_66411;
assign v_66414 = v_66176 | v_66413;
assign v_66417 = v_66175 | v_66416;
assign v_66470 = v_66467 | v_66469;
assign v_66472 = v_66466 | v_66471;
assign v_66474 = v_66464 | v_66473;
assign v_66476 = v_66471 | v_66475;
assign v_66478 = v_66463 | v_66477;
assign v_66480 = v_66461 | v_66479;
assign v_66482 = v_66477 | v_66481;
assign v_66484 = v_66460 | v_66483;
assign v_66486 = v_66458 | v_66485;
assign v_66488 = v_66483 | v_66487;
assign v_66490 = v_66457 | v_66489;
assign v_66492 = v_66455 | v_66491;
assign v_66494 = v_66489 | v_66493;
assign v_66496 = v_66454 | v_66495;
assign v_66498 = v_66452 | v_66497;
assign v_66500 = v_66495 | v_66499;
assign v_66502 = v_66451 | v_66501;
assign v_66504 = v_66449 | v_66503;
assign v_66506 = v_66501 | v_66505;
assign v_66508 = v_66448 | v_66507;
assign v_66510 = v_66446 | v_66509;
assign v_66512 = v_66507 | v_66511;
assign v_66514 = v_66445 | v_66513;
assign v_66516 = v_66443 | v_66515;
assign v_66518 = v_66513 | v_66517;
assign v_66520 = v_66442 | v_66519;
assign v_66522 = v_66440 | v_66521;
assign v_66524 = v_66519 | v_66523;
assign v_66526 = v_66439 | v_66525;
assign v_66528 = v_66437 | v_66527;
assign v_66530 = v_66525 | v_66529;
assign v_66532 = v_66436 | v_66531;
assign v_66534 = v_66434 | v_66533;
assign v_66536 = v_66531 | v_66535;
assign v_66538 = v_66433 | v_66537;
assign v_66540 = v_66431 | v_66539;
assign v_66542 = v_66537 | v_66541;
assign v_66544 = v_66430 | v_66543;
assign v_66546 = v_66428 | v_66545;
assign v_66548 = v_66543 | v_66547;
assign v_66550 = v_66427 | v_66549;
assign v_66552 = v_66425 | v_66551;
assign v_66554 = v_66549 | v_66553;
assign v_66556 = v_66424 | v_66555;
assign v_66558 = v_66422 | v_66557;
assign v_66560 = v_66555 | v_66559;
assign v_66562 = v_66421 | v_66561;
assign v_66564 = v_66419 | v_66563;
assign v_66566 = v_66561 | v_66565;
assign v_66570 = v_66567 | v_66569;
assign v_66577 = v_66466 | v_66576;
assign v_66580 = v_66578 | v_66579;
assign v_66582 = v_66463 | v_66581;
assign v_66585 = v_66583 | v_66584;
assign v_66587 = v_66460 | v_66586;
assign v_66590 = v_66588 | v_66589;
assign v_66592 = v_66457 | v_66591;
assign v_66595 = v_66593 | v_66594;
assign v_66597 = v_66454 | v_66596;
assign v_66600 = v_66598 | v_66599;
assign v_66602 = v_66451 | v_66601;
assign v_66605 = v_66603 | v_66604;
assign v_66607 = v_66448 | v_66606;
assign v_66610 = v_66608 | v_66609;
assign v_66612 = v_66445 | v_66611;
assign v_66615 = v_66613 | v_66614;
assign v_66617 = v_66442 | v_66616;
assign v_66620 = v_66618 | v_66619;
assign v_66622 = v_66439 | v_66621;
assign v_66625 = v_66623 | v_66624;
assign v_66627 = v_66436 | v_66626;
assign v_66630 = v_66628 | v_66629;
assign v_66632 = v_66433 | v_66631;
assign v_66635 = v_66633 | v_66634;
assign v_66637 = v_66430 | v_66636;
assign v_66640 = v_66638 | v_66639;
assign v_66642 = v_66427 | v_66641;
assign v_66645 = v_66643 | v_66644;
assign v_66647 = v_66424 | v_66646;
assign v_66650 = v_66648 | v_66649;
assign v_66652 = v_66421 | v_66651;
assign v_66655 = v_66653 | v_66654;
assign v_66657 = v_66655 | v_66656;
assign v_66660 = v_66418 | v_66659;
assign v_66730 = v_66727 | v_66729;
assign v_66732 = v_66725 | v_66731;
assign v_66734 = v_66723 | v_66733;
assign v_66736 = v_66731 | v_66735;
assign v_66738 = v_66721 | v_66737;
assign v_66740 = v_66719 | v_66739;
assign v_66742 = v_66737 | v_66741;
assign v_66744 = v_66717 | v_66743;
assign v_66746 = v_66715 | v_66745;
assign v_66748 = v_66743 | v_66747;
assign v_66750 = v_66713 | v_66749;
assign v_66752 = v_66711 | v_66751;
assign v_66754 = v_66749 | v_66753;
assign v_66756 = v_66709 | v_66755;
assign v_66758 = v_66707 | v_66757;
assign v_66760 = v_66755 | v_66759;
assign v_66762 = v_66705 | v_66761;
assign v_66764 = v_66703 | v_66763;
assign v_66766 = v_66761 | v_66765;
assign v_66768 = v_66701 | v_66767;
assign v_66770 = v_66699 | v_66769;
assign v_66772 = v_66767 | v_66771;
assign v_66774 = v_66697 | v_66773;
assign v_66776 = v_66695 | v_66775;
assign v_66778 = v_66773 | v_66777;
assign v_66780 = v_66693 | v_66779;
assign v_66782 = v_66691 | v_66781;
assign v_66784 = v_66779 | v_66783;
assign v_66786 = v_66689 | v_66785;
assign v_66788 = v_66687 | v_66787;
assign v_66790 = v_66785 | v_66789;
assign v_66792 = v_66685 | v_66791;
assign v_66794 = v_66683 | v_66793;
assign v_66796 = v_66791 | v_66795;
assign v_66798 = v_66681 | v_66797;
assign v_66800 = v_66679 | v_66799;
assign v_66802 = v_66797 | v_66801;
assign v_66804 = v_66677 | v_66803;
assign v_66806 = v_66674 | v_66805;
assign v_66808 = v_66803 | v_66807;
assign v_66810 = v_66673 | v_66809;
assign v_66812 = v_66670 | v_66811;
assign v_66814 = v_66809 | v_66813;
assign v_66816 = v_66669 | v_66815;
assign v_66818 = v_66666 | v_66817;
assign v_66820 = v_66815 | v_66819;
assign v_66822 = v_66665 | v_66821;
assign v_66824 = v_66662 | v_66823;
assign v_66826 = v_66821 | v_66825;
assign v_66830 = v_66827 | v_66829;
assign v_66837 = v_66725 | v_66836;
assign v_66840 = v_66838 | v_66839;
assign v_66842 = v_66721 | v_66841;
assign v_66845 = v_66843 | v_66844;
assign v_66847 = v_66717 | v_66846;
assign v_66850 = v_66848 | v_66849;
assign v_66852 = v_66713 | v_66851;
assign v_66855 = v_66853 | v_66854;
assign v_66857 = v_66709 | v_66856;
assign v_66860 = v_66858 | v_66859;
assign v_66862 = v_66705 | v_66861;
assign v_66865 = v_66863 | v_66864;
assign v_66867 = v_66701 | v_66866;
assign v_66870 = v_66868 | v_66869;
assign v_66872 = v_66697 | v_66871;
assign v_66875 = v_66873 | v_66874;
assign v_66877 = v_66693 | v_66876;
assign v_66880 = v_66878 | v_66879;
assign v_66882 = v_66689 | v_66881;
assign v_66885 = v_66883 | v_66884;
assign v_66887 = v_66685 | v_66886;
assign v_66890 = v_66888 | v_66889;
assign v_66892 = v_66681 | v_66891;
assign v_66895 = v_66893 | v_66894;
assign v_66897 = v_66677 | v_66896;
assign v_66900 = v_66898 | v_66899;
assign v_66902 = v_66673 | v_66901;
assign v_66905 = v_66903 | v_66904;
assign v_66907 = v_66669 | v_66906;
assign v_66910 = v_66908 | v_66909;
assign v_66912 = v_66665 | v_66911;
assign v_66915 = v_66913 | v_66914;
assign v_66917 = v_66915 | v_66916;
assign v_66920 = v_66661 | v_66919;
assign v_66973 = v_66970 | v_66972;
assign v_66975 = v_66969 | v_66974;
assign v_66977 = v_66967 | v_66976;
assign v_66979 = v_66974 | v_66978;
assign v_66981 = v_66966 | v_66980;
assign v_66983 = v_66964 | v_66982;
assign v_66985 = v_66980 | v_66984;
assign v_66987 = v_66963 | v_66986;
assign v_66989 = v_66961 | v_66988;
assign v_66991 = v_66986 | v_66990;
assign v_66993 = v_66960 | v_66992;
assign v_66995 = v_66958 | v_66994;
assign v_66997 = v_66992 | v_66996;
assign v_66999 = v_66957 | v_66998;
assign v_67001 = v_66955 | v_67000;
assign v_67003 = v_66998 | v_67002;
assign v_67005 = v_66954 | v_67004;
assign v_67007 = v_66952 | v_67006;
assign v_67009 = v_67004 | v_67008;
assign v_67011 = v_66951 | v_67010;
assign v_67013 = v_66949 | v_67012;
assign v_67015 = v_67010 | v_67014;
assign v_67017 = v_66948 | v_67016;
assign v_67019 = v_66946 | v_67018;
assign v_67021 = v_67016 | v_67020;
assign v_67023 = v_66945 | v_67022;
assign v_67025 = v_66943 | v_67024;
assign v_67027 = v_67022 | v_67026;
assign v_67029 = v_66942 | v_67028;
assign v_67031 = v_66940 | v_67030;
assign v_67033 = v_67028 | v_67032;
assign v_67035 = v_66939 | v_67034;
assign v_67037 = v_66937 | v_67036;
assign v_67039 = v_67034 | v_67038;
assign v_67041 = v_66936 | v_67040;
assign v_67043 = v_66934 | v_67042;
assign v_67045 = v_67040 | v_67044;
assign v_67047 = v_66933 | v_67046;
assign v_67049 = v_66931 | v_67048;
assign v_67051 = v_67046 | v_67050;
assign v_67053 = v_66930 | v_67052;
assign v_67055 = v_66928 | v_67054;
assign v_67057 = v_67052 | v_67056;
assign v_67059 = v_66927 | v_67058;
assign v_67061 = v_66925 | v_67060;
assign v_67063 = v_67058 | v_67062;
assign v_67065 = v_66924 | v_67064;
assign v_67067 = v_66922 | v_67066;
assign v_67069 = v_67064 | v_67068;
assign v_67073 = v_67070 | v_67072;
assign v_67080 = v_66969 | v_67079;
assign v_67083 = v_67081 | v_67082;
assign v_67085 = v_66966 | v_67084;
assign v_67088 = v_67086 | v_67087;
assign v_67090 = v_66963 | v_67089;
assign v_67093 = v_67091 | v_67092;
assign v_67095 = v_66960 | v_67094;
assign v_67098 = v_67096 | v_67097;
assign v_67100 = v_66957 | v_67099;
assign v_67103 = v_67101 | v_67102;
assign v_67105 = v_66954 | v_67104;
assign v_67108 = v_67106 | v_67107;
assign v_67110 = v_66951 | v_67109;
assign v_67113 = v_67111 | v_67112;
assign v_67115 = v_66948 | v_67114;
assign v_67118 = v_67116 | v_67117;
assign v_67120 = v_66945 | v_67119;
assign v_67123 = v_67121 | v_67122;
assign v_67125 = v_66942 | v_67124;
assign v_67128 = v_67126 | v_67127;
assign v_67130 = v_66939 | v_67129;
assign v_67133 = v_67131 | v_67132;
assign v_67135 = v_66936 | v_67134;
assign v_67138 = v_67136 | v_67137;
assign v_67140 = v_66933 | v_67139;
assign v_67143 = v_67141 | v_67142;
assign v_67145 = v_66930 | v_67144;
assign v_67148 = v_67146 | v_67147;
assign v_67150 = v_66927 | v_67149;
assign v_67153 = v_67151 | v_67152;
assign v_67155 = v_66924 | v_67154;
assign v_67158 = v_67156 | v_67157;
assign v_67160 = v_67158 | v_67159;
assign v_67163 = v_66921 | v_67162;
assign v_67216 = v_67213 | v_67215;
assign v_67218 = v_67212 | v_67217;
assign v_67220 = v_67210 | v_67219;
assign v_67222 = v_67217 | v_67221;
assign v_67224 = v_67209 | v_67223;
assign v_67226 = v_67207 | v_67225;
assign v_67228 = v_67223 | v_67227;
assign v_67230 = v_67206 | v_67229;
assign v_67232 = v_67204 | v_67231;
assign v_67234 = v_67229 | v_67233;
assign v_67236 = v_67203 | v_67235;
assign v_67238 = v_67201 | v_67237;
assign v_67240 = v_67235 | v_67239;
assign v_67242 = v_67200 | v_67241;
assign v_67244 = v_67198 | v_67243;
assign v_67246 = v_67241 | v_67245;
assign v_67248 = v_67197 | v_67247;
assign v_67250 = v_67195 | v_67249;
assign v_67252 = v_67247 | v_67251;
assign v_67254 = v_67194 | v_67253;
assign v_67256 = v_67192 | v_67255;
assign v_67258 = v_67253 | v_67257;
assign v_67260 = v_67191 | v_67259;
assign v_67262 = v_67189 | v_67261;
assign v_67264 = v_67259 | v_67263;
assign v_67266 = v_67188 | v_67265;
assign v_67268 = v_67186 | v_67267;
assign v_67270 = v_67265 | v_67269;
assign v_67272 = v_67185 | v_67271;
assign v_67274 = v_67183 | v_67273;
assign v_67276 = v_67271 | v_67275;
assign v_67278 = v_67182 | v_67277;
assign v_67280 = v_67180 | v_67279;
assign v_67282 = v_67277 | v_67281;
assign v_67284 = v_67179 | v_67283;
assign v_67286 = v_67177 | v_67285;
assign v_67288 = v_67283 | v_67287;
assign v_67290 = v_67176 | v_67289;
assign v_67292 = v_67174 | v_67291;
assign v_67294 = v_67289 | v_67293;
assign v_67296 = v_67173 | v_67295;
assign v_67298 = v_67171 | v_67297;
assign v_67300 = v_67295 | v_67299;
assign v_67302 = v_67170 | v_67301;
assign v_67304 = v_67168 | v_67303;
assign v_67306 = v_67301 | v_67305;
assign v_67308 = v_67167 | v_67307;
assign v_67310 = v_67165 | v_67309;
assign v_67312 = v_67307 | v_67311;
assign v_67316 = v_67313 | v_67315;
assign v_67323 = v_67212 | v_67322;
assign v_67326 = v_67324 | v_67325;
assign v_67328 = v_67209 | v_67327;
assign v_67331 = v_67329 | v_67330;
assign v_67333 = v_67206 | v_67332;
assign v_67336 = v_67334 | v_67335;
assign v_67338 = v_67203 | v_67337;
assign v_67341 = v_67339 | v_67340;
assign v_67343 = v_67200 | v_67342;
assign v_67346 = v_67344 | v_67345;
assign v_67348 = v_67197 | v_67347;
assign v_67351 = v_67349 | v_67350;
assign v_67353 = v_67194 | v_67352;
assign v_67356 = v_67354 | v_67355;
assign v_67358 = v_67191 | v_67357;
assign v_67361 = v_67359 | v_67360;
assign v_67363 = v_67188 | v_67362;
assign v_67366 = v_67364 | v_67365;
assign v_67368 = v_67185 | v_67367;
assign v_67371 = v_67369 | v_67370;
assign v_67373 = v_67182 | v_67372;
assign v_67376 = v_67374 | v_67375;
assign v_67378 = v_67179 | v_67377;
assign v_67381 = v_67379 | v_67380;
assign v_67383 = v_67176 | v_67382;
assign v_67386 = v_67384 | v_67385;
assign v_67388 = v_67173 | v_67387;
assign v_67391 = v_67389 | v_67390;
assign v_67393 = v_67170 | v_67392;
assign v_67396 = v_67394 | v_67395;
assign v_67398 = v_67167 | v_67397;
assign v_67401 = v_67399 | v_67400;
assign v_67403 = v_67401 | v_67402;
assign v_67406 = v_67164 | v_67405;
assign v_67459 = v_67456 | v_67458;
assign v_67461 = v_67455 | v_67460;
assign v_67463 = v_67453 | v_67462;
assign v_67465 = v_67460 | v_67464;
assign v_67467 = v_67452 | v_67466;
assign v_67469 = v_67450 | v_67468;
assign v_67471 = v_67466 | v_67470;
assign v_67473 = v_67449 | v_67472;
assign v_67475 = v_67447 | v_67474;
assign v_67477 = v_67472 | v_67476;
assign v_67479 = v_67446 | v_67478;
assign v_67481 = v_67444 | v_67480;
assign v_67483 = v_67478 | v_67482;
assign v_67485 = v_67443 | v_67484;
assign v_67487 = v_67441 | v_67486;
assign v_67489 = v_67484 | v_67488;
assign v_67491 = v_67440 | v_67490;
assign v_67493 = v_67438 | v_67492;
assign v_67495 = v_67490 | v_67494;
assign v_67497 = v_67437 | v_67496;
assign v_67499 = v_67435 | v_67498;
assign v_67501 = v_67496 | v_67500;
assign v_67503 = v_67434 | v_67502;
assign v_67505 = v_67432 | v_67504;
assign v_67507 = v_67502 | v_67506;
assign v_67509 = v_67431 | v_67508;
assign v_67511 = v_67429 | v_67510;
assign v_67513 = v_67508 | v_67512;
assign v_67515 = v_67428 | v_67514;
assign v_67517 = v_67426 | v_67516;
assign v_67519 = v_67514 | v_67518;
assign v_67521 = v_67425 | v_67520;
assign v_67523 = v_67423 | v_67522;
assign v_67525 = v_67520 | v_67524;
assign v_67527 = v_67422 | v_67526;
assign v_67529 = v_67420 | v_67528;
assign v_67531 = v_67526 | v_67530;
assign v_67533 = v_67419 | v_67532;
assign v_67535 = v_67417 | v_67534;
assign v_67537 = v_67532 | v_67536;
assign v_67539 = v_67416 | v_67538;
assign v_67541 = v_67414 | v_67540;
assign v_67543 = v_67538 | v_67542;
assign v_67545 = v_67413 | v_67544;
assign v_67547 = v_67411 | v_67546;
assign v_67549 = v_67544 | v_67548;
assign v_67551 = v_67410 | v_67550;
assign v_67553 = v_67408 | v_67552;
assign v_67555 = v_67550 | v_67554;
assign v_67559 = v_67556 | v_67558;
assign v_67566 = v_67455 | v_67565;
assign v_67569 = v_67567 | v_67568;
assign v_67571 = v_67452 | v_67570;
assign v_67574 = v_67572 | v_67573;
assign v_67576 = v_67449 | v_67575;
assign v_67579 = v_67577 | v_67578;
assign v_67581 = v_67446 | v_67580;
assign v_67584 = v_67582 | v_67583;
assign v_67586 = v_67443 | v_67585;
assign v_67589 = v_67587 | v_67588;
assign v_67591 = v_67440 | v_67590;
assign v_67594 = v_67592 | v_67593;
assign v_67596 = v_67437 | v_67595;
assign v_67599 = v_67597 | v_67598;
assign v_67601 = v_67434 | v_67600;
assign v_67604 = v_67602 | v_67603;
assign v_67606 = v_67431 | v_67605;
assign v_67609 = v_67607 | v_67608;
assign v_67611 = v_67428 | v_67610;
assign v_67614 = v_67612 | v_67613;
assign v_67616 = v_67425 | v_67615;
assign v_67619 = v_67617 | v_67618;
assign v_67621 = v_67422 | v_67620;
assign v_67624 = v_67622 | v_67623;
assign v_67626 = v_67419 | v_67625;
assign v_67629 = v_67627 | v_67628;
assign v_67631 = v_67416 | v_67630;
assign v_67634 = v_67632 | v_67633;
assign v_67636 = v_67413 | v_67635;
assign v_67639 = v_67637 | v_67638;
assign v_67641 = v_67410 | v_67640;
assign v_67644 = v_67642 | v_67643;
assign v_67646 = v_67644 | v_67645;
assign v_67649 = v_67407 | v_67648;
assign v_67702 = v_67699 | v_67701;
assign v_67704 = v_67698 | v_67703;
assign v_67706 = v_67696 | v_67705;
assign v_67708 = v_67703 | v_67707;
assign v_67710 = v_67695 | v_67709;
assign v_67712 = v_67693 | v_67711;
assign v_67714 = v_67709 | v_67713;
assign v_67716 = v_67692 | v_67715;
assign v_67718 = v_67690 | v_67717;
assign v_67720 = v_67715 | v_67719;
assign v_67722 = v_67689 | v_67721;
assign v_67724 = v_67687 | v_67723;
assign v_67726 = v_67721 | v_67725;
assign v_67728 = v_67686 | v_67727;
assign v_67730 = v_67684 | v_67729;
assign v_67732 = v_67727 | v_67731;
assign v_67734 = v_67683 | v_67733;
assign v_67736 = v_67681 | v_67735;
assign v_67738 = v_67733 | v_67737;
assign v_67740 = v_67680 | v_67739;
assign v_67742 = v_67678 | v_67741;
assign v_67744 = v_67739 | v_67743;
assign v_67746 = v_67677 | v_67745;
assign v_67748 = v_67675 | v_67747;
assign v_67750 = v_67745 | v_67749;
assign v_67752 = v_67674 | v_67751;
assign v_67754 = v_67672 | v_67753;
assign v_67756 = v_67751 | v_67755;
assign v_67758 = v_67671 | v_67757;
assign v_67760 = v_67669 | v_67759;
assign v_67762 = v_67757 | v_67761;
assign v_67764 = v_67668 | v_67763;
assign v_67766 = v_67666 | v_67765;
assign v_67768 = v_67763 | v_67767;
assign v_67770 = v_67665 | v_67769;
assign v_67772 = v_67663 | v_67771;
assign v_67774 = v_67769 | v_67773;
assign v_67776 = v_67662 | v_67775;
assign v_67778 = v_67660 | v_67777;
assign v_67780 = v_67775 | v_67779;
assign v_67782 = v_67659 | v_67781;
assign v_67784 = v_67657 | v_67783;
assign v_67786 = v_67781 | v_67785;
assign v_67788 = v_67656 | v_67787;
assign v_67790 = v_67654 | v_67789;
assign v_67792 = v_67787 | v_67791;
assign v_67794 = v_67653 | v_67793;
assign v_67796 = v_67651 | v_67795;
assign v_67798 = v_67793 | v_67797;
assign v_67802 = v_67799 | v_67801;
assign v_67809 = v_67698 | v_67808;
assign v_67812 = v_67810 | v_67811;
assign v_67814 = v_67695 | v_67813;
assign v_67817 = v_67815 | v_67816;
assign v_67819 = v_67692 | v_67818;
assign v_67822 = v_67820 | v_67821;
assign v_67824 = v_67689 | v_67823;
assign v_67827 = v_67825 | v_67826;
assign v_67829 = v_67686 | v_67828;
assign v_67832 = v_67830 | v_67831;
assign v_67834 = v_67683 | v_67833;
assign v_67837 = v_67835 | v_67836;
assign v_67839 = v_67680 | v_67838;
assign v_67842 = v_67840 | v_67841;
assign v_67844 = v_67677 | v_67843;
assign v_67847 = v_67845 | v_67846;
assign v_67849 = v_67674 | v_67848;
assign v_67852 = v_67850 | v_67851;
assign v_67854 = v_67671 | v_67853;
assign v_67857 = v_67855 | v_67856;
assign v_67859 = v_67668 | v_67858;
assign v_67862 = v_67860 | v_67861;
assign v_67864 = v_67665 | v_67863;
assign v_67867 = v_67865 | v_67866;
assign v_67869 = v_67662 | v_67868;
assign v_67872 = v_67870 | v_67871;
assign v_67874 = v_67659 | v_67873;
assign v_67877 = v_67875 | v_67876;
assign v_67879 = v_67656 | v_67878;
assign v_67882 = v_67880 | v_67881;
assign v_67884 = v_67653 | v_67883;
assign v_67887 = v_67885 | v_67886;
assign v_67889 = v_67887 | v_67888;
assign v_67892 = v_67650 | v_67891;
assign v_67945 = v_67942 | v_67944;
assign v_67947 = v_67941 | v_67946;
assign v_67949 = v_67939 | v_67948;
assign v_67951 = v_67946 | v_67950;
assign v_67953 = v_67938 | v_67952;
assign v_67955 = v_67936 | v_67954;
assign v_67957 = v_67952 | v_67956;
assign v_67959 = v_67935 | v_67958;
assign v_67961 = v_67933 | v_67960;
assign v_67963 = v_67958 | v_67962;
assign v_67965 = v_67932 | v_67964;
assign v_67967 = v_67930 | v_67966;
assign v_67969 = v_67964 | v_67968;
assign v_67971 = v_67929 | v_67970;
assign v_67973 = v_67927 | v_67972;
assign v_67975 = v_67970 | v_67974;
assign v_67977 = v_67926 | v_67976;
assign v_67979 = v_67924 | v_67978;
assign v_67981 = v_67976 | v_67980;
assign v_67983 = v_67923 | v_67982;
assign v_67985 = v_67921 | v_67984;
assign v_67987 = v_67982 | v_67986;
assign v_67989 = v_67920 | v_67988;
assign v_67991 = v_67918 | v_67990;
assign v_67993 = v_67988 | v_67992;
assign v_67995 = v_67917 | v_67994;
assign v_67997 = v_67915 | v_67996;
assign v_67999 = v_67994 | v_67998;
assign v_68001 = v_67914 | v_68000;
assign v_68003 = v_67912 | v_68002;
assign v_68005 = v_68000 | v_68004;
assign v_68007 = v_67911 | v_68006;
assign v_68009 = v_67909 | v_68008;
assign v_68011 = v_68006 | v_68010;
assign v_68013 = v_67908 | v_68012;
assign v_68015 = v_67906 | v_68014;
assign v_68017 = v_68012 | v_68016;
assign v_68019 = v_67905 | v_68018;
assign v_68021 = v_67903 | v_68020;
assign v_68023 = v_68018 | v_68022;
assign v_68025 = v_67902 | v_68024;
assign v_68027 = v_67900 | v_68026;
assign v_68029 = v_68024 | v_68028;
assign v_68031 = v_67899 | v_68030;
assign v_68033 = v_67897 | v_68032;
assign v_68035 = v_68030 | v_68034;
assign v_68037 = v_67896 | v_68036;
assign v_68039 = v_67894 | v_68038;
assign v_68041 = v_68036 | v_68040;
assign v_68045 = v_68042 | v_68044;
assign v_68052 = v_67941 | v_68051;
assign v_68055 = v_68053 | v_68054;
assign v_68057 = v_67938 | v_68056;
assign v_68060 = v_68058 | v_68059;
assign v_68062 = v_67935 | v_68061;
assign v_68065 = v_68063 | v_68064;
assign v_68067 = v_67932 | v_68066;
assign v_68070 = v_68068 | v_68069;
assign v_68072 = v_67929 | v_68071;
assign v_68075 = v_68073 | v_68074;
assign v_68077 = v_67926 | v_68076;
assign v_68080 = v_68078 | v_68079;
assign v_68082 = v_67923 | v_68081;
assign v_68085 = v_68083 | v_68084;
assign v_68087 = v_67920 | v_68086;
assign v_68090 = v_68088 | v_68089;
assign v_68092 = v_67917 | v_68091;
assign v_68095 = v_68093 | v_68094;
assign v_68097 = v_67914 | v_68096;
assign v_68100 = v_68098 | v_68099;
assign v_68102 = v_67911 | v_68101;
assign v_68105 = v_68103 | v_68104;
assign v_68107 = v_67908 | v_68106;
assign v_68110 = v_68108 | v_68109;
assign v_68112 = v_67905 | v_68111;
assign v_68115 = v_68113 | v_68114;
assign v_68117 = v_67902 | v_68116;
assign v_68120 = v_68118 | v_68119;
assign v_68122 = v_67899 | v_68121;
assign v_68125 = v_68123 | v_68124;
assign v_68127 = v_67896 | v_68126;
assign v_68130 = v_68128 | v_68129;
assign v_68132 = v_68130 | v_68131;
assign v_68135 = v_67893 | v_68134;
assign v_68188 = v_68185 | v_68187;
assign v_68190 = v_68184 | v_68189;
assign v_68192 = v_68182 | v_68191;
assign v_68194 = v_68189 | v_68193;
assign v_68196 = v_68181 | v_68195;
assign v_68198 = v_68179 | v_68197;
assign v_68200 = v_68195 | v_68199;
assign v_68202 = v_68178 | v_68201;
assign v_68204 = v_68176 | v_68203;
assign v_68206 = v_68201 | v_68205;
assign v_68208 = v_68175 | v_68207;
assign v_68210 = v_68173 | v_68209;
assign v_68212 = v_68207 | v_68211;
assign v_68214 = v_68172 | v_68213;
assign v_68216 = v_68170 | v_68215;
assign v_68218 = v_68213 | v_68217;
assign v_68220 = v_68169 | v_68219;
assign v_68222 = v_68167 | v_68221;
assign v_68224 = v_68219 | v_68223;
assign v_68226 = v_68166 | v_68225;
assign v_68228 = v_68164 | v_68227;
assign v_68230 = v_68225 | v_68229;
assign v_68232 = v_68163 | v_68231;
assign v_68234 = v_68161 | v_68233;
assign v_68236 = v_68231 | v_68235;
assign v_68238 = v_68160 | v_68237;
assign v_68240 = v_68158 | v_68239;
assign v_68242 = v_68237 | v_68241;
assign v_68244 = v_68157 | v_68243;
assign v_68246 = v_68155 | v_68245;
assign v_68248 = v_68243 | v_68247;
assign v_68250 = v_68154 | v_68249;
assign v_68252 = v_68152 | v_68251;
assign v_68254 = v_68249 | v_68253;
assign v_68256 = v_68151 | v_68255;
assign v_68258 = v_68149 | v_68257;
assign v_68260 = v_68255 | v_68259;
assign v_68262 = v_68148 | v_68261;
assign v_68264 = v_68146 | v_68263;
assign v_68266 = v_68261 | v_68265;
assign v_68268 = v_68145 | v_68267;
assign v_68270 = v_68143 | v_68269;
assign v_68272 = v_68267 | v_68271;
assign v_68274 = v_68142 | v_68273;
assign v_68276 = v_68140 | v_68275;
assign v_68278 = v_68273 | v_68277;
assign v_68280 = v_68139 | v_68279;
assign v_68282 = v_68137 | v_68281;
assign v_68284 = v_68279 | v_68283;
assign v_68288 = v_68285 | v_68287;
assign v_68295 = v_68184 | v_68294;
assign v_68298 = v_68296 | v_68297;
assign v_68300 = v_68181 | v_68299;
assign v_68303 = v_68301 | v_68302;
assign v_68305 = v_68178 | v_68304;
assign v_68308 = v_68306 | v_68307;
assign v_68310 = v_68175 | v_68309;
assign v_68313 = v_68311 | v_68312;
assign v_68315 = v_68172 | v_68314;
assign v_68318 = v_68316 | v_68317;
assign v_68320 = v_68169 | v_68319;
assign v_68323 = v_68321 | v_68322;
assign v_68325 = v_68166 | v_68324;
assign v_68328 = v_68326 | v_68327;
assign v_68330 = v_68163 | v_68329;
assign v_68333 = v_68331 | v_68332;
assign v_68335 = v_68160 | v_68334;
assign v_68338 = v_68336 | v_68337;
assign v_68340 = v_68157 | v_68339;
assign v_68343 = v_68341 | v_68342;
assign v_68345 = v_68154 | v_68344;
assign v_68348 = v_68346 | v_68347;
assign v_68350 = v_68151 | v_68349;
assign v_68353 = v_68351 | v_68352;
assign v_68355 = v_68148 | v_68354;
assign v_68358 = v_68356 | v_68357;
assign v_68360 = v_68145 | v_68359;
assign v_68363 = v_68361 | v_68362;
assign v_68365 = v_68142 | v_68364;
assign v_68368 = v_68366 | v_68367;
assign v_68370 = v_68139 | v_68369;
assign v_68373 = v_68371 | v_68372;
assign v_68375 = v_68373 | v_68374;
assign v_68378 = v_68136 | v_68377;
assign v_68431 = v_68428 | v_68430;
assign v_68433 = v_68427 | v_68432;
assign v_68435 = v_68425 | v_68434;
assign v_68437 = v_68432 | v_68436;
assign v_68439 = v_68424 | v_68438;
assign v_68441 = v_68422 | v_68440;
assign v_68443 = v_68438 | v_68442;
assign v_68445 = v_68421 | v_68444;
assign v_68447 = v_68419 | v_68446;
assign v_68449 = v_68444 | v_68448;
assign v_68451 = v_68418 | v_68450;
assign v_68453 = v_68416 | v_68452;
assign v_68455 = v_68450 | v_68454;
assign v_68457 = v_68415 | v_68456;
assign v_68459 = v_68413 | v_68458;
assign v_68461 = v_68456 | v_68460;
assign v_68463 = v_68412 | v_68462;
assign v_68465 = v_68410 | v_68464;
assign v_68467 = v_68462 | v_68466;
assign v_68469 = v_68409 | v_68468;
assign v_68471 = v_68407 | v_68470;
assign v_68473 = v_68468 | v_68472;
assign v_68475 = v_68406 | v_68474;
assign v_68477 = v_68404 | v_68476;
assign v_68479 = v_68474 | v_68478;
assign v_68481 = v_68403 | v_68480;
assign v_68483 = v_68401 | v_68482;
assign v_68485 = v_68480 | v_68484;
assign v_68487 = v_68400 | v_68486;
assign v_68489 = v_68398 | v_68488;
assign v_68491 = v_68486 | v_68490;
assign v_68493 = v_68397 | v_68492;
assign v_68495 = v_68395 | v_68494;
assign v_68497 = v_68492 | v_68496;
assign v_68499 = v_68394 | v_68498;
assign v_68501 = v_68392 | v_68500;
assign v_68503 = v_68498 | v_68502;
assign v_68505 = v_68391 | v_68504;
assign v_68507 = v_68389 | v_68506;
assign v_68509 = v_68504 | v_68508;
assign v_68511 = v_68388 | v_68510;
assign v_68513 = v_68386 | v_68512;
assign v_68515 = v_68510 | v_68514;
assign v_68517 = v_68385 | v_68516;
assign v_68519 = v_68383 | v_68518;
assign v_68521 = v_68516 | v_68520;
assign v_68523 = v_68382 | v_68522;
assign v_68525 = v_68380 | v_68524;
assign v_68527 = v_68522 | v_68526;
assign v_68531 = v_68528 | v_68530;
assign v_68538 = v_68427 | v_68537;
assign v_68541 = v_68539 | v_68540;
assign v_68543 = v_68424 | v_68542;
assign v_68546 = v_68544 | v_68545;
assign v_68548 = v_68421 | v_68547;
assign v_68551 = v_68549 | v_68550;
assign v_68553 = v_68418 | v_68552;
assign v_68556 = v_68554 | v_68555;
assign v_68558 = v_68415 | v_68557;
assign v_68561 = v_68559 | v_68560;
assign v_68563 = v_68412 | v_68562;
assign v_68566 = v_68564 | v_68565;
assign v_68568 = v_68409 | v_68567;
assign v_68571 = v_68569 | v_68570;
assign v_68573 = v_68406 | v_68572;
assign v_68576 = v_68574 | v_68575;
assign v_68578 = v_68403 | v_68577;
assign v_68581 = v_68579 | v_68580;
assign v_68583 = v_68400 | v_68582;
assign v_68586 = v_68584 | v_68585;
assign v_68588 = v_68397 | v_68587;
assign v_68591 = v_68589 | v_68590;
assign v_68593 = v_68394 | v_68592;
assign v_68596 = v_68594 | v_68595;
assign v_68598 = v_68391 | v_68597;
assign v_68601 = v_68599 | v_68600;
assign v_68603 = v_68388 | v_68602;
assign v_68606 = v_68604 | v_68605;
assign v_68608 = v_68385 | v_68607;
assign v_68611 = v_68609 | v_68610;
assign v_68613 = v_68382 | v_68612;
assign v_68616 = v_68614 | v_68615;
assign v_68618 = v_68616 | v_68617;
assign v_68621 = v_68379 | v_68620;
assign v_68674 = v_68671 | v_68673;
assign v_68676 = v_68670 | v_68675;
assign v_68678 = v_68668 | v_68677;
assign v_68680 = v_68675 | v_68679;
assign v_68682 = v_68667 | v_68681;
assign v_68684 = v_68665 | v_68683;
assign v_68686 = v_68681 | v_68685;
assign v_68688 = v_68664 | v_68687;
assign v_68690 = v_68662 | v_68689;
assign v_68692 = v_68687 | v_68691;
assign v_68694 = v_68661 | v_68693;
assign v_68696 = v_68659 | v_68695;
assign v_68698 = v_68693 | v_68697;
assign v_68700 = v_68658 | v_68699;
assign v_68702 = v_68656 | v_68701;
assign v_68704 = v_68699 | v_68703;
assign v_68706 = v_68655 | v_68705;
assign v_68708 = v_68653 | v_68707;
assign v_68710 = v_68705 | v_68709;
assign v_68712 = v_68652 | v_68711;
assign v_68714 = v_68650 | v_68713;
assign v_68716 = v_68711 | v_68715;
assign v_68718 = v_68649 | v_68717;
assign v_68720 = v_68647 | v_68719;
assign v_68722 = v_68717 | v_68721;
assign v_68724 = v_68646 | v_68723;
assign v_68726 = v_68644 | v_68725;
assign v_68728 = v_68723 | v_68727;
assign v_68730 = v_68643 | v_68729;
assign v_68732 = v_68641 | v_68731;
assign v_68734 = v_68729 | v_68733;
assign v_68736 = v_68640 | v_68735;
assign v_68738 = v_68638 | v_68737;
assign v_68740 = v_68735 | v_68739;
assign v_68742 = v_68637 | v_68741;
assign v_68744 = v_68635 | v_68743;
assign v_68746 = v_68741 | v_68745;
assign v_68748 = v_68634 | v_68747;
assign v_68750 = v_68632 | v_68749;
assign v_68752 = v_68747 | v_68751;
assign v_68754 = v_68631 | v_68753;
assign v_68756 = v_68629 | v_68755;
assign v_68758 = v_68753 | v_68757;
assign v_68760 = v_68628 | v_68759;
assign v_68762 = v_68626 | v_68761;
assign v_68764 = v_68759 | v_68763;
assign v_68766 = v_68625 | v_68765;
assign v_68768 = v_68623 | v_68767;
assign v_68770 = v_68765 | v_68769;
assign v_68774 = v_68771 | v_68773;
assign v_68781 = v_68670 | v_68780;
assign v_68784 = v_68782 | v_68783;
assign v_68786 = v_68667 | v_68785;
assign v_68789 = v_68787 | v_68788;
assign v_68791 = v_68664 | v_68790;
assign v_68794 = v_68792 | v_68793;
assign v_68796 = v_68661 | v_68795;
assign v_68799 = v_68797 | v_68798;
assign v_68801 = v_68658 | v_68800;
assign v_68804 = v_68802 | v_68803;
assign v_68806 = v_68655 | v_68805;
assign v_68809 = v_68807 | v_68808;
assign v_68811 = v_68652 | v_68810;
assign v_68814 = v_68812 | v_68813;
assign v_68816 = v_68649 | v_68815;
assign v_68819 = v_68817 | v_68818;
assign v_68821 = v_68646 | v_68820;
assign v_68824 = v_68822 | v_68823;
assign v_68826 = v_68643 | v_68825;
assign v_68829 = v_68827 | v_68828;
assign v_68831 = v_68640 | v_68830;
assign v_68834 = v_68832 | v_68833;
assign v_68836 = v_68637 | v_68835;
assign v_68839 = v_68837 | v_68838;
assign v_68841 = v_68634 | v_68840;
assign v_68844 = v_68842 | v_68843;
assign v_68846 = v_68631 | v_68845;
assign v_68849 = v_68847 | v_68848;
assign v_68851 = v_68628 | v_68850;
assign v_68854 = v_68852 | v_68853;
assign v_68856 = v_68625 | v_68855;
assign v_68859 = v_68857 | v_68858;
assign v_68861 = v_68859 | v_68860;
assign v_68864 = v_68622 | v_68863;
assign v_68917 = v_68914 | v_68916;
assign v_68919 = v_68913 | v_68918;
assign v_68921 = v_68911 | v_68920;
assign v_68923 = v_68918 | v_68922;
assign v_68925 = v_68910 | v_68924;
assign v_68927 = v_68908 | v_68926;
assign v_68929 = v_68924 | v_68928;
assign v_68931 = v_68907 | v_68930;
assign v_68933 = v_68905 | v_68932;
assign v_68935 = v_68930 | v_68934;
assign v_68937 = v_68904 | v_68936;
assign v_68939 = v_68902 | v_68938;
assign v_68941 = v_68936 | v_68940;
assign v_68943 = v_68901 | v_68942;
assign v_68945 = v_68899 | v_68944;
assign v_68947 = v_68942 | v_68946;
assign v_68949 = v_68898 | v_68948;
assign v_68951 = v_68896 | v_68950;
assign v_68953 = v_68948 | v_68952;
assign v_68955 = v_68895 | v_68954;
assign v_68957 = v_68893 | v_68956;
assign v_68959 = v_68954 | v_68958;
assign v_68961 = v_68892 | v_68960;
assign v_68963 = v_68890 | v_68962;
assign v_68965 = v_68960 | v_68964;
assign v_68967 = v_68889 | v_68966;
assign v_68969 = v_68887 | v_68968;
assign v_68971 = v_68966 | v_68970;
assign v_68973 = v_68886 | v_68972;
assign v_68975 = v_68884 | v_68974;
assign v_68977 = v_68972 | v_68976;
assign v_68979 = v_68883 | v_68978;
assign v_68981 = v_68881 | v_68980;
assign v_68983 = v_68978 | v_68982;
assign v_68985 = v_68880 | v_68984;
assign v_68987 = v_68878 | v_68986;
assign v_68989 = v_68984 | v_68988;
assign v_68991 = v_68877 | v_68990;
assign v_68993 = v_68875 | v_68992;
assign v_68995 = v_68990 | v_68994;
assign v_68997 = v_68874 | v_68996;
assign v_68999 = v_68872 | v_68998;
assign v_69001 = v_68996 | v_69000;
assign v_69003 = v_68871 | v_69002;
assign v_69005 = v_68869 | v_69004;
assign v_69007 = v_69002 | v_69006;
assign v_69009 = v_68868 | v_69008;
assign v_69011 = v_68866 | v_69010;
assign v_69013 = v_69008 | v_69012;
assign v_69017 = v_69014 | v_69016;
assign v_69024 = v_68913 | v_69023;
assign v_69027 = v_69025 | v_69026;
assign v_69029 = v_68910 | v_69028;
assign v_69032 = v_69030 | v_69031;
assign v_69034 = v_68907 | v_69033;
assign v_69037 = v_69035 | v_69036;
assign v_69039 = v_68904 | v_69038;
assign v_69042 = v_69040 | v_69041;
assign v_69044 = v_68901 | v_69043;
assign v_69047 = v_69045 | v_69046;
assign v_69049 = v_68898 | v_69048;
assign v_69052 = v_69050 | v_69051;
assign v_69054 = v_68895 | v_69053;
assign v_69057 = v_69055 | v_69056;
assign v_69059 = v_68892 | v_69058;
assign v_69062 = v_69060 | v_69061;
assign v_69064 = v_68889 | v_69063;
assign v_69067 = v_69065 | v_69066;
assign v_69069 = v_68886 | v_69068;
assign v_69072 = v_69070 | v_69071;
assign v_69074 = v_68883 | v_69073;
assign v_69077 = v_69075 | v_69076;
assign v_69079 = v_68880 | v_69078;
assign v_69082 = v_69080 | v_69081;
assign v_69084 = v_68877 | v_69083;
assign v_69087 = v_69085 | v_69086;
assign v_69089 = v_68874 | v_69088;
assign v_69092 = v_69090 | v_69091;
assign v_69094 = v_68871 | v_69093;
assign v_69097 = v_69095 | v_69096;
assign v_69099 = v_68868 | v_69098;
assign v_69102 = v_69100 | v_69101;
assign v_69104 = v_69102 | v_69103;
assign v_69107 = v_68865 | v_69106;
assign v_69160 = v_69157 | v_69159;
assign v_69162 = v_69156 | v_69161;
assign v_69164 = v_69154 | v_69163;
assign v_69166 = v_69161 | v_69165;
assign v_69168 = v_69153 | v_69167;
assign v_69170 = v_69151 | v_69169;
assign v_69172 = v_69167 | v_69171;
assign v_69174 = v_69150 | v_69173;
assign v_69176 = v_69148 | v_69175;
assign v_69178 = v_69173 | v_69177;
assign v_69180 = v_69147 | v_69179;
assign v_69182 = v_69145 | v_69181;
assign v_69184 = v_69179 | v_69183;
assign v_69186 = v_69144 | v_69185;
assign v_69188 = v_69142 | v_69187;
assign v_69190 = v_69185 | v_69189;
assign v_69192 = v_69141 | v_69191;
assign v_69194 = v_69139 | v_69193;
assign v_69196 = v_69191 | v_69195;
assign v_69198 = v_69138 | v_69197;
assign v_69200 = v_69136 | v_69199;
assign v_69202 = v_69197 | v_69201;
assign v_69204 = v_69135 | v_69203;
assign v_69206 = v_69133 | v_69205;
assign v_69208 = v_69203 | v_69207;
assign v_69210 = v_69132 | v_69209;
assign v_69212 = v_69130 | v_69211;
assign v_69214 = v_69209 | v_69213;
assign v_69216 = v_69129 | v_69215;
assign v_69218 = v_69127 | v_69217;
assign v_69220 = v_69215 | v_69219;
assign v_69222 = v_69126 | v_69221;
assign v_69224 = v_69124 | v_69223;
assign v_69226 = v_69221 | v_69225;
assign v_69228 = v_69123 | v_69227;
assign v_69230 = v_69121 | v_69229;
assign v_69232 = v_69227 | v_69231;
assign v_69234 = v_69120 | v_69233;
assign v_69236 = v_69118 | v_69235;
assign v_69238 = v_69233 | v_69237;
assign v_69240 = v_69117 | v_69239;
assign v_69242 = v_69115 | v_69241;
assign v_69244 = v_69239 | v_69243;
assign v_69246 = v_69114 | v_69245;
assign v_69248 = v_69112 | v_69247;
assign v_69250 = v_69245 | v_69249;
assign v_69252 = v_69111 | v_69251;
assign v_69254 = v_69109 | v_69253;
assign v_69256 = v_69251 | v_69255;
assign v_69260 = v_69257 | v_69259;
assign v_69267 = v_69156 | v_69266;
assign v_69270 = v_69268 | v_69269;
assign v_69272 = v_69153 | v_69271;
assign v_69275 = v_69273 | v_69274;
assign v_69277 = v_69150 | v_69276;
assign v_69280 = v_69278 | v_69279;
assign v_69282 = v_69147 | v_69281;
assign v_69285 = v_69283 | v_69284;
assign v_69287 = v_69144 | v_69286;
assign v_69290 = v_69288 | v_69289;
assign v_69292 = v_69141 | v_69291;
assign v_69295 = v_69293 | v_69294;
assign v_69297 = v_69138 | v_69296;
assign v_69300 = v_69298 | v_69299;
assign v_69302 = v_69135 | v_69301;
assign v_69305 = v_69303 | v_69304;
assign v_69307 = v_69132 | v_69306;
assign v_69310 = v_69308 | v_69309;
assign v_69312 = v_69129 | v_69311;
assign v_69315 = v_69313 | v_69314;
assign v_69317 = v_69126 | v_69316;
assign v_69320 = v_69318 | v_69319;
assign v_69322 = v_69123 | v_69321;
assign v_69325 = v_69323 | v_69324;
assign v_69327 = v_69120 | v_69326;
assign v_69330 = v_69328 | v_69329;
assign v_69332 = v_69117 | v_69331;
assign v_69335 = v_69333 | v_69334;
assign v_69337 = v_69114 | v_69336;
assign v_69340 = v_69338 | v_69339;
assign v_69342 = v_69111 | v_69341;
assign v_69345 = v_69343 | v_69344;
assign v_69347 = v_69345 | v_69346;
assign v_69350 = v_69108 | v_69349;
assign v_69403 = v_69400 | v_69402;
assign v_69405 = v_69399 | v_69404;
assign v_69407 = v_69397 | v_69406;
assign v_69409 = v_69404 | v_69408;
assign v_69411 = v_69396 | v_69410;
assign v_69413 = v_69394 | v_69412;
assign v_69415 = v_69410 | v_69414;
assign v_69417 = v_69393 | v_69416;
assign v_69419 = v_69391 | v_69418;
assign v_69421 = v_69416 | v_69420;
assign v_69423 = v_69390 | v_69422;
assign v_69425 = v_69388 | v_69424;
assign v_69427 = v_69422 | v_69426;
assign v_69429 = v_69387 | v_69428;
assign v_69431 = v_69385 | v_69430;
assign v_69433 = v_69428 | v_69432;
assign v_69435 = v_69384 | v_69434;
assign v_69437 = v_69382 | v_69436;
assign v_69439 = v_69434 | v_69438;
assign v_69441 = v_69381 | v_69440;
assign v_69443 = v_69379 | v_69442;
assign v_69445 = v_69440 | v_69444;
assign v_69447 = v_69378 | v_69446;
assign v_69449 = v_69376 | v_69448;
assign v_69451 = v_69446 | v_69450;
assign v_69453 = v_69375 | v_69452;
assign v_69455 = v_69373 | v_69454;
assign v_69457 = v_69452 | v_69456;
assign v_69459 = v_69372 | v_69458;
assign v_69461 = v_69370 | v_69460;
assign v_69463 = v_69458 | v_69462;
assign v_69465 = v_69369 | v_69464;
assign v_69467 = v_69367 | v_69466;
assign v_69469 = v_69464 | v_69468;
assign v_69471 = v_69366 | v_69470;
assign v_69473 = v_69364 | v_69472;
assign v_69475 = v_69470 | v_69474;
assign v_69477 = v_69363 | v_69476;
assign v_69479 = v_69361 | v_69478;
assign v_69481 = v_69476 | v_69480;
assign v_69483 = v_69360 | v_69482;
assign v_69485 = v_69358 | v_69484;
assign v_69487 = v_69482 | v_69486;
assign v_69489 = v_69357 | v_69488;
assign v_69491 = v_69355 | v_69490;
assign v_69493 = v_69488 | v_69492;
assign v_69495 = v_69354 | v_69494;
assign v_69497 = v_69352 | v_69496;
assign v_69499 = v_69494 | v_69498;
assign v_69503 = v_69500 | v_69502;
assign v_69510 = v_69399 | v_69509;
assign v_69513 = v_69511 | v_69512;
assign v_69515 = v_69396 | v_69514;
assign v_69518 = v_69516 | v_69517;
assign v_69520 = v_69393 | v_69519;
assign v_69523 = v_69521 | v_69522;
assign v_69525 = v_69390 | v_69524;
assign v_69528 = v_69526 | v_69527;
assign v_69530 = v_69387 | v_69529;
assign v_69533 = v_69531 | v_69532;
assign v_69535 = v_69384 | v_69534;
assign v_69538 = v_69536 | v_69537;
assign v_69540 = v_69381 | v_69539;
assign v_69543 = v_69541 | v_69542;
assign v_69545 = v_69378 | v_69544;
assign v_69548 = v_69546 | v_69547;
assign v_69550 = v_69375 | v_69549;
assign v_69553 = v_69551 | v_69552;
assign v_69555 = v_69372 | v_69554;
assign v_69558 = v_69556 | v_69557;
assign v_69560 = v_69369 | v_69559;
assign v_69563 = v_69561 | v_69562;
assign v_69565 = v_69366 | v_69564;
assign v_69568 = v_69566 | v_69567;
assign v_69570 = v_69363 | v_69569;
assign v_69573 = v_69571 | v_69572;
assign v_69575 = v_69360 | v_69574;
assign v_69578 = v_69576 | v_69577;
assign v_69580 = v_69357 | v_69579;
assign v_69583 = v_69581 | v_69582;
assign v_69585 = v_69354 | v_69584;
assign v_69588 = v_69586 | v_69587;
assign v_69590 = v_69588 | v_69589;
assign v_69593 = v_69351 | v_69592;
assign v_69646 = v_69643 | v_69645;
assign v_69648 = v_69642 | v_69647;
assign v_69650 = v_69640 | v_69649;
assign v_69652 = v_69647 | v_69651;
assign v_69654 = v_69639 | v_69653;
assign v_69656 = v_69637 | v_69655;
assign v_69658 = v_69653 | v_69657;
assign v_69660 = v_69636 | v_69659;
assign v_69662 = v_69634 | v_69661;
assign v_69664 = v_69659 | v_69663;
assign v_69666 = v_69633 | v_69665;
assign v_69668 = v_69631 | v_69667;
assign v_69670 = v_69665 | v_69669;
assign v_69672 = v_69630 | v_69671;
assign v_69674 = v_69628 | v_69673;
assign v_69676 = v_69671 | v_69675;
assign v_69678 = v_69627 | v_69677;
assign v_69680 = v_69625 | v_69679;
assign v_69682 = v_69677 | v_69681;
assign v_69684 = v_69624 | v_69683;
assign v_69686 = v_69622 | v_69685;
assign v_69688 = v_69683 | v_69687;
assign v_69690 = v_69621 | v_69689;
assign v_69692 = v_69619 | v_69691;
assign v_69694 = v_69689 | v_69693;
assign v_69696 = v_69618 | v_69695;
assign v_69698 = v_69616 | v_69697;
assign v_69700 = v_69695 | v_69699;
assign v_69702 = v_69615 | v_69701;
assign v_69704 = v_69613 | v_69703;
assign v_69706 = v_69701 | v_69705;
assign v_69708 = v_69612 | v_69707;
assign v_69710 = v_69610 | v_69709;
assign v_69712 = v_69707 | v_69711;
assign v_69714 = v_69609 | v_69713;
assign v_69716 = v_69607 | v_69715;
assign v_69718 = v_69713 | v_69717;
assign v_69720 = v_69606 | v_69719;
assign v_69722 = v_69604 | v_69721;
assign v_69724 = v_69719 | v_69723;
assign v_69726 = v_69603 | v_69725;
assign v_69728 = v_69601 | v_69727;
assign v_69730 = v_69725 | v_69729;
assign v_69732 = v_69600 | v_69731;
assign v_69734 = v_69598 | v_69733;
assign v_69736 = v_69731 | v_69735;
assign v_69738 = v_69597 | v_69737;
assign v_69740 = v_69595 | v_69739;
assign v_69742 = v_69737 | v_69741;
assign v_69746 = v_69743 | v_69745;
assign v_69753 = v_69642 | v_69752;
assign v_69756 = v_69754 | v_69755;
assign v_69758 = v_69639 | v_69757;
assign v_69761 = v_69759 | v_69760;
assign v_69763 = v_69636 | v_69762;
assign v_69766 = v_69764 | v_69765;
assign v_69768 = v_69633 | v_69767;
assign v_69771 = v_69769 | v_69770;
assign v_69773 = v_69630 | v_69772;
assign v_69776 = v_69774 | v_69775;
assign v_69778 = v_69627 | v_69777;
assign v_69781 = v_69779 | v_69780;
assign v_69783 = v_69624 | v_69782;
assign v_69786 = v_69784 | v_69785;
assign v_69788 = v_69621 | v_69787;
assign v_69791 = v_69789 | v_69790;
assign v_69793 = v_69618 | v_69792;
assign v_69796 = v_69794 | v_69795;
assign v_69798 = v_69615 | v_69797;
assign v_69801 = v_69799 | v_69800;
assign v_69803 = v_69612 | v_69802;
assign v_69806 = v_69804 | v_69805;
assign v_69808 = v_69609 | v_69807;
assign v_69811 = v_69809 | v_69810;
assign v_69813 = v_69606 | v_69812;
assign v_69816 = v_69814 | v_69815;
assign v_69818 = v_69603 | v_69817;
assign v_69821 = v_69819 | v_69820;
assign v_69823 = v_69600 | v_69822;
assign v_69826 = v_69824 | v_69825;
assign v_69828 = v_69597 | v_69827;
assign v_69831 = v_69829 | v_69830;
assign v_69833 = v_69831 | v_69832;
assign v_69836 = v_69594 | v_69835;
assign v_69889 = v_69886 | v_69888;
assign v_69891 = v_69885 | v_69890;
assign v_69893 = v_69883 | v_69892;
assign v_69895 = v_69890 | v_69894;
assign v_69897 = v_69882 | v_69896;
assign v_69899 = v_69880 | v_69898;
assign v_69901 = v_69896 | v_69900;
assign v_69903 = v_69879 | v_69902;
assign v_69905 = v_69877 | v_69904;
assign v_69907 = v_69902 | v_69906;
assign v_69909 = v_69876 | v_69908;
assign v_69911 = v_69874 | v_69910;
assign v_69913 = v_69908 | v_69912;
assign v_69915 = v_69873 | v_69914;
assign v_69917 = v_69871 | v_69916;
assign v_69919 = v_69914 | v_69918;
assign v_69921 = v_69870 | v_69920;
assign v_69923 = v_69868 | v_69922;
assign v_69925 = v_69920 | v_69924;
assign v_69927 = v_69867 | v_69926;
assign v_69929 = v_69865 | v_69928;
assign v_69931 = v_69926 | v_69930;
assign v_69933 = v_69864 | v_69932;
assign v_69935 = v_69862 | v_69934;
assign v_69937 = v_69932 | v_69936;
assign v_69939 = v_69861 | v_69938;
assign v_69941 = v_69859 | v_69940;
assign v_69943 = v_69938 | v_69942;
assign v_69945 = v_69858 | v_69944;
assign v_69947 = v_69856 | v_69946;
assign v_69949 = v_69944 | v_69948;
assign v_69951 = v_69855 | v_69950;
assign v_69953 = v_69853 | v_69952;
assign v_69955 = v_69950 | v_69954;
assign v_69957 = v_69852 | v_69956;
assign v_69959 = v_69850 | v_69958;
assign v_69961 = v_69956 | v_69960;
assign v_69963 = v_69849 | v_69962;
assign v_69965 = v_69847 | v_69964;
assign v_69967 = v_69962 | v_69966;
assign v_69969 = v_69846 | v_69968;
assign v_69971 = v_69844 | v_69970;
assign v_69973 = v_69968 | v_69972;
assign v_69975 = v_69843 | v_69974;
assign v_69977 = v_69841 | v_69976;
assign v_69979 = v_69974 | v_69978;
assign v_69981 = v_69840 | v_69980;
assign v_69983 = v_69838 | v_69982;
assign v_69985 = v_69980 | v_69984;
assign v_69989 = v_69986 | v_69988;
assign v_69996 = v_69885 | v_69995;
assign v_69999 = v_69997 | v_69998;
assign v_70001 = v_69882 | v_70000;
assign v_70004 = v_70002 | v_70003;
assign v_70006 = v_69879 | v_70005;
assign v_70009 = v_70007 | v_70008;
assign v_70011 = v_69876 | v_70010;
assign v_70014 = v_70012 | v_70013;
assign v_70016 = v_69873 | v_70015;
assign v_70019 = v_70017 | v_70018;
assign v_70021 = v_69870 | v_70020;
assign v_70024 = v_70022 | v_70023;
assign v_70026 = v_69867 | v_70025;
assign v_70029 = v_70027 | v_70028;
assign v_70031 = v_69864 | v_70030;
assign v_70034 = v_70032 | v_70033;
assign v_70036 = v_69861 | v_70035;
assign v_70039 = v_70037 | v_70038;
assign v_70041 = v_69858 | v_70040;
assign v_70044 = v_70042 | v_70043;
assign v_70046 = v_69855 | v_70045;
assign v_70049 = v_70047 | v_70048;
assign v_70051 = v_69852 | v_70050;
assign v_70054 = v_70052 | v_70053;
assign v_70056 = v_69849 | v_70055;
assign v_70059 = v_70057 | v_70058;
assign v_70061 = v_69846 | v_70060;
assign v_70064 = v_70062 | v_70063;
assign v_70066 = v_69843 | v_70065;
assign v_70069 = v_70067 | v_70068;
assign v_70071 = v_69840 | v_70070;
assign v_70074 = v_70072 | v_70073;
assign v_70076 = v_70074 | v_70075;
assign v_70079 = v_69837 | v_70078;
assign v_70132 = v_70129 | v_70131;
assign v_70134 = v_70128 | v_70133;
assign v_70136 = v_70126 | v_70135;
assign v_70138 = v_70133 | v_70137;
assign v_70140 = v_70125 | v_70139;
assign v_70142 = v_70123 | v_70141;
assign v_70144 = v_70139 | v_70143;
assign v_70146 = v_70122 | v_70145;
assign v_70148 = v_70120 | v_70147;
assign v_70150 = v_70145 | v_70149;
assign v_70152 = v_70119 | v_70151;
assign v_70154 = v_70117 | v_70153;
assign v_70156 = v_70151 | v_70155;
assign v_70158 = v_70116 | v_70157;
assign v_70160 = v_70114 | v_70159;
assign v_70162 = v_70157 | v_70161;
assign v_70164 = v_70113 | v_70163;
assign v_70166 = v_70111 | v_70165;
assign v_70168 = v_70163 | v_70167;
assign v_70170 = v_70110 | v_70169;
assign v_70172 = v_70108 | v_70171;
assign v_70174 = v_70169 | v_70173;
assign v_70176 = v_70107 | v_70175;
assign v_70178 = v_70105 | v_70177;
assign v_70180 = v_70175 | v_70179;
assign v_70182 = v_70104 | v_70181;
assign v_70184 = v_70102 | v_70183;
assign v_70186 = v_70181 | v_70185;
assign v_70188 = v_70101 | v_70187;
assign v_70190 = v_70099 | v_70189;
assign v_70192 = v_70187 | v_70191;
assign v_70194 = v_70098 | v_70193;
assign v_70196 = v_70096 | v_70195;
assign v_70198 = v_70193 | v_70197;
assign v_70200 = v_70095 | v_70199;
assign v_70202 = v_70093 | v_70201;
assign v_70204 = v_70199 | v_70203;
assign v_70206 = v_70092 | v_70205;
assign v_70208 = v_70090 | v_70207;
assign v_70210 = v_70205 | v_70209;
assign v_70212 = v_70089 | v_70211;
assign v_70214 = v_70087 | v_70213;
assign v_70216 = v_70211 | v_70215;
assign v_70218 = v_70086 | v_70217;
assign v_70220 = v_70084 | v_70219;
assign v_70222 = v_70217 | v_70221;
assign v_70224 = v_70083 | v_70223;
assign v_70226 = v_70081 | v_70225;
assign v_70228 = v_70223 | v_70227;
assign v_70232 = v_70229 | v_70231;
assign v_70239 = v_70128 | v_70238;
assign v_70242 = v_70240 | v_70241;
assign v_70244 = v_70125 | v_70243;
assign v_70247 = v_70245 | v_70246;
assign v_70249 = v_70122 | v_70248;
assign v_70252 = v_70250 | v_70251;
assign v_70254 = v_70119 | v_70253;
assign v_70257 = v_70255 | v_70256;
assign v_70259 = v_70116 | v_70258;
assign v_70262 = v_70260 | v_70261;
assign v_70264 = v_70113 | v_70263;
assign v_70267 = v_70265 | v_70266;
assign v_70269 = v_70110 | v_70268;
assign v_70272 = v_70270 | v_70271;
assign v_70274 = v_70107 | v_70273;
assign v_70277 = v_70275 | v_70276;
assign v_70279 = v_70104 | v_70278;
assign v_70282 = v_70280 | v_70281;
assign v_70284 = v_70101 | v_70283;
assign v_70287 = v_70285 | v_70286;
assign v_70289 = v_70098 | v_70288;
assign v_70292 = v_70290 | v_70291;
assign v_70294 = v_70095 | v_70293;
assign v_70297 = v_70295 | v_70296;
assign v_70299 = v_70092 | v_70298;
assign v_70302 = v_70300 | v_70301;
assign v_70304 = v_70089 | v_70303;
assign v_70307 = v_70305 | v_70306;
assign v_70309 = v_70086 | v_70308;
assign v_70312 = v_70310 | v_70311;
assign v_70314 = v_70083 | v_70313;
assign v_70317 = v_70315 | v_70316;
assign v_70319 = v_70317 | v_70318;
assign v_70322 = v_70080 | v_70321;
assign v_70375 = v_70372 | v_70374;
assign v_70377 = v_70371 | v_70376;
assign v_70379 = v_70369 | v_70378;
assign v_70381 = v_70376 | v_70380;
assign v_70383 = v_70368 | v_70382;
assign v_70385 = v_70366 | v_70384;
assign v_70387 = v_70382 | v_70386;
assign v_70389 = v_70365 | v_70388;
assign v_70391 = v_70363 | v_70390;
assign v_70393 = v_70388 | v_70392;
assign v_70395 = v_70362 | v_70394;
assign v_70397 = v_70360 | v_70396;
assign v_70399 = v_70394 | v_70398;
assign v_70401 = v_70359 | v_70400;
assign v_70403 = v_70357 | v_70402;
assign v_70405 = v_70400 | v_70404;
assign v_70407 = v_70356 | v_70406;
assign v_70409 = v_70354 | v_70408;
assign v_70411 = v_70406 | v_70410;
assign v_70413 = v_70353 | v_70412;
assign v_70415 = v_70351 | v_70414;
assign v_70417 = v_70412 | v_70416;
assign v_70419 = v_70350 | v_70418;
assign v_70421 = v_70348 | v_70420;
assign v_70423 = v_70418 | v_70422;
assign v_70425 = v_70347 | v_70424;
assign v_70427 = v_70345 | v_70426;
assign v_70429 = v_70424 | v_70428;
assign v_70431 = v_70344 | v_70430;
assign v_70433 = v_70342 | v_70432;
assign v_70435 = v_70430 | v_70434;
assign v_70437 = v_70341 | v_70436;
assign v_70439 = v_70339 | v_70438;
assign v_70441 = v_70436 | v_70440;
assign v_70443 = v_70338 | v_70442;
assign v_70445 = v_70336 | v_70444;
assign v_70447 = v_70442 | v_70446;
assign v_70449 = v_70335 | v_70448;
assign v_70451 = v_70333 | v_70450;
assign v_70453 = v_70448 | v_70452;
assign v_70455 = v_70332 | v_70454;
assign v_70457 = v_70330 | v_70456;
assign v_70459 = v_70454 | v_70458;
assign v_70461 = v_70329 | v_70460;
assign v_70463 = v_70327 | v_70462;
assign v_70465 = v_70460 | v_70464;
assign v_70467 = v_70326 | v_70466;
assign v_70469 = v_70324 | v_70468;
assign v_70471 = v_70466 | v_70470;
assign v_70475 = v_70472 | v_70474;
assign v_70482 = v_70371 | v_70481;
assign v_70485 = v_70483 | v_70484;
assign v_70487 = v_70368 | v_70486;
assign v_70490 = v_70488 | v_70489;
assign v_70492 = v_70365 | v_70491;
assign v_70495 = v_70493 | v_70494;
assign v_70497 = v_70362 | v_70496;
assign v_70500 = v_70498 | v_70499;
assign v_70502 = v_70359 | v_70501;
assign v_70505 = v_70503 | v_70504;
assign v_70507 = v_70356 | v_70506;
assign v_70510 = v_70508 | v_70509;
assign v_70512 = v_70353 | v_70511;
assign v_70515 = v_70513 | v_70514;
assign v_70517 = v_70350 | v_70516;
assign v_70520 = v_70518 | v_70519;
assign v_70522 = v_70347 | v_70521;
assign v_70525 = v_70523 | v_70524;
assign v_70527 = v_70344 | v_70526;
assign v_70530 = v_70528 | v_70529;
assign v_70532 = v_70341 | v_70531;
assign v_70535 = v_70533 | v_70534;
assign v_70537 = v_70338 | v_70536;
assign v_70540 = v_70538 | v_70539;
assign v_70542 = v_70335 | v_70541;
assign v_70545 = v_70543 | v_70544;
assign v_70547 = v_70332 | v_70546;
assign v_70550 = v_70548 | v_70549;
assign v_70552 = v_70329 | v_70551;
assign v_70555 = v_70553 | v_70554;
assign v_70557 = v_70326 | v_70556;
assign v_70560 = v_70558 | v_70559;
assign v_70562 = v_70560 | v_70561;
assign v_70565 = v_70323 | v_70564;
assign v_70618 = v_70615 | v_70617;
assign v_70620 = v_70614 | v_70619;
assign v_70622 = v_70612 | v_70621;
assign v_70624 = v_70619 | v_70623;
assign v_70626 = v_70611 | v_70625;
assign v_70628 = v_70609 | v_70627;
assign v_70630 = v_70625 | v_70629;
assign v_70632 = v_70608 | v_70631;
assign v_70634 = v_70606 | v_70633;
assign v_70636 = v_70631 | v_70635;
assign v_70638 = v_70605 | v_70637;
assign v_70640 = v_70603 | v_70639;
assign v_70642 = v_70637 | v_70641;
assign v_70644 = v_70602 | v_70643;
assign v_70646 = v_70600 | v_70645;
assign v_70648 = v_70643 | v_70647;
assign v_70650 = v_70599 | v_70649;
assign v_70652 = v_70597 | v_70651;
assign v_70654 = v_70649 | v_70653;
assign v_70656 = v_70596 | v_70655;
assign v_70658 = v_70594 | v_70657;
assign v_70660 = v_70655 | v_70659;
assign v_70662 = v_70593 | v_70661;
assign v_70664 = v_70591 | v_70663;
assign v_70666 = v_70661 | v_70665;
assign v_70668 = v_70590 | v_70667;
assign v_70670 = v_70588 | v_70669;
assign v_70672 = v_70667 | v_70671;
assign v_70674 = v_70587 | v_70673;
assign v_70676 = v_70585 | v_70675;
assign v_70678 = v_70673 | v_70677;
assign v_70680 = v_70584 | v_70679;
assign v_70682 = v_70582 | v_70681;
assign v_70684 = v_70679 | v_70683;
assign v_70686 = v_70581 | v_70685;
assign v_70688 = v_70579 | v_70687;
assign v_70690 = v_70685 | v_70689;
assign v_70692 = v_70578 | v_70691;
assign v_70694 = v_70576 | v_70693;
assign v_70696 = v_70691 | v_70695;
assign v_70698 = v_70575 | v_70697;
assign v_70700 = v_70573 | v_70699;
assign v_70702 = v_70697 | v_70701;
assign v_70704 = v_70572 | v_70703;
assign v_70706 = v_70570 | v_70705;
assign v_70708 = v_70703 | v_70707;
assign v_70710 = v_70569 | v_70709;
assign v_70712 = v_70567 | v_70711;
assign v_70714 = v_70709 | v_70713;
assign v_70718 = v_70715 | v_70717;
assign v_70725 = v_70614 | v_70724;
assign v_70728 = v_70726 | v_70727;
assign v_70730 = v_70611 | v_70729;
assign v_70733 = v_70731 | v_70732;
assign v_70735 = v_70608 | v_70734;
assign v_70738 = v_70736 | v_70737;
assign v_70740 = v_70605 | v_70739;
assign v_70743 = v_70741 | v_70742;
assign v_70745 = v_70602 | v_70744;
assign v_70748 = v_70746 | v_70747;
assign v_70750 = v_70599 | v_70749;
assign v_70753 = v_70751 | v_70752;
assign v_70755 = v_70596 | v_70754;
assign v_70758 = v_70756 | v_70757;
assign v_70760 = v_70593 | v_70759;
assign v_70763 = v_70761 | v_70762;
assign v_70765 = v_70590 | v_70764;
assign v_70768 = v_70766 | v_70767;
assign v_70770 = v_70587 | v_70769;
assign v_70773 = v_70771 | v_70772;
assign v_70775 = v_70584 | v_70774;
assign v_70778 = v_70776 | v_70777;
assign v_70780 = v_70581 | v_70779;
assign v_70783 = v_70781 | v_70782;
assign v_70785 = v_70578 | v_70784;
assign v_70788 = v_70786 | v_70787;
assign v_70790 = v_70575 | v_70789;
assign v_70793 = v_70791 | v_70792;
assign v_70795 = v_70572 | v_70794;
assign v_70798 = v_70796 | v_70797;
assign v_70800 = v_70569 | v_70799;
assign v_70803 = v_70801 | v_70802;
assign v_70805 = v_70803 | v_70804;
assign v_70808 = v_70566 | v_70807;
assign v_70809 = ~v_4 | v_70808;
assign v_70814 = v_70811 | v_70813;
assign v_70820 = v_70817 | v_70819;
assign v_70828 = v_70825 | v_70827;
assign v_70836 = v_70833 | v_70835;
assign v_70844 = v_70841 | v_70843;
assign v_70852 = v_70849 | v_70851;
assign v_70860 = v_70857 | v_70859;
assign v_70868 = v_70865 | v_70867;
assign v_70876 = v_70873 | v_70875;
assign v_70884 = v_70881 | v_70883;
assign v_70892 = v_70889 | v_70891;
assign v_70900 = v_70897 | v_70899;
assign v_70908 = v_70905 | v_70907;
assign v_70916 = v_70913 | v_70915;
assign v_70924 = v_70921 | v_70923;
assign v_70932 = v_70929 | v_70931;
assign v_70940 = v_70937 | v_70939;
assign v_70948 = v_70945 | v_70947;
assign v_70956 = v_70953 | v_70955;
assign v_70964 = v_70961 | v_70963;
assign v_70972 = v_70969 | v_70971;
assign v_70980 = v_70977 | v_70979;
assign v_70988 = v_70985 | v_70987;
assign v_70996 = v_70993 | v_70995;
assign v_71004 = v_71001 | v_71003;
assign v_71012 = v_71009 | v_71011;
assign v_71020 = v_71017 | v_71019;
assign v_71028 = v_71025 | v_71027;
assign v_71036 = v_71033 | v_71035;
assign v_71044 = v_71041 | v_71043;
assign v_71052 = v_71049 | v_71051;
assign v_71060 = v_71057 | v_71059;
assign v_71068 = v_71065 | v_71067;
assign v_71076 = v_71073 | v_71075;
assign v_71084 = v_71081 | v_71083;
assign v_71092 = v_71089 | v_71091;
assign v_71100 = v_71097 | v_71099;
assign v_71108 = v_71105 | v_71107;
assign v_71116 = v_71113 | v_71115;
assign v_71124 = v_71121 | v_71123;
assign v_71132 = v_71129 | v_71131;
assign v_71140 = v_71137 | v_71139;
assign v_71148 = v_71145 | v_71147;
assign v_71156 = v_71153 | v_71155;
assign v_71164 = v_71161 | v_71163;
assign v_71172 = v_71169 | v_71171;
assign v_71180 = v_71177 | v_71179;
assign v_71188 = v_71185 | v_71187;
assign v_71196 = v_71193 | v_71195;
assign v_71204 = v_71201 | v_71203;
assign v_71212 = v_71209 | v_71211;
assign v_71220 = v_71217 | v_71219;
assign v_71228 = v_71225 | v_71227;
assign v_71236 = v_71233 | v_71235;
assign v_71244 = v_71241 | v_71243;
assign v_71252 = v_71249 | v_71251;
assign v_71260 = v_71257 | v_71259;
assign v_71268 = v_71265 | v_71267;
assign v_71276 = v_71273 | v_71275;
assign v_71284 = v_71281 | v_71283;
assign v_71292 = v_71289 | v_71291;
assign v_71300 = v_71297 | v_71299;
assign v_71308 = v_71305 | v_71307;
assign v_71316 = v_71313 | v_71315;
assign v_71324 = v_71321 | v_71323;
assign v_71332 = v_71329 | v_71331;
assign v_71340 = v_71337 | v_71339;
assign v_71348 = v_71345 | v_71347;
assign v_71356 = v_71353 | v_71355;
assign v_71364 = v_71361 | v_71363;
assign v_71372 = v_71369 | v_71371;
assign v_71380 = v_71377 | v_71379;
assign v_71388 = v_71385 | v_71387;
assign v_71396 = v_71393 | v_71395;
assign v_71404 = v_71401 | v_71403;
assign v_71412 = v_71409 | v_71411;
assign v_71420 = v_71417 | v_71419;
assign v_71428 = v_71425 | v_71427;
assign v_71436 = v_71433 | v_71435;
assign v_71444 = v_71441 | v_71443;
assign v_71452 = v_71449 | v_71451;
assign v_71460 = v_71457 | v_71459;
assign v_71468 = v_71465 | v_71467;
assign v_71476 = v_71473 | v_71475;
assign v_71484 = v_71481 | v_71483;
assign v_71492 = v_71489 | v_71491;
assign v_71500 = v_71497 | v_71499;
assign v_71508 = v_71505 | v_71507;
assign v_71516 = v_71513 | v_71515;
assign v_71524 = v_71521 | v_71523;
assign v_71532 = v_71529 | v_71531;
assign v_71540 = v_71537 | v_71539;
assign v_71548 = v_71545 | v_71547;
assign v_71556 = v_71553 | v_71555;
assign v_71564 = v_71561 | v_71563;
assign v_71572 = v_71569 | v_71571;
assign v_71580 = v_71577 | v_71579;
assign v_71588 = v_71585 | v_71587;
assign v_71596 = v_71593 | v_71595;
assign v_71604 = v_71601 | v_71603;
assign v_71612 = v_71609 | v_71611;
assign v_71620 = v_71617 | v_71619;
assign v_71628 = v_71625 | v_71627;
assign v_71636 = v_71633 | v_71635;
assign v_71644 = v_71641 | v_71643;
assign v_71652 = v_71649 | v_71651;
assign v_71660 = v_71657 | v_71659;
assign v_71668 = v_71665 | v_71667;
assign v_71676 = v_71673 | v_71675;
assign v_71684 = v_71681 | v_71683;
assign v_71692 = v_71689 | v_71691;
assign v_71700 = v_71697 | v_71699;
assign v_71708 = v_71705 | v_71707;
assign v_71716 = v_71713 | v_71715;
assign v_71724 = v_71721 | v_71723;
assign v_71732 = v_71729 | v_71731;
assign v_71740 = v_71737 | v_71739;
assign v_71748 = v_71745 | v_71747;
assign v_71756 = v_71753 | v_71755;
assign v_71764 = v_71761 | v_71763;
assign v_71772 = v_71769 | v_71771;
assign v_71780 = v_71777 | v_71779;
assign v_71788 = v_71785 | v_71787;
assign v_71796 = v_71793 | v_71795;
assign v_71804 = v_71801 | v_71803;
assign v_71812 = v_71809 | v_71811;
assign v_71820 = v_71817 | v_71819;
assign v_71828 = v_71825 | v_71827;
assign v_71836 = v_71833 | v_71835;
assign v_71844 = v_71841 | v_71843;
assign v_71852 = v_71849 | v_71851;
assign v_71860 = v_71857 | v_71859;
assign v_71868 = v_71865 | v_71867;
assign v_71876 = v_71873 | v_71875;
assign v_71884 = v_71881 | v_71883;
assign v_71892 = v_71889 | v_71891;
assign v_71900 = v_71897 | v_71899;
assign v_71908 = v_71905 | v_71907;
assign v_71916 = v_71913 | v_71915;
assign v_71924 = v_71921 | v_71923;
assign v_71932 = v_71929 | v_71931;
assign v_71940 = v_71937 | v_71939;
assign v_71948 = v_71945 | v_71947;
assign v_71956 = v_71953 | v_71955;
assign v_71964 = v_71961 | v_71963;
assign v_71972 = v_71969 | v_71971;
assign v_71980 = v_71977 | v_71979;
assign v_71988 = v_71985 | v_71987;
assign v_71996 = v_71993 | v_71995;
assign v_72004 = v_72001 | v_72003;
assign v_72012 = v_72009 | v_72011;
assign v_72020 = v_72017 | v_72019;
assign v_72028 = v_72025 | v_72027;
assign v_72036 = v_72033 | v_72035;
assign v_72044 = v_72041 | v_72043;
assign v_72052 = v_72049 | v_72051;
assign v_72060 = v_72057 | v_72059;
assign v_72068 = v_72065 | v_72067;
assign v_72076 = v_72073 | v_72075;
assign v_72084 = v_72081 | v_72083;
assign v_72092 = v_72089 | v_72091;
assign v_72100 = v_72097 | v_72099;
assign v_72108 = v_72105 | v_72107;
assign v_72116 = v_72113 | v_72115;
assign v_72124 = v_72121 | v_72123;
assign v_72132 = v_72129 | v_72131;
assign v_72140 = v_72137 | v_72139;
assign v_72148 = v_72145 | v_72147;
assign v_72156 = v_72153 | v_72155;
assign v_72164 = v_72161 | v_72163;
assign v_72172 = v_72169 | v_72171;
assign v_72180 = v_72177 | v_72179;
assign v_72188 = v_72185 | v_72187;
assign v_72196 = v_72193 | v_72195;
assign v_72204 = v_72201 | v_72203;
assign v_72212 = v_72209 | v_72211;
assign v_72220 = v_72217 | v_72219;
assign v_72228 = v_72225 | v_72227;
assign v_72236 = v_72233 | v_72235;
assign v_72244 = v_72241 | v_72243;
assign v_72252 = v_72249 | v_72251;
assign v_72260 = v_72257 | v_72259;
assign v_72268 = v_72265 | v_72267;
assign v_72276 = v_72273 | v_72275;
assign v_72284 = v_72281 | v_72283;
assign v_72292 = v_72289 | v_72291;
assign v_72300 = v_72297 | v_72299;
assign v_72308 = v_72305 | v_72307;
assign v_72316 = v_72313 | v_72315;
assign v_72324 = v_72321 | v_72323;
assign v_72332 = v_72329 | v_72331;
assign v_72340 = v_72337 | v_72339;
assign v_72348 = v_72345 | v_72347;
assign v_72356 = v_72353 | v_72355;
assign v_72364 = v_72361 | v_72363;
assign v_72372 = v_72369 | v_72371;
assign v_72380 = v_72377 | v_72379;
assign v_72388 = v_72385 | v_72387;
assign v_72396 = v_72393 | v_72395;
assign v_72404 = v_72401 | v_72403;
assign v_72412 = v_72409 | v_72411;
assign v_72420 = v_72417 | v_72419;
assign v_72428 = v_72425 | v_72427;
assign v_72436 = v_72433 | v_72435;
assign v_72444 = v_72441 | v_72443;
assign v_72452 = v_72449 | v_72451;
assign v_72460 = v_72457 | v_72459;
assign v_72468 = v_72465 | v_72467;
assign v_72476 = v_72473 | v_72475;
assign v_72484 = v_72481 | v_72483;
assign v_72492 = v_72489 | v_72491;
assign v_72500 = v_72497 | v_72499;
assign v_72508 = v_72505 | v_72507;
assign v_72516 = v_72513 | v_72515;
assign v_72524 = v_72521 | v_72523;
assign v_72532 = v_72529 | v_72531;
assign v_72540 = v_72537 | v_72539;
assign v_72548 = v_72545 | v_72547;
assign v_72556 = v_72553 | v_72555;
assign v_72564 = v_72561 | v_72563;
assign v_72572 = v_72569 | v_72571;
assign v_72580 = v_72577 | v_72579;
assign v_72588 = v_72585 | v_72587;
assign v_72596 = v_72593 | v_72595;
assign v_72604 = v_72601 | v_72603;
assign v_72612 = v_72609 | v_72611;
assign v_72620 = v_72617 | v_72619;
assign v_72628 = v_72625 | v_72627;
assign v_72636 = v_72633 | v_72635;
assign v_72644 = v_72641 | v_72643;
assign v_72652 = v_72649 | v_72651;
assign v_72660 = v_72657 | v_72659;
assign v_72668 = v_72665 | v_72667;
assign v_72676 = v_72673 | v_72675;
assign v_72684 = v_72681 | v_72683;
assign v_72692 = v_72689 | v_72691;
assign v_72700 = v_72697 | v_72699;
assign v_72708 = v_72705 | v_72707;
assign v_72716 = v_72713 | v_72715;
assign v_72724 = v_72721 | v_72723;
assign v_72732 = v_72729 | v_72731;
assign v_72740 = v_72737 | v_72739;
assign v_72748 = v_72745 | v_72747;
assign v_72756 = v_72753 | v_72755;
assign v_72764 = v_72761 | v_72763;
assign v_72772 = v_72769 | v_72771;
assign v_72780 = v_72777 | v_72779;
assign v_72788 = v_72785 | v_72787;
assign v_72796 = v_72793 | v_72795;
assign v_72804 = v_72801 | v_72803;
assign v_72812 = v_72809 | v_72811;
assign v_72820 = v_72817 | v_72819;
assign v_72828 = v_72825 | v_72827;
assign v_72836 = v_72833 | v_72835;
assign v_72844 = v_72841 | v_72843;
assign v_72852 = v_72849 | v_72851;
assign v_72860 = v_72857 | v_72859;
assign v_72868 = v_72865 | v_72867;
assign v_72876 = v_72873 | v_72875;
assign v_72884 = v_72881 | v_72883;
assign v_72892 = v_72889 | v_72891;
assign v_72900 = v_72897 | v_72899;
assign v_72908 = v_72905 | v_72907;
assign v_72916 = v_72913 | v_72915;
assign v_72924 = v_72921 | v_72923;
assign v_72932 = v_72929 | v_72931;
assign v_72940 = v_72937 | v_72939;
assign v_72948 = v_72945 | v_72947;
assign v_72956 = v_72953 | v_72955;
assign v_72964 = v_72961 | v_72963;
assign v_72972 = v_72969 | v_72971;
assign v_72980 = v_72977 | v_72979;
assign v_72988 = v_72985 | v_72987;
assign v_72996 = v_72993 | v_72995;
assign v_73004 = v_73001 | v_73003;
assign v_73012 = v_73009 | v_73011;
assign v_73020 = v_73017 | v_73019;
assign v_73028 = v_73025 | v_73027;
assign v_73036 = v_73033 | v_73035;
assign v_73044 = v_73041 | v_73043;
assign v_73052 = v_73049 | v_73051;
assign v_73060 = v_73057 | v_73059;
assign v_73068 = v_73065 | v_73067;
assign v_73076 = v_73073 | v_73075;
assign v_73084 = v_73081 | v_73083;
assign v_73092 = v_73089 | v_73091;
assign v_73100 = v_73097 | v_73099;
assign v_73108 = v_73105 | v_73107;
assign v_73116 = v_73113 | v_73115;
assign v_73119 = v_4 | v_73118;
assign x_1 = v_3 | v_73122;
assign o_1 = x_1;
endmodule
