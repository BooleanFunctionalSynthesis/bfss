// Generated using findDep.cpp 
module small-swap2-fixpoint-8 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_578, v_579, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_660, v_661, v_662, v_663, v_664, v_665, v_666, v_667, v_668, v_669, v_670, v_671, v_672, v_673, v_674, v_675, v_676, v_677, v_678, v_679, v_680, v_681, v_682, v_683, v_684, v_685, v_686, v_687, v_688, v_689, v_690, v_691, v_692, v_693, v_694, v_695, v_696, v_697, v_698, v_699, v_700, v_701, v_702, v_703, v_704, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_771, v_772, v_773, v_774, v_775, v_776, v_777, v_778, v_779, v_780, v_781, v_782, v_783, v_784, v_785, v_786, v_787, v_788, v_789, v_790, v_791, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_886, v_887, v_888, v_889, v_890, v_891, v_892, v_893, v_894, v_895, v_896, v_897, v_898, v_899, v_900, v_901, v_902, v_903, v_904, v_905, v_906, v_907, v_908, v_909, v_910, v_911, v_912, v_913, v_914, v_915, v_916, v_917, v_918, v_919, v_920, v_921, v_922, v_923, v_924, v_925, v_926, v_927, v_928, v_929, v_930, v_931, v_932, v_933, v_934, v_935, v_936, v_937, v_938, v_939, v_940, v_941, v_942, v_943, v_944, v_945, v_946, v_947, v_948, v_949, v_950, v_951, v_952, v_953, v_954, v_955, v_956, v_957, v_958, v_959, v_960, v_961, v_962, v_963, v_964, v_965, v_966, v_967, v_968, v_969, v_970, v_971, v_972, v_973, v_974, v_975, v_976, v_977, v_978, v_979, v_980, v_981, v_982, v_983, v_984, v_985, v_986, v_987, v_988, v_989, v_990, v_991, v_992, v_993, v_994, v_995, v_996, v_997, v_998, v_999, v_1000, v_1001, v_1002, v_1003, v_1004, v_1005, v_1006, v_1007, v_1008, v_1009, v_1010, v_1011, v_1012, v_1013, v_1014, v_1015, v_1016, v_1017, v_1018, v_1019, v_1020, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_578;
input v_579;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_660;
input v_661;
input v_662;
input v_663;
input v_664;
input v_665;
input v_666;
input v_667;
input v_668;
input v_669;
input v_670;
input v_671;
input v_672;
input v_673;
input v_674;
input v_675;
input v_676;
input v_677;
input v_678;
input v_679;
input v_680;
input v_681;
input v_682;
input v_683;
input v_684;
input v_685;
input v_686;
input v_687;
input v_688;
input v_689;
input v_690;
input v_691;
input v_692;
input v_693;
input v_694;
input v_695;
input v_696;
input v_697;
input v_698;
input v_699;
input v_700;
input v_701;
input v_702;
input v_703;
input v_704;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_771;
input v_772;
input v_773;
input v_774;
input v_775;
input v_776;
input v_777;
input v_778;
input v_779;
input v_780;
input v_781;
input v_782;
input v_783;
input v_784;
input v_785;
input v_786;
input v_787;
input v_788;
input v_789;
input v_790;
input v_791;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_886;
input v_887;
input v_888;
input v_889;
input v_890;
input v_891;
input v_892;
input v_893;
input v_894;
input v_895;
input v_896;
input v_897;
input v_898;
input v_899;
input v_900;
input v_901;
input v_902;
input v_903;
input v_904;
input v_905;
input v_906;
input v_907;
input v_908;
input v_909;
input v_910;
input v_911;
input v_912;
input v_913;
input v_914;
input v_915;
input v_916;
input v_917;
input v_918;
input v_919;
input v_920;
input v_921;
input v_922;
input v_923;
input v_924;
input v_925;
input v_926;
input v_927;
input v_928;
input v_929;
input v_930;
input v_931;
input v_932;
input v_933;
input v_934;
input v_935;
input v_936;
input v_937;
input v_938;
input v_939;
input v_940;
input v_941;
input v_942;
input v_943;
input v_944;
input v_945;
input v_946;
input v_947;
input v_948;
input v_949;
input v_950;
input v_951;
input v_952;
input v_953;
input v_954;
input v_955;
input v_956;
input v_957;
input v_958;
input v_959;
input v_960;
input v_961;
input v_962;
input v_963;
input v_964;
input v_965;
input v_966;
input v_967;
input v_968;
input v_969;
input v_970;
input v_971;
input v_972;
input v_973;
input v_974;
input v_975;
input v_976;
input v_977;
input v_978;
input v_979;
input v_980;
input v_981;
input v_982;
input v_983;
input v_984;
input v_985;
input v_986;
input v_987;
input v_988;
input v_989;
input v_990;
input v_991;
input v_992;
input v_993;
input v_994;
input v_995;
input v_996;
input v_997;
input v_998;
input v_999;
input v_1000;
input v_1001;
input v_1002;
input v_1003;
input v_1004;
input v_1005;
input v_1006;
input v_1007;
input v_1008;
input v_1009;
input v_1010;
input v_1011;
input v_1012;
input v_1013;
input v_1014;
input v_1015;
input v_1016;
input v_1017;
input v_1018;
input v_1019;
input v_1020;
output o_1;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2115;
wire v_2116;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2120;
wire v_2121;
wire v_2122;
wire v_2123;
wire v_2124;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2132;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2136;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2157;
wire v_2158;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2169;
wire v_2170;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2181;
wire v_2182;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2218;
wire v_2219;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2226;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2265;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2362;
wire v_2363;
wire v_2364;
wire v_2365;
wire v_2366;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2371;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2392;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2396;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2640;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2648;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2664;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2680;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2744;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2755;
wire v_2756;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2764;
wire v_2765;
wire v_2766;
wire v_2767;
wire v_2768;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2786;
wire v_2787;
wire v_2788;
wire v_2789;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2795;
wire v_2796;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2804;
wire v_2805;
wire v_2806;
wire v_2807;
wire v_2808;
wire v_2809;
wire v_2810;
wire x_1;
assign v_1021 = v_2505 & v_2506 & v_2507 & v_2508;
assign v_1022 = v_2509 & v_2510 & v_2511 & v_2512;
assign v_1023 = v_2513 & v_2514 & v_2515 & v_2516;
assign v_1024 = v_1021 & v_1022 & v_1023;
assign v_1045 = v_2517 & v_2518 & v_2519 & v_2520;
assign v_1066 = v_2521 & v_2522 & v_2523 & v_2524;
assign v_1087 = v_2525 & v_2526 & v_2527 & v_2528;
assign v_1088 = v_1045 & v_1066 & v_1087;
assign v_1109 = v_2529 & v_2530 & v_2531 & v_2532;
assign v_1130 = v_2533 & v_2534 & v_2535 & v_2536;
assign v_1151 = v_2537 & v_2538 & v_2539 & v_2540;
assign v_1152 = v_1109 & v_1130 & v_1151;
assign v_1173 = v_2541 & v_2542 & v_2543 & v_2544;
assign v_1194 = v_2545 & v_2546 & v_2547 & v_2548;
assign v_1215 = v_2549 & v_2550 & v_2551 & v_2552;
assign v_1216 = v_1173 & v_1194 & v_1215;
assign v_1237 = v_2553 & v_2554 & v_2555 & v_2556;
assign v_1258 = v_2557 & v_2558 & v_2559 & v_2560;
assign v_1279 = v_2561 & v_2562 & v_2563 & v_2564;
assign v_1280 = v_1237 & v_1258 & v_1279;
assign v_1301 = v_2565 & v_2566 & v_2567 & v_2568;
assign v_1322 = v_2569 & v_2570 & v_2571 & v_2572;
assign v_1343 = v_2573 & v_2574 & v_2575 & v_2576;
assign v_1344 = v_1301 & v_1322 & v_1343;
assign v_1365 = v_2577 & v_2578 & v_2579 & v_2580;
assign v_1386 = v_2581 & v_2582 & v_2583 & v_2584;
assign v_1407 = v_2585 & v_2586 & v_2587 & v_2588;
assign v_1408 = v_1365 & v_1386 & v_1407;
assign v_1429 = v_2589 & v_2590 & v_2591 & v_2592;
assign v_1450 = v_2593 & v_2594 & v_2595 & v_2596;
assign v_1471 = v_2597 & v_2598 & v_2599 & v_2600;
assign v_1472 = v_1429 & v_1450 & v_1471;
assign v_1493 = v_2601 & v_2602 & v_2603 & v_2604;
assign v_1514 = v_2605 & v_2606 & v_2607 & v_2608;
assign v_1535 = v_2609 & v_2610 & v_2611 & v_2612;
assign v_1536 = v_1493 & v_1514 & v_1535;
assign v_1537 = v_2613 & v_2614;
assign v_1538 = v_2615 & v_2616 & v_2617 & v_2618;
assign v_1539 = v_2619 & v_2620 & v_2621 & v_2622;
assign v_1540 = v_2623 & v_2624 & v_2625 & v_2626;
assign v_1541 = v_1538 & v_1539 & v_1540;
assign v_1562 = v_2627 & v_2628 & v_2629 & v_2630;
assign v_1583 = v_2631 & v_2632 & v_2633 & v_2634;
assign v_1604 = v_2635 & v_2636 & v_2637 & v_2638;
assign v_1605 = v_1562 & v_1583 & v_1604;
assign v_1626 = v_2639 & v_2640 & v_2641 & v_2642;
assign v_1647 = v_2643 & v_2644 & v_2645 & v_2646;
assign v_1668 = v_2647 & v_2648 & v_2649 & v_2650;
assign v_1669 = v_1626 & v_1647 & v_1668;
assign v_1690 = v_2651 & v_2652 & v_2653 & v_2654;
assign v_1711 = v_2655 & v_2656 & v_2657 & v_2658;
assign v_1732 = v_2659 & v_2660 & v_2661 & v_2662;
assign v_1733 = v_1690 & v_1711 & v_1732;
assign v_1754 = v_2663 & v_2664 & v_2665 & v_2666;
assign v_1775 = v_2667 & v_2668 & v_2669 & v_2670;
assign v_1796 = v_2671 & v_2672 & v_2673 & v_2674;
assign v_1797 = v_1754 & v_1775 & v_1796;
assign v_1818 = v_2675 & v_2676 & v_2677 & v_2678;
assign v_1839 = v_2679 & v_2680 & v_2681 & v_2682;
assign v_1860 = v_2683 & v_2684 & v_2685 & v_2686;
assign v_1861 = v_1818 & v_1839 & v_1860;
assign v_1882 = v_2687 & v_2688 & v_2689 & v_2690;
assign v_1903 = v_2691 & v_2692 & v_2693 & v_2694;
assign v_1924 = v_2695 & v_2696 & v_2697 & v_2698;
assign v_1925 = v_1882 & v_1903 & v_1924;
assign v_1946 = v_2699 & v_2700 & v_2701 & v_2702;
assign v_1967 = v_2703 & v_2704 & v_2705 & v_2706;
assign v_1988 = v_2707 & v_2708 & v_2709 & v_2710;
assign v_1989 = v_1946 & v_1967 & v_1988;
assign v_1990 = v_2711 & v_2712;
assign v_2011 = v_2713 & v_2714 & v_2715 & v_2716;
assign v_2032 = v_2717 & v_2718 & v_2719 & v_2720;
assign v_2053 = v_2721 & v_2722 & v_2723 & v_2724;
assign v_2054 = v_2011 & v_2032 & v_2053;
assign v_2075 = v_2725 & v_2726 & v_2727 & v_2728;
assign v_2096 = v_2729 & v_2730 & v_2731 & v_2732;
assign v_2117 = v_2733 & v_2734 & v_2735 & v_2736;
assign v_2118 = v_2075 & v_2096 & v_2117;
assign v_2139 = v_2737 & v_2738 & v_2739 & v_2740;
assign v_2160 = v_2741 & v_2742 & v_2743 & v_2744;
assign v_2181 = v_2745 & v_2746 & v_2747 & v_2748;
assign v_2182 = v_2139 & v_2160 & v_2181;
assign v_2203 = v_2749 & v_2750 & v_2751 & v_2752;
assign v_2224 = v_2753 & v_2754 & v_2755 & v_2756;
assign v_2245 = v_2757 & v_2758 & v_2759 & v_2760;
assign v_2246 = v_2203 & v_2224 & v_2245;
assign v_2267 = v_2761 & v_2762 & v_2763 & v_2764;
assign v_2288 = v_2765 & v_2766 & v_2767 & v_2768;
assign v_2309 = v_2769 & v_2770 & v_2771 & v_2772;
assign v_2310 = v_2267 & v_2288 & v_2309;
assign v_2331 = v_2773 & v_2774 & v_2775 & v_2776;
assign v_2352 = v_2777 & v_2778 & v_2779 & v_2780;
assign v_2373 = v_2781 & v_2782 & v_2783 & v_2784;
assign v_2374 = v_2331 & v_2352 & v_2373;
assign v_2395 = v_2785 & v_2786 & v_2787 & v_2788;
assign v_2416 = v_2789 & v_2790 & v_2791 & v_2792;
assign v_2437 = v_2793 & v_2794 & v_2795 & v_2796;
assign v_2438 = v_2395 & v_2416 & v_2437;
assign v_2459 = v_2797 & v_2798 & v_2799 & v_2800;
assign v_2480 = v_2801 & v_2802 & v_2803 & v_2804;
assign v_2501 = v_2805 & v_2806 & v_2807 & v_2808;
assign v_2502 = v_2459 & v_2480 & v_2501;
assign v_2504 = v_1990 & v_2503;
assign v_2505 = ~v_2 & ~v_3 & ~v_4 & ~v_5 & ~v_6;
assign v_2506 = ~v_7 & ~v_8 & ~v_9 & ~v_10 & ~v_11;
assign v_2507 = ~v_12 & ~v_13 & ~v_14 & ~v_15 & ~v_16;
assign v_2508 = ~v_17 & ~v_18 & ~v_19 & ~v_20 & v_1;
assign v_2509 = ~v_22 & ~v_24 & ~v_25 & ~v_26 & ~v_27;
assign v_2510 = ~v_28 & ~v_29 & ~v_30 & ~v_31 & ~v_32;
assign v_2511 = ~v_33 & ~v_34 & ~v_35 & ~v_36 & ~v_37;
assign v_2512 = ~v_38 & ~v_39 & ~v_40 & v_21 & v_23;
assign v_2513 = ~v_44 & ~v_45 & ~v_46 & ~v_47 & ~v_48;
assign v_2514 = ~v_49 & ~v_50 & ~v_51 & ~v_52 & ~v_53;
assign v_2515 = ~v_54 & ~v_55 & ~v_56 & ~v_57 & ~v_58;
assign v_2516 = ~v_59 & ~v_60 & v_41 & v_42 & v_43;
assign v_2517 = ~v_1025 & ~v_1026 & ~v_1027 & ~v_1028 & ~v_1029;
assign v_2518 = ~v_1030 & ~v_1031 & ~v_1032 & ~v_1033 & ~v_1034;
assign v_2519 = ~v_1035 & ~v_1036 & ~v_1037 & ~v_1038 & ~v_1039;
assign v_2520 = ~v_1040 & ~v_1041 & ~v_1042 & ~v_1043 & ~v_1044;
assign v_2521 = ~v_1046 & ~v_1047 & ~v_1048 & ~v_1049 & ~v_1050;
assign v_2522 = ~v_1051 & ~v_1052 & ~v_1053 & ~v_1054 & ~v_1055;
assign v_2523 = ~v_1056 & ~v_1057 & ~v_1058 & ~v_1059 & ~v_1060;
assign v_2524 = ~v_1061 & ~v_1062 & ~v_1063 & ~v_1064 & ~v_1065;
assign v_2525 = ~v_1067 & ~v_1068 & ~v_1069 & ~v_1070 & ~v_1071;
assign v_2526 = ~v_1072 & ~v_1073 & ~v_1074 & ~v_1075 & ~v_1076;
assign v_2527 = ~v_1077 & ~v_1078 & ~v_1079 & ~v_1080 & ~v_1081;
assign v_2528 = ~v_1082 & ~v_1083 & ~v_1084 & ~v_1085 & ~v_1086;
assign v_2529 = ~v_1089 & ~v_1090 & ~v_1091 & ~v_1092 & ~v_1093;
assign v_2530 = ~v_1094 & ~v_1095 & ~v_1096 & ~v_1097 & ~v_1098;
assign v_2531 = ~v_1099 & ~v_1100 & ~v_1101 & ~v_1102 & ~v_1103;
assign v_2532 = ~v_1104 & ~v_1105 & ~v_1106 & ~v_1107 & ~v_1108;
assign v_2533 = ~v_1110 & ~v_1111 & ~v_1112 & ~v_1113 & ~v_1114;
assign v_2534 = ~v_1115 & ~v_1116 & ~v_1117 & ~v_1118 & ~v_1119;
assign v_2535 = ~v_1120 & ~v_1121 & ~v_1122 & ~v_1123 & ~v_1124;
assign v_2536 = ~v_1125 & ~v_1126 & ~v_1127 & ~v_1128 & ~v_1129;
assign v_2537 = ~v_1131 & ~v_1132 & ~v_1133 & ~v_1134 & ~v_1135;
assign v_2538 = ~v_1136 & ~v_1137 & ~v_1138 & ~v_1139 & ~v_1140;
assign v_2539 = ~v_1141 & ~v_1142 & ~v_1143 & ~v_1144 & ~v_1145;
assign v_2540 = ~v_1146 & ~v_1147 & ~v_1148 & ~v_1149 & ~v_1150;
assign v_2541 = ~v_1153 & ~v_1154 & ~v_1155 & ~v_1156 & ~v_1157;
assign v_2542 = ~v_1158 & ~v_1159 & ~v_1160 & ~v_1161 & ~v_1162;
assign v_2543 = ~v_1163 & ~v_1164 & ~v_1165 & ~v_1166 & ~v_1167;
assign v_2544 = ~v_1168 & ~v_1169 & ~v_1170 & ~v_1171 & ~v_1172;
assign v_2545 = ~v_1174 & ~v_1175 & ~v_1176 & ~v_1177 & ~v_1178;
assign v_2546 = ~v_1179 & ~v_1180 & ~v_1181 & ~v_1182 & ~v_1183;
assign v_2547 = ~v_1184 & ~v_1185 & ~v_1186 & ~v_1187 & ~v_1188;
assign v_2548 = ~v_1189 & ~v_1190 & ~v_1191 & ~v_1192 & ~v_1193;
assign v_2549 = ~v_1195 & ~v_1196 & ~v_1197 & ~v_1198 & ~v_1199;
assign v_2550 = ~v_1200 & ~v_1201 & ~v_1202 & ~v_1203 & ~v_1204;
assign v_2551 = ~v_1205 & ~v_1206 & ~v_1207 & ~v_1208 & ~v_1209;
assign v_2552 = ~v_1210 & ~v_1211 & ~v_1212 & ~v_1213 & ~v_1214;
assign v_2553 = ~v_1217 & ~v_1218 & ~v_1219 & ~v_1220 & ~v_1221;
assign v_2554 = ~v_1222 & ~v_1223 & ~v_1224 & ~v_1225 & ~v_1226;
assign v_2555 = ~v_1227 & ~v_1228 & ~v_1229 & ~v_1230 & ~v_1231;
assign v_2556 = ~v_1232 & ~v_1233 & ~v_1234 & ~v_1235 & ~v_1236;
assign v_2557 = ~v_1238 & ~v_1239 & ~v_1240 & ~v_1241 & ~v_1242;
assign v_2558 = ~v_1243 & ~v_1244 & ~v_1245 & ~v_1246 & ~v_1247;
assign v_2559 = ~v_1248 & ~v_1249 & ~v_1250 & ~v_1251 & ~v_1252;
assign v_2560 = ~v_1253 & ~v_1254 & ~v_1255 & ~v_1256 & ~v_1257;
assign v_2561 = ~v_1259 & ~v_1260 & ~v_1261 & ~v_1262 & ~v_1263;
assign v_2562 = ~v_1264 & ~v_1265 & ~v_1266 & ~v_1267 & ~v_1268;
assign v_2563 = ~v_1269 & ~v_1270 & ~v_1271 & ~v_1272 & ~v_1273;
assign v_2564 = ~v_1274 & ~v_1275 & ~v_1276 & ~v_1277 & ~v_1278;
assign v_2565 = ~v_1281 & ~v_1282 & ~v_1283 & ~v_1284 & ~v_1285;
assign v_2566 = ~v_1286 & ~v_1287 & ~v_1288 & ~v_1289 & ~v_1290;
assign v_2567 = ~v_1291 & ~v_1292 & ~v_1293 & ~v_1294 & ~v_1295;
assign v_2568 = ~v_1296 & ~v_1297 & ~v_1298 & ~v_1299 & ~v_1300;
assign v_2569 = ~v_1302 & ~v_1303 & ~v_1304 & ~v_1305 & ~v_1306;
assign v_2570 = ~v_1307 & ~v_1308 & ~v_1309 & ~v_1310 & ~v_1311;
assign v_2571 = ~v_1312 & ~v_1313 & ~v_1314 & ~v_1315 & ~v_1316;
assign v_2572 = ~v_1317 & ~v_1318 & ~v_1319 & ~v_1320 & ~v_1321;
assign v_2573 = ~v_1323 & ~v_1324 & ~v_1325 & ~v_1326 & ~v_1327;
assign v_2574 = ~v_1328 & ~v_1329 & ~v_1330 & ~v_1331 & ~v_1332;
assign v_2575 = ~v_1333 & ~v_1334 & ~v_1335 & ~v_1336 & ~v_1337;
assign v_2576 = ~v_1338 & ~v_1339 & ~v_1340 & ~v_1341 & ~v_1342;
assign v_2577 = ~v_1345 & ~v_1346 & ~v_1347 & ~v_1348 & ~v_1349;
assign v_2578 = ~v_1350 & ~v_1351 & ~v_1352 & ~v_1353 & ~v_1354;
assign v_2579 = ~v_1355 & ~v_1356 & ~v_1357 & ~v_1358 & ~v_1359;
assign v_2580 = ~v_1360 & ~v_1361 & ~v_1362 & ~v_1363 & ~v_1364;
assign v_2581 = ~v_1366 & ~v_1367 & ~v_1368 & ~v_1369 & ~v_1370;
assign v_2582 = ~v_1371 & ~v_1372 & ~v_1373 & ~v_1374 & ~v_1375;
assign v_2583 = ~v_1376 & ~v_1377 & ~v_1378 & ~v_1379 & ~v_1380;
assign v_2584 = ~v_1381 & ~v_1382 & ~v_1383 & ~v_1384 & ~v_1385;
assign v_2585 = ~v_1387 & ~v_1388 & ~v_1389 & ~v_1390 & ~v_1391;
assign v_2586 = ~v_1392 & ~v_1393 & ~v_1394 & ~v_1395 & ~v_1396;
assign v_2587 = ~v_1397 & ~v_1398 & ~v_1399 & ~v_1400 & ~v_1401;
assign v_2588 = ~v_1402 & ~v_1403 & ~v_1404 & ~v_1405 & ~v_1406;
assign v_2589 = ~v_1409 & ~v_1410 & ~v_1411 & ~v_1412 & ~v_1413;
assign v_2590 = ~v_1414 & ~v_1415 & ~v_1416 & ~v_1417 & ~v_1418;
assign v_2591 = ~v_1419 & ~v_1420 & ~v_1421 & ~v_1422 & ~v_1423;
assign v_2592 = ~v_1424 & ~v_1425 & ~v_1426 & ~v_1427 & ~v_1428;
assign v_2593 = ~v_1430 & ~v_1431 & ~v_1432 & ~v_1433 & ~v_1434;
assign v_2594 = ~v_1435 & ~v_1436 & ~v_1437 & ~v_1438 & ~v_1439;
assign v_2595 = ~v_1440 & ~v_1441 & ~v_1442 & ~v_1443 & ~v_1444;
assign v_2596 = ~v_1445 & ~v_1446 & ~v_1447 & ~v_1448 & ~v_1449;
assign v_2597 = ~v_1451 & ~v_1452 & ~v_1453 & ~v_1454 & ~v_1455;
assign v_2598 = ~v_1456 & ~v_1457 & ~v_1458 & ~v_1459 & ~v_1460;
assign v_2599 = ~v_1461 & ~v_1462 & ~v_1463 & ~v_1464 & ~v_1465;
assign v_2600 = ~v_1466 & ~v_1467 & ~v_1468 & ~v_1469 & ~v_1470;
assign v_2601 = ~v_1473 & ~v_1474 & ~v_1475 & ~v_1476 & ~v_1477;
assign v_2602 = ~v_1478 & ~v_1479 & ~v_1480 & ~v_1481 & ~v_1482;
assign v_2603 = ~v_1483 & ~v_1484 & ~v_1485 & ~v_1486 & ~v_1487;
assign v_2604 = ~v_1488 & ~v_1489 & ~v_1490 & ~v_1491 & ~v_1492;
assign v_2605 = ~v_1494 & ~v_1495 & ~v_1496 & ~v_1497 & ~v_1498;
assign v_2606 = ~v_1499 & ~v_1500 & ~v_1501 & ~v_1502 & ~v_1503;
assign v_2607 = ~v_1504 & ~v_1505 & ~v_1506 & ~v_1507 & ~v_1508;
assign v_2608 = ~v_1509 & ~v_1510 & ~v_1511 & ~v_1512 & ~v_1513;
assign v_2609 = ~v_1515 & ~v_1516 & ~v_1517 & ~v_1518 & ~v_1519;
assign v_2610 = ~v_1520 & ~v_1521 & ~v_1522 & ~v_1523 & ~v_1524;
assign v_2611 = ~v_1525 & ~v_1526 & ~v_1527 & ~v_1528 & ~v_1529;
assign v_2612 = ~v_1530 & ~v_1531 & ~v_1532 & ~v_1533 & ~v_1534;
assign v_2613 = v_1024 & v_1088 & v_1152 & v_1216 & v_1280;
assign v_2614 = v_1344 & v_1408 & v_1472 & v_1536;
assign v_2615 = ~v_542 & ~v_543 & ~v_544 & ~v_545 & ~v_546;
assign v_2616 = ~v_547 & ~v_548 & ~v_549 & ~v_550 & ~v_551;
assign v_2617 = ~v_552 & ~v_553 & ~v_554 & ~v_555 & ~v_556;
assign v_2618 = ~v_557 & ~v_558 & ~v_559 & ~v_560 & v_541;
assign v_2619 = ~v_562 & ~v_564 & ~v_565 & ~v_566 & ~v_567;
assign v_2620 = ~v_568 & ~v_569 & ~v_570 & ~v_571 & ~v_572;
assign v_2621 = ~v_573 & ~v_574 & ~v_575 & ~v_576 & ~v_577;
assign v_2622 = ~v_578 & ~v_579 & ~v_580 & v_561 & v_563;
assign v_2623 = ~v_584 & ~v_585 & ~v_586 & ~v_587 & ~v_588;
assign v_2624 = ~v_589 & ~v_590 & ~v_591 & ~v_592 & ~v_593;
assign v_2625 = ~v_594 & ~v_595 & ~v_596 & ~v_597 & ~v_598;
assign v_2626 = ~v_599 & ~v_600 & v_581 & v_582 & v_583;
assign v_2627 = ~v_1542 & ~v_1543 & ~v_1544 & ~v_1545 & ~v_1546;
assign v_2628 = ~v_1547 & ~v_1548 & ~v_1549 & ~v_1550 & ~v_1551;
assign v_2629 = ~v_1552 & ~v_1553 & ~v_1554 & ~v_1555 & ~v_1556;
assign v_2630 = ~v_1557 & ~v_1558 & ~v_1559 & ~v_1560 & ~v_1561;
assign v_2631 = ~v_1563 & ~v_1564 & ~v_1565 & ~v_1566 & ~v_1567;
assign v_2632 = ~v_1568 & ~v_1569 & ~v_1570 & ~v_1571 & ~v_1572;
assign v_2633 = ~v_1573 & ~v_1574 & ~v_1575 & ~v_1576 & ~v_1577;
assign v_2634 = ~v_1578 & ~v_1579 & ~v_1580 & ~v_1581 & ~v_1582;
assign v_2635 = ~v_1584 & ~v_1585 & ~v_1586 & ~v_1587 & ~v_1588;
assign v_2636 = ~v_1589 & ~v_1590 & ~v_1591 & ~v_1592 & ~v_1593;
assign v_2637 = ~v_1594 & ~v_1595 & ~v_1596 & ~v_1597 & ~v_1598;
assign v_2638 = ~v_1599 & ~v_1600 & ~v_1601 & ~v_1602 & ~v_1603;
assign v_2639 = ~v_1606 & ~v_1607 & ~v_1608 & ~v_1609 & ~v_1610;
assign v_2640 = ~v_1611 & ~v_1612 & ~v_1613 & ~v_1614 & ~v_1615;
assign v_2641 = ~v_1616 & ~v_1617 & ~v_1618 & ~v_1619 & ~v_1620;
assign v_2642 = ~v_1621 & ~v_1622 & ~v_1623 & ~v_1624 & ~v_1625;
assign v_2643 = ~v_1627 & ~v_1628 & ~v_1629 & ~v_1630 & ~v_1631;
assign v_2644 = ~v_1632 & ~v_1633 & ~v_1634 & ~v_1635 & ~v_1636;
assign v_2645 = ~v_1637 & ~v_1638 & ~v_1639 & ~v_1640 & ~v_1641;
assign v_2646 = ~v_1642 & ~v_1643 & ~v_1644 & ~v_1645 & ~v_1646;
assign v_2647 = ~v_1648 & ~v_1649 & ~v_1650 & ~v_1651 & ~v_1652;
assign v_2648 = ~v_1653 & ~v_1654 & ~v_1655 & ~v_1656 & ~v_1657;
assign v_2649 = ~v_1658 & ~v_1659 & ~v_1660 & ~v_1661 & ~v_1662;
assign v_2650 = ~v_1663 & ~v_1664 & ~v_1665 & ~v_1666 & ~v_1667;
assign v_2651 = ~v_1670 & ~v_1671 & ~v_1672 & ~v_1673 & ~v_1674;
assign v_2652 = ~v_1675 & ~v_1676 & ~v_1677 & ~v_1678 & ~v_1679;
assign v_2653 = ~v_1680 & ~v_1681 & ~v_1682 & ~v_1683 & ~v_1684;
assign v_2654 = ~v_1685 & ~v_1686 & ~v_1687 & ~v_1688 & ~v_1689;
assign v_2655 = ~v_1691 & ~v_1692 & ~v_1693 & ~v_1694 & ~v_1695;
assign v_2656 = ~v_1696 & ~v_1697 & ~v_1698 & ~v_1699 & ~v_1700;
assign v_2657 = ~v_1701 & ~v_1702 & ~v_1703 & ~v_1704 & ~v_1705;
assign v_2658 = ~v_1706 & ~v_1707 & ~v_1708 & ~v_1709 & ~v_1710;
assign v_2659 = ~v_1712 & ~v_1713 & ~v_1714 & ~v_1715 & ~v_1716;
assign v_2660 = ~v_1717 & ~v_1718 & ~v_1719 & ~v_1720 & ~v_1721;
assign v_2661 = ~v_1722 & ~v_1723 & ~v_1724 & ~v_1725 & ~v_1726;
assign v_2662 = ~v_1727 & ~v_1728 & ~v_1729 & ~v_1730 & ~v_1731;
assign v_2663 = ~v_1734 & ~v_1735 & ~v_1736 & ~v_1737 & ~v_1738;
assign v_2664 = ~v_1739 & ~v_1740 & ~v_1741 & ~v_1742 & ~v_1743;
assign v_2665 = ~v_1744 & ~v_1745 & ~v_1746 & ~v_1747 & ~v_1748;
assign v_2666 = ~v_1749 & ~v_1750 & ~v_1751 & ~v_1752 & ~v_1753;
assign v_2667 = ~v_1755 & ~v_1756 & ~v_1757 & ~v_1758 & ~v_1759;
assign v_2668 = ~v_1760 & ~v_1761 & ~v_1762 & ~v_1763 & ~v_1764;
assign v_2669 = ~v_1765 & ~v_1766 & ~v_1767 & ~v_1768 & ~v_1769;
assign v_2670 = ~v_1770 & ~v_1771 & ~v_1772 & ~v_1773 & ~v_1774;
assign v_2671 = ~v_1776 & ~v_1777 & ~v_1778 & ~v_1779 & ~v_1780;
assign v_2672 = ~v_1781 & ~v_1782 & ~v_1783 & ~v_1784 & ~v_1785;
assign v_2673 = ~v_1786 & ~v_1787 & ~v_1788 & ~v_1789 & ~v_1790;
assign v_2674 = ~v_1791 & ~v_1792 & ~v_1793 & ~v_1794 & ~v_1795;
assign v_2675 = ~v_1798 & ~v_1799 & ~v_1800 & ~v_1801 & ~v_1802;
assign v_2676 = ~v_1803 & ~v_1804 & ~v_1805 & ~v_1806 & ~v_1807;
assign v_2677 = ~v_1808 & ~v_1809 & ~v_1810 & ~v_1811 & ~v_1812;
assign v_2678 = ~v_1813 & ~v_1814 & ~v_1815 & ~v_1816 & ~v_1817;
assign v_2679 = ~v_1819 & ~v_1820 & ~v_1821 & ~v_1822 & ~v_1823;
assign v_2680 = ~v_1824 & ~v_1825 & ~v_1826 & ~v_1827 & ~v_1828;
assign v_2681 = ~v_1829 & ~v_1830 & ~v_1831 & ~v_1832 & ~v_1833;
assign v_2682 = ~v_1834 & ~v_1835 & ~v_1836 & ~v_1837 & ~v_1838;
assign v_2683 = ~v_1840 & ~v_1841 & ~v_1842 & ~v_1843 & ~v_1844;
assign v_2684 = ~v_1845 & ~v_1846 & ~v_1847 & ~v_1848 & ~v_1849;
assign v_2685 = ~v_1850 & ~v_1851 & ~v_1852 & ~v_1853 & ~v_1854;
assign v_2686 = ~v_1855 & ~v_1856 & ~v_1857 & ~v_1858 & ~v_1859;
assign v_2687 = ~v_1862 & ~v_1863 & ~v_1864 & ~v_1865 & ~v_1866;
assign v_2688 = ~v_1867 & ~v_1868 & ~v_1869 & ~v_1870 & ~v_1871;
assign v_2689 = ~v_1872 & ~v_1873 & ~v_1874 & ~v_1875 & ~v_1876;
assign v_2690 = ~v_1877 & ~v_1878 & ~v_1879 & ~v_1880 & ~v_1881;
assign v_2691 = ~v_1883 & ~v_1884 & ~v_1885 & ~v_1886 & ~v_1887;
assign v_2692 = ~v_1888 & ~v_1889 & ~v_1890 & ~v_1891 & ~v_1892;
assign v_2693 = ~v_1893 & ~v_1894 & ~v_1895 & ~v_1896 & ~v_1897;
assign v_2694 = ~v_1898 & ~v_1899 & ~v_1900 & ~v_1901 & ~v_1902;
assign v_2695 = ~v_1904 & ~v_1905 & ~v_1906 & ~v_1907 & ~v_1908;
assign v_2696 = ~v_1909 & ~v_1910 & ~v_1911 & ~v_1912 & ~v_1913;
assign v_2697 = ~v_1914 & ~v_1915 & ~v_1916 & ~v_1917 & ~v_1918;
assign v_2698 = ~v_1919 & ~v_1920 & ~v_1921 & ~v_1922 & ~v_1923;
assign v_2699 = ~v_1926 & ~v_1927 & ~v_1928 & ~v_1929 & ~v_1930;
assign v_2700 = ~v_1931 & ~v_1932 & ~v_1933 & ~v_1934 & ~v_1935;
assign v_2701 = ~v_1936 & ~v_1937 & ~v_1938 & ~v_1939 & ~v_1940;
assign v_2702 = ~v_1941 & ~v_1942 & ~v_1943 & ~v_1944 & ~v_1945;
assign v_2703 = ~v_1947 & ~v_1948 & ~v_1949 & ~v_1950 & ~v_1951;
assign v_2704 = ~v_1952 & ~v_1953 & ~v_1954 & ~v_1955 & ~v_1956;
assign v_2705 = ~v_1957 & ~v_1958 & ~v_1959 & ~v_1960 & ~v_1961;
assign v_2706 = ~v_1962 & ~v_1963 & ~v_1964 & ~v_1965 & ~v_1966;
assign v_2707 = ~v_1968 & ~v_1969 & ~v_1970 & ~v_1971 & ~v_1972;
assign v_2708 = ~v_1973 & ~v_1974 & ~v_1975 & ~v_1976 & ~v_1977;
assign v_2709 = ~v_1978 & ~v_1979 & ~v_1980 & ~v_1981 & ~v_1982;
assign v_2710 = ~v_1983 & ~v_1984 & ~v_1985 & ~v_1986 & ~v_1987;
assign v_2711 = v_1541 & v_1605 & v_1669 & v_1733 & v_1797;
assign v_2712 = v_1861 & v_1925 & v_1989;
assign v_2713 = ~v_1991 & ~v_1992 & ~v_1993 & ~v_1994 & ~v_1995;
assign v_2714 = ~v_1996 & ~v_1997 & ~v_1998 & ~v_1999 & ~v_2000;
assign v_2715 = ~v_2001 & ~v_2002 & ~v_2003 & ~v_2004 & ~v_2005;
assign v_2716 = ~v_2006 & ~v_2007 & ~v_2008 & ~v_2009 & ~v_2010;
assign v_2717 = ~v_2012 & ~v_2013 & ~v_2014 & ~v_2015 & ~v_2016;
assign v_2718 = ~v_2017 & ~v_2018 & ~v_2019 & ~v_2020 & ~v_2021;
assign v_2719 = ~v_2022 & ~v_2023 & ~v_2024 & ~v_2025 & ~v_2026;
assign v_2720 = ~v_2027 & ~v_2028 & ~v_2029 & ~v_2030 & ~v_2031;
assign v_2721 = ~v_2033 & ~v_2034 & ~v_2035 & ~v_2036 & ~v_2037;
assign v_2722 = ~v_2038 & ~v_2039 & ~v_2040 & ~v_2041 & ~v_2042;
assign v_2723 = ~v_2043 & ~v_2044 & ~v_2045 & ~v_2046 & ~v_2047;
assign v_2724 = ~v_2048 & ~v_2049 & ~v_2050 & ~v_2051 & ~v_2052;
assign v_2725 = ~v_2055 & ~v_2056 & ~v_2057 & ~v_2058 & ~v_2059;
assign v_2726 = ~v_2060 & ~v_2061 & ~v_2062 & ~v_2063 & ~v_2064;
assign v_2727 = ~v_2065 & ~v_2066 & ~v_2067 & ~v_2068 & ~v_2069;
assign v_2728 = ~v_2070 & ~v_2071 & ~v_2072 & ~v_2073 & ~v_2074;
assign v_2729 = ~v_2076 & ~v_2077 & ~v_2078 & ~v_2079 & ~v_2080;
assign v_2730 = ~v_2081 & ~v_2082 & ~v_2083 & ~v_2084 & ~v_2085;
assign v_2731 = ~v_2086 & ~v_2087 & ~v_2088 & ~v_2089 & ~v_2090;
assign v_2732 = ~v_2091 & ~v_2092 & ~v_2093 & ~v_2094 & ~v_2095;
assign v_2733 = ~v_2097 & ~v_2098 & ~v_2099 & ~v_2100 & ~v_2101;
assign v_2734 = ~v_2102 & ~v_2103 & ~v_2104 & ~v_2105 & ~v_2106;
assign v_2735 = ~v_2107 & ~v_2108 & ~v_2109 & ~v_2110 & ~v_2111;
assign v_2736 = ~v_2112 & ~v_2113 & ~v_2114 & ~v_2115 & ~v_2116;
assign v_2737 = ~v_2119 & ~v_2120 & ~v_2121 & ~v_2122 & ~v_2123;
assign v_2738 = ~v_2124 & ~v_2125 & ~v_2126 & ~v_2127 & ~v_2128;
assign v_2739 = ~v_2129 & ~v_2130 & ~v_2131 & ~v_2132 & ~v_2133;
assign v_2740 = ~v_2134 & ~v_2135 & ~v_2136 & ~v_2137 & ~v_2138;
assign v_2741 = ~v_2140 & ~v_2141 & ~v_2142 & ~v_2143 & ~v_2144;
assign v_2742 = ~v_2145 & ~v_2146 & ~v_2147 & ~v_2148 & ~v_2149;
assign v_2743 = ~v_2150 & ~v_2151 & ~v_2152 & ~v_2153 & ~v_2154;
assign v_2744 = ~v_2155 & ~v_2156 & ~v_2157 & ~v_2158 & ~v_2159;
assign v_2745 = ~v_2161 & ~v_2162 & ~v_2163 & ~v_2164 & ~v_2165;
assign v_2746 = ~v_2166 & ~v_2167 & ~v_2168 & ~v_2169 & ~v_2170;
assign v_2747 = ~v_2171 & ~v_2172 & ~v_2173 & ~v_2174 & ~v_2175;
assign v_2748 = ~v_2176 & ~v_2177 & ~v_2178 & ~v_2179 & ~v_2180;
assign v_2749 = ~v_2183 & ~v_2184 & ~v_2185 & ~v_2186 & ~v_2187;
assign v_2750 = ~v_2188 & ~v_2189 & ~v_2190 & ~v_2191 & ~v_2192;
assign v_2751 = ~v_2193 & ~v_2194 & ~v_2195 & ~v_2196 & ~v_2197;
assign v_2752 = ~v_2198 & ~v_2199 & ~v_2200 & ~v_2201 & ~v_2202;
assign v_2753 = ~v_2204 & ~v_2205 & ~v_2206 & ~v_2207 & ~v_2208;
assign v_2754 = ~v_2209 & ~v_2210 & ~v_2211 & ~v_2212 & ~v_2213;
assign v_2755 = ~v_2214 & ~v_2215 & ~v_2216 & ~v_2217 & ~v_2218;
assign v_2756 = ~v_2219 & ~v_2220 & ~v_2221 & ~v_2222 & ~v_2223;
assign v_2757 = ~v_2225 & ~v_2226 & ~v_2227 & ~v_2228 & ~v_2229;
assign v_2758 = ~v_2230 & ~v_2231 & ~v_2232 & ~v_2233 & ~v_2234;
assign v_2759 = ~v_2235 & ~v_2236 & ~v_2237 & ~v_2238 & ~v_2239;
assign v_2760 = ~v_2240 & ~v_2241 & ~v_2242 & ~v_2243 & ~v_2244;
assign v_2761 = ~v_2247 & ~v_2248 & ~v_2249 & ~v_2250 & ~v_2251;
assign v_2762 = ~v_2252 & ~v_2253 & ~v_2254 & ~v_2255 & ~v_2256;
assign v_2763 = ~v_2257 & ~v_2258 & ~v_2259 & ~v_2260 & ~v_2261;
assign v_2764 = ~v_2262 & ~v_2263 & ~v_2264 & ~v_2265 & ~v_2266;
assign v_2765 = ~v_2268 & ~v_2269 & ~v_2270 & ~v_2271 & ~v_2272;
assign v_2766 = ~v_2273 & ~v_2274 & ~v_2275 & ~v_2276 & ~v_2277;
assign v_2767 = ~v_2278 & ~v_2279 & ~v_2280 & ~v_2281 & ~v_2282;
assign v_2768 = ~v_2283 & ~v_2284 & ~v_2285 & ~v_2286 & ~v_2287;
assign v_2769 = ~v_2289 & ~v_2290 & ~v_2291 & ~v_2292 & ~v_2293;
assign v_2770 = ~v_2294 & ~v_2295 & ~v_2296 & ~v_2297 & ~v_2298;
assign v_2771 = ~v_2299 & ~v_2300 & ~v_2301 & ~v_2302 & ~v_2303;
assign v_2772 = ~v_2304 & ~v_2305 & ~v_2306 & ~v_2307 & ~v_2308;
assign v_2773 = ~v_2311 & ~v_2312 & ~v_2313 & ~v_2314 & ~v_2315;
assign v_2774 = ~v_2316 & ~v_2317 & ~v_2318 & ~v_2319 & ~v_2320;
assign v_2775 = ~v_2321 & ~v_2322 & ~v_2323 & ~v_2324 & ~v_2325;
assign v_2776 = ~v_2326 & ~v_2327 & ~v_2328 & ~v_2329 & ~v_2330;
assign v_2777 = ~v_2332 & ~v_2333 & ~v_2334 & ~v_2335 & ~v_2336;
assign v_2778 = ~v_2337 & ~v_2338 & ~v_2339 & ~v_2340 & ~v_2341;
assign v_2779 = ~v_2342 & ~v_2343 & ~v_2344 & ~v_2345 & ~v_2346;
assign v_2780 = ~v_2347 & ~v_2348 & ~v_2349 & ~v_2350 & ~v_2351;
assign v_2781 = ~v_2353 & ~v_2354 & ~v_2355 & ~v_2356 & ~v_2357;
assign v_2782 = ~v_2358 & ~v_2359 & ~v_2360 & ~v_2361 & ~v_2362;
assign v_2783 = ~v_2363 & ~v_2364 & ~v_2365 & ~v_2366 & ~v_2367;
assign v_2784 = ~v_2368 & ~v_2369 & ~v_2370 & ~v_2371 & ~v_2372;
assign v_2785 = ~v_2375 & ~v_2376 & ~v_2377 & ~v_2378 & ~v_2379;
assign v_2786 = ~v_2380 & ~v_2381 & ~v_2382 & ~v_2383 & ~v_2384;
assign v_2787 = ~v_2385 & ~v_2386 & ~v_2387 & ~v_2388 & ~v_2389;
assign v_2788 = ~v_2390 & ~v_2391 & ~v_2392 & ~v_2393 & ~v_2394;
assign v_2789 = ~v_2396 & ~v_2397 & ~v_2398 & ~v_2399 & ~v_2400;
assign v_2790 = ~v_2401 & ~v_2402 & ~v_2403 & ~v_2404 & ~v_2405;
assign v_2791 = ~v_2406 & ~v_2407 & ~v_2408 & ~v_2409 & ~v_2410;
assign v_2792 = ~v_2411 & ~v_2412 & ~v_2413 & ~v_2414 & ~v_2415;
assign v_2793 = ~v_2417 & ~v_2418 & ~v_2419 & ~v_2420 & ~v_2421;
assign v_2794 = ~v_2422 & ~v_2423 & ~v_2424 & ~v_2425 & ~v_2426;
assign v_2795 = ~v_2427 & ~v_2428 & ~v_2429 & ~v_2430 & ~v_2431;
assign v_2796 = ~v_2432 & ~v_2433 & ~v_2434 & ~v_2435 & ~v_2436;
assign v_2797 = ~v_2439 & ~v_2440 & ~v_2441 & ~v_2442 & ~v_2443;
assign v_2798 = ~v_2444 & ~v_2445 & ~v_2446 & ~v_2447 & ~v_2448;
assign v_2799 = ~v_2449 & ~v_2450 & ~v_2451 & ~v_2452 & ~v_2453;
assign v_2800 = ~v_2454 & ~v_2455 & ~v_2456 & ~v_2457 & ~v_2458;
assign v_2801 = ~v_2460 & ~v_2461 & ~v_2462 & ~v_2463 & ~v_2464;
assign v_2802 = ~v_2465 & ~v_2466 & ~v_2467 & ~v_2468 & ~v_2469;
assign v_2803 = ~v_2470 & ~v_2471 & ~v_2472 & ~v_2473 & ~v_2474;
assign v_2804 = ~v_2475 & ~v_2476 & ~v_2477 & ~v_2478 & ~v_2479;
assign v_2805 = ~v_2481 & ~v_2482 & ~v_2483 & ~v_2484 & ~v_2485;
assign v_2806 = ~v_2486 & ~v_2487 & ~v_2488 & ~v_2489 & ~v_2490;
assign v_2807 = ~v_2491 & ~v_2492 & ~v_2493 & ~v_2494 & ~v_2495;
assign v_2808 = ~v_2496 & ~v_2497 & ~v_2498 & ~v_2499 & ~v_2500;
assign v_2503 = v_2809 | v_2810;
assign v_2809 = v_2054 | v_2118 | v_2182 | v_2246 | v_2310;
assign v_2810 = v_2374 | v_2438 | v_2502;
assign v_1025 = v_21 ^ v_61;
assign v_1026 = v_22 ^ v_62;
assign v_1027 = v_23 ^ v_63;
assign v_1028 = v_24 ^ v_64;
assign v_1029 = v_25 ^ v_65;
assign v_1030 = v_26 ^ v_66;
assign v_1031 = v_27 ^ v_67;
assign v_1032 = v_28 ^ v_68;
assign v_1033 = v_29 ^ v_69;
assign v_1034 = v_30 ^ v_70;
assign v_1035 = v_31 ^ v_71;
assign v_1036 = v_32 ^ v_72;
assign v_1037 = v_33 ^ v_73;
assign v_1038 = v_34 ^ v_74;
assign v_1039 = v_35 ^ v_75;
assign v_1040 = v_36 ^ v_76;
assign v_1041 = v_37 ^ v_77;
assign v_1042 = v_38 ^ v_78;
assign v_1043 = v_39 ^ v_79;
assign v_1044 = v_40 ^ v_80;
assign v_1046 = v_41 ^ v_81;
assign v_1047 = v_42 ^ v_82;
assign v_1048 = v_43 ^ v_83;
assign v_1049 = v_44 ^ v_84;
assign v_1050 = v_45 ^ v_85;
assign v_1051 = v_46 ^ v_86;
assign v_1052 = v_47 ^ v_87;
assign v_1053 = v_48 ^ v_88;
assign v_1054 = v_49 ^ v_89;
assign v_1055 = v_50 ^ v_90;
assign v_1056 = v_51 ^ v_91;
assign v_1057 = v_52 ^ v_92;
assign v_1058 = v_53 ^ v_93;
assign v_1059 = v_54 ^ v_94;
assign v_1060 = v_55 ^ v_95;
assign v_1061 = v_56 ^ v_96;
assign v_1062 = v_57 ^ v_97;
assign v_1063 = v_58 ^ v_98;
assign v_1064 = v_59 ^ v_99;
assign v_1065 = v_60 ^ v_100;
assign v_1067 = v_1 ^ v_101;
assign v_1068 = v_2 ^ v_102;
assign v_1069 = v_3 ^ v_103;
assign v_1070 = v_4 ^ v_104;
assign v_1071 = v_5 ^ v_105;
assign v_1072 = v_6 ^ v_106;
assign v_1073 = v_7 ^ v_107;
assign v_1074 = v_8 ^ v_108;
assign v_1075 = v_9 ^ v_109;
assign v_1076 = v_10 ^ v_110;
assign v_1077 = v_11 ^ v_111;
assign v_1078 = v_12 ^ v_112;
assign v_1079 = v_13 ^ v_113;
assign v_1080 = v_14 ^ v_114;
assign v_1081 = v_15 ^ v_115;
assign v_1082 = v_16 ^ v_116;
assign v_1083 = v_17 ^ v_117;
assign v_1084 = v_18 ^ v_118;
assign v_1085 = v_19 ^ v_119;
assign v_1086 = v_20 ^ v_120;
assign v_1089 = v_81 ^ v_121;
assign v_1090 = v_82 ^ v_122;
assign v_1091 = v_83 ^ v_123;
assign v_1092 = v_84 ^ v_124;
assign v_1093 = v_85 ^ v_125;
assign v_1094 = v_86 ^ v_126;
assign v_1095 = v_87 ^ v_127;
assign v_1096 = v_88 ^ v_128;
assign v_1097 = v_89 ^ v_129;
assign v_1098 = v_90 ^ v_130;
assign v_1099 = v_91 ^ v_131;
assign v_1100 = v_92 ^ v_132;
assign v_1101 = v_93 ^ v_133;
assign v_1102 = v_94 ^ v_134;
assign v_1103 = v_95 ^ v_135;
assign v_1104 = v_96 ^ v_136;
assign v_1105 = v_97 ^ v_137;
assign v_1106 = v_98 ^ v_138;
assign v_1107 = v_99 ^ v_139;
assign v_1108 = v_100 ^ v_140;
assign v_1110 = v_101 ^ v_141;
assign v_1111 = v_102 ^ v_142;
assign v_1112 = v_103 ^ v_143;
assign v_1113 = v_104 ^ v_144;
assign v_1114 = v_105 ^ v_145;
assign v_1115 = v_106 ^ v_146;
assign v_1116 = v_107 ^ v_147;
assign v_1117 = v_108 ^ v_148;
assign v_1118 = v_109 ^ v_149;
assign v_1119 = v_110 ^ v_150;
assign v_1120 = v_111 ^ v_151;
assign v_1121 = v_112 ^ v_152;
assign v_1122 = v_113 ^ v_153;
assign v_1123 = v_114 ^ v_154;
assign v_1124 = v_115 ^ v_155;
assign v_1125 = v_116 ^ v_156;
assign v_1126 = v_117 ^ v_157;
assign v_1127 = v_118 ^ v_158;
assign v_1128 = v_119 ^ v_159;
assign v_1129 = v_120 ^ v_160;
assign v_1131 = v_61 ^ v_161;
assign v_1132 = v_62 ^ v_162;
assign v_1133 = v_63 ^ v_163;
assign v_1134 = v_64 ^ v_164;
assign v_1135 = v_65 ^ v_165;
assign v_1136 = v_66 ^ v_166;
assign v_1137 = v_67 ^ v_167;
assign v_1138 = v_68 ^ v_168;
assign v_1139 = v_69 ^ v_169;
assign v_1140 = v_70 ^ v_170;
assign v_1141 = v_71 ^ v_171;
assign v_1142 = v_72 ^ v_172;
assign v_1143 = v_73 ^ v_173;
assign v_1144 = v_74 ^ v_174;
assign v_1145 = v_75 ^ v_175;
assign v_1146 = v_76 ^ v_176;
assign v_1147 = v_77 ^ v_177;
assign v_1148 = v_78 ^ v_178;
assign v_1149 = v_79 ^ v_179;
assign v_1150 = v_80 ^ v_180;
assign v_1153 = v_141 ^ v_181;
assign v_1154 = v_142 ^ v_182;
assign v_1155 = v_143 ^ v_183;
assign v_1156 = v_144 ^ v_184;
assign v_1157 = v_145 ^ v_185;
assign v_1158 = v_146 ^ v_186;
assign v_1159 = v_147 ^ v_187;
assign v_1160 = v_148 ^ v_188;
assign v_1161 = v_149 ^ v_189;
assign v_1162 = v_150 ^ v_190;
assign v_1163 = v_151 ^ v_191;
assign v_1164 = v_152 ^ v_192;
assign v_1165 = v_153 ^ v_193;
assign v_1166 = v_154 ^ v_194;
assign v_1167 = v_155 ^ v_195;
assign v_1168 = v_156 ^ v_196;
assign v_1169 = v_157 ^ v_197;
assign v_1170 = v_158 ^ v_198;
assign v_1171 = v_159 ^ v_199;
assign v_1172 = v_160 ^ v_200;
assign v_1174 = v_161 ^ v_201;
assign v_1175 = v_162 ^ v_202;
assign v_1176 = v_163 ^ v_203;
assign v_1177 = v_164 ^ v_204;
assign v_1178 = v_165 ^ v_205;
assign v_1179 = v_166 ^ v_206;
assign v_1180 = v_167 ^ v_207;
assign v_1181 = v_168 ^ v_208;
assign v_1182 = v_169 ^ v_209;
assign v_1183 = v_170 ^ v_210;
assign v_1184 = v_171 ^ v_211;
assign v_1185 = v_172 ^ v_212;
assign v_1186 = v_173 ^ v_213;
assign v_1187 = v_174 ^ v_214;
assign v_1188 = v_175 ^ v_215;
assign v_1189 = v_176 ^ v_216;
assign v_1190 = v_177 ^ v_217;
assign v_1191 = v_178 ^ v_218;
assign v_1192 = v_179 ^ v_219;
assign v_1193 = v_180 ^ v_220;
assign v_1195 = v_121 ^ v_221;
assign v_1196 = v_122 ^ v_222;
assign v_1197 = v_123 ^ v_223;
assign v_1198 = v_124 ^ v_224;
assign v_1199 = v_125 ^ v_225;
assign v_1200 = v_126 ^ v_226;
assign v_1201 = v_127 ^ v_227;
assign v_1202 = v_128 ^ v_228;
assign v_1203 = v_129 ^ v_229;
assign v_1204 = v_130 ^ v_230;
assign v_1205 = v_131 ^ v_231;
assign v_1206 = v_132 ^ v_232;
assign v_1207 = v_133 ^ v_233;
assign v_1208 = v_134 ^ v_234;
assign v_1209 = v_135 ^ v_235;
assign v_1210 = v_136 ^ v_236;
assign v_1211 = v_137 ^ v_237;
assign v_1212 = v_138 ^ v_238;
assign v_1213 = v_139 ^ v_239;
assign v_1214 = v_140 ^ v_240;
assign v_1217 = v_201 ^ v_241;
assign v_1218 = v_202 ^ v_242;
assign v_1219 = v_203 ^ v_243;
assign v_1220 = v_204 ^ v_244;
assign v_1221 = v_205 ^ v_245;
assign v_1222 = v_206 ^ v_246;
assign v_1223 = v_207 ^ v_247;
assign v_1224 = v_208 ^ v_248;
assign v_1225 = v_209 ^ v_249;
assign v_1226 = v_210 ^ v_250;
assign v_1227 = v_211 ^ v_251;
assign v_1228 = v_212 ^ v_252;
assign v_1229 = v_213 ^ v_253;
assign v_1230 = v_214 ^ v_254;
assign v_1231 = v_215 ^ v_255;
assign v_1232 = v_216 ^ v_256;
assign v_1233 = v_217 ^ v_257;
assign v_1234 = v_218 ^ v_258;
assign v_1235 = v_219 ^ v_259;
assign v_1236 = v_220 ^ v_260;
assign v_1238 = v_221 ^ v_261;
assign v_1239 = v_222 ^ v_262;
assign v_1240 = v_223 ^ v_263;
assign v_1241 = v_224 ^ v_264;
assign v_1242 = v_225 ^ v_265;
assign v_1243 = v_226 ^ v_266;
assign v_1244 = v_227 ^ v_267;
assign v_1245 = v_228 ^ v_268;
assign v_1246 = v_229 ^ v_269;
assign v_1247 = v_230 ^ v_270;
assign v_1248 = v_231 ^ v_271;
assign v_1249 = v_232 ^ v_272;
assign v_1250 = v_233 ^ v_273;
assign v_1251 = v_234 ^ v_274;
assign v_1252 = v_235 ^ v_275;
assign v_1253 = v_236 ^ v_276;
assign v_1254 = v_237 ^ v_277;
assign v_1255 = v_238 ^ v_278;
assign v_1256 = v_239 ^ v_279;
assign v_1257 = v_240 ^ v_280;
assign v_1259 = v_181 ^ v_281;
assign v_1260 = v_182 ^ v_282;
assign v_1261 = v_183 ^ v_283;
assign v_1262 = v_184 ^ v_284;
assign v_1263 = v_185 ^ v_285;
assign v_1264 = v_186 ^ v_286;
assign v_1265 = v_187 ^ v_287;
assign v_1266 = v_188 ^ v_288;
assign v_1267 = v_189 ^ v_289;
assign v_1268 = v_190 ^ v_290;
assign v_1269 = v_191 ^ v_291;
assign v_1270 = v_192 ^ v_292;
assign v_1271 = v_193 ^ v_293;
assign v_1272 = v_194 ^ v_294;
assign v_1273 = v_195 ^ v_295;
assign v_1274 = v_196 ^ v_296;
assign v_1275 = v_197 ^ v_297;
assign v_1276 = v_198 ^ v_298;
assign v_1277 = v_199 ^ v_299;
assign v_1278 = v_200 ^ v_300;
assign v_1281 = v_261 ^ v_301;
assign v_1282 = v_262 ^ v_302;
assign v_1283 = v_263 ^ v_303;
assign v_1284 = v_264 ^ v_304;
assign v_1285 = v_265 ^ v_305;
assign v_1286 = v_266 ^ v_306;
assign v_1287 = v_267 ^ v_307;
assign v_1288 = v_268 ^ v_308;
assign v_1289 = v_269 ^ v_309;
assign v_1290 = v_270 ^ v_310;
assign v_1291 = v_271 ^ v_311;
assign v_1292 = v_272 ^ v_312;
assign v_1293 = v_273 ^ v_313;
assign v_1294 = v_274 ^ v_314;
assign v_1295 = v_275 ^ v_315;
assign v_1296 = v_276 ^ v_316;
assign v_1297 = v_277 ^ v_317;
assign v_1298 = v_278 ^ v_318;
assign v_1299 = v_279 ^ v_319;
assign v_1300 = v_280 ^ v_320;
assign v_1302 = v_281 ^ v_321;
assign v_1303 = v_282 ^ v_322;
assign v_1304 = v_283 ^ v_323;
assign v_1305 = v_284 ^ v_324;
assign v_1306 = v_285 ^ v_325;
assign v_1307 = v_286 ^ v_326;
assign v_1308 = v_287 ^ v_327;
assign v_1309 = v_288 ^ v_328;
assign v_1310 = v_289 ^ v_329;
assign v_1311 = v_290 ^ v_330;
assign v_1312 = v_291 ^ v_331;
assign v_1313 = v_292 ^ v_332;
assign v_1314 = v_293 ^ v_333;
assign v_1315 = v_294 ^ v_334;
assign v_1316 = v_295 ^ v_335;
assign v_1317 = v_296 ^ v_336;
assign v_1318 = v_297 ^ v_337;
assign v_1319 = v_298 ^ v_338;
assign v_1320 = v_299 ^ v_339;
assign v_1321 = v_300 ^ v_340;
assign v_1323 = v_241 ^ v_341;
assign v_1324 = v_242 ^ v_342;
assign v_1325 = v_243 ^ v_343;
assign v_1326 = v_244 ^ v_344;
assign v_1327 = v_245 ^ v_345;
assign v_1328 = v_246 ^ v_346;
assign v_1329 = v_247 ^ v_347;
assign v_1330 = v_248 ^ v_348;
assign v_1331 = v_249 ^ v_349;
assign v_1332 = v_250 ^ v_350;
assign v_1333 = v_251 ^ v_351;
assign v_1334 = v_252 ^ v_352;
assign v_1335 = v_253 ^ v_353;
assign v_1336 = v_254 ^ v_354;
assign v_1337 = v_255 ^ v_355;
assign v_1338 = v_256 ^ v_356;
assign v_1339 = v_257 ^ v_357;
assign v_1340 = v_258 ^ v_358;
assign v_1341 = v_259 ^ v_359;
assign v_1342 = v_260 ^ v_360;
assign v_1345 = v_321 ^ v_361;
assign v_1346 = v_322 ^ v_362;
assign v_1347 = v_323 ^ v_363;
assign v_1348 = v_324 ^ v_364;
assign v_1349 = v_325 ^ v_365;
assign v_1350 = v_326 ^ v_366;
assign v_1351 = v_327 ^ v_367;
assign v_1352 = v_328 ^ v_368;
assign v_1353 = v_329 ^ v_369;
assign v_1354 = v_330 ^ v_370;
assign v_1355 = v_331 ^ v_371;
assign v_1356 = v_332 ^ v_372;
assign v_1357 = v_333 ^ v_373;
assign v_1358 = v_334 ^ v_374;
assign v_1359 = v_335 ^ v_375;
assign v_1360 = v_336 ^ v_376;
assign v_1361 = v_337 ^ v_377;
assign v_1362 = v_338 ^ v_378;
assign v_1363 = v_339 ^ v_379;
assign v_1364 = v_340 ^ v_380;
assign v_1366 = v_341 ^ v_381;
assign v_1367 = v_342 ^ v_382;
assign v_1368 = v_343 ^ v_383;
assign v_1369 = v_344 ^ v_384;
assign v_1370 = v_345 ^ v_385;
assign v_1371 = v_346 ^ v_386;
assign v_1372 = v_347 ^ v_387;
assign v_1373 = v_348 ^ v_388;
assign v_1374 = v_349 ^ v_389;
assign v_1375 = v_350 ^ v_390;
assign v_1376 = v_351 ^ v_391;
assign v_1377 = v_352 ^ v_392;
assign v_1378 = v_353 ^ v_393;
assign v_1379 = v_354 ^ v_394;
assign v_1380 = v_355 ^ v_395;
assign v_1381 = v_356 ^ v_396;
assign v_1382 = v_357 ^ v_397;
assign v_1383 = v_358 ^ v_398;
assign v_1384 = v_359 ^ v_399;
assign v_1385 = v_360 ^ v_400;
assign v_1387 = v_301 ^ v_401;
assign v_1388 = v_302 ^ v_402;
assign v_1389 = v_303 ^ v_403;
assign v_1390 = v_304 ^ v_404;
assign v_1391 = v_305 ^ v_405;
assign v_1392 = v_306 ^ v_406;
assign v_1393 = v_307 ^ v_407;
assign v_1394 = v_308 ^ v_408;
assign v_1395 = v_309 ^ v_409;
assign v_1396 = v_310 ^ v_410;
assign v_1397 = v_311 ^ v_411;
assign v_1398 = v_312 ^ v_412;
assign v_1399 = v_313 ^ v_413;
assign v_1400 = v_314 ^ v_414;
assign v_1401 = v_315 ^ v_415;
assign v_1402 = v_316 ^ v_416;
assign v_1403 = v_317 ^ v_417;
assign v_1404 = v_318 ^ v_418;
assign v_1405 = v_319 ^ v_419;
assign v_1406 = v_320 ^ v_420;
assign v_1409 = v_381 ^ v_421;
assign v_1410 = v_382 ^ v_422;
assign v_1411 = v_383 ^ v_423;
assign v_1412 = v_384 ^ v_424;
assign v_1413 = v_385 ^ v_425;
assign v_1414 = v_386 ^ v_426;
assign v_1415 = v_387 ^ v_427;
assign v_1416 = v_388 ^ v_428;
assign v_1417 = v_389 ^ v_429;
assign v_1418 = v_390 ^ v_430;
assign v_1419 = v_391 ^ v_431;
assign v_1420 = v_392 ^ v_432;
assign v_1421 = v_393 ^ v_433;
assign v_1422 = v_394 ^ v_434;
assign v_1423 = v_395 ^ v_435;
assign v_1424 = v_396 ^ v_436;
assign v_1425 = v_397 ^ v_437;
assign v_1426 = v_398 ^ v_438;
assign v_1427 = v_399 ^ v_439;
assign v_1428 = v_400 ^ v_440;
assign v_1430 = v_401 ^ v_441;
assign v_1431 = v_402 ^ v_442;
assign v_1432 = v_403 ^ v_443;
assign v_1433 = v_404 ^ v_444;
assign v_1434 = v_405 ^ v_445;
assign v_1435 = v_406 ^ v_446;
assign v_1436 = v_407 ^ v_447;
assign v_1437 = v_408 ^ v_448;
assign v_1438 = v_409 ^ v_449;
assign v_1439 = v_410 ^ v_450;
assign v_1440 = v_411 ^ v_451;
assign v_1441 = v_412 ^ v_452;
assign v_1442 = v_413 ^ v_453;
assign v_1443 = v_414 ^ v_454;
assign v_1444 = v_415 ^ v_455;
assign v_1445 = v_416 ^ v_456;
assign v_1446 = v_417 ^ v_457;
assign v_1447 = v_418 ^ v_458;
assign v_1448 = v_419 ^ v_459;
assign v_1449 = v_420 ^ v_460;
assign v_1451 = v_361 ^ v_461;
assign v_1452 = v_362 ^ v_462;
assign v_1453 = v_363 ^ v_463;
assign v_1454 = v_364 ^ v_464;
assign v_1455 = v_365 ^ v_465;
assign v_1456 = v_366 ^ v_466;
assign v_1457 = v_367 ^ v_467;
assign v_1458 = v_368 ^ v_468;
assign v_1459 = v_369 ^ v_469;
assign v_1460 = v_370 ^ v_470;
assign v_1461 = v_371 ^ v_471;
assign v_1462 = v_372 ^ v_472;
assign v_1463 = v_373 ^ v_473;
assign v_1464 = v_374 ^ v_474;
assign v_1465 = v_375 ^ v_475;
assign v_1466 = v_376 ^ v_476;
assign v_1467 = v_377 ^ v_477;
assign v_1468 = v_378 ^ v_478;
assign v_1469 = v_379 ^ v_479;
assign v_1470 = v_380 ^ v_480;
assign v_1473 = v_441 ^ v_481;
assign v_1474 = v_442 ^ v_482;
assign v_1475 = v_443 ^ v_483;
assign v_1476 = v_444 ^ v_484;
assign v_1477 = v_445 ^ v_485;
assign v_1478 = v_446 ^ v_486;
assign v_1479 = v_447 ^ v_487;
assign v_1480 = v_448 ^ v_488;
assign v_1481 = v_449 ^ v_489;
assign v_1482 = v_450 ^ v_490;
assign v_1483 = v_451 ^ v_491;
assign v_1484 = v_452 ^ v_492;
assign v_1485 = v_453 ^ v_493;
assign v_1486 = v_454 ^ v_494;
assign v_1487 = v_455 ^ v_495;
assign v_1488 = v_456 ^ v_496;
assign v_1489 = v_457 ^ v_497;
assign v_1490 = v_458 ^ v_498;
assign v_1491 = v_459 ^ v_499;
assign v_1492 = v_460 ^ v_500;
assign v_1494 = v_461 ^ v_501;
assign v_1495 = v_462 ^ v_502;
assign v_1496 = v_463 ^ v_503;
assign v_1497 = v_464 ^ v_504;
assign v_1498 = v_465 ^ v_505;
assign v_1499 = v_466 ^ v_506;
assign v_1500 = v_467 ^ v_507;
assign v_1501 = v_468 ^ v_508;
assign v_1502 = v_469 ^ v_509;
assign v_1503 = v_470 ^ v_510;
assign v_1504 = v_471 ^ v_511;
assign v_1505 = v_472 ^ v_512;
assign v_1506 = v_473 ^ v_513;
assign v_1507 = v_474 ^ v_514;
assign v_1508 = v_475 ^ v_515;
assign v_1509 = v_476 ^ v_516;
assign v_1510 = v_477 ^ v_517;
assign v_1511 = v_478 ^ v_518;
assign v_1512 = v_479 ^ v_519;
assign v_1513 = v_480 ^ v_520;
assign v_1515 = v_421 ^ v_521;
assign v_1516 = v_422 ^ v_522;
assign v_1517 = v_423 ^ v_523;
assign v_1518 = v_424 ^ v_524;
assign v_1519 = v_425 ^ v_525;
assign v_1520 = v_426 ^ v_526;
assign v_1521 = v_427 ^ v_527;
assign v_1522 = v_428 ^ v_528;
assign v_1523 = v_429 ^ v_529;
assign v_1524 = v_430 ^ v_530;
assign v_1525 = v_431 ^ v_531;
assign v_1526 = v_432 ^ v_532;
assign v_1527 = v_433 ^ v_533;
assign v_1528 = v_434 ^ v_534;
assign v_1529 = v_435 ^ v_535;
assign v_1530 = v_436 ^ v_536;
assign v_1531 = v_437 ^ v_537;
assign v_1532 = v_438 ^ v_538;
assign v_1533 = v_439 ^ v_539;
assign v_1534 = v_440 ^ v_540;
assign v_1542 = v_561 ^ v_601;
assign v_1543 = v_562 ^ v_602;
assign v_1544 = v_563 ^ v_603;
assign v_1545 = v_564 ^ v_604;
assign v_1546 = v_565 ^ v_605;
assign v_1547 = v_566 ^ v_606;
assign v_1548 = v_567 ^ v_607;
assign v_1549 = v_568 ^ v_608;
assign v_1550 = v_569 ^ v_609;
assign v_1551 = v_570 ^ v_610;
assign v_1552 = v_571 ^ v_611;
assign v_1553 = v_572 ^ v_612;
assign v_1554 = v_573 ^ v_613;
assign v_1555 = v_574 ^ v_614;
assign v_1556 = v_575 ^ v_615;
assign v_1557 = v_576 ^ v_616;
assign v_1558 = v_577 ^ v_617;
assign v_1559 = v_578 ^ v_618;
assign v_1560 = v_579 ^ v_619;
assign v_1561 = v_580 ^ v_620;
assign v_1563 = v_581 ^ v_621;
assign v_1564 = v_582 ^ v_622;
assign v_1565 = v_583 ^ v_623;
assign v_1566 = v_584 ^ v_624;
assign v_1567 = v_585 ^ v_625;
assign v_1568 = v_586 ^ v_626;
assign v_1569 = v_587 ^ v_627;
assign v_1570 = v_588 ^ v_628;
assign v_1571 = v_589 ^ v_629;
assign v_1572 = v_590 ^ v_630;
assign v_1573 = v_591 ^ v_631;
assign v_1574 = v_592 ^ v_632;
assign v_1575 = v_593 ^ v_633;
assign v_1576 = v_594 ^ v_634;
assign v_1577 = v_595 ^ v_635;
assign v_1578 = v_596 ^ v_636;
assign v_1579 = v_597 ^ v_637;
assign v_1580 = v_598 ^ v_638;
assign v_1581 = v_599 ^ v_639;
assign v_1582 = v_600 ^ v_640;
assign v_1584 = v_541 ^ v_641;
assign v_1585 = v_542 ^ v_642;
assign v_1586 = v_543 ^ v_643;
assign v_1587 = v_544 ^ v_644;
assign v_1588 = v_545 ^ v_645;
assign v_1589 = v_546 ^ v_646;
assign v_1590 = v_547 ^ v_647;
assign v_1591 = v_548 ^ v_648;
assign v_1592 = v_549 ^ v_649;
assign v_1593 = v_550 ^ v_650;
assign v_1594 = v_551 ^ v_651;
assign v_1595 = v_552 ^ v_652;
assign v_1596 = v_553 ^ v_653;
assign v_1597 = v_554 ^ v_654;
assign v_1598 = v_555 ^ v_655;
assign v_1599 = v_556 ^ v_656;
assign v_1600 = v_557 ^ v_657;
assign v_1601 = v_558 ^ v_658;
assign v_1602 = v_559 ^ v_659;
assign v_1603 = v_560 ^ v_660;
assign v_1606 = v_621 ^ v_661;
assign v_1607 = v_622 ^ v_662;
assign v_1608 = v_623 ^ v_663;
assign v_1609 = v_624 ^ v_664;
assign v_1610 = v_625 ^ v_665;
assign v_1611 = v_626 ^ v_666;
assign v_1612 = v_627 ^ v_667;
assign v_1613 = v_628 ^ v_668;
assign v_1614 = v_629 ^ v_669;
assign v_1615 = v_630 ^ v_670;
assign v_1616 = v_631 ^ v_671;
assign v_1617 = v_632 ^ v_672;
assign v_1618 = v_633 ^ v_673;
assign v_1619 = v_634 ^ v_674;
assign v_1620 = v_635 ^ v_675;
assign v_1621 = v_636 ^ v_676;
assign v_1622 = v_637 ^ v_677;
assign v_1623 = v_638 ^ v_678;
assign v_1624 = v_639 ^ v_679;
assign v_1625 = v_640 ^ v_680;
assign v_1627 = v_641 ^ v_681;
assign v_1628 = v_642 ^ v_682;
assign v_1629 = v_643 ^ v_683;
assign v_1630 = v_644 ^ v_684;
assign v_1631 = v_645 ^ v_685;
assign v_1632 = v_646 ^ v_686;
assign v_1633 = v_647 ^ v_687;
assign v_1634 = v_648 ^ v_688;
assign v_1635 = v_649 ^ v_689;
assign v_1636 = v_650 ^ v_690;
assign v_1637 = v_651 ^ v_691;
assign v_1638 = v_652 ^ v_692;
assign v_1639 = v_653 ^ v_693;
assign v_1640 = v_654 ^ v_694;
assign v_1641 = v_655 ^ v_695;
assign v_1642 = v_656 ^ v_696;
assign v_1643 = v_657 ^ v_697;
assign v_1644 = v_658 ^ v_698;
assign v_1645 = v_659 ^ v_699;
assign v_1646 = v_660 ^ v_700;
assign v_1648 = v_601 ^ v_701;
assign v_1649 = v_602 ^ v_702;
assign v_1650 = v_603 ^ v_703;
assign v_1651 = v_604 ^ v_704;
assign v_1652 = v_605 ^ v_705;
assign v_1653 = v_606 ^ v_706;
assign v_1654 = v_607 ^ v_707;
assign v_1655 = v_608 ^ v_708;
assign v_1656 = v_609 ^ v_709;
assign v_1657 = v_610 ^ v_710;
assign v_1658 = v_611 ^ v_711;
assign v_1659 = v_612 ^ v_712;
assign v_1660 = v_613 ^ v_713;
assign v_1661 = v_614 ^ v_714;
assign v_1662 = v_615 ^ v_715;
assign v_1663 = v_616 ^ v_716;
assign v_1664 = v_617 ^ v_717;
assign v_1665 = v_618 ^ v_718;
assign v_1666 = v_619 ^ v_719;
assign v_1667 = v_620 ^ v_720;
assign v_1670 = v_681 ^ v_721;
assign v_1671 = v_682 ^ v_722;
assign v_1672 = v_683 ^ v_723;
assign v_1673 = v_684 ^ v_724;
assign v_1674 = v_685 ^ v_725;
assign v_1675 = v_686 ^ v_726;
assign v_1676 = v_687 ^ v_727;
assign v_1677 = v_688 ^ v_728;
assign v_1678 = v_689 ^ v_729;
assign v_1679 = v_690 ^ v_730;
assign v_1680 = v_691 ^ v_731;
assign v_1681 = v_692 ^ v_732;
assign v_1682 = v_693 ^ v_733;
assign v_1683 = v_694 ^ v_734;
assign v_1684 = v_695 ^ v_735;
assign v_1685 = v_696 ^ v_736;
assign v_1686 = v_697 ^ v_737;
assign v_1687 = v_698 ^ v_738;
assign v_1688 = v_699 ^ v_739;
assign v_1689 = v_700 ^ v_740;
assign v_1691 = v_701 ^ v_741;
assign v_1692 = v_702 ^ v_742;
assign v_1693 = v_703 ^ v_743;
assign v_1694 = v_704 ^ v_744;
assign v_1695 = v_705 ^ v_745;
assign v_1696 = v_706 ^ v_746;
assign v_1697 = v_707 ^ v_747;
assign v_1698 = v_708 ^ v_748;
assign v_1699 = v_709 ^ v_749;
assign v_1700 = v_710 ^ v_750;
assign v_1701 = v_711 ^ v_751;
assign v_1702 = v_712 ^ v_752;
assign v_1703 = v_713 ^ v_753;
assign v_1704 = v_714 ^ v_754;
assign v_1705 = v_715 ^ v_755;
assign v_1706 = v_716 ^ v_756;
assign v_1707 = v_717 ^ v_757;
assign v_1708 = v_718 ^ v_758;
assign v_1709 = v_719 ^ v_759;
assign v_1710 = v_720 ^ v_760;
assign v_1712 = v_661 ^ v_761;
assign v_1713 = v_662 ^ v_762;
assign v_1714 = v_663 ^ v_763;
assign v_1715 = v_664 ^ v_764;
assign v_1716 = v_665 ^ v_765;
assign v_1717 = v_666 ^ v_766;
assign v_1718 = v_667 ^ v_767;
assign v_1719 = v_668 ^ v_768;
assign v_1720 = v_669 ^ v_769;
assign v_1721 = v_670 ^ v_770;
assign v_1722 = v_671 ^ v_771;
assign v_1723 = v_672 ^ v_772;
assign v_1724 = v_673 ^ v_773;
assign v_1725 = v_674 ^ v_774;
assign v_1726 = v_675 ^ v_775;
assign v_1727 = v_676 ^ v_776;
assign v_1728 = v_677 ^ v_777;
assign v_1729 = v_678 ^ v_778;
assign v_1730 = v_679 ^ v_779;
assign v_1731 = v_680 ^ v_780;
assign v_1734 = v_741 ^ v_781;
assign v_1735 = v_742 ^ v_782;
assign v_1736 = v_743 ^ v_783;
assign v_1737 = v_744 ^ v_784;
assign v_1738 = v_745 ^ v_785;
assign v_1739 = v_746 ^ v_786;
assign v_1740 = v_747 ^ v_787;
assign v_1741 = v_748 ^ v_788;
assign v_1742 = v_749 ^ v_789;
assign v_1743 = v_750 ^ v_790;
assign v_1744 = v_751 ^ v_791;
assign v_1745 = v_752 ^ v_792;
assign v_1746 = v_753 ^ v_793;
assign v_1747 = v_754 ^ v_794;
assign v_1748 = v_755 ^ v_795;
assign v_1749 = v_756 ^ v_796;
assign v_1750 = v_757 ^ v_797;
assign v_1751 = v_758 ^ v_798;
assign v_1752 = v_759 ^ v_799;
assign v_1753 = v_760 ^ v_800;
assign v_1755 = v_761 ^ v_801;
assign v_1756 = v_762 ^ v_802;
assign v_1757 = v_763 ^ v_803;
assign v_1758 = v_764 ^ v_804;
assign v_1759 = v_765 ^ v_805;
assign v_1760 = v_766 ^ v_806;
assign v_1761 = v_767 ^ v_807;
assign v_1762 = v_768 ^ v_808;
assign v_1763 = v_769 ^ v_809;
assign v_1764 = v_770 ^ v_810;
assign v_1765 = v_771 ^ v_811;
assign v_1766 = v_772 ^ v_812;
assign v_1767 = v_773 ^ v_813;
assign v_1768 = v_774 ^ v_814;
assign v_1769 = v_775 ^ v_815;
assign v_1770 = v_776 ^ v_816;
assign v_1771 = v_777 ^ v_817;
assign v_1772 = v_778 ^ v_818;
assign v_1773 = v_779 ^ v_819;
assign v_1774 = v_780 ^ v_820;
assign v_1776 = v_721 ^ v_821;
assign v_1777 = v_722 ^ v_822;
assign v_1778 = v_723 ^ v_823;
assign v_1779 = v_724 ^ v_824;
assign v_1780 = v_725 ^ v_825;
assign v_1781 = v_726 ^ v_826;
assign v_1782 = v_727 ^ v_827;
assign v_1783 = v_728 ^ v_828;
assign v_1784 = v_729 ^ v_829;
assign v_1785 = v_730 ^ v_830;
assign v_1786 = v_731 ^ v_831;
assign v_1787 = v_732 ^ v_832;
assign v_1788 = v_733 ^ v_833;
assign v_1789 = v_734 ^ v_834;
assign v_1790 = v_735 ^ v_835;
assign v_1791 = v_736 ^ v_836;
assign v_1792 = v_737 ^ v_837;
assign v_1793 = v_738 ^ v_838;
assign v_1794 = v_739 ^ v_839;
assign v_1795 = v_740 ^ v_840;
assign v_1798 = v_801 ^ v_841;
assign v_1799 = v_802 ^ v_842;
assign v_1800 = v_803 ^ v_843;
assign v_1801 = v_804 ^ v_844;
assign v_1802 = v_805 ^ v_845;
assign v_1803 = v_806 ^ v_846;
assign v_1804 = v_807 ^ v_847;
assign v_1805 = v_808 ^ v_848;
assign v_1806 = v_809 ^ v_849;
assign v_1807 = v_810 ^ v_850;
assign v_1808 = v_811 ^ v_851;
assign v_1809 = v_812 ^ v_852;
assign v_1810 = v_813 ^ v_853;
assign v_1811 = v_814 ^ v_854;
assign v_1812 = v_815 ^ v_855;
assign v_1813 = v_816 ^ v_856;
assign v_1814 = v_817 ^ v_857;
assign v_1815 = v_818 ^ v_858;
assign v_1816 = v_819 ^ v_859;
assign v_1817 = v_820 ^ v_860;
assign v_1819 = v_821 ^ v_861;
assign v_1820 = v_822 ^ v_862;
assign v_1821 = v_823 ^ v_863;
assign v_1822 = v_824 ^ v_864;
assign v_1823 = v_825 ^ v_865;
assign v_1824 = v_826 ^ v_866;
assign v_1825 = v_827 ^ v_867;
assign v_1826 = v_828 ^ v_868;
assign v_1827 = v_829 ^ v_869;
assign v_1828 = v_830 ^ v_870;
assign v_1829 = v_831 ^ v_871;
assign v_1830 = v_832 ^ v_872;
assign v_1831 = v_833 ^ v_873;
assign v_1832 = v_834 ^ v_874;
assign v_1833 = v_835 ^ v_875;
assign v_1834 = v_836 ^ v_876;
assign v_1835 = v_837 ^ v_877;
assign v_1836 = v_838 ^ v_878;
assign v_1837 = v_839 ^ v_879;
assign v_1838 = v_840 ^ v_880;
assign v_1840 = v_781 ^ v_881;
assign v_1841 = v_782 ^ v_882;
assign v_1842 = v_783 ^ v_883;
assign v_1843 = v_784 ^ v_884;
assign v_1844 = v_785 ^ v_885;
assign v_1845 = v_786 ^ v_886;
assign v_1846 = v_787 ^ v_887;
assign v_1847 = v_788 ^ v_888;
assign v_1848 = v_789 ^ v_889;
assign v_1849 = v_790 ^ v_890;
assign v_1850 = v_791 ^ v_891;
assign v_1851 = v_792 ^ v_892;
assign v_1852 = v_793 ^ v_893;
assign v_1853 = v_794 ^ v_894;
assign v_1854 = v_795 ^ v_895;
assign v_1855 = v_796 ^ v_896;
assign v_1856 = v_797 ^ v_897;
assign v_1857 = v_798 ^ v_898;
assign v_1858 = v_799 ^ v_899;
assign v_1859 = v_800 ^ v_900;
assign v_1862 = v_861 ^ v_901;
assign v_1863 = v_862 ^ v_902;
assign v_1864 = v_863 ^ v_903;
assign v_1865 = v_864 ^ v_904;
assign v_1866 = v_865 ^ v_905;
assign v_1867 = v_866 ^ v_906;
assign v_1868 = v_867 ^ v_907;
assign v_1869 = v_868 ^ v_908;
assign v_1870 = v_869 ^ v_909;
assign v_1871 = v_870 ^ v_910;
assign v_1872 = v_871 ^ v_911;
assign v_1873 = v_872 ^ v_912;
assign v_1874 = v_873 ^ v_913;
assign v_1875 = v_874 ^ v_914;
assign v_1876 = v_875 ^ v_915;
assign v_1877 = v_876 ^ v_916;
assign v_1878 = v_877 ^ v_917;
assign v_1879 = v_878 ^ v_918;
assign v_1880 = v_879 ^ v_919;
assign v_1881 = v_880 ^ v_920;
assign v_1883 = v_881 ^ v_921;
assign v_1884 = v_882 ^ v_922;
assign v_1885 = v_883 ^ v_923;
assign v_1886 = v_884 ^ v_924;
assign v_1887 = v_885 ^ v_925;
assign v_1888 = v_886 ^ v_926;
assign v_1889 = v_887 ^ v_927;
assign v_1890 = v_888 ^ v_928;
assign v_1891 = v_889 ^ v_929;
assign v_1892 = v_890 ^ v_930;
assign v_1893 = v_891 ^ v_931;
assign v_1894 = v_892 ^ v_932;
assign v_1895 = v_893 ^ v_933;
assign v_1896 = v_894 ^ v_934;
assign v_1897 = v_895 ^ v_935;
assign v_1898 = v_896 ^ v_936;
assign v_1899 = v_897 ^ v_937;
assign v_1900 = v_898 ^ v_938;
assign v_1901 = v_899 ^ v_939;
assign v_1902 = v_900 ^ v_940;
assign v_1904 = v_841 ^ v_941;
assign v_1905 = v_842 ^ v_942;
assign v_1906 = v_843 ^ v_943;
assign v_1907 = v_844 ^ v_944;
assign v_1908 = v_845 ^ v_945;
assign v_1909 = v_846 ^ v_946;
assign v_1910 = v_847 ^ v_947;
assign v_1911 = v_848 ^ v_948;
assign v_1912 = v_849 ^ v_949;
assign v_1913 = v_850 ^ v_950;
assign v_1914 = v_851 ^ v_951;
assign v_1915 = v_852 ^ v_952;
assign v_1916 = v_853 ^ v_953;
assign v_1917 = v_854 ^ v_954;
assign v_1918 = v_855 ^ v_955;
assign v_1919 = v_856 ^ v_956;
assign v_1920 = v_857 ^ v_957;
assign v_1921 = v_858 ^ v_958;
assign v_1922 = v_859 ^ v_959;
assign v_1923 = v_860 ^ v_960;
assign v_1926 = v_921 ^ v_961;
assign v_1927 = v_922 ^ v_962;
assign v_1928 = v_923 ^ v_963;
assign v_1929 = v_924 ^ v_964;
assign v_1930 = v_925 ^ v_965;
assign v_1931 = v_926 ^ v_966;
assign v_1932 = v_927 ^ v_967;
assign v_1933 = v_928 ^ v_968;
assign v_1934 = v_929 ^ v_969;
assign v_1935 = v_930 ^ v_970;
assign v_1936 = v_931 ^ v_971;
assign v_1937 = v_932 ^ v_972;
assign v_1938 = v_933 ^ v_973;
assign v_1939 = v_934 ^ v_974;
assign v_1940 = v_935 ^ v_975;
assign v_1941 = v_936 ^ v_976;
assign v_1942 = v_937 ^ v_977;
assign v_1943 = v_938 ^ v_978;
assign v_1944 = v_939 ^ v_979;
assign v_1945 = v_940 ^ v_980;
assign v_1947 = v_941 ^ v_981;
assign v_1948 = v_942 ^ v_982;
assign v_1949 = v_943 ^ v_983;
assign v_1950 = v_944 ^ v_984;
assign v_1951 = v_945 ^ v_985;
assign v_1952 = v_946 ^ v_986;
assign v_1953 = v_947 ^ v_987;
assign v_1954 = v_948 ^ v_988;
assign v_1955 = v_949 ^ v_989;
assign v_1956 = v_950 ^ v_990;
assign v_1957 = v_951 ^ v_991;
assign v_1958 = v_952 ^ v_992;
assign v_1959 = v_953 ^ v_993;
assign v_1960 = v_954 ^ v_994;
assign v_1961 = v_955 ^ v_995;
assign v_1962 = v_956 ^ v_996;
assign v_1963 = v_957 ^ v_997;
assign v_1964 = v_958 ^ v_998;
assign v_1965 = v_959 ^ v_999;
assign v_1966 = v_960 ^ v_1000;
assign v_1968 = v_901 ^ v_1001;
assign v_1969 = v_902 ^ v_1002;
assign v_1970 = v_903 ^ v_1003;
assign v_1971 = v_904 ^ v_1004;
assign v_1972 = v_905 ^ v_1005;
assign v_1973 = v_906 ^ v_1006;
assign v_1974 = v_907 ^ v_1007;
assign v_1975 = v_908 ^ v_1008;
assign v_1976 = v_909 ^ v_1009;
assign v_1977 = v_910 ^ v_1010;
assign v_1978 = v_911 ^ v_1011;
assign v_1979 = v_912 ^ v_1012;
assign v_1980 = v_913 ^ v_1013;
assign v_1981 = v_914 ^ v_1014;
assign v_1982 = v_915 ^ v_1015;
assign v_1983 = v_916 ^ v_1016;
assign v_1984 = v_917 ^ v_1017;
assign v_1985 = v_918 ^ v_1018;
assign v_1986 = v_919 ^ v_1019;
assign v_1987 = v_920 ^ v_1020;
assign v_1991 = v_541 ^ v_481;
assign v_1992 = v_542 ^ v_482;
assign v_1993 = v_543 ^ v_483;
assign v_1994 = v_544 ^ v_484;
assign v_1995 = v_545 ^ v_485;
assign v_1996 = v_546 ^ v_486;
assign v_1997 = v_547 ^ v_487;
assign v_1998 = v_548 ^ v_488;
assign v_1999 = v_549 ^ v_489;
assign v_2000 = v_550 ^ v_490;
assign v_2001 = v_551 ^ v_491;
assign v_2002 = v_552 ^ v_492;
assign v_2003 = v_553 ^ v_493;
assign v_2004 = v_554 ^ v_494;
assign v_2005 = v_555 ^ v_495;
assign v_2006 = v_556 ^ v_496;
assign v_2007 = v_557 ^ v_497;
assign v_2008 = v_558 ^ v_498;
assign v_2009 = v_559 ^ v_499;
assign v_2010 = v_560 ^ v_500;
assign v_2012 = v_561 ^ v_501;
assign v_2013 = v_562 ^ v_502;
assign v_2014 = v_563 ^ v_503;
assign v_2015 = v_564 ^ v_504;
assign v_2016 = v_565 ^ v_505;
assign v_2017 = v_566 ^ v_506;
assign v_2018 = v_567 ^ v_507;
assign v_2019 = v_568 ^ v_508;
assign v_2020 = v_569 ^ v_509;
assign v_2021 = v_570 ^ v_510;
assign v_2022 = v_571 ^ v_511;
assign v_2023 = v_572 ^ v_512;
assign v_2024 = v_573 ^ v_513;
assign v_2025 = v_574 ^ v_514;
assign v_2026 = v_575 ^ v_515;
assign v_2027 = v_576 ^ v_516;
assign v_2028 = v_577 ^ v_517;
assign v_2029 = v_578 ^ v_518;
assign v_2030 = v_579 ^ v_519;
assign v_2031 = v_580 ^ v_520;
assign v_2033 = v_581 ^ v_521;
assign v_2034 = v_582 ^ v_522;
assign v_2035 = v_583 ^ v_523;
assign v_2036 = v_584 ^ v_524;
assign v_2037 = v_585 ^ v_525;
assign v_2038 = v_586 ^ v_526;
assign v_2039 = v_587 ^ v_527;
assign v_2040 = v_588 ^ v_528;
assign v_2041 = v_589 ^ v_529;
assign v_2042 = v_590 ^ v_530;
assign v_2043 = v_591 ^ v_531;
assign v_2044 = v_592 ^ v_532;
assign v_2045 = v_593 ^ v_533;
assign v_2046 = v_594 ^ v_534;
assign v_2047 = v_595 ^ v_535;
assign v_2048 = v_596 ^ v_536;
assign v_2049 = v_597 ^ v_537;
assign v_2050 = v_598 ^ v_538;
assign v_2051 = v_599 ^ v_539;
assign v_2052 = v_600 ^ v_540;
assign v_2055 = v_601 ^ v_481;
assign v_2056 = v_602 ^ v_482;
assign v_2057 = v_603 ^ v_483;
assign v_2058 = v_604 ^ v_484;
assign v_2059 = v_605 ^ v_485;
assign v_2060 = v_606 ^ v_486;
assign v_2061 = v_607 ^ v_487;
assign v_2062 = v_608 ^ v_488;
assign v_2063 = v_609 ^ v_489;
assign v_2064 = v_610 ^ v_490;
assign v_2065 = v_611 ^ v_491;
assign v_2066 = v_612 ^ v_492;
assign v_2067 = v_613 ^ v_493;
assign v_2068 = v_614 ^ v_494;
assign v_2069 = v_615 ^ v_495;
assign v_2070 = v_616 ^ v_496;
assign v_2071 = v_617 ^ v_497;
assign v_2072 = v_618 ^ v_498;
assign v_2073 = v_619 ^ v_499;
assign v_2074 = v_620 ^ v_500;
assign v_2076 = v_621 ^ v_501;
assign v_2077 = v_622 ^ v_502;
assign v_2078 = v_623 ^ v_503;
assign v_2079 = v_624 ^ v_504;
assign v_2080 = v_625 ^ v_505;
assign v_2081 = v_626 ^ v_506;
assign v_2082 = v_627 ^ v_507;
assign v_2083 = v_628 ^ v_508;
assign v_2084 = v_629 ^ v_509;
assign v_2085 = v_630 ^ v_510;
assign v_2086 = v_631 ^ v_511;
assign v_2087 = v_632 ^ v_512;
assign v_2088 = v_633 ^ v_513;
assign v_2089 = v_634 ^ v_514;
assign v_2090 = v_635 ^ v_515;
assign v_2091 = v_636 ^ v_516;
assign v_2092 = v_637 ^ v_517;
assign v_2093 = v_638 ^ v_518;
assign v_2094 = v_639 ^ v_519;
assign v_2095 = v_640 ^ v_520;
assign v_2097 = v_641 ^ v_521;
assign v_2098 = v_642 ^ v_522;
assign v_2099 = v_643 ^ v_523;
assign v_2100 = v_644 ^ v_524;
assign v_2101 = v_645 ^ v_525;
assign v_2102 = v_646 ^ v_526;
assign v_2103 = v_647 ^ v_527;
assign v_2104 = v_648 ^ v_528;
assign v_2105 = v_649 ^ v_529;
assign v_2106 = v_650 ^ v_530;
assign v_2107 = v_651 ^ v_531;
assign v_2108 = v_652 ^ v_532;
assign v_2109 = v_653 ^ v_533;
assign v_2110 = v_654 ^ v_534;
assign v_2111 = v_655 ^ v_535;
assign v_2112 = v_656 ^ v_536;
assign v_2113 = v_657 ^ v_537;
assign v_2114 = v_658 ^ v_538;
assign v_2115 = v_659 ^ v_539;
assign v_2116 = v_660 ^ v_540;
assign v_2119 = v_661 ^ v_481;
assign v_2120 = v_662 ^ v_482;
assign v_2121 = v_663 ^ v_483;
assign v_2122 = v_664 ^ v_484;
assign v_2123 = v_665 ^ v_485;
assign v_2124 = v_666 ^ v_486;
assign v_2125 = v_667 ^ v_487;
assign v_2126 = v_668 ^ v_488;
assign v_2127 = v_669 ^ v_489;
assign v_2128 = v_670 ^ v_490;
assign v_2129 = v_671 ^ v_491;
assign v_2130 = v_672 ^ v_492;
assign v_2131 = v_673 ^ v_493;
assign v_2132 = v_674 ^ v_494;
assign v_2133 = v_675 ^ v_495;
assign v_2134 = v_676 ^ v_496;
assign v_2135 = v_677 ^ v_497;
assign v_2136 = v_678 ^ v_498;
assign v_2137 = v_679 ^ v_499;
assign v_2138 = v_680 ^ v_500;
assign v_2140 = v_681 ^ v_501;
assign v_2141 = v_682 ^ v_502;
assign v_2142 = v_683 ^ v_503;
assign v_2143 = v_684 ^ v_504;
assign v_2144 = v_685 ^ v_505;
assign v_2145 = v_686 ^ v_506;
assign v_2146 = v_687 ^ v_507;
assign v_2147 = v_688 ^ v_508;
assign v_2148 = v_689 ^ v_509;
assign v_2149 = v_690 ^ v_510;
assign v_2150 = v_691 ^ v_511;
assign v_2151 = v_692 ^ v_512;
assign v_2152 = v_693 ^ v_513;
assign v_2153 = v_694 ^ v_514;
assign v_2154 = v_695 ^ v_515;
assign v_2155 = v_696 ^ v_516;
assign v_2156 = v_697 ^ v_517;
assign v_2157 = v_698 ^ v_518;
assign v_2158 = v_699 ^ v_519;
assign v_2159 = v_700 ^ v_520;
assign v_2161 = v_701 ^ v_521;
assign v_2162 = v_702 ^ v_522;
assign v_2163 = v_703 ^ v_523;
assign v_2164 = v_704 ^ v_524;
assign v_2165 = v_705 ^ v_525;
assign v_2166 = v_706 ^ v_526;
assign v_2167 = v_707 ^ v_527;
assign v_2168 = v_708 ^ v_528;
assign v_2169 = v_709 ^ v_529;
assign v_2170 = v_710 ^ v_530;
assign v_2171 = v_711 ^ v_531;
assign v_2172 = v_712 ^ v_532;
assign v_2173 = v_713 ^ v_533;
assign v_2174 = v_714 ^ v_534;
assign v_2175 = v_715 ^ v_535;
assign v_2176 = v_716 ^ v_536;
assign v_2177 = v_717 ^ v_537;
assign v_2178 = v_718 ^ v_538;
assign v_2179 = v_719 ^ v_539;
assign v_2180 = v_720 ^ v_540;
assign v_2183 = v_721 ^ v_481;
assign v_2184 = v_722 ^ v_482;
assign v_2185 = v_723 ^ v_483;
assign v_2186 = v_724 ^ v_484;
assign v_2187 = v_725 ^ v_485;
assign v_2188 = v_726 ^ v_486;
assign v_2189 = v_727 ^ v_487;
assign v_2190 = v_728 ^ v_488;
assign v_2191 = v_729 ^ v_489;
assign v_2192 = v_730 ^ v_490;
assign v_2193 = v_731 ^ v_491;
assign v_2194 = v_732 ^ v_492;
assign v_2195 = v_733 ^ v_493;
assign v_2196 = v_734 ^ v_494;
assign v_2197 = v_735 ^ v_495;
assign v_2198 = v_736 ^ v_496;
assign v_2199 = v_737 ^ v_497;
assign v_2200 = v_738 ^ v_498;
assign v_2201 = v_739 ^ v_499;
assign v_2202 = v_740 ^ v_500;
assign v_2204 = v_741 ^ v_501;
assign v_2205 = v_742 ^ v_502;
assign v_2206 = v_743 ^ v_503;
assign v_2207 = v_744 ^ v_504;
assign v_2208 = v_745 ^ v_505;
assign v_2209 = v_746 ^ v_506;
assign v_2210 = v_747 ^ v_507;
assign v_2211 = v_748 ^ v_508;
assign v_2212 = v_749 ^ v_509;
assign v_2213 = v_750 ^ v_510;
assign v_2214 = v_751 ^ v_511;
assign v_2215 = v_752 ^ v_512;
assign v_2216 = v_753 ^ v_513;
assign v_2217 = v_754 ^ v_514;
assign v_2218 = v_755 ^ v_515;
assign v_2219 = v_756 ^ v_516;
assign v_2220 = v_757 ^ v_517;
assign v_2221 = v_758 ^ v_518;
assign v_2222 = v_759 ^ v_519;
assign v_2223 = v_760 ^ v_520;
assign v_2225 = v_761 ^ v_521;
assign v_2226 = v_762 ^ v_522;
assign v_2227 = v_763 ^ v_523;
assign v_2228 = v_764 ^ v_524;
assign v_2229 = v_765 ^ v_525;
assign v_2230 = v_766 ^ v_526;
assign v_2231 = v_767 ^ v_527;
assign v_2232 = v_768 ^ v_528;
assign v_2233 = v_769 ^ v_529;
assign v_2234 = v_770 ^ v_530;
assign v_2235 = v_771 ^ v_531;
assign v_2236 = v_772 ^ v_532;
assign v_2237 = v_773 ^ v_533;
assign v_2238 = v_774 ^ v_534;
assign v_2239 = v_775 ^ v_535;
assign v_2240 = v_776 ^ v_536;
assign v_2241 = v_777 ^ v_537;
assign v_2242 = v_778 ^ v_538;
assign v_2243 = v_779 ^ v_539;
assign v_2244 = v_780 ^ v_540;
assign v_2247 = v_781 ^ v_481;
assign v_2248 = v_782 ^ v_482;
assign v_2249 = v_783 ^ v_483;
assign v_2250 = v_784 ^ v_484;
assign v_2251 = v_785 ^ v_485;
assign v_2252 = v_786 ^ v_486;
assign v_2253 = v_787 ^ v_487;
assign v_2254 = v_788 ^ v_488;
assign v_2255 = v_789 ^ v_489;
assign v_2256 = v_790 ^ v_490;
assign v_2257 = v_791 ^ v_491;
assign v_2258 = v_792 ^ v_492;
assign v_2259 = v_793 ^ v_493;
assign v_2260 = v_794 ^ v_494;
assign v_2261 = v_795 ^ v_495;
assign v_2262 = v_796 ^ v_496;
assign v_2263 = v_797 ^ v_497;
assign v_2264 = v_798 ^ v_498;
assign v_2265 = v_799 ^ v_499;
assign v_2266 = v_800 ^ v_500;
assign v_2268 = v_801 ^ v_501;
assign v_2269 = v_802 ^ v_502;
assign v_2270 = v_803 ^ v_503;
assign v_2271 = v_804 ^ v_504;
assign v_2272 = v_805 ^ v_505;
assign v_2273 = v_806 ^ v_506;
assign v_2274 = v_807 ^ v_507;
assign v_2275 = v_808 ^ v_508;
assign v_2276 = v_809 ^ v_509;
assign v_2277 = v_810 ^ v_510;
assign v_2278 = v_811 ^ v_511;
assign v_2279 = v_812 ^ v_512;
assign v_2280 = v_813 ^ v_513;
assign v_2281 = v_814 ^ v_514;
assign v_2282 = v_815 ^ v_515;
assign v_2283 = v_816 ^ v_516;
assign v_2284 = v_817 ^ v_517;
assign v_2285 = v_818 ^ v_518;
assign v_2286 = v_819 ^ v_519;
assign v_2287 = v_820 ^ v_520;
assign v_2289 = v_821 ^ v_521;
assign v_2290 = v_822 ^ v_522;
assign v_2291 = v_823 ^ v_523;
assign v_2292 = v_824 ^ v_524;
assign v_2293 = v_825 ^ v_525;
assign v_2294 = v_826 ^ v_526;
assign v_2295 = v_827 ^ v_527;
assign v_2296 = v_828 ^ v_528;
assign v_2297 = v_829 ^ v_529;
assign v_2298 = v_830 ^ v_530;
assign v_2299 = v_831 ^ v_531;
assign v_2300 = v_832 ^ v_532;
assign v_2301 = v_833 ^ v_533;
assign v_2302 = v_834 ^ v_534;
assign v_2303 = v_835 ^ v_535;
assign v_2304 = v_836 ^ v_536;
assign v_2305 = v_837 ^ v_537;
assign v_2306 = v_838 ^ v_538;
assign v_2307 = v_839 ^ v_539;
assign v_2308 = v_840 ^ v_540;
assign v_2311 = v_841 ^ v_481;
assign v_2312 = v_842 ^ v_482;
assign v_2313 = v_843 ^ v_483;
assign v_2314 = v_844 ^ v_484;
assign v_2315 = v_845 ^ v_485;
assign v_2316 = v_846 ^ v_486;
assign v_2317 = v_847 ^ v_487;
assign v_2318 = v_848 ^ v_488;
assign v_2319 = v_849 ^ v_489;
assign v_2320 = v_850 ^ v_490;
assign v_2321 = v_851 ^ v_491;
assign v_2322 = v_852 ^ v_492;
assign v_2323 = v_853 ^ v_493;
assign v_2324 = v_854 ^ v_494;
assign v_2325 = v_855 ^ v_495;
assign v_2326 = v_856 ^ v_496;
assign v_2327 = v_857 ^ v_497;
assign v_2328 = v_858 ^ v_498;
assign v_2329 = v_859 ^ v_499;
assign v_2330 = v_860 ^ v_500;
assign v_2332 = v_861 ^ v_501;
assign v_2333 = v_862 ^ v_502;
assign v_2334 = v_863 ^ v_503;
assign v_2335 = v_864 ^ v_504;
assign v_2336 = v_865 ^ v_505;
assign v_2337 = v_866 ^ v_506;
assign v_2338 = v_867 ^ v_507;
assign v_2339 = v_868 ^ v_508;
assign v_2340 = v_869 ^ v_509;
assign v_2341 = v_870 ^ v_510;
assign v_2342 = v_871 ^ v_511;
assign v_2343 = v_872 ^ v_512;
assign v_2344 = v_873 ^ v_513;
assign v_2345 = v_874 ^ v_514;
assign v_2346 = v_875 ^ v_515;
assign v_2347 = v_876 ^ v_516;
assign v_2348 = v_877 ^ v_517;
assign v_2349 = v_878 ^ v_518;
assign v_2350 = v_879 ^ v_519;
assign v_2351 = v_880 ^ v_520;
assign v_2353 = v_881 ^ v_521;
assign v_2354 = v_882 ^ v_522;
assign v_2355 = v_883 ^ v_523;
assign v_2356 = v_884 ^ v_524;
assign v_2357 = v_885 ^ v_525;
assign v_2358 = v_886 ^ v_526;
assign v_2359 = v_887 ^ v_527;
assign v_2360 = v_888 ^ v_528;
assign v_2361 = v_889 ^ v_529;
assign v_2362 = v_890 ^ v_530;
assign v_2363 = v_891 ^ v_531;
assign v_2364 = v_892 ^ v_532;
assign v_2365 = v_893 ^ v_533;
assign v_2366 = v_894 ^ v_534;
assign v_2367 = v_895 ^ v_535;
assign v_2368 = v_896 ^ v_536;
assign v_2369 = v_897 ^ v_537;
assign v_2370 = v_898 ^ v_538;
assign v_2371 = v_899 ^ v_539;
assign v_2372 = v_900 ^ v_540;
assign v_2375 = v_901 ^ v_481;
assign v_2376 = v_902 ^ v_482;
assign v_2377 = v_903 ^ v_483;
assign v_2378 = v_904 ^ v_484;
assign v_2379 = v_905 ^ v_485;
assign v_2380 = v_906 ^ v_486;
assign v_2381 = v_907 ^ v_487;
assign v_2382 = v_908 ^ v_488;
assign v_2383 = v_909 ^ v_489;
assign v_2384 = v_910 ^ v_490;
assign v_2385 = v_911 ^ v_491;
assign v_2386 = v_912 ^ v_492;
assign v_2387 = v_913 ^ v_493;
assign v_2388 = v_914 ^ v_494;
assign v_2389 = v_915 ^ v_495;
assign v_2390 = v_916 ^ v_496;
assign v_2391 = v_917 ^ v_497;
assign v_2392 = v_918 ^ v_498;
assign v_2393 = v_919 ^ v_499;
assign v_2394 = v_920 ^ v_500;
assign v_2396 = v_921 ^ v_501;
assign v_2397 = v_922 ^ v_502;
assign v_2398 = v_923 ^ v_503;
assign v_2399 = v_924 ^ v_504;
assign v_2400 = v_925 ^ v_505;
assign v_2401 = v_926 ^ v_506;
assign v_2402 = v_927 ^ v_507;
assign v_2403 = v_928 ^ v_508;
assign v_2404 = v_929 ^ v_509;
assign v_2405 = v_930 ^ v_510;
assign v_2406 = v_931 ^ v_511;
assign v_2407 = v_932 ^ v_512;
assign v_2408 = v_933 ^ v_513;
assign v_2409 = v_934 ^ v_514;
assign v_2410 = v_935 ^ v_515;
assign v_2411 = v_936 ^ v_516;
assign v_2412 = v_937 ^ v_517;
assign v_2413 = v_938 ^ v_518;
assign v_2414 = v_939 ^ v_519;
assign v_2415 = v_940 ^ v_520;
assign v_2417 = v_941 ^ v_521;
assign v_2418 = v_942 ^ v_522;
assign v_2419 = v_943 ^ v_523;
assign v_2420 = v_944 ^ v_524;
assign v_2421 = v_945 ^ v_525;
assign v_2422 = v_946 ^ v_526;
assign v_2423 = v_947 ^ v_527;
assign v_2424 = v_948 ^ v_528;
assign v_2425 = v_949 ^ v_529;
assign v_2426 = v_950 ^ v_530;
assign v_2427 = v_951 ^ v_531;
assign v_2428 = v_952 ^ v_532;
assign v_2429 = v_953 ^ v_533;
assign v_2430 = v_954 ^ v_534;
assign v_2431 = v_955 ^ v_535;
assign v_2432 = v_956 ^ v_536;
assign v_2433 = v_957 ^ v_537;
assign v_2434 = v_958 ^ v_538;
assign v_2435 = v_959 ^ v_539;
assign v_2436 = v_960 ^ v_540;
assign v_2439 = v_961 ^ v_481;
assign v_2440 = v_962 ^ v_482;
assign v_2441 = v_963 ^ v_483;
assign v_2442 = v_964 ^ v_484;
assign v_2443 = v_965 ^ v_485;
assign v_2444 = v_966 ^ v_486;
assign v_2445 = v_967 ^ v_487;
assign v_2446 = v_968 ^ v_488;
assign v_2447 = v_969 ^ v_489;
assign v_2448 = v_970 ^ v_490;
assign v_2449 = v_971 ^ v_491;
assign v_2450 = v_972 ^ v_492;
assign v_2451 = v_973 ^ v_493;
assign v_2452 = v_974 ^ v_494;
assign v_2453 = v_975 ^ v_495;
assign v_2454 = v_976 ^ v_496;
assign v_2455 = v_977 ^ v_497;
assign v_2456 = v_978 ^ v_498;
assign v_2457 = v_979 ^ v_499;
assign v_2458 = v_980 ^ v_500;
assign v_2460 = v_981 ^ v_501;
assign v_2461 = v_982 ^ v_502;
assign v_2462 = v_983 ^ v_503;
assign v_2463 = v_984 ^ v_504;
assign v_2464 = v_985 ^ v_505;
assign v_2465 = v_986 ^ v_506;
assign v_2466 = v_987 ^ v_507;
assign v_2467 = v_988 ^ v_508;
assign v_2468 = v_989 ^ v_509;
assign v_2469 = v_990 ^ v_510;
assign v_2470 = v_991 ^ v_511;
assign v_2471 = v_992 ^ v_512;
assign v_2472 = v_993 ^ v_513;
assign v_2473 = v_994 ^ v_514;
assign v_2474 = v_995 ^ v_515;
assign v_2475 = v_996 ^ v_516;
assign v_2476 = v_997 ^ v_517;
assign v_2477 = v_998 ^ v_518;
assign v_2478 = v_999 ^ v_519;
assign v_2479 = v_1000 ^ v_520;
assign v_2481 = v_1001 ^ v_521;
assign v_2482 = v_1002 ^ v_522;
assign v_2483 = v_1003 ^ v_523;
assign v_2484 = v_1004 ^ v_524;
assign v_2485 = v_1005 ^ v_525;
assign v_2486 = v_1006 ^ v_526;
assign v_2487 = v_1007 ^ v_527;
assign v_2488 = v_1008 ^ v_528;
assign v_2489 = v_1009 ^ v_529;
assign v_2490 = v_1010 ^ v_530;
assign v_2491 = v_1011 ^ v_531;
assign v_2492 = v_1012 ^ v_532;
assign v_2493 = v_1013 ^ v_533;
assign v_2494 = v_1014 ^ v_534;
assign v_2495 = v_1015 ^ v_535;
assign v_2496 = v_1016 ^ v_536;
assign v_2497 = v_1017 ^ v_537;
assign v_2498 = v_1018 ^ v_538;
assign v_2499 = v_1019 ^ v_539;
assign v_2500 = v_1020 ^ v_540;
assign x_1 = v_2504 | ~v_1537;
assign o_1 = x_1;
endmodule
