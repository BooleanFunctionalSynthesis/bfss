// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module bobsynthetic_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37, i_38, i_39, i_40, i_41, i_42, i_43, i_44, i_45, i_46, i_47, i_48, i_49, i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input i_33;
input i_34;
input i_35;
input i_36;
input i_37;
input i_38;
input i_39;
input i_40;
input i_41;
input i_42;
input i_43;
input i_44;
input i_45;
input i_46;
input i_47;
input i_48;
input i_49;
input i_50;
input i_51;
input i_52;
input i_53;
input i_54;
input i_55;
input i_56;
input i_57;
input i_58;
input i_59;
input i_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_2770;
wire n_2771;
wire n_2772;
wire n_2773;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_2790;
wire n_2791;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2796;
wire n_2797;
wire n_2798;
wire n_2799;
wire n_2800;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2808;
wire n_2809;
wire n_2810;
wire n_2811;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2816;
wire n_2817;
wire n_2818;
wire n_2819;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2827;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2832;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2837;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2845;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_2850;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2875;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_2879;
wire n_2880;
wire n_2881;
wire n_2882;
wire n_2883;
wire n_2884;
wire n_2885;
wire n_2886;
wire n_2887;
wire n_2888;
wire n_2889;
wire n_2890;
wire n_2891;
wire n_2892;
wire n_2893;
wire n_2894;
wire n_2895;
wire n_2896;
wire n_2897;
wire n_2898;
wire n_2899;
wire n_2900;
wire n_2901;
wire n_2902;
wire n_2903;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2908;
wire n_2909;
wire n_2910;
wire n_2911;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2923;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2928;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2944;
wire n_2945;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_3069;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_3400;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_3410;
wire n_3411;
wire n_3412;
wire n_3413;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_3428;
wire n_3429;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4038;
wire n_4039;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4125;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire n_4159;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_4178;
wire n_4179;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_4187;
wire n_4188;
wire n_4189;
wire n_4190;
wire n_4191;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_4200;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4216;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_4240;
wire n_4241;
wire n_4242;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire n_4285;
wire n_4286;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4348;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_4790;
wire n_4791;
wire n_4792;
wire n_4793;
wire n_4794;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4803;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
assign n_1 =  x_61 &  x_63;
assign n_2 = ~x_61 & ~x_119;
assign n_3 =  x_61 &  x_119;
assign n_4 = ~n_2 & ~n_3;
assign n_5 = ~x_63 & ~n_4;
assign n_6 = ~n_1 & ~n_5;
assign n_7 =  x_117 & ~n_6;
assign n_8 = ~x_63 &  x_119;
assign n_9 = ~n_2 & ~n_8;
assign n_10 = ~x_117 & ~n_9;
assign n_11 = ~n_7 & ~n_10;
assign n_12 =  x_65 & ~n_11;
assign n_13 = ~x_61 &  x_63;
assign n_14 =  x_119 &  n_13;
assign n_15 =  x_61 & ~x_119;
assign n_16 = ~x_63 &  n_15;
assign n_17 = ~n_14 & ~n_16;
assign n_18 =  x_117 & ~n_17;
assign n_19 = ~x_117 &  n_1;
assign n_20 = ~n_18 & ~n_19;
assign n_21 = ~n_10 &  n_20;
assign n_22 = ~n_7 &  n_21;
assign n_23 = ~n_10 & ~n_22;
assign n_24 = ~x_65 & ~n_23;
assign n_25 = ~n_12 & ~n_24;
assign n_26 =  x_115 & ~n_25;
assign n_27 =  x_65 & ~n_20;
assign n_28 = ~x_65 &  n_7;
assign n_29 = ~n_27 & ~n_28;
assign n_30 = ~n_24 &  n_29;
assign n_31 = ~n_12 &  n_30;
assign n_32 = ~n_24 & ~n_31;
assign n_33 = ~x_115 & ~n_32;
assign n_34 =  x_115 & ~n_29;
assign n_35 = ~x_115 &  n_12;
assign n_36 = ~n_34 & ~n_35;
assign n_37 = ~n_33 &  n_36;
assign n_38 = ~n_26 &  n_37;
assign n_39 =  x_67 & ~n_37;
assign n_40 = ~n_38 & ~n_39;
assign n_41 = ~n_26 & ~n_33;
assign n_42 =  x_67 & ~n_41;
assign n_43 = ~n_33 & ~n_38;
assign n_44 = ~x_67 & ~n_43;
assign n_45 = ~n_42 & ~n_44;
assign n_46 =  x_113 & ~n_45;
assign n_47 = ~x_67 & ~n_26;
assign n_48 =  x_67 &  n_36;
assign n_49 = ~n_47 & ~n_48;
assign n_50 = ~n_44 & ~n_49;
assign n_51 = ~n_42 &  n_50;
assign n_52 = ~n_44 & ~n_51;
assign n_53 = ~x_113 & ~n_52;
assign n_54 = ~n_46 & ~n_53;
assign n_55 =  x_69 & ~n_54;
assign n_56 =  x_113 & ~n_49;
assign n_57 = ~x_113 & ~n_42;
assign n_58 = ~n_56 & ~n_57;
assign n_59 = ~n_53 & ~n_58;
assign n_60 = ~n_46 &  n_59;
assign n_61 = ~n_53 & ~n_60;
assign n_62 = ~x_69 & ~n_61;
assign n_63 = ~n_55 & ~n_62;
assign n_64 =  x_111 & ~n_63;
assign n_65 =  x_69 & ~n_58;
assign n_66 = ~x_69 & ~n_46;
assign n_67 = ~n_65 & ~n_66;
assign n_68 = ~n_62 & ~n_67;
assign n_69 = ~n_55 &  n_68;
assign n_70 = ~n_62 & ~n_69;
assign n_71 = ~x_111 & ~n_70;
assign n_72 = ~n_64 & ~n_71;
assign n_73 =  x_71 & ~n_72;
assign n_74 =  x_111 & ~n_67;
assign n_75 = ~x_111 & ~n_55;
assign n_76 = ~n_74 & ~n_75;
assign n_77 = ~n_71 & ~n_76;
assign n_78 = ~n_64 &  n_77;
assign n_79 = ~n_71 & ~n_78;
assign n_80 = ~x_71 & ~n_79;
assign n_81 = ~n_73 & ~n_80;
assign n_82 =  x_109 & ~n_81;
assign n_83 =  x_71 & ~n_76;
assign n_84 = ~x_71 & ~n_64;
assign n_85 = ~n_83 & ~n_84;
assign n_86 = ~n_80 & ~n_85;
assign n_87 = ~n_73 &  n_86;
assign n_88 = ~n_80 & ~n_87;
assign n_89 = ~x_109 & ~n_88;
assign n_90 = ~n_82 & ~n_89;
assign n_91 =  x_73 & ~n_90;
assign n_92 =  x_109 & ~n_85;
assign n_93 = ~x_109 & ~n_73;
assign n_94 = ~n_92 & ~n_93;
assign n_95 = ~n_89 & ~n_94;
assign n_96 = ~n_82 &  n_95;
assign n_97 = ~n_89 & ~n_96;
assign n_98 = ~x_73 & ~n_97;
assign n_99 = ~n_91 & ~n_98;
assign n_100 =  x_107 & ~n_99;
assign n_101 =  x_73 & ~n_94;
assign n_102 = ~x_73 & ~n_82;
assign n_103 = ~n_101 & ~n_102;
assign n_104 = ~n_98 & ~n_103;
assign n_105 = ~n_91 &  n_104;
assign n_106 = ~n_98 & ~n_105;
assign n_107 = ~x_107 & ~n_106;
assign n_108 = ~n_100 & ~n_107;
assign n_109 =  x_75 & ~n_108;
assign n_110 =  x_107 & ~n_103;
assign n_111 = ~x_107 & ~n_91;
assign n_112 = ~n_110 & ~n_111;
assign n_113 = ~n_107 & ~n_112;
assign n_114 = ~n_100 &  n_113;
assign n_115 = ~n_107 & ~n_114;
assign n_116 = ~x_75 & ~n_115;
assign n_117 = ~n_109 & ~n_116;
assign n_118 =  x_105 & ~n_117;
assign n_119 =  x_75 & ~n_112;
assign n_120 = ~x_75 & ~n_100;
assign n_121 = ~n_119 & ~n_120;
assign n_122 = ~n_116 & ~n_121;
assign n_123 = ~n_109 &  n_122;
assign n_124 = ~n_116 & ~n_123;
assign n_125 = ~x_105 & ~n_124;
assign n_126 = ~n_118 & ~n_125;
assign n_127 =  x_77 & ~n_126;
assign n_128 =  x_105 & ~n_121;
assign n_129 = ~x_105 & ~n_109;
assign n_130 = ~n_128 & ~n_129;
assign n_131 = ~n_125 & ~n_130;
assign n_132 = ~n_118 &  n_131;
assign n_133 = ~n_125 & ~n_132;
assign n_134 = ~x_77 & ~n_133;
assign n_135 = ~n_127 & ~n_134;
assign n_136 =  x_103 & ~n_135;
assign n_137 =  x_77 & ~n_130;
assign n_138 = ~x_77 & ~n_118;
assign n_139 = ~n_137 & ~n_138;
assign n_140 = ~n_134 & ~n_139;
assign n_141 = ~n_127 &  n_140;
assign n_142 = ~n_134 & ~n_141;
assign n_143 = ~x_103 & ~n_142;
assign n_144 = ~n_136 & ~n_143;
assign n_145 =  x_79 & ~n_144;
assign n_146 =  x_103 & ~n_139;
assign n_147 = ~x_103 & ~n_127;
assign n_148 = ~n_146 & ~n_147;
assign n_149 = ~n_143 & ~n_148;
assign n_150 = ~n_136 &  n_149;
assign n_151 = ~n_143 & ~n_150;
assign n_152 = ~x_79 & ~n_151;
assign n_153 = ~n_145 & ~n_152;
assign n_154 =  x_101 & ~n_153;
assign n_155 =  x_79 & ~n_148;
assign n_156 = ~x_79 & ~n_136;
assign n_157 = ~n_155 & ~n_156;
assign n_158 = ~n_152 & ~n_157;
assign n_159 = ~n_145 &  n_158;
assign n_160 = ~n_152 & ~n_159;
assign n_161 = ~x_101 & ~n_160;
assign n_162 = ~n_154 & ~n_161;
assign n_163 =  x_81 & ~n_162;
assign n_164 =  x_101 & ~n_157;
assign n_165 = ~x_101 & ~n_145;
assign n_166 = ~n_164 & ~n_165;
assign n_167 = ~n_161 & ~n_166;
assign n_168 = ~n_154 &  n_167;
assign n_169 = ~n_161 & ~n_168;
assign n_170 = ~x_81 & ~n_169;
assign n_171 = ~n_163 & ~n_170;
assign n_172 =  x_99 & ~n_171;
assign n_173 =  x_81 & ~n_166;
assign n_174 = ~x_81 & ~n_154;
assign n_175 = ~n_173 & ~n_174;
assign n_176 = ~n_170 & ~n_175;
assign n_177 = ~n_163 &  n_176;
assign n_178 = ~n_170 & ~n_177;
assign n_179 = ~x_99 & ~n_178;
assign n_180 = ~n_172 & ~n_179;
assign n_181 =  x_83 & ~n_180;
assign n_182 =  x_99 & ~n_175;
assign n_183 = ~x_99 & ~n_163;
assign n_184 = ~n_182 & ~n_183;
assign n_185 = ~n_179 & ~n_184;
assign n_186 = ~n_172 &  n_185;
assign n_187 = ~n_179 & ~n_186;
assign n_188 = ~x_83 & ~n_187;
assign n_189 = ~n_181 & ~n_188;
assign n_190 =  x_97 & ~n_189;
assign n_191 =  x_83 & ~n_184;
assign n_192 = ~x_83 & ~n_172;
assign n_193 = ~n_191 & ~n_192;
assign n_194 = ~n_188 & ~n_193;
assign n_195 = ~n_181 &  n_194;
assign n_196 = ~n_188 & ~n_195;
assign n_197 = ~x_97 & ~n_196;
assign n_198 = ~n_190 & ~n_197;
assign n_199 =  x_85 & ~n_198;
assign n_200 =  x_97 & ~n_193;
assign n_201 = ~x_97 & ~n_181;
assign n_202 = ~n_200 & ~n_201;
assign n_203 = ~n_197 & ~n_202;
assign n_204 = ~n_190 &  n_203;
assign n_205 = ~n_197 & ~n_204;
assign n_206 = ~x_85 & ~n_205;
assign n_207 = ~n_199 & ~n_206;
assign n_208 =  x_95 & ~n_207;
assign n_209 =  x_85 & ~n_202;
assign n_210 = ~x_85 & ~n_190;
assign n_211 = ~n_209 & ~n_210;
assign n_212 = ~n_206 & ~n_211;
assign n_213 = ~n_199 &  n_212;
assign n_214 = ~n_206 & ~n_213;
assign n_215 = ~x_95 & ~n_214;
assign n_216 = ~n_208 & ~n_215;
assign n_217 =  x_87 & ~n_216;
assign n_218 =  x_95 & ~n_211;
assign n_219 = ~x_95 & ~n_199;
assign n_220 = ~n_218 & ~n_219;
assign n_221 = ~n_215 & ~n_220;
assign n_222 = ~n_208 &  n_221;
assign n_223 = ~n_215 & ~n_222;
assign n_224 = ~x_87 & ~n_223;
assign n_225 = ~n_217 & ~n_224;
assign n_226 =  x_93 & ~n_225;
assign n_227 =  x_87 & ~n_220;
assign n_228 = ~x_87 & ~n_208;
assign n_229 = ~n_227 & ~n_228;
assign n_230 = ~n_224 & ~n_229;
assign n_231 = ~n_217 &  n_230;
assign n_232 = ~n_224 & ~n_231;
assign n_233 = ~x_93 & ~n_232;
assign n_234 = ~n_226 & ~n_233;
assign n_235 =  x_89 & ~n_234;
assign n_236 =  x_93 & ~n_229;
assign n_237 = ~x_93 & ~n_217;
assign n_238 = ~n_236 & ~n_237;
assign n_239 = ~n_233 & ~n_238;
assign n_240 = ~n_226 &  n_239;
assign n_241 = ~n_233 & ~n_240;
assign n_242 = ~x_89 & ~n_241;
assign n_243 = ~n_235 & ~n_242;
assign n_244 =  x_91 & ~n_243;
assign n_245 =  x_89 & ~n_238;
assign n_246 = ~x_89 & ~n_226;
assign n_247 = ~n_245 & ~n_246;
assign n_248 = ~n_242 & ~n_247;
assign n_249 = ~n_235 &  n_248;
assign n_250 = ~n_242 & ~n_249;
assign n_251 = ~x_91 & ~n_250;
assign n_252 = ~n_244 & ~n_251;
assign n_253 =  x_90 & ~n_252;
assign n_254 =  x_91 & ~n_247;
assign n_255 = ~x_91 & ~n_235;
assign n_256 = ~n_254 & ~n_255;
assign n_257 = ~n_251 & ~n_256;
assign n_258 = ~n_244 &  n_257;
assign n_259 = ~n_251 & ~n_258;
assign n_260 = ~x_90 & ~n_259;
assign n_261 = ~n_253 & ~n_260;
assign n_262 =  x_92 & ~n_261;
assign n_263 =  x_90 & ~n_256;
assign n_264 = ~x_90 & ~n_244;
assign n_265 = ~n_263 & ~n_264;
assign n_266 = ~n_260 & ~n_265;
assign n_267 = ~n_253 &  n_266;
assign n_268 = ~n_260 & ~n_267;
assign n_269 = ~x_92 & ~n_268;
assign n_270 = ~n_262 & ~n_269;
assign n_271 =  x_88 & ~n_270;
assign n_272 =  x_92 & ~n_265;
assign n_273 = ~x_92 & ~n_253;
assign n_274 = ~n_272 & ~n_273;
assign n_275 = ~n_269 & ~n_274;
assign n_276 = ~n_262 &  n_275;
assign n_277 = ~n_269 & ~n_276;
assign n_278 = ~x_88 & ~n_277;
assign n_279 = ~n_271 & ~n_278;
assign n_280 =  x_94 & ~n_279;
assign n_281 =  x_88 & ~n_274;
assign n_282 = ~x_88 & ~n_262;
assign n_283 = ~n_281 & ~n_282;
assign n_284 = ~n_278 & ~n_283;
assign n_285 = ~n_271 &  n_284;
assign n_286 = ~n_278 & ~n_285;
assign n_287 = ~x_94 & ~n_286;
assign n_288 = ~n_280 & ~n_287;
assign n_289 =  x_86 & ~n_288;
assign n_290 =  x_94 & ~n_283;
assign n_291 = ~x_94 & ~n_271;
assign n_292 = ~n_290 & ~n_291;
assign n_293 = ~n_287 & ~n_292;
assign n_294 = ~n_280 &  n_293;
assign n_295 = ~n_287 & ~n_294;
assign n_296 = ~x_86 & ~n_295;
assign n_297 = ~n_289 & ~n_296;
assign n_298 =  x_96 & ~n_297;
assign n_299 =  x_86 & ~n_292;
assign n_300 = ~x_86 & ~n_280;
assign n_301 = ~n_299 & ~n_300;
assign n_302 = ~n_296 & ~n_301;
assign n_303 = ~n_289 &  n_302;
assign n_304 = ~n_296 & ~n_303;
assign n_305 = ~x_96 & ~n_304;
assign n_306 = ~n_298 & ~n_305;
assign n_307 =  x_84 & ~n_306;
assign n_308 =  x_96 & ~n_301;
assign n_309 = ~x_96 & ~n_289;
assign n_310 = ~n_308 & ~n_309;
assign n_311 = ~n_305 & ~n_310;
assign n_312 = ~n_298 &  n_311;
assign n_313 = ~n_305 & ~n_312;
assign n_314 = ~x_84 & ~n_313;
assign n_315 = ~n_307 & ~n_314;
assign n_316 =  x_98 & ~n_315;
assign n_317 =  x_84 & ~n_310;
assign n_318 = ~x_84 & ~n_298;
assign n_319 = ~n_317 & ~n_318;
assign n_320 = ~n_314 & ~n_319;
assign n_321 = ~n_307 &  n_320;
assign n_322 = ~n_314 & ~n_321;
assign n_323 = ~x_98 & ~n_322;
assign n_324 = ~n_316 & ~n_323;
assign n_325 =  x_82 & ~n_324;
assign n_326 =  x_98 & ~n_319;
assign n_327 = ~x_98 & ~n_307;
assign n_328 = ~n_326 & ~n_327;
assign n_329 = ~n_323 & ~n_328;
assign n_330 = ~n_316 &  n_329;
assign n_331 = ~n_323 & ~n_330;
assign n_332 = ~x_82 & ~n_331;
assign n_333 = ~n_325 & ~n_332;
assign n_334 =  x_100 & ~n_333;
assign n_335 =  x_82 & ~n_328;
assign n_336 = ~x_82 & ~n_316;
assign n_337 = ~n_335 & ~n_336;
assign n_338 = ~n_332 & ~n_337;
assign n_339 = ~n_325 &  n_338;
assign n_340 = ~n_332 & ~n_339;
assign n_341 = ~x_100 & ~n_340;
assign n_342 = ~n_334 & ~n_341;
assign n_343 =  x_80 & ~n_342;
assign n_344 =  x_100 & ~n_337;
assign n_345 = ~x_100 & ~n_325;
assign n_346 = ~n_344 & ~n_345;
assign n_347 = ~n_341 & ~n_346;
assign n_348 = ~n_334 &  n_347;
assign n_349 = ~n_341 & ~n_348;
assign n_350 = ~x_80 & ~n_349;
assign n_351 = ~n_343 & ~n_350;
assign n_352 =  x_102 & ~n_351;
assign n_353 =  x_80 & ~n_346;
assign n_354 = ~x_80 & ~n_334;
assign n_355 = ~n_353 & ~n_354;
assign n_356 = ~n_350 & ~n_355;
assign n_357 = ~n_343 &  n_356;
assign n_358 = ~n_350 & ~n_357;
assign n_359 = ~x_102 & ~n_358;
assign n_360 = ~n_352 & ~n_359;
assign n_361 =  x_78 & ~n_360;
assign n_362 =  x_102 & ~n_355;
assign n_363 = ~x_102 & ~n_343;
assign n_364 = ~n_362 & ~n_363;
assign n_365 = ~n_359 & ~n_364;
assign n_366 = ~n_352 &  n_365;
assign n_367 = ~n_359 & ~n_366;
assign n_368 = ~x_78 & ~n_367;
assign n_369 = ~n_361 & ~n_368;
assign n_370 =  x_104 & ~n_369;
assign n_371 =  x_78 & ~n_364;
assign n_372 = ~x_78 & ~n_352;
assign n_373 = ~n_371 & ~n_372;
assign n_374 = ~n_368 & ~n_373;
assign n_375 = ~n_361 &  n_374;
assign n_376 = ~n_368 & ~n_375;
assign n_377 = ~x_104 & ~n_376;
assign n_378 = ~n_370 & ~n_377;
assign n_379 =  x_76 & ~n_378;
assign n_380 =  x_104 & ~n_373;
assign n_381 = ~x_104 & ~n_361;
assign n_382 = ~n_380 & ~n_381;
assign n_383 = ~n_377 & ~n_382;
assign n_384 = ~n_370 &  n_383;
assign n_385 = ~n_377 & ~n_384;
assign n_386 = ~x_76 & ~n_385;
assign n_387 = ~n_379 & ~n_386;
assign n_388 =  x_106 & ~n_387;
assign n_389 =  x_76 & ~n_382;
assign n_390 = ~x_76 & ~n_370;
assign n_391 = ~n_389 & ~n_390;
assign n_392 = ~n_386 & ~n_391;
assign n_393 = ~n_379 &  n_392;
assign n_394 = ~n_386 & ~n_393;
assign n_395 = ~x_106 & ~n_394;
assign n_396 = ~n_388 & ~n_395;
assign n_397 =  x_74 & ~n_396;
assign n_398 =  x_106 & ~n_391;
assign n_399 = ~x_106 & ~n_379;
assign n_400 = ~n_398 & ~n_399;
assign n_401 = ~n_395 & ~n_400;
assign n_402 = ~n_388 &  n_401;
assign n_403 = ~n_395 & ~n_402;
assign n_404 = ~x_74 & ~n_403;
assign n_405 = ~n_397 & ~n_404;
assign n_406 =  x_108 & ~n_405;
assign n_407 =  x_74 & ~n_400;
assign n_408 = ~x_74 & ~n_388;
assign n_409 = ~n_407 & ~n_408;
assign n_410 = ~n_404 & ~n_409;
assign n_411 = ~n_397 &  n_410;
assign n_412 = ~n_404 & ~n_411;
assign n_413 = ~x_108 & ~n_412;
assign n_414 = ~n_406 & ~n_413;
assign n_415 =  x_72 & ~n_414;
assign n_416 =  x_108 & ~n_409;
assign n_417 = ~x_108 & ~n_397;
assign n_418 = ~n_416 & ~n_417;
assign n_419 = ~n_413 & ~n_418;
assign n_420 = ~n_406 &  n_419;
assign n_421 = ~n_413 & ~n_420;
assign n_422 = ~x_72 & ~n_421;
assign n_423 = ~n_415 & ~n_422;
assign n_424 =  x_110 & ~n_423;
assign n_425 =  x_72 & ~n_418;
assign n_426 = ~x_72 & ~n_406;
assign n_427 = ~n_425 & ~n_426;
assign n_428 = ~n_422 & ~n_427;
assign n_429 = ~n_415 &  n_428;
assign n_430 = ~n_422 & ~n_429;
assign n_431 = ~x_110 & ~n_430;
assign n_432 = ~n_424 & ~n_431;
assign n_433 =  x_70 & ~n_432;
assign n_434 =  x_110 & ~n_427;
assign n_435 = ~x_110 & ~n_415;
assign n_436 = ~n_434 & ~n_435;
assign n_437 = ~n_431 & ~n_436;
assign n_438 = ~n_424 &  n_437;
assign n_439 = ~n_431 & ~n_438;
assign n_440 = ~x_70 & ~n_439;
assign n_441 = ~n_433 & ~n_440;
assign n_442 =  x_112 & ~n_441;
assign n_443 =  x_70 & ~n_436;
assign n_444 = ~x_70 & ~n_424;
assign n_445 = ~n_443 & ~n_444;
assign n_446 = ~n_440 & ~n_445;
assign n_447 = ~n_433 &  n_446;
assign n_448 = ~n_440 & ~n_447;
assign n_449 = ~x_112 & ~n_448;
assign n_450 = ~n_442 & ~n_449;
assign n_451 =  x_68 & ~n_450;
assign n_452 =  x_112 & ~n_445;
assign n_453 = ~x_112 & ~n_433;
assign n_454 = ~n_452 & ~n_453;
assign n_455 = ~n_449 & ~n_454;
assign n_456 = ~n_442 &  n_455;
assign n_457 = ~n_449 & ~n_456;
assign n_458 = ~x_68 & ~n_457;
assign n_459 = ~n_451 & ~n_458;
assign n_460 =  x_114 & ~n_459;
assign n_461 =  x_68 & ~n_454;
assign n_462 = ~x_68 & ~n_442;
assign n_463 = ~n_461 & ~n_462;
assign n_464 = ~n_458 & ~n_463;
assign n_465 = ~n_451 &  n_464;
assign n_466 = ~n_458 & ~n_465;
assign n_467 = ~x_114 & ~n_466;
assign n_468 = ~n_460 & ~n_467;
assign n_469 =  x_66 & ~n_468;
assign n_470 =  x_114 & ~n_463;
assign n_471 = ~x_114 & ~n_451;
assign n_472 = ~n_470 & ~n_471;
assign n_473 = ~n_467 & ~n_472;
assign n_474 = ~n_460 &  n_473;
assign n_475 = ~n_467 & ~n_474;
assign n_476 = ~x_66 & ~n_475;
assign n_477 = ~n_469 & ~n_476;
assign n_478 =  x_116 & ~n_477;
assign n_479 =  x_66 & ~n_472;
assign n_480 = ~x_66 & ~n_460;
assign n_481 = ~n_479 & ~n_480;
assign n_482 = ~n_476 & ~n_481;
assign n_483 = ~n_469 &  n_482;
assign n_484 = ~n_476 & ~n_483;
assign n_485 = ~x_116 & ~n_484;
assign n_486 =  x_116 & ~n_481;
assign n_487 = ~x_116 & ~n_469;
assign n_488 = ~n_486 & ~n_487;
assign n_489 = ~n_485 & ~n_488;
assign n_490 = ~n_478 &  n_489;
assign n_491 =  x_64 & ~n_489;
assign n_492 = ~n_490 & ~n_491;
assign n_493 =  x_69 & ~n_59;
assign n_494 = ~n_60 & ~n_493;
assign n_495 =  x_66 & ~n_473;
assign n_496 = ~n_474 & ~n_495;
assign n_497 =  x_71 & ~n_77;
assign n_498 = ~n_78 & ~n_497;
assign n_499 =  x_68 & ~n_455;
assign n_500 = ~n_456 & ~n_499;
assign n_501 =  x_73 & ~n_95;
assign n_502 = ~n_96 & ~n_501;
assign n_503 =  x_70 & ~n_437;
assign n_504 = ~n_438 & ~n_503;
assign n_505 =  x_75 & ~n_113;
assign n_506 = ~n_114 & ~n_505;
assign n_507 =  x_72 & ~n_419;
assign n_508 = ~n_420 & ~n_507;
assign n_509 =  x_77 & ~n_131;
assign n_510 = ~n_132 & ~n_509;
assign n_511 =  x_74 & ~n_401;
assign n_512 = ~n_402 & ~n_511;
assign n_513 =  x_79 & ~n_149;
assign n_514 = ~n_150 & ~n_513;
assign n_515 =  x_76 & ~n_383;
assign n_516 = ~n_384 & ~n_515;
assign n_517 =  x_81 & ~n_167;
assign n_518 = ~n_168 & ~n_517;
assign n_519 =  x_78 & ~n_365;
assign n_520 = ~n_366 & ~n_519;
assign n_521 =  x_83 & ~n_185;
assign n_522 = ~n_186 & ~n_521;
assign n_523 =  x_80 & ~n_347;
assign n_524 = ~n_348 & ~n_523;
assign n_525 =  x_85 & ~n_203;
assign n_526 = ~n_204 & ~n_525;
assign n_527 =  x_82 & ~n_329;
assign n_528 = ~n_330 & ~n_527;
assign n_529 =  x_87 & ~n_221;
assign n_530 = ~n_222 & ~n_529;
assign n_531 =  x_84 & ~n_311;
assign n_532 = ~n_312 & ~n_531;
assign n_533 =  x_89 & ~n_239;
assign n_534 = ~n_240 & ~n_533;
assign n_535 =  x_86 & ~n_293;
assign n_536 = ~n_294 & ~n_535;
assign n_537 =  x_90 & ~n_257;
assign n_538 = ~n_258 & ~n_537;
assign n_539 =  x_88 & ~n_275;
assign n_540 = ~n_276 & ~n_539;
assign n_541 =  x_92 & ~n_266;
assign n_542 = ~n_267 & ~n_541;
assign n_543 =  x_94 & ~n_284;
assign n_544 = ~n_285 & ~n_543;
assign n_545 =  x_91 & ~n_248;
assign n_546 = ~n_249 & ~n_545;
assign n_547 =  x_96 & ~n_302;
assign n_548 = ~n_303 & ~n_547;
assign n_549 =  x_93 & ~n_230;
assign n_550 = ~n_231 & ~n_549;
assign n_551 =  x_98 & ~n_320;
assign n_552 = ~n_321 & ~n_551;
assign n_553 =  x_95 & ~n_212;
assign n_554 = ~n_213 & ~n_553;
assign n_555 =  x_100 & ~n_338;
assign n_556 = ~n_339 & ~n_555;
assign n_557 =  x_97 & ~n_194;
assign n_558 = ~n_195 & ~n_557;
assign n_559 =  x_102 & ~n_356;
assign n_560 = ~n_357 & ~n_559;
assign n_561 =  x_99 & ~n_176;
assign n_562 = ~n_177 & ~n_561;
assign n_563 =  x_104 & ~n_374;
assign n_564 = ~n_375 & ~n_563;
assign n_565 =  x_101 & ~n_158;
assign n_566 = ~n_159 & ~n_565;
assign n_567 =  x_106 & ~n_392;
assign n_568 = ~n_393 & ~n_567;
assign n_569 =  x_103 & ~n_140;
assign n_570 = ~n_141 & ~n_569;
assign n_571 =  x_108 & ~n_410;
assign n_572 = ~n_411 & ~n_571;
assign n_573 =  x_105 & ~n_122;
assign n_574 = ~n_123 & ~n_573;
assign n_575 =  x_110 & ~n_428;
assign n_576 = ~n_429 & ~n_575;
assign n_577 =  x_107 & ~n_104;
assign n_578 = ~n_105 & ~n_577;
assign n_579 =  x_112 & ~n_446;
assign n_580 = ~n_447 & ~n_579;
assign n_581 =  x_109 & ~n_86;
assign n_582 = ~n_87 & ~n_581;
assign n_583 =  x_114 & ~n_464;
assign n_584 = ~n_465 & ~n_583;
assign n_585 =  x_111 & ~n_68;
assign n_586 = ~n_69 & ~n_585;
assign n_587 =  x_116 & ~n_482;
assign n_588 = ~n_483 & ~n_587;
assign n_589 =  x_113 & ~n_50;
assign n_590 = ~n_51 & ~n_589;
assign n_591 = ~n_478 & ~n_485;
assign n_592 =  x_64 & ~n_591;
assign n_593 = ~n_485 & ~n_490;
assign n_594 = ~x_64 & ~n_593;
assign n_595 =  x_64 & ~n_488;
assign n_596 = ~x_64 & ~n_478;
assign n_597 = ~n_595 & ~n_596;
assign n_598 = ~n_594 & ~n_597;
assign n_599 = ~n_592 &  n_598;
assign n_600 =  x_118 & ~n_598;
assign n_601 = ~n_599 & ~n_600;
assign n_602 =  x_115 & ~n_30;
assign n_603 = ~n_31 & ~n_602;
assign n_604 = ~n_594 & ~n_599;
assign n_605 = ~x_118 & ~n_604;
assign n_606 = ~n_592 & ~n_594;
assign n_607 =  x_118 & ~n_606;
assign n_608 =  x_118 & ~n_597;
assign n_609 = ~x_118 & ~n_592;
assign n_610 = ~n_608 & ~n_609;
assign n_611 = ~n_605 & ~n_610;
assign n_612 = ~n_607 &  n_611;
assign n_613 = ~n_605 & ~n_612;
assign n_614 = ~x_62 & ~n_613;
assign n_615 = ~n_605 & ~n_607;
assign n_616 =  x_62 & ~n_615;
assign n_617 = ~x_120 & ~n_616;
assign n_618 = ~n_614 &  n_617;
assign n_619 =  x_62 & ~n_610;
assign n_620 = ~x_62 & ~n_607;
assign n_621 = ~n_619 & ~n_620;
assign n_622 = ~n_618 &  n_621;
assign n_623 = ~x_120 & ~n_621;
assign n_624 = ~n_622 & ~n_623;
assign n_625 = ~n_614 & ~n_621;
assign n_626 =  x_120 & ~n_625;
assign n_627 = ~n_616 &  n_625;
assign n_628 = ~n_626 & ~n_627;
assign n_629 = ~n_624 & ~n_628;
assign n_630 = ~n_5 &  n_17;
assign n_631 =  x_117 & ~n_630;
assign n_632 = ~n_1 &  n_630;
assign n_633 = ~n_631 & ~n_632;
assign n_634 =  n_624 &  n_633;
assign n_635 = ~n_624 & ~n_633;
assign n_636 = ~n_634 & ~n_635;
assign n_637 =  n_628 & ~n_636;
assign n_638 = ~n_629 & ~n_637;
assign n_639 = ~n_603 & ~n_638;
assign n_640 = ~n_628 & ~n_633;
assign n_641 =  n_628 &  n_633;
assign n_642 = ~n_640 & ~n_641;
assign n_643 =  n_636 & ~n_642;
assign n_644 =  n_638 & ~n_643;
assign n_645 = ~n_637 & ~n_644;
assign n_646 =  n_603 & ~n_645;
assign n_647 = ~n_639 & ~n_646;
assign n_648 = ~n_601 & ~n_647;
assign n_649 = ~n_603 &  n_643;
assign n_650 =  n_603 &  n_629;
assign n_651 = ~n_649 & ~n_650;
assign n_652 = ~n_646 &  n_651;
assign n_653 = ~n_639 &  n_652;
assign n_654 = ~n_646 & ~n_653;
assign n_655 =  n_601 & ~n_654;
assign n_656 = ~n_648 & ~n_655;
assign n_657 = ~n_590 & ~n_656;
assign n_658 = ~n_601 & ~n_651;
assign n_659 =  n_601 &  n_639;
assign n_660 = ~n_658 & ~n_659;
assign n_661 = ~n_655 &  n_660;
assign n_662 = ~n_648 &  n_661;
assign n_663 = ~n_655 & ~n_662;
assign n_664 =  n_590 & ~n_663;
assign n_665 = ~n_657 & ~n_664;
assign n_666 = ~n_588 & ~n_665;
assign n_667 =  n_590 & ~n_648;
assign n_668 = ~n_590 &  n_660;
assign n_669 = ~n_667 & ~n_668;
assign n_670 = ~n_664 & ~n_669;
assign n_671 = ~n_657 &  n_670;
assign n_672 = ~n_664 & ~n_671;
assign n_673 =  n_588 & ~n_672;
assign n_674 = ~n_666 & ~n_673;
assign n_675 = ~n_586 & ~n_674;
assign n_676 = ~n_588 & ~n_669;
assign n_677 =  n_588 & ~n_657;
assign n_678 = ~n_676 & ~n_677;
assign n_679 = ~n_673 & ~n_678;
assign n_680 = ~n_666 &  n_679;
assign n_681 = ~n_673 & ~n_680;
assign n_682 =  n_586 & ~n_681;
assign n_683 = ~n_675 & ~n_682;
assign n_684 = ~n_584 & ~n_683;
assign n_685 = ~n_586 & ~n_678;
assign n_686 =  n_586 & ~n_666;
assign n_687 = ~n_685 & ~n_686;
assign n_688 = ~n_682 & ~n_687;
assign n_689 = ~n_675 &  n_688;
assign n_690 = ~n_682 & ~n_689;
assign n_691 =  n_584 & ~n_690;
assign n_692 = ~n_684 & ~n_691;
assign n_693 = ~n_582 & ~n_692;
assign n_694 = ~n_584 & ~n_687;
assign n_695 =  n_584 & ~n_675;
assign n_696 = ~n_694 & ~n_695;
assign n_697 = ~n_691 & ~n_696;
assign n_698 = ~n_684 &  n_697;
assign n_699 = ~n_691 & ~n_698;
assign n_700 =  n_582 & ~n_699;
assign n_701 = ~n_693 & ~n_700;
assign n_702 = ~n_580 & ~n_701;
assign n_703 = ~n_582 & ~n_696;
assign n_704 =  n_582 & ~n_684;
assign n_705 = ~n_703 & ~n_704;
assign n_706 = ~n_700 & ~n_705;
assign n_707 = ~n_693 &  n_706;
assign n_708 = ~n_700 & ~n_707;
assign n_709 =  n_580 & ~n_708;
assign n_710 = ~n_702 & ~n_709;
assign n_711 = ~n_578 & ~n_710;
assign n_712 = ~n_580 & ~n_705;
assign n_713 =  n_580 & ~n_693;
assign n_714 = ~n_712 & ~n_713;
assign n_715 = ~n_709 & ~n_714;
assign n_716 = ~n_702 &  n_715;
assign n_717 = ~n_709 & ~n_716;
assign n_718 =  n_578 & ~n_717;
assign n_719 = ~n_711 & ~n_718;
assign n_720 = ~n_576 & ~n_719;
assign n_721 = ~n_578 & ~n_714;
assign n_722 =  n_578 & ~n_702;
assign n_723 = ~n_721 & ~n_722;
assign n_724 = ~n_718 & ~n_723;
assign n_725 = ~n_711 &  n_724;
assign n_726 = ~n_718 & ~n_725;
assign n_727 =  n_576 & ~n_726;
assign n_728 = ~n_720 & ~n_727;
assign n_729 = ~n_574 & ~n_728;
assign n_730 = ~n_576 & ~n_723;
assign n_731 =  n_576 & ~n_711;
assign n_732 = ~n_730 & ~n_731;
assign n_733 = ~n_727 & ~n_732;
assign n_734 = ~n_720 &  n_733;
assign n_735 = ~n_727 & ~n_734;
assign n_736 =  n_574 & ~n_735;
assign n_737 = ~n_729 & ~n_736;
assign n_738 = ~n_572 & ~n_737;
assign n_739 = ~n_574 & ~n_732;
assign n_740 =  n_574 & ~n_720;
assign n_741 = ~n_739 & ~n_740;
assign n_742 = ~n_736 & ~n_741;
assign n_743 = ~n_729 &  n_742;
assign n_744 = ~n_736 & ~n_743;
assign n_745 =  n_572 & ~n_744;
assign n_746 = ~n_738 & ~n_745;
assign n_747 = ~n_570 & ~n_746;
assign n_748 = ~n_572 & ~n_741;
assign n_749 =  n_572 & ~n_729;
assign n_750 = ~n_748 & ~n_749;
assign n_751 = ~n_745 & ~n_750;
assign n_752 = ~n_738 &  n_751;
assign n_753 = ~n_745 & ~n_752;
assign n_754 =  n_570 & ~n_753;
assign n_755 = ~n_747 & ~n_754;
assign n_756 = ~n_568 & ~n_755;
assign n_757 = ~n_570 & ~n_750;
assign n_758 =  n_570 & ~n_738;
assign n_759 = ~n_757 & ~n_758;
assign n_760 = ~n_754 & ~n_759;
assign n_761 = ~n_747 &  n_760;
assign n_762 = ~n_754 & ~n_761;
assign n_763 =  n_568 & ~n_762;
assign n_764 = ~n_756 & ~n_763;
assign n_765 = ~n_566 & ~n_764;
assign n_766 = ~n_568 & ~n_759;
assign n_767 =  n_568 & ~n_747;
assign n_768 = ~n_766 & ~n_767;
assign n_769 = ~n_763 & ~n_768;
assign n_770 = ~n_756 &  n_769;
assign n_771 = ~n_763 & ~n_770;
assign n_772 =  n_566 & ~n_771;
assign n_773 = ~n_765 & ~n_772;
assign n_774 = ~n_564 & ~n_773;
assign n_775 = ~n_566 & ~n_768;
assign n_776 =  n_566 & ~n_756;
assign n_777 = ~n_775 & ~n_776;
assign n_778 = ~n_772 & ~n_777;
assign n_779 = ~n_765 &  n_778;
assign n_780 = ~n_772 & ~n_779;
assign n_781 =  n_564 & ~n_780;
assign n_782 = ~n_774 & ~n_781;
assign n_783 = ~n_562 & ~n_782;
assign n_784 = ~n_564 & ~n_777;
assign n_785 =  n_564 & ~n_765;
assign n_786 = ~n_784 & ~n_785;
assign n_787 = ~n_781 & ~n_786;
assign n_788 = ~n_774 &  n_787;
assign n_789 = ~n_781 & ~n_788;
assign n_790 =  n_562 & ~n_789;
assign n_791 = ~n_783 & ~n_790;
assign n_792 = ~n_560 & ~n_791;
assign n_793 = ~n_562 & ~n_786;
assign n_794 =  n_562 & ~n_774;
assign n_795 = ~n_793 & ~n_794;
assign n_796 = ~n_790 & ~n_795;
assign n_797 = ~n_783 &  n_796;
assign n_798 = ~n_790 & ~n_797;
assign n_799 =  n_560 & ~n_798;
assign n_800 = ~n_792 & ~n_799;
assign n_801 = ~n_558 & ~n_800;
assign n_802 = ~n_560 & ~n_795;
assign n_803 =  n_560 & ~n_783;
assign n_804 = ~n_802 & ~n_803;
assign n_805 = ~n_799 & ~n_804;
assign n_806 = ~n_792 &  n_805;
assign n_807 = ~n_799 & ~n_806;
assign n_808 =  n_558 & ~n_807;
assign n_809 = ~n_801 & ~n_808;
assign n_810 = ~n_556 & ~n_809;
assign n_811 = ~n_558 & ~n_804;
assign n_812 =  n_558 & ~n_792;
assign n_813 = ~n_811 & ~n_812;
assign n_814 = ~n_808 & ~n_813;
assign n_815 = ~n_801 &  n_814;
assign n_816 = ~n_808 & ~n_815;
assign n_817 =  n_556 & ~n_816;
assign n_818 = ~n_810 & ~n_817;
assign n_819 = ~n_554 & ~n_818;
assign n_820 = ~n_556 & ~n_813;
assign n_821 =  n_556 & ~n_801;
assign n_822 = ~n_820 & ~n_821;
assign n_823 = ~n_817 & ~n_822;
assign n_824 = ~n_810 &  n_823;
assign n_825 = ~n_817 & ~n_824;
assign n_826 =  n_554 & ~n_825;
assign n_827 = ~n_819 & ~n_826;
assign n_828 = ~n_552 & ~n_827;
assign n_829 = ~n_554 & ~n_822;
assign n_830 =  n_554 & ~n_810;
assign n_831 = ~n_829 & ~n_830;
assign n_832 = ~n_826 & ~n_831;
assign n_833 = ~n_819 &  n_832;
assign n_834 = ~n_826 & ~n_833;
assign n_835 =  n_552 & ~n_834;
assign n_836 = ~n_828 & ~n_835;
assign n_837 = ~n_550 & ~n_836;
assign n_838 = ~n_552 & ~n_831;
assign n_839 =  n_552 & ~n_819;
assign n_840 = ~n_838 & ~n_839;
assign n_841 = ~n_835 & ~n_840;
assign n_842 = ~n_828 &  n_841;
assign n_843 = ~n_835 & ~n_842;
assign n_844 =  n_550 & ~n_843;
assign n_845 = ~n_837 & ~n_844;
assign n_846 = ~n_548 & ~n_845;
assign n_847 = ~n_550 & ~n_840;
assign n_848 =  n_550 & ~n_828;
assign n_849 = ~n_847 & ~n_848;
assign n_850 = ~n_844 & ~n_849;
assign n_851 = ~n_837 &  n_850;
assign n_852 = ~n_844 & ~n_851;
assign n_853 =  n_548 & ~n_852;
assign n_854 = ~n_846 & ~n_853;
assign n_855 = ~n_546 & ~n_854;
assign n_856 = ~n_548 & ~n_849;
assign n_857 =  n_548 & ~n_837;
assign n_858 = ~n_856 & ~n_857;
assign n_859 = ~n_853 & ~n_858;
assign n_860 = ~n_846 &  n_859;
assign n_861 = ~n_853 & ~n_860;
assign n_862 =  n_546 & ~n_861;
assign n_863 = ~n_855 & ~n_862;
assign n_864 = ~n_544 & ~n_863;
assign n_865 = ~n_546 & ~n_858;
assign n_866 =  n_546 & ~n_846;
assign n_867 = ~n_865 & ~n_866;
assign n_868 = ~n_862 & ~n_867;
assign n_869 = ~n_855 &  n_868;
assign n_870 = ~n_862 & ~n_869;
assign n_871 =  n_544 & ~n_870;
assign n_872 = ~n_864 & ~n_871;
assign n_873 = ~n_542 & ~n_872;
assign n_874 = ~n_544 & ~n_867;
assign n_875 =  n_544 & ~n_855;
assign n_876 = ~n_874 & ~n_875;
assign n_877 = ~n_871 & ~n_876;
assign n_878 = ~n_864 &  n_877;
assign n_879 = ~n_871 & ~n_878;
assign n_880 =  n_542 & ~n_879;
assign n_881 = ~n_873 & ~n_880;
assign n_882 = ~n_540 & ~n_881;
assign n_883 = ~n_542 & ~n_876;
assign n_884 =  n_542 & ~n_864;
assign n_885 = ~n_883 & ~n_884;
assign n_886 = ~n_880 & ~n_885;
assign n_887 = ~n_873 &  n_886;
assign n_888 = ~n_880 & ~n_887;
assign n_889 =  n_540 & ~n_888;
assign n_890 = ~n_882 & ~n_889;
assign n_891 = ~n_538 & ~n_890;
assign n_892 = ~n_540 & ~n_885;
assign n_893 =  n_540 & ~n_873;
assign n_894 = ~n_892 & ~n_893;
assign n_895 = ~n_889 & ~n_894;
assign n_896 = ~n_882 &  n_895;
assign n_897 = ~n_889 & ~n_896;
assign n_898 =  n_538 & ~n_897;
assign n_899 = ~n_891 & ~n_898;
assign n_900 = ~n_536 & ~n_899;
assign n_901 = ~n_538 & ~n_894;
assign n_902 =  n_538 & ~n_882;
assign n_903 = ~n_901 & ~n_902;
assign n_904 = ~n_898 & ~n_903;
assign n_905 = ~n_891 &  n_904;
assign n_906 = ~n_898 & ~n_905;
assign n_907 =  n_536 & ~n_906;
assign n_908 = ~n_900 & ~n_907;
assign n_909 = ~n_534 & ~n_908;
assign n_910 = ~n_536 & ~n_903;
assign n_911 =  n_536 & ~n_891;
assign n_912 = ~n_910 & ~n_911;
assign n_913 = ~n_907 & ~n_912;
assign n_914 = ~n_900 &  n_913;
assign n_915 = ~n_907 & ~n_914;
assign n_916 =  n_534 & ~n_915;
assign n_917 = ~n_909 & ~n_916;
assign n_918 = ~n_532 & ~n_917;
assign n_919 = ~n_534 & ~n_912;
assign n_920 =  n_534 & ~n_900;
assign n_921 = ~n_919 & ~n_920;
assign n_922 = ~n_916 & ~n_921;
assign n_923 = ~n_909 &  n_922;
assign n_924 = ~n_916 & ~n_923;
assign n_925 =  n_532 & ~n_924;
assign n_926 = ~n_918 & ~n_925;
assign n_927 = ~n_530 & ~n_926;
assign n_928 = ~n_532 & ~n_921;
assign n_929 =  n_532 & ~n_909;
assign n_930 = ~n_928 & ~n_929;
assign n_931 = ~n_925 & ~n_930;
assign n_932 = ~n_918 &  n_931;
assign n_933 = ~n_925 & ~n_932;
assign n_934 =  n_530 & ~n_933;
assign n_935 = ~n_927 & ~n_934;
assign n_936 = ~n_528 & ~n_935;
assign n_937 = ~n_530 & ~n_930;
assign n_938 =  n_530 & ~n_918;
assign n_939 = ~n_937 & ~n_938;
assign n_940 = ~n_934 & ~n_939;
assign n_941 = ~n_927 &  n_940;
assign n_942 = ~n_934 & ~n_941;
assign n_943 =  n_528 & ~n_942;
assign n_944 = ~n_936 & ~n_943;
assign n_945 = ~n_526 & ~n_944;
assign n_946 = ~n_528 & ~n_939;
assign n_947 =  n_528 & ~n_927;
assign n_948 = ~n_946 & ~n_947;
assign n_949 = ~n_943 & ~n_948;
assign n_950 = ~n_936 &  n_949;
assign n_951 = ~n_943 & ~n_950;
assign n_952 =  n_526 & ~n_951;
assign n_953 = ~n_945 & ~n_952;
assign n_954 = ~n_524 & ~n_953;
assign n_955 = ~n_526 & ~n_948;
assign n_956 =  n_526 & ~n_936;
assign n_957 = ~n_955 & ~n_956;
assign n_958 = ~n_952 & ~n_957;
assign n_959 = ~n_945 &  n_958;
assign n_960 = ~n_952 & ~n_959;
assign n_961 =  n_524 & ~n_960;
assign n_962 = ~n_954 & ~n_961;
assign n_963 = ~n_522 & ~n_962;
assign n_964 = ~n_524 & ~n_957;
assign n_965 =  n_524 & ~n_945;
assign n_966 = ~n_964 & ~n_965;
assign n_967 = ~n_961 & ~n_966;
assign n_968 = ~n_954 &  n_967;
assign n_969 = ~n_961 & ~n_968;
assign n_970 =  n_522 & ~n_969;
assign n_971 = ~n_963 & ~n_970;
assign n_972 = ~n_520 & ~n_971;
assign n_973 = ~n_522 & ~n_966;
assign n_974 =  n_522 & ~n_954;
assign n_975 = ~n_973 & ~n_974;
assign n_976 = ~n_970 & ~n_975;
assign n_977 = ~n_963 &  n_976;
assign n_978 = ~n_970 & ~n_977;
assign n_979 =  n_520 & ~n_978;
assign n_980 = ~n_972 & ~n_979;
assign n_981 = ~n_518 & ~n_980;
assign n_982 = ~n_520 & ~n_975;
assign n_983 =  n_520 & ~n_963;
assign n_984 = ~n_982 & ~n_983;
assign n_985 = ~n_979 & ~n_984;
assign n_986 = ~n_972 &  n_985;
assign n_987 = ~n_979 & ~n_986;
assign n_988 =  n_518 & ~n_987;
assign n_989 = ~n_981 & ~n_988;
assign n_990 = ~n_516 & ~n_989;
assign n_991 = ~n_518 & ~n_984;
assign n_992 =  n_518 & ~n_972;
assign n_993 = ~n_991 & ~n_992;
assign n_994 = ~n_988 & ~n_993;
assign n_995 = ~n_981 &  n_994;
assign n_996 = ~n_988 & ~n_995;
assign n_997 =  n_516 & ~n_996;
assign n_998 = ~n_990 & ~n_997;
assign n_999 = ~n_514 & ~n_998;
assign n_1000 = ~n_516 & ~n_993;
assign n_1001 =  n_516 & ~n_981;
assign n_1002 = ~n_1000 & ~n_1001;
assign n_1003 = ~n_997 & ~n_1002;
assign n_1004 = ~n_990 &  n_1003;
assign n_1005 = ~n_997 & ~n_1004;
assign n_1006 =  n_514 & ~n_1005;
assign n_1007 = ~n_999 & ~n_1006;
assign n_1008 = ~n_512 & ~n_1007;
assign n_1009 = ~n_514 & ~n_1002;
assign n_1010 =  n_514 & ~n_990;
assign n_1011 = ~n_1009 & ~n_1010;
assign n_1012 = ~n_1006 & ~n_1011;
assign n_1013 = ~n_999 &  n_1012;
assign n_1014 = ~n_1006 & ~n_1013;
assign n_1015 =  n_512 & ~n_1014;
assign n_1016 = ~n_1008 & ~n_1015;
assign n_1017 = ~n_510 & ~n_1016;
assign n_1018 = ~n_512 & ~n_1011;
assign n_1019 =  n_512 & ~n_999;
assign n_1020 = ~n_1018 & ~n_1019;
assign n_1021 = ~n_1015 & ~n_1020;
assign n_1022 = ~n_1008 &  n_1021;
assign n_1023 = ~n_1015 & ~n_1022;
assign n_1024 =  n_510 & ~n_1023;
assign n_1025 = ~n_1017 & ~n_1024;
assign n_1026 = ~n_508 & ~n_1025;
assign n_1027 = ~n_510 & ~n_1020;
assign n_1028 =  n_510 & ~n_1008;
assign n_1029 = ~n_1027 & ~n_1028;
assign n_1030 = ~n_1024 & ~n_1029;
assign n_1031 = ~n_1017 &  n_1030;
assign n_1032 = ~n_1024 & ~n_1031;
assign n_1033 =  n_508 & ~n_1032;
assign n_1034 = ~n_1026 & ~n_1033;
assign n_1035 = ~n_506 & ~n_1034;
assign n_1036 = ~n_508 & ~n_1029;
assign n_1037 =  n_508 & ~n_1017;
assign n_1038 = ~n_1036 & ~n_1037;
assign n_1039 = ~n_1033 & ~n_1038;
assign n_1040 = ~n_1026 &  n_1039;
assign n_1041 = ~n_1033 & ~n_1040;
assign n_1042 =  n_506 & ~n_1041;
assign n_1043 = ~n_1035 & ~n_1042;
assign n_1044 = ~n_504 & ~n_1043;
assign n_1045 = ~n_506 & ~n_1038;
assign n_1046 =  n_506 & ~n_1026;
assign n_1047 = ~n_1045 & ~n_1046;
assign n_1048 = ~n_1042 & ~n_1047;
assign n_1049 = ~n_1035 &  n_1048;
assign n_1050 = ~n_1042 & ~n_1049;
assign n_1051 =  n_504 & ~n_1050;
assign n_1052 = ~n_1044 & ~n_1051;
assign n_1053 = ~n_502 & ~n_1052;
assign n_1054 = ~n_504 & ~n_1047;
assign n_1055 =  n_504 & ~n_1035;
assign n_1056 = ~n_1054 & ~n_1055;
assign n_1057 = ~n_1051 & ~n_1056;
assign n_1058 = ~n_1044 &  n_1057;
assign n_1059 = ~n_1051 & ~n_1058;
assign n_1060 =  n_502 & ~n_1059;
assign n_1061 = ~n_1053 & ~n_1060;
assign n_1062 = ~n_500 & ~n_1061;
assign n_1063 = ~n_502 & ~n_1056;
assign n_1064 =  n_502 & ~n_1044;
assign n_1065 = ~n_1063 & ~n_1064;
assign n_1066 = ~n_1060 & ~n_1065;
assign n_1067 = ~n_1053 &  n_1066;
assign n_1068 = ~n_1060 & ~n_1067;
assign n_1069 =  n_500 & ~n_1068;
assign n_1070 = ~n_1062 & ~n_1069;
assign n_1071 = ~n_498 & ~n_1070;
assign n_1072 = ~n_500 & ~n_1065;
assign n_1073 =  n_500 & ~n_1053;
assign n_1074 = ~n_1072 & ~n_1073;
assign n_1075 = ~n_1069 & ~n_1074;
assign n_1076 = ~n_1062 &  n_1075;
assign n_1077 = ~n_1069 & ~n_1076;
assign n_1078 =  n_498 & ~n_1077;
assign n_1079 = ~n_1071 & ~n_1078;
assign n_1080 = ~n_496 & ~n_1079;
assign n_1081 = ~n_498 & ~n_1074;
assign n_1082 =  n_498 & ~n_1062;
assign n_1083 = ~n_1081 & ~n_1082;
assign n_1084 = ~n_1078 & ~n_1083;
assign n_1085 = ~n_1071 &  n_1084;
assign n_1086 = ~n_1078 & ~n_1085;
assign n_1087 =  n_496 & ~n_1086;
assign n_1088 = ~n_1080 & ~n_1087;
assign n_1089 = ~n_494 & ~n_1088;
assign n_1090 = ~n_496 & ~n_1083;
assign n_1091 =  n_496 & ~n_1071;
assign n_1092 = ~n_1090 & ~n_1091;
assign n_1093 = ~n_1087 & ~n_1092;
assign n_1094 = ~n_1080 &  n_1093;
assign n_1095 = ~n_1087 & ~n_1094;
assign n_1096 =  n_494 & ~n_1095;
assign n_1097 = ~n_1089 & ~n_1096;
assign n_1098 = ~n_492 & ~n_1097;
assign n_1099 = ~n_494 & ~n_1092;
assign n_1100 =  n_494 & ~n_1080;
assign n_1101 = ~n_1099 & ~n_1100;
assign n_1102 = ~n_1096 & ~n_1101;
assign n_1103 = ~n_1089 &  n_1102;
assign n_1104 = ~n_1096 & ~n_1103;
assign n_1105 =  n_492 & ~n_1104;
assign n_1106 = ~n_1098 & ~n_1105;
assign n_1107 = ~n_40 & ~n_1106;
assign n_1108 = ~n_492 & ~n_1101;
assign n_1109 =  n_492 & ~n_1089;
assign n_1110 = ~n_1108 & ~n_1109;
assign n_1111 = ~n_1105 & ~n_1110;
assign n_1112 = ~n_1098 &  n_1111;
assign n_1113 = ~n_1105 & ~n_1112;
assign n_1114 =  n_40 & ~n_1113;
assign n_1115 = ~n_40 & ~n_1110;
assign n_1116 =  n_40 & ~n_1098;
assign n_1117 = ~n_1115 & ~n_1116;
assign n_1118 = ~n_1114 & ~n_1117;
assign n_1119 = ~n_1107 &  n_1118;
assign n_1120 =  x_62 & ~n_611;
assign n_1121 = ~n_612 & ~n_1120;
assign n_1122 = ~n_1118 & ~n_1121;
assign n_1123 = ~n_1119 & ~n_1122;
assign n_1124 = ~n_584 & ~n_688;
assign n_1125 = ~n_689 & ~n_1124;
assign n_1126 = ~n_492 & ~n_1102;
assign n_1127 = ~n_1103 & ~n_1126;
assign n_1128 = ~n_580 & ~n_706;
assign n_1129 = ~n_707 & ~n_1128;
assign n_1130 = ~n_496 & ~n_1084;
assign n_1131 = ~n_1085 & ~n_1130;
assign n_1132 = ~n_576 & ~n_724;
assign n_1133 = ~n_725 & ~n_1132;
assign n_1134 = ~n_500 & ~n_1066;
assign n_1135 = ~n_1067 & ~n_1134;
assign n_1136 = ~n_572 & ~n_742;
assign n_1137 = ~n_743 & ~n_1136;
assign n_1138 = ~n_504 & ~n_1048;
assign n_1139 = ~n_1049 & ~n_1138;
assign n_1140 = ~n_568 & ~n_760;
assign n_1141 = ~n_761 & ~n_1140;
assign n_1142 = ~n_508 & ~n_1030;
assign n_1143 = ~n_1031 & ~n_1142;
assign n_1144 = ~n_564 & ~n_778;
assign n_1145 = ~n_779 & ~n_1144;
assign n_1146 = ~n_512 & ~n_1012;
assign n_1147 = ~n_1013 & ~n_1146;
assign n_1148 = ~n_560 & ~n_796;
assign n_1149 = ~n_797 & ~n_1148;
assign n_1150 = ~n_516 & ~n_994;
assign n_1151 = ~n_995 & ~n_1150;
assign n_1152 = ~n_556 & ~n_814;
assign n_1153 = ~n_815 & ~n_1152;
assign n_1154 = ~n_520 & ~n_976;
assign n_1155 = ~n_977 & ~n_1154;
assign n_1156 = ~n_552 & ~n_832;
assign n_1157 = ~n_833 & ~n_1156;
assign n_1158 = ~n_524 & ~n_958;
assign n_1159 = ~n_959 & ~n_1158;
assign n_1160 = ~n_548 & ~n_850;
assign n_1161 = ~n_851 & ~n_1160;
assign n_1162 = ~n_528 & ~n_940;
assign n_1163 = ~n_941 & ~n_1162;
assign n_1164 = ~n_544 & ~n_868;
assign n_1165 = ~n_869 & ~n_1164;
assign n_1166 = ~n_532 & ~n_922;
assign n_1167 = ~n_923 & ~n_1166;
assign n_1168 = ~n_540 & ~n_886;
assign n_1169 = ~n_887 & ~n_1168;
assign n_1170 = ~n_536 & ~n_904;
assign n_1171 = ~n_905 & ~n_1170;
assign n_1172 = ~n_538 & ~n_895;
assign n_1173 = ~n_896 & ~n_1172;
assign n_1174 = ~n_534 & ~n_913;
assign n_1175 = ~n_914 & ~n_1174;
assign n_1176 = ~n_542 & ~n_877;
assign n_1177 = ~n_878 & ~n_1176;
assign n_1178 = ~n_530 & ~n_931;
assign n_1179 = ~n_932 & ~n_1178;
assign n_1180 = ~n_546 & ~n_859;
assign n_1181 = ~n_860 & ~n_1180;
assign n_1182 = ~n_526 & ~n_949;
assign n_1183 = ~n_950 & ~n_1182;
assign n_1184 = ~n_550 & ~n_841;
assign n_1185 = ~n_842 & ~n_1184;
assign n_1186 = ~n_522 & ~n_967;
assign n_1187 = ~n_968 & ~n_1186;
assign n_1188 = ~n_554 & ~n_823;
assign n_1189 = ~n_824 & ~n_1188;
assign n_1190 = ~n_518 & ~n_985;
assign n_1191 = ~n_986 & ~n_1190;
assign n_1192 = ~n_558 & ~n_805;
assign n_1193 = ~n_806 & ~n_1192;
assign n_1194 = ~n_514 & ~n_1003;
assign n_1195 = ~n_1004 & ~n_1194;
assign n_1196 = ~n_562 & ~n_787;
assign n_1197 = ~n_788 & ~n_1196;
assign n_1198 = ~n_510 & ~n_1021;
assign n_1199 = ~n_1022 & ~n_1198;
assign n_1200 = ~n_566 & ~n_769;
assign n_1201 = ~n_770 & ~n_1200;
assign n_1202 = ~n_506 & ~n_1039;
assign n_1203 = ~n_1040 & ~n_1202;
assign n_1204 = ~n_570 & ~n_751;
assign n_1205 = ~n_752 & ~n_1204;
assign n_1206 = ~n_502 & ~n_1057;
assign n_1207 = ~n_1058 & ~n_1206;
assign n_1208 = ~n_574 & ~n_733;
assign n_1209 = ~n_734 & ~n_1208;
assign n_1210 = ~n_498 & ~n_1075;
assign n_1211 = ~n_1076 & ~n_1210;
assign n_1212 = ~n_578 & ~n_715;
assign n_1213 = ~n_716 & ~n_1212;
assign n_1214 = ~n_494 & ~n_1093;
assign n_1215 = ~n_1094 & ~n_1214;
assign n_1216 = ~n_582 & ~n_697;
assign n_1217 = ~n_698 & ~n_1216;
assign n_1218 = ~n_40 & ~n_1111;
assign n_1219 = ~n_1112 & ~n_1218;
assign n_1220 = ~n_586 & ~n_679;
assign n_1221 = ~n_680 & ~n_1220;
assign n_1222 = ~n_1107 & ~n_1114;
assign n_1223 = ~n_1121 & ~n_1222;
assign n_1224 = ~n_1114 & ~n_1119;
assign n_1225 =  n_1121 & ~n_1224;
assign n_1226 = ~n_1117 & ~n_1121;
assign n_1227 = ~n_1107 &  n_1121;
assign n_1228 = ~n_1226 & ~n_1227;
assign n_1229 = ~n_1225 & ~n_1228;
assign n_1230 = ~n_1223 &  n_1229;
assign n_1231 =  x_65 & ~n_21;
assign n_1232 = ~n_22 & ~n_1231;
assign n_1233 = ~n_1229 & ~n_1232;
assign n_1234 = ~n_1230 & ~n_1233;
assign n_1235 = ~n_590 & ~n_661;
assign n_1236 = ~n_662 & ~n_1235;
assign n_1237 = ~n_616 & ~n_623;
assign n_1238 =  n_616 &  n_623;
assign n_1239 = ~n_1237 & ~n_1238;
assign n_1240 = ~n_614 & ~n_1239;
assign n_1241 = ~n_1225 & ~n_1230;
assign n_1242 =  n_1232 & ~n_1241;
assign n_1243 = ~n_1223 & ~n_1225;
assign n_1244 = ~n_1232 & ~n_1243;
assign n_1245 = ~n_1228 & ~n_1232;
assign n_1246 = ~n_1223 &  n_1232;
assign n_1247 = ~n_1245 & ~n_1246;
assign n_1248 = ~n_1242 & ~n_1247;
assign n_1249 = ~n_1244 &  n_1248;
assign n_1250 = ~n_1242 & ~n_1249;
assign n_1251 =  n_1240 & ~n_1250;
assign n_1252 = ~n_1242 & ~n_1244;
assign n_1253 = ~n_1240 & ~n_1252;
assign n_1254 = ~n_1251 & ~n_1253;
assign n_1255 =  n_1240 & ~n_1244;
assign n_1256 = ~n_1240 & ~n_1247;
assign n_1257 = ~n_1255 & ~n_1256;
assign n_1258 =  n_1254 & ~n_1257;
assign n_1259 = ~n_1251 & ~n_1258;
assign n_1260 = ~n_8 & ~n_15;
assign n_1261 = ~n_1259 & ~n_1260;
assign n_1262 =  n_1253 & ~n_1260;
assign n_1263 =  n_1257 &  n_1260;
assign n_1264 = ~n_1262 & ~n_1263;
assign n_1265 = ~n_1261 &  n_1264;
assign n_1266 = ~n_637 & ~n_643;
assign n_1267 = ~n_603 & ~n_1266;
assign n_1268 = ~n_644 & ~n_1267;
assign n_1269 = ~n_1265 & ~n_1268;
assign n_1270 =  n_1265 &  n_1268;
assign n_1271 = ~n_1269 & ~n_1270;
assign n_1272 =  n_1251 &  n_1260;
assign n_1273 = ~n_1258 & ~n_1263;
assign n_1274 = ~n_1272 &  n_1273;
assign n_1275 = ~n_1271 &  n_1274;
assign n_1276 = ~n_1265 & ~n_1274;
assign n_1277 = ~n_1275 & ~n_1276;
assign n_1278 = ~n_1268 & ~n_1274;
assign n_1279 =  n_1265 & ~n_1278;
assign n_1280 = ~n_1269 & ~n_1279;
assign n_1281 =  n_1277 & ~n_1280;
assign n_1282 = ~n_1275 & ~n_1281;
assign n_1283 =  n_1236 & ~n_1282;
assign n_1284 = ~n_1236 & ~n_1277;
assign n_1285 = ~n_1283 & ~n_1284;
assign n_1286 = ~n_1234 & ~n_1285;
assign n_1287 =  n_1236 &  n_1276;
assign n_1288 = ~n_1236 & ~n_1276;
assign n_1289 =  n_1280 &  n_1288;
assign n_1290 = ~n_1287 & ~n_1289;
assign n_1291 = ~n_1283 &  n_1290;
assign n_1292 = ~n_1284 &  n_1291;
assign n_1293 = ~n_1283 & ~n_1292;
assign n_1294 =  n_1234 & ~n_1293;
assign n_1295 = ~n_1286 & ~n_1294;
assign n_1296 = ~n_1221 & ~n_1295;
assign n_1297 = ~n_1234 & ~n_1290;
assign n_1298 =  n_1234 &  n_1284;
assign n_1299 = ~n_1297 & ~n_1298;
assign n_1300 = ~n_1294 &  n_1299;
assign n_1301 = ~n_1286 &  n_1300;
assign n_1302 = ~n_1294 & ~n_1301;
assign n_1303 =  n_1221 & ~n_1302;
assign n_1304 = ~n_1296 & ~n_1303;
assign n_1305 = ~n_1219 & ~n_1304;
assign n_1306 =  n_1221 & ~n_1286;
assign n_1307 = ~n_1221 &  n_1299;
assign n_1308 = ~n_1306 & ~n_1307;
assign n_1309 = ~n_1303 & ~n_1308;
assign n_1310 = ~n_1296 &  n_1309;
assign n_1311 = ~n_1303 & ~n_1310;
assign n_1312 =  n_1219 & ~n_1311;
assign n_1313 = ~n_1305 & ~n_1312;
assign n_1314 = ~n_1217 & ~n_1313;
assign n_1315 = ~n_1219 & ~n_1308;
assign n_1316 =  n_1219 & ~n_1296;
assign n_1317 = ~n_1315 & ~n_1316;
assign n_1318 = ~n_1312 & ~n_1317;
assign n_1319 = ~n_1305 &  n_1318;
assign n_1320 = ~n_1312 & ~n_1319;
assign n_1321 =  n_1217 & ~n_1320;
assign n_1322 = ~n_1314 & ~n_1321;
assign n_1323 = ~n_1215 & ~n_1322;
assign n_1324 = ~n_1217 & ~n_1317;
assign n_1325 =  n_1217 & ~n_1305;
assign n_1326 = ~n_1324 & ~n_1325;
assign n_1327 = ~n_1321 & ~n_1326;
assign n_1328 = ~n_1314 &  n_1327;
assign n_1329 = ~n_1321 & ~n_1328;
assign n_1330 =  n_1215 & ~n_1329;
assign n_1331 = ~n_1323 & ~n_1330;
assign n_1332 = ~n_1213 & ~n_1331;
assign n_1333 = ~n_1215 & ~n_1326;
assign n_1334 =  n_1215 & ~n_1314;
assign n_1335 = ~n_1333 & ~n_1334;
assign n_1336 = ~n_1330 & ~n_1335;
assign n_1337 = ~n_1323 &  n_1336;
assign n_1338 = ~n_1330 & ~n_1337;
assign n_1339 =  n_1213 & ~n_1338;
assign n_1340 = ~n_1332 & ~n_1339;
assign n_1341 = ~n_1211 & ~n_1340;
assign n_1342 = ~n_1213 & ~n_1335;
assign n_1343 =  n_1213 & ~n_1323;
assign n_1344 = ~n_1342 & ~n_1343;
assign n_1345 = ~n_1339 & ~n_1344;
assign n_1346 = ~n_1332 &  n_1345;
assign n_1347 = ~n_1339 & ~n_1346;
assign n_1348 =  n_1211 & ~n_1347;
assign n_1349 = ~n_1341 & ~n_1348;
assign n_1350 = ~n_1209 & ~n_1349;
assign n_1351 = ~n_1211 & ~n_1344;
assign n_1352 =  n_1211 & ~n_1332;
assign n_1353 = ~n_1351 & ~n_1352;
assign n_1354 = ~n_1348 & ~n_1353;
assign n_1355 = ~n_1341 &  n_1354;
assign n_1356 = ~n_1348 & ~n_1355;
assign n_1357 =  n_1209 & ~n_1356;
assign n_1358 = ~n_1350 & ~n_1357;
assign n_1359 = ~n_1207 & ~n_1358;
assign n_1360 = ~n_1209 & ~n_1353;
assign n_1361 =  n_1209 & ~n_1341;
assign n_1362 = ~n_1360 & ~n_1361;
assign n_1363 = ~n_1357 & ~n_1362;
assign n_1364 = ~n_1350 &  n_1363;
assign n_1365 = ~n_1357 & ~n_1364;
assign n_1366 =  n_1207 & ~n_1365;
assign n_1367 = ~n_1359 & ~n_1366;
assign n_1368 = ~n_1205 & ~n_1367;
assign n_1369 = ~n_1207 & ~n_1362;
assign n_1370 =  n_1207 & ~n_1350;
assign n_1371 = ~n_1369 & ~n_1370;
assign n_1372 = ~n_1366 & ~n_1371;
assign n_1373 = ~n_1359 &  n_1372;
assign n_1374 = ~n_1366 & ~n_1373;
assign n_1375 =  n_1205 & ~n_1374;
assign n_1376 = ~n_1368 & ~n_1375;
assign n_1377 = ~n_1203 & ~n_1376;
assign n_1378 = ~n_1205 & ~n_1371;
assign n_1379 =  n_1205 & ~n_1359;
assign n_1380 = ~n_1378 & ~n_1379;
assign n_1381 = ~n_1375 & ~n_1380;
assign n_1382 = ~n_1368 &  n_1381;
assign n_1383 = ~n_1375 & ~n_1382;
assign n_1384 =  n_1203 & ~n_1383;
assign n_1385 = ~n_1377 & ~n_1384;
assign n_1386 = ~n_1201 & ~n_1385;
assign n_1387 = ~n_1203 & ~n_1380;
assign n_1388 =  n_1203 & ~n_1368;
assign n_1389 = ~n_1387 & ~n_1388;
assign n_1390 = ~n_1384 & ~n_1389;
assign n_1391 = ~n_1377 &  n_1390;
assign n_1392 = ~n_1384 & ~n_1391;
assign n_1393 =  n_1201 & ~n_1392;
assign n_1394 = ~n_1386 & ~n_1393;
assign n_1395 = ~n_1199 & ~n_1394;
assign n_1396 = ~n_1201 & ~n_1389;
assign n_1397 =  n_1201 & ~n_1377;
assign n_1398 = ~n_1396 & ~n_1397;
assign n_1399 = ~n_1393 & ~n_1398;
assign n_1400 = ~n_1386 &  n_1399;
assign n_1401 = ~n_1393 & ~n_1400;
assign n_1402 =  n_1199 & ~n_1401;
assign n_1403 = ~n_1395 & ~n_1402;
assign n_1404 = ~n_1197 & ~n_1403;
assign n_1405 = ~n_1199 & ~n_1398;
assign n_1406 =  n_1199 & ~n_1386;
assign n_1407 = ~n_1405 & ~n_1406;
assign n_1408 = ~n_1402 & ~n_1407;
assign n_1409 = ~n_1395 &  n_1408;
assign n_1410 = ~n_1402 & ~n_1409;
assign n_1411 =  n_1197 & ~n_1410;
assign n_1412 = ~n_1404 & ~n_1411;
assign n_1413 = ~n_1195 & ~n_1412;
assign n_1414 = ~n_1197 & ~n_1407;
assign n_1415 =  n_1197 & ~n_1395;
assign n_1416 = ~n_1414 & ~n_1415;
assign n_1417 = ~n_1411 & ~n_1416;
assign n_1418 = ~n_1404 &  n_1417;
assign n_1419 = ~n_1411 & ~n_1418;
assign n_1420 =  n_1195 & ~n_1419;
assign n_1421 = ~n_1413 & ~n_1420;
assign n_1422 = ~n_1193 & ~n_1421;
assign n_1423 = ~n_1195 & ~n_1416;
assign n_1424 =  n_1195 & ~n_1404;
assign n_1425 = ~n_1423 & ~n_1424;
assign n_1426 = ~n_1420 & ~n_1425;
assign n_1427 = ~n_1413 &  n_1426;
assign n_1428 = ~n_1420 & ~n_1427;
assign n_1429 =  n_1193 & ~n_1428;
assign n_1430 = ~n_1422 & ~n_1429;
assign n_1431 = ~n_1191 & ~n_1430;
assign n_1432 = ~n_1193 & ~n_1425;
assign n_1433 =  n_1193 & ~n_1413;
assign n_1434 = ~n_1432 & ~n_1433;
assign n_1435 = ~n_1429 & ~n_1434;
assign n_1436 = ~n_1422 &  n_1435;
assign n_1437 = ~n_1429 & ~n_1436;
assign n_1438 =  n_1191 & ~n_1437;
assign n_1439 = ~n_1431 & ~n_1438;
assign n_1440 = ~n_1189 & ~n_1439;
assign n_1441 = ~n_1191 & ~n_1434;
assign n_1442 =  n_1191 & ~n_1422;
assign n_1443 = ~n_1441 & ~n_1442;
assign n_1444 = ~n_1438 & ~n_1443;
assign n_1445 = ~n_1431 &  n_1444;
assign n_1446 = ~n_1438 & ~n_1445;
assign n_1447 =  n_1189 & ~n_1446;
assign n_1448 = ~n_1440 & ~n_1447;
assign n_1449 = ~n_1187 & ~n_1448;
assign n_1450 = ~n_1189 & ~n_1443;
assign n_1451 =  n_1189 & ~n_1431;
assign n_1452 = ~n_1450 & ~n_1451;
assign n_1453 = ~n_1447 & ~n_1452;
assign n_1454 = ~n_1440 &  n_1453;
assign n_1455 = ~n_1447 & ~n_1454;
assign n_1456 =  n_1187 & ~n_1455;
assign n_1457 = ~n_1449 & ~n_1456;
assign n_1458 = ~n_1185 & ~n_1457;
assign n_1459 = ~n_1187 & ~n_1452;
assign n_1460 =  n_1187 & ~n_1440;
assign n_1461 = ~n_1459 & ~n_1460;
assign n_1462 = ~n_1456 & ~n_1461;
assign n_1463 = ~n_1449 &  n_1462;
assign n_1464 = ~n_1456 & ~n_1463;
assign n_1465 =  n_1185 & ~n_1464;
assign n_1466 = ~n_1458 & ~n_1465;
assign n_1467 = ~n_1183 & ~n_1466;
assign n_1468 = ~n_1185 & ~n_1461;
assign n_1469 =  n_1185 & ~n_1449;
assign n_1470 = ~n_1468 & ~n_1469;
assign n_1471 = ~n_1465 & ~n_1470;
assign n_1472 = ~n_1458 &  n_1471;
assign n_1473 = ~n_1465 & ~n_1472;
assign n_1474 =  n_1183 & ~n_1473;
assign n_1475 = ~n_1467 & ~n_1474;
assign n_1476 = ~n_1181 & ~n_1475;
assign n_1477 = ~n_1183 & ~n_1470;
assign n_1478 =  n_1183 & ~n_1458;
assign n_1479 = ~n_1477 & ~n_1478;
assign n_1480 = ~n_1474 & ~n_1479;
assign n_1481 = ~n_1467 &  n_1480;
assign n_1482 = ~n_1474 & ~n_1481;
assign n_1483 =  n_1181 & ~n_1482;
assign n_1484 = ~n_1476 & ~n_1483;
assign n_1485 = ~n_1179 & ~n_1484;
assign n_1486 = ~n_1181 & ~n_1479;
assign n_1487 =  n_1181 & ~n_1467;
assign n_1488 = ~n_1486 & ~n_1487;
assign n_1489 = ~n_1483 & ~n_1488;
assign n_1490 = ~n_1476 &  n_1489;
assign n_1491 = ~n_1483 & ~n_1490;
assign n_1492 =  n_1179 & ~n_1491;
assign n_1493 = ~n_1485 & ~n_1492;
assign n_1494 = ~n_1177 & ~n_1493;
assign n_1495 = ~n_1179 & ~n_1488;
assign n_1496 =  n_1179 & ~n_1476;
assign n_1497 = ~n_1495 & ~n_1496;
assign n_1498 = ~n_1492 & ~n_1497;
assign n_1499 = ~n_1485 &  n_1498;
assign n_1500 = ~n_1492 & ~n_1499;
assign n_1501 =  n_1177 & ~n_1500;
assign n_1502 = ~n_1494 & ~n_1501;
assign n_1503 = ~n_1175 & ~n_1502;
assign n_1504 = ~n_1177 & ~n_1497;
assign n_1505 =  n_1177 & ~n_1485;
assign n_1506 = ~n_1504 & ~n_1505;
assign n_1507 = ~n_1501 & ~n_1506;
assign n_1508 = ~n_1494 &  n_1507;
assign n_1509 = ~n_1501 & ~n_1508;
assign n_1510 =  n_1175 & ~n_1509;
assign n_1511 = ~n_1503 & ~n_1510;
assign n_1512 = ~n_1173 & ~n_1511;
assign n_1513 = ~n_1175 & ~n_1506;
assign n_1514 =  n_1175 & ~n_1494;
assign n_1515 = ~n_1513 & ~n_1514;
assign n_1516 = ~n_1510 & ~n_1515;
assign n_1517 = ~n_1503 &  n_1516;
assign n_1518 = ~n_1510 & ~n_1517;
assign n_1519 =  n_1173 & ~n_1518;
assign n_1520 = ~n_1512 & ~n_1519;
assign n_1521 = ~n_1171 & ~n_1520;
assign n_1522 = ~n_1173 & ~n_1515;
assign n_1523 =  n_1173 & ~n_1503;
assign n_1524 = ~n_1522 & ~n_1523;
assign n_1525 = ~n_1519 & ~n_1524;
assign n_1526 = ~n_1512 &  n_1525;
assign n_1527 = ~n_1519 & ~n_1526;
assign n_1528 =  n_1171 & ~n_1527;
assign n_1529 = ~n_1521 & ~n_1528;
assign n_1530 = ~n_1169 & ~n_1529;
assign n_1531 = ~n_1171 & ~n_1524;
assign n_1532 =  n_1171 & ~n_1512;
assign n_1533 = ~n_1531 & ~n_1532;
assign n_1534 = ~n_1528 & ~n_1533;
assign n_1535 = ~n_1521 &  n_1534;
assign n_1536 = ~n_1528 & ~n_1535;
assign n_1537 =  n_1169 & ~n_1536;
assign n_1538 = ~n_1530 & ~n_1537;
assign n_1539 = ~n_1167 & ~n_1538;
assign n_1540 = ~n_1169 & ~n_1533;
assign n_1541 =  n_1169 & ~n_1521;
assign n_1542 = ~n_1540 & ~n_1541;
assign n_1543 = ~n_1537 & ~n_1542;
assign n_1544 = ~n_1530 &  n_1543;
assign n_1545 = ~n_1537 & ~n_1544;
assign n_1546 =  n_1167 & ~n_1545;
assign n_1547 = ~n_1539 & ~n_1546;
assign n_1548 = ~n_1165 & ~n_1547;
assign n_1549 = ~n_1167 & ~n_1542;
assign n_1550 =  n_1167 & ~n_1530;
assign n_1551 = ~n_1549 & ~n_1550;
assign n_1552 = ~n_1546 & ~n_1551;
assign n_1553 = ~n_1539 &  n_1552;
assign n_1554 = ~n_1546 & ~n_1553;
assign n_1555 =  n_1165 & ~n_1554;
assign n_1556 = ~n_1548 & ~n_1555;
assign n_1557 = ~n_1163 & ~n_1556;
assign n_1558 = ~n_1165 & ~n_1551;
assign n_1559 =  n_1165 & ~n_1539;
assign n_1560 = ~n_1558 & ~n_1559;
assign n_1561 = ~n_1555 & ~n_1560;
assign n_1562 = ~n_1548 &  n_1561;
assign n_1563 = ~n_1555 & ~n_1562;
assign n_1564 =  n_1163 & ~n_1563;
assign n_1565 = ~n_1557 & ~n_1564;
assign n_1566 = ~n_1161 & ~n_1565;
assign n_1567 = ~n_1163 & ~n_1560;
assign n_1568 =  n_1163 & ~n_1548;
assign n_1569 = ~n_1567 & ~n_1568;
assign n_1570 = ~n_1564 & ~n_1569;
assign n_1571 = ~n_1557 &  n_1570;
assign n_1572 = ~n_1564 & ~n_1571;
assign n_1573 =  n_1161 & ~n_1572;
assign n_1574 = ~n_1566 & ~n_1573;
assign n_1575 = ~n_1159 & ~n_1574;
assign n_1576 = ~n_1161 & ~n_1569;
assign n_1577 =  n_1161 & ~n_1557;
assign n_1578 = ~n_1576 & ~n_1577;
assign n_1579 = ~n_1573 & ~n_1578;
assign n_1580 = ~n_1566 &  n_1579;
assign n_1581 = ~n_1573 & ~n_1580;
assign n_1582 =  n_1159 & ~n_1581;
assign n_1583 = ~n_1575 & ~n_1582;
assign n_1584 = ~n_1157 & ~n_1583;
assign n_1585 = ~n_1159 & ~n_1578;
assign n_1586 =  n_1159 & ~n_1566;
assign n_1587 = ~n_1585 & ~n_1586;
assign n_1588 = ~n_1582 & ~n_1587;
assign n_1589 = ~n_1575 &  n_1588;
assign n_1590 = ~n_1582 & ~n_1589;
assign n_1591 =  n_1157 & ~n_1590;
assign n_1592 = ~n_1584 & ~n_1591;
assign n_1593 = ~n_1155 & ~n_1592;
assign n_1594 = ~n_1157 & ~n_1587;
assign n_1595 =  n_1157 & ~n_1575;
assign n_1596 = ~n_1594 & ~n_1595;
assign n_1597 = ~n_1591 & ~n_1596;
assign n_1598 = ~n_1584 &  n_1597;
assign n_1599 = ~n_1591 & ~n_1598;
assign n_1600 =  n_1155 & ~n_1599;
assign n_1601 = ~n_1593 & ~n_1600;
assign n_1602 = ~n_1153 & ~n_1601;
assign n_1603 = ~n_1155 & ~n_1596;
assign n_1604 =  n_1155 & ~n_1584;
assign n_1605 = ~n_1603 & ~n_1604;
assign n_1606 = ~n_1600 & ~n_1605;
assign n_1607 = ~n_1593 &  n_1606;
assign n_1608 = ~n_1600 & ~n_1607;
assign n_1609 =  n_1153 & ~n_1608;
assign n_1610 = ~n_1602 & ~n_1609;
assign n_1611 = ~n_1151 & ~n_1610;
assign n_1612 = ~n_1153 & ~n_1605;
assign n_1613 =  n_1153 & ~n_1593;
assign n_1614 = ~n_1612 & ~n_1613;
assign n_1615 = ~n_1609 & ~n_1614;
assign n_1616 = ~n_1602 &  n_1615;
assign n_1617 = ~n_1609 & ~n_1616;
assign n_1618 =  n_1151 & ~n_1617;
assign n_1619 = ~n_1611 & ~n_1618;
assign n_1620 = ~n_1149 & ~n_1619;
assign n_1621 = ~n_1151 & ~n_1614;
assign n_1622 =  n_1151 & ~n_1602;
assign n_1623 = ~n_1621 & ~n_1622;
assign n_1624 = ~n_1618 & ~n_1623;
assign n_1625 = ~n_1611 &  n_1624;
assign n_1626 = ~n_1618 & ~n_1625;
assign n_1627 =  n_1149 & ~n_1626;
assign n_1628 = ~n_1620 & ~n_1627;
assign n_1629 = ~n_1147 & ~n_1628;
assign n_1630 = ~n_1149 & ~n_1623;
assign n_1631 =  n_1149 & ~n_1611;
assign n_1632 = ~n_1630 & ~n_1631;
assign n_1633 = ~n_1627 & ~n_1632;
assign n_1634 = ~n_1620 &  n_1633;
assign n_1635 = ~n_1627 & ~n_1634;
assign n_1636 =  n_1147 & ~n_1635;
assign n_1637 = ~n_1629 & ~n_1636;
assign n_1638 = ~n_1145 & ~n_1637;
assign n_1639 = ~n_1147 & ~n_1632;
assign n_1640 =  n_1147 & ~n_1620;
assign n_1641 = ~n_1639 & ~n_1640;
assign n_1642 = ~n_1636 & ~n_1641;
assign n_1643 = ~n_1629 &  n_1642;
assign n_1644 = ~n_1636 & ~n_1643;
assign n_1645 =  n_1145 & ~n_1644;
assign n_1646 = ~n_1638 & ~n_1645;
assign n_1647 = ~n_1143 & ~n_1646;
assign n_1648 = ~n_1145 & ~n_1641;
assign n_1649 =  n_1145 & ~n_1629;
assign n_1650 = ~n_1648 & ~n_1649;
assign n_1651 = ~n_1645 & ~n_1650;
assign n_1652 = ~n_1638 &  n_1651;
assign n_1653 = ~n_1645 & ~n_1652;
assign n_1654 =  n_1143 & ~n_1653;
assign n_1655 = ~n_1647 & ~n_1654;
assign n_1656 = ~n_1141 & ~n_1655;
assign n_1657 = ~n_1143 & ~n_1650;
assign n_1658 =  n_1143 & ~n_1638;
assign n_1659 = ~n_1657 & ~n_1658;
assign n_1660 = ~n_1654 & ~n_1659;
assign n_1661 = ~n_1647 &  n_1660;
assign n_1662 = ~n_1654 & ~n_1661;
assign n_1663 =  n_1141 & ~n_1662;
assign n_1664 = ~n_1656 & ~n_1663;
assign n_1665 = ~n_1139 & ~n_1664;
assign n_1666 = ~n_1141 & ~n_1659;
assign n_1667 =  n_1141 & ~n_1647;
assign n_1668 = ~n_1666 & ~n_1667;
assign n_1669 = ~n_1663 & ~n_1668;
assign n_1670 = ~n_1656 &  n_1669;
assign n_1671 = ~n_1663 & ~n_1670;
assign n_1672 =  n_1139 & ~n_1671;
assign n_1673 = ~n_1665 & ~n_1672;
assign n_1674 = ~n_1137 & ~n_1673;
assign n_1675 = ~n_1139 & ~n_1668;
assign n_1676 =  n_1139 & ~n_1656;
assign n_1677 = ~n_1675 & ~n_1676;
assign n_1678 = ~n_1672 & ~n_1677;
assign n_1679 = ~n_1665 &  n_1678;
assign n_1680 = ~n_1672 & ~n_1679;
assign n_1681 =  n_1137 & ~n_1680;
assign n_1682 = ~n_1674 & ~n_1681;
assign n_1683 = ~n_1135 & ~n_1682;
assign n_1684 = ~n_1137 & ~n_1677;
assign n_1685 =  n_1137 & ~n_1665;
assign n_1686 = ~n_1684 & ~n_1685;
assign n_1687 = ~n_1681 & ~n_1686;
assign n_1688 = ~n_1674 &  n_1687;
assign n_1689 = ~n_1681 & ~n_1688;
assign n_1690 =  n_1135 & ~n_1689;
assign n_1691 = ~n_1683 & ~n_1690;
assign n_1692 = ~n_1133 & ~n_1691;
assign n_1693 = ~n_1135 & ~n_1686;
assign n_1694 =  n_1135 & ~n_1674;
assign n_1695 = ~n_1693 & ~n_1694;
assign n_1696 = ~n_1690 & ~n_1695;
assign n_1697 = ~n_1683 &  n_1696;
assign n_1698 = ~n_1690 & ~n_1697;
assign n_1699 =  n_1133 & ~n_1698;
assign n_1700 = ~n_1692 & ~n_1699;
assign n_1701 = ~n_1131 & ~n_1700;
assign n_1702 = ~n_1133 & ~n_1695;
assign n_1703 =  n_1133 & ~n_1683;
assign n_1704 = ~n_1702 & ~n_1703;
assign n_1705 = ~n_1699 & ~n_1704;
assign n_1706 = ~n_1692 &  n_1705;
assign n_1707 = ~n_1699 & ~n_1706;
assign n_1708 =  n_1131 & ~n_1707;
assign n_1709 = ~n_1701 & ~n_1708;
assign n_1710 = ~n_1129 & ~n_1709;
assign n_1711 = ~n_1131 & ~n_1704;
assign n_1712 =  n_1131 & ~n_1692;
assign n_1713 = ~n_1711 & ~n_1712;
assign n_1714 = ~n_1708 & ~n_1713;
assign n_1715 = ~n_1701 &  n_1714;
assign n_1716 = ~n_1708 & ~n_1715;
assign n_1717 =  n_1129 & ~n_1716;
assign n_1718 = ~n_1710 & ~n_1717;
assign n_1719 = ~n_1127 & ~n_1718;
assign n_1720 = ~n_1129 & ~n_1713;
assign n_1721 =  n_1129 & ~n_1701;
assign n_1722 = ~n_1720 & ~n_1721;
assign n_1723 = ~n_1717 & ~n_1722;
assign n_1724 = ~n_1710 &  n_1723;
assign n_1725 = ~n_1717 & ~n_1724;
assign n_1726 =  n_1127 & ~n_1725;
assign n_1727 = ~n_1719 & ~n_1726;
assign n_1728 = ~n_1125 & ~n_1727;
assign n_1729 = ~n_1127 & ~n_1722;
assign n_1730 =  n_1127 & ~n_1710;
assign n_1731 = ~n_1729 & ~n_1730;
assign n_1732 = ~n_1726 & ~n_1731;
assign n_1733 = ~n_1719 &  n_1732;
assign n_1734 = ~n_1726 & ~n_1733;
assign n_1735 =  n_1125 & ~n_1734;
assign n_1736 = ~n_1728 & ~n_1735;
assign n_1737 = ~n_1123 & ~n_1736;
assign n_1738 = ~n_1125 & ~n_1731;
assign n_1739 =  n_1125 & ~n_1719;
assign n_1740 = ~n_1738 & ~n_1739;
assign n_1741 = ~n_1123 & ~n_1740;
assign n_1742 =  n_1123 & ~n_1728;
assign n_1743 = ~n_1741 & ~n_1742;
assign n_1744 = ~n_1735 & ~n_1740;
assign n_1745 = ~n_1728 &  n_1744;
assign n_1746 = ~n_1735 & ~n_1745;
assign n_1747 =  n_1123 & ~n_1746;
assign n_1748 = ~n_1743 & ~n_1747;
assign n_1749 = ~n_1737 &  n_1748;
assign n_1750 = ~n_588 & ~n_670;
assign n_1751 = ~n_671 & ~n_1750;
assign n_1752 = ~n_1748 & ~n_1751;
assign n_1753 = ~n_1749 & ~n_1752;
assign n_1754 = ~n_1217 & ~n_1318;
assign n_1755 = ~n_1319 & ~n_1754;
assign n_1756 = ~n_1240 & ~n_1248;
assign n_1757 = ~n_1249 & ~n_1756;
assign n_1758 = ~n_1737 & ~n_1747;
assign n_1759 = ~n_1751 & ~n_1758;
assign n_1760 = ~n_1747 & ~n_1749;
assign n_1761 =  n_1751 & ~n_1760;
assign n_1762 = ~n_1759 & ~n_1761;
assign n_1763 = ~n_1757 & ~n_1762;
assign n_1764 = ~n_1743 & ~n_1751;
assign n_1765 = ~n_1737 &  n_1751;
assign n_1766 = ~n_1764 & ~n_1765;
assign n_1767 = ~n_1757 & ~n_1766;
assign n_1768 =  n_1757 & ~n_1759;
assign n_1769 = ~n_1767 & ~n_1768;
assign n_1770 = ~n_1761 & ~n_1766;
assign n_1771 = ~n_1759 &  n_1770;
assign n_1772 = ~n_1761 & ~n_1771;
assign n_1773 =  n_1757 & ~n_1772;
assign n_1774 = ~n_1769 & ~n_1773;
assign n_1775 = ~n_1763 &  n_1774;
assign n_1776 = ~n_601 & ~n_652;
assign n_1777 = ~n_653 & ~n_1776;
assign n_1778 = ~n_1774 & ~n_1777;
assign n_1779 = ~n_1775 & ~n_1778;
assign n_1780 = ~n_1221 & ~n_1300;
assign n_1781 = ~n_1301 & ~n_1780;
assign n_1782 = ~n_634 & ~n_640;
assign n_1783 = ~n_1254 &  n_1260;
assign n_1784 = ~n_1261 & ~n_1783;
assign n_1785 = ~n_1769 & ~n_1777;
assign n_1786 = ~n_1763 &  n_1777;
assign n_1787 = ~n_1785 & ~n_1786;
assign n_1788 = ~n_1784 & ~n_1787;
assign n_1789 = ~n_1763 & ~n_1773;
assign n_1790 = ~n_1777 & ~n_1789;
assign n_1791 =  n_1784 & ~n_1790;
assign n_1792 = ~n_1788 & ~n_1791;
assign n_1793 = ~n_1773 & ~n_1775;
assign n_1794 =  n_1777 & ~n_1793;
assign n_1795 = ~n_1787 & ~n_1794;
assign n_1796 = ~n_1790 &  n_1795;
assign n_1797 = ~n_1794 & ~n_1796;
assign n_1798 =  n_1784 & ~n_1797;
assign n_1799 = ~n_1792 & ~n_1798;
assign n_1800 = ~n_1782 & ~n_1799;
assign n_1801 = ~n_1790 & ~n_1794;
assign n_1802 = ~n_1784 & ~n_1801;
assign n_1803 = ~n_1798 & ~n_1802;
assign n_1804 = ~n_1792 &  n_1803;
assign n_1805 = ~n_1800 & ~n_1804;
assign n_1806 = ~n_1782 & ~n_1792;
assign n_1807 =  n_1782 &  n_1792;
assign n_1808 = ~n_1806 & ~n_1807;
assign n_1809 = ~n_1236 &  n_1275;
assign n_1810 = ~n_1289 & ~n_1809;
assign n_1811 = ~n_1281 &  n_1810;
assign n_1812 = ~n_1808 &  n_1811;
assign n_1813 =  n_1808 & ~n_1811;
assign n_1814 = ~n_1812 & ~n_1813;
assign n_1815 =  n_1805 & ~n_1814;
assign n_1816 = ~n_1805 & ~n_1806;
assign n_1817 = ~n_1815 & ~n_1816;
assign n_1818 = ~n_1781 & ~n_1817;
assign n_1819 = ~n_1805 & ~n_1811;
assign n_1820 =  n_1805 &  n_1811;
assign n_1821 = ~n_1819 & ~n_1820;
assign n_1822 =  n_1814 & ~n_1821;
assign n_1823 =  n_1817 & ~n_1822;
assign n_1824 = ~n_1815 & ~n_1823;
assign n_1825 =  n_1781 & ~n_1824;
assign n_1826 = ~n_1818 & ~n_1825;
assign n_1827 = ~n_1779 & ~n_1826;
assign n_1828 = ~n_1781 &  n_1822;
assign n_1829 =  n_1781 &  n_1816;
assign n_1830 = ~n_1828 & ~n_1829;
assign n_1831 = ~n_1825 &  n_1830;
assign n_1832 = ~n_1818 &  n_1831;
assign n_1833 = ~n_1825 & ~n_1832;
assign n_1834 =  n_1779 & ~n_1833;
assign n_1835 = ~n_1827 & ~n_1834;
assign n_1836 = ~n_1755 & ~n_1835;
assign n_1837 = ~n_1779 & ~n_1830;
assign n_1838 =  n_1779 &  n_1818;
assign n_1839 = ~n_1837 & ~n_1838;
assign n_1840 = ~n_1834 &  n_1839;
assign n_1841 = ~n_1827 &  n_1840;
assign n_1842 = ~n_1834 & ~n_1841;
assign n_1843 =  n_1755 & ~n_1842;
assign n_1844 = ~n_1836 & ~n_1843;
assign n_1845 = ~n_1753 & ~n_1844;
assign n_1846 =  n_1755 & ~n_1827;
assign n_1847 = ~n_1755 &  n_1839;
assign n_1848 = ~n_1846 & ~n_1847;
assign n_1849 = ~n_1843 & ~n_1848;
assign n_1850 = ~n_1836 &  n_1849;
assign n_1851 = ~n_1843 & ~n_1850;
assign n_1852 =  n_1753 & ~n_1851;
assign n_1853 = ~n_1753 & ~n_1848;
assign n_1854 =  n_1753 & ~n_1836;
assign n_1855 = ~n_1853 & ~n_1854;
assign n_1856 = ~n_1852 & ~n_1855;
assign n_1857 = ~n_1845 &  n_1856;
assign n_1858 = ~n_1213 & ~n_1336;
assign n_1859 = ~n_1337 & ~n_1858;
assign n_1860 = ~n_1856 & ~n_1859;
assign n_1861 = ~n_1857 & ~n_1860;
assign n_1862 = ~n_1784 & ~n_1795;
assign n_1863 = ~n_1796 & ~n_1862;
assign n_1864 = ~n_1219 & ~n_1309;
assign n_1865 = ~n_1310 & ~n_1864;
assign n_1866 = ~n_1757 & ~n_1770;
assign n_1867 = ~n_1771 & ~n_1866;
assign n_1868 = ~n_1215 & ~n_1327;
assign n_1869 = ~n_1328 & ~n_1868;
assign n_1870 = ~n_1123 & ~n_1744;
assign n_1871 = ~n_1745 & ~n_1870;
assign n_1872 = ~n_1211 & ~n_1345;
assign n_1873 = ~n_1346 & ~n_1872;
assign n_1874 = ~n_1127 & ~n_1723;
assign n_1875 = ~n_1724 & ~n_1874;
assign n_1876 = ~n_1207 & ~n_1363;
assign n_1877 = ~n_1364 & ~n_1876;
assign n_1878 = ~n_1131 & ~n_1705;
assign n_1879 = ~n_1706 & ~n_1878;
assign n_1880 = ~n_1203 & ~n_1381;
assign n_1881 = ~n_1382 & ~n_1880;
assign n_1882 = ~n_1135 & ~n_1687;
assign n_1883 = ~n_1688 & ~n_1882;
assign n_1884 = ~n_1199 & ~n_1399;
assign n_1885 = ~n_1400 & ~n_1884;
assign n_1886 = ~n_1139 & ~n_1669;
assign n_1887 = ~n_1670 & ~n_1886;
assign n_1888 = ~n_1195 & ~n_1417;
assign n_1889 = ~n_1418 & ~n_1888;
assign n_1890 = ~n_1143 & ~n_1651;
assign n_1891 = ~n_1652 & ~n_1890;
assign n_1892 = ~n_1191 & ~n_1435;
assign n_1893 = ~n_1436 & ~n_1892;
assign n_1894 = ~n_1147 & ~n_1633;
assign n_1895 = ~n_1634 & ~n_1894;
assign n_1896 = ~n_1187 & ~n_1453;
assign n_1897 = ~n_1454 & ~n_1896;
assign n_1898 = ~n_1151 & ~n_1615;
assign n_1899 = ~n_1616 & ~n_1898;
assign n_1900 = ~n_1183 & ~n_1471;
assign n_1901 = ~n_1472 & ~n_1900;
assign n_1902 = ~n_1155 & ~n_1597;
assign n_1903 = ~n_1598 & ~n_1902;
assign n_1904 = ~n_1179 & ~n_1489;
assign n_1905 = ~n_1490 & ~n_1904;
assign n_1906 = ~n_1159 & ~n_1579;
assign n_1907 = ~n_1580 & ~n_1906;
assign n_1908 = ~n_1175 & ~n_1507;
assign n_1909 = ~n_1508 & ~n_1908;
assign n_1910 = ~n_1163 & ~n_1561;
assign n_1911 = ~n_1562 & ~n_1910;
assign n_1912 = ~n_1171 & ~n_1525;
assign n_1913 = ~n_1526 & ~n_1912;
assign n_1914 = ~n_1167 & ~n_1543;
assign n_1915 = ~n_1544 & ~n_1914;
assign n_1916 = ~n_1169 & ~n_1534;
assign n_1917 = ~n_1535 & ~n_1916;
assign n_1918 = ~n_1165 & ~n_1552;
assign n_1919 = ~n_1553 & ~n_1918;
assign n_1920 = ~n_1173 & ~n_1516;
assign n_1921 = ~n_1517 & ~n_1920;
assign n_1922 = ~n_1161 & ~n_1570;
assign n_1923 = ~n_1571 & ~n_1922;
assign n_1924 = ~n_1177 & ~n_1498;
assign n_1925 = ~n_1499 & ~n_1924;
assign n_1926 = ~n_1157 & ~n_1588;
assign n_1927 = ~n_1589 & ~n_1926;
assign n_1928 = ~n_1181 & ~n_1480;
assign n_1929 = ~n_1481 & ~n_1928;
assign n_1930 = ~n_1153 & ~n_1606;
assign n_1931 = ~n_1607 & ~n_1930;
assign n_1932 = ~n_1185 & ~n_1462;
assign n_1933 = ~n_1463 & ~n_1932;
assign n_1934 = ~n_1149 & ~n_1624;
assign n_1935 = ~n_1625 & ~n_1934;
assign n_1936 = ~n_1189 & ~n_1444;
assign n_1937 = ~n_1445 & ~n_1936;
assign n_1938 = ~n_1145 & ~n_1642;
assign n_1939 = ~n_1643 & ~n_1938;
assign n_1940 = ~n_1193 & ~n_1426;
assign n_1941 = ~n_1427 & ~n_1940;
assign n_1942 = ~n_1141 & ~n_1660;
assign n_1943 = ~n_1661 & ~n_1942;
assign n_1944 = ~n_1197 & ~n_1408;
assign n_1945 = ~n_1409 & ~n_1944;
assign n_1946 = ~n_1137 & ~n_1678;
assign n_1947 = ~n_1679 & ~n_1946;
assign n_1948 = ~n_1201 & ~n_1390;
assign n_1949 = ~n_1391 & ~n_1948;
assign n_1950 = ~n_1133 & ~n_1696;
assign n_1951 = ~n_1697 & ~n_1950;
assign n_1952 = ~n_1205 & ~n_1372;
assign n_1953 = ~n_1373 & ~n_1952;
assign n_1954 = ~n_1129 & ~n_1714;
assign n_1955 = ~n_1715 & ~n_1954;
assign n_1956 = ~n_1209 & ~n_1354;
assign n_1957 = ~n_1355 & ~n_1956;
assign n_1958 = ~n_1125 & ~n_1732;
assign n_1959 = ~n_1733 & ~n_1958;
assign n_1960 = ~n_1845 & ~n_1852;
assign n_1961 = ~n_1859 & ~n_1960;
assign n_1962 = ~n_1852 & ~n_1857;
assign n_1963 =  n_1859 & ~n_1962;
assign n_1964 = ~n_1961 & ~n_1963;
assign n_1965 = ~n_1959 & ~n_1964;
assign n_1966 = ~n_1855 & ~n_1859;
assign n_1967 = ~n_1845 &  n_1859;
assign n_1968 = ~n_1966 & ~n_1967;
assign n_1969 = ~n_1963 & ~n_1968;
assign n_1970 = ~n_1961 &  n_1969;
assign n_1971 = ~n_1963 & ~n_1970;
assign n_1972 =  n_1959 & ~n_1971;
assign n_1973 = ~n_1965 & ~n_1972;
assign n_1974 = ~n_1957 & ~n_1973;
assign n_1975 = ~n_1959 & ~n_1968;
assign n_1976 =  n_1959 & ~n_1961;
assign n_1977 = ~n_1975 & ~n_1976;
assign n_1978 = ~n_1972 & ~n_1977;
assign n_1979 = ~n_1965 &  n_1978;
assign n_1980 = ~n_1972 & ~n_1979;
assign n_1981 =  n_1957 & ~n_1980;
assign n_1982 = ~n_1974 & ~n_1981;
assign n_1983 = ~n_1955 & ~n_1982;
assign n_1984 = ~n_1957 & ~n_1977;
assign n_1985 =  n_1957 & ~n_1965;
assign n_1986 = ~n_1984 & ~n_1985;
assign n_1987 = ~n_1981 & ~n_1986;
assign n_1988 = ~n_1974 &  n_1987;
assign n_1989 = ~n_1981 & ~n_1988;
assign n_1990 =  n_1955 & ~n_1989;
assign n_1991 = ~n_1983 & ~n_1990;
assign n_1992 = ~n_1953 & ~n_1991;
assign n_1993 = ~n_1955 & ~n_1986;
assign n_1994 =  n_1955 & ~n_1974;
assign n_1995 = ~n_1993 & ~n_1994;
assign n_1996 = ~n_1990 & ~n_1995;
assign n_1997 = ~n_1983 &  n_1996;
assign n_1998 = ~n_1990 & ~n_1997;
assign n_1999 =  n_1953 & ~n_1998;
assign n_2000 = ~n_1992 & ~n_1999;
assign n_2001 = ~n_1951 & ~n_2000;
assign n_2002 = ~n_1953 & ~n_1995;
assign n_2003 =  n_1953 & ~n_1983;
assign n_2004 = ~n_2002 & ~n_2003;
assign n_2005 = ~n_1999 & ~n_2004;
assign n_2006 = ~n_1992 &  n_2005;
assign n_2007 = ~n_1999 & ~n_2006;
assign n_2008 =  n_1951 & ~n_2007;
assign n_2009 = ~n_2001 & ~n_2008;
assign n_2010 = ~n_1949 & ~n_2009;
assign n_2011 = ~n_1951 & ~n_2004;
assign n_2012 =  n_1951 & ~n_1992;
assign n_2013 = ~n_2011 & ~n_2012;
assign n_2014 = ~n_2008 & ~n_2013;
assign n_2015 = ~n_2001 &  n_2014;
assign n_2016 = ~n_2008 & ~n_2015;
assign n_2017 =  n_1949 & ~n_2016;
assign n_2018 = ~n_2010 & ~n_2017;
assign n_2019 = ~n_1947 & ~n_2018;
assign n_2020 = ~n_1949 & ~n_2013;
assign n_2021 =  n_1949 & ~n_2001;
assign n_2022 = ~n_2020 & ~n_2021;
assign n_2023 = ~n_2017 & ~n_2022;
assign n_2024 = ~n_2010 &  n_2023;
assign n_2025 = ~n_2017 & ~n_2024;
assign n_2026 =  n_1947 & ~n_2025;
assign n_2027 = ~n_2019 & ~n_2026;
assign n_2028 = ~n_1945 & ~n_2027;
assign n_2029 = ~n_1947 & ~n_2022;
assign n_2030 =  n_1947 & ~n_2010;
assign n_2031 = ~n_2029 & ~n_2030;
assign n_2032 = ~n_2026 & ~n_2031;
assign n_2033 = ~n_2019 &  n_2032;
assign n_2034 = ~n_2026 & ~n_2033;
assign n_2035 =  n_1945 & ~n_2034;
assign n_2036 = ~n_2028 & ~n_2035;
assign n_2037 = ~n_1943 & ~n_2036;
assign n_2038 = ~n_1945 & ~n_2031;
assign n_2039 =  n_1945 & ~n_2019;
assign n_2040 = ~n_2038 & ~n_2039;
assign n_2041 = ~n_2035 & ~n_2040;
assign n_2042 = ~n_2028 &  n_2041;
assign n_2043 = ~n_2035 & ~n_2042;
assign n_2044 =  n_1943 & ~n_2043;
assign n_2045 = ~n_2037 & ~n_2044;
assign n_2046 = ~n_1941 & ~n_2045;
assign n_2047 = ~n_1943 & ~n_2040;
assign n_2048 =  n_1943 & ~n_2028;
assign n_2049 = ~n_2047 & ~n_2048;
assign n_2050 = ~n_2044 & ~n_2049;
assign n_2051 = ~n_2037 &  n_2050;
assign n_2052 = ~n_2044 & ~n_2051;
assign n_2053 =  n_1941 & ~n_2052;
assign n_2054 = ~n_2046 & ~n_2053;
assign n_2055 = ~n_1939 & ~n_2054;
assign n_2056 = ~n_1941 & ~n_2049;
assign n_2057 =  n_1941 & ~n_2037;
assign n_2058 = ~n_2056 & ~n_2057;
assign n_2059 = ~n_2053 & ~n_2058;
assign n_2060 = ~n_2046 &  n_2059;
assign n_2061 = ~n_2053 & ~n_2060;
assign n_2062 =  n_1939 & ~n_2061;
assign n_2063 = ~n_2055 & ~n_2062;
assign n_2064 = ~n_1937 & ~n_2063;
assign n_2065 = ~n_1939 & ~n_2058;
assign n_2066 =  n_1939 & ~n_2046;
assign n_2067 = ~n_2065 & ~n_2066;
assign n_2068 = ~n_2062 & ~n_2067;
assign n_2069 = ~n_2055 &  n_2068;
assign n_2070 = ~n_2062 & ~n_2069;
assign n_2071 =  n_1937 & ~n_2070;
assign n_2072 = ~n_2064 & ~n_2071;
assign n_2073 = ~n_1935 & ~n_2072;
assign n_2074 = ~n_1937 & ~n_2067;
assign n_2075 =  n_1937 & ~n_2055;
assign n_2076 = ~n_2074 & ~n_2075;
assign n_2077 = ~n_2071 & ~n_2076;
assign n_2078 = ~n_2064 &  n_2077;
assign n_2079 = ~n_2071 & ~n_2078;
assign n_2080 =  n_1935 & ~n_2079;
assign n_2081 = ~n_2073 & ~n_2080;
assign n_2082 = ~n_1933 & ~n_2081;
assign n_2083 = ~n_1935 & ~n_2076;
assign n_2084 =  n_1935 & ~n_2064;
assign n_2085 = ~n_2083 & ~n_2084;
assign n_2086 = ~n_2080 & ~n_2085;
assign n_2087 = ~n_2073 &  n_2086;
assign n_2088 = ~n_2080 & ~n_2087;
assign n_2089 =  n_1933 & ~n_2088;
assign n_2090 = ~n_2082 & ~n_2089;
assign n_2091 = ~n_1931 & ~n_2090;
assign n_2092 = ~n_1933 & ~n_2085;
assign n_2093 =  n_1933 & ~n_2073;
assign n_2094 = ~n_2092 & ~n_2093;
assign n_2095 = ~n_2089 & ~n_2094;
assign n_2096 = ~n_2082 &  n_2095;
assign n_2097 = ~n_2089 & ~n_2096;
assign n_2098 =  n_1931 & ~n_2097;
assign n_2099 = ~n_2091 & ~n_2098;
assign n_2100 = ~n_1929 & ~n_2099;
assign n_2101 = ~n_1931 & ~n_2094;
assign n_2102 =  n_1931 & ~n_2082;
assign n_2103 = ~n_2101 & ~n_2102;
assign n_2104 = ~n_2098 & ~n_2103;
assign n_2105 = ~n_2091 &  n_2104;
assign n_2106 = ~n_2098 & ~n_2105;
assign n_2107 =  n_1929 & ~n_2106;
assign n_2108 = ~n_2100 & ~n_2107;
assign n_2109 = ~n_1927 & ~n_2108;
assign n_2110 = ~n_1929 & ~n_2103;
assign n_2111 =  n_1929 & ~n_2091;
assign n_2112 = ~n_2110 & ~n_2111;
assign n_2113 = ~n_2107 & ~n_2112;
assign n_2114 = ~n_2100 &  n_2113;
assign n_2115 = ~n_2107 & ~n_2114;
assign n_2116 =  n_1927 & ~n_2115;
assign n_2117 = ~n_2109 & ~n_2116;
assign n_2118 = ~n_1925 & ~n_2117;
assign n_2119 = ~n_1927 & ~n_2112;
assign n_2120 =  n_1927 & ~n_2100;
assign n_2121 = ~n_2119 & ~n_2120;
assign n_2122 = ~n_2116 & ~n_2121;
assign n_2123 = ~n_2109 &  n_2122;
assign n_2124 = ~n_2116 & ~n_2123;
assign n_2125 =  n_1925 & ~n_2124;
assign n_2126 = ~n_2118 & ~n_2125;
assign n_2127 = ~n_1923 & ~n_2126;
assign n_2128 = ~n_1925 & ~n_2121;
assign n_2129 =  n_1925 & ~n_2109;
assign n_2130 = ~n_2128 & ~n_2129;
assign n_2131 = ~n_2125 & ~n_2130;
assign n_2132 = ~n_2118 &  n_2131;
assign n_2133 = ~n_2125 & ~n_2132;
assign n_2134 =  n_1923 & ~n_2133;
assign n_2135 = ~n_2127 & ~n_2134;
assign n_2136 = ~n_1921 & ~n_2135;
assign n_2137 = ~n_1923 & ~n_2130;
assign n_2138 =  n_1923 & ~n_2118;
assign n_2139 = ~n_2137 & ~n_2138;
assign n_2140 = ~n_2134 & ~n_2139;
assign n_2141 = ~n_2127 &  n_2140;
assign n_2142 = ~n_2134 & ~n_2141;
assign n_2143 =  n_1921 & ~n_2142;
assign n_2144 = ~n_2136 & ~n_2143;
assign n_2145 = ~n_1919 & ~n_2144;
assign n_2146 = ~n_1921 & ~n_2139;
assign n_2147 =  n_1921 & ~n_2127;
assign n_2148 = ~n_2146 & ~n_2147;
assign n_2149 = ~n_2143 & ~n_2148;
assign n_2150 = ~n_2136 &  n_2149;
assign n_2151 = ~n_2143 & ~n_2150;
assign n_2152 =  n_1919 & ~n_2151;
assign n_2153 = ~n_2145 & ~n_2152;
assign n_2154 = ~n_1917 & ~n_2153;
assign n_2155 = ~n_1919 & ~n_2148;
assign n_2156 =  n_1919 & ~n_2136;
assign n_2157 = ~n_2155 & ~n_2156;
assign n_2158 = ~n_2152 & ~n_2157;
assign n_2159 = ~n_2145 &  n_2158;
assign n_2160 = ~n_2152 & ~n_2159;
assign n_2161 =  n_1917 & ~n_2160;
assign n_2162 = ~n_2154 & ~n_2161;
assign n_2163 = ~n_1915 & ~n_2162;
assign n_2164 = ~n_1917 & ~n_2157;
assign n_2165 =  n_1917 & ~n_2145;
assign n_2166 = ~n_2164 & ~n_2165;
assign n_2167 = ~n_2161 & ~n_2166;
assign n_2168 = ~n_2154 &  n_2167;
assign n_2169 = ~n_2161 & ~n_2168;
assign n_2170 =  n_1915 & ~n_2169;
assign n_2171 = ~n_2163 & ~n_2170;
assign n_2172 = ~n_1913 & ~n_2171;
assign n_2173 = ~n_1915 & ~n_2166;
assign n_2174 =  n_1915 & ~n_2154;
assign n_2175 = ~n_2173 & ~n_2174;
assign n_2176 = ~n_2170 & ~n_2175;
assign n_2177 = ~n_2163 &  n_2176;
assign n_2178 = ~n_2170 & ~n_2177;
assign n_2179 =  n_1913 & ~n_2178;
assign n_2180 = ~n_2172 & ~n_2179;
assign n_2181 = ~n_1911 & ~n_2180;
assign n_2182 = ~n_1913 & ~n_2175;
assign n_2183 =  n_1913 & ~n_2163;
assign n_2184 = ~n_2182 & ~n_2183;
assign n_2185 = ~n_2179 & ~n_2184;
assign n_2186 = ~n_2172 &  n_2185;
assign n_2187 = ~n_2179 & ~n_2186;
assign n_2188 =  n_1911 & ~n_2187;
assign n_2189 = ~n_2181 & ~n_2188;
assign n_2190 = ~n_1909 & ~n_2189;
assign n_2191 = ~n_1911 & ~n_2184;
assign n_2192 =  n_1911 & ~n_2172;
assign n_2193 = ~n_2191 & ~n_2192;
assign n_2194 = ~n_2188 & ~n_2193;
assign n_2195 = ~n_2181 &  n_2194;
assign n_2196 = ~n_2188 & ~n_2195;
assign n_2197 =  n_1909 & ~n_2196;
assign n_2198 = ~n_2190 & ~n_2197;
assign n_2199 = ~n_1907 & ~n_2198;
assign n_2200 = ~n_1909 & ~n_2193;
assign n_2201 =  n_1909 & ~n_2181;
assign n_2202 = ~n_2200 & ~n_2201;
assign n_2203 = ~n_2197 & ~n_2202;
assign n_2204 = ~n_2190 &  n_2203;
assign n_2205 = ~n_2197 & ~n_2204;
assign n_2206 =  n_1907 & ~n_2205;
assign n_2207 = ~n_2199 & ~n_2206;
assign n_2208 = ~n_1905 & ~n_2207;
assign n_2209 = ~n_1907 & ~n_2202;
assign n_2210 =  n_1907 & ~n_2190;
assign n_2211 = ~n_2209 & ~n_2210;
assign n_2212 = ~n_2206 & ~n_2211;
assign n_2213 = ~n_2199 &  n_2212;
assign n_2214 = ~n_2206 & ~n_2213;
assign n_2215 =  n_1905 & ~n_2214;
assign n_2216 = ~n_2208 & ~n_2215;
assign n_2217 = ~n_1903 & ~n_2216;
assign n_2218 = ~n_1905 & ~n_2211;
assign n_2219 =  n_1905 & ~n_2199;
assign n_2220 = ~n_2218 & ~n_2219;
assign n_2221 = ~n_2215 & ~n_2220;
assign n_2222 = ~n_2208 &  n_2221;
assign n_2223 = ~n_2215 & ~n_2222;
assign n_2224 =  n_1903 & ~n_2223;
assign n_2225 = ~n_2217 & ~n_2224;
assign n_2226 = ~n_1901 & ~n_2225;
assign n_2227 = ~n_1903 & ~n_2220;
assign n_2228 =  n_1903 & ~n_2208;
assign n_2229 = ~n_2227 & ~n_2228;
assign n_2230 = ~n_2224 & ~n_2229;
assign n_2231 = ~n_2217 &  n_2230;
assign n_2232 = ~n_2224 & ~n_2231;
assign n_2233 =  n_1901 & ~n_2232;
assign n_2234 = ~n_2226 & ~n_2233;
assign n_2235 = ~n_1899 & ~n_2234;
assign n_2236 = ~n_1901 & ~n_2229;
assign n_2237 =  n_1901 & ~n_2217;
assign n_2238 = ~n_2236 & ~n_2237;
assign n_2239 = ~n_2233 & ~n_2238;
assign n_2240 = ~n_2226 &  n_2239;
assign n_2241 = ~n_2233 & ~n_2240;
assign n_2242 =  n_1899 & ~n_2241;
assign n_2243 = ~n_2235 & ~n_2242;
assign n_2244 = ~n_1897 & ~n_2243;
assign n_2245 = ~n_1899 & ~n_2238;
assign n_2246 =  n_1899 & ~n_2226;
assign n_2247 = ~n_2245 & ~n_2246;
assign n_2248 = ~n_2242 & ~n_2247;
assign n_2249 = ~n_2235 &  n_2248;
assign n_2250 = ~n_2242 & ~n_2249;
assign n_2251 =  n_1897 & ~n_2250;
assign n_2252 = ~n_2244 & ~n_2251;
assign n_2253 = ~n_1895 & ~n_2252;
assign n_2254 = ~n_1897 & ~n_2247;
assign n_2255 =  n_1897 & ~n_2235;
assign n_2256 = ~n_2254 & ~n_2255;
assign n_2257 = ~n_2251 & ~n_2256;
assign n_2258 = ~n_2244 &  n_2257;
assign n_2259 = ~n_2251 & ~n_2258;
assign n_2260 =  n_1895 & ~n_2259;
assign n_2261 = ~n_2253 & ~n_2260;
assign n_2262 = ~n_1893 & ~n_2261;
assign n_2263 = ~n_1895 & ~n_2256;
assign n_2264 =  n_1895 & ~n_2244;
assign n_2265 = ~n_2263 & ~n_2264;
assign n_2266 = ~n_2260 & ~n_2265;
assign n_2267 = ~n_2253 &  n_2266;
assign n_2268 = ~n_2260 & ~n_2267;
assign n_2269 =  n_1893 & ~n_2268;
assign n_2270 = ~n_2262 & ~n_2269;
assign n_2271 = ~n_1891 & ~n_2270;
assign n_2272 = ~n_1893 & ~n_2265;
assign n_2273 =  n_1893 & ~n_2253;
assign n_2274 = ~n_2272 & ~n_2273;
assign n_2275 = ~n_2269 & ~n_2274;
assign n_2276 = ~n_2262 &  n_2275;
assign n_2277 = ~n_2269 & ~n_2276;
assign n_2278 =  n_1891 & ~n_2277;
assign n_2279 = ~n_2271 & ~n_2278;
assign n_2280 = ~n_1889 & ~n_2279;
assign n_2281 = ~n_1891 & ~n_2274;
assign n_2282 =  n_1891 & ~n_2262;
assign n_2283 = ~n_2281 & ~n_2282;
assign n_2284 = ~n_2278 & ~n_2283;
assign n_2285 = ~n_2271 &  n_2284;
assign n_2286 = ~n_2278 & ~n_2285;
assign n_2287 =  n_1889 & ~n_2286;
assign n_2288 = ~n_2280 & ~n_2287;
assign n_2289 = ~n_1887 & ~n_2288;
assign n_2290 = ~n_1889 & ~n_2283;
assign n_2291 =  n_1889 & ~n_2271;
assign n_2292 = ~n_2290 & ~n_2291;
assign n_2293 = ~n_2287 & ~n_2292;
assign n_2294 = ~n_2280 &  n_2293;
assign n_2295 = ~n_2287 & ~n_2294;
assign n_2296 =  n_1887 & ~n_2295;
assign n_2297 = ~n_2289 & ~n_2296;
assign n_2298 = ~n_1885 & ~n_2297;
assign n_2299 = ~n_1887 & ~n_2292;
assign n_2300 =  n_1887 & ~n_2280;
assign n_2301 = ~n_2299 & ~n_2300;
assign n_2302 = ~n_2296 & ~n_2301;
assign n_2303 = ~n_2289 &  n_2302;
assign n_2304 = ~n_2296 & ~n_2303;
assign n_2305 =  n_1885 & ~n_2304;
assign n_2306 = ~n_2298 & ~n_2305;
assign n_2307 = ~n_1883 & ~n_2306;
assign n_2308 = ~n_1885 & ~n_2301;
assign n_2309 =  n_1885 & ~n_2289;
assign n_2310 = ~n_2308 & ~n_2309;
assign n_2311 = ~n_2305 & ~n_2310;
assign n_2312 = ~n_2298 &  n_2311;
assign n_2313 = ~n_2305 & ~n_2312;
assign n_2314 =  n_1883 & ~n_2313;
assign n_2315 = ~n_2307 & ~n_2314;
assign n_2316 = ~n_1881 & ~n_2315;
assign n_2317 = ~n_1883 & ~n_2310;
assign n_2318 =  n_1883 & ~n_2298;
assign n_2319 = ~n_2317 & ~n_2318;
assign n_2320 = ~n_2314 & ~n_2319;
assign n_2321 = ~n_2307 &  n_2320;
assign n_2322 = ~n_2314 & ~n_2321;
assign n_2323 =  n_1881 & ~n_2322;
assign n_2324 = ~n_2316 & ~n_2323;
assign n_2325 = ~n_1879 & ~n_2324;
assign n_2326 = ~n_1881 & ~n_2319;
assign n_2327 =  n_1881 & ~n_2307;
assign n_2328 = ~n_2326 & ~n_2327;
assign n_2329 = ~n_2323 & ~n_2328;
assign n_2330 = ~n_2316 &  n_2329;
assign n_2331 = ~n_2323 & ~n_2330;
assign n_2332 =  n_1879 & ~n_2331;
assign n_2333 = ~n_2325 & ~n_2332;
assign n_2334 = ~n_1877 & ~n_2333;
assign n_2335 = ~n_1879 & ~n_2328;
assign n_2336 =  n_1879 & ~n_2316;
assign n_2337 = ~n_2335 & ~n_2336;
assign n_2338 = ~n_2332 & ~n_2337;
assign n_2339 = ~n_2325 &  n_2338;
assign n_2340 = ~n_2332 & ~n_2339;
assign n_2341 =  n_1877 & ~n_2340;
assign n_2342 = ~n_2334 & ~n_2341;
assign n_2343 = ~n_1875 & ~n_2342;
assign n_2344 = ~n_1877 & ~n_2337;
assign n_2345 =  n_1877 & ~n_2325;
assign n_2346 = ~n_2344 & ~n_2345;
assign n_2347 = ~n_2341 & ~n_2346;
assign n_2348 = ~n_2334 &  n_2347;
assign n_2349 = ~n_2341 & ~n_2348;
assign n_2350 =  n_1875 & ~n_2349;
assign n_2351 = ~n_2343 & ~n_2350;
assign n_2352 = ~n_1873 & ~n_2351;
assign n_2353 = ~n_1875 & ~n_2346;
assign n_2354 =  n_1875 & ~n_2334;
assign n_2355 = ~n_2353 & ~n_2354;
assign n_2356 = ~n_2350 & ~n_2355;
assign n_2357 = ~n_2343 &  n_2356;
assign n_2358 = ~n_2350 & ~n_2357;
assign n_2359 =  n_1873 & ~n_2358;
assign n_2360 = ~n_2352 & ~n_2359;
assign n_2361 = ~n_1871 & ~n_2360;
assign n_2362 = ~n_1873 & ~n_2355;
assign n_2363 =  n_1873 & ~n_2343;
assign n_2364 = ~n_2362 & ~n_2363;
assign n_2365 = ~n_2359 & ~n_2364;
assign n_2366 = ~n_2352 &  n_2365;
assign n_2367 = ~n_2359 & ~n_2366;
assign n_2368 =  n_1871 & ~n_2367;
assign n_2369 = ~n_2361 & ~n_2368;
assign n_2370 = ~n_1869 & ~n_2369;
assign n_2371 = ~n_1871 & ~n_2364;
assign n_2372 =  n_1871 & ~n_2352;
assign n_2373 = ~n_2371 & ~n_2372;
assign n_2374 = ~n_2368 & ~n_2373;
assign n_2375 = ~n_2361 &  n_2374;
assign n_2376 = ~n_2368 & ~n_2375;
assign n_2377 =  n_1869 & ~n_2376;
assign n_2378 = ~n_2370 & ~n_2377;
assign n_2379 = ~n_1867 & ~n_2378;
assign n_2380 = ~n_1869 & ~n_2373;
assign n_2381 =  n_1869 & ~n_2361;
assign n_2382 = ~n_2380 & ~n_2381;
assign n_2383 = ~n_2377 & ~n_2382;
assign n_2384 = ~n_2370 &  n_2383;
assign n_2385 = ~n_2377 & ~n_2384;
assign n_2386 =  n_1867 & ~n_2385;
assign n_2387 = ~n_2379 & ~n_2386;
assign n_2388 = ~n_1865 & ~n_2387;
assign n_2389 = ~n_1867 & ~n_2382;
assign n_2390 =  n_1867 & ~n_2370;
assign n_2391 = ~n_2389 & ~n_2390;
assign n_2392 = ~n_2386 & ~n_2391;
assign n_2393 = ~n_2379 &  n_2392;
assign n_2394 = ~n_2386 & ~n_2393;
assign n_2395 =  n_1865 & ~n_2394;
assign n_2396 = ~n_2388 & ~n_2395;
assign n_2397 = ~n_1863 & ~n_2396;
assign n_2398 = ~n_1865 & ~n_2391;
assign n_2399 =  n_1865 & ~n_2379;
assign n_2400 = ~n_2398 & ~n_2399;
assign n_2401 = ~n_2395 & ~n_2400;
assign n_2402 = ~n_2388 &  n_2401;
assign n_2403 = ~n_2395 & ~n_2402;
assign n_2404 =  n_1863 & ~n_2403;
assign n_2405 = ~n_1863 & ~n_2400;
assign n_2406 =  n_1863 & ~n_2388;
assign n_2407 = ~n_2405 & ~n_2406;
assign n_2408 = ~n_2404 & ~n_2407;
assign n_2409 = ~n_2397 &  n_2408;
assign n_2410 = ~n_1234 & ~n_1291;
assign n_2411 = ~n_1292 & ~n_2410;
assign n_2412 = ~n_2408 & ~n_2411;
assign n_2413 = ~n_2409 & ~n_2412;
assign n_2414 = ~n_1755 & ~n_1840;
assign n_2415 = ~n_1841 & ~n_2414;
assign n_2416 = ~n_1270 & ~n_1278;
assign n_2417 =  n_1782 &  n_1799;
assign n_2418 = ~n_1802 &  n_2417;
assign n_2419 = ~n_1803 & ~n_2417;
assign n_2420 = ~n_2418 & ~n_2419;
assign n_2421 = ~n_2404 & ~n_2409;
assign n_2422 =  n_2411 & ~n_2421;
assign n_2423 = ~n_2397 & ~n_2404;
assign n_2424 = ~n_2411 & ~n_2423;
assign n_2425 = ~n_2407 & ~n_2411;
assign n_2426 = ~n_2397 &  n_2411;
assign n_2427 = ~n_2425 & ~n_2426;
assign n_2428 = ~n_2422 & ~n_2427;
assign n_2429 = ~n_2424 &  n_2428;
assign n_2430 = ~n_2422 & ~n_2429;
assign n_2431 =  n_2420 & ~n_2430;
assign n_2432 = ~n_2416 &  n_2431;
assign n_2433 = ~n_2422 & ~n_2424;
assign n_2434 = ~n_2420 & ~n_2433;
assign n_2435 = ~n_2431 & ~n_2434;
assign n_2436 = ~n_2420 & ~n_2427;
assign n_2437 =  n_2420 & ~n_2424;
assign n_2438 = ~n_2436 & ~n_2437;
assign n_2439 =  n_2435 & ~n_2438;
assign n_2440 = ~n_2416 &  n_2438;
assign n_2441 = ~n_2439 & ~n_2440;
assign n_2442 = ~n_2432 &  n_2441;
assign n_2443 = ~n_2431 & ~n_2439;
assign n_2444 =  n_2416 & ~n_2443;
assign n_2445 =  n_2416 &  n_2434;
assign n_2446 = ~n_2440 & ~n_2445;
assign n_2447 = ~n_2444 &  n_2446;
assign n_2448 = ~n_1815 & ~n_1822;
assign n_2449 = ~n_1781 & ~n_2448;
assign n_2450 = ~n_1823 & ~n_2449;
assign n_2451 = ~n_2447 & ~n_2450;
assign n_2452 =  n_2447 &  n_2450;
assign n_2453 = ~n_2451 & ~n_2452;
assign n_2454 =  n_2442 & ~n_2453;
assign n_2455 = ~n_2442 & ~n_2447;
assign n_2456 = ~n_2454 & ~n_2455;
assign n_2457 = ~n_2442 & ~n_2450;
assign n_2458 =  n_2447 & ~n_2457;
assign n_2459 = ~n_2451 & ~n_2455;
assign n_2460 = ~n_2458 &  n_2459;
assign n_2461 =  n_2456 & ~n_2460;
assign n_2462 = ~n_2454 & ~n_2461;
assign n_2463 =  n_2415 & ~n_2462;
assign n_2464 = ~n_2415 & ~n_2456;
assign n_2465 = ~n_2463 & ~n_2464;
assign n_2466 = ~n_2415 & ~n_2460;
assign n_2467 =  n_2415 & ~n_2455;
assign n_2468 = ~n_2466 & ~n_2467;
assign n_2469 =  n_2465 & ~n_2468;
assign n_2470 = ~n_2463 & ~n_2469;
assign n_2471 =  n_2413 & ~n_2470;
assign n_2472 = ~n_1861 &  n_2471;
assign n_2473 = ~n_2413 & ~n_2465;
assign n_2474 = ~n_2471 & ~n_2473;
assign n_2475 = ~n_2413 &  n_2468;
assign n_2476 =  n_2413 &  n_2464;
assign n_2477 = ~n_2475 & ~n_2476;
assign n_2478 =  n_2474 &  n_2477;
assign n_2479 = ~n_1861 & ~n_2477;
assign n_2480 = ~n_2478 & ~n_2479;
assign n_2481 = ~n_2472 &  n_2480;
assign n_2482 = ~n_1865 & ~n_2392;
assign n_2483 = ~n_2393 & ~n_2482;
assign n_2484 = ~n_2471 & ~n_2478;
assign n_2485 =  n_1861 & ~n_2484;
assign n_2486 = ~n_2483 &  n_2485;
assign n_2487 = ~n_1861 & ~n_2474;
assign n_2488 = ~n_2485 & ~n_2487;
assign n_2489 =  n_1861 &  n_2473;
assign n_2490 = ~n_2479 & ~n_2489;
assign n_2491 =  n_2488 &  n_2490;
assign n_2492 = ~n_2483 & ~n_2490;
assign n_2493 = ~n_2491 & ~n_2492;
assign n_2494 = ~n_2486 &  n_2493;
assign n_2495 = ~x_80 & ~x_81;
assign n_2496 = ~x_82 & ~x_83;
assign n_2497 =  n_2495 &  n_2496;
assign n_2498 = ~x_76 & ~x_77;
assign n_2499 = ~x_78 & ~x_79;
assign n_2500 =  n_2498 &  n_2499;
assign n_2501 =  n_2497 &  n_2500;
assign n_2502 = ~x_88 & ~x_89;
assign n_2503 = ~x_90 & ~x_91;
assign n_2504 =  n_2502 &  n_2503;
assign n_2505 = ~x_84 & ~x_85;
assign n_2506 = ~x_86 & ~x_87;
assign n_2507 =  n_2505 &  n_2506;
assign n_2508 =  n_2504 &  n_2507;
assign n_2509 =  n_2501 &  n_2508;
assign n_2510 = ~x_64 & ~x_65;
assign n_2511 = ~x_66 & ~x_67;
assign n_2512 =  n_2510 &  n_2511;
assign n_2513 = ~x_62 & ~x_63;
assign n_2514 =  n_2 &  n_2513;
assign n_2515 =  n_2512 &  n_2514;
assign n_2516 = ~x_72 & ~x_73;
assign n_2517 = ~x_74 & ~x_75;
assign n_2518 =  n_2516 &  n_2517;
assign n_2519 = ~x_68 & ~x_69;
assign n_2520 = ~x_70 & ~x_71;
assign n_2521 =  n_2519 &  n_2520;
assign n_2522 =  n_2518 &  n_2521;
assign n_2523 =  n_2515 &  n_2522;
assign n_2524 =  n_2509 &  n_2523;
assign n_2525 = ~x_116 & ~x_117;
assign n_2526 = ~x_118 & ~x_120;
assign n_2527 =  n_2525 &  n_2526;
assign n_2528 = ~x_112 & ~x_113;
assign n_2529 = ~x_114 & ~x_115;
assign n_2530 =  n_2528 &  n_2529;
assign n_2531 = ~x_108 & ~x_109;
assign n_2532 = ~x_110 & ~x_111;
assign n_2533 =  n_2531 &  n_2532;
assign n_2534 =  n_2530 &  n_2533;
assign n_2535 =  n_2527 &  n_2534;
assign n_2536 = ~x_96 & ~x_97;
assign n_2537 = ~x_98 & ~x_99;
assign n_2538 =  n_2536 &  n_2537;
assign n_2539 = ~x_92 & ~x_93;
assign n_2540 = ~x_94 & ~x_95;
assign n_2541 =  n_2539 &  n_2540;
assign n_2542 =  n_2538 &  n_2541;
assign n_2543 = ~x_104 & ~x_105;
assign n_2544 = ~x_106 & ~x_107;
assign n_2545 =  n_2543 &  n_2544;
assign n_2546 = ~x_100 & ~x_101;
assign n_2547 = ~x_102 & ~x_103;
assign n_2548 =  n_2546 &  n_2547;
assign n_2549 =  n_2545 &  n_2548;
assign n_2550 =  n_2542 &  n_2549;
assign n_2551 =  n_2535 &  n_2550;
assign n_2552 =  n_2524 &  n_2551;
assign n_2553 = ~n_1957 & ~n_1978;
assign n_2554 = ~n_1979 & ~n_2553;
assign n_2555 = ~n_2485 & ~n_2491;
assign n_2556 =  n_2483 & ~n_2555;
assign n_2557 = ~n_2554 &  n_2556;
assign n_2558 = ~n_2483 & ~n_2488;
assign n_2559 = ~n_2556 & ~n_2558;
assign n_2560 =  n_2483 &  n_2487;
assign n_2561 = ~n_2492 & ~n_2560;
assign n_2562 =  n_2559 &  n_2561;
assign n_2563 = ~n_2554 & ~n_2561;
assign n_2564 = ~n_2562 & ~n_2563;
assign n_2565 = ~n_2557 &  n_2564;
assign n_2566 = ~n_2552 & ~n_2565;
assign n_2567 = ~n_1869 & ~n_2374;
assign n_2568 = ~n_2375 & ~n_2567;
assign n_2569 = ~n_2556 & ~n_2562;
assign n_2570 =  n_2554 & ~n_2569;
assign n_2571 = ~n_2568 &  n_2570;
assign n_2572 = ~n_2554 & ~n_2559;
assign n_2573 = ~n_2570 & ~n_2572;
assign n_2574 =  n_2554 &  n_2558;
assign n_2575 = ~n_2563 & ~n_2574;
assign n_2576 =  n_2573 &  n_2575;
assign n_2577 = ~n_2568 & ~n_2575;
assign n_2578 = ~n_2576 & ~n_2577;
assign n_2579 = ~n_2571 &  n_2578;
assign n_2580 = ~n_1953 & ~n_1996;
assign n_2581 = ~n_1997 & ~n_2580;
assign n_2582 = ~n_2570 & ~n_2576;
assign n_2583 =  n_2568 & ~n_2582;
assign n_2584 = ~n_2581 &  n_2583;
assign n_2585 = ~n_2568 & ~n_2573;
assign n_2586 = ~n_2583 & ~n_2585;
assign n_2587 =  n_2568 &  n_2572;
assign n_2588 = ~n_2577 & ~n_2587;
assign n_2589 =  n_2586 &  n_2588;
assign n_2590 = ~n_2581 & ~n_2588;
assign n_2591 = ~n_2589 & ~n_2590;
assign n_2592 = ~n_2584 &  n_2591;
assign n_2593 = ~n_1873 & ~n_2356;
assign n_2594 = ~n_2357 & ~n_2593;
assign n_2595 = ~n_2583 & ~n_2589;
assign n_2596 =  n_2581 & ~n_2595;
assign n_2597 = ~n_2594 &  n_2596;
assign n_2598 = ~n_2581 & ~n_2586;
assign n_2599 = ~n_2596 & ~n_2598;
assign n_2600 =  n_2581 &  n_2585;
assign n_2601 = ~n_2590 & ~n_2600;
assign n_2602 =  n_2599 &  n_2601;
assign n_2603 = ~n_2594 & ~n_2601;
assign n_2604 = ~n_2602 & ~n_2603;
assign n_2605 = ~n_2597 &  n_2604;
assign n_2606 = ~n_1949 & ~n_2014;
assign n_2607 = ~n_2015 & ~n_2606;
assign n_2608 = ~n_2596 & ~n_2602;
assign n_2609 =  n_2594 & ~n_2608;
assign n_2610 = ~n_2607 &  n_2609;
assign n_2611 = ~n_2594 & ~n_2599;
assign n_2612 = ~n_2609 & ~n_2611;
assign n_2613 =  n_2594 &  n_2598;
assign n_2614 = ~n_2603 & ~n_2613;
assign n_2615 =  n_2612 &  n_2614;
assign n_2616 = ~n_2607 & ~n_2614;
assign n_2617 = ~n_2615 & ~n_2616;
assign n_2618 = ~n_2610 &  n_2617;
assign n_2619 = ~n_1877 & ~n_2338;
assign n_2620 = ~n_2339 & ~n_2619;
assign n_2621 = ~n_2609 & ~n_2615;
assign n_2622 =  n_2607 & ~n_2621;
assign n_2623 = ~n_2620 &  n_2622;
assign n_2624 = ~n_2607 & ~n_2612;
assign n_2625 = ~n_2622 & ~n_2624;
assign n_2626 =  n_2607 &  n_2611;
assign n_2627 = ~n_2616 & ~n_2626;
assign n_2628 =  n_2625 &  n_2627;
assign n_2629 = ~n_2620 & ~n_2627;
assign n_2630 = ~n_2628 & ~n_2629;
assign n_2631 = ~n_2623 &  n_2630;
assign n_2632 = ~n_1945 & ~n_2032;
assign n_2633 = ~n_2033 & ~n_2632;
assign n_2634 = ~n_2622 & ~n_2628;
assign n_2635 =  n_2620 & ~n_2634;
assign n_2636 = ~n_2633 &  n_2635;
assign n_2637 = ~n_2620 & ~n_2625;
assign n_2638 = ~n_2635 & ~n_2637;
assign n_2639 =  n_2620 &  n_2624;
assign n_2640 = ~n_2629 & ~n_2639;
assign n_2641 =  n_2638 &  n_2640;
assign n_2642 = ~n_2633 & ~n_2640;
assign n_2643 = ~n_2641 & ~n_2642;
assign n_2644 = ~n_2636 &  n_2643;
assign n_2645 = ~n_1881 & ~n_2320;
assign n_2646 = ~n_2321 & ~n_2645;
assign n_2647 = ~n_2635 & ~n_2641;
assign n_2648 =  n_2633 & ~n_2647;
assign n_2649 = ~n_2646 &  n_2648;
assign n_2650 = ~n_2633 & ~n_2638;
assign n_2651 = ~n_2648 & ~n_2650;
assign n_2652 =  n_2633 &  n_2637;
assign n_2653 = ~n_2642 & ~n_2652;
assign n_2654 =  n_2651 &  n_2653;
assign n_2655 = ~n_2646 & ~n_2653;
assign n_2656 = ~n_2654 & ~n_2655;
assign n_2657 = ~n_2649 &  n_2656;
assign n_2658 = ~n_1941 & ~n_2050;
assign n_2659 = ~n_2051 & ~n_2658;
assign n_2660 = ~n_2648 & ~n_2654;
assign n_2661 =  n_2646 & ~n_2660;
assign n_2662 = ~n_2659 &  n_2661;
assign n_2663 = ~n_2646 & ~n_2651;
assign n_2664 = ~n_2661 & ~n_2663;
assign n_2665 =  n_2646 &  n_2650;
assign n_2666 = ~n_2655 & ~n_2665;
assign n_2667 =  n_2664 &  n_2666;
assign n_2668 = ~n_2659 & ~n_2666;
assign n_2669 = ~n_2667 & ~n_2668;
assign n_2670 = ~n_2662 &  n_2669;
assign n_2671 = ~n_1885 & ~n_2302;
assign n_2672 = ~n_2303 & ~n_2671;
assign n_2673 = ~n_2661 & ~n_2667;
assign n_2674 =  n_2659 & ~n_2673;
assign n_2675 = ~n_2672 &  n_2674;
assign n_2676 = ~n_2659 & ~n_2664;
assign n_2677 = ~n_2674 & ~n_2676;
assign n_2678 =  n_2659 &  n_2663;
assign n_2679 = ~n_2668 & ~n_2678;
assign n_2680 =  n_2677 &  n_2679;
assign n_2681 = ~n_2672 & ~n_2679;
assign n_2682 = ~n_2680 & ~n_2681;
assign n_2683 = ~n_2675 &  n_2682;
assign n_2684 = ~n_1937 & ~n_2068;
assign n_2685 = ~n_2069 & ~n_2684;
assign n_2686 = ~n_2674 & ~n_2680;
assign n_2687 =  n_2672 & ~n_2686;
assign n_2688 = ~n_2685 &  n_2687;
assign n_2689 = ~n_2672 & ~n_2677;
assign n_2690 = ~n_2687 & ~n_2689;
assign n_2691 =  n_2672 &  n_2676;
assign n_2692 = ~n_2681 & ~n_2691;
assign n_2693 =  n_2690 &  n_2692;
assign n_2694 = ~n_2685 & ~n_2692;
assign n_2695 = ~n_2693 & ~n_2694;
assign n_2696 = ~n_2688 &  n_2695;
assign n_2697 = ~n_1889 & ~n_2284;
assign n_2698 = ~n_2285 & ~n_2697;
assign n_2699 = ~n_2687 & ~n_2693;
assign n_2700 =  n_2685 & ~n_2699;
assign n_2701 = ~n_2698 &  n_2700;
assign n_2702 = ~n_2685 & ~n_2690;
assign n_2703 = ~n_2700 & ~n_2702;
assign n_2704 =  n_2685 &  n_2689;
assign n_2705 = ~n_2694 & ~n_2704;
assign n_2706 =  n_2703 &  n_2705;
assign n_2707 = ~n_2698 & ~n_2705;
assign n_2708 = ~n_2706 & ~n_2707;
assign n_2709 = ~n_2701 &  n_2708;
assign n_2710 = ~n_1933 & ~n_2086;
assign n_2711 = ~n_2087 & ~n_2710;
assign n_2712 = ~n_2700 & ~n_2706;
assign n_2713 =  n_2698 & ~n_2712;
assign n_2714 = ~n_2711 &  n_2713;
assign n_2715 = ~n_2698 & ~n_2703;
assign n_2716 = ~n_2713 & ~n_2715;
assign n_2717 =  n_2698 &  n_2702;
assign n_2718 = ~n_2707 & ~n_2717;
assign n_2719 =  n_2716 &  n_2718;
assign n_2720 = ~n_2711 & ~n_2718;
assign n_2721 = ~n_2719 & ~n_2720;
assign n_2722 = ~n_2714 &  n_2721;
assign n_2723 = ~n_1893 & ~n_2266;
assign n_2724 = ~n_2267 & ~n_2723;
assign n_2725 = ~n_2713 & ~n_2719;
assign n_2726 =  n_2711 & ~n_2725;
assign n_2727 = ~n_2724 &  n_2726;
assign n_2728 = ~n_2711 & ~n_2716;
assign n_2729 = ~n_2726 & ~n_2728;
assign n_2730 =  n_2711 &  n_2715;
assign n_2731 = ~n_2720 & ~n_2730;
assign n_2732 =  n_2729 &  n_2731;
assign n_2733 = ~n_2724 & ~n_2731;
assign n_2734 = ~n_2732 & ~n_2733;
assign n_2735 = ~n_2727 &  n_2734;
assign n_2736 = ~n_1929 & ~n_2104;
assign n_2737 = ~n_2105 & ~n_2736;
assign n_2738 = ~n_2726 & ~n_2732;
assign n_2739 =  n_2724 & ~n_2738;
assign n_2740 = ~n_2737 &  n_2739;
assign n_2741 = ~n_2724 & ~n_2729;
assign n_2742 = ~n_2739 & ~n_2741;
assign n_2743 =  n_2724 &  n_2728;
assign n_2744 = ~n_2733 & ~n_2743;
assign n_2745 =  n_2742 &  n_2744;
assign n_2746 = ~n_2737 & ~n_2744;
assign n_2747 = ~n_2745 & ~n_2746;
assign n_2748 = ~n_2740 &  n_2747;
assign n_2749 = ~n_1897 & ~n_2248;
assign n_2750 = ~n_2249 & ~n_2749;
assign n_2751 = ~n_2739 & ~n_2745;
assign n_2752 =  n_2737 & ~n_2751;
assign n_2753 = ~n_2750 &  n_2752;
assign n_2754 = ~n_2737 & ~n_2742;
assign n_2755 = ~n_2752 & ~n_2754;
assign n_2756 =  n_2737 &  n_2741;
assign n_2757 = ~n_2746 & ~n_2756;
assign n_2758 =  n_2755 &  n_2757;
assign n_2759 = ~n_2750 & ~n_2757;
assign n_2760 = ~n_2758 & ~n_2759;
assign n_2761 = ~n_2753 &  n_2760;
assign n_2762 = ~n_1925 & ~n_2122;
assign n_2763 = ~n_2123 & ~n_2762;
assign n_2764 = ~n_2752 & ~n_2758;
assign n_2765 =  n_2750 & ~n_2764;
assign n_2766 = ~n_2763 &  n_2765;
assign n_2767 = ~n_2750 & ~n_2755;
assign n_2768 = ~n_2765 & ~n_2767;
assign n_2769 =  n_2750 &  n_2754;
assign n_2770 = ~n_2759 & ~n_2769;
assign n_2771 =  n_2768 &  n_2770;
assign n_2772 = ~n_2763 & ~n_2770;
assign n_2773 = ~n_2771 & ~n_2772;
assign n_2774 = ~n_2766 &  n_2773;
assign n_2775 = ~n_1901 & ~n_2230;
assign n_2776 = ~n_2231 & ~n_2775;
assign n_2777 = ~n_2765 & ~n_2771;
assign n_2778 =  n_2763 & ~n_2777;
assign n_2779 = ~n_2776 &  n_2778;
assign n_2780 = ~n_2763 & ~n_2768;
assign n_2781 = ~n_2778 & ~n_2780;
assign n_2782 =  n_2763 &  n_2767;
assign n_2783 = ~n_2772 & ~n_2782;
assign n_2784 =  n_2781 &  n_2783;
assign n_2785 = ~n_2776 & ~n_2783;
assign n_2786 = ~n_2784 & ~n_2785;
assign n_2787 = ~n_2779 &  n_2786;
assign n_2788 = ~n_1921 & ~n_2140;
assign n_2789 = ~n_2141 & ~n_2788;
assign n_2790 = ~n_2778 & ~n_2784;
assign n_2791 =  n_2776 & ~n_2790;
assign n_2792 = ~n_2789 &  n_2791;
assign n_2793 = ~n_2776 & ~n_2781;
assign n_2794 = ~n_2791 & ~n_2793;
assign n_2795 =  n_2776 &  n_2780;
assign n_2796 = ~n_2785 & ~n_2795;
assign n_2797 =  n_2794 &  n_2796;
assign n_2798 = ~n_2789 & ~n_2796;
assign n_2799 = ~n_2797 & ~n_2798;
assign n_2800 = ~n_2792 &  n_2799;
assign n_2801 = ~n_1905 & ~n_2212;
assign n_2802 = ~n_2213 & ~n_2801;
assign n_2803 = ~n_2791 & ~n_2797;
assign n_2804 =  n_2789 & ~n_2803;
assign n_2805 = ~n_2802 &  n_2804;
assign n_2806 = ~n_2789 & ~n_2794;
assign n_2807 = ~n_2804 & ~n_2806;
assign n_2808 =  n_2789 &  n_2793;
assign n_2809 = ~n_2798 & ~n_2808;
assign n_2810 =  n_2807 &  n_2809;
assign n_2811 = ~n_2802 & ~n_2809;
assign n_2812 = ~n_2810 & ~n_2811;
assign n_2813 = ~n_2805 &  n_2812;
assign n_2814 = ~n_1917 & ~n_2158;
assign n_2815 = ~n_2159 & ~n_2814;
assign n_2816 = ~n_2804 & ~n_2810;
assign n_2817 =  n_2802 & ~n_2816;
assign n_2818 = ~n_2815 &  n_2817;
assign n_2819 = ~n_2802 & ~n_2807;
assign n_2820 = ~n_2817 & ~n_2819;
assign n_2821 =  n_2802 &  n_2806;
assign n_2822 = ~n_2811 & ~n_2821;
assign n_2823 =  n_2820 &  n_2822;
assign n_2824 = ~n_2815 & ~n_2822;
assign n_2825 = ~n_2823 & ~n_2824;
assign n_2826 = ~n_2818 &  n_2825;
assign n_2827 = ~n_1909 & ~n_2194;
assign n_2828 = ~n_2195 & ~n_2827;
assign n_2829 = ~n_2817 & ~n_2823;
assign n_2830 =  n_2815 & ~n_2829;
assign n_2831 = ~n_2828 &  n_2830;
assign n_2832 = ~n_2815 & ~n_2820;
assign n_2833 = ~n_2830 & ~n_2832;
assign n_2834 =  n_2815 &  n_2819;
assign n_2835 = ~n_2824 & ~n_2834;
assign n_2836 =  n_2833 &  n_2835;
assign n_2837 = ~n_2828 & ~n_2835;
assign n_2838 = ~n_2836 & ~n_2837;
assign n_2839 = ~n_2831 &  n_2838;
assign n_2840 = ~n_1913 & ~n_2176;
assign n_2841 = ~n_2177 & ~n_2840;
assign n_2842 = ~n_2830 & ~n_2836;
assign n_2843 =  n_2828 & ~n_2842;
assign n_2844 = ~n_2841 &  n_2843;
assign n_2845 = ~n_2828 & ~n_2833;
assign n_2846 = ~n_2843 & ~n_2845;
assign n_2847 =  n_2828 &  n_2832;
assign n_2848 = ~n_2837 & ~n_2847;
assign n_2849 =  n_2846 &  n_2848;
assign n_2850 = ~n_2841 & ~n_2848;
assign n_2851 = ~n_2849 & ~n_2850;
assign n_2852 = ~n_2844 &  n_2851;
assign n_2853 = ~n_1911 & ~n_2185;
assign n_2854 = ~n_2186 & ~n_2853;
assign n_2855 = ~n_2843 & ~n_2849;
assign n_2856 =  n_2841 & ~n_2855;
assign n_2857 = ~n_2854 &  n_2856;
assign n_2858 = ~n_2841 & ~n_2846;
assign n_2859 = ~n_2856 & ~n_2858;
assign n_2860 =  n_2841 &  n_2845;
assign n_2861 = ~n_2850 & ~n_2860;
assign n_2862 =  n_2859 &  n_2861;
assign n_2863 = ~n_2854 & ~n_2861;
assign n_2864 = ~n_2862 & ~n_2863;
assign n_2865 = ~n_2857 &  n_2864;
assign n_2866 = ~n_1915 & ~n_2167;
assign n_2867 = ~n_2168 & ~n_2866;
assign n_2868 = ~n_2856 & ~n_2862;
assign n_2869 =  n_2854 & ~n_2868;
assign n_2870 = ~n_2867 &  n_2869;
assign n_2871 = ~n_2854 & ~n_2859;
assign n_2872 = ~n_2869 & ~n_2871;
assign n_2873 =  n_2854 &  n_2858;
assign n_2874 = ~n_2863 & ~n_2873;
assign n_2875 =  n_2872 &  n_2874;
assign n_2876 = ~n_2867 & ~n_2874;
assign n_2877 = ~n_2875 & ~n_2876;
assign n_2878 = ~n_2870 &  n_2877;
assign n_2879 = ~n_1907 & ~n_2203;
assign n_2880 = ~n_2204 & ~n_2879;
assign n_2881 = ~n_2869 & ~n_2875;
assign n_2882 =  n_2867 & ~n_2881;
assign n_2883 = ~n_2880 &  n_2882;
assign n_2884 = ~n_2867 & ~n_2872;
assign n_2885 = ~n_2882 & ~n_2884;
assign n_2886 =  n_2867 &  n_2871;
assign n_2887 = ~n_2876 & ~n_2886;
assign n_2888 =  n_2885 &  n_2887;
assign n_2889 = ~n_2880 & ~n_2887;
assign n_2890 = ~n_2888 & ~n_2889;
assign n_2891 = ~n_2883 &  n_2890;
assign n_2892 = ~n_1919 & ~n_2149;
assign n_2893 = ~n_2150 & ~n_2892;
assign n_2894 = ~n_2882 & ~n_2888;
assign n_2895 =  n_2880 & ~n_2894;
assign n_2896 = ~n_2893 &  n_2895;
assign n_2897 = ~n_2880 & ~n_2885;
assign n_2898 = ~n_2895 & ~n_2897;
assign n_2899 =  n_2880 &  n_2884;
assign n_2900 = ~n_2889 & ~n_2899;
assign n_2901 =  n_2898 &  n_2900;
assign n_2902 = ~n_2893 & ~n_2900;
assign n_2903 = ~n_2901 & ~n_2902;
assign n_2904 = ~n_2896 &  n_2903;
assign n_2905 = ~n_1903 & ~n_2221;
assign n_2906 = ~n_2222 & ~n_2905;
assign n_2907 = ~n_2895 & ~n_2901;
assign n_2908 =  n_2893 & ~n_2907;
assign n_2909 = ~n_2906 &  n_2908;
assign n_2910 = ~n_2893 & ~n_2898;
assign n_2911 = ~n_2908 & ~n_2910;
assign n_2912 =  n_2893 &  n_2897;
assign n_2913 = ~n_2902 & ~n_2912;
assign n_2914 =  n_2911 &  n_2913;
assign n_2915 = ~n_2906 & ~n_2913;
assign n_2916 = ~n_2914 & ~n_2915;
assign n_2917 = ~n_2909 &  n_2916;
assign n_2918 = ~n_1923 & ~n_2131;
assign n_2919 = ~n_2132 & ~n_2918;
assign n_2920 = ~n_2908 & ~n_2914;
assign n_2921 =  n_2906 & ~n_2920;
assign n_2922 = ~n_2919 &  n_2921;
assign n_2923 = ~n_2906 & ~n_2911;
assign n_2924 = ~n_2921 & ~n_2923;
assign n_2925 =  n_2906 &  n_2910;
assign n_2926 = ~n_2915 & ~n_2925;
assign n_2927 =  n_2924 &  n_2926;
assign n_2928 = ~n_2919 & ~n_2926;
assign n_2929 = ~n_2927 & ~n_2928;
assign n_2930 = ~n_2922 &  n_2929;
assign n_2931 = ~n_1899 & ~n_2239;
assign n_2932 = ~n_2240 & ~n_2931;
assign n_2933 = ~n_2921 & ~n_2927;
assign n_2934 =  n_2919 & ~n_2933;
assign n_2935 = ~n_2932 &  n_2934;
assign n_2936 = ~n_2919 & ~n_2924;
assign n_2937 = ~n_2934 & ~n_2936;
assign n_2938 =  n_2919 &  n_2923;
assign n_2939 = ~n_2928 & ~n_2938;
assign n_2940 =  n_2937 &  n_2939;
assign n_2941 = ~n_2932 & ~n_2939;
assign n_2942 = ~n_2940 & ~n_2941;
assign n_2943 = ~n_2935 &  n_2942;
assign n_2944 = ~n_1927 & ~n_2113;
assign n_2945 = ~n_2114 & ~n_2944;
assign n_2946 = ~n_2934 & ~n_2940;
assign n_2947 =  n_2932 & ~n_2946;
assign n_2948 = ~n_2945 &  n_2947;
assign n_2949 = ~n_2932 & ~n_2937;
assign n_2950 = ~n_2947 & ~n_2949;
assign n_2951 =  n_2932 &  n_2936;
assign n_2952 = ~n_2941 & ~n_2951;
assign n_2953 =  n_2950 &  n_2952;
assign n_2954 = ~n_2945 & ~n_2952;
assign n_2955 = ~n_2953 & ~n_2954;
assign n_2956 = ~n_2948 &  n_2955;
assign n_2957 = ~n_1895 & ~n_2257;
assign n_2958 = ~n_2258 & ~n_2957;
assign n_2959 = ~n_2947 & ~n_2953;
assign n_2960 =  n_2945 & ~n_2959;
assign n_2961 = ~n_2958 &  n_2960;
assign n_2962 = ~n_2945 & ~n_2950;
assign n_2963 = ~n_2960 & ~n_2962;
assign n_2964 =  n_2945 &  n_2949;
assign n_2965 = ~n_2954 & ~n_2964;
assign n_2966 =  n_2963 &  n_2965;
assign n_2967 = ~n_2958 & ~n_2965;
assign n_2968 = ~n_2966 & ~n_2967;
assign n_2969 = ~n_2961 &  n_2968;
assign n_2970 = ~n_1931 & ~n_2095;
assign n_2971 = ~n_2096 & ~n_2970;
assign n_2972 = ~n_2960 & ~n_2966;
assign n_2973 =  n_2958 & ~n_2972;
assign n_2974 = ~n_2971 &  n_2973;
assign n_2975 = ~n_2958 & ~n_2963;
assign n_2976 = ~n_2973 & ~n_2975;
assign n_2977 =  n_2958 &  n_2962;
assign n_2978 = ~n_2967 & ~n_2977;
assign n_2979 =  n_2976 &  n_2978;
assign n_2980 = ~n_2971 & ~n_2978;
assign n_2981 = ~n_2979 & ~n_2980;
assign n_2982 = ~n_2974 &  n_2981;
assign n_2983 = ~n_1891 & ~n_2275;
assign n_2984 = ~n_2276 & ~n_2983;
assign n_2985 = ~n_2973 & ~n_2979;
assign n_2986 =  n_2971 & ~n_2985;
assign n_2987 = ~n_2984 &  n_2986;
assign n_2988 = ~n_2971 & ~n_2976;
assign n_2989 = ~n_2986 & ~n_2988;
assign n_2990 =  n_2971 &  n_2975;
assign n_2991 = ~n_2980 & ~n_2990;
assign n_2992 =  n_2989 &  n_2991;
assign n_2993 = ~n_2984 & ~n_2991;
assign n_2994 = ~n_2992 & ~n_2993;
assign n_2995 = ~n_2987 &  n_2994;
assign n_2996 = ~n_1935 & ~n_2077;
assign n_2997 = ~n_2078 & ~n_2996;
assign n_2998 = ~n_2986 & ~n_2992;
assign n_2999 =  n_2984 & ~n_2998;
assign n_3000 = ~n_2997 &  n_2999;
assign n_3001 = ~n_2984 & ~n_2989;
assign n_3002 = ~n_2999 & ~n_3001;
assign n_3003 =  n_2984 &  n_2988;
assign n_3004 = ~n_2993 & ~n_3003;
assign n_3005 =  n_3002 &  n_3004;
assign n_3006 = ~n_2997 & ~n_3004;
assign n_3007 = ~n_3005 & ~n_3006;
assign n_3008 = ~n_3000 &  n_3007;
assign n_3009 = ~n_1887 & ~n_2293;
assign n_3010 = ~n_2294 & ~n_3009;
assign n_3011 = ~n_2999 & ~n_3005;
assign n_3012 =  n_2997 & ~n_3011;
assign n_3013 = ~n_3010 &  n_3012;
assign n_3014 = ~n_2997 & ~n_3002;
assign n_3015 = ~n_3012 & ~n_3014;
assign n_3016 =  n_2997 &  n_3001;
assign n_3017 = ~n_3006 & ~n_3016;
assign n_3018 =  n_3015 &  n_3017;
assign n_3019 = ~n_3010 & ~n_3017;
assign n_3020 = ~n_3018 & ~n_3019;
assign n_3021 = ~n_3013 &  n_3020;
assign n_3022 = ~n_1939 & ~n_2059;
assign n_3023 = ~n_2060 & ~n_3022;
assign n_3024 = ~n_3012 & ~n_3018;
assign n_3025 =  n_3010 & ~n_3024;
assign n_3026 = ~n_3023 &  n_3025;
assign n_3027 = ~n_3010 & ~n_3015;
assign n_3028 = ~n_3025 & ~n_3027;
assign n_3029 =  n_3010 &  n_3014;
assign n_3030 = ~n_3019 & ~n_3029;
assign n_3031 =  n_3028 &  n_3030;
assign n_3032 = ~n_3023 & ~n_3030;
assign n_3033 = ~n_3031 & ~n_3032;
assign n_3034 = ~n_3026 &  n_3033;
assign n_3035 = ~n_1883 & ~n_2311;
assign n_3036 = ~n_2312 & ~n_3035;
assign n_3037 = ~n_3025 & ~n_3031;
assign n_3038 =  n_3023 & ~n_3037;
assign n_3039 = ~n_3036 &  n_3038;
assign n_3040 = ~n_3023 & ~n_3028;
assign n_3041 = ~n_3038 & ~n_3040;
assign n_3042 =  n_3023 &  n_3027;
assign n_3043 = ~n_3032 & ~n_3042;
assign n_3044 =  n_3041 &  n_3043;
assign n_3045 = ~n_3036 & ~n_3043;
assign n_3046 = ~n_3044 & ~n_3045;
assign n_3047 = ~n_3039 &  n_3046;
assign n_3048 = ~n_1943 & ~n_2041;
assign n_3049 = ~n_2042 & ~n_3048;
assign n_3050 = ~n_3038 & ~n_3044;
assign n_3051 =  n_3036 & ~n_3050;
assign n_3052 = ~n_3049 &  n_3051;
assign n_3053 = ~n_3036 & ~n_3041;
assign n_3054 = ~n_3051 & ~n_3053;
assign n_3055 =  n_3036 &  n_3040;
assign n_3056 = ~n_3045 & ~n_3055;
assign n_3057 =  n_3054 &  n_3056;
assign n_3058 = ~n_3049 & ~n_3056;
assign n_3059 = ~n_3057 & ~n_3058;
assign n_3060 = ~n_3052 &  n_3059;
assign n_3061 = ~n_1879 & ~n_2329;
assign n_3062 = ~n_2330 & ~n_3061;
assign n_3063 = ~n_3051 & ~n_3057;
assign n_3064 =  n_3049 & ~n_3063;
assign n_3065 = ~n_3062 &  n_3064;
assign n_3066 = ~n_3049 & ~n_3054;
assign n_3067 = ~n_3064 & ~n_3066;
assign n_3068 =  n_3049 &  n_3053;
assign n_3069 = ~n_3058 & ~n_3068;
assign n_3070 =  n_3067 &  n_3069;
assign n_3071 = ~n_3062 & ~n_3069;
assign n_3072 = ~n_3070 & ~n_3071;
assign n_3073 = ~n_3065 &  n_3072;
assign n_3074 = ~n_1947 & ~n_2023;
assign n_3075 = ~n_2024 & ~n_3074;
assign n_3076 = ~n_3064 & ~n_3070;
assign n_3077 =  n_3062 & ~n_3076;
assign n_3078 = ~n_3075 &  n_3077;
assign n_3079 = ~n_3062 & ~n_3067;
assign n_3080 = ~n_3077 & ~n_3079;
assign n_3081 =  n_3062 &  n_3066;
assign n_3082 = ~n_3071 & ~n_3081;
assign n_3083 =  n_3080 &  n_3082;
assign n_3084 = ~n_3075 & ~n_3082;
assign n_3085 = ~n_3083 & ~n_3084;
assign n_3086 = ~n_3078 &  n_3085;
assign n_3087 = ~n_1875 & ~n_2347;
assign n_3088 = ~n_2348 & ~n_3087;
assign n_3089 = ~n_3077 & ~n_3083;
assign n_3090 =  n_3075 & ~n_3089;
assign n_3091 = ~n_3088 &  n_3090;
assign n_3092 = ~n_3075 & ~n_3080;
assign n_3093 = ~n_3090 & ~n_3092;
assign n_3094 =  n_3075 &  n_3079;
assign n_3095 = ~n_3084 & ~n_3094;
assign n_3096 =  n_3093 &  n_3095;
assign n_3097 = ~n_3088 & ~n_3095;
assign n_3098 = ~n_3096 & ~n_3097;
assign n_3099 = ~n_3091 &  n_3098;
assign n_3100 = ~n_1951 & ~n_2005;
assign n_3101 = ~n_2006 & ~n_3100;
assign n_3102 = ~n_3090 & ~n_3096;
assign n_3103 =  n_3088 & ~n_3102;
assign n_3104 = ~n_3101 &  n_3103;
assign n_3105 = ~n_3088 & ~n_3093;
assign n_3106 = ~n_3103 & ~n_3105;
assign n_3107 =  n_3088 &  n_3092;
assign n_3108 = ~n_3097 & ~n_3107;
assign n_3109 =  n_3106 &  n_3108;
assign n_3110 = ~n_3101 & ~n_3108;
assign n_3111 = ~n_3109 & ~n_3110;
assign n_3112 = ~n_3104 &  n_3111;
assign n_3113 = ~n_1871 & ~n_2365;
assign n_3114 = ~n_2366 & ~n_3113;
assign n_3115 = ~n_3103 & ~n_3109;
assign n_3116 =  n_3101 & ~n_3115;
assign n_3117 = ~n_3114 &  n_3116;
assign n_3118 = ~n_3101 & ~n_3106;
assign n_3119 = ~n_3116 & ~n_3118;
assign n_3120 =  n_3101 &  n_3105;
assign n_3121 = ~n_3110 & ~n_3120;
assign n_3122 =  n_3119 &  n_3121;
assign n_3123 = ~n_3114 & ~n_3121;
assign n_3124 = ~n_3122 & ~n_3123;
assign n_3125 = ~n_3117 &  n_3124;
assign n_3126 = ~n_1955 & ~n_1987;
assign n_3127 = ~n_1988 & ~n_3126;
assign n_3128 = ~n_3116 & ~n_3122;
assign n_3129 =  n_3114 & ~n_3128;
assign n_3130 = ~n_3127 &  n_3129;
assign n_3131 = ~n_3114 & ~n_3119;
assign n_3132 = ~n_3129 & ~n_3131;
assign n_3133 =  n_3114 &  n_3118;
assign n_3134 = ~n_3123 & ~n_3133;
assign n_3135 =  n_3132 &  n_3134;
assign n_3136 = ~n_3127 & ~n_3134;
assign n_3137 = ~n_3135 & ~n_3136;
assign n_3138 = ~n_3130 &  n_3137;
assign n_3139 = ~n_1867 & ~n_2383;
assign n_3140 = ~n_2384 & ~n_3139;
assign n_3141 = ~n_3129 & ~n_3135;
assign n_3142 =  n_3127 & ~n_3141;
assign n_3143 = ~n_3140 &  n_3142;
assign n_3144 = ~n_3127 & ~n_3132;
assign n_3145 = ~n_3142 & ~n_3144;
assign n_3146 =  n_3127 &  n_3131;
assign n_3147 = ~n_3136 & ~n_3146;
assign n_3148 =  n_3145 &  n_3147;
assign n_3149 = ~n_3140 & ~n_3147;
assign n_3150 = ~n_3148 & ~n_3149;
assign n_3151 = ~n_3143 &  n_3150;
assign n_3152 = ~n_2552 & ~n_3151;
assign n_3153 = ~n_1959 & ~n_1969;
assign n_3154 = ~n_1970 & ~n_3153;
assign n_3155 = ~n_3142 & ~n_3148;
assign n_3156 =  n_3140 & ~n_3155;
assign n_3157 = ~n_3154 &  n_3156;
assign n_3158 = ~n_3140 & ~n_3145;
assign n_3159 = ~n_3156 & ~n_3158;
assign n_3160 =  n_3140 &  n_3144;
assign n_3161 = ~n_3149 & ~n_3160;
assign n_3162 =  n_3159 &  n_3161;
assign n_3163 = ~n_3154 & ~n_3161;
assign n_3164 = ~n_3162 & ~n_3163;
assign n_3165 = ~n_3157 &  n_3164;
assign n_3166 = ~n_1863 & ~n_2401;
assign n_3167 = ~n_2402 & ~n_3166;
assign n_3168 = ~n_3156 & ~n_3162;
assign n_3169 =  n_3154 & ~n_3168;
assign n_3170 = ~n_3167 &  n_3169;
assign n_3171 = ~n_3154 & ~n_3159;
assign n_3172 = ~n_3169 & ~n_3171;
assign n_3173 =  n_3154 &  n_3158;
assign n_3174 = ~n_3163 & ~n_3173;
assign n_3175 =  n_3172 &  n_3174;
assign n_3176 = ~n_3167 & ~n_3174;
assign n_3177 = ~n_3175 & ~n_3176;
assign n_3178 = ~n_3170 &  n_3177;
assign n_3179 = ~n_1753 & ~n_1849;
assign n_3180 = ~n_1850 & ~n_3179;
assign n_3181 = ~n_3169 & ~n_3175;
assign n_3182 =  n_3167 & ~n_3181;
assign n_3183 = ~n_3180 &  n_3182;
assign n_3184 = ~n_3167 & ~n_3172;
assign n_3185 = ~n_3182 & ~n_3184;
assign n_3186 =  n_3167 &  n_3171;
assign n_3187 = ~n_3176 & ~n_3186;
assign n_3188 =  n_3185 &  n_3187;
assign n_3189 = ~n_3180 & ~n_3187;
assign n_3190 = ~n_3188 & ~n_3189;
assign n_3191 = ~n_3183 &  n_3190;
assign n_3192 = ~n_2552 & ~n_3191;
assign n_3193 = ~n_2420 & ~n_2428;
assign n_3194 = ~n_2429 & ~n_3193;
assign n_3195 = ~n_3182 & ~n_3188;
assign n_3196 =  n_3180 & ~n_3195;
assign n_3197 = ~n_3194 &  n_3196;
assign n_3198 = ~n_3180 & ~n_3185;
assign n_3199 = ~n_3196 & ~n_3198;
assign n_3200 =  n_3180 &  n_3184;
assign n_3201 = ~n_3189 & ~n_3200;
assign n_3202 =  n_3199 &  n_3201;
assign n_3203 = ~n_3194 & ~n_3201;
assign n_3204 = ~n_3202 & ~n_3203;
assign n_3205 = ~n_3197 &  n_3204;
assign n_3206 = ~n_1779 & ~n_1831;
assign n_3207 = ~n_1832 & ~n_3206;
assign n_3208 = ~n_3196 & ~n_3202;
assign n_3209 =  n_3194 & ~n_3208;
assign n_3210 = ~n_3207 &  n_3209;
assign n_3211 = ~n_3194 & ~n_3199;
assign n_3212 = ~n_3209 & ~n_3211;
assign n_3213 =  n_3194 &  n_3198;
assign n_3214 = ~n_3203 & ~n_3213;
assign n_3215 =  n_3212 &  n_3214;
assign n_3216 = ~n_3207 & ~n_3214;
assign n_3217 = ~n_3215 & ~n_3216;
assign n_3218 = ~n_3210 &  n_3217;
assign n_3219 = ~n_2552 & ~n_3218;
assign n_3220 = ~n_2416 & ~n_2435;
assign n_3221 = ~n_2444 & ~n_3220;
assign n_3222 = ~n_3209 & ~n_3215;
assign n_3223 =  n_3207 & ~n_3222;
assign n_3224 = ~n_3221 &  n_3223;
assign n_3225 = ~n_3207 & ~n_3212;
assign n_3226 = ~n_3223 & ~n_3225;
assign n_3227 =  n_3207 &  n_3211;
assign n_3228 = ~n_3216 & ~n_3227;
assign n_3229 =  n_3226 &  n_3228;
assign n_3230 = ~n_3221 & ~n_3228;
assign n_3231 = ~n_3229 & ~n_3230;
assign n_3232 = ~n_3224 &  n_3231;
assign n_3233 = ~n_1812 & ~n_1819;
assign n_3234 = ~n_3221 & ~n_3226;
assign n_3235 = ~n_3223 & ~n_3229;
assign n_3236 =  n_3221 & ~n_3235;
assign n_3237 = ~n_3234 & ~n_3236;
assign n_3238 =  n_3221 &  n_3225;
assign n_3239 = ~n_3230 & ~n_3238;
assign n_3240 =  n_3237 &  n_3239;
assign n_3241 =  n_3233 &  n_3240;
assign n_3242 = ~n_3232 &  n_3241;
assign n_3243 =  n_3219 &  n_3242;
assign n_3244 = ~n_3205 &  n_3243;
assign n_3245 =  n_3192 &  n_3244;
assign n_3246 = ~n_3178 &  n_3245;
assign n_3247 = ~n_3165 &  n_3246;
assign n_3248 =  n_3152 &  n_3247;
assign n_3249 = ~n_3138 &  n_3248;
assign n_3250 = ~n_3125 &  n_3249;
assign n_3251 = ~n_3112 &  n_3250;
assign n_3252 = ~n_3099 &  n_3251;
assign n_3253 = ~n_3086 &  n_3252;
assign n_3254 = ~n_3073 &  n_3253;
assign n_3255 = ~n_3060 &  n_3254;
assign n_3256 = ~n_3047 &  n_3255;
assign n_3257 = ~n_3034 &  n_3256;
assign n_3258 = ~n_3021 &  n_3257;
assign n_3259 = ~n_3008 &  n_3258;
assign n_3260 = ~n_2995 &  n_3259;
assign n_3261 = ~n_2982 &  n_3260;
assign n_3262 = ~n_2969 &  n_3261;
assign n_3263 = ~n_2956 &  n_3262;
assign n_3264 = ~n_2943 &  n_3263;
assign n_3265 = ~n_2930 &  n_3264;
assign n_3266 = ~n_2917 &  n_3265;
assign n_3267 = ~n_2904 &  n_3266;
assign n_3268 = ~n_2891 &  n_3267;
assign n_3269 = ~n_2878 &  n_3268;
assign n_3270 = ~n_2865 &  n_3269;
assign n_3271 = ~n_2852 &  n_3270;
assign n_3272 = ~n_2839 &  n_3271;
assign n_3273 = ~n_2826 &  n_3272;
assign n_3274 = ~n_2813 &  n_3273;
assign n_3275 = ~n_2800 &  n_3274;
assign n_3276 = ~n_2787 &  n_3275;
assign n_3277 = ~n_2774 &  n_3276;
assign n_3278 = ~n_2761 &  n_3277;
assign n_3279 = ~n_2748 &  n_3278;
assign n_3280 = ~n_2735 &  n_3279;
assign n_3281 = ~n_2722 &  n_3280;
assign n_3282 = ~n_2709 &  n_3281;
assign n_3283 = ~n_2696 &  n_3282;
assign n_3284 = ~n_2683 &  n_3283;
assign n_3285 = ~n_2670 &  n_3284;
assign n_3286 = ~n_2657 &  n_3285;
assign n_3287 = ~n_2644 &  n_3286;
assign n_3288 = ~n_2631 &  n_3287;
assign n_3289 = ~n_2618 &  n_3288;
assign n_3290 = ~n_2605 &  n_3289;
assign n_3291 = ~n_2592 &  n_3290;
assign n_3292 = ~n_2579 &  n_3291;
assign n_3293 =  n_2566 &  n_3292;
assign n_3294 = ~n_2494 &  n_3293;
assign n_3295 = ~n_2481 &  n_3294;
assign n_3296 =  n_2481 & ~n_3294;
assign n_3297 = ~n_3295 & ~n_3296;
assign n_3298 =  i_57 & ~n_3297;
assign n_3299 =  n_2494 & ~n_3293;
assign n_3300 = ~n_3294 & ~n_3299;
assign n_3301 = ~i_56 &  n_3300;
assign n_3302 =  i_56 & ~n_3300;
assign n_3303 = ~n_2566 & ~n_3292;
assign n_3304 = ~n_3293 & ~n_3303;
assign n_3305 = ~i_55 &  n_3304;
assign n_3306 =  i_55 & ~n_3304;
assign n_3307 =  n_2579 & ~n_3291;
assign n_3308 = ~n_3292 & ~n_3307;
assign n_3309 = ~i_54 &  n_3308;
assign n_3310 =  i_54 & ~n_3308;
assign n_3311 =  n_2592 & ~n_3290;
assign n_3312 = ~n_3291 & ~n_3311;
assign n_3313 = ~i_53 &  n_3312;
assign n_3314 =  i_53 & ~n_3312;
assign n_3315 =  n_2605 & ~n_3289;
assign n_3316 = ~n_3290 & ~n_3315;
assign n_3317 = ~i_52 &  n_3316;
assign n_3318 =  i_52 & ~n_3316;
assign n_3319 =  n_2618 & ~n_3288;
assign n_3320 = ~n_3289 & ~n_3319;
assign n_3321 = ~i_51 &  n_3320;
assign n_3322 =  i_51 & ~n_3320;
assign n_3323 =  n_2631 & ~n_3287;
assign n_3324 = ~n_3288 & ~n_3323;
assign n_3325 = ~i_50 &  n_3324;
assign n_3326 =  i_50 & ~n_3324;
assign n_3327 =  n_2644 & ~n_3286;
assign n_3328 = ~n_3287 & ~n_3327;
assign n_3329 = ~i_49 &  n_3328;
assign n_3330 =  i_49 & ~n_3328;
assign n_3331 =  n_2657 & ~n_3285;
assign n_3332 = ~n_3286 & ~n_3331;
assign n_3333 = ~i_48 &  n_3332;
assign n_3334 =  i_48 & ~n_3332;
assign n_3335 =  n_2670 & ~n_3284;
assign n_3336 = ~n_3285 & ~n_3335;
assign n_3337 = ~i_47 &  n_3336;
assign n_3338 =  i_47 & ~n_3336;
assign n_3339 =  n_2683 & ~n_3283;
assign n_3340 = ~n_3284 & ~n_3339;
assign n_3341 = ~i_46 &  n_3340;
assign n_3342 =  i_46 & ~n_3340;
assign n_3343 =  n_2696 & ~n_3282;
assign n_3344 = ~n_3283 & ~n_3343;
assign n_3345 = ~i_45 &  n_3344;
assign n_3346 =  i_45 & ~n_3344;
assign n_3347 =  n_2709 & ~n_3281;
assign n_3348 = ~n_3282 & ~n_3347;
assign n_3349 = ~i_44 &  n_3348;
assign n_3350 =  i_44 & ~n_3348;
assign n_3351 =  n_2722 & ~n_3280;
assign n_3352 = ~n_3281 & ~n_3351;
assign n_3353 = ~i_43 &  n_3352;
assign n_3354 =  i_43 & ~n_3352;
assign n_3355 =  n_2735 & ~n_3279;
assign n_3356 = ~n_3280 & ~n_3355;
assign n_3357 = ~i_42 &  n_3356;
assign n_3358 =  i_42 & ~n_3356;
assign n_3359 =  n_2748 & ~n_3278;
assign n_3360 = ~n_3279 & ~n_3359;
assign n_3361 = ~i_41 &  n_3360;
assign n_3362 =  i_41 & ~n_3360;
assign n_3363 =  n_2761 & ~n_3277;
assign n_3364 = ~n_3278 & ~n_3363;
assign n_3365 = ~i_40 &  n_3364;
assign n_3366 =  i_40 & ~n_3364;
assign n_3367 =  n_2774 & ~n_3276;
assign n_3368 = ~n_3277 & ~n_3367;
assign n_3369 = ~i_39 &  n_3368;
assign n_3370 =  i_39 & ~n_3368;
assign n_3371 =  n_2787 & ~n_3275;
assign n_3372 = ~n_3276 & ~n_3371;
assign n_3373 = ~i_38 &  n_3372;
assign n_3374 =  i_38 & ~n_3372;
assign n_3375 =  n_2800 & ~n_3274;
assign n_3376 = ~n_3275 & ~n_3375;
assign n_3377 = ~i_37 &  n_3376;
assign n_3378 =  i_37 & ~n_3376;
assign n_3379 =  n_2813 & ~n_3273;
assign n_3380 = ~n_3274 & ~n_3379;
assign n_3381 = ~i_36 &  n_3380;
assign n_3382 =  i_36 & ~n_3380;
assign n_3383 =  n_2826 & ~n_3272;
assign n_3384 = ~n_3273 & ~n_3383;
assign n_3385 = ~i_35 &  n_3384;
assign n_3386 =  i_35 & ~n_3384;
assign n_3387 =  n_2839 & ~n_3271;
assign n_3388 = ~n_3272 & ~n_3387;
assign n_3389 = ~i_34 &  n_3388;
assign n_3390 =  i_34 & ~n_3388;
assign n_3391 =  n_2852 & ~n_3270;
assign n_3392 = ~n_3271 & ~n_3391;
assign n_3393 = ~i_33 &  n_3392;
assign n_3394 =  i_33 & ~n_3392;
assign n_3395 =  n_2865 & ~n_3269;
assign n_3396 = ~n_3270 & ~n_3395;
assign n_3397 = ~i_32 &  n_3396;
assign n_3398 =  i_32 & ~n_3396;
assign n_3399 =  n_2878 & ~n_3268;
assign n_3400 = ~n_3269 & ~n_3399;
assign n_3401 = ~i_31 &  n_3400;
assign n_3402 =  i_31 & ~n_3400;
assign n_3403 =  n_2891 & ~n_3267;
assign n_3404 = ~n_3268 & ~n_3403;
assign n_3405 = ~i_30 &  n_3404;
assign n_3406 =  i_30 & ~n_3404;
assign n_3407 =  n_2904 & ~n_3266;
assign n_3408 = ~n_3267 & ~n_3407;
assign n_3409 = ~i_29 &  n_3408;
assign n_3410 =  i_29 & ~n_3408;
assign n_3411 =  n_2917 & ~n_3265;
assign n_3412 = ~n_3266 & ~n_3411;
assign n_3413 = ~i_28 &  n_3412;
assign n_3414 =  i_28 & ~n_3412;
assign n_3415 =  n_2930 & ~n_3264;
assign n_3416 = ~n_3265 & ~n_3415;
assign n_3417 = ~i_27 &  n_3416;
assign n_3418 =  i_27 & ~n_3416;
assign n_3419 =  n_2943 & ~n_3263;
assign n_3420 = ~n_3264 & ~n_3419;
assign n_3421 = ~i_26 &  n_3420;
assign n_3422 =  i_26 & ~n_3420;
assign n_3423 =  n_2956 & ~n_3262;
assign n_3424 = ~n_3263 & ~n_3423;
assign n_3425 = ~i_25 &  n_3424;
assign n_3426 =  i_25 & ~n_3424;
assign n_3427 =  n_2969 & ~n_3261;
assign n_3428 = ~n_3262 & ~n_3427;
assign n_3429 = ~i_24 &  n_3428;
assign n_3430 =  i_24 & ~n_3428;
assign n_3431 =  n_2982 & ~n_3260;
assign n_3432 = ~n_3261 & ~n_3431;
assign n_3433 = ~i_23 &  n_3432;
assign n_3434 =  i_23 & ~n_3432;
assign n_3435 =  n_2995 & ~n_3259;
assign n_3436 = ~n_3260 & ~n_3435;
assign n_3437 = ~i_22 &  n_3436;
assign n_3438 =  i_22 & ~n_3436;
assign n_3439 =  n_3008 & ~n_3258;
assign n_3440 = ~n_3259 & ~n_3439;
assign n_3441 = ~i_21 &  n_3440;
assign n_3442 =  i_21 & ~n_3440;
assign n_3443 =  n_3021 & ~n_3257;
assign n_3444 = ~n_3258 & ~n_3443;
assign n_3445 = ~i_20 &  n_3444;
assign n_3446 =  i_20 & ~n_3444;
assign n_3447 =  n_3034 & ~n_3256;
assign n_3448 = ~n_3257 & ~n_3447;
assign n_3449 = ~i_19 &  n_3448;
assign n_3450 =  i_19 & ~n_3448;
assign n_3451 =  n_3047 & ~n_3255;
assign n_3452 = ~n_3256 & ~n_3451;
assign n_3453 = ~i_18 &  n_3452;
assign n_3454 =  i_18 & ~n_3452;
assign n_3455 =  n_3060 & ~n_3254;
assign n_3456 = ~n_3255 & ~n_3455;
assign n_3457 = ~i_17 &  n_3456;
assign n_3458 =  i_17 & ~n_3456;
assign n_3459 =  n_3073 & ~n_3253;
assign n_3460 = ~n_3254 & ~n_3459;
assign n_3461 = ~i_16 &  n_3460;
assign n_3462 =  i_16 & ~n_3460;
assign n_3463 =  n_3086 & ~n_3252;
assign n_3464 = ~n_3253 & ~n_3463;
assign n_3465 = ~i_15 &  n_3464;
assign n_3466 =  i_15 & ~n_3464;
assign n_3467 =  n_3099 & ~n_3251;
assign n_3468 = ~n_3252 & ~n_3467;
assign n_3469 = ~i_14 &  n_3468;
assign n_3470 =  i_14 & ~n_3468;
assign n_3471 =  n_3112 & ~n_3250;
assign n_3472 = ~n_3251 & ~n_3471;
assign n_3473 = ~i_13 &  n_3472;
assign n_3474 =  i_13 & ~n_3472;
assign n_3475 =  n_3125 & ~n_3249;
assign n_3476 = ~n_3250 & ~n_3475;
assign n_3477 = ~i_12 &  n_3476;
assign n_3478 =  i_12 & ~n_3476;
assign n_3479 =  n_3138 & ~n_3248;
assign n_3480 = ~n_3249 & ~n_3479;
assign n_3481 = ~i_11 &  n_3480;
assign n_3482 =  i_11 & ~n_3480;
assign n_3483 = ~n_3152 & ~n_3247;
assign n_3484 = ~n_3248 & ~n_3483;
assign n_3485 = ~i_10 &  n_3484;
assign n_3486 =  i_10 & ~n_3484;
assign n_3487 =  n_3165 & ~n_3246;
assign n_3488 = ~n_3247 & ~n_3487;
assign n_3489 = ~i_9 &  n_3488;
assign n_3490 =  i_9 & ~n_3488;
assign n_3491 =  n_3178 & ~n_3245;
assign n_3492 = ~n_3246 & ~n_3491;
assign n_3493 = ~i_8 &  n_3492;
assign n_3494 =  i_8 & ~n_3492;
assign n_3495 = ~n_3192 & ~n_3244;
assign n_3496 = ~n_3245 & ~n_3495;
assign n_3497 = ~i_7 &  n_3496;
assign n_3498 =  i_7 & ~n_3496;
assign n_3499 =  n_3205 & ~n_3243;
assign n_3500 = ~n_3244 & ~n_3499;
assign n_3501 = ~i_6 &  n_3500;
assign n_3502 =  i_6 & ~n_3500;
assign n_3503 = ~n_3219 & ~n_3242;
assign n_3504 = ~n_3243 & ~n_3503;
assign n_3505 = ~i_5 &  n_3504;
assign n_3506 =  i_5 & ~n_3504;
assign n_3507 =  n_3232 & ~n_3241;
assign n_3508 = ~n_3242 & ~n_3507;
assign n_3509 = ~i_4 &  n_3508;
assign n_3510 =  i_4 & ~n_3508;
assign n_3511 = ~n_3233 &  n_3240;
assign n_3512 = ~n_3233 & ~n_3239;
assign n_3513 = ~n_3236 & ~n_3512;
assign n_3514 = ~n_3511 &  n_3513;
assign n_3515 = ~i_3 & ~n_3514;
assign n_3516 = ~n_3236 & ~n_3240;
assign n_3517 =  n_3233 & ~n_3516;
assign n_3518 =  n_3233 &  n_3234;
assign n_3519 = ~n_3512 & ~n_3518;
assign n_3520 = ~n_3517 &  n_3519;
assign n_3521 = ~n_2552 & ~n_3520;
assign n_3522 =  i_1 &  n_3521;
assign n_3523 = ~i_2 & ~n_3522;
assign n_3524 = ~n_3233 & ~n_3237;
assign n_3525 = ~n_3517 &  n_3521;
assign n_3526 = ~n_3524 & ~n_3525;
assign n_3527 = ~n_3523 &  n_3526;
assign n_3528 =  i_3 &  n_3514;
assign n_3529 =  i_2 &  n_3522;
assign n_3530 = ~n_3528 & ~n_3529;
assign n_3531 = ~n_3527 &  n_3530;
assign n_3532 = ~n_3515 & ~n_3531;
assign n_3533 = ~n_3510 & ~n_3532;
assign n_3534 = ~n_3509 & ~n_3533;
assign n_3535 = ~n_3506 & ~n_3534;
assign n_3536 = ~n_3505 & ~n_3535;
assign n_3537 = ~n_3502 & ~n_3536;
assign n_3538 = ~n_3501 & ~n_3537;
assign n_3539 = ~n_3498 & ~n_3538;
assign n_3540 = ~n_3497 & ~n_3539;
assign n_3541 = ~n_3494 & ~n_3540;
assign n_3542 = ~n_3493 & ~n_3541;
assign n_3543 = ~n_3490 & ~n_3542;
assign n_3544 = ~n_3489 & ~n_3543;
assign n_3545 = ~n_3486 & ~n_3544;
assign n_3546 = ~n_3485 & ~n_3545;
assign n_3547 = ~n_3482 & ~n_3546;
assign n_3548 = ~n_3481 & ~n_3547;
assign n_3549 = ~n_3478 & ~n_3548;
assign n_3550 = ~n_3477 & ~n_3549;
assign n_3551 = ~n_3474 & ~n_3550;
assign n_3552 = ~n_3473 & ~n_3551;
assign n_3553 = ~n_3470 & ~n_3552;
assign n_3554 = ~n_3469 & ~n_3553;
assign n_3555 = ~n_3466 & ~n_3554;
assign n_3556 = ~n_3465 & ~n_3555;
assign n_3557 = ~n_3462 & ~n_3556;
assign n_3558 = ~n_3461 & ~n_3557;
assign n_3559 = ~n_3458 & ~n_3558;
assign n_3560 = ~n_3457 & ~n_3559;
assign n_3561 = ~n_3454 & ~n_3560;
assign n_3562 = ~n_3453 & ~n_3561;
assign n_3563 = ~n_3450 & ~n_3562;
assign n_3564 = ~n_3449 & ~n_3563;
assign n_3565 = ~n_3446 & ~n_3564;
assign n_3566 = ~n_3445 & ~n_3565;
assign n_3567 = ~n_3442 & ~n_3566;
assign n_3568 = ~n_3441 & ~n_3567;
assign n_3569 = ~n_3438 & ~n_3568;
assign n_3570 = ~n_3437 & ~n_3569;
assign n_3571 = ~n_3434 & ~n_3570;
assign n_3572 = ~n_3433 & ~n_3571;
assign n_3573 = ~n_3430 & ~n_3572;
assign n_3574 = ~n_3429 & ~n_3573;
assign n_3575 = ~n_3426 & ~n_3574;
assign n_3576 = ~n_3425 & ~n_3575;
assign n_3577 = ~n_3422 & ~n_3576;
assign n_3578 = ~n_3421 & ~n_3577;
assign n_3579 = ~n_3418 & ~n_3578;
assign n_3580 = ~n_3417 & ~n_3579;
assign n_3581 = ~n_3414 & ~n_3580;
assign n_3582 = ~n_3413 & ~n_3581;
assign n_3583 = ~n_3410 & ~n_3582;
assign n_3584 = ~n_3409 & ~n_3583;
assign n_3585 = ~n_3406 & ~n_3584;
assign n_3586 = ~n_3405 & ~n_3585;
assign n_3587 = ~n_3402 & ~n_3586;
assign n_3588 = ~n_3401 & ~n_3587;
assign n_3589 = ~n_3398 & ~n_3588;
assign n_3590 = ~n_3397 & ~n_3589;
assign n_3591 = ~n_3394 & ~n_3590;
assign n_3592 = ~n_3393 & ~n_3591;
assign n_3593 = ~n_3390 & ~n_3592;
assign n_3594 = ~n_3389 & ~n_3593;
assign n_3595 = ~n_3386 & ~n_3594;
assign n_3596 = ~n_3385 & ~n_3595;
assign n_3597 = ~n_3382 & ~n_3596;
assign n_3598 = ~n_3381 & ~n_3597;
assign n_3599 = ~n_3378 & ~n_3598;
assign n_3600 = ~n_3377 & ~n_3599;
assign n_3601 = ~n_3374 & ~n_3600;
assign n_3602 = ~n_3373 & ~n_3601;
assign n_3603 = ~n_3370 & ~n_3602;
assign n_3604 = ~n_3369 & ~n_3603;
assign n_3605 = ~n_3366 & ~n_3604;
assign n_3606 = ~n_3365 & ~n_3605;
assign n_3607 = ~n_3362 & ~n_3606;
assign n_3608 = ~n_3361 & ~n_3607;
assign n_3609 = ~n_3358 & ~n_3608;
assign n_3610 = ~n_3357 & ~n_3609;
assign n_3611 = ~n_3354 & ~n_3610;
assign n_3612 = ~n_3353 & ~n_3611;
assign n_3613 = ~n_3350 & ~n_3612;
assign n_3614 = ~n_3349 & ~n_3613;
assign n_3615 = ~n_3346 & ~n_3614;
assign n_3616 = ~n_3345 & ~n_3615;
assign n_3617 = ~n_3342 & ~n_3616;
assign n_3618 = ~n_3341 & ~n_3617;
assign n_3619 = ~n_3338 & ~n_3618;
assign n_3620 = ~n_3337 & ~n_3619;
assign n_3621 = ~n_3334 & ~n_3620;
assign n_3622 = ~n_3333 & ~n_3621;
assign n_3623 = ~n_3330 & ~n_3622;
assign n_3624 = ~n_3329 & ~n_3623;
assign n_3625 = ~n_3326 & ~n_3624;
assign n_3626 = ~n_3325 & ~n_3625;
assign n_3627 = ~n_3322 & ~n_3626;
assign n_3628 = ~n_3321 & ~n_3627;
assign n_3629 = ~n_3318 & ~n_3628;
assign n_3630 = ~n_3317 & ~n_3629;
assign n_3631 = ~n_3314 & ~n_3630;
assign n_3632 = ~n_3313 & ~n_3631;
assign n_3633 = ~n_3310 & ~n_3632;
assign n_3634 = ~n_3309 & ~n_3633;
assign n_3635 = ~n_3306 & ~n_3634;
assign n_3636 = ~n_3305 & ~n_3635;
assign n_3637 = ~n_3302 & ~n_3636;
assign n_3638 = ~n_3301 & ~n_3637;
assign n_3639 = ~n_3298 & ~n_3638;
assign n_3640 = ~i_57 &  n_3297;
assign n_3641 = ~n_2413 &  n_2463;
assign n_3642 = ~n_2469 & ~n_2475;
assign n_3643 = ~n_3641 &  n_3642;
assign n_3644 = ~n_2552 & ~n_3643;
assign n_3645 =  n_3295 &  n_3644;
assign n_3646 = ~n_3295 & ~n_3644;
assign n_3647 = ~n_3645 & ~n_3646;
assign n_3648 = ~i_58 &  n_3647;
assign n_3649 = ~n_3640 & ~n_3648;
assign n_3650 = ~n_3639 &  n_3649;
assign n_3651 =  i_58 & ~n_3647;
assign n_3652 = ~n_2454 & ~n_2460;
assign n_3653 = ~n_2415 & ~n_3652;
assign n_3654 = ~n_2461 & ~n_3653;
assign n_3655 =  n_3645 & ~n_3654;
assign n_3656 = ~n_2552 & ~n_3654;
assign n_3657 = ~n_3645 & ~n_3656;
assign n_3658 = ~n_3655 & ~n_3657;
assign n_3659 =  i_59 & ~n_3658;
assign n_3660 = ~n_3651 & ~n_3659;
assign n_3661 = ~n_3650 &  n_3660;
assign n_3662 = ~i_59 &  n_3658;
assign n_3663 = ~n_2452 & ~n_2457;
assign n_3664 = ~n_2552 & ~n_3663;
assign n_3665 = ~n_3655 &  n_3664;
assign n_3666 =  n_3655 & ~n_3664;
assign n_3667 = ~n_3665 & ~n_3666;
assign n_3668 = ~i_60 & ~n_3667;
assign n_3669 = ~n_3662 & ~n_3668;
assign n_3670 = ~n_3661 &  n_3669;
assign n_3671 = ~i_11 & ~i_12;
assign n_3672 = ~i_13 & ~i_14;
assign n_3673 = ~i_15 & ~i_16;
assign n_3674 =  n_3672 &  n_3673;
assign n_3675 =  n_3671 &  n_3674;
assign n_3676 = ~i_21 & ~i_22;
assign n_3677 = ~i_23 & ~i_24;
assign n_3678 =  n_3676 &  n_3677;
assign n_3679 = ~i_17 & ~i_18;
assign n_3680 = ~i_19 & ~i_20;
assign n_3681 =  n_3679 &  n_3680;
assign n_3682 =  n_3678 &  n_3681;
assign n_3683 = ~i_29 & ~i_30;
assign n_3684 = ~i_31 & ~i_32;
assign n_3685 =  n_3683 &  n_3684;
assign n_3686 = ~i_25 & ~i_26;
assign n_3687 = ~i_27 & ~i_28;
assign n_3688 =  n_3686 &  n_3687;
assign n_3689 =  n_3685 &  n_3688;
assign n_3690 =  n_3682 &  n_3689;
assign n_3691 =  n_3675 &  n_3690;
assign n_3692 = ~i_57 & ~i_58;
assign n_3693 = ~i_59 & ~i_60;
assign n_3694 =  n_3692 &  n_3693;
assign n_3695 = ~i_53 & ~i_54;
assign n_3696 = ~i_55 & ~i_56;
assign n_3697 =  n_3695 &  n_3696;
assign n_3698 = ~i_49 & ~i_50;
assign n_3699 = ~i_51 & ~i_52;
assign n_3700 =  n_3698 &  n_3699;
assign n_3701 =  n_3697 &  n_3700;
assign n_3702 =  n_3694 &  n_3701;
assign n_3703 = ~i_37 & ~i_38;
assign n_3704 = ~i_39 & ~i_40;
assign n_3705 =  n_3703 &  n_3704;
assign n_3706 = ~i_33 & ~i_34;
assign n_3707 = ~i_35 & ~i_36;
assign n_3708 =  n_3706 &  n_3707;
assign n_3709 =  n_3705 &  n_3708;
assign n_3710 = ~i_45 & ~i_46;
assign n_3711 = ~i_47 & ~i_48;
assign n_3712 =  n_3710 &  n_3711;
assign n_3713 = ~i_41 & ~i_42;
assign n_3714 = ~i_43 & ~i_44;
assign n_3715 =  n_3713 &  n_3714;
assign n_3716 =  n_3712 &  n_3715;
assign n_3717 =  n_3709 &  n_3716;
assign n_3718 =  n_3702 &  n_3717;
assign n_3719 =  n_3691 &  n_3718;
assign n_3720 = ~n_3670 &  n_3719;
assign n_3721 =  i_9 &  n_3720;
assign n_3722 =  i_10 &  n_3720;
assign n_3723 =  i_8 &  n_3720;
assign n_3724 = ~n_3722 & ~n_3723;
assign n_3725 = ~n_3721 &  n_3724;
assign n_3726 = ~i_1 & ~i_2;
assign n_3727 =  n_3720 & ~n_3726;
assign n_3728 =  i_3 &  n_3720;
assign n_3729 = ~n_3727 & ~n_3728;
assign n_3730 =  i_6 &  n_3720;
assign n_3731 =  i_4 &  n_3720;
assign n_3732 = ~n_3730 & ~n_3731;
assign n_3733 =  i_5 &  n_3720;
assign n_3734 =  i_7 &  n_3720;
assign n_3735 = ~n_3733 & ~n_3734;
assign n_3736 =  n_3732 &  n_3735;
assign n_3737 =  n_3729 &  n_3736;
assign n_3738 =  n_3725 &  n_3737;
assign n_3739 =  i_1 &  i_3;
assign n_3740 =  n_3727 & ~n_3739;
assign n_3741 =  i_2 &  n_3720;
assign n_3742 =  i_1 &  n_3741;
assign n_3743 =  i_3 &  n_3727;
assign n_3744 = ~n_3742 &  n_3743;
assign n_3745 = ~i_3 &  n_3742;
assign n_3746 = ~n_3745 & ~n_3729;
assign n_3747 = ~n_3744 &  n_3746;
assign n_3748 =  n_3740 &  n_3747;
assign n_3749 = ~n_3747 & ~n_3731;
assign n_3750 = ~n_3748 & ~n_3749;
assign n_3751 = ~n_3740 &  n_3731;
assign n_3752 = ~i_4 &  n_3740;
assign n_3753 = ~n_3751 & ~n_3752;
assign n_3754 =  n_3747 & ~n_3753;
assign n_3755 = ~n_3747 &  n_3753;
assign n_3756 = ~n_3754 & ~n_3755;
assign n_3757 =  n_3750 & ~n_3756;
assign n_3758 =  n_3756 &  n_3733;
assign n_3759 = ~n_3757 & ~n_3758;
assign n_3760 = ~n_3730 & ~n_3759;
assign n_3761 =  n_3730 &  n_3759;
assign n_3762 = ~n_3760 & ~n_3761;
assign n_3763 = ~n_3750 &  n_3756;
assign n_3764 = ~n_3757 & ~n_3763;
assign n_3765 =  n_3733 & ~n_3764;
assign n_3766 = ~n_3733 &  n_3764;
assign n_3767 = ~n_3765 & ~n_3766;
assign n_3768 =  n_3762 & ~n_3767;
assign n_3769 = ~n_3762 &  n_3767;
assign n_3770 = ~n_3768 & ~n_3769;
assign n_3771 = ~n_3730 & ~n_3765;
assign n_3772 = ~n_3766 & ~n_3771;
assign n_3773 = ~n_3770 & ~n_3772;
assign n_3774 =  n_3770 & ~n_3734;
assign n_3775 = ~n_3773 & ~n_3774;
assign n_3776 = ~n_3723 &  n_3775;
assign n_3777 =  n_3723 & ~n_3775;
assign n_3778 = ~n_3776 & ~n_3777;
assign n_3779 = ~n_3770 &  n_3734;
assign n_3780 = ~n_3774 & ~n_3779;
assign n_3781 = ~n_3772 & ~n_3780;
assign n_3782 =  n_3772 &  n_3780;
assign n_3783 = ~n_3781 & ~n_3782;
assign n_3784 =  n_3778 & ~n_3783;
assign n_3785 = ~n_3778 &  n_3783;
assign n_3786 = ~n_3784 & ~n_3785;
assign n_3787 = ~n_3723 & ~n_3783;
assign n_3788 = ~n_3775 &  n_3783;
assign n_3789 = ~n_3787 & ~n_3788;
assign n_3790 =  n_3786 &  n_3789;
assign n_3791 = ~n_3786 &  n_3721;
assign n_3792 = ~n_3790 & ~n_3791;
assign n_3793 = ~n_3722 & ~n_3792;
assign n_3794 =  n_3722 &  n_3792;
assign n_3795 = ~n_3793 & ~n_3794;
assign n_3796 = ~n_3786 & ~n_3789;
assign n_3797 = ~n_3790 & ~n_3796;
assign n_3798 =  n_3721 & ~n_3797;
assign n_3799 = ~n_3721 &  n_3797;
assign n_3800 = ~n_3798 & ~n_3799;
assign n_3801 =  n_3795 & ~n_3800;
assign n_3802 = ~n_3795 &  n_3800;
assign n_3803 = ~n_3801 & ~n_3802;
assign n_3804 = ~i_9 &  n_3797;
assign n_3805 = ~n_3722 & ~n_3798;
assign n_3806 = ~n_3804 & ~n_3805;
assign n_3807 =  n_3803 & ~n_3806;
assign n_3808 = ~n_3803 & ~n_3806;
assign n_3809 =  n_3792 &  n_3800;
assign n_3810 = ~n_3793 & ~n_3809;
assign n_3811 = ~n_3748 & ~n_3751;
assign n_3812 =  n_3759 &  n_3767;
assign n_3813 = ~n_3760 & ~n_3812;
assign n_3814 =  n_3811 & ~n_3813;
assign n_3815 = ~n_3811 &  n_3813;
assign n_3816 = ~n_3814 & ~n_3815;
assign n_3817 =  n_3807 & ~n_3816;
assign n_3818 = ~n_3776 & ~n_3781;
assign n_3819 =  n_3816 & ~n_3818;
assign n_3820 = ~n_3817 & ~n_3819;
assign n_3821 =  n_3807 &  n_3814;
assign n_3822 =  n_3818 &  n_3821;
assign n_3823 = ~n_3811 & ~n_3818;
assign n_3824 = ~n_3807 &  n_3823;
assign n_3825 = ~n_3816 & ~n_3824;
assign n_3826 = ~n_3822 &  n_3825;
assign n_3827 = ~n_3820 &  n_3826;
assign n_3828 =  n_3820 & ~n_3826;
assign n_3829 = ~n_3827 & ~n_3828;
assign n_3830 =  n_3810 &  n_3829;
assign n_3831 =  n_3807 & ~n_3830;
assign n_3832 = ~n_3810 & ~n_3829;
assign n_3833 =  n_3831 & ~n_3832;
assign n_3834 = ~n_3810 & ~n_3826;
assign n_3835 = ~n_3827 & ~n_3834;
assign n_3836 =  n_3833 & ~n_3835;
assign n_3837 =  n_3722 & ~n_3800;
assign n_3838 = ~n_3809 & ~n_3837;
assign n_3839 = ~n_3807 &  n_3810;
assign n_3840 = ~n_3828 &  n_3839;
assign n_3841 =  n_3835 & ~n_3840;
assign n_3842 = ~n_3833 &  n_3841;
assign n_3843 = ~n_3807 &  n_3815;
assign n_3844 =  n_3807 & ~n_3815;
assign n_3845 = ~n_3814 & ~n_3844;
assign n_3846 = ~n_3843 &  n_3845;
assign n_3847 = ~n_3821 & ~n_3846;
assign n_3848 =  n_3818 &  n_3847;
assign n_3849 = ~n_3807 &  n_3818;
assign n_3850 = ~n_3843 & ~n_3849;
assign n_3851 = ~n_3810 & ~n_3850;
assign n_3852 = ~n_3848 &  n_3851;
assign n_3853 = ~n_3836 & ~n_3852;
assign n_3854 = ~n_3842 &  n_3853;
assign n_3855 =  n_3838 &  n_3854;
assign n_3856 = ~n_3831 & ~n_3852;
assign n_3857 = ~n_3838 & ~n_3854;
assign n_3858 =  n_3856 & ~n_3857;
assign n_3859 = ~n_3855 &  n_3858;
assign n_3860 = ~n_3836 & ~n_3859;
assign n_3861 =  n_3808 & ~n_3860;
assign n_3862 = ~n_3831 &  n_3854;
assign n_3863 =  n_3807 & ~n_3838;
assign n_3864 = ~n_3862 &  n_3863;
assign n_3865 = ~n_3808 & ~n_3864;
assign n_3866 = ~n_3836 & ~n_3865;
assign n_3867 = ~n_3861 &  n_3866;
assign n_3868 =  n_3789 & ~n_3721;
assign n_3869 = ~n_3796 & ~n_3868;
assign n_3870 =  n_3859 &  n_3865;
assign n_3871 = ~n_3856 &  n_3857;
assign n_3872 =  n_3864 & ~n_3871;
assign n_3873 = ~n_3859 &  n_3872;
assign n_3874 = ~n_3836 & ~n_3873;
assign n_3875 = ~n_3870 &  n_3874;
assign n_3876 = ~n_3869 & ~n_3875;
assign n_3877 =  n_3869 &  n_3875;
assign n_3878 = ~n_3876 & ~n_3877;
assign n_3879 = ~n_3867 &  n_3878;
assign n_3880 =  n_3867 & ~n_3878;
assign n_3881 = ~n_3879 & ~n_3880;
assign n_3882 = ~n_3807 & ~n_3881;
assign n_3883 = ~n_3867 &  n_3876;
assign n_3884 = ~n_3873 & ~n_3883;
assign n_3885 = ~n_3882 &  n_3884;
assign n_3886 = ~n_3867 & ~n_3869;
assign n_3887 =  n_3875 &  n_3886;
assign n_3888 = ~n_3873 & ~n_3886;
assign n_3889 =  n_3807 & ~n_3888;
assign n_3890 =  n_3881 &  n_3889;
assign n_3891 = ~n_3887 & ~n_3890;
assign n_3892 = ~n_3885 &  n_3891;
assign n_3893 =  n_3867 & ~n_3875;
assign n_3894 = ~n_3869 &  n_3893;
assign n_3895 =  n_3892 &  n_3894;
assign n_3896 =  n_3772 &  n_3734;
assign n_3897 = ~n_3773 & ~n_3896;
assign n_3898 =  n_3891 & ~n_3894;
assign n_3899 = ~n_3897 &  n_3898;
assign n_3900 = ~n_3895 & ~n_3899;
assign n_3901 =  n_3897 & ~n_3892;
assign n_3902 = ~n_3901 & ~n_3894;
assign n_3903 =  n_3885 &  n_3898;
assign n_3904 = ~n_3903 & ~n_3895;
assign n_3905 = ~n_3897 &  n_3904;
assign n_3906 =  n_3897 & ~n_3904;
assign n_3907 = ~n_3905 & ~n_3906;
assign n_3908 = ~n_3902 & ~n_3907;
assign n_3909 =  n_3807 &  n_3907;
assign n_3910 = ~n_3908 & ~n_3909;
assign n_3911 = ~n_3807 &  n_3902;
assign n_3912 =  n_3807 & ~n_3902;
assign n_3913 = ~n_3911 & ~n_3912;
assign n_3914 =  n_3907 &  n_3913;
assign n_3915 = ~n_3907 & ~n_3913;
assign n_3916 = ~n_3914 & ~n_3915;
assign n_3917 = ~n_3910 & ~n_3916;
assign n_3918 =  n_3750 & ~n_3733;
assign n_3919 = ~n_3763 & ~n_3918;
assign n_3920 =  n_3910 &  n_3919;
assign n_3921 = ~n_3917 & ~n_3920;
assign n_3922 =  n_3818 &  n_3845;
assign n_3923 = ~n_3821 & ~n_3922;
assign n_3924 = ~n_3741 & ~n_3728;
assign n_3925 = ~n_3742 & ~n_3924;
assign n_3926 =  n_3910 &  n_3916;
assign n_3927 = ~n_3917 & ~n_3926;
assign n_3928 = ~n_3919 & ~n_3927;
assign n_3929 =  n_3807 & ~n_3928;
assign n_3930 =  n_3919 &  n_3927;
assign n_3931 = ~n_3928 & ~n_3930;
assign n_3932 =  n_3916 & ~n_3919;
assign n_3933 = ~n_3807 & ~n_3932;
assign n_3934 = ~n_3931 &  n_3933;
assign n_3935 = ~n_3929 & ~n_3934;
assign n_3936 =  n_3925 & ~n_3935;
assign n_3937 = ~n_3917 & ~n_3932;
assign n_3938 =  n_3807 & ~n_3937;
assign n_3939 = ~n_3933 & ~n_3938;
assign n_3940 =  n_3931 & ~n_3939;
assign n_3941 = ~n_3931 &  n_3939;
assign n_3942 = ~n_3940 & ~n_3941;
assign n_3943 = ~n_3925 &  n_3942;
assign n_3944 = ~n_3936 & ~n_3943;
assign n_3945 = ~n_3807 &  n_3813;
assign n_3946 =  n_3807 &  n_3811;
assign n_3947 = ~n_3945 & ~n_3946;
assign n_3948 =  n_3944 &  n_3947;
assign n_3949 = ~n_3944 & ~n_3947;
assign n_3950 = ~n_3948 & ~n_3949;
assign n_3951 =  n_3923 & ~n_3950;
assign n_3952 = ~n_3923 &  n_3950;
assign n_3953 = ~n_3951 & ~n_3952;
assign n_3954 =  n_3935 & ~n_3942;
assign n_3955 = ~n_3947 & ~n_3954;
assign n_3956 = ~n_3943 & ~n_3955;
assign n_3957 =  n_3953 &  n_3956;
assign n_3958 = ~n_3953 & ~n_3956;
assign n_3959 = ~n_3957 & ~n_3958;
assign n_3960 =  n_3921 & ~n_3959;
assign n_3961 = ~n_3949 & ~n_3956;
assign n_3962 = ~n_3951 & ~n_3961;
assign n_3963 = ~n_3958 & ~n_3962;
assign n_3964 = ~n_3960 & ~n_3963;
assign n_3965 =  n_3810 &  n_3820;
assign n_3966 = ~n_3827 & ~n_3965;
assign n_3967 =  n_3964 & ~n_3966;
assign n_3968 = ~n_3964 &  n_3966;
assign n_3969 = ~n_3967 & ~n_3968;
assign n_3970 = ~n_3921 &  n_3959;
assign n_3971 = ~n_3960 & ~n_3970;
assign n_3972 = ~n_3962 & ~n_3971;
assign n_3973 =  n_3962 &  n_3971;
assign n_3974 = ~n_3972 & ~n_3973;
assign n_3975 =  n_3969 &  n_3974;
assign n_3976 = ~n_3969 & ~n_3974;
assign n_3977 = ~n_3975 & ~n_3976;
assign n_3978 = ~n_3900 &  n_3977;
assign n_3979 = ~n_3964 & ~n_3972;
assign n_3980 =  n_3966 & ~n_3974;
assign n_3981 = ~n_3979 & ~n_3980;
assign n_3982 = ~n_3977 & ~n_3981;
assign n_3983 = ~n_3978 & ~n_3982;
assign n_3984 =  n_3838 &  n_3856;
assign n_3985 = ~n_3838 & ~n_3856;
assign n_3986 = ~n_3984 & ~n_3985;
assign n_3987 = ~n_3857 & ~n_3986;
assign n_3988 =  n_3983 & ~n_3987;
assign n_3989 = ~n_3877 & ~n_3893;
assign n_3990 =  n_3900 & ~n_3977;
assign n_3991 = ~n_3978 & ~n_3990;
assign n_3992 =  n_3981 &  n_3991;
assign n_3993 = ~n_3981 & ~n_3991;
assign n_3994 = ~n_3992 & ~n_3993;
assign n_3995 = ~n_3987 & ~n_3994;
assign n_3996 =  n_3977 & ~n_3981;
assign n_3997 = ~n_3990 & ~n_3996;
assign n_3998 = ~n_3993 & ~n_3997;
assign n_3999 = ~n_3995 & ~n_3998;
assign n_4000 = ~n_3989 &  n_3999;
assign n_4001 = ~n_3988 & ~n_4000;
assign n_4002 = ~n_3983 &  n_3987;
assign n_4003 = ~n_3988 & ~n_3989;
assign n_4004 = ~n_4002 & ~n_4003;
assign n_4005 =  n_3989 & ~n_3999;
assign n_4006 = ~n_4000 & ~n_4005;
assign n_4007 = ~n_4002 & ~n_3988;
assign n_4008 =  n_4006 &  n_4007;
assign n_4009 = ~n_4006 & ~n_4007;
assign n_4010 = ~n_4008 & ~n_4009;
assign n_4011 =  n_4004 & ~n_4010;
assign n_4012 = ~n_3807 & ~n_3852;
assign n_4013 =  n_3857 &  n_4012;
assign n_4014 = ~n_3836 & ~n_4013;
assign n_4015 =  n_4010 & ~n_4014;
assign n_4016 = ~n_4011 & ~n_4015;
assign n_4017 = ~n_3861 & ~n_3866;
assign n_4018 =  n_4016 & ~n_4017;
assign n_4019 = ~n_4004 &  n_4014;
assign n_4020 =  n_4004 & ~n_4014;
assign n_4021 = ~n_4019 & ~n_4020;
assign n_4022 =  n_4010 &  n_4021;
assign n_4023 = ~n_4010 & ~n_4021;
assign n_4024 = ~n_4022 & ~n_4023;
assign n_4025 = ~n_4016 &  n_4017;
assign n_4026 = ~n_4024 &  n_4025;
assign n_4027 = ~n_4018 & ~n_4026;
assign n_4028 = ~n_3807 &  n_3884;
assign n_4029 = ~n_3887 & ~n_3894;
assign n_4030 = ~n_4028 &  n_4029;
assign n_4031 =  n_4018 &  n_4024;
assign n_4032 =  n_4016 & ~n_4024;
assign n_4033 =  n_4017 &  n_4032;
assign n_4034 = ~n_4031 & ~n_4033;
assign n_4035 =  n_4024 &  n_4025;
assign n_4036 =  n_4034 & ~n_4035;
assign n_4037 =  n_3836 &  n_4036;
assign n_4038 =  n_4030 & ~n_4037;
assign n_4039 =  n_3836 & ~n_4036;
assign n_4040 = ~n_3836 &  n_3865;
assign n_4041 = ~n_4032 &  n_4040;
assign n_4042 =  n_4036 &  n_4041;
assign n_4043 = ~n_4039 & ~n_4042;
assign n_4044 =  n_3871 & ~n_4037;
assign n_4045 =  n_3807 &  n_3937;
assign n_4046 = ~n_3928 & ~n_4045;
assign n_4047 = ~n_3908 & ~n_3911;
assign n_4048 = ~n_3871 & ~n_4034;
assign n_4049 = ~n_3836 &  n_3871;
assign n_4050 =  n_4034 &  n_4049;
assign n_4051 = ~n_4048 & ~n_4050;
assign n_4052 = ~n_4039 &  n_4051;
assign n_4053 = ~n_4052 &  n_4030;
assign n_4054 = ~n_4053 & ~n_4037;
assign n_4055 = ~n_4034 &  n_4049;
assign n_4056 = ~n_4039 & ~n_4055;
assign n_4057 =  n_3807 &  n_3832;
assign n_4058 = ~n_3807 &  n_3835;
assign n_4059 = ~n_3852 & ~n_4058;
assign n_4060 = ~n_4057 &  n_4059;
assign n_4061 =  n_4056 & ~n_4060;
assign n_4062 =  n_4052 & ~n_4030;
assign n_4063 =  n_4054 & ~n_4062;
assign n_4064 =  n_4061 & ~n_4063;
assign n_4065 = ~n_4054 &  n_4064;
assign n_4066 =  n_4054 &  n_4061;
assign n_4067 =  n_4063 &  n_4066;
assign n_4068 =  n_4056 &  n_4060;
assign n_4069 =  n_4062 &  n_4068;
assign n_4070 = ~n_4039 & ~n_4069;
assign n_4071 = ~n_4067 &  n_4070;
assign n_4072 = ~n_4065 &  n_4071;
assign n_4073 =  n_4047 & ~n_4072;
assign n_4074 =  n_4063 &  n_4068;
assign n_4075 = ~n_4054 &  n_4068;
assign n_4076 = ~n_4039 & ~n_4075;
assign n_4077 = ~n_4074 &  n_4076;
assign n_4078 = ~n_4065 &  n_4077;
assign n_4079 =  n_4072 & ~n_4078;
assign n_4080 = ~n_4073 & ~n_4079;
assign n_4081 = ~n_3818 & ~n_3847;
assign n_4082 =  n_3850 & ~n_4081;
assign n_4083 = ~n_4047 &  n_4072;
assign n_4084 = ~n_4073 & ~n_4083;
assign n_4085 =  n_4078 &  n_4084;
assign n_4086 = ~n_4078 & ~n_4084;
assign n_4087 = ~n_4085 & ~n_4086;
assign n_4088 =  n_4082 & ~n_4087;
assign n_4089 = ~n_4082 &  n_4087;
assign n_4090 = ~n_4088 & ~n_4089;
assign n_4091 =  n_4080 &  n_4090;
assign n_4092 = ~n_4080 & ~n_4090;
assign n_4093 = ~n_4091 & ~n_4092;
assign n_4094 =  n_4046 & ~n_4093;
assign n_4095 = ~n_4080 & ~n_4086;
assign n_4096 = ~n_4088 & ~n_4095;
assign n_4097 = ~n_4092 & ~n_4096;
assign n_4098 = ~n_4094 & ~n_4097;
assign n_4099 = ~n_4046 &  n_4096;
assign n_4100 =  n_4046 & ~n_4096;
assign n_4101 = ~n_4099 & ~n_4100;
assign n_4102 = ~n_4093 &  n_4101;
assign n_4103 =  n_4093 & ~n_4101;
assign n_4104 = ~n_4102 & ~n_4103;
assign n_4105 = ~n_4098 & ~n_4104;
assign n_4106 =  n_3807 & ~n_3814;
assign n_4107 =  n_4098 & ~n_4106;
assign n_4108 = ~n_4105 & ~n_4107;
assign n_4109 = ~n_3807 &  n_3811;
assign n_4110 =  n_4104 &  n_4106;
assign n_4111 = ~n_4105 & ~n_4110;
assign n_4112 = ~n_4098 &  n_4106;
assign n_4113 = ~n_4107 & ~n_4112;
assign n_4114 =  n_4104 &  n_4113;
assign n_4115 = ~n_4104 & ~n_4113;
assign n_4116 = ~n_4114 & ~n_4115;
assign n_4117 = ~n_4111 & ~n_4116;
assign n_4118 =  n_4111 &  n_4116;
assign n_4119 = ~n_4117 & ~n_4118;
assign n_4120 = ~n_3925 &  n_3935;
assign n_4121 = ~n_3936 & ~n_4120;
assign n_4122 =  n_3942 &  n_4121;
assign n_4123 = ~n_3942 & ~n_4121;
assign n_4124 = ~n_4122 & ~n_4123;
assign n_4125 = ~n_4119 & ~n_4124;
assign n_4126 =  n_4119 &  n_4124;
assign n_4127 = ~n_4125 & ~n_4126;
assign n_4128 = ~n_4109 &  n_4127;
assign n_4129 = ~n_3923 &  n_3956;
assign n_4130 = ~n_3961 & ~n_4129;
assign n_4131 = ~n_4125 & ~n_4130;
assign n_4132 = ~n_4128 & ~n_4131;
assign n_4133 =  n_4116 & ~n_4124;
assign n_4134 = ~n_4117 & ~n_4133;
assign n_4135 =  n_4109 &  n_4134;
assign n_4136 = ~n_4128 & ~n_4135;
assign n_4137 = ~n_4130 &  n_4136;
assign n_4138 = ~n_4125 &  n_4130;
assign n_4139 = ~n_4136 &  n_4138;
assign n_4140 = ~n_4137 & ~n_4139;
assign n_4141 = ~n_4132 &  n_4140;
assign n_4142 = ~n_3967 & ~n_3979;
assign n_4143 = ~n_4142 & ~n_4140;
assign n_4144 = ~n_4141 & ~n_4143;
assign n_4145 =  n_4108 &  n_4144;
assign n_4146 =  n_3987 &  n_3997;
assign n_4147 = ~n_3998 & ~n_4146;
assign n_4148 = ~n_4108 & ~n_4144;
assign n_4149 = ~n_4145 & ~n_4148;
assign n_4150 =  n_4147 &  n_4149;
assign n_4151 = ~n_4145 & ~n_4150;
assign n_4152 = ~n_4147 & ~n_4149;
assign n_4153 = ~n_4150 & ~n_4152;
assign n_4154 =  n_4132 & ~n_4140;
assign n_4155 = ~n_4141 & ~n_4154;
assign n_4156 = ~n_4142 & ~n_4155;
assign n_4157 =  n_4142 &  n_4155;
assign n_4158 = ~n_4157 & ~n_4108;
assign n_4159 = ~n_4156 & ~n_4158;
assign n_4160 =  n_4153 & ~n_4159;
assign n_4161 = ~n_4153 &  n_4159;
assign n_4162 = ~n_4160 & ~n_4161;
assign n_4163 = ~n_4151 &  n_4162;
assign n_4164 =  n_4080 & ~n_4082;
assign n_4165 = ~n_4095 & ~n_4164;
assign n_4166 = ~n_4162 &  n_4165;
assign n_4167 = ~n_4163 & ~n_4166;
assign n_4168 = ~n_4011 & ~n_4019;
assign n_4169 =  n_4162 & ~n_4165;
assign n_4170 = ~n_4166 & ~n_4169;
assign n_4171 =  n_4151 &  n_4170;
assign n_4172 = ~n_4151 & ~n_4170;
assign n_4173 = ~n_4171 & ~n_4172;
assign n_4174 =  n_4168 & ~n_4173;
assign n_4175 = ~n_4168 &  n_4173;
assign n_4176 = ~n_4174 & ~n_4175;
assign n_4177 = ~n_4167 & ~n_4176;
assign n_4178 =  n_4167 &  n_4176;
assign n_4179 = ~n_4177 & ~n_4178;
assign n_4180 = ~n_4172 & ~n_4167;
assign n_4181 = ~n_4174 & ~n_4180;
assign n_4182 = ~n_4066 & ~n_4075;
assign n_4183 = ~n_4064 &  n_4182;
assign n_4184 =  n_4181 & ~n_4183;
assign n_4185 = ~n_4181 &  n_4183;
assign n_4186 = ~n_4184 & ~n_4185;
assign n_4187 =  n_4179 &  n_4186;
assign n_4188 = ~n_4179 & ~n_4186;
assign n_4189 = ~n_4187 & ~n_4188;
assign n_4190 = ~n_4035 &  n_4189;
assign n_4191 = ~n_4181 & ~n_4177;
assign n_4192 =  n_4183 & ~n_4179;
assign n_4193 = ~n_4191 & ~n_4192;
assign n_4194 = ~n_4193 & ~n_4189;
assign n_4195 = ~n_4190 & ~n_4194;
assign n_4196 =  n_4044 & ~n_4195;
assign n_4197 = ~n_4044 &  n_4195;
assign n_4198 = ~n_4196 & ~n_4197;
assign n_4199 =  n_4035 & ~n_4189;
assign n_4200 = ~n_4190 & ~n_4199;
assign n_4201 = ~n_4193 & ~n_4200;
assign n_4202 = ~n_4193 &  n_4189;
assign n_4203 = ~n_4199 & ~n_4202;
assign n_4204 = ~n_4201 & ~n_4203;
assign n_4205 =  n_4193 &  n_4200;
assign n_4206 = ~n_4201 & ~n_4205;
assign n_4207 =  n_4044 & ~n_4206;
assign n_4208 = ~n_4204 & ~n_4207;
assign n_4209 = ~n_4198 &  n_4208;
assign n_4210 = ~n_4039 & ~n_4209;
assign n_4211 = ~n_4043 & ~n_4210;
assign n_4212 = ~n_4038 & ~n_4211;
assign n_4213 =  n_4042 & ~n_4209;
assign n_4214 =  n_4039 & ~n_4198;
assign n_4215 =  n_4043 &  n_4209;
assign n_4216 = ~n_4214 & ~n_4215;
assign n_4217 = ~n_4213 &  n_4216;
assign n_4218 =  n_4212 & ~n_4217;
assign n_4219 =  n_4038 &  n_4211;
assign n_4220 = ~n_4212 &  n_4217;
assign n_4221 = ~n_4219 &  n_4220;
assign n_4222 = ~n_4214 & ~n_4221;
assign n_4223 = ~n_4218 &  n_4222;
assign n_4224 =  n_4027 & ~n_4223;
assign n_4225 =  n_4043 &  n_4216;
assign n_4226 = ~n_4212 & ~n_4225;
assign n_4227 =  n_4222 &  n_4226;
assign n_4228 = ~n_4224 & ~n_4227;
assign n_4229 = ~n_4047 &  n_4078;
assign n_4230 = ~n_4079 & ~n_4229;
assign n_4231 = ~n_4027 &  n_4223;
assign n_4232 = ~n_4224 & ~n_4231;
assign n_4233 =  n_4226 & ~n_4232;
assign n_4234 = ~n_4226 &  n_4232;
assign n_4235 = ~n_4233 & ~n_4234;
assign n_4236 =  n_4230 & ~n_4235;
assign n_4237 = ~n_4230 &  n_4235;
assign n_4238 = ~n_4236 & ~n_4237;
assign n_4239 =  n_4228 &  n_4238;
assign n_4240 = ~n_4228 & ~n_4238;
assign n_4241 = ~n_4239 & ~n_4240;
assign n_4242 =  n_4001 & ~n_4241;
assign n_4243 = ~n_4228 & ~n_4233;
assign n_4244 = ~n_4243 & ~n_4236;
assign n_4245 = ~n_4240 & ~n_4244;
assign n_4246 = ~n_4242 & ~n_4245;
assign n_4247 = ~n_4001 &  n_4244;
assign n_4248 =  n_4001 & ~n_4244;
assign n_4249 = ~n_4247 & ~n_4248;
assign n_4250 =  n_4241 &  n_4249;
assign n_4251 = ~n_4241 & ~n_4249;
assign n_4252 = ~n_4250 & ~n_4251;
assign n_4253 = ~n_4246 &  n_4252;
assign n_4254 = ~n_4097 & ~n_4099;
assign n_4255 = ~n_4252 &  n_4254;
assign n_4256 = ~n_4253 & ~n_4255;
assign n_4257 =  n_4246 & ~n_4254;
assign n_4258 = ~n_4246 &  n_4254;
assign n_4259 = ~n_4257 & ~n_4258;
assign n_4260 =  n_4252 &  n_4259;
assign n_4261 = ~n_4252 & ~n_4259;
assign n_4262 = ~n_4260 & ~n_4261;
assign n_4263 = ~n_4256 &  n_4262;
assign n_4264 =  n_3900 &  n_3981;
assign n_4265 = ~n_3982 & ~n_4264;
assign n_4266 = ~n_4262 & ~n_4265;
assign n_4267 = ~n_4263 & ~n_4266;
assign n_4268 =  n_4256 &  n_4265;
assign n_4269 = ~n_4256 & ~n_4265;
assign n_4270 = ~n_4268 & ~n_4269;
assign n_4271 =  n_4262 &  n_4270;
assign n_4272 = ~n_4262 & ~n_4270;
assign n_4273 = ~n_4271 & ~n_4272;
assign n_4274 = ~n_4267 &  n_4273;
assign n_4275 =  n_4111 &  n_4124;
assign n_4276 = ~n_4117 & ~n_4275;
assign n_4277 = ~n_4273 &  n_4276;
assign n_4278 = ~n_4274 & ~n_4277;
assign n_4279 =  n_4267 & ~n_4276;
assign n_4280 = ~n_4267 &  n_4276;
assign n_4281 = ~n_4279 & ~n_4280;
assign n_4282 =  n_4273 &  n_4281;
assign n_4283 = ~n_4273 & ~n_4281;
assign n_4284 = ~n_4282 & ~n_4283;
assign n_4285 = ~n_4278 &  n_4284;
assign n_4286 = ~n_3921 &  n_3962;
assign n_4287 = ~n_3963 & ~n_4286;
assign n_4288 =  n_4287 & ~n_4284;
assign n_4289 = ~n_4285 & ~n_4288;
assign n_4290 =  n_4109 & ~n_4127;
assign n_4291 = ~n_4128 & ~n_4290;
assign n_4292 =  n_4134 &  n_4291;
assign n_4293 = ~n_4134 & ~n_4291;
assign n_4294 = ~n_4292 & ~n_4293;
assign n_4295 =  n_4278 & ~n_4287;
assign n_4296 = ~n_4278 &  n_4287;
assign n_4297 = ~n_4295 & ~n_4296;
assign n_4298 =  n_4284 &  n_4297;
assign n_4299 = ~n_4284 & ~n_4297;
assign n_4300 = ~n_4298 & ~n_4299;
assign n_4301 =  n_4294 & ~n_4300;
assign n_4302 = ~n_4294 &  n_4300;
assign n_4303 = ~n_4301 & ~n_4302;
assign n_4304 = ~n_4289 & ~n_4303;
assign n_4305 = ~n_4289 &  n_4300;
assign n_4306 = ~n_4301 & ~n_4305;
assign n_4307 = ~n_4304 & ~n_4306;
assign n_4308 = ~n_3943 &  n_3955;
assign n_4309 =  n_3947 &  n_3954;
assign n_4310 = ~n_3936 & ~n_4309;
assign n_4311 = ~n_4308 &  n_4310;
assign n_4312 = ~n_4311 &  n_4306;
assign n_4313 = ~n_4307 & ~n_4312;
assign n_4314 =  n_4142 &  n_4132;
assign n_4315 = ~n_4141 & ~n_4314;
assign n_4316 =  n_4315 & ~n_4312;
assign n_4317 = ~n_4313 & ~n_4316;
assign n_4318 =  n_4289 &  n_4303;
assign n_4319 = ~n_4304 & ~n_4318;
assign n_4320 = ~n_4319 &  n_4311;
assign n_4321 =  n_4315 & ~n_4307;
assign n_4322 = ~n_4320 &  n_4321;
assign n_4323 = ~n_4317 & ~n_4322;
assign n_4324 = ~n_3738 & ~n_4323;
assign n_4325 =  x_120 &  n_4324;
assign n_4326 = ~x_120 & ~n_4324;
assign n_4327 = ~n_4325 & ~n_4326;
assign n_4328 = ~n_4142 &  n_4140;
assign n_4329 = ~n_4154 & ~n_4328;
assign n_4330 = ~n_4108 & ~n_4329;
assign n_4331 = ~n_4157 & ~n_4330;
assign n_4332 =  n_4151 & ~n_4165;
assign n_4333 = ~n_4163 & ~n_4332;
assign n_4334 = ~n_4184 & ~n_4191;
assign n_4335 =  n_4203 & ~n_4044;
assign n_4336 = ~n_4204 & ~n_4335;
assign n_4337 =  n_4228 & ~n_4230;
assign n_4338 = ~n_4243 & ~n_4337;
assign n_4339 = ~n_4043 &  n_4217;
assign n_4340 = ~n_4212 & ~n_4339;
assign n_4341 = ~n_4214 &  n_4340;
assign n_4342 = ~n_4263 & ~n_4268;
assign n_4343 = ~n_4295 & ~n_4285;
assign n_4344 = ~n_4320 & ~n_4321;
assign n_4345 = ~n_4320 & ~n_4307;
assign n_4346 = ~n_4315 & ~n_4313;
assign n_4347 = ~n_4321 & ~n_4346;
assign n_4348 = ~n_4345 & ~n_4347;
assign n_4349 = ~n_4320 & ~n_4316;
assign n_4350 = ~n_4346 &  n_4349;
assign n_4351 = ~n_4348 & ~n_4350;
assign n_4352 = ~n_4344 &  n_4351;
assign n_4353 = ~n_4147 & ~n_4159;
assign n_4354 = ~n_4145 & ~n_4353;
assign n_4355 = ~n_4351 &  n_4354;
assign n_4356 = ~n_4352 & ~n_4355;
assign n_4357 =  n_4344 & ~n_4354;
assign n_4358 = ~n_4344 &  n_4354;
assign n_4359 = ~n_4357 & ~n_4358;
assign n_4360 =  n_4351 &  n_4359;
assign n_4361 = ~n_4351 & ~n_4359;
assign n_4362 = ~n_4360 & ~n_4361;
assign n_4363 = ~n_4356 &  n_4362;
assign n_4364 =  n_4356 & ~n_4362;
assign n_4365 = ~n_4363 & ~n_4364;
assign n_4366 =  n_4343 & ~n_4365;
assign n_4367 = ~n_4343 &  n_4365;
assign n_4368 = ~n_4366 & ~n_4367;
assign n_4369 = ~n_4168 &  n_4167;
assign n_4370 = ~n_4180 & ~n_4369;
assign n_4371 =  n_4343 & ~n_4362;
assign n_4372 = ~n_4363 & ~n_4371;
assign n_4373 = ~n_4370 &  n_4372;
assign n_4374 =  n_4370 & ~n_4372;
assign n_4375 = ~n_4373 & ~n_4374;
assign n_4376 =  n_4368 & ~n_4375;
assign n_4377 = ~n_4368 &  n_4375;
assign n_4378 = ~n_4376 & ~n_4377;
assign n_4379 =  n_4342 & ~n_4378;
assign n_4380 = ~n_4342 &  n_4378;
assign n_4381 = ~n_4379 & ~n_4380;
assign n_4382 = ~n_4366 & ~n_4370;
assign n_4383 = ~n_4367 & ~n_4382;
assign n_4384 =  n_4381 & ~n_4383;
assign n_4385 = ~n_4381 &  n_4383;
assign n_4386 = ~n_4384 & ~n_4385;
assign n_4387 = ~n_4035 &  n_4193;
assign n_4388 = ~n_4202 & ~n_4387;
assign n_4389 =  n_4378 &  n_4383;
assign n_4390 = ~n_4379 & ~n_4389;
assign n_4391 = ~n_4388 &  n_4390;
assign n_4392 =  n_4388 & ~n_4390;
assign n_4393 = ~n_4391 & ~n_4392;
assign n_4394 =  n_4386 & ~n_4393;
assign n_4395 = ~n_4386 &  n_4393;
assign n_4396 = ~n_4394 & ~n_4395;
assign n_4397 = ~n_4386 &  n_4388;
assign n_4398 = ~n_4385 & ~n_4390;
assign n_4399 = ~n_4397 & ~n_4398;
assign n_4400 = ~n_4245 & ~n_4247;
assign n_4401 =  n_4399 & ~n_4400;
assign n_4402 = ~n_4399 &  n_4400;
assign n_4403 = ~n_4401 & ~n_4402;
assign n_4404 =  n_4396 &  n_4403;
assign n_4405 = ~n_4396 & ~n_4403;
assign n_4406 = ~n_4404 & ~n_4405;
assign n_4407 = ~n_4396 & ~n_4399;
assign n_4408 =  n_4396 &  n_4400;
assign n_4409 = ~n_4407 & ~n_4408;
assign n_4410 = ~n_4198 & ~n_4208;
assign n_4411 =  n_4409 & ~n_4410;
assign n_4412 = ~n_4409 &  n_4410;
assign n_4413 = ~n_4411 & ~n_4412;
assign n_4414 =  n_4406 &  n_4413;
assign n_4415 = ~n_4406 & ~n_4413;
assign n_4416 = ~n_4414 & ~n_4415;
assign n_4417 = ~n_4406 & ~n_4409;
assign n_4418 =  n_4406 &  n_4410;
assign n_4419 = ~n_4417 & ~n_4418;
assign n_4420 = ~n_4027 & ~n_4226;
assign n_4421 = ~n_4227 & ~n_4420;
assign n_4422 = ~n_4419 &  n_4421;
assign n_4423 =  n_4416 &  n_4422;
assign n_4424 =  n_4419 & ~n_4421;
assign n_4425 =  n_4416 &  n_4424;
assign n_4426 = ~n_4416 & ~n_4424;
assign n_4427 = ~n_4425 & ~n_4426;
assign n_4428 = ~n_4416 & ~n_4419;
assign n_4429 =  n_4421 &  n_4428;
assign n_4430 = ~n_4427 & ~n_4429;
assign n_4431 = ~n_4423 & ~n_4430;
assign n_4432 =  n_4214 & ~n_4431;
assign n_4433 =  n_4416 &  n_4419;
assign n_4434 = ~n_4428 & ~n_4433;
assign n_4435 = ~n_4424 & ~n_4434;
assign n_4436 = ~n_4432 & ~n_4435;
assign n_4437 =  n_4039 &  n_4198;
assign n_4438 = ~n_4043 & ~n_4437;
assign n_4439 =  n_4436 &  n_4438;
assign n_4440 = ~n_4214 &  n_4435;
assign n_4441 =  n_4431 &  n_4440;
assign n_4442 = ~n_4430 & ~n_4432;
assign n_4443 = ~n_4441 &  n_4442;
assign n_4444 =  n_4439 &  n_4443;
assign n_4445 =  n_4436 & ~n_4438;
assign n_4446 = ~n_4443 &  n_4445;
assign n_4447 = ~n_4444 & ~n_4446;
assign n_4448 = ~n_4432 &  n_4447;
assign n_4449 = ~n_4341 &  n_4448;
assign n_4450 =  n_4341 & ~n_4447;
assign n_4451 = ~n_4214 & ~n_4450;
assign n_4452 = ~n_4039 & ~n_4198;
assign n_4453 = ~n_4437 & ~n_4452;
assign n_4454 = ~n_4208 &  n_4453;
assign n_4455 =  n_4451 & ~n_4454;
assign n_4456 = ~n_4449 &  n_4455;
assign n_4457 =  n_4214 &  n_4448;
assign n_4458 =  n_4449 &  n_4454;
assign n_4459 = ~n_4457 &  n_4458;
assign n_4460 = ~n_4432 & ~n_4450;
assign n_4461 = ~n_4459 &  n_4460;
assign n_4462 = ~n_4456 &  n_4461;
assign n_4463 =  n_4338 & ~n_4462;
assign n_4464 = ~n_4338 &  n_4462;
assign n_4465 = ~n_4463 & ~n_4464;
assign n_4466 = ~n_4449 &  n_4454;
assign n_4467 =  n_4451 & ~n_4466;
assign n_4468 =  n_4465 &  n_4467;
assign n_4469 = ~n_4465 & ~n_4467;
assign n_4470 = ~n_4468 & ~n_4469;
assign n_4471 =  n_4336 & ~n_4470;
assign n_4472 =  n_4461 & ~n_4467;
assign n_4473 = ~n_4463 & ~n_4472;
assign n_4474 = ~n_4469 & ~n_4473;
assign n_4475 = ~n_4471 & ~n_4474;
assign n_4476 = ~n_4253 & ~n_4257;
assign n_4477 = ~n_4336 &  n_4473;
assign n_4478 =  n_4336 & ~n_4473;
assign n_4479 = ~n_4477 & ~n_4478;
assign n_4480 =  n_4470 &  n_4479;
assign n_4481 = ~n_4470 & ~n_4479;
assign n_4482 = ~n_4480 & ~n_4481;
assign n_4483 = ~n_4476 &  n_4482;
assign n_4484 =  n_4476 & ~n_4482;
assign n_4485 = ~n_4483 & ~n_4484;
assign n_4486 =  n_4475 &  n_4485;
assign n_4487 = ~n_4475 & ~n_4485;
assign n_4488 = ~n_4486 & ~n_4487;
assign n_4489 =  n_4334 & ~n_4488;
assign n_4490 = ~n_4475 &  n_4482;
assign n_4491 = ~n_4484 & ~n_4490;
assign n_4492 = ~n_4487 & ~n_4491;
assign n_4493 = ~n_4489 & ~n_4492;
assign n_4494 = ~n_4274 & ~n_4279;
assign n_4495 = ~n_4475 & ~n_4482;
assign n_4496 = ~n_4483 & ~n_4495;
assign n_4497 =  n_4334 &  n_4496;
assign n_4498 = ~n_4334 & ~n_4496;
assign n_4499 = ~n_4497 & ~n_4498;
assign n_4500 =  n_4494 &  n_4499;
assign n_4501 = ~n_4494 & ~n_4499;
assign n_4502 = ~n_4500 & ~n_4501;
assign n_4503 =  n_4493 & ~n_4502;
assign n_4504 = ~n_4493 &  n_4502;
assign n_4505 = ~n_4503 & ~n_4504;
assign n_4506 =  n_4333 &  n_4505;
assign n_4507 = ~n_4497 & ~n_4500;
assign n_4508 = ~n_4505 & ~n_4507;
assign n_4509 = ~n_4506 & ~n_4508;
assign n_4510 =  n_4289 & ~n_4294;
assign n_4511 = ~n_4305 & ~n_4510;
assign n_4512 = ~n_4333 & ~n_4505;
assign n_4513 = ~n_4506 & ~n_4512;
assign n_4514 =  n_4507 &  n_4513;
assign n_4515 = ~n_4507 & ~n_4513;
assign n_4516 = ~n_4514 & ~n_4515;
assign n_4517 =  n_4511 & ~n_4516;
assign n_4518 = ~n_4511 &  n_4516;
assign n_4519 = ~n_4517 & ~n_4518;
assign n_4520 =  n_4509 &  n_4519;
assign n_4521 = ~n_4509 & ~n_4519;
assign n_4522 = ~n_4520 & ~n_4521;
assign n_4523 =  n_4331 & ~n_4522;
assign n_4524 = ~n_4509 & ~n_4515;
assign n_4525 = ~n_4517 & ~n_4524;
assign n_4526 = ~n_4521 & ~n_4525;
assign n_4527 = ~n_4523 & ~n_4526;
assign n_4528 = ~n_4331 &  n_4525;
assign n_4529 =  n_4331 & ~n_4525;
assign n_4530 = ~n_4528 & ~n_4529;
assign n_4531 =  n_4522 &  n_4530;
assign n_4532 = ~n_4522 & ~n_4530;
assign n_4533 = ~n_4531 & ~n_4532;
assign n_4534 = ~n_4527 &  n_4533;
assign n_4535 =  n_4527 & ~n_4533;
assign n_4536 = ~n_4534 & ~n_4535;
assign n_4537 =  n_4319 & ~n_4311;
assign n_4538 = ~n_4320 & ~n_4537;
assign n_4539 =  n_4306 &  n_4538;
assign n_4540 = ~n_4306 & ~n_4538;
assign n_4541 = ~n_4539 & ~n_4540;
assign n_4542 =  n_4536 & ~n_4541;
assign n_4543 = ~n_4536 &  n_4541;
assign n_4544 = ~n_4542 & ~n_4543;
assign n_4545 = ~n_4128 &  n_4131;
assign n_4546 =  n_4125 &  n_4130;
assign n_4547 = ~n_4135 & ~n_4546;
assign n_4548 = ~n_4545 &  n_4547;
assign n_4549 = ~n_4533 &  n_4541;
assign n_4550 = ~n_4534 & ~n_4549;
assign n_4551 = ~n_4548 &  n_4550;
assign n_4552 =  n_4548 & ~n_4550;
assign n_4553 = ~n_4551 & ~n_4552;
assign n_4554 =  n_4544 & ~n_4553;
assign n_4555 = ~n_4544 &  n_4553;
assign n_4556 = ~n_4554 & ~n_4555;
assign n_4557 = ~n_3738 & ~n_4556;
assign n_4558 =  x_119 &  n_4557;
assign n_4559 = ~x_119 & ~n_4557;
assign n_4560 = ~n_4558 & ~n_4559;
assign n_4561 = ~n_4343 &  n_4356;
assign n_4562 = ~n_4363 & ~n_4561;
assign n_4563 =  x_118 & ~n_4562;
assign n_4564 = ~x_118 &  n_4562;
assign n_4565 = ~n_4563 & ~n_4564;
assign n_4566 =  n_4527 & ~n_4541;
assign n_4567 = ~n_4534 & ~n_4566;
assign n_4568 = ~n_3738 & ~n_4567;
assign n_4569 =  x_117 &  n_4568;
assign n_4570 = ~x_117 & ~n_4568;
assign n_4571 = ~n_4569 & ~n_4570;
assign n_4572 = ~n_4342 & ~n_4383;
assign n_4573 = ~n_4389 & ~n_4572;
assign n_4574 = ~n_3738 & ~n_4573;
assign n_4575 =  x_116 &  n_4574;
assign n_4576 = ~x_116 & ~n_4574;
assign n_4577 = ~n_4575 & ~n_4576;
assign n_4578 =  n_4509 & ~n_4511;
assign n_4579 = ~n_4524 & ~n_4578;
assign n_4580 =  x_115 & ~n_4579;
assign n_4581 = ~x_115 &  n_4579;
assign n_4582 = ~n_4580 & ~n_4581;
assign n_4583 = ~n_4401 & ~n_4407;
assign n_4584 = ~n_3738 & ~n_4583;
assign n_4585 =  x_114 &  n_4584;
assign n_4586 = ~x_114 & ~n_4584;
assign n_4587 = ~n_4585 & ~n_4586;
assign n_4588 =  n_4493 & ~n_4494;
assign n_4589 = ~n_4497 & ~n_4588;
assign n_4590 =  x_113 & ~n_4589;
assign n_4591 = ~x_113 &  n_4589;
assign n_4592 = ~n_4590 & ~n_4591;
assign n_4593 = ~n_4424 & ~n_4429;
assign n_4594 = ~n_3738 & ~n_4593;
assign n_4595 =  x_112 &  n_4594;
assign n_4596 = ~x_112 & ~n_4594;
assign n_4597 = ~n_4595 & ~n_4596;
assign n_4598 =  n_4475 & ~n_4476;
assign n_4599 = ~n_4490 & ~n_4598;
assign n_4600 =  x_111 & ~n_4599;
assign n_4601 = ~x_111 &  n_4599;
assign n_4602 = ~n_4600 & ~n_4601;
assign n_4603 = ~n_4445 & ~n_4457;
assign n_4604 = ~n_3738 & ~n_4603;
assign n_4605 =  x_110 &  n_4604;
assign n_4606 = ~x_110 & ~n_4604;
assign n_4607 = ~n_4605 & ~n_4606;
assign n_4608 = ~n_4338 &  n_4467;
assign n_4609 = ~n_4472 & ~n_4608;
assign n_4610 = ~n_3738 & ~n_4609;
assign n_4611 =  x_109 &  n_4610;
assign n_4612 = ~x_109 & ~n_4610;
assign n_4613 = ~n_4611 & ~n_4612;
assign n_4614 = ~n_4432 & ~n_4439;
assign n_4615 =  n_4447 & ~n_4614;
assign n_4616 = ~n_3738 & ~n_4615;
assign n_4617 =  x_108 &  n_4616;
assign n_4618 = ~x_108 & ~n_4616;
assign n_4619 = ~n_4617 & ~n_4618;
assign n_4620 =  n_4340 & ~n_4457;
assign n_4621 = ~n_3738 & ~n_4620;
assign n_4622 =  x_107 &  n_4621;
assign n_4623 = ~x_107 & ~n_4621;
assign n_4624 = ~n_4622 & ~n_4623;
assign n_4625 = ~n_4432 & ~n_3738;
assign n_4626 =  x_106 &  n_4625;
assign n_4627 = ~x_106 & ~n_4625;
assign n_4628 = ~n_4626 & ~n_4627;
assign n_4629 =  x_105 &  n_4625;
assign n_4630 = ~x_105 & ~n_4625;
assign n_4631 = ~n_4629 & ~n_4630;
assign n_4632 =  x_104 &  n_4625;
assign n_4633 = ~x_104 & ~n_4625;
assign n_4634 = ~n_4632 & ~n_4633;
assign n_4635 =  x_103 &  n_4625;
assign n_4636 = ~x_103 & ~n_4625;
assign n_4637 = ~n_4635 & ~n_4636;
assign n_4638 =  x_102 &  n_4625;
assign n_4639 = ~x_102 & ~n_4625;
assign n_4640 = ~n_4638 & ~n_4639;
assign n_4641 =  x_101 &  n_4625;
assign n_4642 = ~x_101 & ~n_4625;
assign n_4643 = ~n_4641 & ~n_4642;
assign n_4644 =  x_100 &  n_4625;
assign n_4645 = ~x_100 & ~n_4625;
assign n_4646 = ~n_4644 & ~n_4645;
assign n_4647 =  x_99 &  n_4625;
assign n_4648 = ~x_99 & ~n_4625;
assign n_4649 = ~n_4647 & ~n_4648;
assign n_4650 =  x_98 &  n_4625;
assign n_4651 = ~x_98 & ~n_4625;
assign n_4652 = ~n_4650 & ~n_4651;
assign n_4653 =  x_97 &  n_4625;
assign n_4654 = ~x_97 & ~n_4625;
assign n_4655 = ~n_4653 & ~n_4654;
assign n_4656 =  x_96 &  n_4625;
assign n_4657 = ~x_96 & ~n_4625;
assign n_4658 = ~n_4656 & ~n_4657;
assign n_4659 =  x_95 &  n_4625;
assign n_4660 = ~x_95 & ~n_4625;
assign n_4661 = ~n_4659 & ~n_4660;
assign n_4662 =  x_94 &  n_4625;
assign n_4663 = ~x_94 & ~n_4625;
assign n_4664 = ~n_4662 & ~n_4663;
assign n_4665 =  x_93 &  n_4625;
assign n_4666 = ~x_93 & ~n_4625;
assign n_4667 = ~n_4665 & ~n_4666;
assign n_4668 =  x_92 &  n_4625;
assign n_4669 = ~x_92 & ~n_4625;
assign n_4670 = ~n_4668 & ~n_4669;
assign n_4671 =  x_91 &  n_4625;
assign n_4672 = ~x_91 & ~n_4625;
assign n_4673 = ~n_4671 & ~n_4672;
assign n_4674 =  x_90 &  n_4625;
assign n_4675 = ~x_90 & ~n_4625;
assign n_4676 = ~n_4674 & ~n_4675;
assign n_4677 =  x_89 &  n_4625;
assign n_4678 = ~x_89 & ~n_4625;
assign n_4679 = ~n_4677 & ~n_4678;
assign n_4680 =  x_88 &  n_4625;
assign n_4681 = ~x_88 & ~n_4625;
assign n_4682 = ~n_4680 & ~n_4681;
assign n_4683 =  x_87 &  n_4625;
assign n_4684 = ~x_87 & ~n_4625;
assign n_4685 = ~n_4683 & ~n_4684;
assign n_4686 =  x_86 &  n_4625;
assign n_4687 = ~x_86 & ~n_4625;
assign n_4688 = ~n_4686 & ~n_4687;
assign n_4689 =  x_85 &  n_4625;
assign n_4690 = ~x_85 & ~n_4625;
assign n_4691 = ~n_4689 & ~n_4690;
assign n_4692 =  x_84 &  n_4625;
assign n_4693 = ~x_84 & ~n_4625;
assign n_4694 = ~n_4692 & ~n_4693;
assign n_4695 =  x_83 &  n_4625;
assign n_4696 = ~x_83 & ~n_4625;
assign n_4697 = ~n_4695 & ~n_4696;
assign n_4698 =  x_82 &  n_4625;
assign n_4699 = ~x_82 & ~n_4625;
assign n_4700 = ~n_4698 & ~n_4699;
assign n_4701 =  x_81 &  n_4625;
assign n_4702 = ~x_81 & ~n_4625;
assign n_4703 = ~n_4701 & ~n_4702;
assign n_4704 =  x_80 &  n_4625;
assign n_4705 = ~x_80 & ~n_4625;
assign n_4706 = ~n_4704 & ~n_4705;
assign n_4707 =  x_79 &  n_4625;
assign n_4708 = ~x_79 & ~n_4625;
assign n_4709 = ~n_4707 & ~n_4708;
assign n_4710 =  x_78 &  n_4625;
assign n_4711 = ~x_78 & ~n_4625;
assign n_4712 = ~n_4710 & ~n_4711;
assign n_4713 =  x_77 &  n_4625;
assign n_4714 = ~x_77 & ~n_4625;
assign n_4715 = ~n_4713 & ~n_4714;
assign n_4716 =  x_76 &  n_4625;
assign n_4717 = ~x_76 & ~n_4625;
assign n_4718 = ~n_4716 & ~n_4717;
assign n_4719 =  x_75 &  n_4625;
assign n_4720 = ~x_75 & ~n_4625;
assign n_4721 = ~n_4719 & ~n_4720;
assign n_4722 =  x_74 &  n_4625;
assign n_4723 = ~x_74 & ~n_4625;
assign n_4724 = ~n_4722 & ~n_4723;
assign n_4725 =  n_4454 & ~n_4457;
assign n_4726 = ~n_3738 & ~n_4725;
assign n_4727 =  x_73 &  n_4726;
assign n_4728 = ~x_73 & ~n_4726;
assign n_4729 = ~n_4727 & ~n_4728;
assign n_4730 = ~n_4436 &  n_4438;
assign n_4731 = ~n_4443 &  n_4730;
assign n_4732 = ~n_3738 & ~n_4731;
assign n_4733 =  x_72 &  n_4732;
assign n_4734 = ~x_72 & ~n_4732;
assign n_4735 = ~n_4733 & ~n_4734;
assign n_4736 = ~n_4474 & ~n_4477;
assign n_4737 = ~n_3738 & ~n_4736;
assign n_4738 =  x_71 &  n_4737;
assign n_4739 = ~x_71 & ~n_4737;
assign n_4740 = ~n_4738 & ~n_4739;
assign n_4741 = ~n_4423 & ~n_3738;
assign n_4742 =  x_70 &  n_4741;
assign n_4743 = ~x_70 & ~n_4741;
assign n_4744 = ~n_4742 & ~n_4743;
assign n_4745 = ~n_4334 &  n_4491;
assign n_4746 = ~n_4492 & ~n_4745;
assign n_4747 = ~n_3738 & ~n_4746;
assign n_4748 =  x_69 &  n_4747;
assign n_4749 = ~x_69 & ~n_4747;
assign n_4750 = ~n_4748 & ~n_4749;
assign n_4751 = ~n_4411 & ~n_4417;
assign n_4752 = ~n_3738 & ~n_4751;
assign n_4753 =  x_68 &  n_4752;
assign n_4754 = ~x_68 & ~n_4752;
assign n_4755 = ~n_4753 & ~n_4754;
assign n_4756 = ~n_4333 &  n_4507;
assign n_4757 = ~n_4508 & ~n_4756;
assign n_4758 = ~n_3738 & ~n_4757;
assign n_4759 =  x_67 &  n_4758;
assign n_4760 = ~x_67 & ~n_4758;
assign n_4761 = ~n_4759 & ~n_4760;
assign n_4762 = ~n_4391 & ~n_4398;
assign n_4763 = ~n_3738 & ~n_4762;
assign n_4764 =  x_66 &  n_4763;
assign n_4765 = ~x_66 & ~n_4763;
assign n_4766 = ~n_4764 & ~n_4765;
assign n_4767 = ~n_4526 & ~n_4528;
assign n_4768 =  x_65 & ~n_4767;
assign n_4769 = ~x_65 &  n_4767;
assign n_4770 = ~n_4768 & ~n_4769;
assign n_4771 = ~n_4366 & ~n_4373;
assign n_4772 = ~n_3738 & ~n_4771;
assign n_4773 =  x_64 &  n_4772;
assign n_4774 = ~x_64 & ~n_4772;
assign n_4775 = ~n_4773 & ~n_4774;
assign n_4776 = ~n_4543 & ~n_4551;
assign n_4777 =  x_63 & ~n_4776;
assign n_4778 = ~x_63 &  n_4776;
assign n_4779 = ~n_4777 & ~n_4778;
assign n_4780 = ~n_4543 & ~n_4548;
assign n_4781 = ~n_4542 & ~n_4780;
assign n_4782 =  x_61 &  n_4781;
assign n_4783 = ~x_61 & ~n_4781;
assign n_4784 = ~n_4782 & ~n_4783;
assign n_4785 = ~n_4352 & ~n_4357;
assign n_4786 = ~n_4785 & ~n_3738;
assign n_4787 =  x_62 &  n_4786;
assign n_4788 = ~x_62 & ~n_4786;
assign n_4789 = ~n_4787 & ~n_4788;
assign n_4790 = ~n_4784 & ~n_4789;
assign n_4791 = ~n_4779 &  n_4790;
assign n_4792 = ~n_4775 &  n_4791;
assign n_4793 = ~n_4770 &  n_4792;
assign n_4794 = ~n_4766 &  n_4793;
assign n_4795 = ~n_4761 &  n_4794;
assign n_4796 = ~n_4755 &  n_4795;
assign n_4797 = ~n_4750 &  n_4796;
assign n_4798 = ~n_4744 &  n_4797;
assign n_4799 = ~n_4740 &  n_4798;
assign n_4800 = ~n_4735 &  n_4799;
assign n_4801 = ~n_4729 &  n_4800;
assign n_4802 = ~n_4724 &  n_4801;
assign n_4803 = ~n_4721 &  n_4802;
assign n_4804 = ~n_4718 &  n_4803;
assign n_4805 = ~n_4715 &  n_4804;
assign n_4806 = ~n_4712 &  n_4805;
assign n_4807 = ~n_4709 &  n_4806;
assign n_4808 = ~n_4706 &  n_4807;
assign n_4809 = ~n_4703 &  n_4808;
assign n_4810 = ~n_4700 &  n_4809;
assign n_4811 = ~n_4697 &  n_4810;
assign n_4812 = ~n_4694 &  n_4811;
assign n_4813 = ~n_4691 &  n_4812;
assign n_4814 = ~n_4688 &  n_4813;
assign n_4815 = ~n_4685 &  n_4814;
assign n_4816 = ~n_4682 &  n_4815;
assign n_4817 = ~n_4679 &  n_4816;
assign n_4818 = ~n_4676 &  n_4817;
assign n_4819 = ~n_4673 &  n_4818;
assign n_4820 = ~n_4670 &  n_4819;
assign n_4821 = ~n_4667 &  n_4820;
assign n_4822 = ~n_4664 &  n_4821;
assign n_4823 = ~n_4661 &  n_4822;
assign n_4824 = ~n_4658 &  n_4823;
assign n_4825 = ~n_4655 &  n_4824;
assign n_4826 = ~n_4652 &  n_4825;
assign n_4827 = ~n_4649 &  n_4826;
assign n_4828 = ~n_4646 &  n_4827;
assign n_4829 = ~n_4643 &  n_4828;
assign n_4830 = ~n_4640 &  n_4829;
assign n_4831 = ~n_4637 &  n_4830;
assign n_4832 = ~n_4634 &  n_4831;
assign n_4833 = ~n_4631 &  n_4832;
assign n_4834 = ~n_4628 &  n_4833;
assign n_4835 = ~n_4624 &  n_4834;
assign n_4836 = ~n_4619 &  n_4835;
assign n_4837 = ~n_4613 &  n_4836;
assign n_4838 = ~n_4607 &  n_4837;
assign n_4839 = ~n_4602 &  n_4838;
assign n_4840 = ~n_4597 &  n_4839;
assign n_4841 = ~n_4592 &  n_4840;
assign n_4842 = ~n_4587 &  n_4841;
assign n_4843 = ~n_4582 &  n_4842;
assign n_4844 = ~n_4577 &  n_4843;
assign n_4845 = ~n_4571 &  n_4844;
assign n_4846 = ~n_4565 &  n_4845;
assign n_4847 = ~n_4560 &  n_4846;
assign n_4848 = ~n_4327 &  n_4847;
assign o_1 = ~n_4848;
endmodule

