// Generated using findDep.cpp 
module trueque_query42_1344n (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_55, v_56, v_57, v_58, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_20, v_44, v_54, v_59, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_266, v_267, v_268, v_269, v_270, v_271, v_273, v_274, v_275, v_276, v_277, v_278, v_280, v_281, v_282, v_284, v_285, v_286, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_296, v_297, v_298, v_300, v_301, v_302, v_304, v_305, v_306, v_308, v_309, v_310, v_312, v_313, v_314, v_316, v_317, v_318, v_320, v_321, v_322, v_324, v_325, v_326, v_328, v_329, v_330, v_331, v_332, v_333, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_55;
input v_56;
input v_57;
input v_58;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_20;
input v_44;
input v_54;
input v_59;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_280;
input v_281;
input v_282;
input v_284;
input v_285;
input v_286;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_296;
input v_297;
input v_298;
input v_300;
input v_301;
input v_302;
input v_304;
input v_305;
input v_306;
input v_308;
input v_309;
input v_310;
input v_312;
input v_313;
input v_314;
input v_316;
input v_317;
input v_318;
input v_320;
input v_321;
input v_322;
input v_324;
input v_325;
input v_326;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
output o_1;
wire v_241;
wire v_265;
wire v_272;
wire v_279;
wire v_283;
wire v_287;
wire v_295;
wire v_299;
wire v_303;
wire v_307;
wire v_311;
wire v_315;
wire v_319;
wire v_323;
wire v_327;
wire v_334;
wire v_335;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
assign v_335 = 0;
assign v_334 = 0;
assign v_327 = 0;
assign v_323 = 0;
assign v_319 = 0;
assign v_315 = 0;
assign v_311 = 0;
assign v_307 = 0;
assign v_303 = 0;
assign v_299 = 0;
assign v_295 = 0;
assign v_287 = 0;
assign v_283 = 0;
assign v_279 = 0;
assign v_272 = 0;
assign v_265 = 0;
assign v_241 = 0;
assign x_1 = v_5 | v_4 | v_6 | v_3 | v_2 | v_1 | ~v_240 | ~v_239 | ~v_333;
assign x_2 = v_333 | ~v_332;
assign x_3 = v_333 | ~v_293;
assign x_4 = v_333 | ~v_263;
assign x_5 = v_333 | ~v_237;
assign x_6 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_331 | v_332;
assign x_7 = v_331 | ~v_328;
assign x_8 = v_331 | ~v_329;
assign x_9 = v_331 | ~v_330;
assign x_10 = v_32 | v_38 | v_33 | v_35 | v_37 | v_36 | v_34 | ~v_149 | ~v_148 | ~v_99 | ~v_98 | v_330;
assign x_11 = v_25 | v_24 | v_23 | v_28 | v_29 | v_27 | v_26 | ~v_146 | ~v_145 | ~v_94 | ~v_93 | v_329;
assign x_12 = v_13 | v_19 | v_18 | v_17 | v_16 | v_15 | v_14 | ~v_143 | ~v_142 | ~v_89 | ~v_88 | v_328;
assign x_13 = v_5 | v_4 | v_3 | v_2 | v_1 | v_66 | ~v_240 | ~v_239 | ~v_326;
assign x_14 = v_326 | ~v_324;
assign x_15 = v_326 | ~v_325;
assign x_16 = v_326 | ~v_266;
assign x_17 = v_326 | ~v_210;
assign x_18 = v_326 | ~v_211;
assign x_19 = v_326 | ~v_267;
assign x_20 = v_326 | ~v_212;
assign x_21 = ~v_222 | ~v_218 | v_325;
assign x_22 = ~v_258 | ~v_254 | v_324;
assign x_23 = v_4 | v_6 | v_3 | v_2 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_322;
assign x_24 = v_322 | ~v_320;
assign x_25 = v_322 | ~v_321;
assign x_26 = v_322 | ~v_186;
assign x_27 = v_322 | ~v_195;
assign x_28 = v_322 | ~v_196;
assign x_29 = v_322 | ~v_197;
assign x_30 = v_322 | ~v_198;
assign x_31 = ~v_218 | ~v_250 | v_321;
assign x_32 = ~v_236 | ~v_258 | v_320;
assign x_33 = v_5 | v_4 | v_6 | v_3 | v_2 | v_65 | ~v_240 | ~v_239 | ~v_318;
assign x_34 = v_318 | ~v_316;
assign x_35 = v_318 | ~v_317;
assign x_36 = v_318 | ~v_227;
assign x_37 = v_318 | ~v_232;
assign x_38 = v_318 | ~v_233;
assign x_39 = v_318 | ~v_234;
assign x_40 = v_318 | ~v_235;
assign x_41 = ~v_262 | ~v_199 | v_317;
assign x_42 = ~v_275 | ~v_218 | v_316;
assign x_43 = v_5 | v_4 | v_3 | v_2 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_314;
assign x_44 = v_314 | ~v_312;
assign x_45 = v_314 | ~v_313;
assign x_46 = v_314 | ~v_209;
assign x_47 = v_314 | ~v_214;
assign x_48 = v_314 | ~v_215;
assign x_49 = v_314 | ~v_216;
assign x_50 = v_314 | ~v_217;
assign x_51 = ~v_254 | ~v_199 | v_313;
assign x_52 = ~v_236 | ~v_268 | v_312;
assign x_53 = v_4 | v_6 | v_3 | v_2 | v_1 | v_66 | ~v_240 | ~v_239 | ~v_310;
assign x_54 = v_310 | ~v_308;
assign x_55 = v_310 | ~v_309;
assign x_56 = v_310 | ~v_256;
assign x_57 = v_310 | ~v_187;
assign x_58 = v_310 | ~v_188;
assign x_59 = v_310 | ~v_257;
assign x_60 = v_310 | ~v_189;
assign x_61 = ~v_222 | ~v_199 | v_309;
assign x_62 = ~v_268 | ~v_250 | v_308;
assign x_63 = v_5 | v_6 | v_3 | v_2 | v_1 | v_66 | ~v_240 | ~v_239 | ~v_306;
assign x_64 = v_306 | ~v_304;
assign x_65 = v_306 | ~v_305;
assign x_66 = v_306 | ~v_114;
assign x_67 = v_306 | ~v_135;
assign x_68 = v_306 | ~v_220;
assign x_69 = v_306 | ~v_221;
assign x_70 = v_306 | ~v_140;
assign x_71 = ~v_258 | ~v_173 | v_305;
assign x_72 = ~v_268 | ~v_204 | v_304;
assign x_73 = v_5 | v_6 | v_2 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_302;
assign x_74 = v_302 | ~v_300;
assign x_75 = v_302 | ~v_301;
assign x_76 = v_302 | ~v_201;
assign x_77 = v_302 | ~v_203;
assign x_78 = v_302 | ~v_157;
assign x_79 = v_302 | ~v_162;
assign x_80 = v_302 | ~v_163;
assign x_81 = ~v_250 | ~v_173 | v_301;
assign x_82 = ~v_222 | ~v_275 | v_300;
assign x_83 = v_5 | v_4 | v_6 | v_2 | v_1 | v_65 | ~v_240 | ~v_239 | ~v_298;
assign x_84 = v_298 | ~v_296;
assign x_85 = v_298 | ~v_297;
assign x_86 = v_298 | ~v_273;
assign x_87 = v_298 | ~v_274;
assign x_88 = v_298 | ~v_223;
assign x_89 = v_298 | ~v_224;
assign x_90 = v_298 | ~v_225;
assign x_91 = ~v_236 | ~v_204 | v_297;
assign x_92 = ~v_262 | ~v_250 | v_296;
assign x_93 = v_5 | v_4 | v_2 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_294;
assign x_94 = v_294 | ~v_292;
assign x_95 = v_294 | ~v_255;
assign x_96 = v_294 | ~v_219;
assign x_97 = v_294 | ~v_293;
assign x_98 = ~v_275 | ~v_268 | v_293;
assign x_99 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_291 | v_292;
assign x_100 = v_291 | ~v_288;
assign x_101 = v_291 | ~v_289;
assign x_102 = v_291 | ~v_290;
assign x_103 = v_32 | v_38 | v_35 | v_37 | v_36 | v_53 | v_49 | ~v_132 | ~v_131 | ~v_122 | ~v_121 | v_290;
assign x_104 = v_23 | v_28 | v_29 | v_27 | v_26 | v_52 | v_46 | ~v_129 | ~v_128 | ~v_119 | ~v_118 | v_289;
assign x_105 = v_13 | v_19 | v_18 | v_17 | v_16 | v_51 | v_42 | ~v_126 | ~v_125 | ~v_116 | ~v_115 | v_288;
assign x_106 = v_4 | v_6 | v_2 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_286;
assign x_107 = v_286 | ~v_284;
assign x_108 = v_286 | ~v_285;
assign x_109 = v_286 | ~v_247;
assign x_110 = v_286 | ~v_249;
assign x_111 = v_286 | ~v_178;
assign x_112 = v_286 | ~v_179;
assign x_113 = v_286 | ~v_180;
assign x_114 = ~v_199 | ~v_204 | v_285;
assign x_115 = ~v_258 | ~v_275 | v_284;
assign x_116 = v_5 | v_6 | v_3 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_282;
assign x_117 = v_282 | ~v_280;
assign x_118 = v_282 | ~v_281;
assign x_119 = v_282 | ~v_152;
assign x_120 = v_282 | ~v_169;
assign x_121 = v_282 | ~v_170;
assign x_122 = v_282 | ~v_171;
assign x_123 = v_282 | ~v_172;
assign x_124 = ~v_254 | ~v_204 | v_281;
assign x_125 = ~v_222 | ~v_262 | v_280;
assign x_126 = v_5 | v_4 | v_6 | v_3 | v_1 | v_65 | ~v_240 | ~v_239 | ~v_278;
assign x_127 = v_278 | ~v_276;
assign x_128 = v_278 | ~v_277;
assign x_129 = v_278 | ~v_259;
assign x_130 = v_278 | ~v_261;
assign x_131 = v_278 | ~v_228;
assign x_132 = v_278 | ~v_229;
assign x_133 = v_278 | ~v_230;
assign x_134 = ~v_236 | ~v_173 | v_277;
assign x_135 = ~v_275 | ~v_254 | v_276;
assign x_136 = v_275 | ~v_273;
assign x_137 = v_275 | ~v_274;
assign x_138 = v_275 | ~v_223;
assign x_139 = v_275 | ~v_224;
assign x_140 = v_275 | ~v_225;
assign x_141 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_260 | ~v_134 | v_274;
assign x_142 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_231 | ~v_156 | v_273;
assign x_143 = v_5 | v_4 | v_3 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_271;
assign x_144 = v_271 | ~v_269;
assign x_145 = v_271 | ~v_270;
assign x_146 = v_271 | ~v_252;
assign x_147 = v_271 | ~v_253;
assign x_148 = v_271 | ~v_205;
assign x_149 = v_271 | ~v_206;
assign x_150 = v_271 | ~v_207;
assign x_151 = ~v_218 | ~v_173 | v_270;
assign x_152 = ~v_262 | ~v_268 | v_269;
assign x_153 = v_268 | ~v_266;
assign x_154 = v_268 | ~v_210;
assign x_155 = v_268 | ~v_211;
assign x_156 = v_268 | ~v_267;
assign x_157 = v_268 | ~v_212;
assign x_158 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_139 | ~v_251 | v_267;
assign x_159 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_103 | ~v_208 | v_266;
assign x_160 = v_4 | v_6 | v_3 | v_1 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_264;
assign x_161 = v_264 | ~v_246;
assign x_162 = v_264 | ~v_200;
assign x_163 = v_264 | ~v_255;
assign x_164 = v_264 | ~v_263;
assign x_165 = ~v_262 | ~v_258 | v_263;
assign x_166 = v_262 | ~v_259;
assign x_167 = v_262 | ~v_261;
assign x_168 = v_262 | ~v_228;
assign x_169 = v_262 | ~v_229;
assign x_170 = v_262 | ~v_230;
assign x_171 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_260 | ~v_113 | v_261;
assign x_172 = v_260 | ~v_233;
assign x_173 = v_260 | ~v_234;
assign x_174 = v_260 | ~v_235;
assign x_175 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_168 | ~v_226 | v_259;
assign x_176 = v_258 | ~v_256;
assign x_177 = v_258 | ~v_187;
assign x_178 = v_258 | ~v_188;
assign x_179 = v_258 | ~v_257;
assign x_180 = v_258 | ~v_189;
assign x_181 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_139 | ~v_248 | v_257;
assign x_182 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_124 | ~v_181 | v_256;
assign x_183 = ~v_254 | ~v_250 | v_255;
assign x_184 = v_254 | ~v_252;
assign x_185 = v_254 | ~v_253;
assign x_186 = v_254 | ~v_205;
assign x_187 = v_254 | ~v_206;
assign x_188 = v_254 | ~v_207;
assign x_189 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | ~v_213 | v_253;
assign x_190 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_113 | ~v_251 | v_252;
assign x_191 = v_251 | ~v_215;
assign x_192 = v_251 | ~v_216;
assign x_193 = v_251 | ~v_217;
assign x_194 = v_250 | ~v_247;
assign x_195 = v_250 | ~v_249;
assign x_196 = v_250 | ~v_178;
assign x_197 = v_250 | ~v_179;
assign x_198 = v_250 | ~v_180;
assign x_199 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_134 | ~v_248 | v_249;
assign x_200 = v_248 | ~v_196;
assign x_201 = v_248 | ~v_197;
assign x_202 = v_248 | ~v_198;
assign x_203 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_190 | v_247;
assign x_204 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_245 | v_246;
assign x_205 = v_245 | ~v_242;
assign x_206 = v_245 | ~v_243;
assign x_207 = v_245 | ~v_244;
assign x_208 = v_32 | v_38 | v_35 | v_37 | v_36 | v_53 | v_49 | ~v_101 | ~v_100 | ~v_111 | ~v_110 | v_244;
assign x_209 = v_23 | v_28 | v_29 | v_27 | v_26 | v_52 | v_46 | ~v_96 | ~v_95 | ~v_108 | ~v_107 | v_243;
assign x_210 = v_13 | v_19 | v_18 | v_17 | v_16 | v_51 | v_42 | ~v_91 | ~v_90 | ~v_105 | ~v_104 | v_242;
assign x_211 = v_5 | v_6 | v_3 | v_2 | v_66 | v_65 | ~v_240 | ~v_239 | ~v_238;
assign x_212 = v_240 | ~v_65;
assign x_213 = v_240 | ~v_3;
assign x_214 = v_240 | ~v_2;
assign x_215 = v_240 | ~v_1;
assign x_216 = v_239 | ~v_66;
assign x_217 = v_239 | ~v_6;
assign x_218 = v_239 | ~v_5;
assign x_219 = v_239 | ~v_4;
assign x_220 = v_238 | ~v_87;
assign x_221 = v_238 | ~v_200;
assign x_222 = v_238 | ~v_219;
assign x_223 = v_238 | ~v_237;
assign x_224 = ~v_236 | ~v_222 | v_237;
assign x_225 = v_236 | ~v_227;
assign x_226 = v_236 | ~v_232;
assign x_227 = v_236 | ~v_233;
assign x_228 = v_236 | ~v_234;
assign x_229 = v_236 | ~v_235;
assign x_230 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | v_235;
assign x_231 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_151 | v_234;
assign x_232 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_185 | v_233;
assign x_233 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_231 | v_232;
assign x_234 = v_231 | ~v_228;
assign x_235 = v_231 | ~v_229;
assign x_236 = v_231 | ~v_230;
assign x_237 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | v_230;
assign x_238 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_113 | v_229;
assign x_239 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_168 | v_228;
assign x_240 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | ~v_226 | v_227;
assign x_241 = v_226 | ~v_223;
assign x_242 = v_226 | ~v_224;
assign x_243 = v_226 | ~v_225;
assign x_244 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | v_225;
assign x_245 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | ~v_156 | v_224;
assign x_246 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_134 | v_223;
assign x_247 = v_222 | ~v_114;
assign x_248 = v_222 | ~v_135;
assign x_249 = v_222 | ~v_220;
assign x_250 = v_222 | ~v_221;
assign x_251 = v_222 | ~v_140;
assign x_252 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_164 | ~v_124 | v_221;
assign x_253 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_202 | ~v_103 | v_220;
assign x_254 = ~v_218 | ~v_204 | v_219;
assign x_255 = v_218 | ~v_209;
assign x_256 = v_218 | ~v_214;
assign x_257 = v_218 | ~v_215;
assign x_258 = v_218 | ~v_216;
assign x_259 = v_218 | ~v_217;
assign x_260 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | v_217;
assign x_261 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_124 | v_216;
assign x_262 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_168 | v_215;
assign x_263 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_213 | v_214;
assign x_264 = v_213 | ~v_210;
assign x_265 = v_213 | ~v_211;
assign x_266 = v_213 | ~v_212;
assign x_267 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_124 | v_212;
assign x_268 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | ~v_139 | v_211;
assign x_269 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_168 | ~v_103 | v_210;
assign x_270 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_208 | v_209;
assign x_271 = v_208 | ~v_205;
assign x_272 = v_208 | ~v_206;
assign x_273 = v_208 | ~v_207;
assign x_274 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_168 | v_207;
assign x_275 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | ~v_124 | v_206;
assign x_276 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | ~v_113 | v_205;
assign x_277 = v_204 | ~v_201;
assign x_278 = v_204 | ~v_203;
assign x_279 = v_204 | ~v_157;
assign x_280 = v_204 | ~v_162;
assign x_281 = v_204 | ~v_163;
assign x_282 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_156 | ~v_202 | v_203;
assign x_283 = v_202 | ~v_170;
assign x_284 = v_202 | ~v_171;
assign x_285 = v_202 | ~v_172;
assign x_286 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_141 | v_201;
assign x_287 = ~v_199 | ~v_173 | v_200;
assign x_288 = v_199 | ~v_186;
assign x_289 = v_199 | ~v_195;
assign x_290 = v_199 | ~v_196;
assign x_291 = v_199 | ~v_197;
assign x_292 = v_199 | ~v_198;
assign x_293 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | v_198;
assign x_294 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_103 | v_197;
assign x_295 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | ~v_156 | v_196;
assign x_296 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_194 | ~v_190 | v_195;
assign x_297 = v_194 | ~v_191;
assign x_298 = v_194 | ~v_192;
assign x_299 = v_194 | ~v_193;
assign x_300 = v_38 | v_37 | v_36 | v_34 | v_53 | v_48 | v_64 | ~v_80 | ~v_79 | ~v_149 | ~v_148 | v_193;
assign x_301 = v_25 | v_28 | v_29 | v_27 | v_52 | v_45 | v_63 | ~v_75 | ~v_74 | ~v_146 | ~v_145 | v_192;
assign x_302 = v_19 | v_18 | v_17 | v_15 | v_51 | v_62 | v_41 | ~v_68 | ~v_67 | ~v_143 | ~v_142 | v_191;
assign x_303 = v_190 | ~v_187;
assign x_304 = v_190 | ~v_188;
assign x_305 = v_190 | ~v_189;
assign x_306 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_103 | v_189;
assign x_307 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_139 | v_188;
assign x_308 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_156 | ~v_124 | v_187;
assign x_309 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_185 | ~v_181 | v_186;
assign x_310 = v_185 | ~v_182;
assign x_311 = v_185 | ~v_183;
assign x_312 = v_185 | ~v_184;
assign x_313 = v_38 | v_37 | v_36 | v_53 | v_49 | v_48 | v_64 | ~v_80 | ~v_79 | ~v_122 | ~v_121 | v_184;
assign x_314 = v_28 | v_29 | v_27 | v_52 | v_46 | v_45 | v_63 | ~v_75 | ~v_74 | ~v_119 | ~v_118 | v_183;
assign x_315 = v_19 | v_18 | v_17 | v_51 | v_62 | v_42 | v_41 | ~v_68 | ~v_67 | ~v_116 | ~v_115 | v_182;
assign x_316 = v_181 | ~v_178;
assign x_317 = v_181 | ~v_179;
assign x_318 = v_181 | ~v_180;
assign x_319 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_156 | v_180;
assign x_320 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_103 | v_179;
assign x_321 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_177 | ~v_134 | v_178;
assign x_322 = v_177 | ~v_174;
assign x_323 = v_177 | ~v_175;
assign x_324 = v_177 | ~v_176;
assign x_325 = v_37 | v_36 | v_53 | v_49 | v_48 | v_64 | v_57 | ~v_80 | ~v_79 | ~v_101 | ~v_100 | v_176;
assign x_326 = v_28 | v_27 | v_56 | v_52 | v_46 | v_45 | v_63 | ~v_75 | ~v_74 | ~v_96 | ~v_95 | v_175;
assign x_327 = v_18 | v_17 | v_55 | v_51 | v_62 | v_42 | v_41 | ~v_91 | ~v_90 | ~v_68 | ~v_67 | v_174;
assign x_328 = v_173 | ~v_152;
assign x_329 = v_173 | ~v_169;
assign x_330 = v_173 | ~v_170;
assign x_331 = v_173 | ~v_171;
assign x_332 = v_173 | ~v_172;
assign x_333 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_113 | v_172;
assign x_334 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | ~v_139 | v_171;
assign x_335 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_168 | ~v_134 | v_170;
assign x_336 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_168 | ~v_164 | v_169;
assign x_337 = v_168 | ~v_165;
assign x_338 = v_168 | ~v_166;
assign x_339 = v_168 | ~v_167;
assign x_340 = v_35 | v_37 | v_36 | v_53 | v_49 | v_48 | v_57 | ~v_111 | ~v_110 | ~v_122 | ~v_121 | v_167;
assign x_341 = v_28 | v_27 | v_26 | v_56 | v_52 | v_46 | v_45 | ~v_108 | ~v_107 | ~v_119 | ~v_118 | v_166;
assign x_342 = v_18 | v_17 | v_16 | v_55 | v_51 | v_42 | v_41 | ~v_105 | ~v_104 | ~v_116 | ~v_115 | v_165;
assign x_343 = v_164 | ~v_157;
assign x_344 = v_164 | ~v_162;
assign x_345 = v_164 | ~v_163;
assign x_346 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_134 | v_163;
assign x_347 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_161 | ~v_139 | v_162;
assign x_348 = v_161 | ~v_158;
assign x_349 = v_161 | ~v_159;
assign x_350 = v_161 | ~v_160;
assign x_351 = v_35 | v_37 | v_36 | v_34 | v_53 | v_48 | v_57 | ~v_149 | ~v_148 | ~v_132 | ~v_131 | v_160;
assign x_352 = v_25 | v_28 | v_27 | v_26 | v_56 | v_52 | v_45 | ~v_146 | ~v_145 | ~v_129 | ~v_128 | v_159;
assign x_353 = v_18 | v_17 | v_16 | v_15 | v_55 | v_51 | v_41 | ~v_143 | ~v_142 | ~v_126 | ~v_125 | v_158;
assign x_354 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_113 | ~v_156 | v_157;
assign x_355 = v_156 | ~v_153;
assign x_356 = v_156 | ~v_154;
assign x_357 = v_156 | ~v_155;
assign x_358 = v_38 | v_35 | v_36 | v_53 | v_50 | v_49 | v_48 | ~v_101 | ~v_100 | ~v_132 | ~v_131 | v_155;
assign x_359 = v_29 | v_27 | v_26 | v_52 | v_46 | v_45 | v_47 | ~v_96 | ~v_95 | ~v_129 | ~v_128 | v_154;
assign x_360 = v_19 | v_17 | v_16 | v_51 | v_43 | v_42 | v_41 | ~v_91 | ~v_90 | ~v_126 | ~v_125 | v_153;
assign x_361 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_151 | ~v_141 | v_152;
assign x_362 = v_151 | ~v_144;
assign x_363 = v_151 | ~v_147;
assign x_364 = v_151 | ~v_150;
assign x_365 = v_38 | v_35 | v_37 | v_36 | v_34 | v_53 | v_48 | ~v_149 | ~v_148 | ~v_111 | ~v_110 | v_150;
assign x_366 = v_149 | v_40;
assign x_367 = v_149 | v_20;
assign x_368 = v_148 | v_39;
assign x_369 = v_148 | ~v_20;
assign x_370 = v_25 | v_28 | v_29 | v_27 | v_26 | v_52 | v_45 | ~v_146 | ~v_145 | ~v_108 | ~v_107 | v_147;
assign x_371 = v_146 | v_31;
assign x_372 = v_146 | v_20;
assign x_373 = v_145 | v_30;
assign x_374 = v_145 | ~v_20;
assign x_375 = v_19 | v_18 | v_17 | v_16 | v_15 | v_51 | v_41 | ~v_143 | ~v_142 | ~v_105 | ~v_104 | v_144;
assign x_376 = v_143 | v_20;
assign x_377 = v_143 | v_22;
assign x_378 = v_142 | v_21;
assign x_379 = v_142 | ~v_20;
assign x_380 = v_141 | ~v_114;
assign x_381 = v_141 | ~v_135;
assign x_382 = v_141 | ~v_140;
assign x_383 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_139 | v_140;
assign x_384 = v_139 | ~v_136;
assign x_385 = v_139 | ~v_137;
assign x_386 = v_139 | ~v_138;
assign x_387 = v_38 | v_33 | v_35 | v_37 | v_61 | v_49 | v_48 | ~v_78 | ~v_77 | ~v_99 | ~v_98 | v_138;
assign x_388 = v_24 | v_28 | v_29 | v_26 | v_46 | v_45 | v_60 | ~v_73 | ~v_72 | ~v_94 | ~v_93 | v_137;
assign x_389 = v_19 | v_18 | v_16 | v_14 | v_58 | v_42 | v_41 | ~v_70 | ~v_69 | ~v_89 | ~v_88 | v_136;
assign x_390 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_134 | ~v_124 | v_135;
assign x_391 = v_134 | ~v_127;
assign x_392 = v_134 | ~v_130;
assign x_393 = v_134 | ~v_133;
assign x_394 = v_38 | v_35 | v_37 | v_53 | v_61 | v_49 | v_48 | ~v_132 | ~v_131 | ~v_78 | ~v_77 | v_133;
assign x_395 = v_132 | v_44;
assign x_396 = v_132 | v_12;
assign x_397 = v_131 | ~v_44;
assign x_398 = v_131 | v_9;
assign x_399 = v_28 | v_29 | v_26 | v_52 | v_46 | v_45 | v_60 | ~v_129 | ~v_128 | ~v_73 | ~v_72 | v_130;
assign x_400 = v_129 | v_44;
assign x_401 = v_129 | v_10;
assign x_402 = v_128 | ~v_44;
assign x_403 = v_128 | v_8;
assign x_404 = v_19 | v_18 | v_16 | v_51 | v_58 | v_42 | v_41 | ~v_70 | ~v_69 | ~v_126 | ~v_125 | v_127;
assign x_405 = v_126 | v_44;
assign x_406 = v_126 | v_11;
assign x_407 = v_125 | ~v_44;
assign x_408 = v_125 | v_7;
assign x_409 = v_124 | ~v_117;
assign x_410 = v_124 | ~v_120;
assign x_411 = v_124 | ~v_123;
assign x_412 = v_38 | v_33 | v_35 | v_36 | v_50 | v_49 | v_48 | ~v_122 | ~v_121 | ~v_99 | ~v_98 | v_123;
assign x_413 = v_122 | v_44;
assign x_414 = v_122 | v_40;
assign x_415 = v_121 | ~v_44;
assign x_416 = v_121 | v_39;
assign x_417 = v_24 | v_29 | v_27 | v_26 | v_46 | v_45 | v_47 | ~v_119 | ~v_118 | ~v_94 | ~v_93 | v_120;
assign x_418 = v_119 | v_44;
assign x_419 = v_119 | v_31;
assign x_420 = v_118 | ~v_44;
assign x_421 = v_118 | v_30;
assign x_422 = v_19 | v_17 | v_16 | v_14 | v_43 | v_42 | v_41 | ~v_116 | ~v_115 | ~v_89 | ~v_88 | v_117;
assign x_423 = v_116 | v_44;
assign x_424 = v_116 | v_22;
assign x_425 = v_115 | ~v_44;
assign x_426 = v_115 | v_21;
assign x_427 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_113 | ~v_103 | v_114;
assign x_428 = v_113 | ~v_106;
assign x_429 = v_113 | ~v_109;
assign x_430 = v_113 | ~v_112;
assign x_431 = v_38 | v_35 | v_53 | v_61 | v_50 | v_49 | v_48 | ~v_111 | ~v_110 | ~v_78 | ~v_77 | v_112;
assign x_432 = v_111 | v_54;
assign x_433 = v_111 | v_12;
assign x_434 = v_110 | ~v_54;
assign x_435 = v_110 | v_9;
assign x_436 = v_29 | v_26 | v_52 | v_46 | v_45 | v_60 | v_47 | ~v_108 | ~v_107 | ~v_73 | ~v_72 | v_109;
assign x_437 = v_108 | v_54;
assign x_438 = v_108 | v_10;
assign x_439 = v_107 | ~v_54;
assign x_440 = v_107 | v_8;
assign x_441 = v_19 | v_16 | v_51 | v_43 | v_58 | v_42 | v_41 | ~v_70 | ~v_69 | ~v_105 | ~v_104 | v_106;
assign x_442 = v_105 | v_54;
assign x_443 = v_105 | v_11;
assign x_444 = v_104 | ~v_54;
assign x_445 = v_104 | v_7;
assign x_446 = v_103 | ~v_92;
assign x_447 = v_103 | ~v_97;
assign x_448 = v_103 | ~v_102;
assign x_449 = v_38 | v_33 | v_35 | v_37 | v_36 | v_49 | v_48 | ~v_101 | ~v_100 | ~v_99 | ~v_98 | v_102;
assign x_450 = v_101 | v_40;
assign x_451 = v_101 | v_54;
assign x_452 = v_100 | ~v_54;
assign x_453 = v_100 | v_39;
assign x_454 = v_99 | v_12;
assign x_455 = v_99 | v_20;
assign x_456 = v_98 | v_9;
assign x_457 = v_98 | ~v_20;
assign x_458 = v_24 | v_28 | v_29 | v_27 | v_26 | v_46 | v_45 | ~v_96 | ~v_95 | ~v_94 | ~v_93 | v_97;
assign x_459 = v_96 | v_54;
assign x_460 = v_96 | v_31;
assign x_461 = v_95 | ~v_54;
assign x_462 = v_95 | v_30;
assign x_463 = v_94 | v_10;
assign x_464 = v_94 | v_20;
assign x_465 = v_93 | v_8;
assign x_466 = v_93 | ~v_20;
assign x_467 = v_19 | v_18 | v_17 | v_16 | v_14 | v_42 | v_41 | ~v_91 | ~v_90 | ~v_89 | ~v_88 | v_92;
assign x_468 = v_91 | ~v_54;
assign x_469 = v_91 | v_21;
assign x_470 = v_90 | v_54;
assign x_471 = v_90 | v_22;
assign x_472 = v_89 | v_11;
assign x_473 = v_89 | v_20;
assign x_474 = v_88 | v_7;
assign x_475 = v_88 | ~v_20;
assign x_476 = ~v_86 | ~v_85 | ~v_84 | ~v_83 | ~v_82 | v_87;
assign x_477 = v_86 | v_8;
assign x_478 = v_86 | ~v_7;
assign x_479 = v_85 | v_9;
assign x_480 = v_85 | ~v_8;
assign x_481 = v_84 | v_11;
assign x_482 = v_84 | ~v_10;
assign x_483 = v_83 | v_10;
assign x_484 = v_83 | ~v_12;
assign x_485 = v_82 | ~v_71;
assign x_486 = v_82 | ~v_76;
assign x_487 = v_82 | ~v_81;
assign x_488 = v_32 | v_38 | v_37 | v_53 | v_61 | v_49 | v_64 | ~v_80 | ~v_79 | ~v_78 | ~v_77 | v_81;
assign x_489 = v_80 | v_59;
assign x_490 = v_80 | v_12;
assign x_491 = v_79 | ~v_59;
assign x_492 = v_79 | v_9;
assign x_493 = v_78 | v_59;
assign x_494 = v_78 | v_40;
assign x_495 = v_77 | ~v_59;
assign x_496 = v_77 | v_39;
assign x_497 = v_23 | v_28 | v_29 | v_52 | v_46 | v_63 | v_60 | ~v_75 | ~v_74 | ~v_73 | ~v_72 | v_76;
assign x_498 = v_75 | v_59;
assign x_499 = v_75 | v_10;
assign x_500 = v_74 | ~v_59;
assign x_501 = v_74 | v_8;
assign x_502 = v_73 | v_59;
assign x_503 = v_73 | v_31;
assign x_504 = v_72 | ~v_59;
assign x_505 = v_72 | v_30;
assign x_506 = v_13 | v_19 | v_18 | v_51 | v_62 | v_58 | v_42 | ~v_70 | ~v_69 | ~v_68 | ~v_67 | v_71;
assign x_507 = v_70 | v_59;
assign x_508 = v_70 | v_22;
assign x_509 = v_69 | ~v_59;
assign x_510 = v_69 | v_21;
assign x_511 = v_68 | v_59;
assign x_512 = v_68 | v_11;
assign x_513 = v_67 | ~v_59;
assign x_514 = v_67 | v_7;
assign x_515 = x_1 & x_2;
assign x_516 = x_3 & x_4;
assign x_517 = x_515 & x_516;
assign x_518 = x_5 & x_6;
assign x_519 = x_7 & x_8;
assign x_520 = x_518 & x_519;
assign x_521 = x_517 & x_520;
assign x_522 = x_9 & x_10;
assign x_523 = x_11 & x_12;
assign x_524 = x_522 & x_523;
assign x_525 = x_13 & x_14;
assign x_526 = x_15 & x_16;
assign x_527 = x_525 & x_526;
assign x_528 = x_524 & x_527;
assign x_529 = x_521 & x_528;
assign x_530 = x_17 & x_18;
assign x_531 = x_19 & x_20;
assign x_532 = x_530 & x_531;
assign x_533 = x_21 & x_22;
assign x_534 = x_23 & x_24;
assign x_535 = x_533 & x_534;
assign x_536 = x_532 & x_535;
assign x_537 = x_25 & x_26;
assign x_538 = x_27 & x_28;
assign x_539 = x_537 & x_538;
assign x_540 = x_29 & x_30;
assign x_541 = x_31 & x_32;
assign x_542 = x_540 & x_541;
assign x_543 = x_539 & x_542;
assign x_544 = x_536 & x_543;
assign x_545 = x_529 & x_544;
assign x_546 = x_33 & x_34;
assign x_547 = x_35 & x_36;
assign x_548 = x_546 & x_547;
assign x_549 = x_37 & x_38;
assign x_550 = x_39 & x_40;
assign x_551 = x_549 & x_550;
assign x_552 = x_548 & x_551;
assign x_553 = x_41 & x_42;
assign x_554 = x_43 & x_44;
assign x_555 = x_553 & x_554;
assign x_556 = x_45 & x_46;
assign x_557 = x_47 & x_48;
assign x_558 = x_556 & x_557;
assign x_559 = x_555 & x_558;
assign x_560 = x_552 & x_559;
assign x_561 = x_49 & x_50;
assign x_562 = x_51 & x_52;
assign x_563 = x_561 & x_562;
assign x_564 = x_53 & x_54;
assign x_565 = x_55 & x_56;
assign x_566 = x_564 & x_565;
assign x_567 = x_563 & x_566;
assign x_568 = x_57 & x_58;
assign x_569 = x_59 & x_60;
assign x_570 = x_568 & x_569;
assign x_571 = x_61 & x_62;
assign x_572 = x_63 & x_64;
assign x_573 = x_571 & x_572;
assign x_574 = x_570 & x_573;
assign x_575 = x_567 & x_574;
assign x_576 = x_560 & x_575;
assign x_577 = x_545 & x_576;
assign x_578 = x_65 & x_66;
assign x_579 = x_67 & x_68;
assign x_580 = x_578 & x_579;
assign x_581 = x_69 & x_70;
assign x_582 = x_71 & x_72;
assign x_583 = x_581 & x_582;
assign x_584 = x_580 & x_583;
assign x_585 = x_73 & x_74;
assign x_586 = x_75 & x_76;
assign x_587 = x_585 & x_586;
assign x_588 = x_77 & x_78;
assign x_589 = x_79 & x_80;
assign x_590 = x_588 & x_589;
assign x_591 = x_587 & x_590;
assign x_592 = x_584 & x_591;
assign x_593 = x_81 & x_82;
assign x_594 = x_83 & x_84;
assign x_595 = x_593 & x_594;
assign x_596 = x_85 & x_86;
assign x_597 = x_87 & x_88;
assign x_598 = x_596 & x_597;
assign x_599 = x_595 & x_598;
assign x_600 = x_89 & x_90;
assign x_601 = x_91 & x_92;
assign x_602 = x_600 & x_601;
assign x_603 = x_93 & x_94;
assign x_604 = x_95 & x_96;
assign x_605 = x_603 & x_604;
assign x_606 = x_602 & x_605;
assign x_607 = x_599 & x_606;
assign x_608 = x_592 & x_607;
assign x_609 = x_97 & x_98;
assign x_610 = x_99 & x_100;
assign x_611 = x_609 & x_610;
assign x_612 = x_101 & x_102;
assign x_613 = x_103 & x_104;
assign x_614 = x_612 & x_613;
assign x_615 = x_611 & x_614;
assign x_616 = x_105 & x_106;
assign x_617 = x_107 & x_108;
assign x_618 = x_616 & x_617;
assign x_619 = x_109 & x_110;
assign x_620 = x_111 & x_112;
assign x_621 = x_619 & x_620;
assign x_622 = x_618 & x_621;
assign x_623 = x_615 & x_622;
assign x_624 = x_113 & x_114;
assign x_625 = x_115 & x_116;
assign x_626 = x_624 & x_625;
assign x_627 = x_117 & x_118;
assign x_628 = x_119 & x_120;
assign x_629 = x_627 & x_628;
assign x_630 = x_626 & x_629;
assign x_631 = x_121 & x_122;
assign x_632 = x_123 & x_124;
assign x_633 = x_631 & x_632;
assign x_634 = x_125 & x_126;
assign x_635 = x_127 & x_128;
assign x_636 = x_634 & x_635;
assign x_637 = x_633 & x_636;
assign x_638 = x_630 & x_637;
assign x_639 = x_623 & x_638;
assign x_640 = x_608 & x_639;
assign x_641 = x_577 & x_640;
assign x_642 = x_129 & x_130;
assign x_643 = x_131 & x_132;
assign x_644 = x_642 & x_643;
assign x_645 = x_133 & x_134;
assign x_646 = x_135 & x_136;
assign x_647 = x_645 & x_646;
assign x_648 = x_644 & x_647;
assign x_649 = x_137 & x_138;
assign x_650 = x_139 & x_140;
assign x_651 = x_649 & x_650;
assign x_652 = x_141 & x_142;
assign x_653 = x_143 & x_144;
assign x_654 = x_652 & x_653;
assign x_655 = x_651 & x_654;
assign x_656 = x_648 & x_655;
assign x_657 = x_145 & x_146;
assign x_658 = x_147 & x_148;
assign x_659 = x_657 & x_658;
assign x_660 = x_149 & x_150;
assign x_661 = x_151 & x_152;
assign x_662 = x_660 & x_661;
assign x_663 = x_659 & x_662;
assign x_664 = x_153 & x_154;
assign x_665 = x_155 & x_156;
assign x_666 = x_664 & x_665;
assign x_667 = x_157 & x_158;
assign x_668 = x_159 & x_160;
assign x_669 = x_667 & x_668;
assign x_670 = x_666 & x_669;
assign x_671 = x_663 & x_670;
assign x_672 = x_656 & x_671;
assign x_673 = x_161 & x_162;
assign x_674 = x_163 & x_164;
assign x_675 = x_673 & x_674;
assign x_676 = x_165 & x_166;
assign x_677 = x_167 & x_168;
assign x_678 = x_676 & x_677;
assign x_679 = x_675 & x_678;
assign x_680 = x_169 & x_170;
assign x_681 = x_171 & x_172;
assign x_682 = x_680 & x_681;
assign x_683 = x_173 & x_174;
assign x_684 = x_175 & x_176;
assign x_685 = x_683 & x_684;
assign x_686 = x_682 & x_685;
assign x_687 = x_679 & x_686;
assign x_688 = x_177 & x_178;
assign x_689 = x_179 & x_180;
assign x_690 = x_688 & x_689;
assign x_691 = x_181 & x_182;
assign x_692 = x_183 & x_184;
assign x_693 = x_691 & x_692;
assign x_694 = x_690 & x_693;
assign x_695 = x_185 & x_186;
assign x_696 = x_187 & x_188;
assign x_697 = x_695 & x_696;
assign x_698 = x_189 & x_190;
assign x_699 = x_191 & x_192;
assign x_700 = x_698 & x_699;
assign x_701 = x_697 & x_700;
assign x_702 = x_694 & x_701;
assign x_703 = x_687 & x_702;
assign x_704 = x_672 & x_703;
assign x_705 = x_193 & x_194;
assign x_706 = x_195 & x_196;
assign x_707 = x_705 & x_706;
assign x_708 = x_197 & x_198;
assign x_709 = x_199 & x_200;
assign x_710 = x_708 & x_709;
assign x_711 = x_707 & x_710;
assign x_712 = x_201 & x_202;
assign x_713 = x_203 & x_204;
assign x_714 = x_712 & x_713;
assign x_715 = x_205 & x_206;
assign x_716 = x_207 & x_208;
assign x_717 = x_715 & x_716;
assign x_718 = x_714 & x_717;
assign x_719 = x_711 & x_718;
assign x_720 = x_209 & x_210;
assign x_721 = x_211 & x_212;
assign x_722 = x_720 & x_721;
assign x_723 = x_213 & x_214;
assign x_724 = x_215 & x_216;
assign x_725 = x_723 & x_724;
assign x_726 = x_722 & x_725;
assign x_727 = x_217 & x_218;
assign x_728 = x_219 & x_220;
assign x_729 = x_727 & x_728;
assign x_730 = x_221 & x_222;
assign x_731 = x_223 & x_224;
assign x_732 = x_730 & x_731;
assign x_733 = x_729 & x_732;
assign x_734 = x_726 & x_733;
assign x_735 = x_719 & x_734;
assign x_736 = x_225 & x_226;
assign x_737 = x_227 & x_228;
assign x_738 = x_736 & x_737;
assign x_739 = x_229 & x_230;
assign x_740 = x_231 & x_232;
assign x_741 = x_739 & x_740;
assign x_742 = x_738 & x_741;
assign x_743 = x_233 & x_234;
assign x_744 = x_235 & x_236;
assign x_745 = x_743 & x_744;
assign x_746 = x_237 & x_238;
assign x_747 = x_239 & x_240;
assign x_748 = x_746 & x_747;
assign x_749 = x_745 & x_748;
assign x_750 = x_742 & x_749;
assign x_751 = x_241 & x_242;
assign x_752 = x_243 & x_244;
assign x_753 = x_751 & x_752;
assign x_754 = x_245 & x_246;
assign x_755 = x_247 & x_248;
assign x_756 = x_754 & x_755;
assign x_757 = x_753 & x_756;
assign x_758 = x_249 & x_250;
assign x_759 = x_251 & x_252;
assign x_760 = x_758 & x_759;
assign x_761 = x_253 & x_254;
assign x_762 = x_256 & x_257;
assign x_763 = x_255 & x_762;
assign x_764 = x_761 & x_763;
assign x_765 = x_760 & x_764;
assign x_766 = x_757 & x_765;
assign x_767 = x_750 & x_766;
assign x_768 = x_735 & x_767;
assign x_769 = x_704 & x_768;
assign x_770 = x_641 & x_769;
assign x_771 = x_258 & x_259;
assign x_772 = x_260 & x_261;
assign x_773 = x_771 & x_772;
assign x_774 = x_262 & x_263;
assign x_775 = x_264 & x_265;
assign x_776 = x_774 & x_775;
assign x_777 = x_773 & x_776;
assign x_778 = x_266 & x_267;
assign x_779 = x_268 & x_269;
assign x_780 = x_778 & x_779;
assign x_781 = x_270 & x_271;
assign x_782 = x_272 & x_273;
assign x_783 = x_781 & x_782;
assign x_784 = x_780 & x_783;
assign x_785 = x_777 & x_784;
assign x_786 = x_274 & x_275;
assign x_787 = x_276 & x_277;
assign x_788 = x_786 & x_787;
assign x_789 = x_278 & x_279;
assign x_790 = x_280 & x_281;
assign x_791 = x_789 & x_790;
assign x_792 = x_788 & x_791;
assign x_793 = x_282 & x_283;
assign x_794 = x_284 & x_285;
assign x_795 = x_793 & x_794;
assign x_796 = x_286 & x_287;
assign x_797 = x_288 & x_289;
assign x_798 = x_796 & x_797;
assign x_799 = x_795 & x_798;
assign x_800 = x_792 & x_799;
assign x_801 = x_785 & x_800;
assign x_802 = x_290 & x_291;
assign x_803 = x_292 & x_293;
assign x_804 = x_802 & x_803;
assign x_805 = x_294 & x_295;
assign x_806 = x_296 & x_297;
assign x_807 = x_805 & x_806;
assign x_808 = x_804 & x_807;
assign x_809 = x_298 & x_299;
assign x_810 = x_300 & x_301;
assign x_811 = x_809 & x_810;
assign x_812 = x_302 & x_303;
assign x_813 = x_304 & x_305;
assign x_814 = x_812 & x_813;
assign x_815 = x_811 & x_814;
assign x_816 = x_808 & x_815;
assign x_817 = x_306 & x_307;
assign x_818 = x_308 & x_309;
assign x_819 = x_817 & x_818;
assign x_820 = x_310 & x_311;
assign x_821 = x_312 & x_313;
assign x_822 = x_820 & x_821;
assign x_823 = x_819 & x_822;
assign x_824 = x_314 & x_315;
assign x_825 = x_316 & x_317;
assign x_826 = x_824 & x_825;
assign x_827 = x_318 & x_319;
assign x_828 = x_320 & x_321;
assign x_829 = x_827 & x_828;
assign x_830 = x_826 & x_829;
assign x_831 = x_823 & x_830;
assign x_832 = x_816 & x_831;
assign x_833 = x_801 & x_832;
assign x_834 = x_322 & x_323;
assign x_835 = x_324 & x_325;
assign x_836 = x_834 & x_835;
assign x_837 = x_326 & x_327;
assign x_838 = x_328 & x_329;
assign x_839 = x_837 & x_838;
assign x_840 = x_836 & x_839;
assign x_841 = x_330 & x_331;
assign x_842 = x_332 & x_333;
assign x_843 = x_841 & x_842;
assign x_844 = x_334 & x_335;
assign x_845 = x_336 & x_337;
assign x_846 = x_844 & x_845;
assign x_847 = x_843 & x_846;
assign x_848 = x_840 & x_847;
assign x_849 = x_338 & x_339;
assign x_850 = x_340 & x_341;
assign x_851 = x_849 & x_850;
assign x_852 = x_342 & x_343;
assign x_853 = x_344 & x_345;
assign x_854 = x_852 & x_853;
assign x_855 = x_851 & x_854;
assign x_856 = x_346 & x_347;
assign x_857 = x_348 & x_349;
assign x_858 = x_856 & x_857;
assign x_859 = x_350 & x_351;
assign x_860 = x_352 & x_353;
assign x_861 = x_859 & x_860;
assign x_862 = x_858 & x_861;
assign x_863 = x_855 & x_862;
assign x_864 = x_848 & x_863;
assign x_865 = x_354 & x_355;
assign x_866 = x_356 & x_357;
assign x_867 = x_865 & x_866;
assign x_868 = x_358 & x_359;
assign x_869 = x_360 & x_361;
assign x_870 = x_868 & x_869;
assign x_871 = x_867 & x_870;
assign x_872 = x_362 & x_363;
assign x_873 = x_364 & x_365;
assign x_874 = x_872 & x_873;
assign x_875 = x_366 & x_367;
assign x_876 = x_368 & x_369;
assign x_877 = x_875 & x_876;
assign x_878 = x_874 & x_877;
assign x_879 = x_871 & x_878;
assign x_880 = x_370 & x_371;
assign x_881 = x_372 & x_373;
assign x_882 = x_880 & x_881;
assign x_883 = x_374 & x_375;
assign x_884 = x_376 & x_377;
assign x_885 = x_883 & x_884;
assign x_886 = x_882 & x_885;
assign x_887 = x_378 & x_379;
assign x_888 = x_380 & x_381;
assign x_889 = x_887 & x_888;
assign x_890 = x_382 & x_383;
assign x_891 = x_384 & x_385;
assign x_892 = x_890 & x_891;
assign x_893 = x_889 & x_892;
assign x_894 = x_886 & x_893;
assign x_895 = x_879 & x_894;
assign x_896 = x_864 & x_895;
assign x_897 = x_833 & x_896;
assign x_898 = x_386 & x_387;
assign x_899 = x_388 & x_389;
assign x_900 = x_898 & x_899;
assign x_901 = x_390 & x_391;
assign x_902 = x_392 & x_393;
assign x_903 = x_901 & x_902;
assign x_904 = x_900 & x_903;
assign x_905 = x_394 & x_395;
assign x_906 = x_396 & x_397;
assign x_907 = x_905 & x_906;
assign x_908 = x_398 & x_399;
assign x_909 = x_400 & x_401;
assign x_910 = x_908 & x_909;
assign x_911 = x_907 & x_910;
assign x_912 = x_904 & x_911;
assign x_913 = x_402 & x_403;
assign x_914 = x_404 & x_405;
assign x_915 = x_913 & x_914;
assign x_916 = x_406 & x_407;
assign x_917 = x_408 & x_409;
assign x_918 = x_916 & x_917;
assign x_919 = x_915 & x_918;
assign x_920 = x_410 & x_411;
assign x_921 = x_412 & x_413;
assign x_922 = x_920 & x_921;
assign x_923 = x_414 & x_415;
assign x_924 = x_416 & x_417;
assign x_925 = x_923 & x_924;
assign x_926 = x_922 & x_925;
assign x_927 = x_919 & x_926;
assign x_928 = x_912 & x_927;
assign x_929 = x_418 & x_419;
assign x_930 = x_420 & x_421;
assign x_931 = x_929 & x_930;
assign x_932 = x_422 & x_423;
assign x_933 = x_424 & x_425;
assign x_934 = x_932 & x_933;
assign x_935 = x_931 & x_934;
assign x_936 = x_426 & x_427;
assign x_937 = x_428 & x_429;
assign x_938 = x_936 & x_937;
assign x_939 = x_430 & x_431;
assign x_940 = x_432 & x_433;
assign x_941 = x_939 & x_940;
assign x_942 = x_938 & x_941;
assign x_943 = x_935 & x_942;
assign x_944 = x_434 & x_435;
assign x_945 = x_436 & x_437;
assign x_946 = x_944 & x_945;
assign x_947 = x_438 & x_439;
assign x_948 = x_440 & x_441;
assign x_949 = x_947 & x_948;
assign x_950 = x_946 & x_949;
assign x_951 = x_442 & x_443;
assign x_952 = x_444 & x_445;
assign x_953 = x_951 & x_952;
assign x_954 = x_446 & x_447;
assign x_955 = x_448 & x_449;
assign x_956 = x_954 & x_955;
assign x_957 = x_953 & x_956;
assign x_958 = x_950 & x_957;
assign x_959 = x_943 & x_958;
assign x_960 = x_928 & x_959;
assign x_961 = x_450 & x_451;
assign x_962 = x_452 & x_453;
assign x_963 = x_961 & x_962;
assign x_964 = x_454 & x_455;
assign x_965 = x_456 & x_457;
assign x_966 = x_964 & x_965;
assign x_967 = x_963 & x_966;
assign x_968 = x_458 & x_459;
assign x_969 = x_460 & x_461;
assign x_970 = x_968 & x_969;
assign x_971 = x_462 & x_463;
assign x_972 = x_464 & x_465;
assign x_973 = x_971 & x_972;
assign x_974 = x_970 & x_973;
assign x_975 = x_967 & x_974;
assign x_976 = x_466 & x_467;
assign x_977 = x_468 & x_469;
assign x_978 = x_976 & x_977;
assign x_979 = x_470 & x_471;
assign x_980 = x_472 & x_473;
assign x_981 = x_979 & x_980;
assign x_982 = x_978 & x_981;
assign x_983 = x_474 & x_475;
assign x_984 = x_476 & x_477;
assign x_985 = x_983 & x_984;
assign x_986 = x_478 & x_479;
assign x_987 = x_480 & x_481;
assign x_988 = x_986 & x_987;
assign x_989 = x_985 & x_988;
assign x_990 = x_982 & x_989;
assign x_991 = x_975 & x_990;
assign x_992 = x_482 & x_483;
assign x_993 = x_484 & x_485;
assign x_994 = x_992 & x_993;
assign x_995 = x_486 & x_487;
assign x_996 = x_488 & x_489;
assign x_997 = x_995 & x_996;
assign x_998 = x_994 & x_997;
assign x_999 = x_490 & x_491;
assign x_1000 = x_492 & x_493;
assign x_1001 = x_999 & x_1000;
assign x_1002 = x_494 & x_495;
assign x_1003 = x_496 & x_497;
assign x_1004 = x_1002 & x_1003;
assign x_1005 = x_1001 & x_1004;
assign x_1006 = x_998 & x_1005;
assign x_1007 = x_498 & x_499;
assign x_1008 = x_500 & x_501;
assign x_1009 = x_1007 & x_1008;
assign x_1010 = x_502 & x_503;
assign x_1011 = x_504 & x_505;
assign x_1012 = x_1010 & x_1011;
assign x_1013 = x_1009 & x_1012;
assign x_1014 = x_506 & x_507;
assign x_1015 = x_508 & x_509;
assign x_1016 = x_1014 & x_1015;
assign x_1017 = x_510 & x_511;
assign x_1018 = x_513 & x_514;
assign x_1019 = x_512 & x_1018;
assign x_1020 = x_1017 & x_1019;
assign x_1021 = x_1016 & x_1020;
assign x_1022 = x_1013 & x_1021;
assign x_1023 = x_1006 & x_1022;
assign x_1024 = x_991 & x_1023;
assign x_1025 = x_960 & x_1024;
assign x_1026 = x_897 & x_1025;
assign x_1027 = x_770 & x_1026;
assign o_1 = x_1027;
endmodule
